module basic_2500_25000_3000_100_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_1725,In_1472);
xnor U1 (N_1,In_2087,In_835);
nand U2 (N_2,In_354,In_2363);
xor U3 (N_3,In_2413,In_261);
nor U4 (N_4,In_2390,In_1397);
nand U5 (N_5,In_125,In_484);
nor U6 (N_6,In_398,In_2038);
xor U7 (N_7,In_37,In_1242);
xor U8 (N_8,In_2311,In_2392);
xor U9 (N_9,In_1356,In_478);
or U10 (N_10,In_2252,In_625);
nor U11 (N_11,In_608,In_492);
xnor U12 (N_12,In_2318,In_2456);
and U13 (N_13,In_485,In_95);
xnor U14 (N_14,In_2253,In_327);
or U15 (N_15,In_1502,In_833);
nor U16 (N_16,In_2387,In_2463);
nor U17 (N_17,In_100,In_1048);
and U18 (N_18,In_1793,In_1375);
or U19 (N_19,In_1171,In_70);
nor U20 (N_20,In_1929,In_1453);
and U21 (N_21,In_2012,In_1214);
nand U22 (N_22,In_449,In_1314);
nor U23 (N_23,In_181,In_2435);
nand U24 (N_24,In_1713,In_2420);
xor U25 (N_25,In_1054,In_29);
and U26 (N_26,In_1534,In_2427);
xnor U27 (N_27,In_2141,In_2182);
or U28 (N_28,In_961,In_1252);
or U29 (N_29,In_1404,In_2186);
nor U30 (N_30,In_992,In_62);
nor U31 (N_31,In_204,In_1238);
or U32 (N_32,In_1794,In_513);
xor U33 (N_33,In_136,In_291);
xor U34 (N_34,In_2351,In_1703);
or U35 (N_35,In_1352,In_378);
and U36 (N_36,In_236,In_1056);
nand U37 (N_37,In_1531,In_1824);
xor U38 (N_38,In_1983,In_2349);
and U39 (N_39,In_940,In_2411);
xnor U40 (N_40,In_477,In_375);
and U41 (N_41,In_1648,In_493);
or U42 (N_42,In_1973,In_616);
xor U43 (N_43,In_182,In_345);
and U44 (N_44,In_247,In_1445);
nand U45 (N_45,In_69,In_2088);
and U46 (N_46,In_800,In_1051);
nand U47 (N_47,In_138,In_2019);
or U48 (N_48,In_83,In_166);
nor U49 (N_49,In_1190,In_1550);
or U50 (N_50,In_1295,In_429);
nor U51 (N_51,In_1627,In_682);
nand U52 (N_52,In_830,In_1717);
nand U53 (N_53,In_2256,In_698);
and U54 (N_54,In_299,In_917);
xor U55 (N_55,In_1920,In_688);
nor U56 (N_56,In_338,In_788);
nor U57 (N_57,In_984,In_1165);
or U58 (N_58,In_67,In_1264);
or U59 (N_59,In_1077,In_920);
xor U60 (N_60,In_2477,In_42);
and U61 (N_61,In_1278,In_171);
nand U62 (N_62,In_2377,In_1290);
xor U63 (N_63,In_2434,In_733);
and U64 (N_64,In_503,In_1387);
nor U65 (N_65,In_1057,In_2319);
xnor U66 (N_66,In_1718,In_832);
nand U67 (N_67,In_599,In_1912);
xnor U68 (N_68,In_1811,In_740);
nor U69 (N_69,In_2379,In_1766);
and U70 (N_70,In_849,In_1667);
and U71 (N_71,In_2028,In_875);
nand U72 (N_72,In_1932,In_2224);
xnor U73 (N_73,In_1828,In_1331);
and U74 (N_74,In_164,In_1910);
nor U75 (N_75,In_490,In_16);
and U76 (N_76,In_922,In_1598);
or U77 (N_77,In_1343,In_930);
or U78 (N_78,In_1741,In_2286);
and U79 (N_79,In_2417,In_2400);
nand U80 (N_80,In_1711,In_1976);
nand U81 (N_81,In_679,In_1805);
and U82 (N_82,In_1095,In_1186);
or U83 (N_83,In_1353,In_284);
nand U84 (N_84,In_315,In_2350);
nand U85 (N_85,In_75,In_1599);
and U86 (N_86,In_1306,In_2086);
nand U87 (N_87,In_1587,In_318);
xnor U88 (N_88,In_1956,In_604);
and U89 (N_89,In_1755,In_794);
or U90 (N_90,In_280,In_115);
nand U91 (N_91,In_656,In_854);
or U92 (N_92,In_749,In_1770);
nor U93 (N_93,In_1359,In_1562);
nand U94 (N_94,In_2037,In_2083);
xor U95 (N_95,In_887,In_691);
nand U96 (N_96,In_512,In_2187);
nand U97 (N_97,In_1651,In_133);
or U98 (N_98,In_2484,In_1427);
xor U99 (N_99,In_1887,In_147);
xor U100 (N_100,In_1132,In_663);
nand U101 (N_101,In_489,In_560);
or U102 (N_102,In_1998,In_1560);
xnor U103 (N_103,In_2073,In_947);
and U104 (N_104,In_1913,In_841);
nand U105 (N_105,In_1880,In_798);
nor U106 (N_106,In_1151,In_633);
nand U107 (N_107,In_266,In_2448);
or U108 (N_108,In_1437,In_2061);
and U109 (N_109,In_593,In_1742);
and U110 (N_110,In_1287,In_1954);
xor U111 (N_111,In_2218,In_1854);
xnor U112 (N_112,In_1644,In_729);
nor U113 (N_113,In_1737,In_127);
xnor U114 (N_114,In_1544,In_2231);
or U115 (N_115,In_1324,In_389);
xnor U116 (N_116,In_1832,In_205);
or U117 (N_117,In_1175,In_2174);
nor U118 (N_118,In_714,In_1941);
nand U119 (N_119,In_1873,In_846);
nor U120 (N_120,In_996,In_797);
xor U121 (N_121,In_1201,In_844);
and U122 (N_122,In_488,In_1779);
and U123 (N_123,In_46,In_1342);
xnor U124 (N_124,In_767,In_2245);
nand U125 (N_125,In_1628,In_2120);
or U126 (N_126,In_114,In_458);
nor U127 (N_127,In_1181,In_1421);
or U128 (N_128,In_758,In_4);
and U129 (N_129,In_1698,In_9);
nor U130 (N_130,In_1303,In_1650);
and U131 (N_131,In_2100,In_592);
nor U132 (N_132,In_594,In_1645);
xnor U133 (N_133,In_2402,In_1149);
nor U134 (N_134,In_1184,In_1402);
or U135 (N_135,In_1921,In_421);
and U136 (N_136,In_1567,In_1552);
nand U137 (N_137,In_240,In_1809);
xor U138 (N_138,In_1559,In_1726);
nor U139 (N_139,In_1035,In_859);
nor U140 (N_140,In_1507,In_1194);
nand U141 (N_141,In_1441,In_827);
or U142 (N_142,In_239,In_660);
and U143 (N_143,In_649,In_1394);
xnor U144 (N_144,In_1274,In_600);
and U145 (N_145,In_200,In_1169);
xnor U146 (N_146,In_1189,In_562);
or U147 (N_147,In_793,In_2122);
xnor U148 (N_148,In_207,In_1623);
xnor U149 (N_149,In_2323,In_2391);
xor U150 (N_150,In_172,In_2489);
or U151 (N_151,In_402,In_1112);
or U152 (N_152,In_233,In_2238);
and U153 (N_153,In_2166,In_523);
xor U154 (N_154,In_1503,In_1275);
nand U155 (N_155,In_476,In_215);
nor U156 (N_156,In_748,In_2431);
and U157 (N_157,In_313,In_908);
nor U158 (N_158,In_547,In_1928);
and U159 (N_159,In_1422,In_1757);
xor U160 (N_160,In_2084,In_2326);
and U161 (N_161,In_823,In_2382);
and U162 (N_162,In_1866,In_1480);
or U163 (N_163,In_1838,In_71);
and U164 (N_164,In_2446,In_2273);
xnor U165 (N_165,In_861,In_2276);
xor U166 (N_166,In_2135,In_435);
and U167 (N_167,In_694,In_231);
nor U168 (N_168,In_2490,In_1449);
nor U169 (N_169,In_1075,In_1923);
xor U170 (N_170,In_807,In_550);
or U171 (N_171,In_1037,In_54);
xor U172 (N_172,In_736,In_659);
or U173 (N_173,In_122,In_287);
xnor U174 (N_174,In_993,In_746);
and U175 (N_175,In_1597,In_331);
and U176 (N_176,In_583,In_410);
or U177 (N_177,In_2486,In_955);
nand U178 (N_178,In_2176,In_966);
nand U179 (N_179,In_2030,In_451);
nand U180 (N_180,In_1145,In_1443);
or U181 (N_181,In_2219,In_1886);
or U182 (N_182,In_787,In_2430);
xnor U183 (N_183,In_774,In_637);
or U184 (N_184,In_310,In_2107);
and U185 (N_185,In_1801,In_2254);
or U186 (N_186,In_2004,In_622);
nand U187 (N_187,In_198,In_1549);
nand U188 (N_188,In_2188,In_1355);
nor U189 (N_189,In_2171,In_1438);
or U190 (N_190,In_1256,In_301);
and U191 (N_191,In_1787,In_1951);
nand U192 (N_192,In_2094,In_415);
or U193 (N_193,In_704,In_1364);
or U194 (N_194,In_194,In_584);
nor U195 (N_195,In_1494,In_1752);
nand U196 (N_196,In_1827,In_1140);
nor U197 (N_197,In_1647,In_53);
nand U198 (N_198,In_498,In_1895);
or U199 (N_199,In_2184,In_350);
or U200 (N_200,In_712,In_2447);
nand U201 (N_201,In_469,In_474);
or U202 (N_202,In_564,In_1868);
xor U203 (N_203,In_1918,In_641);
nand U204 (N_204,In_2185,In_99);
nor U205 (N_205,In_819,In_408);
and U206 (N_206,In_103,In_143);
or U207 (N_207,In_915,In_2263);
nand U208 (N_208,In_921,In_1191);
xnor U209 (N_209,In_817,In_1780);
nand U210 (N_210,In_586,In_699);
or U211 (N_211,In_668,In_1875);
xnor U212 (N_212,In_2112,In_874);
xnor U213 (N_213,In_153,In_1116);
nand U214 (N_214,In_860,In_615);
nand U215 (N_215,In_268,In_452);
xor U216 (N_216,In_2381,In_59);
and U217 (N_217,In_686,In_1401);
nand U218 (N_218,In_282,In_1831);
or U219 (N_219,In_1059,In_2370);
and U220 (N_220,In_1909,In_1043);
and U221 (N_221,In_1685,In_1509);
or U222 (N_222,In_1596,In_1601);
and U223 (N_223,In_2396,In_804);
xnor U224 (N_224,In_72,In_442);
and U225 (N_225,In_169,In_1150);
or U226 (N_226,In_2475,In_697);
and U227 (N_227,In_2007,In_362);
and U228 (N_228,In_145,In_579);
nand U229 (N_229,In_480,In_837);
and U230 (N_230,In_782,In_971);
xor U231 (N_231,In_270,In_1984);
xnor U232 (N_232,In_339,In_1336);
or U233 (N_233,In_1411,In_188);
and U234 (N_234,In_130,In_1781);
xnor U235 (N_235,In_2343,In_277);
and U236 (N_236,In_1891,In_1620);
nor U237 (N_237,In_385,In_1152);
xor U238 (N_238,In_1136,In_2146);
nor U239 (N_239,In_1608,In_1296);
xnor U240 (N_240,In_1800,In_356);
or U241 (N_241,In_1329,In_872);
or U242 (N_242,In_1989,In_2029);
or U243 (N_243,In_471,In_2241);
xnor U244 (N_244,In_1046,In_332);
or U245 (N_245,In_2167,In_2214);
or U246 (N_246,In_2246,In_776);
nor U247 (N_247,In_1847,In_86);
nor U248 (N_248,In_1864,In_1313);
xor U249 (N_249,In_1374,In_2156);
and U250 (N_250,In_92,In_806);
nand U251 (N_251,In_413,In_2488);
nand U252 (N_252,In_2358,In_991);
nand U253 (N_253,In_700,In_1055);
nand U254 (N_254,In_1734,N_45);
xnor U255 (N_255,In_927,In_1486);
or U256 (N_256,In_191,In_1396);
nor U257 (N_257,In_2419,In_945);
nand U258 (N_258,In_718,In_1814);
nor U259 (N_259,In_1273,In_1241);
nor U260 (N_260,In_2281,In_2287);
and U261 (N_261,In_348,N_173);
nor U262 (N_262,In_960,In_454);
nand U263 (N_263,In_1257,In_1916);
or U264 (N_264,In_689,In_1460);
or U265 (N_265,In_2069,In_2236);
or U266 (N_266,In_1553,In_1829);
and U267 (N_267,In_1395,In_1100);
xor U268 (N_268,N_120,In_420);
and U269 (N_269,In_717,In_811);
nand U270 (N_270,In_2126,In_2162);
or U271 (N_271,In_245,In_1749);
nand U272 (N_272,N_123,In_981);
nor U273 (N_273,N_124,In_329);
or U274 (N_274,In_211,In_627);
and U275 (N_275,N_203,In_40);
nor U276 (N_276,In_2406,In_724);
or U277 (N_277,N_59,In_680);
or U278 (N_278,In_1641,In_610);
and U279 (N_279,In_1450,In_1782);
nand U280 (N_280,In_1690,In_1898);
and U281 (N_281,In_1533,In_1930);
and U282 (N_282,In_1985,In_1247);
nor U283 (N_283,N_243,In_2106);
nand U284 (N_284,In_1993,In_2438);
nand U285 (N_285,N_74,In_274);
xor U286 (N_286,In_1992,In_1939);
xnor U287 (N_287,In_324,In_664);
nand U288 (N_288,In_1610,In_2117);
nor U289 (N_289,In_1488,In_1052);
or U290 (N_290,In_225,In_1423);
or U291 (N_291,In_713,In_1936);
xnor U292 (N_292,In_1272,N_189);
or U293 (N_293,In_1268,In_1218);
and U294 (N_294,In_1677,N_241);
or U295 (N_295,In_1915,In_2157);
and U296 (N_296,In_383,In_1351);
nand U297 (N_297,In_973,In_901);
nor U298 (N_298,In_2242,In_696);
xnor U299 (N_299,In_2204,In_1777);
or U300 (N_300,In_2476,In_507);
or U301 (N_301,In_453,In_431);
or U302 (N_302,In_246,In_1361);
or U303 (N_303,In_1840,In_1520);
nor U304 (N_304,In_1662,In_1636);
nor U305 (N_305,In_588,In_1068);
nand U306 (N_306,In_1638,In_2074);
xnor U307 (N_307,In_19,N_145);
nand U308 (N_308,In_2,In_109);
or U309 (N_309,In_1029,In_2398);
or U310 (N_310,In_1468,In_1282);
xnor U311 (N_311,In_2054,In_2329);
nand U312 (N_312,In_692,In_256);
and U313 (N_313,In_1861,In_1119);
and U314 (N_314,In_1018,In_1117);
and U315 (N_315,In_1906,N_150);
nor U316 (N_316,N_153,In_791);
nor U317 (N_317,In_886,In_2334);
nand U318 (N_318,In_1061,In_1721);
nand U319 (N_319,In_578,In_851);
and U320 (N_320,In_1090,In_2123);
nand U321 (N_321,In_2403,In_1366);
nand U322 (N_322,In_710,In_352);
and U323 (N_323,In_909,In_496);
nand U324 (N_324,In_755,In_2441);
xor U325 (N_325,In_1889,In_896);
nand U326 (N_326,In_906,In_1894);
nand U327 (N_327,In_73,In_384);
and U328 (N_328,In_538,In_2330);
nor U329 (N_329,In_1826,In_1491);
nor U330 (N_330,In_1373,In_1530);
and U331 (N_331,In_1626,In_1978);
or U332 (N_332,In_235,In_1340);
xnor U333 (N_333,In_987,In_305);
xor U334 (N_334,In_866,In_2255);
nand U335 (N_335,In_2362,In_654);
xnor U336 (N_336,In_263,In_1473);
or U337 (N_337,In_2017,In_2493);
or U338 (N_338,In_141,N_7);
nand U339 (N_339,N_55,In_939);
nand U340 (N_340,N_249,In_977);
xor U341 (N_341,In_1196,In_693);
nor U342 (N_342,In_568,In_1934);
nand U343 (N_343,In_1842,In_2309);
or U344 (N_344,In_303,N_16);
or U345 (N_345,In_2453,In_1876);
nand U346 (N_346,In_2366,In_1542);
nor U347 (N_347,In_2217,In_1413);
or U348 (N_348,In_366,In_1591);
nor U349 (N_349,In_89,In_2132);
nand U350 (N_350,In_187,In_1694);
or U351 (N_351,In_1695,N_90);
xor U352 (N_352,In_742,In_1419);
nor U353 (N_353,In_1511,In_559);
nor U354 (N_354,In_1806,In_1341);
or U355 (N_355,In_1323,In_910);
nor U356 (N_356,In_30,In_31);
or U357 (N_357,In_370,N_180);
nand U358 (N_358,In_737,N_198);
and U359 (N_359,In_1935,N_148);
nand U360 (N_360,In_2058,In_49);
nand U361 (N_361,In_64,In_1231);
and U362 (N_362,In_1668,In_197);
and U363 (N_363,In_555,In_862);
nor U364 (N_364,In_2344,In_646);
nor U365 (N_365,In_630,In_2429);
nand U366 (N_366,In_1762,In_2144);
or U367 (N_367,In_1783,In_1253);
nand U368 (N_368,In_1848,In_1281);
xor U369 (N_369,In_706,In_1316);
and U370 (N_370,In_1094,In_1461);
or U371 (N_371,In_1229,In_213);
xnor U372 (N_372,N_25,In_897);
nand U373 (N_373,In_1672,In_1674);
nor U374 (N_374,In_543,In_20);
nor U375 (N_375,In_893,In_1269);
or U376 (N_376,In_1379,In_2280);
or U377 (N_377,In_1344,In_294);
nand U378 (N_378,In_1129,In_825);
or U379 (N_379,In_2203,In_2057);
xnor U380 (N_380,In_1967,In_222);
nor U381 (N_381,In_361,In_1250);
nand U382 (N_382,In_2405,In_1870);
or U383 (N_383,In_1408,In_751);
xnor U384 (N_384,In_934,N_33);
nor U385 (N_385,In_903,In_2364);
nand U386 (N_386,In_482,In_26);
xnor U387 (N_387,In_1643,N_34);
xnor U388 (N_388,In_1288,N_222);
nand U389 (N_389,In_1631,In_417);
nor U390 (N_390,In_1266,In_1592);
nor U391 (N_391,In_1528,In_781);
or U392 (N_392,N_113,In_192);
or U393 (N_393,In_1154,In_1877);
xor U394 (N_394,In_1174,N_218);
nand U395 (N_395,In_177,In_1362);
or U396 (N_396,In_533,In_669);
and U397 (N_397,N_245,In_443);
nand U398 (N_398,In_1161,In_2418);
and U399 (N_399,In_1334,In_1772);
nor U400 (N_400,In_1882,In_790);
nor U401 (N_401,In_161,In_2320);
and U402 (N_402,In_473,In_2006);
or U403 (N_403,In_2265,In_1399);
xnor U404 (N_404,In_146,In_390);
or U405 (N_405,In_1455,In_1004);
nand U406 (N_406,In_1086,In_2016);
nand U407 (N_407,N_129,In_936);
nor U408 (N_408,In_320,In_2258);
nor U409 (N_409,In_2491,In_1433);
nor U410 (N_410,In_45,In_1869);
and U411 (N_411,In_1944,In_502);
or U412 (N_412,In_1153,In_2227);
or U413 (N_413,In_944,In_2481);
or U414 (N_414,In_1859,In_1697);
nand U415 (N_415,In_1237,In_2365);
nor U416 (N_416,In_184,In_926);
xor U417 (N_417,In_253,In_1042);
xor U418 (N_418,N_65,In_2394);
xnor U419 (N_419,In_553,N_61);
nand U420 (N_420,In_796,In_1865);
and U421 (N_421,In_620,In_1529);
nor U422 (N_422,N_149,In_2439);
xnor U423 (N_423,In_2230,N_171);
nand U424 (N_424,In_35,In_2210);
or U425 (N_425,In_1118,N_117);
nor U426 (N_426,In_997,In_708);
nor U427 (N_427,In_1255,In_2416);
or U428 (N_428,In_1028,In_1157);
or U429 (N_429,In_1791,In_1710);
nor U430 (N_430,In_1147,In_720);
nor U431 (N_431,In_1065,In_386);
or U432 (N_432,In_1409,In_2047);
and U433 (N_433,In_60,In_2115);
nand U434 (N_434,In_2353,In_1872);
nor U435 (N_435,In_238,In_1945);
or U436 (N_436,In_1837,In_1008);
or U437 (N_437,In_1588,N_71);
nor U438 (N_438,In_1893,In_2040);
nand U439 (N_439,In_1195,N_146);
xnor U440 (N_440,In_108,In_2015);
nand U441 (N_441,In_914,In_1492);
nand U442 (N_442,In_2189,In_1280);
xor U443 (N_443,N_98,In_74);
or U444 (N_444,In_175,In_1927);
or U445 (N_445,In_363,N_48);
or U446 (N_446,In_119,In_970);
nor U447 (N_447,In_1962,In_1758);
nor U448 (N_448,In_818,In_942);
xnor U449 (N_449,In_1270,In_1576);
and U450 (N_450,In_1309,In_2172);
or U451 (N_451,In_152,In_2498);
nor U452 (N_452,In_1763,N_137);
and U453 (N_453,N_230,In_2000);
and U454 (N_454,In_179,N_209);
or U455 (N_455,In_2164,In_497);
xnor U456 (N_456,In_567,In_1234);
nand U457 (N_457,In_2397,In_769);
and U458 (N_458,In_400,In_2150);
xnor U459 (N_459,N_62,In_1133);
xnor U460 (N_460,In_190,In_1416);
and U461 (N_461,In_836,In_2033);
or U462 (N_462,In_2426,In_761);
nor U463 (N_463,In_2148,In_387);
or U464 (N_464,In_393,In_2243);
nor U465 (N_465,In_333,In_657);
nor U466 (N_466,In_965,In_1570);
and U467 (N_467,In_80,In_2262);
nand U468 (N_468,In_1011,In_2361);
nand U469 (N_469,In_217,N_96);
and U470 (N_470,In_1302,In_1245);
xor U471 (N_471,In_1629,In_1818);
nand U472 (N_472,In_173,In_1510);
and U473 (N_473,In_2485,In_544);
xnor U474 (N_474,In_2314,In_1977);
nor U475 (N_475,In_13,In_2315);
xor U476 (N_476,In_1982,In_530);
xor U477 (N_477,In_2295,In_570);
nand U478 (N_478,In_838,In_1289);
nand U479 (N_479,In_809,In_1271);
nand U480 (N_480,In_2010,In_1774);
nand U481 (N_481,In_557,In_2371);
xor U482 (N_482,In_1386,N_75);
and U483 (N_483,In_340,In_414);
and U484 (N_484,In_468,N_161);
and U485 (N_485,In_956,In_1217);
nor U486 (N_486,In_1834,In_199);
and U487 (N_487,In_1384,In_2298);
nor U488 (N_488,In_515,In_1463);
or U489 (N_489,In_1032,In_681);
and U490 (N_490,In_349,N_225);
xor U491 (N_491,In_756,In_63);
or U492 (N_492,In_1543,In_980);
xor U493 (N_493,In_2163,In_1160);
nor U494 (N_494,In_7,In_1084);
or U495 (N_495,In_1988,In_1205);
or U496 (N_496,In_2465,In_2445);
nor U497 (N_497,In_719,In_1412);
xor U498 (N_498,In_1911,In_1566);
or U499 (N_499,In_810,In_401);
nand U500 (N_500,N_331,N_217);
and U501 (N_501,In_165,In_309);
nand U502 (N_502,N_464,N_69);
or U503 (N_503,In_2451,N_40);
and U504 (N_504,In_78,N_359);
nor U505 (N_505,In_229,In_1370);
and U506 (N_506,N_379,In_1292);
nand U507 (N_507,In_1203,In_1568);
nand U508 (N_508,In_526,N_99);
or U509 (N_509,In_1501,N_57);
nand U510 (N_510,In_609,In_163);
nor U511 (N_511,N_393,In_2303);
or U512 (N_512,N_58,In_463);
and U513 (N_513,In_1613,In_396);
nor U514 (N_514,In_2399,In_2283);
nand U515 (N_515,N_274,In_953);
or U516 (N_516,In_1328,N_485);
and U517 (N_517,In_1579,In_962);
or U518 (N_518,N_477,In_2108);
and U519 (N_519,N_499,N_315);
nor U520 (N_520,N_496,In_1446);
or U521 (N_521,In_982,In_1310);
or U522 (N_522,In_904,In_342);
xnor U523 (N_523,In_1709,In_890);
xor U524 (N_524,In_799,In_426);
nor U525 (N_525,N_265,N_104);
nor U526 (N_526,N_338,In_1222);
xnor U527 (N_527,In_446,In_684);
xor U528 (N_528,In_157,In_1689);
xnor U529 (N_529,In_210,In_2317);
and U530 (N_530,In_2032,N_490);
nand U531 (N_531,In_597,In_816);
or U532 (N_532,In_1406,In_404);
and U533 (N_533,In_1213,In_1702);
nor U534 (N_534,In_1914,In_2197);
and U535 (N_535,N_406,In_1000);
or U536 (N_536,N_303,N_448);
nand U537 (N_537,In_448,In_1047);
nor U538 (N_538,In_2023,In_1661);
nand U539 (N_539,In_856,In_2143);
or U540 (N_540,In_2008,N_368);
nand U541 (N_541,In_556,In_2178);
xor U542 (N_542,In_1676,In_2065);
xnor U543 (N_543,In_1952,In_2462);
nor U544 (N_544,N_407,In_167);
nand U545 (N_545,In_1745,In_687);
xor U546 (N_546,In_2114,In_2332);
or U547 (N_547,In_1917,In_1123);
and U548 (N_548,In_358,In_2410);
or U549 (N_549,In_551,In_201);
and U550 (N_550,N_176,N_323);
and U551 (N_551,In_643,N_95);
xnor U552 (N_552,In_1489,In_1701);
or U553 (N_553,N_400,In_1808);
nor U554 (N_554,In_1197,N_437);
xnor U555 (N_555,In_1283,In_869);
xor U556 (N_556,In_1815,N_262);
or U557 (N_557,In_506,In_1810);
and U558 (N_558,In_2293,N_233);
nand U559 (N_559,In_466,In_28);
nand U560 (N_560,In_1448,In_128);
or U561 (N_561,In_1058,In_1320);
xnor U562 (N_562,In_1159,In_1192);
xnor U563 (N_563,In_2239,In_432);
xnor U564 (N_564,In_722,In_2234);
or U565 (N_565,In_590,N_174);
and U566 (N_566,In_1768,N_494);
or U567 (N_567,N_28,In_185);
nand U568 (N_568,In_1822,In_2357);
and U569 (N_569,In_754,N_362);
nor U570 (N_570,In_1788,In_159);
nand U571 (N_571,In_1746,In_1541);
or U572 (N_572,N_264,In_1655);
or U573 (N_573,In_937,In_1949);
and U574 (N_574,In_1104,In_1739);
and U575 (N_575,In_780,In_690);
and U576 (N_576,In_472,In_1955);
and U577 (N_577,N_435,In_2160);
nor U578 (N_578,In_1512,In_1462);
nor U579 (N_579,In_2289,In_1753);
and U580 (N_580,In_1010,N_498);
xnor U581 (N_581,In_2421,In_2125);
nor U582 (N_582,In_2341,In_1972);
nor U583 (N_583,In_269,N_237);
xnor U584 (N_584,In_2044,In_539);
nand U585 (N_585,In_242,In_1033);
or U586 (N_586,In_2408,In_2376);
xnor U587 (N_587,N_8,N_219);
and U588 (N_588,In_427,In_1518);
xor U589 (N_589,In_1182,In_1947);
nand U590 (N_590,In_33,In_1960);
xor U591 (N_591,N_272,N_326);
or U592 (N_592,N_351,N_155);
and U593 (N_593,N_416,In_725);
and U594 (N_594,In_1821,N_430);
and U595 (N_595,In_1429,In_475);
and U596 (N_596,In_617,In_1407);
nor U597 (N_597,N_227,In_2389);
and U598 (N_598,In_2104,In_678);
and U599 (N_599,In_2452,N_109);
and U600 (N_600,In_1339,In_805);
or U601 (N_601,In_1064,In_2333);
and U602 (N_602,In_2240,N_409);
xnor U603 (N_603,In_581,In_347);
nand U604 (N_604,In_2313,N_91);
xnor U605 (N_605,In_1958,In_1500);
nand U606 (N_606,In_1139,In_881);
xor U607 (N_607,In_2221,In_1435);
xnor U608 (N_608,In_2312,In_998);
xnor U609 (N_609,In_1693,In_1071);
and U610 (N_610,In_1586,In_1521);
and U611 (N_611,In_2205,In_450);
xnor U612 (N_612,In_1896,In_360);
nor U613 (N_613,In_2466,N_125);
and U614 (N_614,In_38,In_2066);
or U615 (N_615,N_22,In_531);
and U616 (N_616,In_1966,N_370);
or U617 (N_617,In_1796,In_1425);
nand U618 (N_618,In_1277,In_372);
or U619 (N_619,N_342,In_193);
nand U620 (N_620,In_243,In_1922);
or U621 (N_621,In_1110,In_2247);
and U622 (N_622,In_1073,In_1714);
nand U623 (N_623,In_554,In_440);
xnor U624 (N_624,N_186,In_22);
nor U625 (N_625,N_160,In_1759);
and U626 (N_626,In_1513,In_1456);
or U627 (N_627,In_328,In_316);
nand U628 (N_628,N_236,In_2031);
nand U629 (N_629,In_1036,N_486);
and U630 (N_630,In_1551,In_2278);
xor U631 (N_631,N_77,N_248);
nor U632 (N_632,In_950,In_647);
xnor U633 (N_633,In_1858,N_27);
nor U634 (N_634,In_624,N_472);
nor U635 (N_635,N_221,In_2051);
nand U636 (N_636,In_2422,In_304);
and U637 (N_637,In_1202,In_1483);
and U638 (N_638,In_911,In_843);
nand U639 (N_639,In_1091,In_802);
xor U640 (N_640,In_1120,N_41);
nor U641 (N_641,In_2374,In_1142);
xor U642 (N_642,In_36,In_892);
xor U643 (N_643,In_1226,In_2461);
nand U644 (N_644,N_369,In_1803);
nor U645 (N_645,In_752,In_655);
xor U646 (N_646,In_397,In_1111);
or U647 (N_647,In_14,In_2018);
or U648 (N_648,In_777,In_2222);
nor U649 (N_649,In_81,In_1957);
nor U650 (N_650,N_88,N_115);
and U651 (N_651,N_478,In_1569);
and U652 (N_652,In_216,N_80);
and U653 (N_653,In_412,In_1617);
and U654 (N_654,In_10,In_848);
nor U655 (N_655,In_1571,In_220);
or U656 (N_656,In_1078,In_296);
or U657 (N_657,In_425,In_1107);
nor U658 (N_658,In_129,In_158);
or U659 (N_659,N_103,In_1675);
or U660 (N_660,In_1009,In_1736);
or U661 (N_661,In_779,In_262);
nand U662 (N_662,In_27,In_1790);
nor U663 (N_663,In_2152,N_78);
xnor U664 (N_664,In_335,In_969);
nor U665 (N_665,N_10,N_341);
xor U666 (N_666,N_101,In_371);
nor U667 (N_667,In_771,N_210);
xor U668 (N_668,In_1884,In_822);
nor U669 (N_669,In_2140,In_1664);
and U670 (N_670,In_2270,In_2471);
nand U671 (N_671,In_662,N_162);
or U672 (N_672,In_1167,In_598);
nor U673 (N_673,In_509,N_373);
nand U674 (N_674,In_2175,In_2348);
xnor U675 (N_675,In_650,N_310);
nand U676 (N_676,In_380,In_2424);
nor U677 (N_677,In_2212,In_501);
and U678 (N_678,In_1346,In_828);
xnor U679 (N_679,N_330,In_334);
and U680 (N_680,N_97,In_208);
nand U681 (N_681,In_1385,In_2068);
nor U682 (N_682,In_1497,N_455);
xnor U683 (N_683,In_1254,In_2264);
xnor U684 (N_684,In_377,In_628);
xnor U685 (N_685,In_1444,In_1938);
or U686 (N_686,In_1633,In_785);
nor U687 (N_687,In_632,In_1856);
xor U688 (N_688,In_1602,N_159);
and U689 (N_689,N_355,In_44);
xor U690 (N_690,In_2181,In_436);
and U691 (N_691,In_1581,N_347);
nor U692 (N_692,In_1144,N_242);
nor U693 (N_693,In_2131,In_2168);
or U694 (N_694,In_1686,N_216);
or U695 (N_695,In_1162,In_618);
xor U696 (N_696,In_1680,In_2352);
nor U697 (N_697,In_2036,In_249);
xor U698 (N_698,N_247,N_223);
nor U699 (N_699,N_51,In_1496);
or U700 (N_700,In_2354,N_357);
nand U701 (N_701,N_328,In_1901);
xor U702 (N_702,N_287,In_524);
and U703 (N_703,In_259,In_278);
nand U704 (N_704,N_483,In_941);
nor U705 (N_705,In_1981,In_739);
nor U706 (N_706,N_276,In_1430);
and U707 (N_707,In_1424,In_101);
nor U708 (N_708,In_260,N_489);
and U709 (N_709,In_1611,N_291);
nor U710 (N_710,In_135,N_319);
xor U711 (N_711,In_2099,In_1115);
nor U712 (N_712,In_732,In_1652);
xor U713 (N_713,In_1322,N_110);
or U714 (N_714,In_566,In_2213);
or U715 (N_715,In_2450,In_1687);
nand U716 (N_716,In_839,In_1499);
or U717 (N_717,In_2492,In_1209);
xnor U718 (N_718,In_826,In_2482);
or U719 (N_719,In_1249,N_6);
or U720 (N_720,N_306,In_721);
and U721 (N_721,In_1258,In_2056);
nor U722 (N_722,In_56,In_1126);
nor U723 (N_723,In_1158,In_1639);
and U724 (N_724,In_2201,In_1622);
nand U725 (N_725,N_68,In_1548);
nor U726 (N_726,N_23,N_100);
nor U727 (N_727,N_383,N_302);
nor U728 (N_728,In_403,In_978);
nor U729 (N_729,In_2440,In_117);
nor U730 (N_730,In_2025,In_1614);
xor U731 (N_731,In_563,In_745);
nand U732 (N_732,In_1700,In_1);
and U733 (N_733,In_626,In_2412);
and U734 (N_734,In_1558,N_366);
nor U735 (N_735,N_349,In_2401);
and U736 (N_736,In_1795,In_1007);
nor U737 (N_737,In_1669,In_2198);
nand U738 (N_738,In_1925,In_1001);
nand U739 (N_739,N_201,In_2191);
or U740 (N_740,N_497,In_521);
nor U741 (N_741,In_1959,In_3);
nand U742 (N_742,In_1414,N_444);
nand U743 (N_743,N_190,In_1575);
xor U744 (N_744,In_1506,In_1475);
xor U745 (N_745,In_311,In_351);
and U746 (N_746,In_946,In_949);
or U747 (N_747,In_529,In_2169);
and U748 (N_748,In_1225,In_1557);
xor U749 (N_749,In_2211,In_2116);
nor U750 (N_750,In_6,In_571);
xor U751 (N_751,In_587,N_651);
xor U752 (N_752,In_381,In_439);
or U753 (N_753,In_2078,In_801);
xnor U754 (N_754,In_783,In_1211);
or U755 (N_755,N_337,In_1715);
nor U756 (N_756,N_538,N_364);
nor U757 (N_757,N_495,In_214);
or U758 (N_758,In_1418,N_715);
xnor U759 (N_759,In_1580,In_1846);
nor U760 (N_760,N_134,In_1660);
or U761 (N_761,N_53,N_621);
or U762 (N_762,In_1593,N_92);
nand U763 (N_763,In_576,In_1653);
or U764 (N_764,N_743,In_2096);
or U765 (N_765,In_1199,In_2369);
nand U766 (N_766,In_252,N_76);
nor U767 (N_767,N_457,N_420);
or U768 (N_768,N_574,N_471);
and U769 (N_769,N_545,N_573);
xor U770 (N_770,N_718,In_2005);
and U771 (N_771,In_221,In_273);
nand U772 (N_772,N_377,In_2497);
xnor U773 (N_773,In_65,In_1476);
nor U774 (N_774,In_2460,In_392);
nor U775 (N_775,In_885,In_1267);
or U776 (N_776,In_1179,In_1775);
xnor U777 (N_777,In_1235,N_639);
and U778 (N_778,N_313,N_659);
xnor U779 (N_779,In_104,In_2328);
nand U780 (N_780,In_1712,In_1744);
xnor U781 (N_781,N_352,In_1885);
nand U782 (N_782,In_79,In_1498);
or U783 (N_783,N_417,In_379);
nand U784 (N_784,In_1584,N_292);
or U785 (N_785,In_855,In_82);
or U786 (N_786,In_1484,In_676);
and U787 (N_787,In_1330,N_592);
nor U788 (N_788,In_894,N_402);
xnor U789 (N_789,In_156,In_1092);
and U790 (N_790,In_741,In_808);
xnor U791 (N_791,In_923,N_181);
nor U792 (N_792,In_281,In_1556);
nor U793 (N_793,In_137,In_1371);
or U794 (N_794,N_532,N_589);
or U795 (N_795,In_2124,In_2165);
xnor U796 (N_796,N_695,N_169);
xnor U797 (N_797,N_256,In_1798);
xnor U798 (N_798,In_1263,In_1773);
nand U799 (N_799,In_2055,In_2455);
nor U800 (N_800,N_157,In_1649);
nor U801 (N_801,N_44,In_812);
and U802 (N_802,In_1097,N_511);
nand U803 (N_803,In_857,In_433);
xor U804 (N_804,N_37,N_662);
xnor U805 (N_805,In_527,N_428);
and U806 (N_806,In_948,N_132);
nor U807 (N_807,In_459,N_403);
and U808 (N_808,In_409,N_587);
xor U809 (N_809,In_1223,In_883);
xnor U810 (N_810,In_1970,In_964);
nand U811 (N_811,In_1845,In_2072);
xor U812 (N_812,In_1176,In_382);
and U813 (N_813,In_487,N_597);
or U814 (N_814,In_357,In_1761);
and U815 (N_815,In_1079,N_493);
nor U816 (N_816,N_73,N_672);
and U817 (N_817,N_660,In_1378);
or U818 (N_818,In_297,In_1027);
nand U819 (N_819,In_516,N_127);
and U820 (N_820,N_726,In_2153);
xor U821 (N_821,In_1621,N_322);
or U822 (N_822,In_1716,In_623);
or U823 (N_823,N_530,In_1538);
nor U824 (N_824,N_636,N_723);
nor U825 (N_825,N_4,N_454);
xor U826 (N_826,In_1319,In_2118);
xnor U827 (N_827,N_655,N_481);
nor U828 (N_828,N_567,In_1508);
nand U829 (N_829,N_588,In_1367);
or U830 (N_830,In_2409,N_513);
nor U831 (N_831,In_968,N_193);
xnor U832 (N_832,In_1083,N_544);
nand U833 (N_833,In_870,N_590);
nor U834 (N_834,In_495,In_734);
xor U835 (N_835,In_1789,In_2428);
or U836 (N_836,In_2147,In_251);
xnor U837 (N_837,In_1148,In_743);
nand U838 (N_838,In_715,In_1312);
and U839 (N_839,In_1350,N_559);
nor U840 (N_840,In_1299,In_1216);
nand U841 (N_841,In_1457,In_1632);
xor U842 (N_842,In_2375,In_255);
nor U843 (N_843,In_1410,N_2);
or U844 (N_844,N_183,In_1670);
or U845 (N_845,In_1085,In_341);
nand U846 (N_846,In_988,In_2404);
and U847 (N_847,In_1166,In_867);
and U848 (N_848,In_1839,N_721);
or U849 (N_849,N_24,N_84);
or U850 (N_850,In_2105,In_2291);
xnor U851 (N_851,In_1540,N_244);
and U852 (N_852,In_2046,In_32);
and U853 (N_853,In_2337,N_467);
nand U854 (N_854,In_2048,N_595);
xor U855 (N_855,In_2080,In_406);
nand U856 (N_856,In_499,In_2284);
xor U857 (N_857,N_623,In_97);
or U858 (N_858,In_1019,In_289);
and U859 (N_859,In_612,In_353);
or U860 (N_860,N_126,In_1380);
or U861 (N_861,In_279,N_657);
and U862 (N_862,N_488,N_235);
nand U863 (N_863,N_165,In_12);
xor U864 (N_864,N_576,In_1971);
and U865 (N_865,In_2101,N_543);
nand U866 (N_866,N_131,In_884);
xor U867 (N_867,In_150,N_554);
and U868 (N_868,In_1881,In_2288);
xnor U869 (N_869,In_636,In_1997);
or U870 (N_870,In_728,In_760);
nor U871 (N_871,N_273,In_2155);
nand U872 (N_872,In_975,N_270);
and U873 (N_873,In_467,In_1365);
xnor U874 (N_874,In_2003,In_428);
nor U875 (N_875,In_2050,In_1844);
nand U876 (N_876,N_484,In_1812);
and U877 (N_877,In_1890,In_196);
and U878 (N_878,N_667,N_617);
or U879 (N_879,N_410,N_586);
nor U880 (N_880,N_424,N_604);
or U881 (N_881,N_534,N_474);
or U882 (N_882,In_1817,In_2384);
and U883 (N_883,In_2127,In_1504);
nor U884 (N_884,In_2053,N_681);
xor U885 (N_885,In_234,In_683);
and U886 (N_886,In_738,In_326);
and U887 (N_887,In_1733,In_1465);
xnor U888 (N_888,In_1867,N_111);
nand U889 (N_889,N_329,N_246);
nor U890 (N_890,N_376,In_1005);
nor U891 (N_891,In_2136,N_569);
nor U892 (N_892,In_1996,In_368);
and U893 (N_893,In_93,N_482);
xor U894 (N_894,In_1262,In_954);
or U895 (N_895,N_507,N_215);
nand U896 (N_896,N_197,N_81);
or U897 (N_897,In_131,In_1096);
xnor U898 (N_898,N_466,In_1603);
and U899 (N_899,In_455,In_186);
nor U900 (N_900,In_2139,In_2215);
xor U901 (N_901,In_52,In_202);
nor U902 (N_902,N_468,In_873);
nand U903 (N_903,In_951,In_842);
nor U904 (N_904,In_784,N_675);
xnor U905 (N_905,N_282,In_2042);
nor U906 (N_906,In_1751,In_1681);
nor U907 (N_907,N_213,In_541);
nor U908 (N_908,In_154,In_520);
and U909 (N_909,N_656,In_891);
xor U910 (N_910,N_185,In_405);
and U911 (N_911,In_1729,N_685);
nand U912 (N_912,N_143,In_1616);
and U913 (N_913,In_479,In_644);
xor U914 (N_914,In_2266,In_434);
nor U915 (N_915,In_1493,N_187);
xnor U916 (N_916,In_580,In_2347);
or U917 (N_917,N_422,In_1180);
or U918 (N_918,N_427,N_324);
xor U919 (N_919,In_1168,In_388);
xnor U920 (N_920,In_5,In_1979);
or U921 (N_921,In_606,N_611);
and U922 (N_922,In_2302,N_348);
nand U923 (N_923,N_434,N_729);
xnor U924 (N_924,In_344,N_456);
nand U925 (N_925,N_480,In_224);
nor U926 (N_926,In_2368,In_1705);
nand U927 (N_927,N_740,In_1526);
or U928 (N_928,In_994,In_2202);
xor U929 (N_929,N_654,N_503);
or U930 (N_930,N_696,In_1415);
xnor U931 (N_931,N_378,In_546);
or U932 (N_932,In_1053,In_561);
nor U933 (N_933,N_112,In_534);
xnor U934 (N_934,In_2035,In_1391);
nand U935 (N_935,In_2180,In_1943);
and U936 (N_936,N_50,In_1585);
nor U937 (N_937,In_250,In_1539);
nand U938 (N_938,In_416,N_555);
nor U939 (N_939,In_876,N_311);
nor U940 (N_940,N_533,In_359);
and U941 (N_941,N_297,In_2495);
or U942 (N_942,In_2292,N_314);
nor U943 (N_943,In_1337,In_766);
nor U944 (N_944,In_757,N_519);
and U945 (N_945,In_460,N_354);
or U946 (N_946,In_1565,In_336);
xnor U947 (N_947,In_552,In_189);
xor U948 (N_948,In_441,In_2290);
and U949 (N_949,In_1673,In_707);
or U950 (N_950,N_372,N_460);
or U951 (N_951,N_316,In_2437);
or U952 (N_952,N_698,N_644);
xnor U953 (N_953,N_177,In_288);
and U954 (N_954,In_1634,In_711);
xnor U955 (N_955,In_847,In_702);
nand U956 (N_956,In_2244,In_1102);
and U957 (N_957,In_1785,In_1470);
nor U958 (N_958,N_281,In_1933);
or U959 (N_959,N_375,In_66);
and U960 (N_960,In_2308,In_1926);
and U961 (N_961,In_271,N_140);
nand U962 (N_962,In_1469,N_575);
xnor U963 (N_963,In_2085,In_1624);
and U964 (N_964,In_795,In_58);
and U965 (N_965,In_2200,N_54);
nor U966 (N_966,In_1134,In_2161);
and U967 (N_967,In_149,In_1942);
or U968 (N_968,In_548,In_1398);
nor U969 (N_969,In_573,In_2195);
xor U970 (N_970,In_2316,N_652);
or U971 (N_971,N_31,N_463);
nand U972 (N_972,N_358,In_2233);
nor U973 (N_973,N_266,In_789);
and U974 (N_974,N_491,N_299);
nand U975 (N_975,In_763,N_42);
xor U976 (N_976,In_254,N_650);
nor U977 (N_977,In_1604,In_1722);
and U978 (N_978,In_2209,In_1754);
xor U979 (N_979,N_89,In_258);
and U980 (N_980,In_264,In_1062);
nand U981 (N_981,N_607,N_649);
nor U982 (N_982,In_1802,In_465);
and U983 (N_983,In_23,In_1907);
nor U984 (N_984,In_1230,In_1345);
xor U985 (N_985,In_1684,In_1246);
and U986 (N_986,N_212,N_114);
xor U987 (N_987,In_464,In_979);
nor U988 (N_988,N_361,In_1368);
xor U989 (N_989,N_431,N_234);
and U990 (N_990,N_625,N_705);
and U991 (N_991,In_1321,N_350);
and U992 (N_992,N_459,In_1114);
xor U993 (N_993,In_585,N_433);
and U994 (N_994,In_1573,In_1305);
nor U995 (N_995,N_398,In_228);
xor U996 (N_996,N_746,In_50);
and U997 (N_997,In_1961,N_564);
and U998 (N_998,N_139,N_142);
nand U999 (N_999,In_102,In_2467);
or U1000 (N_1000,N_928,In_1663);
xor U1001 (N_1001,N_736,N_207);
xnor U1002 (N_1002,In_1383,In_272);
or U1003 (N_1003,In_1400,N_194);
or U1004 (N_1004,In_661,N_745);
nand U1005 (N_1005,In_2338,In_1014);
and U1006 (N_1006,In_907,N_948);
or U1007 (N_1007,In_1308,In_267);
and U1008 (N_1008,In_483,N_295);
nand U1009 (N_1009,In_1349,N_699);
xnor U1010 (N_1010,In_935,In_438);
or U1011 (N_1011,N_811,N_570);
nor U1012 (N_1012,In_486,In_1431);
nor U1013 (N_1013,In_2380,N_790);
and U1014 (N_1014,N_419,In_85);
nand U1015 (N_1015,N_756,In_1578);
xor U1016 (N_1016,N_881,N_815);
nand U1017 (N_1017,In_1732,N_970);
nor U1018 (N_1018,N_11,In_1108);
and U1019 (N_1019,In_1900,N_500);
or U1020 (N_1020,N_582,In_1239);
or U1021 (N_1021,N_548,In_2367);
nor U1022 (N_1022,In_1640,In_549);
or U1023 (N_1023,In_1113,In_8);
and U1024 (N_1024,N_211,In_1393);
nand U1025 (N_1025,In_653,In_1170);
or U1026 (N_1026,In_91,N_462);
or U1027 (N_1027,In_84,In_1517);
nand U1028 (N_1028,In_2190,In_1595);
nor U1029 (N_1029,In_1076,In_508);
or U1030 (N_1030,N_845,N_732);
and U1031 (N_1031,In_1555,In_1523);
or U1032 (N_1032,In_542,In_2013);
or U1033 (N_1033,N_676,In_2296);
xnor U1034 (N_1034,In_1044,N_268);
nor U1035 (N_1035,In_638,N_747);
xnor U1036 (N_1036,In_1991,In_2478);
nor U1037 (N_1037,In_518,In_1707);
nor U1038 (N_1038,In_391,In_1505);
nor U1039 (N_1039,N_794,N_761);
and U1040 (N_1040,In_1743,N_166);
nand U1041 (N_1041,N_759,N_20);
xor U1042 (N_1042,In_821,N_154);
or U1043 (N_1043,N_767,In_792);
or U1044 (N_1044,N_653,In_2442);
nor U1045 (N_1045,In_1730,In_77);
nor U1046 (N_1046,In_1771,In_2192);
and U1047 (N_1047,N_72,N_365);
nand U1048 (N_1048,In_1106,N_848);
nor U1049 (N_1049,N_240,N_5);
or U1050 (N_1050,In_118,In_2464);
and U1051 (N_1051,N_918,In_1968);
or U1052 (N_1052,In_1187,N_620);
or U1053 (N_1053,In_1855,N_933);
or U1054 (N_1054,In_447,In_1276);
xnor U1055 (N_1055,In_1026,In_300);
nand U1056 (N_1056,In_1953,In_155);
xor U1057 (N_1057,N_753,In_2009);
or U1058 (N_1058,N_325,In_2049);
xor U1059 (N_1059,N_285,N_867);
xnor U1060 (N_1060,N_439,N_188);
nor U1061 (N_1061,N_541,In_1388);
and U1062 (N_1062,In_113,N_757);
nand U1063 (N_1063,In_2022,In_2199);
or U1064 (N_1064,In_2041,In_1006);
or U1065 (N_1065,N_563,N_831);
xnor U1066 (N_1066,In_2071,N_516);
xnor U1067 (N_1067,In_317,N_476);
nand U1068 (N_1068,In_1124,N_885);
xnor U1069 (N_1069,N_445,N_175);
nand U1070 (N_1070,N_844,N_606);
and U1071 (N_1071,In_1067,In_665);
xnor U1072 (N_1072,N_637,In_1738);
or U1073 (N_1073,In_1023,In_1354);
nor U1074 (N_1074,N_260,N_164);
and U1075 (N_1075,In_577,N_825);
nor U1076 (N_1076,N_388,N_118);
xor U1077 (N_1077,In_2274,In_286);
nor U1078 (N_1078,In_2378,N_751);
and U1079 (N_1079,In_2271,N_996);
nor U1080 (N_1080,In_1524,In_1760);
nor U1081 (N_1081,In_2110,In_2469);
and U1082 (N_1082,In_2237,In_1173);
nand U1083 (N_1083,In_1440,In_2496);
and U1084 (N_1084,N_624,N_977);
xnor U1085 (N_1085,In_223,N_791);
and U1086 (N_1086,N_784,In_2128);
or U1087 (N_1087,In_2310,In_2340);
nand U1088 (N_1088,N_271,N_713);
or U1089 (N_1089,N_128,N_926);
xnor U1090 (N_1090,N_722,In_2067);
nor U1091 (N_1091,N_551,In_1487);
nor U1092 (N_1092,N_731,N_613);
xnor U1093 (N_1093,In_677,N_773);
nor U1094 (N_1094,In_958,N_897);
and U1095 (N_1095,N_49,In_1082);
nand U1096 (N_1096,In_1317,In_1688);
nand U1097 (N_1097,In_2137,In_1020);
xnor U1098 (N_1098,In_1458,N_778);
and U1099 (N_1099,N_214,In_1125);
and U1100 (N_1100,N_749,In_244);
nand U1101 (N_1101,N_941,N_911);
nor U1102 (N_1102,N_924,N_980);
nand U1103 (N_1103,In_139,N_560);
xor U1104 (N_1104,In_1093,In_1074);
and U1105 (N_1105,In_522,N_878);
or U1106 (N_1106,N_279,N_395);
nor U1107 (N_1107,N_907,In_2407);
or U1108 (N_1108,N_141,N_988);
nor U1109 (N_1109,In_2260,N_305);
or U1110 (N_1110,In_2479,In_2415);
nor U1111 (N_1111,In_430,N_46);
or U1112 (N_1112,In_1950,N_631);
nand U1113 (N_1113,In_629,In_1537);
and U1114 (N_1114,In_1778,In_2331);
nor U1115 (N_1115,In_1731,N_922);
or U1116 (N_1116,In_919,N_807);
or U1117 (N_1117,In_290,In_1016);
xor U1118 (N_1118,In_1109,N_906);
or U1119 (N_1119,N_967,In_1704);
nand U1120 (N_1120,In_1041,In_1490);
nand U1121 (N_1121,In_1227,N_738);
xor U1122 (N_1122,N_994,In_999);
nand U1123 (N_1123,In_582,In_1220);
or U1124 (N_1124,In_1069,In_2268);
xor U1125 (N_1125,In_1224,In_824);
nand U1126 (N_1126,In_2062,In_1678);
xor U1127 (N_1127,N_339,N_254);
and U1128 (N_1128,N_208,N_813);
xnor U1129 (N_1129,In_1756,N_429);
or U1130 (N_1130,In_1335,In_1590);
nor U1131 (N_1131,N_577,In_1924);
nand U1132 (N_1132,In_2208,N_981);
or U1133 (N_1133,In_2002,N_716);
nor U1134 (N_1134,In_670,N_678);
nor U1135 (N_1135,N_979,N_701);
nor U1136 (N_1136,N_635,In_709);
or U1137 (N_1137,N_987,N_733);
and U1138 (N_1138,In_865,N_944);
nor U1139 (N_1139,N_777,In_2142);
or U1140 (N_1140,N_808,In_770);
nor U1141 (N_1141,N_399,In_232);
or U1142 (N_1142,N_340,In_1261);
or U1143 (N_1143,N_43,N_571);
and U1144 (N_1144,N_724,N_797);
nand U1145 (N_1145,In_174,In_2356);
nor U1146 (N_1146,N_810,In_2070);
and U1147 (N_1147,N_990,In_671);
nor U1148 (N_1148,In_1699,In_878);
or U1149 (N_1149,In_1215,N_605);
nand U1150 (N_1150,N_786,N_998);
nor U1151 (N_1151,In_1439,In_517);
xor U1152 (N_1152,N_891,N_321);
or U1153 (N_1153,N_130,N_397);
and U1154 (N_1154,In_1219,N_156);
or U1155 (N_1155,N_492,In_716);
xnor U1156 (N_1156,In_1360,In_1902);
nor U1157 (N_1157,In_106,N_294);
or U1158 (N_1158,N_286,N_556);
nand U1159 (N_1159,In_1851,In_237);
xnor U1160 (N_1160,In_2121,N_799);
xor U1161 (N_1161,In_1477,N_334);
nand U1162 (N_1162,In_422,In_1060);
and U1163 (N_1163,In_1974,N_983);
xnor U1164 (N_1164,In_2443,N_816);
xnor U1165 (N_1165,In_195,N_930);
and U1166 (N_1166,N_847,In_536);
nor U1167 (N_1167,N_547,N_785);
nand U1168 (N_1168,In_1606,In_323);
or U1169 (N_1169,N_144,N_381);
xnor U1170 (N_1170,In_330,N_835);
xnor U1171 (N_1171,In_2102,N_204);
and U1172 (N_1172,N_572,In_68);
nor U1173 (N_1173,N_958,In_470);
nand U1174 (N_1174,In_1127,In_2494);
or U1175 (N_1175,In_2206,In_461);
or U1176 (N_1176,In_1748,N_250);
nand U1177 (N_1177,In_21,N_971);
or U1178 (N_1178,N_296,In_1637);
and U1179 (N_1179,In_820,N_568);
and U1180 (N_1180,N_895,In_1420);
nand U1181 (N_1181,In_2001,N_510);
nor U1182 (N_1182,In_1240,N_682);
and U1183 (N_1183,N_982,N_951);
nand U1184 (N_1184,N_823,In_1405);
nor U1185 (N_1185,In_369,N_261);
and U1186 (N_1186,In_1291,In_1089);
nand U1187 (N_1187,In_212,In_34);
nand U1188 (N_1188,N_939,In_744);
and U1189 (N_1189,In_1428,In_500);
nand U1190 (N_1190,In_1447,N_883);
or U1191 (N_1191,In_1857,N_107);
and U1192 (N_1192,N_601,In_2436);
and U1193 (N_1193,In_96,In_938);
or U1194 (N_1194,N_594,N_451);
and U1195 (N_1195,In_727,In_1482);
nor U1196 (N_1196,In_110,In_2220);
and U1197 (N_1197,N_367,In_1635);
nand U1198 (N_1198,N_1,In_1063);
nor U1199 (N_1199,N_765,N_509);
and U1200 (N_1200,In_1233,N_857);
xor U1201 (N_1201,In_1615,N_935);
xor U1202 (N_1202,N_889,In_1609);
and U1203 (N_1203,In_1692,N_36);
and U1204 (N_1204,In_1904,In_1141);
nand U1205 (N_1205,In_642,In_528);
nand U1206 (N_1206,N_638,In_511);
nor U1207 (N_1207,In_1002,In_2225);
xor U1208 (N_1208,N_228,N_683);
xor U1209 (N_1209,N_677,In_1087);
or U1210 (N_1210,In_322,N_608);
and U1211 (N_1211,N_934,In_1363);
nand U1212 (N_1212,In_2277,In_1740);
and U1213 (N_1213,In_1980,N_628);
nand U1214 (N_1214,N_238,In_308);
and U1215 (N_1215,N_993,N_630);
and U1216 (N_1216,In_845,N_663);
and U1217 (N_1217,In_1577,In_1903);
and U1218 (N_1218,N_838,N_909);
and U1219 (N_1219,In_1459,In_2269);
nand U1220 (N_1220,N_855,N_833);
xnor U1221 (N_1221,In_1833,In_888);
and U1222 (N_1222,In_2257,N_943);
and U1223 (N_1223,In_1326,In_1804);
and U1224 (N_1224,In_1485,N_814);
or U1225 (N_1225,In_1583,In_1478);
nand U1226 (N_1226,N_854,N_642);
xor U1227 (N_1227,In_2459,N_449);
and U1228 (N_1228,In_2359,In_226);
and U1229 (N_1229,In_1849,In_1536);
and U1230 (N_1230,In_2145,N_557);
nand U1231 (N_1231,In_2342,In_1656);
nand U1232 (N_1232,N_371,In_2414);
and U1233 (N_1233,In_2111,N_106);
nor U1234 (N_1234,In_2259,N_972);
xnor U1235 (N_1235,N_562,In_773);
xnor U1236 (N_1236,In_537,In_1193);
nand U1237 (N_1237,In_1679,In_976);
nand U1238 (N_1238,In_1105,N_206);
or U1239 (N_1239,In_863,In_731);
xnor U1240 (N_1240,In_1919,N_879);
and U1241 (N_1241,N_404,In_1212);
xnor U1242 (N_1242,N_775,In_778);
or U1243 (N_1243,N_865,N_229);
or U1244 (N_1244,N_550,In_1454);
nand U1245 (N_1245,N_565,N_346);
nand U1246 (N_1246,In_2052,In_1764);
xor U1247 (N_1247,N_824,N_647);
and U1248 (N_1248,In_1691,In_55);
and U1249 (N_1249,In_611,In_2261);
nand U1250 (N_1250,In_2299,In_2306);
and U1251 (N_1251,N_253,N_1130);
and U1252 (N_1252,In_1358,In_2109);
xor U1253 (N_1253,N_748,In_1735);
nor U1254 (N_1254,In_241,N_1222);
nand U1255 (N_1255,N_750,In_298);
nand U1256 (N_1256,N_30,N_822);
or U1257 (N_1257,In_1905,In_1101);
nand U1258 (N_1258,In_306,N_684);
nand U1259 (N_1259,In_2282,N_1146);
nor U1260 (N_1260,N_793,N_405);
or U1261 (N_1261,In_1285,N_744);
and U1262 (N_1262,N_300,N_692);
or U1263 (N_1263,N_93,In_1723);
or U1264 (N_1264,N_1097,In_2499);
or U1265 (N_1265,N_633,N_634);
or U1266 (N_1266,N_135,N_1075);
and U1267 (N_1267,In_868,N_871);
and U1268 (N_1268,In_321,N_940);
and U1269 (N_1269,N_553,In_1467);
nor U1270 (N_1270,In_419,In_667);
nand U1271 (N_1271,In_2249,In_834);
xnor U1272 (N_1272,N_389,N_290);
nand U1273 (N_1273,N_1005,N_788);
nand U1274 (N_1274,N_664,In_695);
nor U1275 (N_1275,N_714,N_1206);
nand U1276 (N_1276,In_2011,N_852);
or U1277 (N_1277,In_2226,N_717);
nand U1278 (N_1278,In_1516,In_88);
and U1279 (N_1279,In_1260,In_1995);
or U1280 (N_1280,N_26,In_2458);
or U1281 (N_1281,N_758,N_999);
and U1282 (N_1282,N_789,N_1122);
and U1283 (N_1283,N_1216,N_742);
nor U1284 (N_1284,N_1169,N_458);
and U1285 (N_1285,N_1175,N_385);
and U1286 (N_1286,N_1007,N_1118);
and U1287 (N_1287,In_1696,N_1162);
nand U1288 (N_1288,In_2235,N_304);
nor U1289 (N_1289,N_1208,N_317);
and U1290 (N_1290,In_803,N_191);
xnor U1291 (N_1291,N_1243,In_1892);
nand U1292 (N_1292,N_390,In_813);
nor U1293 (N_1293,In_1003,N_936);
nor U1294 (N_1294,In_120,N_1151);
xnor U1295 (N_1295,N_712,N_1084);
nand U1296 (N_1296,N_730,In_276);
nand U1297 (N_1297,N_1209,In_424);
xnor U1298 (N_1298,In_1204,In_2267);
nor U1299 (N_1299,In_61,In_1871);
nor U1300 (N_1300,In_15,N_163);
and U1301 (N_1301,In_2425,N_1159);
nor U1302 (N_1302,N_1137,In_1682);
xnor U1303 (N_1303,In_1024,In_2059);
nor U1304 (N_1304,In_1720,N_1114);
nor U1305 (N_1305,N_668,N_475);
and U1306 (N_1306,In_957,In_621);
xnor U1307 (N_1307,In_2097,In_640);
or U1308 (N_1308,In_2077,N_917);
and U1309 (N_1309,N_179,N_473);
or U1310 (N_1310,In_1547,N_309);
nand U1311 (N_1311,N_392,In_514);
or U1312 (N_1312,N_1198,In_1948);
nand U1313 (N_1313,N_283,In_1297);
nand U1314 (N_1314,N_1049,In_575);
or U1315 (N_1315,In_2301,N_552);
nor U1316 (N_1316,In_2324,N_1183);
and U1317 (N_1317,In_2248,N_946);
nand U1318 (N_1318,In_0,In_206);
nor U1319 (N_1319,In_1080,In_762);
nor U1320 (N_1320,In_2138,In_407);
and U1321 (N_1321,N_345,In_1646);
nor U1322 (N_1322,N_769,N_1157);
xor U1323 (N_1323,In_2093,N_1141);
nand U1324 (N_1324,N_527,N_1132);
nor U1325 (N_1325,N_87,N_1152);
or U1326 (N_1326,N_646,N_754);
nand U1327 (N_1327,N_1036,In_1300);
nand U1328 (N_1328,N_413,N_1013);
nand U1329 (N_1329,In_2024,N_591);
nand U1330 (N_1330,In_1098,N_184);
nor U1331 (N_1331,In_596,In_2020);
nand U1332 (N_1332,In_1304,In_376);
nor U1333 (N_1333,In_1338,N_356);
xor U1334 (N_1334,In_607,N_529);
and U1335 (N_1335,In_723,N_1020);
nand U1336 (N_1336,In_283,N_839);
and U1337 (N_1337,N_232,In_1031);
and U1338 (N_1338,In_444,In_1908);
nand U1339 (N_1339,N_1133,N_963);
and U1340 (N_1340,N_384,N_856);
or U1341 (N_1341,In_2480,N_17);
nand U1342 (N_1342,In_1519,N_780);
or U1343 (N_1343,In_2251,In_545);
nand U1344 (N_1344,In_248,In_39);
or U1345 (N_1345,N_752,In_1937);
nor U1346 (N_1346,In_1434,In_1874);
nand U1347 (N_1347,N_252,N_259);
nand U1348 (N_1348,In_2339,N_707);
xor U1349 (N_1349,N_566,N_826);
xor U1350 (N_1350,N_846,N_658);
or U1351 (N_1351,In_995,In_2449);
or U1352 (N_1352,In_1835,In_2090);
and U1353 (N_1353,N_1088,In_1030);
or U1354 (N_1354,In_952,N_258);
or U1355 (N_1355,In_1072,N_293);
or U1356 (N_1356,N_1149,N_945);
nor U1357 (N_1357,In_2064,N_955);
xor U1358 (N_1358,N_861,In_1206);
or U1359 (N_1359,N_205,N_1102);
xnor U1360 (N_1360,In_2091,In_1039);
nor U1361 (N_1361,N_446,In_1769);
and U1362 (N_1362,N_986,N_600);
nand U1363 (N_1363,N_1078,In_302);
and U1364 (N_1364,N_819,In_111);
xor U1365 (N_1365,In_1284,In_852);
xnor U1366 (N_1366,N_19,In_1293);
nor U1367 (N_1367,N_645,In_307);
xnor U1368 (N_1368,In_491,In_51);
nand U1369 (N_1369,N_1032,In_2194);
nand U1370 (N_1370,N_870,N_172);
nor U1371 (N_1371,In_1103,N_411);
nor U1372 (N_1372,N_616,N_688);
nand U1373 (N_1373,In_1563,In_619);
nor U1374 (N_1374,N_278,N_851);
xnor U1375 (N_1375,In_1807,N_1226);
nor U1376 (N_1376,N_1120,In_1099);
and U1377 (N_1377,N_1012,N_1034);
or U1378 (N_1378,N_1172,N_709);
or U1379 (N_1379,In_1452,In_1369);
or U1380 (N_1380,In_558,N_952);
and U1381 (N_1381,In_1765,N_843);
or U1382 (N_1382,In_2360,N_1037);
nor U1383 (N_1383,In_1665,N_916);
xnor U1384 (N_1384,In_1040,In_343);
nand U1385 (N_1385,N_1030,N_1143);
and U1386 (N_1386,In_203,In_462);
xnor U1387 (N_1387,In_959,N_643);
xor U1388 (N_1388,In_90,N_942);
nor U1389 (N_1389,N_336,N_522);
nor U1390 (N_1390,In_1301,In_913);
or U1391 (N_1391,N_487,In_1146);
nor U1392 (N_1392,In_112,N_122);
xor U1393 (N_1393,N_734,N_894);
and U1394 (N_1394,N_670,N_1031);
or U1395 (N_1395,N_1213,In_1843);
nor U1396 (N_1396,N_774,In_2193);
xnor U1397 (N_1397,N_968,In_2468);
nor U1398 (N_1398,N_360,In_2026);
or U1399 (N_1399,In_1025,In_1853);
xor U1400 (N_1400,N_720,In_1719);
nor U1401 (N_1401,N_1015,N_1077);
and U1402 (N_1402,N_1135,In_2372);
and U1403 (N_1403,In_1128,N_436);
and U1404 (N_1404,N_517,N_641);
nand U1405 (N_1405,N_779,N_1153);
nand U1406 (N_1406,N_612,In_2275);
or U1407 (N_1407,N_903,N_829);
and U1408 (N_1408,In_963,N_461);
and U1409 (N_1409,In_747,N_502);
and U1410 (N_1410,In_1862,In_1825);
nor U1411 (N_1411,N_453,In_437);
xnor U1412 (N_1412,In_1658,N_593);
or U1413 (N_1413,N_196,N_1022);
nand U1414 (N_1414,In_603,N_170);
nand U1415 (N_1415,In_1545,N_795);
and U1416 (N_1416,N_1192,N_1223);
nand U1417 (N_1417,N_969,In_98);
nand U1418 (N_1418,N_596,N_1204);
or U1419 (N_1419,N_1188,N_842);
or U1420 (N_1420,N_526,N_1167);
xnor U1421 (N_1421,In_364,N_710);
nand U1422 (N_1422,N_39,In_986);
xor U1423 (N_1423,N_1124,In_1860);
or U1424 (N_1424,N_380,N_812);
and U1425 (N_1425,N_168,N_919);
xor U1426 (N_1426,In_1836,In_1466);
nor U1427 (N_1427,In_2060,In_1965);
and U1428 (N_1428,N_536,In_2089);
nand U1429 (N_1429,In_148,N_1083);
xor U1430 (N_1430,In_2473,N_1112);
or U1431 (N_1431,N_973,N_277);
and U1432 (N_1432,N_1017,In_325);
and U1433 (N_1433,N_1073,N_67);
nor U1434 (N_1434,In_2232,In_94);
nor U1435 (N_1435,In_2173,N_1045);
nand U1436 (N_1436,In_105,N_974);
or U1437 (N_1437,In_648,N_158);
nor U1438 (N_1438,N_618,N_686);
and U1439 (N_1439,In_2130,In_395);
nor U1440 (N_1440,In_2098,In_140);
or U1441 (N_1441,N_912,N_1029);
nand U1442 (N_1442,N_1134,In_293);
nand U1443 (N_1443,N_1072,In_853);
or U1444 (N_1444,In_43,In_1532);
nand U1445 (N_1445,N_1046,N_13);
or U1446 (N_1446,N_1074,In_905);
and U1447 (N_1447,In_510,In_1792);
nand U1448 (N_1448,In_2014,N_1246);
nand U1449 (N_1449,In_735,N_1047);
and U1450 (N_1450,In_1417,In_895);
nor U1451 (N_1451,In_1830,In_871);
nand U1452 (N_1452,N_447,N_1139);
xor U1453 (N_1453,In_1311,In_672);
nor U1454 (N_1454,N_450,N_609);
nand U1455 (N_1455,N_18,In_1012);
xnor U1456 (N_1456,In_1841,In_519);
or U1457 (N_1457,N_1147,In_879);
nand U1458 (N_1458,In_1671,In_2179);
and U1459 (N_1459,N_1160,N_1190);
and U1460 (N_1460,N_307,N_991);
and U1461 (N_1461,N_1052,In_457);
nor U1462 (N_1462,In_1750,In_2345);
and U1463 (N_1463,In_2472,In_312);
xor U1464 (N_1464,In_2045,N_116);
xnor U1465 (N_1465,N_828,N_521);
nor U1466 (N_1466,In_1021,N_515);
or U1467 (N_1467,In_1333,In_1708);
and U1468 (N_1468,N_1006,N_394);
or U1469 (N_1469,In_1038,N_739);
or U1470 (N_1470,In_1630,N_1035);
or U1471 (N_1471,N_927,In_614);
or U1472 (N_1472,N_1055,In_285);
nand U1473 (N_1473,N_83,N_1248);
and U1474 (N_1474,In_18,N_764);
nand U1475 (N_1475,In_1706,N_694);
nand U1476 (N_1476,N_626,N_1203);
nor U1477 (N_1477,N_501,In_227);
and U1478 (N_1478,In_230,In_257);
or U1479 (N_1479,In_1535,N_1249);
xnor U1480 (N_1480,In_764,In_1897);
xor U1481 (N_1481,In_639,In_2454);
nor U1482 (N_1482,In_2207,N_766);
or U1483 (N_1483,In_505,In_1786);
and U1484 (N_1484,N_962,In_1210);
nand U1485 (N_1485,N_1123,In_2223);
and U1486 (N_1486,In_925,N_711);
or U1487 (N_1487,N_192,N_56);
nor U1488 (N_1488,In_2336,N_52);
nor U1489 (N_1489,N_558,N_1024);
and U1490 (N_1490,N_1110,In_2297);
and U1491 (N_1491,In_673,In_337);
xnor U1492 (N_1492,N_1026,In_2393);
nand U1493 (N_1493,In_365,N_1071);
nor U1494 (N_1494,N_869,N_363);
nand U1495 (N_1495,In_916,N_1009);
nor U1496 (N_1496,N_423,N_549);
or U1497 (N_1497,N_267,N_1179);
or U1498 (N_1498,In_1236,In_1990);
xnor U1499 (N_1499,N_875,In_2151);
xor U1500 (N_1500,In_2432,N_432);
or U1501 (N_1501,N_771,N_531);
or U1502 (N_1502,N_1476,In_1969);
and U1503 (N_1503,N_1241,In_1683);
or U1504 (N_1504,N_1418,N_1388);
xnor U1505 (N_1505,N_798,N_1451);
nor U1506 (N_1506,N_1490,In_1198);
nor U1507 (N_1507,N_1351,In_635);
nand U1508 (N_1508,In_1248,N_1438);
nor U1509 (N_1509,N_1283,N_687);
or U1510 (N_1510,N_288,N_1367);
or U1511 (N_1511,N_1416,N_1401);
nor U1512 (N_1512,In_183,N_284);
nor U1513 (N_1513,N_414,In_1221);
nor U1514 (N_1514,N_1497,N_1091);
nor U1515 (N_1515,N_1063,N_1376);
nor U1516 (N_1516,In_701,In_1659);
or U1517 (N_1517,N_602,N_1312);
nand U1518 (N_1518,N_1311,N_440);
nand U1519 (N_1519,N_901,N_1419);
xnor U1520 (N_1520,In_1554,In_1315);
nor U1521 (N_1521,In_1899,N_864);
xnor U1522 (N_1522,In_932,N_1033);
or U1523 (N_1523,N_1268,N_1194);
nand U1524 (N_1524,N_1420,In_2034);
xor U1525 (N_1525,In_2158,N_1483);
nor U1526 (N_1526,In_76,N_1323);
and U1527 (N_1527,In_928,In_1426);
nand U1528 (N_1528,N_1285,N_1040);
nor U1529 (N_1529,N_1089,N_1325);
and U1530 (N_1530,In_399,In_1799);
nor U1531 (N_1531,N_1079,N_442);
nand U1532 (N_1532,In_1813,N_1329);
nand U1533 (N_1533,N_1291,In_613);
and U1534 (N_1534,N_1349,N_1446);
nand U1535 (N_1535,N_1273,N_382);
xor U1536 (N_1536,In_481,N_1253);
nand U1537 (N_1537,N_1095,In_2082);
or U1538 (N_1538,N_1021,N_679);
or U1539 (N_1539,N_1409,N_1044);
nand U1540 (N_1540,In_1879,In_2304);
and U1541 (N_1541,N_1193,N_1441);
nand U1542 (N_1542,N_47,N_1413);
or U1543 (N_1543,N_1065,N_1061);
nand U1544 (N_1544,N_866,In_1121);
xor U1545 (N_1545,In_864,N_1062);
nor U1546 (N_1546,N_836,N_850);
or U1547 (N_1547,In_1081,N_1019);
nor U1548 (N_1548,N_1184,N_965);
nor U1549 (N_1549,N_1341,In_1940);
xor U1550 (N_1550,In_1964,In_880);
and U1551 (N_1551,N_858,N_1227);
and U1552 (N_1552,N_1290,N_741);
nor U1553 (N_1553,In_1963,In_2294);
xor U1554 (N_1554,N_1433,N_776);
and U1555 (N_1555,N_1302,N_1173);
or U1556 (N_1556,N_985,In_1619);
and U1557 (N_1557,N_452,N_1308);
nand U1558 (N_1558,N_1176,N_697);
and U1559 (N_1559,In_753,N_1058);
xor U1560 (N_1560,N_1229,N_1106);
xor U1561 (N_1561,N_893,N_1200);
nand U1562 (N_1562,In_569,N_949);
nor U1563 (N_1563,N_220,In_1357);
or U1564 (N_1564,N_1010,N_441);
nand U1565 (N_1565,N_479,In_1618);
nor U1566 (N_1566,N_257,N_1424);
and U1567 (N_1567,N_1472,N_1452);
or U1568 (N_1568,N_1333,N_1038);
xor U1569 (N_1569,N_102,N_915);
or U1570 (N_1570,N_1181,In_705);
xor U1571 (N_1571,N_1251,N_231);
nor U1572 (N_1572,N_1086,N_1426);
xor U1573 (N_1573,N_470,N_953);
xor U1574 (N_1574,In_107,In_2307);
and U1575 (N_1575,N_1491,In_275);
xnor U1576 (N_1576,N_333,In_943);
nand U1577 (N_1577,N_318,In_1156);
and U1578 (N_1578,N_1379,N_1450);
and U1579 (N_1579,In_1377,N_1318);
nand U1580 (N_1580,N_1131,N_167);
xnor U1581 (N_1581,N_1344,N_251);
xor U1582 (N_1582,In_2228,N_1165);
xnor U1583 (N_1583,N_94,N_1279);
xor U1584 (N_1584,N_886,N_900);
nand U1585 (N_1585,N_1166,N_1324);
nand U1586 (N_1586,N_224,N_1076);
and U1587 (N_1587,In_645,N_787);
xnor U1588 (N_1588,N_1328,N_1001);
and U1589 (N_1589,N_119,N_704);
xnor U1590 (N_1590,N_1008,N_666);
nand U1591 (N_1591,N_772,N_1396);
or U1592 (N_1592,N_1468,N_905);
and U1593 (N_1593,In_1034,N_583);
nor U1594 (N_1594,N_950,N_1295);
nand U1595 (N_1595,In_535,N_1070);
or U1596 (N_1596,N_540,In_525);
and U1597 (N_1597,In_1451,In_2346);
nand U1598 (N_1598,N_1210,In_170);
or U1599 (N_1599,In_2119,N_1048);
nand U1600 (N_1600,N_1358,N_1464);
nor U1601 (N_1601,In_87,In_877);
or U1602 (N_1602,In_967,N_975);
xnor U1603 (N_1603,N_1060,In_176);
xor U1604 (N_1604,N_1392,N_1207);
xnor U1605 (N_1605,In_134,N_581);
xor U1606 (N_1606,In_209,N_147);
nor U1607 (N_1607,N_29,N_884);
nand U1608 (N_1608,N_1202,N_1305);
and U1609 (N_1609,N_1386,In_2063);
nand U1610 (N_1610,In_2183,N_1057);
and U1611 (N_1611,In_418,N_1185);
and U1612 (N_1612,N_9,N_801);
nor U1613 (N_1613,N_1108,N_876);
nor U1614 (N_1614,N_877,N_1163);
or U1615 (N_1615,In_2103,N_438);
nand U1616 (N_1616,N_512,N_426);
and U1617 (N_1617,N_1039,N_849);
nand U1618 (N_1618,N_1025,N_1125);
xnor U1619 (N_1619,In_1188,N_1477);
or U1620 (N_1620,N_1014,N_1199);
xor U1621 (N_1621,N_584,N_387);
and U1622 (N_1622,N_585,N_1469);
xnor U1623 (N_1623,In_1050,N_1066);
and U1624 (N_1624,N_671,In_730);
or U1625 (N_1625,N_1064,In_1727);
nand U1626 (N_1626,N_335,N_1339);
xnor U1627 (N_1627,N_1069,In_1642);
xor U1628 (N_1628,N_1460,N_1197);
nor U1629 (N_1629,N_1360,N_1427);
xnor U1630 (N_1630,N_755,N_1050);
nor U1631 (N_1631,In_160,N_85);
or U1632 (N_1632,N_1042,N_1319);
xor U1633 (N_1633,N_1443,N_1320);
nand U1634 (N_1634,In_2474,N_535);
nand U1635 (N_1635,In_1163,N_1087);
or U1636 (N_1636,In_423,In_1185);
nor U1637 (N_1637,N_1275,N_1321);
xnor U1638 (N_1638,In_2149,N_868);
nand U1639 (N_1639,In_2043,N_1140);
nand U1640 (N_1640,N_1447,N_1489);
xor U1641 (N_1641,N_1380,In_314);
xor U1642 (N_1642,N_1437,In_319);
nand U1643 (N_1643,N_640,N_1431);
xnor U1644 (N_1644,In_1797,In_1654);
and U1645 (N_1645,In_374,N_966);
nor U1646 (N_1646,N_1458,N_1090);
nor U1647 (N_1647,N_1331,N_1082);
xor U1648 (N_1648,N_1394,In_2386);
nand U1649 (N_1649,In_1607,N_925);
nand U1650 (N_1650,N_255,N_64);
and U1651 (N_1651,In_2355,N_1359);
xnor U1652 (N_1652,N_880,N_1068);
and U1653 (N_1653,N_82,In_2300);
nand U1654 (N_1654,N_1264,N_1436);
or U1655 (N_1655,In_1265,N_627);
xor U1656 (N_1656,N_1067,N_1486);
nand U1657 (N_1657,N_1316,N_1309);
or U1658 (N_1658,N_1459,N_1205);
nor U1659 (N_1659,N_1170,N_1286);
and U1660 (N_1660,N_1422,N_938);
nand U1661 (N_1661,In_1243,N_1299);
nor U1662 (N_1662,In_2433,N_1189);
nor U1663 (N_1663,In_2487,In_2039);
or U1664 (N_1664,N_152,N_1094);
or U1665 (N_1665,N_79,N_518);
and U1666 (N_1666,N_344,N_1369);
xor U1667 (N_1667,N_904,N_1115);
nor U1668 (N_1668,N_1177,N_504);
nor U1669 (N_1669,N_1317,N_514);
nor U1670 (N_1670,N_1332,In_589);
nor U1671 (N_1671,N_1465,N_1393);
and U1672 (N_1672,In_1131,N_632);
nand U1673 (N_1673,In_2373,N_1211);
nor U1674 (N_1674,N_1093,N_690);
or U1675 (N_1675,N_308,In_1122);
xor U1676 (N_1676,In_1850,In_1767);
or U1677 (N_1677,N_508,N_1098);
or U1678 (N_1678,N_1355,N_834);
xor U1679 (N_1679,N_386,N_728);
nor U1680 (N_1680,N_465,N_1003);
and U1681 (N_1681,N_762,N_301);
xor U1682 (N_1682,In_634,In_1325);
or U1683 (N_1683,N_226,N_289);
xnor U1684 (N_1684,N_1399,N_1363);
or U1685 (N_1685,N_1256,In_132);
xnor U1686 (N_1686,N_1187,N_505);
or U1687 (N_1687,N_1265,In_831);
xor U1688 (N_1688,N_809,N_0);
or U1689 (N_1689,N_546,In_17);
and U1690 (N_1690,In_814,N_1276);
nand U1691 (N_1691,N_1154,N_1493);
and U1692 (N_1692,In_2385,In_889);
xnor U1693 (N_1693,N_821,In_898);
nor U1694 (N_1694,N_806,N_1053);
nand U1695 (N_1695,N_1148,In_355);
or U1696 (N_1696,N_1330,N_937);
or U1697 (N_1697,N_691,In_601);
nand U1698 (N_1698,N_60,N_908);
xor U1699 (N_1699,N_1298,In_41);
and U1700 (N_1700,N_320,N_768);
and U1701 (N_1701,In_989,In_1464);
xor U1702 (N_1702,In_2216,N_525);
xor U1703 (N_1703,N_853,N_1100);
or U1704 (N_1704,N_920,N_1336);
or U1705 (N_1705,In_2423,N_1129);
xor U1706 (N_1706,In_631,In_1471);
or U1707 (N_1707,N_599,In_786);
or U1708 (N_1708,N_1113,N_1281);
nand U1709 (N_1709,In_1657,N_200);
nand U1710 (N_1710,N_1111,N_802);
nand U1711 (N_1711,In_2321,N_1269);
or U1712 (N_1712,N_1307,N_506);
and U1713 (N_1713,In_1823,In_2133);
and U1714 (N_1714,N_1326,In_1600);
and U1715 (N_1715,N_995,In_765);
nand U1716 (N_1716,N_1384,N_1121);
or U1717 (N_1717,N_1397,In_1259);
nor U1718 (N_1718,N_1480,N_182);
and U1719 (N_1719,N_1410,N_1196);
nand U1720 (N_1720,N_1284,In_1376);
and U1721 (N_1721,N_1252,N_1186);
nor U1722 (N_1722,In_162,In_1442);
xnor U1723 (N_1723,N_961,In_2075);
or U1724 (N_1724,N_629,In_652);
nand U1725 (N_1725,N_1417,In_1820);
nor U1726 (N_1726,In_990,N_1250);
and U1727 (N_1727,N_421,In_1819);
or U1728 (N_1728,N_1288,N_669);
nand U1729 (N_1729,N_796,N_1385);
xnor U1730 (N_1730,In_1481,N_1470);
or U1731 (N_1731,In_1728,In_1582);
or U1732 (N_1732,N_887,N_133);
nor U1733 (N_1733,In_124,N_520);
or U1734 (N_1734,N_1406,N_1429);
nor U1735 (N_1735,N_239,In_1177);
or U1736 (N_1736,N_1212,N_781);
nor U1737 (N_1737,N_32,N_863);
xnor U1738 (N_1738,N_1375,N_1377);
xnor U1739 (N_1739,N_38,In_1172);
xor U1740 (N_1740,N_280,N_1056);
nor U1741 (N_1741,N_1408,N_408);
nand U1742 (N_1742,N_700,N_1345);
nand U1743 (N_1743,N_1293,In_685);
nand U1744 (N_1744,In_1318,N_1145);
nor U1745 (N_1745,N_614,N_1168);
nand U1746 (N_1746,In_1138,N_1244);
xnor U1747 (N_1747,N_1411,N_1220);
or U1748 (N_1748,N_1439,N_727);
or U1749 (N_1749,N_931,N_899);
nand U1750 (N_1750,N_1322,N_1662);
and U1751 (N_1751,N_957,N_1582);
xnor U1752 (N_1752,N_1280,In_2327);
nor U1753 (N_1753,In_772,N_1671);
nand U1754 (N_1754,N_1218,N_902);
and U1755 (N_1755,N_1520,N_1271);
nor U1756 (N_1756,In_265,In_1390);
and U1757 (N_1757,In_47,N_1368);
nor U1758 (N_1758,N_1018,N_1555);
and U1759 (N_1759,In_983,N_412);
or U1760 (N_1760,N_804,In_456);
and U1761 (N_1761,In_924,In_1572);
nand U1762 (N_1762,N_396,N_622);
xnor U1763 (N_1763,N_1736,In_1986);
nand U1764 (N_1764,In_48,N_1715);
and U1765 (N_1765,N_1402,In_1017);
nand U1766 (N_1766,In_2170,N_561);
xnor U1767 (N_1767,N_1613,In_2027);
or U1768 (N_1768,N_1737,In_658);
and U1769 (N_1769,N_1623,N_615);
nand U1770 (N_1770,N_1575,In_394);
or U1771 (N_1771,N_1407,N_1335);
or U1772 (N_1772,In_219,N_1652);
nor U1773 (N_1773,N_1563,N_1627);
nor U1774 (N_1774,N_1586,N_1557);
or U1775 (N_1775,In_151,In_591);
nor U1776 (N_1776,In_1612,N_542);
xnor U1777 (N_1777,N_1138,In_1625);
and U1778 (N_1778,N_1542,N_578);
or U1779 (N_1779,N_539,N_1658);
nor U1780 (N_1780,N_1104,N_1714);
xor U1781 (N_1781,N_1466,N_1716);
or U1782 (N_1782,N_1667,N_1703);
nor U1783 (N_1783,N_1618,In_1232);
and U1784 (N_1784,N_298,In_1088);
or U1785 (N_1785,N_1315,N_1434);
or U1786 (N_1786,In_2457,N_1721);
or U1787 (N_1787,N_1664,N_1301);
and U1788 (N_1788,N_1641,In_775);
nand U1789 (N_1789,In_1863,N_1303);
nand U1790 (N_1790,N_1538,In_1994);
nand U1791 (N_1791,N_1730,In_1347);
or U1792 (N_1792,N_1105,In_1987);
nor U1793 (N_1793,N_1292,N_1690);
and U1794 (N_1794,N_1266,N_1027);
or U1795 (N_1795,In_1049,N_1605);
nand U1796 (N_1796,In_1432,In_1474);
and U1797 (N_1797,N_1556,N_1741);
nor U1798 (N_1798,N_1372,N_1735);
nand U1799 (N_1799,In_750,N_1746);
nor U1800 (N_1800,N_1503,N_708);
nor U1801 (N_1801,N_890,N_1548);
nand U1802 (N_1802,N_1574,In_168);
nor U1803 (N_1803,N_872,N_1707);
nor U1804 (N_1804,N_1686,In_900);
nand U1805 (N_1805,N_1004,N_1601);
or U1806 (N_1806,In_768,N_1245);
nor U1807 (N_1807,N_1622,N_1373);
nand U1808 (N_1808,In_2196,N_1215);
nor U1809 (N_1809,In_295,N_1545);
or U1810 (N_1810,N_1708,In_1888);
or U1811 (N_1811,In_1045,In_180);
xor U1812 (N_1812,N_1041,N_524);
nor U1813 (N_1813,N_1569,N_1632);
nor U1814 (N_1814,In_1228,N_1588);
xnor U1815 (N_1815,N_1553,In_2250);
or U1816 (N_1816,N_1640,N_1531);
or U1817 (N_1817,N_832,In_142);
xnor U1818 (N_1818,N_1495,In_218);
or U1819 (N_1819,In_918,In_974);
nor U1820 (N_1820,In_602,N_1092);
or U1821 (N_1821,N_1231,N_1423);
and U1822 (N_1822,N_1442,N_1648);
nand U1823 (N_1823,N_1677,N_1156);
nand U1824 (N_1824,N_1565,N_1107);
nand U1825 (N_1825,In_1130,N_1258);
nor U1826 (N_1826,N_1513,N_136);
nand U1827 (N_1827,In_1066,In_292);
and U1828 (N_1828,N_1722,N_1725);
xnor U1829 (N_1829,N_1705,N_1454);
nand U1830 (N_1830,N_1161,N_1539);
xnor U1831 (N_1831,N_1572,N_1544);
nand U1832 (N_1832,N_1614,In_1332);
nor U1833 (N_1833,In_1251,N_1382);
nand U1834 (N_1834,N_1362,N_888);
nor U1835 (N_1835,N_1585,N_1547);
and U1836 (N_1836,N_1238,In_494);
and U1837 (N_1837,N_1011,In_116);
or U1838 (N_1838,In_1931,N_1383);
and U1839 (N_1839,N_693,In_1495);
and U1840 (N_1840,N_1612,N_1679);
nand U1841 (N_1841,N_401,N_1356);
and U1842 (N_1842,N_1566,N_1475);
nand U1843 (N_1843,N_1698,N_1590);
xnor U1844 (N_1844,N_1661,N_976);
nand U1845 (N_1845,N_1561,N_1164);
nor U1846 (N_1846,N_1235,In_1479);
nand U1847 (N_1847,N_1381,N_1691);
xor U1848 (N_1848,N_12,N_896);
or U1849 (N_1849,N_1711,N_1537);
xnor U1850 (N_1850,In_933,N_1484);
and U1851 (N_1851,N_1479,N_1720);
nor U1852 (N_1852,N_1467,In_2129);
nor U1853 (N_1853,N_648,N_1517);
or U1854 (N_1854,N_1519,N_1415);
nor U1855 (N_1855,In_1589,N_66);
nor U1856 (N_1856,N_603,N_1158);
nand U1857 (N_1857,N_1655,N_1278);
nor U1858 (N_1858,N_1499,N_1270);
and U1859 (N_1859,N_121,N_837);
xor U1860 (N_1860,N_1174,N_3);
or U1861 (N_1861,N_1444,N_1254);
or U1862 (N_1862,In_2325,In_1200);
nor U1863 (N_1863,N_312,N_770);
xnor U1864 (N_1864,In_2322,N_1099);
nand U1865 (N_1865,In_1279,N_1535);
nand U1866 (N_1866,N_1678,N_1260);
nor U1867 (N_1867,In_858,N_929);
nor U1868 (N_1868,N_1660,N_269);
or U1869 (N_1869,N_1602,N_859);
xor U1870 (N_1870,N_1682,In_144);
nand U1871 (N_1871,N_1366,N_1233);
xor U1872 (N_1872,N_1630,N_1554);
and U1873 (N_1873,In_1605,N_959);
nand U1874 (N_1874,N_1217,N_1103);
xnor U1875 (N_1875,N_1370,N_960);
and U1876 (N_1876,N_1259,N_1313);
or U1877 (N_1877,N_1603,N_1558);
xnor U1878 (N_1878,N_882,N_1665);
nand U1879 (N_1879,N_1435,N_1609);
xor U1880 (N_1880,In_1070,In_25);
and U1881 (N_1881,N_1456,N_805);
xnor U1882 (N_1882,N_1304,N_1471);
or U1883 (N_1883,N_353,N_1727);
nor U1884 (N_1884,N_1533,In_1514);
or U1885 (N_1885,N_1619,N_1621);
and U1886 (N_1886,N_528,N_873);
nand U1887 (N_1887,N_1414,In_1666);
nand U1888 (N_1888,N_1743,In_902);
and U1889 (N_1889,N_1559,N_15);
or U1890 (N_1890,N_1257,N_1593);
or U1891 (N_1891,N_1272,In_759);
xnor U1892 (N_1892,N_1680,N_841);
nor U1893 (N_1893,N_1732,N_1506);
xor U1894 (N_1894,N_1668,In_595);
nand U1895 (N_1895,N_1262,N_1550);
nand U1896 (N_1896,N_1631,N_1527);
nor U1897 (N_1897,N_1549,N_921);
xnor U1898 (N_1898,N_1371,N_1389);
or U1899 (N_1899,In_2159,N_1263);
xnor U1900 (N_1900,N_1002,In_1164);
nand U1901 (N_1901,N_374,N_1738);
or U1902 (N_1902,N_792,N_1546);
xnor U1903 (N_1903,In_1724,N_1051);
xnor U1904 (N_1904,N_860,N_1432);
xor U1905 (N_1905,N_1023,In_1776);
nor U1906 (N_1906,N_1717,N_735);
nand U1907 (N_1907,In_574,In_445);
or U1908 (N_1908,In_605,N_956);
nand U1909 (N_1909,In_1015,N_1643);
nor U1910 (N_1910,N_1532,In_1436);
or U1911 (N_1911,N_763,N_1724);
and U1912 (N_1912,N_443,N_1028);
xor U1913 (N_1913,In_2279,In_1527);
nor U1914 (N_1914,N_14,In_1525);
and U1915 (N_1915,In_1564,N_1338);
nor U1916 (N_1916,N_1525,N_1669);
or U1917 (N_1917,N_1144,N_610);
xor U1918 (N_1918,N_1731,N_1054);
or U1919 (N_1919,N_1342,N_537);
xor U1920 (N_1920,N_1155,N_1522);
nand U1921 (N_1921,N_1224,N_1214);
xor U1922 (N_1922,In_532,N_1718);
or U1923 (N_1923,In_2076,N_1400);
nand U1924 (N_1924,N_1749,N_1314);
and U1925 (N_1925,N_619,N_1182);
nand U1926 (N_1926,N_1560,In_2335);
and U1927 (N_1927,N_21,N_1608);
or U1928 (N_1928,In_504,N_1742);
nor U1929 (N_1929,N_1693,N_1504);
xnor U1930 (N_1930,N_1508,N_1530);
xnor U1931 (N_1931,N_1629,N_1702);
or U1932 (N_1932,N_997,N_1043);
xnor U1933 (N_1933,In_121,N_1310);
or U1934 (N_1934,N_1096,In_1784);
or U1935 (N_1935,N_1639,In_1561);
or U1936 (N_1936,In_178,N_1576);
nand U1937 (N_1937,N_1142,N_1353);
nand U1938 (N_1938,N_1412,N_579);
nor U1939 (N_1939,N_1567,N_1390);
nor U1940 (N_1940,N_1287,In_346);
or U1941 (N_1941,N_1694,N_1516);
nand U1942 (N_1942,N_1500,N_1541);
or U1943 (N_1943,In_2305,N_1455);
xnor U1944 (N_1944,N_1116,N_1403);
nand U1945 (N_1945,N_1620,In_1022);
nor U1946 (N_1946,In_1178,N_1511);
or U1947 (N_1947,In_1137,N_1536);
nand U1948 (N_1948,N_1697,N_343);
or U1949 (N_1949,In_931,N_910);
nand U1950 (N_1950,N_1606,N_580);
nor U1951 (N_1951,N_263,N_782);
and U1952 (N_1952,N_1463,N_1599);
nor U1953 (N_1953,N_1242,In_1594);
xnor U1954 (N_1954,N_665,N_1568);
xor U1955 (N_1955,N_1670,In_1522);
or U1956 (N_1956,N_725,N_1126);
nand U1957 (N_1957,N_1663,N_689);
nor U1958 (N_1958,N_1117,N_1178);
and U1959 (N_1959,N_1580,N_978);
nand U1960 (N_1960,In_2092,N_702);
nand U1961 (N_1961,N_1085,N_1604);
nand U1962 (N_1962,N_1745,N_1699);
or U1963 (N_1963,N_1352,N_1666);
nand U1964 (N_1964,N_1597,N_1482);
nand U1965 (N_1965,N_1591,N_1267);
or U1966 (N_1966,N_1729,N_1685);
nand U1967 (N_1967,N_1706,N_1357);
or U1968 (N_1968,N_391,N_1481);
or U1969 (N_1969,In_2395,In_1155);
nor U1970 (N_1970,N_1616,N_1228);
and U1971 (N_1971,In_1546,In_24);
and U1972 (N_1972,N_63,N_1696);
nand U1973 (N_1973,N_1642,In_2134);
nor U1974 (N_1974,N_820,In_57);
and U1975 (N_1975,N_1347,In_2383);
and U1976 (N_1976,In_850,N_1421);
and U1977 (N_1977,In_2081,N_1201);
or U1978 (N_1978,In_2095,N_418);
xor U1979 (N_1979,N_1296,N_1637);
nor U1980 (N_1980,N_1564,N_1523);
nand U1981 (N_1981,N_661,N_1650);
and U1982 (N_1982,N_425,N_1695);
xor U1983 (N_1983,N_1551,N_1261);
nor U1984 (N_1984,N_1404,N_332);
xor U1985 (N_1985,N_105,N_1700);
and U1986 (N_1986,N_1119,N_1587);
nand U1987 (N_1987,N_1128,N_1171);
nor U1988 (N_1988,N_1225,N_1628);
xnor U1989 (N_1989,N_1348,N_1692);
and U1990 (N_1990,In_126,N_1577);
nor U1991 (N_1991,In_675,N_1635);
and U1992 (N_1992,In_2154,N_151);
and U1993 (N_1993,N_1644,N_1710);
nor U1994 (N_1994,N_1221,In_2388);
nand U1995 (N_1995,N_1440,In_1975);
or U1996 (N_1996,In_1392,N_1688);
or U1997 (N_1997,N_1374,N_1649);
xnor U1998 (N_1998,N_1704,N_1405);
and U1999 (N_1999,In_11,N_1728);
xnor U2000 (N_2000,N_1498,N_1340);
xnor U2001 (N_2001,N_1759,N_1886);
nand U2002 (N_2002,N_992,N_1906);
and U2003 (N_2003,N_1768,N_1734);
or U2004 (N_2004,N_1733,N_1996);
nand U2005 (N_2005,N_1816,In_1307);
nor U2006 (N_2006,N_1988,N_1835);
nor U2007 (N_2007,N_1867,In_1381);
nor U2008 (N_2008,N_737,In_674);
or U2009 (N_2009,In_1298,N_1756);
xnor U2010 (N_2010,N_1877,N_1944);
nand U2011 (N_2011,N_1391,In_899);
xor U2012 (N_2012,N_1930,N_947);
nand U2013 (N_2013,N_1846,In_1747);
xor U2014 (N_2014,N_1956,N_1998);
nand U2015 (N_2015,N_1769,In_2470);
nor U2016 (N_2016,N_1935,N_1552);
xor U2017 (N_2017,N_1136,N_1780);
and U2018 (N_2018,N_1774,N_827);
xor U2019 (N_2019,In_1999,N_1750);
nand U2020 (N_2020,N_1921,N_1684);
and U2021 (N_2021,N_1878,N_1818);
nor U2022 (N_2022,N_1573,In_726);
nor U2023 (N_2023,In_2483,N_1817);
xnor U2024 (N_2024,N_830,N_1795);
or U2025 (N_2025,N_1236,N_1961);
xor U2026 (N_2026,N_1758,N_1989);
nor U2027 (N_2027,N_1681,N_1453);
or U2028 (N_2028,N_1457,N_1925);
xnor U2029 (N_2029,In_2113,N_1740);
nor U2030 (N_2030,N_1127,N_1943);
or U2031 (N_2031,N_1501,N_1723);
nand U2032 (N_2032,N_1751,In_1208);
nand U2033 (N_2033,N_1462,N_1689);
nand U2034 (N_2034,N_1350,N_1346);
and U2035 (N_2035,N_1739,N_1109);
nand U2036 (N_2036,N_1845,N_1888);
and U2037 (N_2037,N_1654,N_108);
nand U2038 (N_2038,N_1981,N_1870);
nand U2039 (N_2039,N_1924,N_1364);
xor U2040 (N_2040,N_1327,N_1625);
xor U2041 (N_2041,In_1389,In_1348);
and U2042 (N_2042,N_1918,N_1802);
nor U2043 (N_2043,N_1887,N_1809);
nor U2044 (N_2044,In_1883,N_1920);
or U2045 (N_2045,N_1861,N_1792);
or U2046 (N_2046,N_1529,In_912);
nor U2047 (N_2047,N_1826,N_1945);
nand U2048 (N_2048,N_1581,N_1297);
or U2049 (N_2049,N_1959,N_1847);
or U2050 (N_2050,N_1974,N_1873);
nor U2051 (N_2051,N_1940,N_1496);
or U2052 (N_2052,N_1584,In_411);
or U2053 (N_2053,N_1713,N_1687);
nor U2054 (N_2054,N_1815,N_1882);
nand U2055 (N_2055,N_1855,N_1928);
or U2056 (N_2056,N_1783,N_1844);
nor U2057 (N_2057,N_86,N_1800);
or U2058 (N_2058,N_1953,N_1274);
nor U2059 (N_2059,In_1143,N_1594);
xor U2060 (N_2060,N_1838,N_1907);
nor U2061 (N_2061,N_1822,N_1819);
and U2062 (N_2062,N_1827,N_1801);
xnor U2063 (N_2063,N_1595,N_818);
nand U2064 (N_2064,N_1823,N_1191);
xnor U2065 (N_2065,N_1796,N_1808);
nor U2066 (N_2066,N_1828,N_674);
nand U2067 (N_2067,N_1999,N_1980);
and U2068 (N_2068,N_1596,N_1675);
nand U2069 (N_2069,In_1327,N_1647);
xnor U2070 (N_2070,N_1534,N_1398);
nand U2071 (N_2071,N_1866,N_1987);
nand U2072 (N_2072,N_1934,N_1915);
xnor U2073 (N_2073,N_1954,N_1748);
xor U2074 (N_2074,N_1448,N_1230);
or U2075 (N_2075,N_1910,N_1791);
and U2076 (N_2076,N_1645,N_1488);
nor U2077 (N_2077,N_138,N_1430);
and U2078 (N_2078,N_1851,N_1785);
nor U2079 (N_2079,N_984,N_1395);
xor U2080 (N_2080,N_1101,N_1651);
nand U2081 (N_2081,N_1806,N_1150);
nand U2082 (N_2082,In_1135,N_673);
nor U2083 (N_2083,N_1387,N_1636);
nand U2084 (N_2084,N_1903,N_1653);
nand U2085 (N_2085,N_1803,N_1365);
or U2086 (N_2086,N_1948,N_1813);
nor U2087 (N_2087,N_1937,In_929);
or U2088 (N_2088,N_1676,N_760);
nor U2089 (N_2089,N_1965,N_1868);
xnor U2090 (N_2090,N_892,In_123);
nand U2091 (N_2091,N_1884,N_923);
nor U2092 (N_2092,N_1832,N_1294);
and U2093 (N_2093,N_1957,N_1805);
nand U2094 (N_2094,In_540,N_1247);
xnor U2095 (N_2095,In_1286,N_1841);
nand U2096 (N_2096,N_1219,N_1902);
nand U2097 (N_2097,N_1991,In_829);
xnor U2098 (N_2098,N_1782,N_1983);
xor U2099 (N_2099,In_985,N_1709);
or U2100 (N_2100,N_1521,N_1939);
nor U2101 (N_2101,N_1842,N_1000);
xnor U2102 (N_2102,N_703,N_1081);
or U2103 (N_2103,In_1013,N_1757);
or U2104 (N_2104,N_1747,N_1829);
and U2105 (N_2105,In_1294,N_1834);
xor U2106 (N_2106,N_1760,N_199);
xor U2107 (N_2107,N_1994,N_1840);
nor U2108 (N_2108,N_1839,N_1914);
xor U2109 (N_2109,N_989,N_1674);
or U2110 (N_2110,N_1787,N_1909);
xor U2111 (N_2111,N_1428,N_1899);
nor U2112 (N_2112,N_1626,In_840);
nor U2113 (N_2113,N_1277,N_1874);
nand U2114 (N_2114,N_1485,N_1646);
or U2115 (N_2115,In_2021,N_1820);
xnor U2116 (N_2116,In_972,N_1719);
nor U2117 (N_2117,N_1973,N_1853);
xor U2118 (N_2118,N_1509,In_1574);
nor U2119 (N_2119,N_1080,N_1872);
nor U2120 (N_2120,N_1922,N_1528);
xor U2121 (N_2121,N_1255,N_1833);
or U2122 (N_2122,N_1885,N_1814);
and U2123 (N_2123,N_1334,N_1967);
xnor U2124 (N_2124,N_1337,In_2177);
nand U2125 (N_2125,N_1512,N_70);
xor U2126 (N_2126,N_1510,N_1990);
nor U2127 (N_2127,N_1793,N_1672);
or U2128 (N_2128,N_1978,N_1797);
and U2129 (N_2129,N_1790,N_874);
and U2130 (N_2130,In_1852,N_1600);
nand U2131 (N_2131,N_1811,N_914);
xor U2132 (N_2132,N_1540,N_1962);
or U2133 (N_2133,In_2079,N_1180);
nand U2134 (N_2134,N_1610,N_1753);
nand U2135 (N_2135,N_1657,N_1863);
or U2136 (N_2136,N_1778,N_1972);
nand U2137 (N_2137,N_1240,N_1781);
xnor U2138 (N_2138,N_1615,N_803);
and U2139 (N_2139,N_1726,N_1570);
xnor U2140 (N_2140,N_1300,N_1779);
and U2141 (N_2141,In_1382,N_1964);
and U2142 (N_2142,N_1995,N_1857);
and U2143 (N_2143,In_1372,N_1761);
and U2144 (N_2144,N_1354,N_1836);
nor U2145 (N_2145,N_1869,N_1788);
and U2146 (N_2146,N_1938,In_2229);
or U2147 (N_2147,N_1982,N_1786);
and U2148 (N_2148,N_1908,N_1970);
nand U2149 (N_2149,N_1898,N_275);
xor U2150 (N_2150,In_1244,N_1889);
and U2151 (N_2151,N_1856,N_1963);
or U2152 (N_2152,N_1232,N_1583);
nand U2153 (N_2153,N_1449,N_1712);
nor U2154 (N_2154,N_1848,N_1871);
or U2155 (N_2155,N_415,N_1744);
nand U2156 (N_2156,N_1656,N_862);
or U2157 (N_2157,N_1473,N_1977);
nand U2158 (N_2158,N_1518,In_1816);
nand U2159 (N_2159,N_1879,N_1762);
xor U2160 (N_2160,N_1239,N_1986);
nor U2161 (N_2161,N_1897,N_195);
nand U2162 (N_2162,N_1425,N_1282);
or U2163 (N_2163,N_1775,N_1904);
nor U2164 (N_2164,In_1515,N_954);
and U2165 (N_2165,N_1772,N_1810);
and U2166 (N_2166,N_1985,N_1890);
nor U2167 (N_2167,N_1850,N_1950);
nor U2168 (N_2168,In_1878,N_1969);
or U2169 (N_2169,N_1936,In_1207);
xnor U2170 (N_2170,In_572,N_1752);
and U2171 (N_2171,N_1579,N_1952);
or U2172 (N_2172,N_932,N_1875);
or U2173 (N_2173,N_1824,N_1754);
nor U2174 (N_2174,N_1016,N_1932);
xor U2175 (N_2175,N_1865,N_1854);
or U2176 (N_2176,N_1755,N_1773);
and U2177 (N_2177,N_783,N_1378);
nand U2178 (N_2178,N_1234,N_1912);
xor U2179 (N_2179,In_651,N_1638);
nand U2180 (N_2180,N_178,N_1843);
nor U2181 (N_2181,N_1942,N_706);
xor U2182 (N_2182,N_1578,In_373);
and U2183 (N_2183,N_1931,N_1502);
and U2184 (N_2184,N_1895,N_1997);
or U2185 (N_2185,N_1976,N_1860);
xnor U2186 (N_2186,N_1852,In_1403);
or U2187 (N_2187,In_1183,N_1951);
or U2188 (N_2188,N_327,N_719);
and U2189 (N_2189,N_1767,N_1487);
nand U2190 (N_2190,N_1592,N_1917);
and U2191 (N_2191,N_800,N_1825);
xor U2192 (N_2192,N_1289,N_1900);
and U2193 (N_2193,N_1505,N_1633);
xnor U2194 (N_2194,N_1896,In_2272);
and U2195 (N_2195,N_1807,N_817);
or U2196 (N_2196,N_1831,N_1617);
or U2197 (N_2197,N_1911,N_1514);
nand U2198 (N_2198,N_1798,N_1905);
nor U2199 (N_2199,N_1993,N_1927);
or U2200 (N_2200,N_1763,In_367);
or U2201 (N_2201,N_1673,N_1492);
nor U2202 (N_2202,N_1916,N_1804);
and U2203 (N_2203,N_1923,N_1821);
xor U2204 (N_2204,N_1611,In_815);
nand U2205 (N_2205,In_2285,N_1876);
or U2206 (N_2206,N_1858,N_1919);
or U2207 (N_2207,N_1361,N_1933);
nor U2208 (N_2208,N_1949,N_1812);
nand U2209 (N_2209,N_1958,In_1946);
nor U2210 (N_2210,N_1901,N_1883);
and U2211 (N_2211,N_1975,N_1893);
xor U2212 (N_2212,N_680,N_1634);
xnor U2213 (N_2213,N_1894,N_1195);
and U2214 (N_2214,N_469,N_1794);
xor U2215 (N_2215,N_1789,N_1237);
and U2216 (N_2216,N_1598,N_1571);
nor U2217 (N_2217,N_1926,N_1929);
nor U2218 (N_2218,N_1445,N_1955);
and U2219 (N_2219,N_1859,In_565);
or U2220 (N_2220,N_1971,N_1984);
and U2221 (N_2221,N_1837,N_1765);
nor U2222 (N_2222,N_1777,N_1764);
xor U2223 (N_2223,N_1880,In_666);
nand U2224 (N_2224,N_898,N_1799);
xor U2225 (N_2225,N_1960,N_1562);
and U2226 (N_2226,N_1526,N_202);
and U2227 (N_2227,N_1515,N_1892);
xor U2228 (N_2228,N_1891,In_882);
and U2229 (N_2229,N_1589,N_840);
nand U2230 (N_2230,N_1864,N_1776);
nand U2231 (N_2231,N_1941,N_1624);
xnor U2232 (N_2232,N_1966,N_1478);
xor U2233 (N_2233,In_703,N_1659);
or U2234 (N_2234,N_1306,N_1343);
or U2235 (N_2235,N_1946,N_1507);
nor U2236 (N_2236,N_1683,N_1543);
and U2237 (N_2237,N_1524,N_1701);
and U2238 (N_2238,N_598,N_1968);
xnor U2239 (N_2239,N_1913,N_1881);
nor U2240 (N_2240,N_1830,N_1784);
and U2241 (N_2241,N_1771,N_1474);
and U2242 (N_2242,N_1947,N_913);
or U2243 (N_2243,N_35,In_2444);
or U2244 (N_2244,N_1992,N_1494);
nand U2245 (N_2245,N_1607,N_1461);
or U2246 (N_2246,N_1862,N_1059);
or U2247 (N_2247,N_964,N_523);
nor U2248 (N_2248,N_1766,N_1849);
nand U2249 (N_2249,N_1979,N_1770);
nor U2250 (N_2250,N_2116,N_2073);
nor U2251 (N_2251,N_2172,N_2204);
nor U2252 (N_2252,N_2156,N_2144);
or U2253 (N_2253,N_2131,N_2135);
nand U2254 (N_2254,N_2235,N_2036);
xor U2255 (N_2255,N_2142,N_2200);
or U2256 (N_2256,N_2115,N_2063);
or U2257 (N_2257,N_2234,N_2082);
and U2258 (N_2258,N_2193,N_2205);
nor U2259 (N_2259,N_2199,N_2242);
and U2260 (N_2260,N_2168,N_2220);
and U2261 (N_2261,N_2202,N_2231);
or U2262 (N_2262,N_2025,N_2097);
xor U2263 (N_2263,N_2146,N_2019);
xor U2264 (N_2264,N_2008,N_2004);
or U2265 (N_2265,N_2195,N_2171);
and U2266 (N_2266,N_2068,N_2108);
nor U2267 (N_2267,N_2033,N_2112);
nand U2268 (N_2268,N_2027,N_2048);
nand U2269 (N_2269,N_2192,N_2028);
nor U2270 (N_2270,N_2100,N_2133);
nor U2271 (N_2271,N_2159,N_2088);
nor U2272 (N_2272,N_2249,N_2130);
or U2273 (N_2273,N_2218,N_2143);
and U2274 (N_2274,N_2087,N_2189);
and U2275 (N_2275,N_2011,N_2080);
xnor U2276 (N_2276,N_2103,N_2085);
and U2277 (N_2277,N_2024,N_2094);
or U2278 (N_2278,N_2107,N_2099);
nor U2279 (N_2279,N_2118,N_2150);
nor U2280 (N_2280,N_2122,N_2084);
and U2281 (N_2281,N_2244,N_2182);
nand U2282 (N_2282,N_2240,N_2003);
nor U2283 (N_2283,N_2006,N_2104);
xnor U2284 (N_2284,N_2232,N_2213);
and U2285 (N_2285,N_2002,N_2201);
nor U2286 (N_2286,N_2058,N_2092);
nor U2287 (N_2287,N_2055,N_2208);
xor U2288 (N_2288,N_2059,N_2022);
or U2289 (N_2289,N_2061,N_2226);
and U2290 (N_2290,N_2225,N_2123);
nor U2291 (N_2291,N_2209,N_2247);
and U2292 (N_2292,N_2186,N_2134);
or U2293 (N_2293,N_2190,N_2187);
nor U2294 (N_2294,N_2158,N_2132);
nand U2295 (N_2295,N_2045,N_2046);
or U2296 (N_2296,N_2090,N_2236);
nand U2297 (N_2297,N_2009,N_2096);
or U2298 (N_2298,N_2203,N_2042);
xnor U2299 (N_2299,N_2185,N_2018);
or U2300 (N_2300,N_2161,N_2160);
or U2301 (N_2301,N_2173,N_2117);
nand U2302 (N_2302,N_2215,N_2217);
xnor U2303 (N_2303,N_2044,N_2238);
nor U2304 (N_2304,N_2015,N_2081);
nor U2305 (N_2305,N_2020,N_2248);
nor U2306 (N_2306,N_2219,N_2050);
or U2307 (N_2307,N_2149,N_2105);
or U2308 (N_2308,N_2210,N_2109);
or U2309 (N_2309,N_2040,N_2223);
nand U2310 (N_2310,N_2167,N_2141);
or U2311 (N_2311,N_2089,N_2222);
nand U2312 (N_2312,N_2120,N_2023);
and U2313 (N_2313,N_2239,N_2164);
or U2314 (N_2314,N_2121,N_2165);
xnor U2315 (N_2315,N_2211,N_2031);
xnor U2316 (N_2316,N_2153,N_2066);
nor U2317 (N_2317,N_2060,N_2154);
nand U2318 (N_2318,N_2111,N_2157);
or U2319 (N_2319,N_2224,N_2162);
xnor U2320 (N_2320,N_2245,N_2075);
nand U2321 (N_2321,N_2214,N_2098);
xor U2322 (N_2322,N_2072,N_2083);
and U2323 (N_2323,N_2183,N_2125);
and U2324 (N_2324,N_2110,N_2145);
or U2325 (N_2325,N_2140,N_2169);
xor U2326 (N_2326,N_2188,N_2126);
nor U2327 (N_2327,N_2039,N_2207);
or U2328 (N_2328,N_2101,N_2032);
nand U2329 (N_2329,N_2102,N_2013);
xnor U2330 (N_2330,N_2137,N_2037);
nor U2331 (N_2331,N_2127,N_2166);
nand U2332 (N_2332,N_2012,N_2014);
xor U2333 (N_2333,N_2197,N_2049);
nand U2334 (N_2334,N_2181,N_2147);
and U2335 (N_2335,N_2091,N_2206);
nor U2336 (N_2336,N_2128,N_2151);
and U2337 (N_2337,N_2148,N_2001);
nor U2338 (N_2338,N_2095,N_2228);
xnor U2339 (N_2339,N_2191,N_2106);
and U2340 (N_2340,N_2176,N_2079);
or U2341 (N_2341,N_2233,N_2065);
and U2342 (N_2342,N_2051,N_2180);
xor U2343 (N_2343,N_2227,N_2124);
nand U2344 (N_2344,N_2067,N_2071);
or U2345 (N_2345,N_2170,N_2139);
xor U2346 (N_2346,N_2005,N_2056);
nand U2347 (N_2347,N_2212,N_2076);
nand U2348 (N_2348,N_2177,N_2074);
nand U2349 (N_2349,N_2155,N_2163);
xnor U2350 (N_2350,N_2041,N_2174);
xor U2351 (N_2351,N_2119,N_2216);
or U2352 (N_2352,N_2047,N_2000);
or U2353 (N_2353,N_2038,N_2198);
nand U2354 (N_2354,N_2007,N_2069);
xnor U2355 (N_2355,N_2184,N_2054);
nor U2356 (N_2356,N_2179,N_2017);
and U2357 (N_2357,N_2077,N_2070);
nor U2358 (N_2358,N_2064,N_2196);
nor U2359 (N_2359,N_2016,N_2021);
nor U2360 (N_2360,N_2152,N_2114);
nand U2361 (N_2361,N_2026,N_2053);
xor U2362 (N_2362,N_2052,N_2243);
nor U2363 (N_2363,N_2230,N_2062);
or U2364 (N_2364,N_2138,N_2194);
nor U2365 (N_2365,N_2129,N_2078);
xnor U2366 (N_2366,N_2246,N_2241);
xor U2367 (N_2367,N_2229,N_2221);
nor U2368 (N_2368,N_2237,N_2030);
or U2369 (N_2369,N_2136,N_2113);
or U2370 (N_2370,N_2093,N_2057);
and U2371 (N_2371,N_2035,N_2175);
nor U2372 (N_2372,N_2178,N_2029);
nor U2373 (N_2373,N_2034,N_2086);
nor U2374 (N_2374,N_2043,N_2010);
nand U2375 (N_2375,N_2083,N_2194);
nand U2376 (N_2376,N_2111,N_2179);
and U2377 (N_2377,N_2035,N_2214);
and U2378 (N_2378,N_2243,N_2211);
nor U2379 (N_2379,N_2093,N_2037);
and U2380 (N_2380,N_2085,N_2157);
nand U2381 (N_2381,N_2203,N_2075);
nor U2382 (N_2382,N_2037,N_2117);
nor U2383 (N_2383,N_2095,N_2009);
and U2384 (N_2384,N_2100,N_2192);
or U2385 (N_2385,N_2239,N_2094);
xor U2386 (N_2386,N_2145,N_2083);
nor U2387 (N_2387,N_2148,N_2034);
xnor U2388 (N_2388,N_2000,N_2094);
and U2389 (N_2389,N_2143,N_2028);
nand U2390 (N_2390,N_2125,N_2029);
nand U2391 (N_2391,N_2019,N_2203);
nand U2392 (N_2392,N_2115,N_2137);
or U2393 (N_2393,N_2197,N_2176);
or U2394 (N_2394,N_2169,N_2026);
nand U2395 (N_2395,N_2085,N_2008);
nand U2396 (N_2396,N_2053,N_2205);
and U2397 (N_2397,N_2205,N_2119);
xor U2398 (N_2398,N_2092,N_2118);
and U2399 (N_2399,N_2005,N_2203);
xnor U2400 (N_2400,N_2074,N_2117);
nand U2401 (N_2401,N_2090,N_2175);
nor U2402 (N_2402,N_2150,N_2139);
nor U2403 (N_2403,N_2163,N_2209);
and U2404 (N_2404,N_2046,N_2041);
and U2405 (N_2405,N_2188,N_2132);
or U2406 (N_2406,N_2043,N_2210);
or U2407 (N_2407,N_2005,N_2237);
nor U2408 (N_2408,N_2044,N_2220);
or U2409 (N_2409,N_2183,N_2122);
and U2410 (N_2410,N_2231,N_2045);
or U2411 (N_2411,N_2146,N_2158);
and U2412 (N_2412,N_2084,N_2138);
xnor U2413 (N_2413,N_2146,N_2094);
or U2414 (N_2414,N_2209,N_2169);
or U2415 (N_2415,N_2132,N_2242);
nand U2416 (N_2416,N_2039,N_2120);
nor U2417 (N_2417,N_2128,N_2131);
nand U2418 (N_2418,N_2015,N_2068);
nand U2419 (N_2419,N_2233,N_2012);
nand U2420 (N_2420,N_2108,N_2228);
nor U2421 (N_2421,N_2074,N_2038);
and U2422 (N_2422,N_2180,N_2061);
or U2423 (N_2423,N_2138,N_2007);
nor U2424 (N_2424,N_2089,N_2142);
xor U2425 (N_2425,N_2240,N_2150);
and U2426 (N_2426,N_2151,N_2019);
and U2427 (N_2427,N_2230,N_2216);
or U2428 (N_2428,N_2144,N_2137);
nand U2429 (N_2429,N_2124,N_2051);
nor U2430 (N_2430,N_2138,N_2160);
nor U2431 (N_2431,N_2233,N_2114);
xor U2432 (N_2432,N_2138,N_2001);
nor U2433 (N_2433,N_2241,N_2025);
nor U2434 (N_2434,N_2165,N_2053);
and U2435 (N_2435,N_2051,N_2216);
nand U2436 (N_2436,N_2082,N_2165);
or U2437 (N_2437,N_2036,N_2155);
or U2438 (N_2438,N_2084,N_2153);
nor U2439 (N_2439,N_2203,N_2028);
nor U2440 (N_2440,N_2171,N_2177);
nor U2441 (N_2441,N_2103,N_2078);
xnor U2442 (N_2442,N_2007,N_2223);
nor U2443 (N_2443,N_2219,N_2212);
xnor U2444 (N_2444,N_2084,N_2121);
xor U2445 (N_2445,N_2030,N_2050);
and U2446 (N_2446,N_2008,N_2121);
nor U2447 (N_2447,N_2146,N_2047);
xnor U2448 (N_2448,N_2202,N_2065);
xor U2449 (N_2449,N_2073,N_2042);
or U2450 (N_2450,N_2132,N_2061);
nand U2451 (N_2451,N_2144,N_2073);
and U2452 (N_2452,N_2068,N_2209);
and U2453 (N_2453,N_2145,N_2241);
nand U2454 (N_2454,N_2161,N_2158);
xnor U2455 (N_2455,N_2116,N_2244);
xnor U2456 (N_2456,N_2004,N_2014);
nor U2457 (N_2457,N_2187,N_2095);
nand U2458 (N_2458,N_2093,N_2205);
nor U2459 (N_2459,N_2108,N_2002);
or U2460 (N_2460,N_2010,N_2140);
and U2461 (N_2461,N_2033,N_2049);
or U2462 (N_2462,N_2193,N_2110);
or U2463 (N_2463,N_2054,N_2135);
nand U2464 (N_2464,N_2041,N_2176);
or U2465 (N_2465,N_2015,N_2108);
or U2466 (N_2466,N_2045,N_2024);
and U2467 (N_2467,N_2119,N_2244);
xor U2468 (N_2468,N_2038,N_2205);
or U2469 (N_2469,N_2046,N_2022);
xnor U2470 (N_2470,N_2205,N_2076);
nor U2471 (N_2471,N_2202,N_2093);
nor U2472 (N_2472,N_2069,N_2222);
nor U2473 (N_2473,N_2160,N_2066);
nand U2474 (N_2474,N_2037,N_2219);
nand U2475 (N_2475,N_2007,N_2056);
or U2476 (N_2476,N_2102,N_2197);
or U2477 (N_2477,N_2026,N_2156);
or U2478 (N_2478,N_2008,N_2088);
nor U2479 (N_2479,N_2229,N_2095);
nand U2480 (N_2480,N_2174,N_2226);
nor U2481 (N_2481,N_2002,N_2022);
or U2482 (N_2482,N_2099,N_2084);
nand U2483 (N_2483,N_2000,N_2174);
or U2484 (N_2484,N_2091,N_2221);
or U2485 (N_2485,N_2219,N_2242);
xnor U2486 (N_2486,N_2000,N_2126);
or U2487 (N_2487,N_2175,N_2131);
or U2488 (N_2488,N_2160,N_2050);
nor U2489 (N_2489,N_2146,N_2218);
xnor U2490 (N_2490,N_2143,N_2153);
nor U2491 (N_2491,N_2196,N_2227);
or U2492 (N_2492,N_2011,N_2177);
nand U2493 (N_2493,N_2038,N_2214);
xnor U2494 (N_2494,N_2174,N_2236);
nand U2495 (N_2495,N_2198,N_2016);
nor U2496 (N_2496,N_2041,N_2137);
xor U2497 (N_2497,N_2088,N_2209);
nor U2498 (N_2498,N_2125,N_2015);
and U2499 (N_2499,N_2111,N_2012);
xor U2500 (N_2500,N_2308,N_2404);
and U2501 (N_2501,N_2412,N_2419);
nor U2502 (N_2502,N_2341,N_2487);
nand U2503 (N_2503,N_2336,N_2290);
and U2504 (N_2504,N_2455,N_2461);
nand U2505 (N_2505,N_2267,N_2431);
and U2506 (N_2506,N_2390,N_2491);
and U2507 (N_2507,N_2459,N_2470);
or U2508 (N_2508,N_2330,N_2298);
and U2509 (N_2509,N_2362,N_2281);
nand U2510 (N_2510,N_2474,N_2493);
nor U2511 (N_2511,N_2306,N_2424);
nand U2512 (N_2512,N_2282,N_2492);
or U2513 (N_2513,N_2383,N_2477);
xnor U2514 (N_2514,N_2460,N_2415);
nand U2515 (N_2515,N_2387,N_2452);
and U2516 (N_2516,N_2269,N_2483);
xor U2517 (N_2517,N_2399,N_2413);
or U2518 (N_2518,N_2319,N_2328);
nand U2519 (N_2519,N_2378,N_2488);
xnor U2520 (N_2520,N_2454,N_2498);
nand U2521 (N_2521,N_2349,N_2266);
and U2522 (N_2522,N_2482,N_2253);
xnor U2523 (N_2523,N_2379,N_2329);
nor U2524 (N_2524,N_2311,N_2406);
nand U2525 (N_2525,N_2261,N_2439);
nor U2526 (N_2526,N_2370,N_2258);
or U2527 (N_2527,N_2497,N_2352);
and U2528 (N_2528,N_2393,N_2361);
nand U2529 (N_2529,N_2337,N_2490);
or U2530 (N_2530,N_2275,N_2360);
and U2531 (N_2531,N_2421,N_2475);
nand U2532 (N_2532,N_2458,N_2473);
nor U2533 (N_2533,N_2438,N_2429);
xor U2534 (N_2534,N_2320,N_2372);
or U2535 (N_2535,N_2323,N_2397);
nor U2536 (N_2536,N_2277,N_2448);
xor U2537 (N_2537,N_2398,N_2440);
xnor U2538 (N_2538,N_2268,N_2289);
xor U2539 (N_2539,N_2292,N_2381);
and U2540 (N_2540,N_2433,N_2254);
or U2541 (N_2541,N_2446,N_2280);
nor U2542 (N_2542,N_2380,N_2449);
or U2543 (N_2543,N_2297,N_2316);
or U2544 (N_2544,N_2436,N_2392);
and U2545 (N_2545,N_2420,N_2351);
nand U2546 (N_2546,N_2367,N_2462);
nor U2547 (N_2547,N_2312,N_2386);
or U2548 (N_2548,N_2284,N_2447);
nand U2549 (N_2549,N_2400,N_2407);
xnor U2550 (N_2550,N_2279,N_2340);
nand U2551 (N_2551,N_2366,N_2444);
xnor U2552 (N_2552,N_2355,N_2434);
xor U2553 (N_2553,N_2276,N_2423);
or U2554 (N_2554,N_2302,N_2485);
nor U2555 (N_2555,N_2287,N_2356);
or U2556 (N_2556,N_2382,N_2403);
xor U2557 (N_2557,N_2283,N_2295);
or U2558 (N_2558,N_2377,N_2263);
xor U2559 (N_2559,N_2375,N_2405);
nand U2560 (N_2560,N_2499,N_2293);
nand U2561 (N_2561,N_2469,N_2478);
nand U2562 (N_2562,N_2343,N_2486);
or U2563 (N_2563,N_2384,N_2481);
nand U2564 (N_2564,N_2385,N_2451);
or U2565 (N_2565,N_2318,N_2411);
and U2566 (N_2566,N_2408,N_2476);
and U2567 (N_2567,N_2395,N_2394);
xor U2568 (N_2568,N_2358,N_2315);
and U2569 (N_2569,N_2354,N_2494);
xor U2570 (N_2570,N_2346,N_2489);
or U2571 (N_2571,N_2296,N_2314);
and U2572 (N_2572,N_2286,N_2442);
nand U2573 (N_2573,N_2456,N_2332);
nor U2574 (N_2574,N_2285,N_2317);
nand U2575 (N_2575,N_2402,N_2274);
nand U2576 (N_2576,N_2305,N_2270);
and U2577 (N_2577,N_2376,N_2472);
nor U2578 (N_2578,N_2432,N_2288);
nor U2579 (N_2579,N_2425,N_2414);
or U2580 (N_2580,N_2291,N_2333);
nor U2581 (N_2581,N_2278,N_2310);
nor U2582 (N_2582,N_2327,N_2445);
xor U2583 (N_2583,N_2331,N_2353);
and U2584 (N_2584,N_2322,N_2410);
xnor U2585 (N_2585,N_2260,N_2338);
xor U2586 (N_2586,N_2401,N_2495);
xnor U2587 (N_2587,N_2363,N_2437);
and U2588 (N_2588,N_2365,N_2443);
xnor U2589 (N_2589,N_2304,N_2427);
nor U2590 (N_2590,N_2441,N_2435);
and U2591 (N_2591,N_2391,N_2422);
nand U2592 (N_2592,N_2428,N_2465);
xor U2593 (N_2593,N_2373,N_2453);
nand U2594 (N_2594,N_2457,N_2344);
nor U2595 (N_2595,N_2264,N_2303);
or U2596 (N_2596,N_2479,N_2388);
and U2597 (N_2597,N_2307,N_2321);
or U2598 (N_2598,N_2300,N_2309);
nor U2599 (N_2599,N_2409,N_2335);
or U2600 (N_2600,N_2334,N_2357);
or U2601 (N_2601,N_2345,N_2259);
nor U2602 (N_2602,N_2313,N_2466);
and U2603 (N_2603,N_2426,N_2496);
or U2604 (N_2604,N_2262,N_2271);
or U2605 (N_2605,N_2299,N_2250);
or U2606 (N_2606,N_2471,N_2256);
nand U2607 (N_2607,N_2430,N_2467);
and U2608 (N_2608,N_2364,N_2416);
or U2609 (N_2609,N_2468,N_2294);
nand U2610 (N_2610,N_2369,N_2368);
xor U2611 (N_2611,N_2464,N_2348);
xor U2612 (N_2612,N_2484,N_2339);
xor U2613 (N_2613,N_2418,N_2347);
and U2614 (N_2614,N_2301,N_2324);
nor U2615 (N_2615,N_2396,N_2251);
nor U2616 (N_2616,N_2359,N_2350);
nand U2617 (N_2617,N_2389,N_2255);
and U2618 (N_2618,N_2265,N_2326);
or U2619 (N_2619,N_2374,N_2371);
xor U2620 (N_2620,N_2450,N_2257);
nand U2621 (N_2621,N_2252,N_2273);
and U2622 (N_2622,N_2417,N_2325);
nand U2623 (N_2623,N_2463,N_2272);
nand U2624 (N_2624,N_2480,N_2342);
nor U2625 (N_2625,N_2465,N_2299);
and U2626 (N_2626,N_2480,N_2493);
xnor U2627 (N_2627,N_2349,N_2466);
and U2628 (N_2628,N_2488,N_2465);
or U2629 (N_2629,N_2313,N_2292);
xor U2630 (N_2630,N_2250,N_2385);
nand U2631 (N_2631,N_2273,N_2412);
nor U2632 (N_2632,N_2299,N_2348);
or U2633 (N_2633,N_2259,N_2304);
xor U2634 (N_2634,N_2387,N_2402);
and U2635 (N_2635,N_2439,N_2473);
nand U2636 (N_2636,N_2462,N_2317);
nand U2637 (N_2637,N_2316,N_2298);
nand U2638 (N_2638,N_2481,N_2310);
or U2639 (N_2639,N_2379,N_2437);
or U2640 (N_2640,N_2420,N_2418);
nor U2641 (N_2641,N_2438,N_2405);
nor U2642 (N_2642,N_2404,N_2487);
nor U2643 (N_2643,N_2437,N_2265);
xnor U2644 (N_2644,N_2443,N_2271);
nand U2645 (N_2645,N_2459,N_2484);
xor U2646 (N_2646,N_2290,N_2425);
nand U2647 (N_2647,N_2358,N_2263);
nand U2648 (N_2648,N_2314,N_2294);
xor U2649 (N_2649,N_2422,N_2462);
nor U2650 (N_2650,N_2310,N_2384);
nor U2651 (N_2651,N_2288,N_2485);
xor U2652 (N_2652,N_2419,N_2398);
nor U2653 (N_2653,N_2434,N_2255);
or U2654 (N_2654,N_2395,N_2377);
or U2655 (N_2655,N_2492,N_2258);
xnor U2656 (N_2656,N_2257,N_2278);
xor U2657 (N_2657,N_2371,N_2464);
and U2658 (N_2658,N_2446,N_2487);
xor U2659 (N_2659,N_2329,N_2335);
nand U2660 (N_2660,N_2316,N_2347);
or U2661 (N_2661,N_2326,N_2266);
nand U2662 (N_2662,N_2284,N_2478);
and U2663 (N_2663,N_2302,N_2321);
xor U2664 (N_2664,N_2410,N_2253);
xor U2665 (N_2665,N_2250,N_2262);
and U2666 (N_2666,N_2444,N_2496);
xor U2667 (N_2667,N_2328,N_2489);
nand U2668 (N_2668,N_2455,N_2305);
nor U2669 (N_2669,N_2473,N_2495);
nor U2670 (N_2670,N_2294,N_2414);
nor U2671 (N_2671,N_2366,N_2395);
nor U2672 (N_2672,N_2491,N_2471);
and U2673 (N_2673,N_2382,N_2321);
or U2674 (N_2674,N_2420,N_2262);
xnor U2675 (N_2675,N_2263,N_2461);
nand U2676 (N_2676,N_2426,N_2381);
nand U2677 (N_2677,N_2403,N_2277);
nor U2678 (N_2678,N_2418,N_2488);
nor U2679 (N_2679,N_2338,N_2393);
and U2680 (N_2680,N_2401,N_2346);
xnor U2681 (N_2681,N_2333,N_2284);
xor U2682 (N_2682,N_2371,N_2352);
nand U2683 (N_2683,N_2264,N_2387);
nand U2684 (N_2684,N_2384,N_2277);
xnor U2685 (N_2685,N_2479,N_2449);
nor U2686 (N_2686,N_2436,N_2472);
nand U2687 (N_2687,N_2471,N_2375);
and U2688 (N_2688,N_2365,N_2258);
nor U2689 (N_2689,N_2341,N_2397);
or U2690 (N_2690,N_2271,N_2384);
xnor U2691 (N_2691,N_2268,N_2312);
or U2692 (N_2692,N_2457,N_2328);
and U2693 (N_2693,N_2314,N_2465);
nor U2694 (N_2694,N_2482,N_2471);
nand U2695 (N_2695,N_2483,N_2259);
xnor U2696 (N_2696,N_2457,N_2373);
and U2697 (N_2697,N_2340,N_2388);
nor U2698 (N_2698,N_2325,N_2361);
nor U2699 (N_2699,N_2461,N_2311);
xnor U2700 (N_2700,N_2440,N_2361);
nor U2701 (N_2701,N_2423,N_2452);
nor U2702 (N_2702,N_2254,N_2460);
and U2703 (N_2703,N_2318,N_2368);
xor U2704 (N_2704,N_2463,N_2424);
and U2705 (N_2705,N_2303,N_2353);
xor U2706 (N_2706,N_2400,N_2327);
nor U2707 (N_2707,N_2463,N_2343);
and U2708 (N_2708,N_2286,N_2445);
and U2709 (N_2709,N_2345,N_2415);
nand U2710 (N_2710,N_2478,N_2401);
and U2711 (N_2711,N_2464,N_2490);
nor U2712 (N_2712,N_2464,N_2406);
nor U2713 (N_2713,N_2426,N_2497);
and U2714 (N_2714,N_2312,N_2445);
nand U2715 (N_2715,N_2251,N_2485);
xor U2716 (N_2716,N_2283,N_2365);
or U2717 (N_2717,N_2268,N_2498);
nand U2718 (N_2718,N_2416,N_2343);
or U2719 (N_2719,N_2399,N_2250);
or U2720 (N_2720,N_2428,N_2367);
nand U2721 (N_2721,N_2304,N_2464);
nand U2722 (N_2722,N_2361,N_2457);
nor U2723 (N_2723,N_2366,N_2293);
nor U2724 (N_2724,N_2359,N_2411);
and U2725 (N_2725,N_2391,N_2360);
nand U2726 (N_2726,N_2303,N_2400);
and U2727 (N_2727,N_2442,N_2423);
nand U2728 (N_2728,N_2371,N_2392);
nor U2729 (N_2729,N_2305,N_2265);
and U2730 (N_2730,N_2294,N_2293);
nand U2731 (N_2731,N_2424,N_2358);
and U2732 (N_2732,N_2266,N_2319);
nor U2733 (N_2733,N_2353,N_2397);
or U2734 (N_2734,N_2362,N_2443);
xnor U2735 (N_2735,N_2471,N_2326);
xor U2736 (N_2736,N_2475,N_2283);
and U2737 (N_2737,N_2431,N_2359);
and U2738 (N_2738,N_2429,N_2309);
and U2739 (N_2739,N_2310,N_2275);
xnor U2740 (N_2740,N_2349,N_2315);
nand U2741 (N_2741,N_2391,N_2264);
nand U2742 (N_2742,N_2383,N_2440);
and U2743 (N_2743,N_2256,N_2291);
or U2744 (N_2744,N_2352,N_2466);
and U2745 (N_2745,N_2434,N_2400);
and U2746 (N_2746,N_2304,N_2401);
nor U2747 (N_2747,N_2430,N_2343);
or U2748 (N_2748,N_2467,N_2399);
and U2749 (N_2749,N_2276,N_2437);
nor U2750 (N_2750,N_2507,N_2688);
and U2751 (N_2751,N_2578,N_2685);
nand U2752 (N_2752,N_2530,N_2577);
nand U2753 (N_2753,N_2535,N_2658);
nor U2754 (N_2754,N_2711,N_2721);
and U2755 (N_2755,N_2651,N_2720);
nand U2756 (N_2756,N_2616,N_2654);
and U2757 (N_2757,N_2727,N_2678);
or U2758 (N_2758,N_2510,N_2573);
nor U2759 (N_2759,N_2526,N_2705);
and U2760 (N_2760,N_2565,N_2701);
nor U2761 (N_2761,N_2714,N_2520);
xor U2762 (N_2762,N_2504,N_2503);
nor U2763 (N_2763,N_2562,N_2514);
and U2764 (N_2764,N_2704,N_2706);
or U2765 (N_2765,N_2517,N_2634);
nand U2766 (N_2766,N_2724,N_2686);
nor U2767 (N_2767,N_2670,N_2675);
and U2768 (N_2768,N_2622,N_2599);
xnor U2769 (N_2769,N_2603,N_2738);
nor U2770 (N_2770,N_2570,N_2659);
and U2771 (N_2771,N_2544,N_2575);
nand U2772 (N_2772,N_2615,N_2619);
and U2773 (N_2773,N_2627,N_2630);
nor U2774 (N_2774,N_2568,N_2723);
nand U2775 (N_2775,N_2555,N_2591);
xnor U2776 (N_2776,N_2687,N_2657);
xnor U2777 (N_2777,N_2653,N_2700);
nor U2778 (N_2778,N_2600,N_2731);
xnor U2779 (N_2779,N_2676,N_2744);
nor U2780 (N_2780,N_2741,N_2640);
nor U2781 (N_2781,N_2518,N_2743);
xnor U2782 (N_2782,N_2585,N_2529);
nor U2783 (N_2783,N_2666,N_2541);
nor U2784 (N_2784,N_2549,N_2574);
nand U2785 (N_2785,N_2583,N_2702);
nand U2786 (N_2786,N_2710,N_2642);
xnor U2787 (N_2787,N_2542,N_2554);
or U2788 (N_2788,N_2669,N_2602);
xnor U2789 (N_2789,N_2604,N_2652);
nand U2790 (N_2790,N_2594,N_2567);
nand U2791 (N_2791,N_2580,N_2749);
or U2792 (N_2792,N_2635,N_2537);
and U2793 (N_2793,N_2643,N_2560);
nand U2794 (N_2794,N_2601,N_2558);
xor U2795 (N_2795,N_2709,N_2733);
nor U2796 (N_2796,N_2672,N_2610);
nand U2797 (N_2797,N_2536,N_2725);
or U2798 (N_2798,N_2547,N_2552);
and U2799 (N_2799,N_2606,N_2716);
nor U2800 (N_2800,N_2695,N_2563);
nand U2801 (N_2801,N_2543,N_2506);
and U2802 (N_2802,N_2621,N_2508);
nor U2803 (N_2803,N_2671,N_2501);
or U2804 (N_2804,N_2690,N_2538);
xnor U2805 (N_2805,N_2728,N_2689);
nand U2806 (N_2806,N_2628,N_2593);
nand U2807 (N_2807,N_2557,N_2715);
xor U2808 (N_2808,N_2605,N_2590);
nor U2809 (N_2809,N_2532,N_2735);
nand U2810 (N_2810,N_2699,N_2650);
or U2811 (N_2811,N_2674,N_2533);
and U2812 (N_2812,N_2553,N_2645);
and U2813 (N_2813,N_2729,N_2588);
or U2814 (N_2814,N_2747,N_2667);
xor U2815 (N_2815,N_2608,N_2697);
nor U2816 (N_2816,N_2511,N_2668);
xor U2817 (N_2817,N_2637,N_2717);
xor U2818 (N_2818,N_2513,N_2664);
or U2819 (N_2819,N_2556,N_2576);
or U2820 (N_2820,N_2661,N_2726);
nor U2821 (N_2821,N_2730,N_2523);
or U2822 (N_2822,N_2748,N_2665);
xor U2823 (N_2823,N_2561,N_2703);
nor U2824 (N_2824,N_2698,N_2649);
or U2825 (N_2825,N_2719,N_2519);
and U2826 (N_2826,N_2680,N_2713);
nand U2827 (N_2827,N_2631,N_2647);
and U2828 (N_2828,N_2629,N_2569);
nand U2829 (N_2829,N_2586,N_2626);
nor U2830 (N_2830,N_2636,N_2582);
nand U2831 (N_2831,N_2527,N_2641);
and U2832 (N_2832,N_2732,N_2540);
nand U2833 (N_2833,N_2522,N_2596);
and U2834 (N_2834,N_2740,N_2679);
nor U2835 (N_2835,N_2559,N_2739);
xnor U2836 (N_2836,N_2681,N_2572);
nand U2837 (N_2837,N_2592,N_2742);
nor U2838 (N_2838,N_2548,N_2581);
xor U2839 (N_2839,N_2648,N_2623);
nor U2840 (N_2840,N_2525,N_2673);
nand U2841 (N_2841,N_2737,N_2589);
or U2842 (N_2842,N_2595,N_2618);
nor U2843 (N_2843,N_2745,N_2683);
or U2844 (N_2844,N_2597,N_2662);
and U2845 (N_2845,N_2515,N_2505);
nor U2846 (N_2846,N_2696,N_2613);
nor U2847 (N_2847,N_2620,N_2663);
nand U2848 (N_2848,N_2546,N_2571);
nor U2849 (N_2849,N_2611,N_2660);
or U2850 (N_2850,N_2551,N_2692);
nor U2851 (N_2851,N_2639,N_2587);
nor U2852 (N_2852,N_2584,N_2694);
or U2853 (N_2853,N_2579,N_2656);
nor U2854 (N_2854,N_2682,N_2609);
xor U2855 (N_2855,N_2655,N_2718);
or U2856 (N_2856,N_2617,N_2545);
nor U2857 (N_2857,N_2691,N_2707);
and U2858 (N_2858,N_2677,N_2644);
xor U2859 (N_2859,N_2638,N_2633);
nand U2860 (N_2860,N_2624,N_2612);
and U2861 (N_2861,N_2722,N_2598);
nand U2862 (N_2862,N_2734,N_2566);
xor U2863 (N_2863,N_2500,N_2693);
nor U2864 (N_2864,N_2708,N_2632);
and U2865 (N_2865,N_2502,N_2684);
or U2866 (N_2866,N_2607,N_2512);
nor U2867 (N_2867,N_2539,N_2746);
nand U2868 (N_2868,N_2521,N_2736);
and U2869 (N_2869,N_2516,N_2524);
nand U2870 (N_2870,N_2531,N_2646);
xor U2871 (N_2871,N_2550,N_2625);
or U2872 (N_2872,N_2614,N_2564);
xnor U2873 (N_2873,N_2712,N_2528);
and U2874 (N_2874,N_2509,N_2534);
or U2875 (N_2875,N_2636,N_2540);
xor U2876 (N_2876,N_2676,N_2508);
xor U2877 (N_2877,N_2709,N_2677);
and U2878 (N_2878,N_2626,N_2569);
nor U2879 (N_2879,N_2647,N_2663);
nand U2880 (N_2880,N_2507,N_2727);
xor U2881 (N_2881,N_2583,N_2715);
xor U2882 (N_2882,N_2643,N_2653);
or U2883 (N_2883,N_2745,N_2740);
nor U2884 (N_2884,N_2548,N_2593);
or U2885 (N_2885,N_2726,N_2503);
and U2886 (N_2886,N_2501,N_2708);
xnor U2887 (N_2887,N_2635,N_2581);
or U2888 (N_2888,N_2587,N_2681);
nand U2889 (N_2889,N_2568,N_2699);
nor U2890 (N_2890,N_2636,N_2630);
nand U2891 (N_2891,N_2732,N_2665);
xor U2892 (N_2892,N_2573,N_2675);
and U2893 (N_2893,N_2742,N_2598);
xnor U2894 (N_2894,N_2607,N_2721);
nor U2895 (N_2895,N_2580,N_2501);
and U2896 (N_2896,N_2561,N_2539);
xor U2897 (N_2897,N_2575,N_2624);
or U2898 (N_2898,N_2569,N_2739);
xor U2899 (N_2899,N_2552,N_2708);
nand U2900 (N_2900,N_2530,N_2555);
xnor U2901 (N_2901,N_2565,N_2666);
xor U2902 (N_2902,N_2613,N_2561);
or U2903 (N_2903,N_2581,N_2678);
or U2904 (N_2904,N_2626,N_2719);
and U2905 (N_2905,N_2528,N_2627);
and U2906 (N_2906,N_2556,N_2508);
xor U2907 (N_2907,N_2503,N_2594);
or U2908 (N_2908,N_2629,N_2533);
nor U2909 (N_2909,N_2709,N_2729);
xor U2910 (N_2910,N_2535,N_2599);
xor U2911 (N_2911,N_2702,N_2710);
or U2912 (N_2912,N_2722,N_2717);
nor U2913 (N_2913,N_2670,N_2555);
nor U2914 (N_2914,N_2708,N_2541);
nand U2915 (N_2915,N_2582,N_2595);
nand U2916 (N_2916,N_2531,N_2676);
and U2917 (N_2917,N_2711,N_2631);
or U2918 (N_2918,N_2652,N_2662);
nand U2919 (N_2919,N_2651,N_2551);
nand U2920 (N_2920,N_2684,N_2632);
and U2921 (N_2921,N_2663,N_2730);
nor U2922 (N_2922,N_2595,N_2612);
or U2923 (N_2923,N_2528,N_2520);
nor U2924 (N_2924,N_2561,N_2508);
nor U2925 (N_2925,N_2700,N_2617);
nand U2926 (N_2926,N_2702,N_2551);
xor U2927 (N_2927,N_2705,N_2627);
nand U2928 (N_2928,N_2515,N_2583);
nand U2929 (N_2929,N_2652,N_2634);
and U2930 (N_2930,N_2553,N_2646);
xnor U2931 (N_2931,N_2554,N_2520);
nor U2932 (N_2932,N_2673,N_2591);
nor U2933 (N_2933,N_2533,N_2561);
or U2934 (N_2934,N_2724,N_2550);
xnor U2935 (N_2935,N_2657,N_2533);
and U2936 (N_2936,N_2594,N_2504);
and U2937 (N_2937,N_2550,N_2624);
nand U2938 (N_2938,N_2649,N_2729);
xnor U2939 (N_2939,N_2662,N_2688);
xor U2940 (N_2940,N_2739,N_2551);
or U2941 (N_2941,N_2584,N_2659);
nor U2942 (N_2942,N_2682,N_2588);
nor U2943 (N_2943,N_2654,N_2646);
xnor U2944 (N_2944,N_2745,N_2641);
nor U2945 (N_2945,N_2615,N_2710);
and U2946 (N_2946,N_2642,N_2726);
xnor U2947 (N_2947,N_2668,N_2595);
nand U2948 (N_2948,N_2667,N_2622);
and U2949 (N_2949,N_2522,N_2546);
and U2950 (N_2950,N_2737,N_2644);
or U2951 (N_2951,N_2574,N_2742);
nand U2952 (N_2952,N_2725,N_2643);
xnor U2953 (N_2953,N_2644,N_2587);
and U2954 (N_2954,N_2680,N_2553);
and U2955 (N_2955,N_2537,N_2647);
nand U2956 (N_2956,N_2635,N_2747);
xnor U2957 (N_2957,N_2585,N_2510);
or U2958 (N_2958,N_2685,N_2715);
and U2959 (N_2959,N_2721,N_2744);
nor U2960 (N_2960,N_2519,N_2570);
nor U2961 (N_2961,N_2638,N_2579);
and U2962 (N_2962,N_2637,N_2534);
xor U2963 (N_2963,N_2580,N_2696);
and U2964 (N_2964,N_2646,N_2742);
xor U2965 (N_2965,N_2588,N_2629);
nand U2966 (N_2966,N_2592,N_2715);
xnor U2967 (N_2967,N_2696,N_2726);
xor U2968 (N_2968,N_2659,N_2525);
xor U2969 (N_2969,N_2596,N_2741);
and U2970 (N_2970,N_2556,N_2629);
xor U2971 (N_2971,N_2693,N_2507);
nor U2972 (N_2972,N_2697,N_2525);
xnor U2973 (N_2973,N_2621,N_2520);
and U2974 (N_2974,N_2600,N_2736);
or U2975 (N_2975,N_2532,N_2662);
or U2976 (N_2976,N_2627,N_2731);
and U2977 (N_2977,N_2612,N_2576);
nor U2978 (N_2978,N_2747,N_2653);
nor U2979 (N_2979,N_2591,N_2598);
nor U2980 (N_2980,N_2503,N_2738);
nand U2981 (N_2981,N_2546,N_2701);
or U2982 (N_2982,N_2599,N_2586);
or U2983 (N_2983,N_2623,N_2525);
nor U2984 (N_2984,N_2506,N_2692);
and U2985 (N_2985,N_2567,N_2631);
nand U2986 (N_2986,N_2598,N_2680);
nor U2987 (N_2987,N_2721,N_2652);
nand U2988 (N_2988,N_2645,N_2506);
and U2989 (N_2989,N_2512,N_2552);
xnor U2990 (N_2990,N_2589,N_2672);
nand U2991 (N_2991,N_2736,N_2719);
and U2992 (N_2992,N_2661,N_2557);
or U2993 (N_2993,N_2727,N_2611);
and U2994 (N_2994,N_2581,N_2716);
nor U2995 (N_2995,N_2734,N_2505);
nand U2996 (N_2996,N_2631,N_2644);
xnor U2997 (N_2997,N_2566,N_2500);
nor U2998 (N_2998,N_2535,N_2520);
and U2999 (N_2999,N_2609,N_2570);
nor U3000 (N_3000,N_2846,N_2818);
nor U3001 (N_3001,N_2841,N_2976);
and U3002 (N_3002,N_2861,N_2986);
nand U3003 (N_3003,N_2888,N_2899);
xor U3004 (N_3004,N_2822,N_2914);
xor U3005 (N_3005,N_2840,N_2813);
and U3006 (N_3006,N_2837,N_2919);
nor U3007 (N_3007,N_2759,N_2898);
or U3008 (N_3008,N_2950,N_2956);
and U3009 (N_3009,N_2804,N_2904);
nor U3010 (N_3010,N_2913,N_2799);
nor U3011 (N_3011,N_2912,N_2808);
or U3012 (N_3012,N_2996,N_2774);
or U3013 (N_3013,N_2894,N_2847);
or U3014 (N_3014,N_2869,N_2827);
and U3015 (N_3015,N_2762,N_2926);
xnor U3016 (N_3016,N_2990,N_2892);
xor U3017 (N_3017,N_2787,N_2961);
xor U3018 (N_3018,N_2911,N_2770);
and U3019 (N_3019,N_2987,N_2811);
nor U3020 (N_3020,N_2887,N_2854);
or U3021 (N_3021,N_2865,N_2821);
or U3022 (N_3022,N_2973,N_2751);
xor U3023 (N_3023,N_2766,N_2975);
and U3024 (N_3024,N_2983,N_2752);
or U3025 (N_3025,N_2997,N_2929);
or U3026 (N_3026,N_2858,N_2842);
nand U3027 (N_3027,N_2817,N_2864);
and U3028 (N_3028,N_2793,N_2809);
or U3029 (N_3029,N_2944,N_2848);
xnor U3030 (N_3030,N_2834,N_2939);
nand U3031 (N_3031,N_2977,N_2853);
and U3032 (N_3032,N_2930,N_2931);
xnor U3033 (N_3033,N_2962,N_2844);
or U3034 (N_3034,N_2897,N_2937);
nor U3035 (N_3035,N_2924,N_2768);
xor U3036 (N_3036,N_2780,N_2843);
xor U3037 (N_3037,N_2958,N_2825);
xnor U3038 (N_3038,N_2984,N_2871);
nand U3039 (N_3039,N_2773,N_2771);
nand U3040 (N_3040,N_2850,N_2985);
xnor U3041 (N_3041,N_2935,N_2932);
xor U3042 (N_3042,N_2891,N_2775);
xor U3043 (N_3043,N_2796,N_2948);
and U3044 (N_3044,N_2807,N_2862);
and U3045 (N_3045,N_2765,N_2832);
and U3046 (N_3046,N_2826,N_2873);
nand U3047 (N_3047,N_2916,N_2943);
or U3048 (N_3048,N_2802,N_2782);
xnor U3049 (N_3049,N_2810,N_2798);
or U3050 (N_3050,N_2951,N_2978);
nor U3051 (N_3051,N_2905,N_2790);
nand U3052 (N_3052,N_2814,N_2758);
nand U3053 (N_3053,N_2880,N_2828);
or U3054 (N_3054,N_2901,N_2785);
or U3055 (N_3055,N_2886,N_2941);
or U3056 (N_3056,N_2815,N_2957);
and U3057 (N_3057,N_2812,N_2872);
or U3058 (N_3058,N_2945,N_2753);
or U3059 (N_3059,N_2791,N_2801);
nand U3060 (N_3060,N_2903,N_2769);
nor U3061 (N_3061,N_2927,N_2794);
xor U3062 (N_3062,N_2750,N_2761);
and U3063 (N_3063,N_2756,N_2893);
nand U3064 (N_3064,N_2972,N_2920);
nor U3065 (N_3065,N_2884,N_2999);
nor U3066 (N_3066,N_2772,N_2797);
nor U3067 (N_3067,N_2934,N_2868);
nand U3068 (N_3068,N_2788,N_2806);
xnor U3069 (N_3069,N_2767,N_2980);
and U3070 (N_3070,N_2860,N_2786);
nand U3071 (N_3071,N_2917,N_2968);
nor U3072 (N_3072,N_2795,N_2778);
nor U3073 (N_3073,N_2967,N_2838);
nor U3074 (N_3074,N_2857,N_2994);
nand U3075 (N_3075,N_2960,N_2895);
nand U3076 (N_3076,N_2874,N_2942);
nor U3077 (N_3077,N_2907,N_2852);
or U3078 (N_3078,N_2969,N_2974);
or U3079 (N_3079,N_2993,N_2882);
nand U3080 (N_3080,N_2982,N_2877);
nand U3081 (N_3081,N_2763,N_2781);
or U3082 (N_3082,N_2866,N_2953);
or U3083 (N_3083,N_2764,N_2900);
nor U3084 (N_3084,N_2839,N_2940);
and U3085 (N_3085,N_2889,N_2776);
nor U3086 (N_3086,N_2836,N_2835);
and U3087 (N_3087,N_2979,N_2779);
nand U3088 (N_3088,N_2792,N_2760);
or U3089 (N_3089,N_2970,N_2921);
and U3090 (N_3090,N_2959,N_2928);
nand U3091 (N_3091,N_2964,N_2923);
or U3092 (N_3092,N_2824,N_2754);
and U3093 (N_3093,N_2981,N_2954);
nor U3094 (N_3094,N_2902,N_2820);
nor U3095 (N_3095,N_2816,N_2949);
nand U3096 (N_3096,N_2896,N_2925);
or U3097 (N_3097,N_2805,N_2876);
or U3098 (N_3098,N_2915,N_2933);
and U3099 (N_3099,N_2831,N_2789);
nand U3100 (N_3100,N_2890,N_2946);
nand U3101 (N_3101,N_2856,N_2881);
nand U3102 (N_3102,N_2885,N_2823);
xnor U3103 (N_3103,N_2908,N_2784);
xnor U3104 (N_3104,N_2906,N_2879);
or U3105 (N_3105,N_2938,N_2995);
xnor U3106 (N_3106,N_2851,N_2936);
or U3107 (N_3107,N_2803,N_2988);
nor U3108 (N_3108,N_2845,N_2965);
nor U3109 (N_3109,N_2875,N_2829);
nand U3110 (N_3110,N_2991,N_2998);
or U3111 (N_3111,N_2909,N_2755);
nand U3112 (N_3112,N_2966,N_2819);
or U3113 (N_3113,N_2878,N_2952);
xor U3114 (N_3114,N_2922,N_2918);
or U3115 (N_3115,N_2955,N_2963);
xor U3116 (N_3116,N_2910,N_2830);
nor U3117 (N_3117,N_2863,N_2855);
xnor U3118 (N_3118,N_2859,N_2883);
and U3119 (N_3119,N_2867,N_2971);
and U3120 (N_3120,N_2800,N_2947);
nor U3121 (N_3121,N_2992,N_2833);
or U3122 (N_3122,N_2757,N_2989);
nand U3123 (N_3123,N_2777,N_2849);
nor U3124 (N_3124,N_2783,N_2870);
or U3125 (N_3125,N_2850,N_2996);
nand U3126 (N_3126,N_2810,N_2968);
or U3127 (N_3127,N_2945,N_2994);
nand U3128 (N_3128,N_2952,N_2959);
nor U3129 (N_3129,N_2927,N_2911);
and U3130 (N_3130,N_2866,N_2832);
xnor U3131 (N_3131,N_2905,N_2870);
nor U3132 (N_3132,N_2791,N_2782);
nand U3133 (N_3133,N_2963,N_2832);
or U3134 (N_3134,N_2891,N_2799);
or U3135 (N_3135,N_2834,N_2981);
nand U3136 (N_3136,N_2973,N_2924);
and U3137 (N_3137,N_2785,N_2918);
or U3138 (N_3138,N_2789,N_2775);
or U3139 (N_3139,N_2957,N_2876);
nand U3140 (N_3140,N_2942,N_2986);
or U3141 (N_3141,N_2971,N_2889);
xor U3142 (N_3142,N_2776,N_2933);
and U3143 (N_3143,N_2937,N_2816);
and U3144 (N_3144,N_2787,N_2893);
nor U3145 (N_3145,N_2846,N_2853);
nand U3146 (N_3146,N_2806,N_2922);
xor U3147 (N_3147,N_2759,N_2952);
nor U3148 (N_3148,N_2933,N_2875);
xnor U3149 (N_3149,N_2930,N_2900);
or U3150 (N_3150,N_2766,N_2957);
and U3151 (N_3151,N_2924,N_2790);
nor U3152 (N_3152,N_2784,N_2973);
and U3153 (N_3153,N_2918,N_2945);
xor U3154 (N_3154,N_2911,N_2814);
or U3155 (N_3155,N_2972,N_2915);
nand U3156 (N_3156,N_2892,N_2894);
nand U3157 (N_3157,N_2907,N_2876);
and U3158 (N_3158,N_2933,N_2780);
nand U3159 (N_3159,N_2787,N_2840);
nand U3160 (N_3160,N_2818,N_2963);
nand U3161 (N_3161,N_2823,N_2796);
nand U3162 (N_3162,N_2818,N_2815);
and U3163 (N_3163,N_2801,N_2977);
xor U3164 (N_3164,N_2989,N_2891);
nand U3165 (N_3165,N_2843,N_2851);
and U3166 (N_3166,N_2819,N_2751);
or U3167 (N_3167,N_2931,N_2915);
and U3168 (N_3168,N_2831,N_2752);
xnor U3169 (N_3169,N_2918,N_2881);
and U3170 (N_3170,N_2924,N_2899);
xor U3171 (N_3171,N_2816,N_2772);
nand U3172 (N_3172,N_2871,N_2951);
and U3173 (N_3173,N_2798,N_2940);
xnor U3174 (N_3174,N_2895,N_2874);
nor U3175 (N_3175,N_2800,N_2969);
or U3176 (N_3176,N_2973,N_2951);
xnor U3177 (N_3177,N_2865,N_2997);
nand U3178 (N_3178,N_2906,N_2943);
and U3179 (N_3179,N_2853,N_2839);
nor U3180 (N_3180,N_2813,N_2992);
or U3181 (N_3181,N_2952,N_2974);
nand U3182 (N_3182,N_2782,N_2896);
nand U3183 (N_3183,N_2997,N_2752);
or U3184 (N_3184,N_2828,N_2832);
nor U3185 (N_3185,N_2896,N_2991);
nand U3186 (N_3186,N_2861,N_2823);
or U3187 (N_3187,N_2874,N_2889);
nand U3188 (N_3188,N_2935,N_2989);
or U3189 (N_3189,N_2782,N_2915);
xnor U3190 (N_3190,N_2999,N_2982);
nand U3191 (N_3191,N_2835,N_2887);
and U3192 (N_3192,N_2961,N_2816);
and U3193 (N_3193,N_2864,N_2799);
or U3194 (N_3194,N_2908,N_2875);
and U3195 (N_3195,N_2982,N_2870);
xor U3196 (N_3196,N_2972,N_2764);
and U3197 (N_3197,N_2844,N_2994);
xor U3198 (N_3198,N_2840,N_2992);
and U3199 (N_3199,N_2942,N_2814);
and U3200 (N_3200,N_2938,N_2890);
xor U3201 (N_3201,N_2838,N_2841);
nor U3202 (N_3202,N_2965,N_2975);
and U3203 (N_3203,N_2778,N_2777);
xnor U3204 (N_3204,N_2840,N_2998);
and U3205 (N_3205,N_2775,N_2767);
xor U3206 (N_3206,N_2941,N_2975);
and U3207 (N_3207,N_2865,N_2820);
nand U3208 (N_3208,N_2894,N_2909);
or U3209 (N_3209,N_2757,N_2769);
and U3210 (N_3210,N_2922,N_2798);
xnor U3211 (N_3211,N_2776,N_2784);
xnor U3212 (N_3212,N_2916,N_2951);
xnor U3213 (N_3213,N_2798,N_2854);
nor U3214 (N_3214,N_2849,N_2768);
nor U3215 (N_3215,N_2934,N_2930);
nand U3216 (N_3216,N_2852,N_2861);
nor U3217 (N_3217,N_2827,N_2751);
nor U3218 (N_3218,N_2957,N_2984);
xnor U3219 (N_3219,N_2855,N_2839);
nor U3220 (N_3220,N_2919,N_2954);
nand U3221 (N_3221,N_2905,N_2762);
and U3222 (N_3222,N_2880,N_2923);
nand U3223 (N_3223,N_2944,N_2820);
or U3224 (N_3224,N_2912,N_2763);
and U3225 (N_3225,N_2972,N_2844);
nor U3226 (N_3226,N_2813,N_2851);
nor U3227 (N_3227,N_2991,N_2911);
nor U3228 (N_3228,N_2999,N_2772);
or U3229 (N_3229,N_2783,N_2985);
or U3230 (N_3230,N_2808,N_2904);
or U3231 (N_3231,N_2758,N_2900);
nor U3232 (N_3232,N_2853,N_2829);
and U3233 (N_3233,N_2936,N_2900);
or U3234 (N_3234,N_2801,N_2802);
nand U3235 (N_3235,N_2961,N_2883);
or U3236 (N_3236,N_2877,N_2835);
nor U3237 (N_3237,N_2825,N_2944);
nor U3238 (N_3238,N_2875,N_2805);
xnor U3239 (N_3239,N_2858,N_2905);
or U3240 (N_3240,N_2999,N_2775);
xor U3241 (N_3241,N_2829,N_2804);
nor U3242 (N_3242,N_2904,N_2806);
or U3243 (N_3243,N_2842,N_2900);
nor U3244 (N_3244,N_2963,N_2760);
and U3245 (N_3245,N_2837,N_2853);
nand U3246 (N_3246,N_2929,N_2841);
nor U3247 (N_3247,N_2884,N_2963);
nor U3248 (N_3248,N_2792,N_2931);
and U3249 (N_3249,N_2971,N_2986);
nand U3250 (N_3250,N_3000,N_3006);
or U3251 (N_3251,N_3063,N_3091);
and U3252 (N_3252,N_3004,N_3179);
xnor U3253 (N_3253,N_3078,N_3147);
xnor U3254 (N_3254,N_3047,N_3244);
nor U3255 (N_3255,N_3022,N_3068);
nand U3256 (N_3256,N_3053,N_3216);
and U3257 (N_3257,N_3046,N_3086);
and U3258 (N_3258,N_3090,N_3180);
nor U3259 (N_3259,N_3101,N_3247);
nor U3260 (N_3260,N_3083,N_3201);
nand U3261 (N_3261,N_3059,N_3113);
xnor U3262 (N_3262,N_3164,N_3187);
nand U3263 (N_3263,N_3036,N_3248);
nand U3264 (N_3264,N_3211,N_3028);
and U3265 (N_3265,N_3055,N_3002);
or U3266 (N_3266,N_3171,N_3104);
xor U3267 (N_3267,N_3027,N_3225);
nor U3268 (N_3268,N_3190,N_3238);
nand U3269 (N_3269,N_3135,N_3117);
and U3270 (N_3270,N_3197,N_3156);
nor U3271 (N_3271,N_3108,N_3057);
nor U3272 (N_3272,N_3110,N_3152);
nand U3273 (N_3273,N_3070,N_3178);
and U3274 (N_3274,N_3048,N_3043);
and U3275 (N_3275,N_3236,N_3010);
xnor U3276 (N_3276,N_3231,N_3125);
xor U3277 (N_3277,N_3212,N_3160);
or U3278 (N_3278,N_3207,N_3120);
xor U3279 (N_3279,N_3195,N_3208);
nand U3280 (N_3280,N_3126,N_3194);
nor U3281 (N_3281,N_3039,N_3232);
and U3282 (N_3282,N_3073,N_3162);
nor U3283 (N_3283,N_3122,N_3051);
xor U3284 (N_3284,N_3230,N_3054);
nor U3285 (N_3285,N_3155,N_3132);
nand U3286 (N_3286,N_3173,N_3058);
and U3287 (N_3287,N_3242,N_3204);
nand U3288 (N_3288,N_3089,N_3030);
nand U3289 (N_3289,N_3102,N_3243);
or U3290 (N_3290,N_3001,N_3150);
and U3291 (N_3291,N_3013,N_3129);
xnor U3292 (N_3292,N_3097,N_3241);
nor U3293 (N_3293,N_3200,N_3228);
and U3294 (N_3294,N_3050,N_3192);
or U3295 (N_3295,N_3032,N_3154);
nor U3296 (N_3296,N_3141,N_3240);
and U3297 (N_3297,N_3174,N_3134);
nor U3298 (N_3298,N_3069,N_3100);
xor U3299 (N_3299,N_3014,N_3109);
and U3300 (N_3300,N_3021,N_3220);
and U3301 (N_3301,N_3191,N_3144);
and U3302 (N_3302,N_3139,N_3214);
and U3303 (N_3303,N_3075,N_3016);
nor U3304 (N_3304,N_3119,N_3092);
nor U3305 (N_3305,N_3081,N_3062);
nor U3306 (N_3306,N_3093,N_3177);
or U3307 (N_3307,N_3217,N_3052);
and U3308 (N_3308,N_3105,N_3193);
and U3309 (N_3309,N_3015,N_3229);
nor U3310 (N_3310,N_3095,N_3170);
nand U3311 (N_3311,N_3157,N_3245);
nand U3312 (N_3312,N_3219,N_3088);
nand U3313 (N_3313,N_3153,N_3224);
nand U3314 (N_3314,N_3168,N_3018);
xnor U3315 (N_3315,N_3094,N_3202);
nor U3316 (N_3316,N_3085,N_3246);
nand U3317 (N_3317,N_3124,N_3056);
xnor U3318 (N_3318,N_3060,N_3146);
or U3319 (N_3319,N_3040,N_3133);
nor U3320 (N_3320,N_3106,N_3033);
nor U3321 (N_3321,N_3138,N_3218);
xnor U3322 (N_3322,N_3035,N_3082);
or U3323 (N_3323,N_3130,N_3128);
nand U3324 (N_3324,N_3042,N_3034);
or U3325 (N_3325,N_3025,N_3096);
nand U3326 (N_3326,N_3103,N_3199);
nor U3327 (N_3327,N_3136,N_3067);
nor U3328 (N_3328,N_3205,N_3115);
or U3329 (N_3329,N_3223,N_3080);
nor U3330 (N_3330,N_3038,N_3041);
or U3331 (N_3331,N_3143,N_3003);
and U3332 (N_3332,N_3099,N_3076);
nor U3333 (N_3333,N_3196,N_3142);
xnor U3334 (N_3334,N_3118,N_3175);
or U3335 (N_3335,N_3031,N_3221);
nand U3336 (N_3336,N_3061,N_3227);
nor U3337 (N_3337,N_3186,N_3017);
nand U3338 (N_3338,N_3163,N_3098);
or U3339 (N_3339,N_3049,N_3234);
nor U3340 (N_3340,N_3176,N_3007);
nor U3341 (N_3341,N_3249,N_3233);
nor U3342 (N_3342,N_3158,N_3020);
or U3343 (N_3343,N_3222,N_3084);
or U3344 (N_3344,N_3184,N_3107);
xnor U3345 (N_3345,N_3206,N_3169);
nor U3346 (N_3346,N_3127,N_3065);
and U3347 (N_3347,N_3114,N_3209);
xnor U3348 (N_3348,N_3181,N_3044);
nor U3349 (N_3349,N_3005,N_3198);
nand U3350 (N_3350,N_3116,N_3066);
xnor U3351 (N_3351,N_3210,N_3019);
or U3352 (N_3352,N_3182,N_3188);
or U3353 (N_3353,N_3145,N_3009);
xor U3354 (N_3354,N_3165,N_3226);
or U3355 (N_3355,N_3213,N_3074);
nand U3356 (N_3356,N_3183,N_3166);
and U3357 (N_3357,N_3149,N_3077);
or U3358 (N_3358,N_3123,N_3215);
nand U3359 (N_3359,N_3026,N_3189);
nand U3360 (N_3360,N_3012,N_3237);
xor U3361 (N_3361,N_3079,N_3023);
or U3362 (N_3362,N_3045,N_3159);
nor U3363 (N_3363,N_3185,N_3172);
nand U3364 (N_3364,N_3024,N_3203);
or U3365 (N_3365,N_3161,N_3111);
and U3366 (N_3366,N_3235,N_3071);
and U3367 (N_3367,N_3029,N_3064);
nand U3368 (N_3368,N_3011,N_3131);
and U3369 (N_3369,N_3137,N_3167);
and U3370 (N_3370,N_3140,N_3037);
or U3371 (N_3371,N_3121,N_3148);
and U3372 (N_3372,N_3008,N_3112);
xnor U3373 (N_3373,N_3239,N_3087);
nand U3374 (N_3374,N_3151,N_3072);
xnor U3375 (N_3375,N_3069,N_3124);
and U3376 (N_3376,N_3015,N_3179);
nor U3377 (N_3377,N_3154,N_3214);
or U3378 (N_3378,N_3052,N_3095);
or U3379 (N_3379,N_3215,N_3168);
nor U3380 (N_3380,N_3025,N_3146);
or U3381 (N_3381,N_3024,N_3060);
nand U3382 (N_3382,N_3151,N_3184);
nand U3383 (N_3383,N_3035,N_3150);
xnor U3384 (N_3384,N_3036,N_3167);
and U3385 (N_3385,N_3133,N_3196);
nand U3386 (N_3386,N_3128,N_3071);
nor U3387 (N_3387,N_3039,N_3245);
nor U3388 (N_3388,N_3233,N_3001);
nor U3389 (N_3389,N_3169,N_3030);
and U3390 (N_3390,N_3147,N_3125);
or U3391 (N_3391,N_3184,N_3003);
nor U3392 (N_3392,N_3189,N_3019);
nand U3393 (N_3393,N_3049,N_3224);
xnor U3394 (N_3394,N_3165,N_3233);
nor U3395 (N_3395,N_3088,N_3024);
xor U3396 (N_3396,N_3190,N_3162);
nor U3397 (N_3397,N_3150,N_3013);
xnor U3398 (N_3398,N_3109,N_3022);
or U3399 (N_3399,N_3170,N_3045);
nor U3400 (N_3400,N_3182,N_3117);
nor U3401 (N_3401,N_3089,N_3231);
nand U3402 (N_3402,N_3171,N_3144);
and U3403 (N_3403,N_3066,N_3156);
nor U3404 (N_3404,N_3060,N_3243);
nor U3405 (N_3405,N_3022,N_3234);
nor U3406 (N_3406,N_3126,N_3130);
or U3407 (N_3407,N_3098,N_3160);
or U3408 (N_3408,N_3157,N_3219);
nor U3409 (N_3409,N_3044,N_3249);
xnor U3410 (N_3410,N_3043,N_3079);
nor U3411 (N_3411,N_3195,N_3078);
xnor U3412 (N_3412,N_3058,N_3214);
nand U3413 (N_3413,N_3144,N_3045);
or U3414 (N_3414,N_3083,N_3008);
nand U3415 (N_3415,N_3234,N_3016);
nand U3416 (N_3416,N_3232,N_3144);
xnor U3417 (N_3417,N_3225,N_3010);
nor U3418 (N_3418,N_3234,N_3094);
xor U3419 (N_3419,N_3081,N_3160);
nor U3420 (N_3420,N_3075,N_3081);
nand U3421 (N_3421,N_3060,N_3158);
nor U3422 (N_3422,N_3086,N_3030);
or U3423 (N_3423,N_3132,N_3224);
nor U3424 (N_3424,N_3144,N_3025);
xnor U3425 (N_3425,N_3026,N_3237);
nor U3426 (N_3426,N_3023,N_3046);
nand U3427 (N_3427,N_3174,N_3051);
and U3428 (N_3428,N_3206,N_3125);
nor U3429 (N_3429,N_3168,N_3245);
nor U3430 (N_3430,N_3208,N_3166);
and U3431 (N_3431,N_3151,N_3168);
nand U3432 (N_3432,N_3246,N_3078);
or U3433 (N_3433,N_3128,N_3131);
nor U3434 (N_3434,N_3107,N_3078);
or U3435 (N_3435,N_3225,N_3235);
and U3436 (N_3436,N_3011,N_3110);
and U3437 (N_3437,N_3116,N_3097);
and U3438 (N_3438,N_3058,N_3077);
xor U3439 (N_3439,N_3034,N_3074);
nand U3440 (N_3440,N_3045,N_3016);
nand U3441 (N_3441,N_3073,N_3091);
or U3442 (N_3442,N_3079,N_3016);
xor U3443 (N_3443,N_3131,N_3248);
or U3444 (N_3444,N_3047,N_3118);
nand U3445 (N_3445,N_3067,N_3204);
nand U3446 (N_3446,N_3243,N_3240);
xor U3447 (N_3447,N_3117,N_3033);
or U3448 (N_3448,N_3190,N_3203);
nor U3449 (N_3449,N_3120,N_3200);
or U3450 (N_3450,N_3069,N_3197);
and U3451 (N_3451,N_3080,N_3041);
xor U3452 (N_3452,N_3235,N_3227);
and U3453 (N_3453,N_3203,N_3046);
xnor U3454 (N_3454,N_3035,N_3226);
xor U3455 (N_3455,N_3138,N_3185);
nor U3456 (N_3456,N_3177,N_3014);
nand U3457 (N_3457,N_3020,N_3006);
nand U3458 (N_3458,N_3033,N_3024);
nor U3459 (N_3459,N_3173,N_3139);
nand U3460 (N_3460,N_3086,N_3236);
nand U3461 (N_3461,N_3167,N_3070);
xor U3462 (N_3462,N_3215,N_3214);
xor U3463 (N_3463,N_3198,N_3029);
nand U3464 (N_3464,N_3001,N_3011);
xnor U3465 (N_3465,N_3051,N_3207);
nor U3466 (N_3466,N_3231,N_3134);
or U3467 (N_3467,N_3038,N_3134);
or U3468 (N_3468,N_3063,N_3222);
or U3469 (N_3469,N_3160,N_3216);
nand U3470 (N_3470,N_3044,N_3007);
xor U3471 (N_3471,N_3038,N_3025);
or U3472 (N_3472,N_3049,N_3227);
and U3473 (N_3473,N_3186,N_3008);
nand U3474 (N_3474,N_3165,N_3156);
or U3475 (N_3475,N_3091,N_3029);
xor U3476 (N_3476,N_3165,N_3079);
or U3477 (N_3477,N_3216,N_3027);
and U3478 (N_3478,N_3152,N_3092);
and U3479 (N_3479,N_3153,N_3174);
and U3480 (N_3480,N_3023,N_3230);
and U3481 (N_3481,N_3197,N_3099);
nor U3482 (N_3482,N_3232,N_3054);
nand U3483 (N_3483,N_3109,N_3084);
nand U3484 (N_3484,N_3019,N_3010);
or U3485 (N_3485,N_3098,N_3103);
xor U3486 (N_3486,N_3211,N_3225);
nor U3487 (N_3487,N_3142,N_3106);
and U3488 (N_3488,N_3183,N_3071);
nand U3489 (N_3489,N_3178,N_3062);
and U3490 (N_3490,N_3189,N_3120);
nor U3491 (N_3491,N_3213,N_3217);
nand U3492 (N_3492,N_3247,N_3133);
nand U3493 (N_3493,N_3053,N_3155);
and U3494 (N_3494,N_3141,N_3241);
xor U3495 (N_3495,N_3094,N_3171);
nor U3496 (N_3496,N_3034,N_3157);
xor U3497 (N_3497,N_3037,N_3024);
xor U3498 (N_3498,N_3178,N_3212);
nor U3499 (N_3499,N_3046,N_3237);
nand U3500 (N_3500,N_3358,N_3335);
or U3501 (N_3501,N_3303,N_3301);
and U3502 (N_3502,N_3275,N_3319);
nor U3503 (N_3503,N_3419,N_3296);
or U3504 (N_3504,N_3267,N_3459);
or U3505 (N_3505,N_3450,N_3321);
nor U3506 (N_3506,N_3449,N_3368);
xor U3507 (N_3507,N_3422,N_3351);
xnor U3508 (N_3508,N_3436,N_3452);
or U3509 (N_3509,N_3417,N_3426);
nand U3510 (N_3510,N_3435,N_3390);
nand U3511 (N_3511,N_3377,N_3388);
nor U3512 (N_3512,N_3376,N_3408);
nor U3513 (N_3513,N_3424,N_3473);
or U3514 (N_3514,N_3256,N_3372);
nand U3515 (N_3515,N_3265,N_3404);
or U3516 (N_3516,N_3345,N_3280);
xor U3517 (N_3517,N_3298,N_3400);
and U3518 (N_3518,N_3464,N_3279);
and U3519 (N_3519,N_3340,N_3357);
or U3520 (N_3520,N_3409,N_3371);
and U3521 (N_3521,N_3258,N_3457);
and U3522 (N_3522,N_3297,N_3441);
or U3523 (N_3523,N_3446,N_3468);
nand U3524 (N_3524,N_3407,N_3339);
and U3525 (N_3525,N_3255,N_3437);
nor U3526 (N_3526,N_3363,N_3268);
xor U3527 (N_3527,N_3289,N_3427);
xor U3528 (N_3528,N_3291,N_3253);
and U3529 (N_3529,N_3315,N_3308);
or U3530 (N_3530,N_3278,N_3329);
xor U3531 (N_3531,N_3325,N_3485);
and U3532 (N_3532,N_3354,N_3391);
nor U3533 (N_3533,N_3385,N_3471);
or U3534 (N_3534,N_3346,N_3284);
or U3535 (N_3535,N_3412,N_3314);
or U3536 (N_3536,N_3487,N_3359);
or U3537 (N_3537,N_3469,N_3430);
or U3538 (N_3538,N_3332,N_3456);
and U3539 (N_3539,N_3271,N_3344);
xnor U3540 (N_3540,N_3310,N_3250);
xor U3541 (N_3541,N_3387,N_3465);
nor U3542 (N_3542,N_3270,N_3378);
nor U3543 (N_3543,N_3432,N_3482);
or U3544 (N_3544,N_3431,N_3402);
nor U3545 (N_3545,N_3496,N_3286);
nor U3546 (N_3546,N_3294,N_3269);
nand U3547 (N_3547,N_3331,N_3293);
nor U3548 (N_3548,N_3444,N_3475);
or U3549 (N_3549,N_3379,N_3277);
nor U3550 (N_3550,N_3369,N_3304);
and U3551 (N_3551,N_3395,N_3466);
nand U3552 (N_3552,N_3397,N_3343);
nand U3553 (N_3553,N_3341,N_3266);
nor U3554 (N_3554,N_3361,N_3484);
xor U3555 (N_3555,N_3347,N_3367);
nor U3556 (N_3556,N_3495,N_3491);
or U3557 (N_3557,N_3324,N_3313);
and U3558 (N_3558,N_3362,N_3477);
nor U3559 (N_3559,N_3383,N_3418);
or U3560 (N_3560,N_3393,N_3366);
and U3561 (N_3561,N_3440,N_3492);
nand U3562 (N_3562,N_3447,N_3396);
and U3563 (N_3563,N_3272,N_3423);
nor U3564 (N_3564,N_3474,N_3411);
and U3565 (N_3565,N_3445,N_3406);
xor U3566 (N_3566,N_3288,N_3499);
nand U3567 (N_3567,N_3416,N_3476);
xor U3568 (N_3568,N_3264,N_3355);
xor U3569 (N_3569,N_3311,N_3306);
xnor U3570 (N_3570,N_3300,N_3348);
and U3571 (N_3571,N_3413,N_3338);
or U3572 (N_3572,N_3285,N_3323);
or U3573 (N_3573,N_3403,N_3458);
xnor U3574 (N_3574,N_3330,N_3480);
xor U3575 (N_3575,N_3489,N_3382);
or U3576 (N_3576,N_3381,N_3420);
and U3577 (N_3577,N_3394,N_3454);
xor U3578 (N_3578,N_3439,N_3320);
nor U3579 (N_3579,N_3467,N_3259);
nand U3580 (N_3580,N_3318,N_3360);
or U3581 (N_3581,N_3282,N_3494);
xnor U3582 (N_3582,N_3398,N_3290);
and U3583 (N_3583,N_3380,N_3251);
nor U3584 (N_3584,N_3352,N_3453);
and U3585 (N_3585,N_3309,N_3317);
nand U3586 (N_3586,N_3442,N_3356);
and U3587 (N_3587,N_3305,N_3299);
xnor U3588 (N_3588,N_3287,N_3262);
and U3589 (N_3589,N_3333,N_3448);
nor U3590 (N_3590,N_3302,N_3336);
xor U3591 (N_3591,N_3334,N_3254);
xnor U3592 (N_3592,N_3373,N_3488);
nand U3593 (N_3593,N_3370,N_3433);
xor U3594 (N_3594,N_3364,N_3461);
nand U3595 (N_3595,N_3281,N_3425);
nor U3596 (N_3596,N_3392,N_3405);
nand U3597 (N_3597,N_3415,N_3292);
xor U3598 (N_3598,N_3337,N_3438);
and U3599 (N_3599,N_3316,N_3498);
nand U3600 (N_3600,N_3326,N_3274);
or U3601 (N_3601,N_3327,N_3328);
nor U3602 (N_3602,N_3462,N_3257);
nand U3603 (N_3603,N_3401,N_3283);
nand U3604 (N_3604,N_3463,N_3443);
xnor U3605 (N_3605,N_3389,N_3307);
and U3606 (N_3606,N_3261,N_3276);
xnor U3607 (N_3607,N_3399,N_3429);
and U3608 (N_3608,N_3342,N_3490);
nand U3609 (N_3609,N_3350,N_3479);
nor U3610 (N_3610,N_3493,N_3451);
and U3611 (N_3611,N_3470,N_3428);
nand U3612 (N_3612,N_3263,N_3252);
nor U3613 (N_3613,N_3478,N_3455);
and U3614 (N_3614,N_3472,N_3349);
nor U3615 (N_3615,N_3260,N_3410);
nor U3616 (N_3616,N_3384,N_3365);
nor U3617 (N_3617,N_3295,N_3374);
nor U3618 (N_3618,N_3486,N_3386);
or U3619 (N_3619,N_3481,N_3414);
nand U3620 (N_3620,N_3312,N_3322);
nor U3621 (N_3621,N_3421,N_3483);
and U3622 (N_3622,N_3375,N_3460);
xor U3623 (N_3623,N_3353,N_3434);
xor U3624 (N_3624,N_3497,N_3273);
and U3625 (N_3625,N_3267,N_3250);
xor U3626 (N_3626,N_3406,N_3260);
nand U3627 (N_3627,N_3362,N_3486);
nand U3628 (N_3628,N_3419,N_3336);
and U3629 (N_3629,N_3326,N_3354);
xnor U3630 (N_3630,N_3497,N_3443);
and U3631 (N_3631,N_3284,N_3358);
or U3632 (N_3632,N_3277,N_3355);
nor U3633 (N_3633,N_3316,N_3380);
xnor U3634 (N_3634,N_3327,N_3458);
nand U3635 (N_3635,N_3446,N_3377);
and U3636 (N_3636,N_3281,N_3299);
nor U3637 (N_3637,N_3396,N_3491);
or U3638 (N_3638,N_3462,N_3438);
and U3639 (N_3639,N_3253,N_3391);
and U3640 (N_3640,N_3295,N_3365);
or U3641 (N_3641,N_3415,N_3489);
nor U3642 (N_3642,N_3439,N_3464);
or U3643 (N_3643,N_3485,N_3372);
nand U3644 (N_3644,N_3497,N_3339);
nand U3645 (N_3645,N_3367,N_3314);
nand U3646 (N_3646,N_3317,N_3304);
or U3647 (N_3647,N_3442,N_3325);
nor U3648 (N_3648,N_3255,N_3428);
or U3649 (N_3649,N_3335,N_3474);
or U3650 (N_3650,N_3354,N_3287);
xor U3651 (N_3651,N_3268,N_3451);
nand U3652 (N_3652,N_3401,N_3379);
xor U3653 (N_3653,N_3459,N_3269);
and U3654 (N_3654,N_3449,N_3480);
nor U3655 (N_3655,N_3281,N_3289);
nand U3656 (N_3656,N_3433,N_3309);
xor U3657 (N_3657,N_3360,N_3452);
or U3658 (N_3658,N_3452,N_3433);
xor U3659 (N_3659,N_3321,N_3373);
nor U3660 (N_3660,N_3273,N_3489);
xnor U3661 (N_3661,N_3305,N_3269);
and U3662 (N_3662,N_3264,N_3278);
nor U3663 (N_3663,N_3472,N_3297);
xnor U3664 (N_3664,N_3473,N_3277);
nor U3665 (N_3665,N_3471,N_3382);
nor U3666 (N_3666,N_3435,N_3441);
nand U3667 (N_3667,N_3423,N_3495);
or U3668 (N_3668,N_3460,N_3443);
xor U3669 (N_3669,N_3336,N_3470);
and U3670 (N_3670,N_3251,N_3442);
and U3671 (N_3671,N_3425,N_3310);
nand U3672 (N_3672,N_3290,N_3366);
and U3673 (N_3673,N_3351,N_3313);
nand U3674 (N_3674,N_3425,N_3433);
and U3675 (N_3675,N_3386,N_3348);
and U3676 (N_3676,N_3364,N_3387);
or U3677 (N_3677,N_3404,N_3312);
xnor U3678 (N_3678,N_3404,N_3485);
or U3679 (N_3679,N_3463,N_3324);
and U3680 (N_3680,N_3288,N_3424);
or U3681 (N_3681,N_3384,N_3320);
xor U3682 (N_3682,N_3395,N_3484);
nor U3683 (N_3683,N_3363,N_3320);
and U3684 (N_3684,N_3467,N_3338);
xor U3685 (N_3685,N_3434,N_3320);
or U3686 (N_3686,N_3485,N_3334);
and U3687 (N_3687,N_3467,N_3313);
and U3688 (N_3688,N_3341,N_3453);
and U3689 (N_3689,N_3463,N_3438);
and U3690 (N_3690,N_3302,N_3290);
nor U3691 (N_3691,N_3284,N_3364);
nand U3692 (N_3692,N_3321,N_3423);
and U3693 (N_3693,N_3305,N_3252);
and U3694 (N_3694,N_3328,N_3315);
or U3695 (N_3695,N_3263,N_3487);
nand U3696 (N_3696,N_3317,N_3383);
nand U3697 (N_3697,N_3322,N_3454);
xor U3698 (N_3698,N_3420,N_3262);
nand U3699 (N_3699,N_3463,N_3255);
or U3700 (N_3700,N_3273,N_3301);
xnor U3701 (N_3701,N_3308,N_3283);
xor U3702 (N_3702,N_3481,N_3326);
and U3703 (N_3703,N_3351,N_3296);
nand U3704 (N_3704,N_3280,N_3366);
nand U3705 (N_3705,N_3339,N_3482);
or U3706 (N_3706,N_3292,N_3385);
xor U3707 (N_3707,N_3441,N_3367);
nand U3708 (N_3708,N_3454,N_3325);
or U3709 (N_3709,N_3354,N_3498);
nor U3710 (N_3710,N_3404,N_3432);
and U3711 (N_3711,N_3442,N_3473);
nor U3712 (N_3712,N_3343,N_3361);
xor U3713 (N_3713,N_3295,N_3420);
nor U3714 (N_3714,N_3296,N_3293);
nor U3715 (N_3715,N_3427,N_3473);
nand U3716 (N_3716,N_3251,N_3462);
or U3717 (N_3717,N_3352,N_3282);
and U3718 (N_3718,N_3458,N_3477);
and U3719 (N_3719,N_3255,N_3351);
or U3720 (N_3720,N_3499,N_3455);
nand U3721 (N_3721,N_3290,N_3374);
and U3722 (N_3722,N_3298,N_3474);
xnor U3723 (N_3723,N_3300,N_3290);
xor U3724 (N_3724,N_3436,N_3270);
or U3725 (N_3725,N_3367,N_3469);
or U3726 (N_3726,N_3410,N_3404);
and U3727 (N_3727,N_3395,N_3479);
xor U3728 (N_3728,N_3321,N_3433);
nand U3729 (N_3729,N_3496,N_3270);
nand U3730 (N_3730,N_3441,N_3422);
or U3731 (N_3731,N_3286,N_3359);
nand U3732 (N_3732,N_3314,N_3358);
and U3733 (N_3733,N_3484,N_3306);
or U3734 (N_3734,N_3430,N_3466);
xor U3735 (N_3735,N_3413,N_3341);
nor U3736 (N_3736,N_3385,N_3281);
nand U3737 (N_3737,N_3373,N_3344);
and U3738 (N_3738,N_3449,N_3427);
xnor U3739 (N_3739,N_3463,N_3277);
or U3740 (N_3740,N_3374,N_3497);
xor U3741 (N_3741,N_3304,N_3474);
nor U3742 (N_3742,N_3431,N_3359);
nor U3743 (N_3743,N_3292,N_3283);
or U3744 (N_3744,N_3481,N_3295);
xor U3745 (N_3745,N_3394,N_3343);
or U3746 (N_3746,N_3272,N_3378);
or U3747 (N_3747,N_3300,N_3390);
nor U3748 (N_3748,N_3297,N_3471);
or U3749 (N_3749,N_3468,N_3343);
or U3750 (N_3750,N_3678,N_3570);
nand U3751 (N_3751,N_3704,N_3749);
nand U3752 (N_3752,N_3553,N_3727);
nand U3753 (N_3753,N_3594,N_3710);
and U3754 (N_3754,N_3630,N_3605);
or U3755 (N_3755,N_3644,N_3662);
and U3756 (N_3756,N_3574,N_3646);
xor U3757 (N_3757,N_3683,N_3546);
nand U3758 (N_3758,N_3706,N_3712);
xnor U3759 (N_3759,N_3691,N_3622);
nor U3760 (N_3760,N_3746,N_3620);
or U3761 (N_3761,N_3522,N_3533);
nand U3762 (N_3762,N_3659,N_3614);
nor U3763 (N_3763,N_3571,N_3545);
nor U3764 (N_3764,N_3550,N_3603);
nand U3765 (N_3765,N_3618,N_3657);
or U3766 (N_3766,N_3668,N_3509);
nor U3767 (N_3767,N_3627,N_3557);
xnor U3768 (N_3768,N_3588,N_3673);
nand U3769 (N_3769,N_3578,N_3529);
xnor U3770 (N_3770,N_3548,N_3595);
nand U3771 (N_3771,N_3699,N_3591);
nor U3772 (N_3772,N_3613,N_3608);
xor U3773 (N_3773,N_3601,N_3525);
xnor U3774 (N_3774,N_3607,N_3516);
xor U3775 (N_3775,N_3701,N_3676);
or U3776 (N_3776,N_3742,N_3667);
and U3777 (N_3777,N_3636,N_3530);
nor U3778 (N_3778,N_3711,N_3729);
nor U3779 (N_3779,N_3737,N_3590);
or U3780 (N_3780,N_3584,N_3615);
and U3781 (N_3781,N_3625,N_3649);
nand U3782 (N_3782,N_3521,N_3652);
and U3783 (N_3783,N_3748,N_3563);
or U3784 (N_3784,N_3599,N_3573);
nand U3785 (N_3785,N_3558,N_3684);
nor U3786 (N_3786,N_3747,N_3628);
nor U3787 (N_3787,N_3612,N_3585);
nand U3788 (N_3788,N_3566,N_3515);
or U3789 (N_3789,N_3726,N_3554);
or U3790 (N_3790,N_3645,N_3643);
xnor U3791 (N_3791,N_3587,N_3555);
and U3792 (N_3792,N_3739,N_3617);
or U3793 (N_3793,N_3675,N_3561);
xor U3794 (N_3794,N_3559,N_3709);
and U3795 (N_3795,N_3682,N_3718);
and U3796 (N_3796,N_3592,N_3536);
xor U3797 (N_3797,N_3695,N_3689);
or U3798 (N_3798,N_3549,N_3671);
nor U3799 (N_3799,N_3518,N_3565);
and U3800 (N_3800,N_3621,N_3714);
and U3801 (N_3801,N_3661,N_3735);
xor U3802 (N_3802,N_3506,N_3586);
and U3803 (N_3803,N_3688,N_3740);
nor U3804 (N_3804,N_3719,N_3696);
nor U3805 (N_3805,N_3531,N_3653);
or U3806 (N_3806,N_3505,N_3564);
xor U3807 (N_3807,N_3519,N_3744);
xnor U3808 (N_3808,N_3686,N_3654);
nand U3809 (N_3809,N_3658,N_3543);
xnor U3810 (N_3810,N_3582,N_3637);
nor U3811 (N_3811,N_3725,N_3743);
nand U3812 (N_3812,N_3631,N_3513);
and U3813 (N_3813,N_3647,N_3579);
or U3814 (N_3814,N_3745,N_3732);
and U3815 (N_3815,N_3641,N_3639);
xnor U3816 (N_3816,N_3532,N_3619);
or U3817 (N_3817,N_3560,N_3730);
or U3818 (N_3818,N_3656,N_3523);
xor U3819 (N_3819,N_3700,N_3716);
or U3820 (N_3820,N_3634,N_3514);
xnor U3821 (N_3821,N_3538,N_3537);
or U3822 (N_3822,N_3508,N_3660);
and U3823 (N_3823,N_3604,N_3542);
nand U3824 (N_3824,N_3524,N_3694);
nor U3825 (N_3825,N_3648,N_3504);
xnor U3826 (N_3826,N_3741,N_3674);
or U3827 (N_3827,N_3650,N_3633);
nor U3828 (N_3828,N_3562,N_3534);
nand U3829 (N_3829,N_3707,N_3670);
or U3830 (N_3830,N_3611,N_3581);
and U3831 (N_3831,N_3517,N_3567);
nor U3832 (N_3832,N_3677,N_3723);
nor U3833 (N_3833,N_3609,N_3552);
and U3834 (N_3834,N_3501,N_3717);
nand U3835 (N_3835,N_3593,N_3596);
and U3836 (N_3836,N_3575,N_3512);
nand U3837 (N_3837,N_3663,N_3669);
nor U3838 (N_3838,N_3640,N_3572);
and U3839 (N_3839,N_3638,N_3728);
nand U3840 (N_3840,N_3629,N_3526);
or U3841 (N_3841,N_3527,N_3721);
nand U3842 (N_3842,N_3708,N_3540);
and U3843 (N_3843,N_3606,N_3734);
xor U3844 (N_3844,N_3502,N_3507);
or U3845 (N_3845,N_3693,N_3597);
and U3846 (N_3846,N_3568,N_3713);
xnor U3847 (N_3847,N_3528,N_3642);
nor U3848 (N_3848,N_3635,N_3626);
xnor U3849 (N_3849,N_3722,N_3510);
or U3850 (N_3850,N_3705,N_3632);
xnor U3851 (N_3851,N_3598,N_3580);
or U3852 (N_3852,N_3583,N_3616);
or U3853 (N_3853,N_3544,N_3623);
and U3854 (N_3854,N_3535,N_3511);
xor U3855 (N_3855,N_3500,N_3503);
or U3856 (N_3856,N_3731,N_3520);
or U3857 (N_3857,N_3738,N_3551);
nand U3858 (N_3858,N_3679,N_3733);
nand U3859 (N_3859,N_3539,N_3724);
xnor U3860 (N_3860,N_3692,N_3541);
nand U3861 (N_3861,N_3720,N_3576);
xor U3862 (N_3862,N_3624,N_3697);
nand U3863 (N_3863,N_3547,N_3685);
nand U3864 (N_3864,N_3680,N_3651);
or U3865 (N_3865,N_3664,N_3589);
and U3866 (N_3866,N_3602,N_3610);
nor U3867 (N_3867,N_3655,N_3556);
nor U3868 (N_3868,N_3703,N_3600);
xor U3869 (N_3869,N_3569,N_3715);
or U3870 (N_3870,N_3690,N_3665);
or U3871 (N_3871,N_3736,N_3672);
nor U3872 (N_3872,N_3702,N_3681);
nor U3873 (N_3873,N_3687,N_3698);
or U3874 (N_3874,N_3577,N_3666);
nand U3875 (N_3875,N_3640,N_3556);
nand U3876 (N_3876,N_3733,N_3637);
or U3877 (N_3877,N_3739,N_3613);
nor U3878 (N_3878,N_3672,N_3686);
xor U3879 (N_3879,N_3717,N_3668);
xor U3880 (N_3880,N_3688,N_3721);
nor U3881 (N_3881,N_3702,N_3583);
or U3882 (N_3882,N_3617,N_3590);
xor U3883 (N_3883,N_3575,N_3694);
nor U3884 (N_3884,N_3564,N_3617);
nand U3885 (N_3885,N_3681,N_3591);
or U3886 (N_3886,N_3720,N_3722);
nor U3887 (N_3887,N_3668,N_3533);
nor U3888 (N_3888,N_3572,N_3536);
nor U3889 (N_3889,N_3623,N_3653);
xor U3890 (N_3890,N_3597,N_3567);
xor U3891 (N_3891,N_3719,N_3745);
nor U3892 (N_3892,N_3699,N_3541);
nor U3893 (N_3893,N_3735,N_3539);
nor U3894 (N_3894,N_3674,N_3544);
or U3895 (N_3895,N_3731,N_3589);
nor U3896 (N_3896,N_3654,N_3657);
or U3897 (N_3897,N_3746,N_3691);
nand U3898 (N_3898,N_3662,N_3660);
or U3899 (N_3899,N_3575,N_3624);
nand U3900 (N_3900,N_3622,N_3589);
nand U3901 (N_3901,N_3551,N_3644);
nor U3902 (N_3902,N_3615,N_3712);
nor U3903 (N_3903,N_3746,N_3524);
and U3904 (N_3904,N_3598,N_3723);
and U3905 (N_3905,N_3728,N_3688);
nor U3906 (N_3906,N_3583,N_3740);
or U3907 (N_3907,N_3557,N_3741);
or U3908 (N_3908,N_3682,N_3642);
nor U3909 (N_3909,N_3587,N_3724);
or U3910 (N_3910,N_3683,N_3681);
and U3911 (N_3911,N_3616,N_3657);
nand U3912 (N_3912,N_3530,N_3570);
nor U3913 (N_3913,N_3641,N_3668);
and U3914 (N_3914,N_3732,N_3743);
or U3915 (N_3915,N_3565,N_3653);
or U3916 (N_3916,N_3648,N_3528);
or U3917 (N_3917,N_3582,N_3697);
and U3918 (N_3918,N_3731,N_3670);
xnor U3919 (N_3919,N_3595,N_3538);
nor U3920 (N_3920,N_3746,N_3517);
nand U3921 (N_3921,N_3558,N_3699);
nand U3922 (N_3922,N_3538,N_3576);
xor U3923 (N_3923,N_3649,N_3711);
nand U3924 (N_3924,N_3645,N_3642);
or U3925 (N_3925,N_3506,N_3507);
and U3926 (N_3926,N_3520,N_3588);
nand U3927 (N_3927,N_3548,N_3577);
xnor U3928 (N_3928,N_3709,N_3665);
xor U3929 (N_3929,N_3715,N_3502);
nand U3930 (N_3930,N_3662,N_3712);
and U3931 (N_3931,N_3670,N_3570);
and U3932 (N_3932,N_3559,N_3510);
nand U3933 (N_3933,N_3668,N_3536);
or U3934 (N_3934,N_3688,N_3715);
and U3935 (N_3935,N_3659,N_3545);
and U3936 (N_3936,N_3653,N_3567);
xnor U3937 (N_3937,N_3613,N_3698);
xor U3938 (N_3938,N_3556,N_3674);
nand U3939 (N_3939,N_3737,N_3655);
xnor U3940 (N_3940,N_3524,N_3564);
nand U3941 (N_3941,N_3632,N_3713);
nor U3942 (N_3942,N_3568,N_3537);
nand U3943 (N_3943,N_3689,N_3656);
nor U3944 (N_3944,N_3529,N_3712);
or U3945 (N_3945,N_3637,N_3639);
nor U3946 (N_3946,N_3597,N_3608);
nand U3947 (N_3947,N_3627,N_3625);
nand U3948 (N_3948,N_3616,N_3570);
nand U3949 (N_3949,N_3745,N_3646);
nor U3950 (N_3950,N_3675,N_3588);
or U3951 (N_3951,N_3532,N_3540);
or U3952 (N_3952,N_3675,N_3696);
or U3953 (N_3953,N_3738,N_3745);
nand U3954 (N_3954,N_3726,N_3688);
xor U3955 (N_3955,N_3718,N_3520);
nor U3956 (N_3956,N_3604,N_3737);
nor U3957 (N_3957,N_3612,N_3646);
nand U3958 (N_3958,N_3704,N_3526);
xnor U3959 (N_3959,N_3586,N_3576);
nor U3960 (N_3960,N_3624,N_3703);
xnor U3961 (N_3961,N_3580,N_3657);
xnor U3962 (N_3962,N_3616,N_3747);
nand U3963 (N_3963,N_3616,N_3607);
nand U3964 (N_3964,N_3596,N_3671);
or U3965 (N_3965,N_3531,N_3677);
xnor U3966 (N_3966,N_3687,N_3523);
and U3967 (N_3967,N_3712,N_3562);
and U3968 (N_3968,N_3674,N_3548);
nand U3969 (N_3969,N_3514,N_3550);
xor U3970 (N_3970,N_3668,N_3590);
or U3971 (N_3971,N_3601,N_3539);
xnor U3972 (N_3972,N_3684,N_3696);
and U3973 (N_3973,N_3627,N_3517);
or U3974 (N_3974,N_3567,N_3668);
nand U3975 (N_3975,N_3541,N_3508);
or U3976 (N_3976,N_3570,N_3745);
nor U3977 (N_3977,N_3651,N_3535);
xor U3978 (N_3978,N_3633,N_3624);
and U3979 (N_3979,N_3511,N_3678);
nand U3980 (N_3980,N_3538,N_3706);
or U3981 (N_3981,N_3583,N_3582);
and U3982 (N_3982,N_3507,N_3584);
nand U3983 (N_3983,N_3559,N_3692);
or U3984 (N_3984,N_3622,N_3539);
nand U3985 (N_3985,N_3618,N_3706);
and U3986 (N_3986,N_3660,N_3640);
or U3987 (N_3987,N_3530,N_3593);
nand U3988 (N_3988,N_3555,N_3616);
and U3989 (N_3989,N_3557,N_3550);
nor U3990 (N_3990,N_3543,N_3665);
and U3991 (N_3991,N_3743,N_3642);
nor U3992 (N_3992,N_3590,N_3680);
nor U3993 (N_3993,N_3585,N_3554);
nor U3994 (N_3994,N_3560,N_3705);
or U3995 (N_3995,N_3686,N_3565);
or U3996 (N_3996,N_3723,N_3517);
or U3997 (N_3997,N_3689,N_3609);
or U3998 (N_3998,N_3652,N_3579);
nor U3999 (N_3999,N_3632,N_3536);
xnor U4000 (N_4000,N_3840,N_3988);
and U4001 (N_4001,N_3784,N_3806);
xnor U4002 (N_4002,N_3895,N_3877);
or U4003 (N_4003,N_3880,N_3925);
xor U4004 (N_4004,N_3957,N_3845);
and U4005 (N_4005,N_3930,N_3859);
and U4006 (N_4006,N_3766,N_3832);
or U4007 (N_4007,N_3756,N_3808);
or U4008 (N_4008,N_3935,N_3867);
nand U4009 (N_4009,N_3800,N_3862);
and U4010 (N_4010,N_3922,N_3948);
nand U4011 (N_4011,N_3855,N_3952);
xnor U4012 (N_4012,N_3753,N_3975);
nand U4013 (N_4013,N_3803,N_3940);
and U4014 (N_4014,N_3857,N_3819);
nor U4015 (N_4015,N_3900,N_3906);
nand U4016 (N_4016,N_3834,N_3913);
or U4017 (N_4017,N_3780,N_3983);
and U4018 (N_4018,N_3951,N_3801);
or U4019 (N_4019,N_3821,N_3762);
nor U4020 (N_4020,N_3882,N_3782);
or U4021 (N_4021,N_3865,N_3890);
xor U4022 (N_4022,N_3994,N_3998);
nand U4023 (N_4023,N_3751,N_3933);
and U4024 (N_4024,N_3968,N_3807);
and U4025 (N_4025,N_3879,N_3770);
or U4026 (N_4026,N_3868,N_3854);
or U4027 (N_4027,N_3896,N_3934);
and U4028 (N_4028,N_3897,N_3969);
or U4029 (N_4029,N_3781,N_3919);
or U4030 (N_4030,N_3822,N_3920);
and U4031 (N_4031,N_3873,N_3778);
nor U4032 (N_4032,N_3804,N_3851);
nor U4033 (N_4033,N_3826,N_3980);
nor U4034 (N_4034,N_3899,N_3908);
xor U4035 (N_4035,N_3964,N_3771);
or U4036 (N_4036,N_3966,N_3984);
and U4037 (N_4037,N_3829,N_3789);
and U4038 (N_4038,N_3788,N_3838);
and U4039 (N_4039,N_3786,N_3767);
nor U4040 (N_4040,N_3946,N_3950);
xor U4041 (N_4041,N_3811,N_3949);
nor U4042 (N_4042,N_3870,N_3985);
nand U4043 (N_4043,N_3905,N_3765);
nand U4044 (N_4044,N_3961,N_3792);
nor U4045 (N_4045,N_3907,N_3953);
nand U4046 (N_4046,N_3939,N_3818);
and U4047 (N_4047,N_3777,N_3794);
nor U4048 (N_4048,N_3866,N_3912);
and U4049 (N_4049,N_3881,N_3790);
nor U4050 (N_4050,N_3978,N_3760);
xnor U4051 (N_4051,N_3916,N_3847);
xnor U4052 (N_4052,N_3996,N_3885);
xnor U4053 (N_4053,N_3901,N_3954);
nor U4054 (N_4054,N_3918,N_3893);
or U4055 (N_4055,N_3944,N_3763);
nor U4056 (N_4056,N_3850,N_3843);
nor U4057 (N_4057,N_3926,N_3904);
and U4058 (N_4058,N_3837,N_3871);
or U4059 (N_4059,N_3962,N_3960);
nor U4060 (N_4060,N_3755,N_3924);
nand U4061 (N_4061,N_3772,N_3793);
nor U4062 (N_4062,N_3970,N_3973);
nor U4063 (N_4063,N_3750,N_3999);
xor U4064 (N_4064,N_3945,N_3846);
nand U4065 (N_4065,N_3863,N_3997);
and U4066 (N_4066,N_3910,N_3989);
nand U4067 (N_4067,N_3842,N_3974);
nand U4068 (N_4068,N_3848,N_3884);
and U4069 (N_4069,N_3936,N_3991);
or U4070 (N_4070,N_3956,N_3785);
nor U4071 (N_4071,N_3827,N_3835);
nor U4072 (N_4072,N_3876,N_3887);
nand U4073 (N_4073,N_3982,N_3820);
nand U4074 (N_4074,N_3754,N_3815);
nand U4075 (N_4075,N_3776,N_3764);
nor U4076 (N_4076,N_3883,N_3909);
nor U4077 (N_4077,N_3987,N_3813);
xnor U4078 (N_4078,N_3932,N_3959);
or U4079 (N_4079,N_3903,N_3955);
xor U4080 (N_4080,N_3894,N_3856);
nand U4081 (N_4081,N_3931,N_3824);
nor U4082 (N_4082,N_3878,N_3779);
nor U4083 (N_4083,N_3927,N_3875);
xor U4084 (N_4084,N_3937,N_3796);
or U4085 (N_4085,N_3928,N_3942);
or U4086 (N_4086,N_3849,N_3993);
nor U4087 (N_4087,N_3810,N_3830);
nor U4088 (N_4088,N_3795,N_3990);
nor U4089 (N_4089,N_3947,N_3773);
xor U4090 (N_4090,N_3938,N_3774);
xnor U4091 (N_4091,N_3891,N_3823);
nor U4092 (N_4092,N_3943,N_3844);
or U4093 (N_4093,N_3941,N_3825);
xnor U4094 (N_4094,N_3972,N_3965);
and U4095 (N_4095,N_3787,N_3967);
nor U4096 (N_4096,N_3992,N_3981);
or U4097 (N_4097,N_3802,N_3977);
or U4098 (N_4098,N_3995,N_3915);
or U4099 (N_4099,N_3963,N_3914);
nand U4100 (N_4100,N_3864,N_3836);
nor U4101 (N_4101,N_3828,N_3869);
nor U4102 (N_4102,N_3917,N_3757);
nand U4103 (N_4103,N_3759,N_3911);
or U4104 (N_4104,N_3791,N_3783);
or U4105 (N_4105,N_3979,N_3775);
nor U4106 (N_4106,N_3860,N_3817);
or U4107 (N_4107,N_3923,N_3902);
and U4108 (N_4108,N_3976,N_3858);
and U4109 (N_4109,N_3889,N_3814);
nand U4110 (N_4110,N_3886,N_3861);
nor U4111 (N_4111,N_3833,N_3971);
or U4112 (N_4112,N_3986,N_3768);
nand U4113 (N_4113,N_3816,N_3841);
or U4114 (N_4114,N_3799,N_3809);
xnor U4115 (N_4115,N_3761,N_3852);
xnor U4116 (N_4116,N_3853,N_3797);
nand U4117 (N_4117,N_3839,N_3752);
xnor U4118 (N_4118,N_3798,N_3929);
or U4119 (N_4119,N_3758,N_3769);
and U4120 (N_4120,N_3874,N_3812);
nand U4121 (N_4121,N_3958,N_3805);
nand U4122 (N_4122,N_3921,N_3872);
or U4123 (N_4123,N_3888,N_3892);
and U4124 (N_4124,N_3831,N_3898);
nor U4125 (N_4125,N_3997,N_3949);
xnor U4126 (N_4126,N_3851,N_3948);
and U4127 (N_4127,N_3756,N_3772);
or U4128 (N_4128,N_3967,N_3872);
nor U4129 (N_4129,N_3899,N_3756);
xnor U4130 (N_4130,N_3750,N_3915);
xnor U4131 (N_4131,N_3948,N_3989);
nand U4132 (N_4132,N_3955,N_3933);
and U4133 (N_4133,N_3945,N_3791);
and U4134 (N_4134,N_3986,N_3850);
xnor U4135 (N_4135,N_3962,N_3833);
or U4136 (N_4136,N_3769,N_3754);
nor U4137 (N_4137,N_3903,N_3926);
or U4138 (N_4138,N_3883,N_3926);
nand U4139 (N_4139,N_3953,N_3912);
xnor U4140 (N_4140,N_3981,N_3834);
xnor U4141 (N_4141,N_3939,N_3804);
nand U4142 (N_4142,N_3781,N_3998);
nor U4143 (N_4143,N_3868,N_3812);
xnor U4144 (N_4144,N_3913,N_3890);
and U4145 (N_4145,N_3850,N_3851);
or U4146 (N_4146,N_3904,N_3831);
xor U4147 (N_4147,N_3993,N_3759);
nor U4148 (N_4148,N_3760,N_3983);
or U4149 (N_4149,N_3923,N_3916);
and U4150 (N_4150,N_3842,N_3831);
nor U4151 (N_4151,N_3770,N_3863);
nand U4152 (N_4152,N_3894,N_3893);
nor U4153 (N_4153,N_3891,N_3868);
nor U4154 (N_4154,N_3968,N_3997);
xnor U4155 (N_4155,N_3845,N_3882);
nor U4156 (N_4156,N_3824,N_3946);
or U4157 (N_4157,N_3938,N_3952);
xor U4158 (N_4158,N_3943,N_3856);
or U4159 (N_4159,N_3987,N_3784);
nand U4160 (N_4160,N_3967,N_3751);
nor U4161 (N_4161,N_3878,N_3809);
xnor U4162 (N_4162,N_3990,N_3775);
nor U4163 (N_4163,N_3790,N_3780);
nor U4164 (N_4164,N_3962,N_3912);
or U4165 (N_4165,N_3755,N_3868);
nor U4166 (N_4166,N_3866,N_3808);
xor U4167 (N_4167,N_3750,N_3779);
or U4168 (N_4168,N_3968,N_3826);
nand U4169 (N_4169,N_3855,N_3832);
or U4170 (N_4170,N_3822,N_3828);
and U4171 (N_4171,N_3799,N_3993);
or U4172 (N_4172,N_3929,N_3901);
nand U4173 (N_4173,N_3761,N_3960);
xnor U4174 (N_4174,N_3862,N_3832);
nor U4175 (N_4175,N_3792,N_3827);
xor U4176 (N_4176,N_3790,N_3800);
nand U4177 (N_4177,N_3914,N_3872);
or U4178 (N_4178,N_3769,N_3911);
or U4179 (N_4179,N_3877,N_3918);
or U4180 (N_4180,N_3761,N_3858);
nor U4181 (N_4181,N_3839,N_3890);
nor U4182 (N_4182,N_3904,N_3766);
xnor U4183 (N_4183,N_3987,N_3859);
and U4184 (N_4184,N_3887,N_3856);
nor U4185 (N_4185,N_3992,N_3892);
nand U4186 (N_4186,N_3866,N_3916);
nand U4187 (N_4187,N_3799,N_3857);
xnor U4188 (N_4188,N_3847,N_3805);
xor U4189 (N_4189,N_3981,N_3777);
and U4190 (N_4190,N_3882,N_3871);
or U4191 (N_4191,N_3839,N_3849);
and U4192 (N_4192,N_3764,N_3998);
xnor U4193 (N_4193,N_3924,N_3975);
and U4194 (N_4194,N_3779,N_3906);
and U4195 (N_4195,N_3875,N_3774);
nand U4196 (N_4196,N_3842,N_3800);
or U4197 (N_4197,N_3846,N_3951);
or U4198 (N_4198,N_3822,N_3769);
xor U4199 (N_4199,N_3946,N_3819);
or U4200 (N_4200,N_3872,N_3851);
nor U4201 (N_4201,N_3824,N_3812);
or U4202 (N_4202,N_3750,N_3812);
and U4203 (N_4203,N_3823,N_3947);
nand U4204 (N_4204,N_3951,N_3898);
nand U4205 (N_4205,N_3972,N_3863);
and U4206 (N_4206,N_3888,N_3958);
and U4207 (N_4207,N_3977,N_3912);
or U4208 (N_4208,N_3846,N_3758);
and U4209 (N_4209,N_3977,N_3797);
xnor U4210 (N_4210,N_3841,N_3979);
nor U4211 (N_4211,N_3782,N_3883);
nor U4212 (N_4212,N_3976,N_3787);
nor U4213 (N_4213,N_3799,N_3813);
and U4214 (N_4214,N_3980,N_3831);
xnor U4215 (N_4215,N_3794,N_3944);
or U4216 (N_4216,N_3965,N_3896);
or U4217 (N_4217,N_3848,N_3801);
or U4218 (N_4218,N_3832,N_3948);
or U4219 (N_4219,N_3796,N_3820);
nor U4220 (N_4220,N_3958,N_3926);
xnor U4221 (N_4221,N_3849,N_3900);
nand U4222 (N_4222,N_3805,N_3837);
and U4223 (N_4223,N_3794,N_3955);
and U4224 (N_4224,N_3831,N_3779);
nor U4225 (N_4225,N_3975,N_3814);
nand U4226 (N_4226,N_3976,N_3996);
and U4227 (N_4227,N_3999,N_3987);
or U4228 (N_4228,N_3864,N_3756);
nor U4229 (N_4229,N_3754,N_3757);
nor U4230 (N_4230,N_3930,N_3952);
or U4231 (N_4231,N_3896,N_3899);
or U4232 (N_4232,N_3857,N_3946);
xor U4233 (N_4233,N_3937,N_3964);
and U4234 (N_4234,N_3821,N_3891);
or U4235 (N_4235,N_3839,N_3913);
xnor U4236 (N_4236,N_3820,N_3967);
nor U4237 (N_4237,N_3965,N_3884);
or U4238 (N_4238,N_3995,N_3850);
nor U4239 (N_4239,N_3941,N_3752);
and U4240 (N_4240,N_3952,N_3934);
nand U4241 (N_4241,N_3990,N_3825);
nand U4242 (N_4242,N_3929,N_3994);
xor U4243 (N_4243,N_3972,N_3841);
nand U4244 (N_4244,N_3913,N_3974);
and U4245 (N_4245,N_3954,N_3969);
xnor U4246 (N_4246,N_3815,N_3898);
nor U4247 (N_4247,N_3891,N_3914);
and U4248 (N_4248,N_3985,N_3907);
nor U4249 (N_4249,N_3864,N_3868);
xnor U4250 (N_4250,N_4100,N_4067);
nand U4251 (N_4251,N_4203,N_4059);
and U4252 (N_4252,N_4160,N_4217);
nor U4253 (N_4253,N_4185,N_4164);
or U4254 (N_4254,N_4231,N_4032);
and U4255 (N_4255,N_4183,N_4145);
xnor U4256 (N_4256,N_4248,N_4001);
or U4257 (N_4257,N_4037,N_4191);
and U4258 (N_4258,N_4193,N_4036);
or U4259 (N_4259,N_4058,N_4192);
and U4260 (N_4260,N_4149,N_4107);
and U4261 (N_4261,N_4009,N_4008);
nor U4262 (N_4262,N_4152,N_4043);
and U4263 (N_4263,N_4233,N_4177);
or U4264 (N_4264,N_4092,N_4179);
nor U4265 (N_4265,N_4141,N_4096);
and U4266 (N_4266,N_4053,N_4035);
and U4267 (N_4267,N_4181,N_4031);
nor U4268 (N_4268,N_4065,N_4155);
xor U4269 (N_4269,N_4225,N_4218);
xnor U4270 (N_4270,N_4243,N_4024);
nand U4271 (N_4271,N_4212,N_4010);
or U4272 (N_4272,N_4121,N_4077);
xnor U4273 (N_4273,N_4049,N_4142);
nor U4274 (N_4274,N_4219,N_4097);
and U4275 (N_4275,N_4169,N_4029);
and U4276 (N_4276,N_4200,N_4040);
xnor U4277 (N_4277,N_4144,N_4020);
nor U4278 (N_4278,N_4112,N_4066);
xor U4279 (N_4279,N_4108,N_4197);
or U4280 (N_4280,N_4114,N_4028);
or U4281 (N_4281,N_4237,N_4215);
nand U4282 (N_4282,N_4165,N_4126);
and U4283 (N_4283,N_4079,N_4073);
xor U4284 (N_4284,N_4161,N_4245);
nor U4285 (N_4285,N_4041,N_4115);
nand U4286 (N_4286,N_4015,N_4137);
or U4287 (N_4287,N_4188,N_4175);
or U4288 (N_4288,N_4125,N_4202);
xnor U4289 (N_4289,N_4246,N_4054);
nand U4290 (N_4290,N_4083,N_4147);
nor U4291 (N_4291,N_4078,N_4006);
and U4292 (N_4292,N_4148,N_4071);
xnor U4293 (N_4293,N_4017,N_4012);
and U4294 (N_4294,N_4234,N_4135);
nand U4295 (N_4295,N_4195,N_4194);
nor U4296 (N_4296,N_4146,N_4238);
and U4297 (N_4297,N_4076,N_4176);
nor U4298 (N_4298,N_4064,N_4063);
and U4299 (N_4299,N_4180,N_4089);
nand U4300 (N_4300,N_4127,N_4047);
or U4301 (N_4301,N_4061,N_4099);
nand U4302 (N_4302,N_4232,N_4023);
nand U4303 (N_4303,N_4018,N_4124);
nor U4304 (N_4304,N_4004,N_4174);
nand U4305 (N_4305,N_4226,N_4038);
or U4306 (N_4306,N_4060,N_4143);
nand U4307 (N_4307,N_4014,N_4025);
nand U4308 (N_4308,N_4221,N_4241);
nand U4309 (N_4309,N_4207,N_4211);
and U4310 (N_4310,N_4138,N_4156);
xor U4311 (N_4311,N_4206,N_4044);
nand U4312 (N_4312,N_4209,N_4210);
nand U4313 (N_4313,N_4201,N_4110);
or U4314 (N_4314,N_4190,N_4111);
nand U4315 (N_4315,N_4055,N_4187);
and U4316 (N_4316,N_4122,N_4132);
xor U4317 (N_4317,N_4056,N_4227);
or U4318 (N_4318,N_4204,N_4003);
and U4319 (N_4319,N_4046,N_4074);
nor U4320 (N_4320,N_4062,N_4139);
nor U4321 (N_4321,N_4042,N_4088);
or U4322 (N_4322,N_4158,N_4198);
nand U4323 (N_4323,N_4222,N_4033);
nor U4324 (N_4324,N_4172,N_4171);
nor U4325 (N_4325,N_4216,N_4048);
nor U4326 (N_4326,N_4068,N_4189);
nor U4327 (N_4327,N_4151,N_4186);
or U4328 (N_4328,N_4109,N_4080);
xor U4329 (N_4329,N_4094,N_4095);
and U4330 (N_4330,N_4090,N_4235);
nor U4331 (N_4331,N_4085,N_4205);
and U4332 (N_4332,N_4220,N_4057);
nor U4333 (N_4333,N_4000,N_4118);
nor U4334 (N_4334,N_4199,N_4166);
and U4335 (N_4335,N_4123,N_4120);
nor U4336 (N_4336,N_4104,N_4022);
nor U4337 (N_4337,N_4223,N_4236);
or U4338 (N_4338,N_4091,N_4051);
or U4339 (N_4339,N_4136,N_4228);
nor U4340 (N_4340,N_4106,N_4178);
nand U4341 (N_4341,N_4184,N_4229);
nor U4342 (N_4342,N_4240,N_4101);
nor U4343 (N_4343,N_4103,N_4117);
and U4344 (N_4344,N_4247,N_4070);
and U4345 (N_4345,N_4154,N_4116);
xor U4346 (N_4346,N_4167,N_4011);
and U4347 (N_4347,N_4130,N_4129);
or U4348 (N_4348,N_4239,N_4150);
nor U4349 (N_4349,N_4196,N_4013);
nand U4350 (N_4350,N_4050,N_4069);
nor U4351 (N_4351,N_4045,N_4249);
xor U4352 (N_4352,N_4159,N_4016);
nand U4353 (N_4353,N_4081,N_4027);
or U4354 (N_4354,N_4168,N_4026);
nand U4355 (N_4355,N_4093,N_4170);
nor U4356 (N_4356,N_4105,N_4087);
and U4357 (N_4357,N_4208,N_4162);
nand U4358 (N_4358,N_4052,N_4039);
or U4359 (N_4359,N_4086,N_4230);
or U4360 (N_4360,N_4102,N_4157);
nand U4361 (N_4361,N_4007,N_4082);
nand U4362 (N_4362,N_4213,N_4244);
and U4363 (N_4363,N_4098,N_4214);
xnor U4364 (N_4364,N_4134,N_4128);
and U4365 (N_4365,N_4119,N_4173);
xnor U4366 (N_4366,N_4075,N_4242);
xor U4367 (N_4367,N_4182,N_4019);
nor U4368 (N_4368,N_4072,N_4021);
or U4369 (N_4369,N_4034,N_4113);
xor U4370 (N_4370,N_4002,N_4153);
nor U4371 (N_4371,N_4005,N_4131);
and U4372 (N_4372,N_4163,N_4133);
xor U4373 (N_4373,N_4084,N_4224);
nand U4374 (N_4374,N_4030,N_4140);
nand U4375 (N_4375,N_4001,N_4031);
nand U4376 (N_4376,N_4226,N_4112);
nor U4377 (N_4377,N_4191,N_4062);
nand U4378 (N_4378,N_4174,N_4243);
nand U4379 (N_4379,N_4150,N_4066);
or U4380 (N_4380,N_4089,N_4078);
nand U4381 (N_4381,N_4094,N_4006);
nand U4382 (N_4382,N_4086,N_4216);
or U4383 (N_4383,N_4155,N_4168);
xnor U4384 (N_4384,N_4100,N_4062);
nor U4385 (N_4385,N_4154,N_4002);
nor U4386 (N_4386,N_4170,N_4134);
nor U4387 (N_4387,N_4195,N_4063);
nand U4388 (N_4388,N_4148,N_4031);
and U4389 (N_4389,N_4051,N_4020);
and U4390 (N_4390,N_4081,N_4186);
nand U4391 (N_4391,N_4140,N_4158);
xnor U4392 (N_4392,N_4134,N_4183);
and U4393 (N_4393,N_4229,N_4227);
and U4394 (N_4394,N_4057,N_4036);
nor U4395 (N_4395,N_4045,N_4155);
xnor U4396 (N_4396,N_4201,N_4187);
and U4397 (N_4397,N_4073,N_4112);
and U4398 (N_4398,N_4045,N_4037);
or U4399 (N_4399,N_4130,N_4049);
and U4400 (N_4400,N_4126,N_4248);
and U4401 (N_4401,N_4059,N_4044);
xnor U4402 (N_4402,N_4223,N_4116);
nor U4403 (N_4403,N_4042,N_4064);
xor U4404 (N_4404,N_4073,N_4010);
nor U4405 (N_4405,N_4035,N_4165);
or U4406 (N_4406,N_4036,N_4246);
nor U4407 (N_4407,N_4103,N_4220);
and U4408 (N_4408,N_4117,N_4033);
and U4409 (N_4409,N_4000,N_4221);
or U4410 (N_4410,N_4122,N_4200);
and U4411 (N_4411,N_4228,N_4126);
or U4412 (N_4412,N_4053,N_4015);
or U4413 (N_4413,N_4175,N_4241);
nand U4414 (N_4414,N_4058,N_4110);
nand U4415 (N_4415,N_4044,N_4186);
nand U4416 (N_4416,N_4220,N_4009);
and U4417 (N_4417,N_4019,N_4247);
nor U4418 (N_4418,N_4156,N_4048);
xor U4419 (N_4419,N_4128,N_4063);
xnor U4420 (N_4420,N_4022,N_4084);
nand U4421 (N_4421,N_4055,N_4060);
and U4422 (N_4422,N_4047,N_4045);
or U4423 (N_4423,N_4230,N_4241);
xor U4424 (N_4424,N_4234,N_4050);
xor U4425 (N_4425,N_4239,N_4054);
or U4426 (N_4426,N_4076,N_4088);
or U4427 (N_4427,N_4167,N_4201);
and U4428 (N_4428,N_4094,N_4047);
and U4429 (N_4429,N_4210,N_4091);
or U4430 (N_4430,N_4202,N_4078);
nor U4431 (N_4431,N_4176,N_4234);
nor U4432 (N_4432,N_4037,N_4117);
or U4433 (N_4433,N_4114,N_4239);
and U4434 (N_4434,N_4138,N_4099);
and U4435 (N_4435,N_4239,N_4108);
and U4436 (N_4436,N_4101,N_4234);
nor U4437 (N_4437,N_4164,N_4193);
nor U4438 (N_4438,N_4030,N_4219);
xnor U4439 (N_4439,N_4159,N_4109);
nand U4440 (N_4440,N_4122,N_4245);
xnor U4441 (N_4441,N_4054,N_4101);
xor U4442 (N_4442,N_4091,N_4168);
and U4443 (N_4443,N_4153,N_4214);
and U4444 (N_4444,N_4192,N_4066);
and U4445 (N_4445,N_4210,N_4198);
or U4446 (N_4446,N_4245,N_4040);
xor U4447 (N_4447,N_4036,N_4167);
nand U4448 (N_4448,N_4234,N_4074);
nand U4449 (N_4449,N_4002,N_4234);
and U4450 (N_4450,N_4014,N_4198);
or U4451 (N_4451,N_4125,N_4010);
xor U4452 (N_4452,N_4212,N_4186);
xnor U4453 (N_4453,N_4041,N_4151);
nor U4454 (N_4454,N_4070,N_4176);
nor U4455 (N_4455,N_4088,N_4001);
and U4456 (N_4456,N_4134,N_4008);
or U4457 (N_4457,N_4143,N_4217);
nor U4458 (N_4458,N_4086,N_4245);
and U4459 (N_4459,N_4116,N_4100);
or U4460 (N_4460,N_4169,N_4000);
nor U4461 (N_4461,N_4029,N_4083);
and U4462 (N_4462,N_4033,N_4094);
xnor U4463 (N_4463,N_4225,N_4223);
nand U4464 (N_4464,N_4142,N_4071);
xor U4465 (N_4465,N_4228,N_4032);
nand U4466 (N_4466,N_4040,N_4093);
and U4467 (N_4467,N_4211,N_4034);
xor U4468 (N_4468,N_4170,N_4091);
and U4469 (N_4469,N_4080,N_4069);
nand U4470 (N_4470,N_4222,N_4239);
or U4471 (N_4471,N_4203,N_4164);
and U4472 (N_4472,N_4163,N_4218);
and U4473 (N_4473,N_4067,N_4003);
and U4474 (N_4474,N_4204,N_4109);
nor U4475 (N_4475,N_4164,N_4141);
and U4476 (N_4476,N_4200,N_4217);
nor U4477 (N_4477,N_4155,N_4189);
or U4478 (N_4478,N_4193,N_4030);
nand U4479 (N_4479,N_4202,N_4080);
xnor U4480 (N_4480,N_4149,N_4045);
xor U4481 (N_4481,N_4166,N_4206);
nor U4482 (N_4482,N_4058,N_4147);
nor U4483 (N_4483,N_4242,N_4236);
and U4484 (N_4484,N_4035,N_4083);
xor U4485 (N_4485,N_4068,N_4002);
and U4486 (N_4486,N_4245,N_4049);
nor U4487 (N_4487,N_4207,N_4128);
nand U4488 (N_4488,N_4224,N_4214);
xor U4489 (N_4489,N_4071,N_4186);
and U4490 (N_4490,N_4235,N_4039);
nor U4491 (N_4491,N_4040,N_4098);
or U4492 (N_4492,N_4155,N_4094);
xnor U4493 (N_4493,N_4190,N_4052);
nand U4494 (N_4494,N_4198,N_4146);
and U4495 (N_4495,N_4151,N_4241);
or U4496 (N_4496,N_4188,N_4180);
and U4497 (N_4497,N_4230,N_4227);
nor U4498 (N_4498,N_4084,N_4028);
nand U4499 (N_4499,N_4015,N_4075);
or U4500 (N_4500,N_4429,N_4361);
or U4501 (N_4501,N_4489,N_4312);
or U4502 (N_4502,N_4399,N_4390);
nand U4503 (N_4503,N_4292,N_4480);
xor U4504 (N_4504,N_4403,N_4466);
and U4505 (N_4505,N_4263,N_4442);
or U4506 (N_4506,N_4273,N_4449);
xor U4507 (N_4507,N_4290,N_4401);
xnor U4508 (N_4508,N_4421,N_4369);
nor U4509 (N_4509,N_4254,N_4323);
nor U4510 (N_4510,N_4419,N_4345);
nand U4511 (N_4511,N_4357,N_4391);
xnor U4512 (N_4512,N_4294,N_4495);
and U4513 (N_4513,N_4430,N_4383);
nor U4514 (N_4514,N_4309,N_4306);
or U4515 (N_4515,N_4291,N_4415);
nand U4516 (N_4516,N_4253,N_4343);
nor U4517 (N_4517,N_4439,N_4258);
xnor U4518 (N_4518,N_4493,N_4264);
or U4519 (N_4519,N_4420,N_4285);
and U4520 (N_4520,N_4423,N_4293);
nand U4521 (N_4521,N_4494,N_4354);
xnor U4522 (N_4522,N_4307,N_4365);
nor U4523 (N_4523,N_4251,N_4479);
xnor U4524 (N_4524,N_4454,N_4470);
xnor U4525 (N_4525,N_4404,N_4327);
nand U4526 (N_4526,N_4339,N_4431);
or U4527 (N_4527,N_4485,N_4368);
xor U4528 (N_4528,N_4341,N_4378);
nor U4529 (N_4529,N_4408,N_4372);
or U4530 (N_4530,N_4370,N_4464);
and U4531 (N_4531,N_4358,N_4409);
or U4532 (N_4532,N_4407,N_4487);
xnor U4533 (N_4533,N_4392,N_4475);
nor U4534 (N_4534,N_4481,N_4299);
and U4535 (N_4535,N_4266,N_4458);
xnor U4536 (N_4536,N_4308,N_4333);
or U4537 (N_4537,N_4387,N_4396);
or U4538 (N_4538,N_4256,N_4482);
nor U4539 (N_4539,N_4313,N_4448);
nor U4540 (N_4540,N_4355,N_4320);
nand U4541 (N_4541,N_4305,N_4400);
nor U4542 (N_4542,N_4297,N_4255);
or U4543 (N_4543,N_4433,N_4463);
or U4544 (N_4544,N_4301,N_4283);
or U4545 (N_4545,N_4321,N_4456);
xnor U4546 (N_4546,N_4284,N_4270);
or U4547 (N_4547,N_4328,N_4498);
or U4548 (N_4548,N_4318,N_4418);
nand U4549 (N_4549,N_4286,N_4348);
xnor U4550 (N_4550,N_4478,N_4324);
nor U4551 (N_4551,N_4296,N_4440);
or U4552 (N_4552,N_4278,N_4451);
xor U4553 (N_4553,N_4468,N_4304);
and U4554 (N_4554,N_4269,N_4364);
nand U4555 (N_4555,N_4337,N_4311);
or U4556 (N_4556,N_4406,N_4484);
xor U4557 (N_4557,N_4434,N_4385);
xnor U4558 (N_4558,N_4252,N_4259);
or U4559 (N_4559,N_4257,N_4474);
or U4560 (N_4560,N_4362,N_4267);
nor U4561 (N_4561,N_4347,N_4332);
and U4562 (N_4562,N_4422,N_4492);
nor U4563 (N_4563,N_4367,N_4444);
and U4564 (N_4564,N_4336,N_4386);
nand U4565 (N_4565,N_4435,N_4426);
nor U4566 (N_4566,N_4317,N_4402);
nor U4567 (N_4567,N_4413,N_4486);
nor U4568 (N_4568,N_4425,N_4340);
and U4569 (N_4569,N_4374,N_4289);
nor U4570 (N_4570,N_4462,N_4282);
or U4571 (N_4571,N_4315,N_4428);
or U4572 (N_4572,N_4325,N_4342);
nand U4573 (N_4573,N_4471,N_4265);
nand U4574 (N_4574,N_4295,N_4310);
nor U4575 (N_4575,N_4319,N_4376);
xnor U4576 (N_4576,N_4352,N_4268);
or U4577 (N_4577,N_4344,N_4443);
nand U4578 (N_4578,N_4488,N_4395);
nand U4579 (N_4579,N_4334,N_4473);
and U4580 (N_4580,N_4363,N_4329);
nor U4581 (N_4581,N_4350,N_4459);
xor U4582 (N_4582,N_4465,N_4398);
nor U4583 (N_4583,N_4445,N_4476);
or U4584 (N_4584,N_4436,N_4346);
and U4585 (N_4585,N_4490,N_4497);
nand U4586 (N_4586,N_4394,N_4316);
nand U4587 (N_4587,N_4447,N_4349);
xor U4588 (N_4588,N_4359,N_4427);
and U4589 (N_4589,N_4446,N_4483);
and U4590 (N_4590,N_4262,N_4300);
xnor U4591 (N_4591,N_4441,N_4393);
nand U4592 (N_4592,N_4450,N_4380);
or U4593 (N_4593,N_4330,N_4360);
nor U4594 (N_4594,N_4275,N_4460);
and U4595 (N_4595,N_4303,N_4260);
and U4596 (N_4596,N_4280,N_4276);
or U4597 (N_4597,N_4371,N_4277);
and U4598 (N_4598,N_4417,N_4373);
xor U4599 (N_4599,N_4437,N_4331);
nor U4600 (N_4600,N_4377,N_4353);
xor U4601 (N_4601,N_4261,N_4432);
xnor U4602 (N_4602,N_4410,N_4414);
or U4603 (N_4603,N_4384,N_4298);
xor U4604 (N_4604,N_4379,N_4499);
xnor U4605 (N_4605,N_4287,N_4416);
and U4606 (N_4606,N_4338,N_4438);
nor U4607 (N_4607,N_4351,N_4457);
nor U4608 (N_4608,N_4335,N_4455);
nor U4609 (N_4609,N_4389,N_4412);
and U4610 (N_4610,N_4477,N_4272);
nor U4611 (N_4611,N_4366,N_4469);
or U4612 (N_4612,N_4397,N_4381);
and U4613 (N_4613,N_4461,N_4382);
nand U4614 (N_4614,N_4411,N_4288);
nand U4615 (N_4615,N_4274,N_4271);
and U4616 (N_4616,N_4314,N_4375);
nand U4617 (N_4617,N_4472,N_4302);
or U4618 (N_4618,N_4424,N_4491);
xnor U4619 (N_4619,N_4467,N_4452);
nor U4620 (N_4620,N_4322,N_4279);
and U4621 (N_4621,N_4496,N_4356);
nor U4622 (N_4622,N_4405,N_4281);
or U4623 (N_4623,N_4326,N_4250);
and U4624 (N_4624,N_4388,N_4453);
nand U4625 (N_4625,N_4476,N_4322);
nand U4626 (N_4626,N_4271,N_4362);
or U4627 (N_4627,N_4355,N_4357);
nor U4628 (N_4628,N_4388,N_4420);
xor U4629 (N_4629,N_4495,N_4394);
nor U4630 (N_4630,N_4402,N_4454);
nor U4631 (N_4631,N_4334,N_4437);
xnor U4632 (N_4632,N_4470,N_4429);
xor U4633 (N_4633,N_4303,N_4320);
nor U4634 (N_4634,N_4340,N_4254);
nand U4635 (N_4635,N_4254,N_4296);
xnor U4636 (N_4636,N_4400,N_4413);
xnor U4637 (N_4637,N_4426,N_4367);
nor U4638 (N_4638,N_4388,N_4347);
xor U4639 (N_4639,N_4410,N_4256);
nor U4640 (N_4640,N_4379,N_4474);
xor U4641 (N_4641,N_4322,N_4444);
and U4642 (N_4642,N_4383,N_4489);
xor U4643 (N_4643,N_4460,N_4320);
nand U4644 (N_4644,N_4363,N_4487);
xor U4645 (N_4645,N_4258,N_4373);
xor U4646 (N_4646,N_4304,N_4374);
nand U4647 (N_4647,N_4380,N_4253);
or U4648 (N_4648,N_4256,N_4291);
xnor U4649 (N_4649,N_4397,N_4377);
or U4650 (N_4650,N_4403,N_4327);
and U4651 (N_4651,N_4442,N_4324);
nor U4652 (N_4652,N_4383,N_4300);
nand U4653 (N_4653,N_4314,N_4457);
and U4654 (N_4654,N_4281,N_4412);
or U4655 (N_4655,N_4318,N_4456);
and U4656 (N_4656,N_4264,N_4266);
and U4657 (N_4657,N_4402,N_4458);
nand U4658 (N_4658,N_4468,N_4339);
nand U4659 (N_4659,N_4354,N_4488);
xor U4660 (N_4660,N_4275,N_4312);
and U4661 (N_4661,N_4410,N_4406);
nor U4662 (N_4662,N_4358,N_4277);
nor U4663 (N_4663,N_4422,N_4357);
or U4664 (N_4664,N_4353,N_4274);
or U4665 (N_4665,N_4306,N_4388);
and U4666 (N_4666,N_4365,N_4415);
xor U4667 (N_4667,N_4408,N_4407);
and U4668 (N_4668,N_4352,N_4403);
xor U4669 (N_4669,N_4337,N_4264);
or U4670 (N_4670,N_4320,N_4439);
and U4671 (N_4671,N_4257,N_4260);
and U4672 (N_4672,N_4299,N_4451);
xnor U4673 (N_4673,N_4262,N_4383);
nor U4674 (N_4674,N_4380,N_4471);
and U4675 (N_4675,N_4422,N_4425);
or U4676 (N_4676,N_4402,N_4330);
xnor U4677 (N_4677,N_4320,N_4312);
and U4678 (N_4678,N_4278,N_4468);
and U4679 (N_4679,N_4265,N_4441);
nor U4680 (N_4680,N_4495,N_4291);
and U4681 (N_4681,N_4375,N_4457);
and U4682 (N_4682,N_4374,N_4290);
or U4683 (N_4683,N_4410,N_4259);
and U4684 (N_4684,N_4257,N_4334);
nand U4685 (N_4685,N_4329,N_4320);
nor U4686 (N_4686,N_4470,N_4338);
or U4687 (N_4687,N_4358,N_4372);
nor U4688 (N_4688,N_4330,N_4317);
nor U4689 (N_4689,N_4470,N_4335);
nand U4690 (N_4690,N_4272,N_4357);
and U4691 (N_4691,N_4312,N_4311);
or U4692 (N_4692,N_4335,N_4485);
and U4693 (N_4693,N_4261,N_4328);
nor U4694 (N_4694,N_4353,N_4283);
nand U4695 (N_4695,N_4400,N_4353);
nand U4696 (N_4696,N_4320,N_4282);
nor U4697 (N_4697,N_4399,N_4317);
and U4698 (N_4698,N_4498,N_4471);
or U4699 (N_4699,N_4453,N_4317);
nor U4700 (N_4700,N_4361,N_4368);
xnor U4701 (N_4701,N_4466,N_4462);
nand U4702 (N_4702,N_4434,N_4420);
or U4703 (N_4703,N_4404,N_4448);
and U4704 (N_4704,N_4452,N_4458);
nor U4705 (N_4705,N_4356,N_4413);
and U4706 (N_4706,N_4488,N_4343);
xnor U4707 (N_4707,N_4461,N_4451);
nand U4708 (N_4708,N_4446,N_4470);
nor U4709 (N_4709,N_4266,N_4341);
xnor U4710 (N_4710,N_4265,N_4253);
or U4711 (N_4711,N_4436,N_4428);
or U4712 (N_4712,N_4477,N_4294);
and U4713 (N_4713,N_4464,N_4346);
or U4714 (N_4714,N_4260,N_4280);
or U4715 (N_4715,N_4440,N_4307);
xnor U4716 (N_4716,N_4254,N_4436);
nand U4717 (N_4717,N_4407,N_4348);
nor U4718 (N_4718,N_4466,N_4273);
or U4719 (N_4719,N_4391,N_4351);
or U4720 (N_4720,N_4469,N_4421);
xor U4721 (N_4721,N_4405,N_4344);
nand U4722 (N_4722,N_4329,N_4365);
xor U4723 (N_4723,N_4330,N_4462);
nor U4724 (N_4724,N_4405,N_4430);
nand U4725 (N_4725,N_4478,N_4382);
and U4726 (N_4726,N_4430,N_4340);
and U4727 (N_4727,N_4278,N_4410);
nor U4728 (N_4728,N_4345,N_4261);
nand U4729 (N_4729,N_4302,N_4283);
or U4730 (N_4730,N_4282,N_4461);
xnor U4731 (N_4731,N_4442,N_4299);
nand U4732 (N_4732,N_4321,N_4449);
nor U4733 (N_4733,N_4250,N_4343);
xor U4734 (N_4734,N_4492,N_4351);
xnor U4735 (N_4735,N_4422,N_4377);
nor U4736 (N_4736,N_4430,N_4325);
or U4737 (N_4737,N_4387,N_4391);
nor U4738 (N_4738,N_4358,N_4414);
and U4739 (N_4739,N_4484,N_4414);
nor U4740 (N_4740,N_4294,N_4485);
xnor U4741 (N_4741,N_4472,N_4252);
and U4742 (N_4742,N_4289,N_4342);
nand U4743 (N_4743,N_4485,N_4493);
and U4744 (N_4744,N_4392,N_4423);
and U4745 (N_4745,N_4342,N_4410);
or U4746 (N_4746,N_4316,N_4254);
or U4747 (N_4747,N_4378,N_4262);
and U4748 (N_4748,N_4432,N_4313);
xnor U4749 (N_4749,N_4269,N_4455);
xnor U4750 (N_4750,N_4703,N_4666);
xor U4751 (N_4751,N_4532,N_4739);
nor U4752 (N_4752,N_4691,N_4597);
xnor U4753 (N_4753,N_4717,N_4573);
nor U4754 (N_4754,N_4614,N_4700);
and U4755 (N_4755,N_4671,N_4587);
xnor U4756 (N_4756,N_4540,N_4521);
or U4757 (N_4757,N_4629,N_4694);
or U4758 (N_4758,N_4716,N_4543);
or U4759 (N_4759,N_4569,N_4565);
nand U4760 (N_4760,N_4509,N_4709);
and U4761 (N_4761,N_4680,N_4648);
nor U4762 (N_4762,N_4737,N_4743);
and U4763 (N_4763,N_4676,N_4530);
nand U4764 (N_4764,N_4539,N_4708);
xor U4765 (N_4765,N_4675,N_4502);
xnor U4766 (N_4766,N_4704,N_4622);
xor U4767 (N_4767,N_4541,N_4625);
and U4768 (N_4768,N_4747,N_4658);
and U4769 (N_4769,N_4729,N_4731);
nor U4770 (N_4770,N_4600,N_4672);
xnor U4771 (N_4771,N_4613,N_4715);
and U4772 (N_4772,N_4526,N_4511);
nand U4773 (N_4773,N_4746,N_4713);
nand U4774 (N_4774,N_4665,N_4711);
nand U4775 (N_4775,N_4523,N_4664);
xor U4776 (N_4776,N_4542,N_4536);
nand U4777 (N_4777,N_4682,N_4669);
xor U4778 (N_4778,N_4619,N_4514);
nand U4779 (N_4779,N_4673,N_4590);
xor U4780 (N_4780,N_4533,N_4645);
or U4781 (N_4781,N_4566,N_4524);
and U4782 (N_4782,N_4531,N_4537);
and U4783 (N_4783,N_4544,N_4608);
nand U4784 (N_4784,N_4688,N_4618);
xor U4785 (N_4785,N_4630,N_4535);
and U4786 (N_4786,N_4506,N_4635);
or U4787 (N_4787,N_4563,N_4670);
nor U4788 (N_4788,N_4574,N_4726);
nor U4789 (N_4789,N_4576,N_4609);
nand U4790 (N_4790,N_4545,N_4702);
nand U4791 (N_4791,N_4685,N_4607);
or U4792 (N_4792,N_4741,N_4561);
xor U4793 (N_4793,N_4518,N_4722);
nand U4794 (N_4794,N_4549,N_4560);
or U4795 (N_4795,N_4616,N_4571);
and U4796 (N_4796,N_4749,N_4677);
nand U4797 (N_4797,N_4697,N_4686);
and U4798 (N_4798,N_4744,N_4695);
and U4799 (N_4799,N_4552,N_4551);
or U4800 (N_4800,N_4628,N_4718);
xnor U4801 (N_4801,N_4554,N_4657);
nand U4802 (N_4802,N_4605,N_4577);
nand U4803 (N_4803,N_4662,N_4647);
or U4804 (N_4804,N_4620,N_4707);
or U4805 (N_4805,N_4701,N_4712);
xnor U4806 (N_4806,N_4699,N_4516);
and U4807 (N_4807,N_4723,N_4719);
or U4808 (N_4808,N_4710,N_4683);
or U4809 (N_4809,N_4568,N_4681);
nor U4810 (N_4810,N_4621,N_4519);
and U4811 (N_4811,N_4660,N_4599);
xor U4812 (N_4812,N_4646,N_4558);
or U4813 (N_4813,N_4734,N_4684);
or U4814 (N_4814,N_4730,N_4627);
nand U4815 (N_4815,N_4735,N_4617);
or U4816 (N_4816,N_4725,N_4546);
xor U4817 (N_4817,N_4742,N_4556);
nor U4818 (N_4818,N_4594,N_4606);
and U4819 (N_4819,N_4693,N_4583);
or U4820 (N_4820,N_4668,N_4650);
nand U4821 (N_4821,N_4612,N_4529);
nand U4822 (N_4822,N_4637,N_4557);
xor U4823 (N_4823,N_4689,N_4534);
xnor U4824 (N_4824,N_4632,N_4570);
xor U4825 (N_4825,N_4667,N_4538);
or U4826 (N_4826,N_4692,N_4522);
and U4827 (N_4827,N_4659,N_4639);
and U4828 (N_4828,N_4624,N_4596);
nor U4829 (N_4829,N_4508,N_4513);
nand U4830 (N_4830,N_4733,N_4728);
or U4831 (N_4831,N_4661,N_4575);
and U4832 (N_4832,N_4643,N_4732);
nor U4833 (N_4833,N_4698,N_4527);
and U4834 (N_4834,N_4520,N_4591);
nor U4835 (N_4835,N_4623,N_4525);
and U4836 (N_4836,N_4602,N_4548);
and U4837 (N_4837,N_4515,N_4553);
and U4838 (N_4838,N_4564,N_4640);
xor U4839 (N_4839,N_4585,N_4651);
nand U4840 (N_4840,N_4567,N_4679);
nand U4841 (N_4841,N_4690,N_4641);
and U4842 (N_4842,N_4696,N_4510);
nand U4843 (N_4843,N_4503,N_4736);
and U4844 (N_4844,N_4721,N_4500);
nand U4845 (N_4845,N_4572,N_4663);
and U4846 (N_4846,N_4626,N_4604);
nand U4847 (N_4847,N_4582,N_4595);
xor U4848 (N_4848,N_4652,N_4738);
and U4849 (N_4849,N_4745,N_4610);
and U4850 (N_4850,N_4611,N_4517);
nand U4851 (N_4851,N_4588,N_4649);
xor U4852 (N_4852,N_4727,N_4580);
xnor U4853 (N_4853,N_4592,N_4501);
xor U4854 (N_4854,N_4547,N_4636);
nand U4855 (N_4855,N_4528,N_4642);
and U4856 (N_4856,N_4579,N_4714);
nand U4857 (N_4857,N_4720,N_4705);
xor U4858 (N_4858,N_4601,N_4654);
nor U4859 (N_4859,N_4593,N_4512);
and U4860 (N_4860,N_4724,N_4507);
and U4861 (N_4861,N_4559,N_4578);
and U4862 (N_4862,N_4634,N_4504);
nor U4863 (N_4863,N_4740,N_4589);
and U4864 (N_4864,N_4603,N_4653);
nand U4865 (N_4865,N_4550,N_4748);
xnor U4866 (N_4866,N_4555,N_4633);
xnor U4867 (N_4867,N_4631,N_4638);
nand U4868 (N_4868,N_4505,N_4562);
and U4869 (N_4869,N_4581,N_4674);
xnor U4870 (N_4870,N_4678,N_4656);
nand U4871 (N_4871,N_4644,N_4706);
nand U4872 (N_4872,N_4586,N_4687);
xor U4873 (N_4873,N_4598,N_4655);
nor U4874 (N_4874,N_4615,N_4584);
nor U4875 (N_4875,N_4603,N_4549);
nor U4876 (N_4876,N_4542,N_4583);
and U4877 (N_4877,N_4570,N_4720);
and U4878 (N_4878,N_4613,N_4704);
xor U4879 (N_4879,N_4556,N_4603);
xor U4880 (N_4880,N_4571,N_4559);
or U4881 (N_4881,N_4530,N_4613);
and U4882 (N_4882,N_4540,N_4716);
and U4883 (N_4883,N_4643,N_4699);
xor U4884 (N_4884,N_4721,N_4743);
nor U4885 (N_4885,N_4549,N_4677);
xor U4886 (N_4886,N_4662,N_4674);
and U4887 (N_4887,N_4696,N_4525);
nand U4888 (N_4888,N_4659,N_4557);
or U4889 (N_4889,N_4527,N_4625);
xnor U4890 (N_4890,N_4570,N_4599);
nand U4891 (N_4891,N_4580,N_4749);
nor U4892 (N_4892,N_4542,N_4655);
xor U4893 (N_4893,N_4630,N_4621);
or U4894 (N_4894,N_4685,N_4638);
nor U4895 (N_4895,N_4665,N_4620);
nor U4896 (N_4896,N_4583,N_4551);
and U4897 (N_4897,N_4739,N_4658);
nor U4898 (N_4898,N_4514,N_4733);
nor U4899 (N_4899,N_4554,N_4568);
or U4900 (N_4900,N_4562,N_4729);
or U4901 (N_4901,N_4718,N_4721);
nor U4902 (N_4902,N_4675,N_4627);
nand U4903 (N_4903,N_4580,N_4544);
nand U4904 (N_4904,N_4747,N_4554);
and U4905 (N_4905,N_4500,N_4524);
nand U4906 (N_4906,N_4685,N_4695);
and U4907 (N_4907,N_4503,N_4740);
nand U4908 (N_4908,N_4503,N_4643);
or U4909 (N_4909,N_4593,N_4737);
and U4910 (N_4910,N_4586,N_4562);
or U4911 (N_4911,N_4677,N_4678);
and U4912 (N_4912,N_4520,N_4705);
xor U4913 (N_4913,N_4621,N_4728);
and U4914 (N_4914,N_4725,N_4691);
or U4915 (N_4915,N_4632,N_4549);
nor U4916 (N_4916,N_4668,N_4517);
or U4917 (N_4917,N_4582,N_4594);
nand U4918 (N_4918,N_4510,N_4695);
or U4919 (N_4919,N_4530,N_4555);
or U4920 (N_4920,N_4664,N_4737);
or U4921 (N_4921,N_4663,N_4571);
nor U4922 (N_4922,N_4674,N_4584);
nor U4923 (N_4923,N_4624,N_4620);
and U4924 (N_4924,N_4676,N_4510);
xnor U4925 (N_4925,N_4716,N_4732);
and U4926 (N_4926,N_4602,N_4545);
nor U4927 (N_4927,N_4571,N_4611);
xor U4928 (N_4928,N_4713,N_4693);
nor U4929 (N_4929,N_4659,N_4743);
and U4930 (N_4930,N_4681,N_4544);
nor U4931 (N_4931,N_4735,N_4565);
and U4932 (N_4932,N_4641,N_4639);
nand U4933 (N_4933,N_4638,N_4661);
or U4934 (N_4934,N_4544,N_4529);
or U4935 (N_4935,N_4690,N_4542);
or U4936 (N_4936,N_4537,N_4593);
and U4937 (N_4937,N_4741,N_4564);
xnor U4938 (N_4938,N_4640,N_4606);
or U4939 (N_4939,N_4685,N_4599);
nand U4940 (N_4940,N_4541,N_4682);
or U4941 (N_4941,N_4745,N_4698);
and U4942 (N_4942,N_4598,N_4662);
xnor U4943 (N_4943,N_4551,N_4604);
and U4944 (N_4944,N_4631,N_4562);
xor U4945 (N_4945,N_4620,N_4677);
xnor U4946 (N_4946,N_4593,N_4708);
and U4947 (N_4947,N_4611,N_4555);
or U4948 (N_4948,N_4654,N_4505);
or U4949 (N_4949,N_4507,N_4662);
xor U4950 (N_4950,N_4581,N_4625);
xnor U4951 (N_4951,N_4640,N_4747);
nor U4952 (N_4952,N_4715,N_4724);
nand U4953 (N_4953,N_4699,N_4738);
nor U4954 (N_4954,N_4671,N_4682);
nor U4955 (N_4955,N_4571,N_4657);
xor U4956 (N_4956,N_4640,N_4522);
xnor U4957 (N_4957,N_4513,N_4684);
nand U4958 (N_4958,N_4651,N_4598);
nor U4959 (N_4959,N_4587,N_4711);
xnor U4960 (N_4960,N_4601,N_4589);
nor U4961 (N_4961,N_4644,N_4511);
xor U4962 (N_4962,N_4514,N_4627);
nand U4963 (N_4963,N_4661,N_4603);
xor U4964 (N_4964,N_4665,N_4732);
and U4965 (N_4965,N_4704,N_4682);
nor U4966 (N_4966,N_4520,N_4603);
xor U4967 (N_4967,N_4649,N_4716);
and U4968 (N_4968,N_4704,N_4511);
and U4969 (N_4969,N_4505,N_4742);
nor U4970 (N_4970,N_4673,N_4655);
nand U4971 (N_4971,N_4702,N_4583);
xnor U4972 (N_4972,N_4503,N_4589);
xor U4973 (N_4973,N_4564,N_4541);
xnor U4974 (N_4974,N_4584,N_4566);
or U4975 (N_4975,N_4626,N_4713);
or U4976 (N_4976,N_4680,N_4569);
nand U4977 (N_4977,N_4679,N_4634);
or U4978 (N_4978,N_4600,N_4541);
nor U4979 (N_4979,N_4710,N_4733);
nor U4980 (N_4980,N_4719,N_4604);
nor U4981 (N_4981,N_4522,N_4547);
or U4982 (N_4982,N_4743,N_4720);
nand U4983 (N_4983,N_4640,N_4745);
and U4984 (N_4984,N_4722,N_4539);
nand U4985 (N_4985,N_4666,N_4617);
nor U4986 (N_4986,N_4529,N_4548);
nor U4987 (N_4987,N_4519,N_4684);
and U4988 (N_4988,N_4709,N_4585);
and U4989 (N_4989,N_4717,N_4607);
and U4990 (N_4990,N_4629,N_4647);
xnor U4991 (N_4991,N_4501,N_4585);
and U4992 (N_4992,N_4618,N_4624);
nand U4993 (N_4993,N_4511,N_4699);
nor U4994 (N_4994,N_4573,N_4535);
nand U4995 (N_4995,N_4680,N_4687);
xor U4996 (N_4996,N_4747,N_4527);
nand U4997 (N_4997,N_4696,N_4658);
xor U4998 (N_4998,N_4676,N_4555);
and U4999 (N_4999,N_4745,N_4676);
nor U5000 (N_5000,N_4852,N_4797);
nor U5001 (N_5001,N_4764,N_4891);
xor U5002 (N_5002,N_4854,N_4816);
and U5003 (N_5003,N_4970,N_4840);
xor U5004 (N_5004,N_4796,N_4956);
or U5005 (N_5005,N_4899,N_4998);
nand U5006 (N_5006,N_4974,N_4966);
or U5007 (N_5007,N_4777,N_4980);
xor U5008 (N_5008,N_4786,N_4909);
xnor U5009 (N_5009,N_4914,N_4976);
nor U5010 (N_5010,N_4948,N_4905);
nand U5011 (N_5011,N_4911,N_4856);
and U5012 (N_5012,N_4865,N_4757);
nand U5013 (N_5013,N_4935,N_4947);
nor U5014 (N_5014,N_4773,N_4874);
or U5015 (N_5015,N_4879,N_4822);
nor U5016 (N_5016,N_4754,N_4996);
nor U5017 (N_5017,N_4919,N_4913);
or U5018 (N_5018,N_4812,N_4761);
or U5019 (N_5019,N_4983,N_4807);
and U5020 (N_5020,N_4964,N_4861);
nand U5021 (N_5021,N_4760,N_4779);
nor U5022 (N_5022,N_4939,N_4782);
and U5023 (N_5023,N_4982,N_4994);
xnor U5024 (N_5024,N_4768,N_4863);
and U5025 (N_5025,N_4787,N_4804);
and U5026 (N_5026,N_4850,N_4907);
or U5027 (N_5027,N_4972,N_4938);
nand U5028 (N_5028,N_4903,N_4927);
nor U5029 (N_5029,N_4835,N_4892);
nor U5030 (N_5030,N_4873,N_4770);
nor U5031 (N_5031,N_4987,N_4924);
nor U5032 (N_5032,N_4989,N_4886);
or U5033 (N_5033,N_4851,N_4900);
and U5034 (N_5034,N_4944,N_4951);
and U5035 (N_5035,N_4867,N_4817);
nand U5036 (N_5036,N_4933,N_4876);
or U5037 (N_5037,N_4803,N_4834);
xor U5038 (N_5038,N_4908,N_4792);
nand U5039 (N_5039,N_4890,N_4884);
and U5040 (N_5040,N_4862,N_4774);
nand U5041 (N_5041,N_4842,N_4758);
nand U5042 (N_5042,N_4928,N_4898);
or U5043 (N_5043,N_4940,N_4853);
or U5044 (N_5044,N_4870,N_4753);
xnor U5045 (N_5045,N_4778,N_4950);
nor U5046 (N_5046,N_4751,N_4963);
or U5047 (N_5047,N_4820,N_4794);
xor U5048 (N_5048,N_4801,N_4789);
nor U5049 (N_5049,N_4859,N_4755);
or U5050 (N_5050,N_4946,N_4825);
or U5051 (N_5051,N_4831,N_4915);
xor U5052 (N_5052,N_4783,N_4941);
nand U5053 (N_5053,N_4858,N_4769);
nor U5054 (N_5054,N_4889,N_4750);
or U5055 (N_5055,N_4847,N_4893);
and U5056 (N_5056,N_4772,N_4866);
nand U5057 (N_5057,N_4781,N_4988);
nor U5058 (N_5058,N_4918,N_4979);
xor U5059 (N_5059,N_4828,N_4780);
or U5060 (N_5060,N_4916,N_4930);
xnor U5061 (N_5061,N_4836,N_4810);
and U5062 (N_5062,N_4910,N_4855);
xnor U5063 (N_5063,N_4776,N_4981);
nor U5064 (N_5064,N_4882,N_4798);
or U5065 (N_5065,N_4881,N_4971);
nand U5066 (N_5066,N_4895,N_4826);
or U5067 (N_5067,N_4906,N_4921);
xnor U5068 (N_5068,N_4997,N_4857);
or U5069 (N_5069,N_4992,N_4811);
xnor U5070 (N_5070,N_4880,N_4894);
and U5071 (N_5071,N_4993,N_4759);
or U5072 (N_5072,N_4845,N_4942);
nor U5073 (N_5073,N_4917,N_4849);
and U5074 (N_5074,N_4766,N_4985);
nor U5075 (N_5075,N_4967,N_4958);
nor U5076 (N_5076,N_4809,N_4814);
nor U5077 (N_5077,N_4923,N_4756);
nor U5078 (N_5078,N_4832,N_4922);
and U5079 (N_5079,N_4969,N_4827);
and U5080 (N_5080,N_4975,N_4815);
nor U5081 (N_5081,N_4839,N_4959);
or U5082 (N_5082,N_4868,N_4788);
xor U5083 (N_5083,N_4945,N_4878);
nor U5084 (N_5084,N_4830,N_4841);
or U5085 (N_5085,N_4800,N_4833);
or U5086 (N_5086,N_4965,N_4912);
xor U5087 (N_5087,N_4937,N_4837);
xnor U5088 (N_5088,N_4901,N_4795);
xnor U5089 (N_5089,N_4843,N_4805);
xor U5090 (N_5090,N_4821,N_4943);
xnor U5091 (N_5091,N_4936,N_4799);
nand U5092 (N_5092,N_4883,N_4888);
nand U5093 (N_5093,N_4869,N_4860);
and U5094 (N_5094,N_4961,N_4990);
nand U5095 (N_5095,N_4864,N_4818);
nand U5096 (N_5096,N_4877,N_4875);
nor U5097 (N_5097,N_4791,N_4765);
nand U5098 (N_5098,N_4806,N_4931);
nor U5099 (N_5099,N_4885,N_4986);
nor U5100 (N_5100,N_4793,N_4784);
or U5101 (N_5101,N_4926,N_4819);
nor U5102 (N_5102,N_4952,N_4846);
nand U5103 (N_5103,N_4844,N_4872);
nand U5104 (N_5104,N_4762,N_4897);
nor U5105 (N_5105,N_4932,N_4999);
xnor U5106 (N_5106,N_4978,N_4763);
xnor U5107 (N_5107,N_4968,N_4813);
nand U5108 (N_5108,N_4848,N_4871);
or U5109 (N_5109,N_4902,N_4995);
xor U5110 (N_5110,N_4954,N_4949);
and U5111 (N_5111,N_4790,N_4808);
and U5112 (N_5112,N_4838,N_4896);
xor U5113 (N_5113,N_4962,N_4991);
or U5114 (N_5114,N_4955,N_4960);
xor U5115 (N_5115,N_4785,N_4752);
or U5116 (N_5116,N_4920,N_4977);
and U5117 (N_5117,N_4771,N_4904);
nor U5118 (N_5118,N_4824,N_4973);
or U5119 (N_5119,N_4775,N_4984);
xor U5120 (N_5120,N_4929,N_4829);
or U5121 (N_5121,N_4767,N_4925);
or U5122 (N_5122,N_4953,N_4934);
xor U5123 (N_5123,N_4823,N_4887);
nor U5124 (N_5124,N_4802,N_4957);
and U5125 (N_5125,N_4776,N_4982);
xor U5126 (N_5126,N_4897,N_4768);
or U5127 (N_5127,N_4846,N_4826);
nand U5128 (N_5128,N_4996,N_4761);
nor U5129 (N_5129,N_4826,N_4919);
nor U5130 (N_5130,N_4794,N_4915);
nand U5131 (N_5131,N_4802,N_4900);
and U5132 (N_5132,N_4774,N_4832);
xor U5133 (N_5133,N_4964,N_4802);
nand U5134 (N_5134,N_4779,N_4987);
nor U5135 (N_5135,N_4938,N_4947);
nand U5136 (N_5136,N_4750,N_4877);
nand U5137 (N_5137,N_4943,N_4843);
and U5138 (N_5138,N_4962,N_4920);
nand U5139 (N_5139,N_4818,N_4838);
nand U5140 (N_5140,N_4907,N_4756);
xor U5141 (N_5141,N_4761,N_4765);
nand U5142 (N_5142,N_4864,N_4930);
nor U5143 (N_5143,N_4981,N_4844);
nor U5144 (N_5144,N_4805,N_4999);
nand U5145 (N_5145,N_4972,N_4873);
or U5146 (N_5146,N_4967,N_4926);
nor U5147 (N_5147,N_4964,N_4917);
or U5148 (N_5148,N_4888,N_4907);
and U5149 (N_5149,N_4973,N_4842);
or U5150 (N_5150,N_4905,N_4755);
xor U5151 (N_5151,N_4846,N_4753);
or U5152 (N_5152,N_4998,N_4902);
or U5153 (N_5153,N_4998,N_4856);
and U5154 (N_5154,N_4998,N_4822);
and U5155 (N_5155,N_4975,N_4808);
nand U5156 (N_5156,N_4955,N_4779);
nand U5157 (N_5157,N_4964,N_4898);
and U5158 (N_5158,N_4953,N_4782);
xor U5159 (N_5159,N_4970,N_4772);
nor U5160 (N_5160,N_4854,N_4928);
or U5161 (N_5161,N_4766,N_4944);
xnor U5162 (N_5162,N_4750,N_4897);
and U5163 (N_5163,N_4822,N_4767);
nor U5164 (N_5164,N_4901,N_4905);
nor U5165 (N_5165,N_4926,N_4843);
nor U5166 (N_5166,N_4820,N_4968);
nor U5167 (N_5167,N_4778,N_4815);
or U5168 (N_5168,N_4907,N_4806);
or U5169 (N_5169,N_4830,N_4998);
or U5170 (N_5170,N_4806,N_4942);
or U5171 (N_5171,N_4970,N_4961);
nor U5172 (N_5172,N_4963,N_4875);
nand U5173 (N_5173,N_4923,N_4853);
nor U5174 (N_5174,N_4999,N_4900);
and U5175 (N_5175,N_4894,N_4814);
and U5176 (N_5176,N_4939,N_4977);
and U5177 (N_5177,N_4826,N_4953);
nand U5178 (N_5178,N_4940,N_4947);
xnor U5179 (N_5179,N_4767,N_4986);
nor U5180 (N_5180,N_4778,N_4951);
nand U5181 (N_5181,N_4756,N_4899);
xor U5182 (N_5182,N_4887,N_4826);
or U5183 (N_5183,N_4755,N_4993);
nor U5184 (N_5184,N_4879,N_4767);
nand U5185 (N_5185,N_4877,N_4820);
or U5186 (N_5186,N_4804,N_4987);
and U5187 (N_5187,N_4882,N_4850);
and U5188 (N_5188,N_4978,N_4839);
nand U5189 (N_5189,N_4971,N_4875);
nand U5190 (N_5190,N_4937,N_4868);
xnor U5191 (N_5191,N_4882,N_4941);
nor U5192 (N_5192,N_4983,N_4948);
xor U5193 (N_5193,N_4776,N_4927);
or U5194 (N_5194,N_4817,N_4787);
xor U5195 (N_5195,N_4996,N_4888);
and U5196 (N_5196,N_4955,N_4939);
xnor U5197 (N_5197,N_4915,N_4912);
and U5198 (N_5198,N_4871,N_4847);
and U5199 (N_5199,N_4834,N_4950);
and U5200 (N_5200,N_4824,N_4965);
nand U5201 (N_5201,N_4843,N_4928);
nor U5202 (N_5202,N_4901,N_4780);
nand U5203 (N_5203,N_4985,N_4767);
or U5204 (N_5204,N_4949,N_4993);
and U5205 (N_5205,N_4920,N_4837);
and U5206 (N_5206,N_4776,N_4870);
or U5207 (N_5207,N_4759,N_4995);
nand U5208 (N_5208,N_4840,N_4763);
nor U5209 (N_5209,N_4779,N_4788);
nor U5210 (N_5210,N_4827,N_4955);
or U5211 (N_5211,N_4849,N_4869);
xnor U5212 (N_5212,N_4990,N_4831);
xor U5213 (N_5213,N_4893,N_4873);
xnor U5214 (N_5214,N_4971,N_4946);
nand U5215 (N_5215,N_4919,N_4915);
or U5216 (N_5216,N_4925,N_4842);
xor U5217 (N_5217,N_4954,N_4989);
and U5218 (N_5218,N_4939,N_4850);
nor U5219 (N_5219,N_4862,N_4909);
nor U5220 (N_5220,N_4887,N_4988);
xor U5221 (N_5221,N_4806,N_4846);
or U5222 (N_5222,N_4856,N_4927);
or U5223 (N_5223,N_4865,N_4903);
nor U5224 (N_5224,N_4752,N_4834);
and U5225 (N_5225,N_4766,N_4761);
and U5226 (N_5226,N_4792,N_4796);
nand U5227 (N_5227,N_4899,N_4812);
and U5228 (N_5228,N_4841,N_4979);
nand U5229 (N_5229,N_4776,N_4912);
nor U5230 (N_5230,N_4874,N_4830);
nor U5231 (N_5231,N_4777,N_4934);
nor U5232 (N_5232,N_4978,N_4960);
and U5233 (N_5233,N_4774,N_4968);
nand U5234 (N_5234,N_4907,N_4777);
or U5235 (N_5235,N_4777,N_4921);
xnor U5236 (N_5236,N_4986,N_4770);
and U5237 (N_5237,N_4926,N_4993);
nand U5238 (N_5238,N_4852,N_4804);
nand U5239 (N_5239,N_4848,N_4891);
nor U5240 (N_5240,N_4842,N_4787);
nor U5241 (N_5241,N_4814,N_4880);
and U5242 (N_5242,N_4751,N_4885);
or U5243 (N_5243,N_4983,N_4910);
xor U5244 (N_5244,N_4913,N_4793);
and U5245 (N_5245,N_4875,N_4902);
nand U5246 (N_5246,N_4888,N_4840);
xnor U5247 (N_5247,N_4795,N_4756);
xor U5248 (N_5248,N_4922,N_4756);
nor U5249 (N_5249,N_4763,N_4936);
or U5250 (N_5250,N_5049,N_5014);
nor U5251 (N_5251,N_5013,N_5079);
xor U5252 (N_5252,N_5153,N_5159);
or U5253 (N_5253,N_5133,N_5088);
nor U5254 (N_5254,N_5228,N_5199);
or U5255 (N_5255,N_5018,N_5230);
or U5256 (N_5256,N_5192,N_5032);
nor U5257 (N_5257,N_5148,N_5016);
nor U5258 (N_5258,N_5236,N_5074);
nand U5259 (N_5259,N_5132,N_5068);
or U5260 (N_5260,N_5034,N_5080);
xor U5261 (N_5261,N_5248,N_5063);
nor U5262 (N_5262,N_5136,N_5090);
nand U5263 (N_5263,N_5067,N_5029);
nand U5264 (N_5264,N_5023,N_5006);
nor U5265 (N_5265,N_5000,N_5007);
and U5266 (N_5266,N_5096,N_5163);
and U5267 (N_5267,N_5117,N_5108);
xnor U5268 (N_5268,N_5036,N_5167);
nand U5269 (N_5269,N_5008,N_5186);
nor U5270 (N_5270,N_5211,N_5065);
xnor U5271 (N_5271,N_5202,N_5051);
xnor U5272 (N_5272,N_5245,N_5205);
nand U5273 (N_5273,N_5046,N_5095);
and U5274 (N_5274,N_5247,N_5178);
nor U5275 (N_5275,N_5077,N_5235);
xnor U5276 (N_5276,N_5098,N_5191);
nor U5277 (N_5277,N_5081,N_5062);
nor U5278 (N_5278,N_5113,N_5213);
and U5279 (N_5279,N_5047,N_5224);
and U5280 (N_5280,N_5076,N_5086);
or U5281 (N_5281,N_5200,N_5085);
and U5282 (N_5282,N_5229,N_5028);
nor U5283 (N_5283,N_5212,N_5035);
xnor U5284 (N_5284,N_5075,N_5188);
nand U5285 (N_5285,N_5233,N_5050);
or U5286 (N_5286,N_5160,N_5243);
and U5287 (N_5287,N_5165,N_5135);
xor U5288 (N_5288,N_5138,N_5196);
xor U5289 (N_5289,N_5058,N_5037);
and U5290 (N_5290,N_5183,N_5091);
nand U5291 (N_5291,N_5151,N_5118);
xnor U5292 (N_5292,N_5209,N_5115);
nor U5293 (N_5293,N_5154,N_5126);
and U5294 (N_5294,N_5082,N_5112);
and U5295 (N_5295,N_5119,N_5227);
nor U5296 (N_5296,N_5124,N_5206);
nor U5297 (N_5297,N_5048,N_5149);
nand U5298 (N_5298,N_5187,N_5194);
or U5299 (N_5299,N_5231,N_5130);
or U5300 (N_5300,N_5240,N_5141);
nor U5301 (N_5301,N_5182,N_5177);
and U5302 (N_5302,N_5109,N_5170);
xnor U5303 (N_5303,N_5131,N_5114);
and U5304 (N_5304,N_5122,N_5015);
or U5305 (N_5305,N_5166,N_5104);
or U5306 (N_5306,N_5190,N_5221);
xor U5307 (N_5307,N_5070,N_5005);
or U5308 (N_5308,N_5217,N_5110);
xor U5309 (N_5309,N_5164,N_5021);
nor U5310 (N_5310,N_5173,N_5222);
xor U5311 (N_5311,N_5057,N_5030);
nor U5312 (N_5312,N_5127,N_5041);
xnor U5313 (N_5313,N_5094,N_5137);
and U5314 (N_5314,N_5161,N_5175);
and U5315 (N_5315,N_5121,N_5054);
xnor U5316 (N_5316,N_5234,N_5142);
or U5317 (N_5317,N_5061,N_5020);
nand U5318 (N_5318,N_5176,N_5225);
and U5319 (N_5319,N_5146,N_5214);
and U5320 (N_5320,N_5218,N_5026);
xnor U5321 (N_5321,N_5140,N_5155);
or U5322 (N_5322,N_5125,N_5134);
xnor U5323 (N_5323,N_5105,N_5107);
nor U5324 (N_5324,N_5093,N_5128);
or U5325 (N_5325,N_5197,N_5027);
nor U5326 (N_5326,N_5017,N_5189);
xnor U5327 (N_5327,N_5003,N_5180);
nor U5328 (N_5328,N_5203,N_5147);
nand U5329 (N_5329,N_5195,N_5038);
nand U5330 (N_5330,N_5071,N_5204);
nand U5331 (N_5331,N_5210,N_5056);
nor U5332 (N_5332,N_5123,N_5042);
nor U5333 (N_5333,N_5162,N_5089);
xor U5334 (N_5334,N_5156,N_5208);
nor U5335 (N_5335,N_5242,N_5179);
and U5336 (N_5336,N_5066,N_5073);
xnor U5337 (N_5337,N_5100,N_5011);
or U5338 (N_5338,N_5040,N_5168);
nand U5339 (N_5339,N_5169,N_5207);
nand U5340 (N_5340,N_5078,N_5241);
xnor U5341 (N_5341,N_5060,N_5039);
nor U5342 (N_5342,N_5201,N_5216);
and U5343 (N_5343,N_5244,N_5193);
and U5344 (N_5344,N_5106,N_5174);
nand U5345 (N_5345,N_5084,N_5022);
nand U5346 (N_5346,N_5150,N_5097);
nor U5347 (N_5347,N_5055,N_5145);
nor U5348 (N_5348,N_5045,N_5215);
nor U5349 (N_5349,N_5157,N_5219);
nand U5350 (N_5350,N_5246,N_5239);
or U5351 (N_5351,N_5198,N_5072);
and U5352 (N_5352,N_5010,N_5158);
nor U5353 (N_5353,N_5143,N_5238);
nand U5354 (N_5354,N_5009,N_5181);
xnor U5355 (N_5355,N_5099,N_5043);
or U5356 (N_5356,N_5024,N_5083);
xnor U5357 (N_5357,N_5012,N_5087);
or U5358 (N_5358,N_5139,N_5249);
nand U5359 (N_5359,N_5092,N_5059);
nor U5360 (N_5360,N_5111,N_5031);
and U5361 (N_5361,N_5025,N_5052);
xor U5362 (N_5362,N_5232,N_5103);
nor U5363 (N_5363,N_5069,N_5223);
nor U5364 (N_5364,N_5144,N_5171);
and U5365 (N_5365,N_5120,N_5001);
xnor U5366 (N_5366,N_5064,N_5237);
nand U5367 (N_5367,N_5116,N_5152);
xor U5368 (N_5368,N_5004,N_5101);
nor U5369 (N_5369,N_5129,N_5102);
or U5370 (N_5370,N_5220,N_5044);
xor U5371 (N_5371,N_5019,N_5185);
nor U5372 (N_5372,N_5172,N_5226);
or U5373 (N_5373,N_5053,N_5002);
and U5374 (N_5374,N_5184,N_5033);
and U5375 (N_5375,N_5145,N_5085);
and U5376 (N_5376,N_5099,N_5067);
xor U5377 (N_5377,N_5052,N_5236);
or U5378 (N_5378,N_5212,N_5067);
and U5379 (N_5379,N_5217,N_5198);
nand U5380 (N_5380,N_5166,N_5113);
nand U5381 (N_5381,N_5209,N_5192);
xor U5382 (N_5382,N_5013,N_5135);
nand U5383 (N_5383,N_5048,N_5195);
nor U5384 (N_5384,N_5244,N_5180);
nor U5385 (N_5385,N_5106,N_5230);
and U5386 (N_5386,N_5174,N_5082);
nor U5387 (N_5387,N_5133,N_5101);
and U5388 (N_5388,N_5149,N_5210);
nand U5389 (N_5389,N_5014,N_5130);
nand U5390 (N_5390,N_5197,N_5046);
and U5391 (N_5391,N_5179,N_5171);
or U5392 (N_5392,N_5041,N_5164);
nand U5393 (N_5393,N_5022,N_5121);
xnor U5394 (N_5394,N_5010,N_5247);
xnor U5395 (N_5395,N_5012,N_5223);
and U5396 (N_5396,N_5192,N_5170);
nor U5397 (N_5397,N_5123,N_5065);
or U5398 (N_5398,N_5181,N_5087);
or U5399 (N_5399,N_5165,N_5013);
nand U5400 (N_5400,N_5102,N_5091);
or U5401 (N_5401,N_5218,N_5172);
xnor U5402 (N_5402,N_5073,N_5247);
and U5403 (N_5403,N_5140,N_5184);
xnor U5404 (N_5404,N_5095,N_5015);
or U5405 (N_5405,N_5133,N_5066);
xnor U5406 (N_5406,N_5153,N_5213);
nand U5407 (N_5407,N_5092,N_5161);
xnor U5408 (N_5408,N_5071,N_5180);
xor U5409 (N_5409,N_5030,N_5022);
xor U5410 (N_5410,N_5176,N_5171);
and U5411 (N_5411,N_5131,N_5036);
nand U5412 (N_5412,N_5014,N_5167);
nor U5413 (N_5413,N_5230,N_5150);
nor U5414 (N_5414,N_5200,N_5204);
nand U5415 (N_5415,N_5140,N_5005);
xnor U5416 (N_5416,N_5022,N_5059);
xnor U5417 (N_5417,N_5164,N_5183);
nand U5418 (N_5418,N_5134,N_5158);
or U5419 (N_5419,N_5066,N_5164);
nor U5420 (N_5420,N_5236,N_5230);
and U5421 (N_5421,N_5071,N_5006);
xnor U5422 (N_5422,N_5095,N_5080);
nor U5423 (N_5423,N_5196,N_5060);
xor U5424 (N_5424,N_5086,N_5112);
xnor U5425 (N_5425,N_5153,N_5002);
and U5426 (N_5426,N_5016,N_5180);
xor U5427 (N_5427,N_5129,N_5075);
or U5428 (N_5428,N_5059,N_5237);
xnor U5429 (N_5429,N_5235,N_5240);
nor U5430 (N_5430,N_5052,N_5226);
or U5431 (N_5431,N_5103,N_5125);
nand U5432 (N_5432,N_5224,N_5206);
or U5433 (N_5433,N_5233,N_5216);
nor U5434 (N_5434,N_5241,N_5015);
or U5435 (N_5435,N_5169,N_5135);
and U5436 (N_5436,N_5053,N_5113);
nor U5437 (N_5437,N_5148,N_5060);
nor U5438 (N_5438,N_5121,N_5085);
or U5439 (N_5439,N_5032,N_5098);
nor U5440 (N_5440,N_5087,N_5213);
nand U5441 (N_5441,N_5139,N_5059);
nor U5442 (N_5442,N_5194,N_5023);
xor U5443 (N_5443,N_5234,N_5148);
nor U5444 (N_5444,N_5041,N_5046);
nand U5445 (N_5445,N_5150,N_5158);
and U5446 (N_5446,N_5011,N_5063);
nor U5447 (N_5447,N_5031,N_5189);
nor U5448 (N_5448,N_5056,N_5076);
xnor U5449 (N_5449,N_5163,N_5028);
nor U5450 (N_5450,N_5241,N_5179);
or U5451 (N_5451,N_5061,N_5234);
nand U5452 (N_5452,N_5114,N_5069);
or U5453 (N_5453,N_5119,N_5190);
nor U5454 (N_5454,N_5032,N_5089);
and U5455 (N_5455,N_5128,N_5209);
and U5456 (N_5456,N_5052,N_5058);
nor U5457 (N_5457,N_5244,N_5034);
xnor U5458 (N_5458,N_5011,N_5013);
nand U5459 (N_5459,N_5162,N_5034);
and U5460 (N_5460,N_5206,N_5157);
nand U5461 (N_5461,N_5022,N_5027);
nand U5462 (N_5462,N_5078,N_5081);
xnor U5463 (N_5463,N_5227,N_5072);
and U5464 (N_5464,N_5026,N_5094);
nor U5465 (N_5465,N_5106,N_5049);
xor U5466 (N_5466,N_5043,N_5131);
nand U5467 (N_5467,N_5229,N_5149);
and U5468 (N_5468,N_5241,N_5019);
or U5469 (N_5469,N_5114,N_5119);
nand U5470 (N_5470,N_5195,N_5190);
nor U5471 (N_5471,N_5152,N_5058);
nand U5472 (N_5472,N_5017,N_5211);
nor U5473 (N_5473,N_5194,N_5135);
nand U5474 (N_5474,N_5032,N_5127);
nor U5475 (N_5475,N_5221,N_5205);
nand U5476 (N_5476,N_5228,N_5040);
nor U5477 (N_5477,N_5242,N_5002);
nor U5478 (N_5478,N_5178,N_5155);
nand U5479 (N_5479,N_5228,N_5039);
nor U5480 (N_5480,N_5170,N_5232);
xnor U5481 (N_5481,N_5056,N_5112);
nand U5482 (N_5482,N_5224,N_5173);
and U5483 (N_5483,N_5141,N_5091);
xor U5484 (N_5484,N_5055,N_5038);
xnor U5485 (N_5485,N_5057,N_5224);
nor U5486 (N_5486,N_5229,N_5241);
nor U5487 (N_5487,N_5168,N_5165);
nand U5488 (N_5488,N_5175,N_5217);
nand U5489 (N_5489,N_5065,N_5102);
or U5490 (N_5490,N_5028,N_5013);
and U5491 (N_5491,N_5055,N_5054);
nand U5492 (N_5492,N_5140,N_5105);
nor U5493 (N_5493,N_5061,N_5128);
or U5494 (N_5494,N_5130,N_5071);
nor U5495 (N_5495,N_5080,N_5248);
xor U5496 (N_5496,N_5226,N_5108);
nor U5497 (N_5497,N_5115,N_5116);
nand U5498 (N_5498,N_5104,N_5171);
or U5499 (N_5499,N_5022,N_5206);
and U5500 (N_5500,N_5497,N_5479);
and U5501 (N_5501,N_5441,N_5344);
nand U5502 (N_5502,N_5380,N_5256);
and U5503 (N_5503,N_5404,N_5393);
and U5504 (N_5504,N_5449,N_5397);
and U5505 (N_5505,N_5467,N_5407);
or U5506 (N_5506,N_5294,N_5286);
or U5507 (N_5507,N_5364,N_5465);
xor U5508 (N_5508,N_5260,N_5428);
nor U5509 (N_5509,N_5492,N_5399);
or U5510 (N_5510,N_5496,N_5346);
nor U5511 (N_5511,N_5369,N_5480);
and U5512 (N_5512,N_5445,N_5386);
xnor U5513 (N_5513,N_5471,N_5403);
or U5514 (N_5514,N_5491,N_5468);
nand U5515 (N_5515,N_5297,N_5341);
nor U5516 (N_5516,N_5388,N_5405);
nor U5517 (N_5517,N_5318,N_5427);
nor U5518 (N_5518,N_5422,N_5265);
and U5519 (N_5519,N_5466,N_5335);
xor U5520 (N_5520,N_5308,N_5410);
nand U5521 (N_5521,N_5322,N_5412);
nand U5522 (N_5522,N_5377,N_5320);
or U5523 (N_5523,N_5330,N_5283);
nand U5524 (N_5524,N_5462,N_5278);
or U5525 (N_5525,N_5316,N_5400);
or U5526 (N_5526,N_5332,N_5423);
and U5527 (N_5527,N_5257,N_5359);
nor U5528 (N_5528,N_5334,N_5448);
and U5529 (N_5529,N_5474,N_5317);
xnor U5530 (N_5530,N_5355,N_5319);
and U5531 (N_5531,N_5337,N_5374);
or U5532 (N_5532,N_5424,N_5284);
xor U5533 (N_5533,N_5362,N_5457);
nor U5534 (N_5534,N_5280,N_5490);
nor U5535 (N_5535,N_5326,N_5383);
xor U5536 (N_5536,N_5347,N_5487);
and U5537 (N_5537,N_5387,N_5343);
or U5538 (N_5538,N_5455,N_5444);
nor U5539 (N_5539,N_5498,N_5494);
nor U5540 (N_5540,N_5477,N_5372);
xnor U5541 (N_5541,N_5357,N_5287);
xor U5542 (N_5542,N_5483,N_5253);
nand U5543 (N_5543,N_5370,N_5327);
xnor U5544 (N_5544,N_5430,N_5349);
and U5545 (N_5545,N_5434,N_5406);
nor U5546 (N_5546,N_5361,N_5481);
nor U5547 (N_5547,N_5440,N_5459);
nand U5548 (N_5548,N_5255,N_5447);
nor U5549 (N_5549,N_5266,N_5458);
and U5550 (N_5550,N_5351,N_5415);
nand U5551 (N_5551,N_5360,N_5476);
and U5552 (N_5552,N_5421,N_5478);
xnor U5553 (N_5553,N_5276,N_5254);
xnor U5554 (N_5554,N_5385,N_5358);
xnor U5555 (N_5555,N_5352,N_5270);
or U5556 (N_5556,N_5398,N_5268);
nand U5557 (N_5557,N_5273,N_5464);
and U5558 (N_5558,N_5435,N_5301);
and U5559 (N_5559,N_5391,N_5281);
xor U5560 (N_5560,N_5438,N_5356);
or U5561 (N_5561,N_5271,N_5413);
or U5562 (N_5562,N_5470,N_5321);
or U5563 (N_5563,N_5315,N_5417);
or U5564 (N_5564,N_5371,N_5473);
and U5565 (N_5565,N_5396,N_5432);
nand U5566 (N_5566,N_5354,N_5456);
and U5567 (N_5567,N_5279,N_5488);
nand U5568 (N_5568,N_5461,N_5310);
and U5569 (N_5569,N_5258,N_5433);
xor U5570 (N_5570,N_5418,N_5302);
xor U5571 (N_5571,N_5451,N_5314);
and U5572 (N_5572,N_5442,N_5416);
nor U5573 (N_5573,N_5298,N_5311);
xor U5574 (N_5574,N_5420,N_5296);
nor U5575 (N_5575,N_5267,N_5402);
or U5576 (N_5576,N_5325,N_5378);
or U5577 (N_5577,N_5363,N_5251);
nand U5578 (N_5578,N_5304,N_5290);
or U5579 (N_5579,N_5408,N_5323);
or U5580 (N_5580,N_5307,N_5475);
nor U5581 (N_5581,N_5437,N_5300);
and U5582 (N_5582,N_5382,N_5431);
or U5583 (N_5583,N_5379,N_5259);
nor U5584 (N_5584,N_5485,N_5489);
or U5585 (N_5585,N_5472,N_5252);
xnor U5586 (N_5586,N_5285,N_5450);
xnor U5587 (N_5587,N_5384,N_5342);
nor U5588 (N_5588,N_5375,N_5365);
xor U5589 (N_5589,N_5469,N_5373);
nand U5590 (N_5590,N_5401,N_5493);
nor U5591 (N_5591,N_5460,N_5295);
nor U5592 (N_5592,N_5324,N_5312);
nor U5593 (N_5593,N_5272,N_5436);
nand U5594 (N_5594,N_5275,N_5446);
nand U5595 (N_5595,N_5305,N_5348);
or U5596 (N_5596,N_5338,N_5495);
nand U5597 (N_5597,N_5443,N_5282);
nand U5598 (N_5598,N_5261,N_5339);
and U5599 (N_5599,N_5381,N_5453);
nand U5600 (N_5600,N_5414,N_5429);
nor U5601 (N_5601,N_5264,N_5292);
nor U5602 (N_5602,N_5313,N_5367);
or U5603 (N_5603,N_5329,N_5353);
and U5604 (N_5604,N_5395,N_5288);
or U5605 (N_5605,N_5499,N_5389);
nand U5606 (N_5606,N_5486,N_5439);
xor U5607 (N_5607,N_5303,N_5331);
xor U5608 (N_5608,N_5293,N_5250);
xnor U5609 (N_5609,N_5336,N_5291);
nand U5610 (N_5610,N_5309,N_5333);
nor U5611 (N_5611,N_5376,N_5299);
and U5612 (N_5612,N_5392,N_5289);
or U5613 (N_5613,N_5394,N_5366);
and U5614 (N_5614,N_5484,N_5368);
or U5615 (N_5615,N_5328,N_5426);
and U5616 (N_5616,N_5274,N_5454);
nand U5617 (N_5617,N_5345,N_5350);
and U5618 (N_5618,N_5409,N_5340);
or U5619 (N_5619,N_5482,N_5390);
xnor U5620 (N_5620,N_5425,N_5306);
and U5621 (N_5621,N_5411,N_5263);
nor U5622 (N_5622,N_5262,N_5277);
xor U5623 (N_5623,N_5452,N_5269);
nor U5624 (N_5624,N_5419,N_5463);
and U5625 (N_5625,N_5316,N_5355);
and U5626 (N_5626,N_5266,N_5479);
nand U5627 (N_5627,N_5351,N_5371);
and U5628 (N_5628,N_5465,N_5358);
or U5629 (N_5629,N_5435,N_5267);
or U5630 (N_5630,N_5252,N_5313);
xnor U5631 (N_5631,N_5436,N_5494);
nand U5632 (N_5632,N_5356,N_5398);
and U5633 (N_5633,N_5418,N_5428);
nor U5634 (N_5634,N_5278,N_5481);
nor U5635 (N_5635,N_5411,N_5291);
or U5636 (N_5636,N_5460,N_5357);
and U5637 (N_5637,N_5337,N_5425);
or U5638 (N_5638,N_5347,N_5273);
xor U5639 (N_5639,N_5293,N_5354);
and U5640 (N_5640,N_5253,N_5447);
xor U5641 (N_5641,N_5487,N_5399);
xnor U5642 (N_5642,N_5494,N_5275);
and U5643 (N_5643,N_5365,N_5483);
nand U5644 (N_5644,N_5268,N_5300);
and U5645 (N_5645,N_5321,N_5308);
xor U5646 (N_5646,N_5254,N_5350);
or U5647 (N_5647,N_5415,N_5381);
and U5648 (N_5648,N_5256,N_5374);
nand U5649 (N_5649,N_5356,N_5335);
xnor U5650 (N_5650,N_5349,N_5451);
nand U5651 (N_5651,N_5400,N_5469);
nor U5652 (N_5652,N_5307,N_5489);
nand U5653 (N_5653,N_5288,N_5463);
or U5654 (N_5654,N_5390,N_5265);
nor U5655 (N_5655,N_5493,N_5488);
and U5656 (N_5656,N_5395,N_5397);
and U5657 (N_5657,N_5493,N_5419);
or U5658 (N_5658,N_5374,N_5349);
xnor U5659 (N_5659,N_5307,N_5254);
or U5660 (N_5660,N_5495,N_5324);
nor U5661 (N_5661,N_5352,N_5413);
nor U5662 (N_5662,N_5324,N_5458);
and U5663 (N_5663,N_5322,N_5310);
nor U5664 (N_5664,N_5460,N_5371);
nand U5665 (N_5665,N_5274,N_5331);
xor U5666 (N_5666,N_5344,N_5253);
and U5667 (N_5667,N_5393,N_5389);
nand U5668 (N_5668,N_5295,N_5326);
nor U5669 (N_5669,N_5345,N_5436);
xnor U5670 (N_5670,N_5408,N_5479);
nor U5671 (N_5671,N_5296,N_5472);
nor U5672 (N_5672,N_5497,N_5458);
and U5673 (N_5673,N_5330,N_5369);
nand U5674 (N_5674,N_5325,N_5405);
and U5675 (N_5675,N_5467,N_5428);
and U5676 (N_5676,N_5493,N_5478);
and U5677 (N_5677,N_5403,N_5353);
xor U5678 (N_5678,N_5379,N_5331);
nor U5679 (N_5679,N_5494,N_5332);
xor U5680 (N_5680,N_5406,N_5256);
nor U5681 (N_5681,N_5470,N_5484);
nand U5682 (N_5682,N_5350,N_5382);
nand U5683 (N_5683,N_5438,N_5467);
or U5684 (N_5684,N_5304,N_5375);
xnor U5685 (N_5685,N_5340,N_5424);
xor U5686 (N_5686,N_5341,N_5426);
or U5687 (N_5687,N_5368,N_5306);
nand U5688 (N_5688,N_5447,N_5431);
nand U5689 (N_5689,N_5289,N_5391);
nand U5690 (N_5690,N_5319,N_5290);
and U5691 (N_5691,N_5392,N_5261);
or U5692 (N_5692,N_5272,N_5302);
xor U5693 (N_5693,N_5399,N_5421);
xnor U5694 (N_5694,N_5316,N_5498);
xnor U5695 (N_5695,N_5464,N_5482);
nor U5696 (N_5696,N_5338,N_5481);
nor U5697 (N_5697,N_5282,N_5484);
nand U5698 (N_5698,N_5495,N_5427);
nor U5699 (N_5699,N_5393,N_5401);
nand U5700 (N_5700,N_5443,N_5451);
xor U5701 (N_5701,N_5413,N_5387);
nand U5702 (N_5702,N_5497,N_5430);
nand U5703 (N_5703,N_5458,N_5396);
nor U5704 (N_5704,N_5461,N_5371);
or U5705 (N_5705,N_5405,N_5418);
xor U5706 (N_5706,N_5319,N_5447);
or U5707 (N_5707,N_5346,N_5319);
xnor U5708 (N_5708,N_5420,N_5387);
nand U5709 (N_5709,N_5325,N_5334);
and U5710 (N_5710,N_5397,N_5311);
or U5711 (N_5711,N_5491,N_5461);
nand U5712 (N_5712,N_5436,N_5489);
and U5713 (N_5713,N_5385,N_5340);
xor U5714 (N_5714,N_5346,N_5384);
nor U5715 (N_5715,N_5459,N_5252);
nor U5716 (N_5716,N_5359,N_5479);
xnor U5717 (N_5717,N_5257,N_5488);
nand U5718 (N_5718,N_5330,N_5473);
and U5719 (N_5719,N_5289,N_5362);
and U5720 (N_5720,N_5499,N_5344);
and U5721 (N_5721,N_5260,N_5348);
and U5722 (N_5722,N_5498,N_5292);
or U5723 (N_5723,N_5405,N_5463);
nor U5724 (N_5724,N_5309,N_5395);
nor U5725 (N_5725,N_5341,N_5347);
nand U5726 (N_5726,N_5378,N_5348);
or U5727 (N_5727,N_5410,N_5317);
or U5728 (N_5728,N_5472,N_5448);
nor U5729 (N_5729,N_5298,N_5476);
or U5730 (N_5730,N_5446,N_5344);
nor U5731 (N_5731,N_5473,N_5414);
and U5732 (N_5732,N_5279,N_5309);
or U5733 (N_5733,N_5436,N_5432);
and U5734 (N_5734,N_5454,N_5350);
nand U5735 (N_5735,N_5267,N_5343);
nor U5736 (N_5736,N_5253,N_5469);
or U5737 (N_5737,N_5409,N_5382);
xor U5738 (N_5738,N_5371,N_5409);
or U5739 (N_5739,N_5370,N_5401);
or U5740 (N_5740,N_5320,N_5280);
xnor U5741 (N_5741,N_5398,N_5407);
and U5742 (N_5742,N_5259,N_5413);
and U5743 (N_5743,N_5315,N_5300);
and U5744 (N_5744,N_5341,N_5476);
nor U5745 (N_5745,N_5379,N_5455);
nand U5746 (N_5746,N_5280,N_5257);
nor U5747 (N_5747,N_5285,N_5410);
nor U5748 (N_5748,N_5454,N_5306);
or U5749 (N_5749,N_5335,N_5359);
xor U5750 (N_5750,N_5636,N_5577);
or U5751 (N_5751,N_5743,N_5615);
nand U5752 (N_5752,N_5661,N_5508);
and U5753 (N_5753,N_5638,N_5557);
nand U5754 (N_5754,N_5620,N_5626);
and U5755 (N_5755,N_5655,N_5512);
and U5756 (N_5756,N_5528,N_5540);
or U5757 (N_5757,N_5598,N_5574);
nand U5758 (N_5758,N_5618,N_5728);
and U5759 (N_5759,N_5503,N_5710);
or U5760 (N_5760,N_5610,N_5741);
nor U5761 (N_5761,N_5525,N_5732);
or U5762 (N_5762,N_5699,N_5719);
and U5763 (N_5763,N_5734,N_5599);
or U5764 (N_5764,N_5602,N_5568);
or U5765 (N_5765,N_5742,N_5644);
and U5766 (N_5766,N_5652,N_5562);
and U5767 (N_5767,N_5647,N_5749);
xor U5768 (N_5768,N_5679,N_5666);
xnor U5769 (N_5769,N_5695,N_5544);
nand U5770 (N_5770,N_5531,N_5546);
and U5771 (N_5771,N_5648,N_5507);
nand U5772 (N_5772,N_5663,N_5646);
or U5773 (N_5773,N_5736,N_5642);
nor U5774 (N_5774,N_5502,N_5706);
nor U5775 (N_5775,N_5549,N_5583);
xor U5776 (N_5776,N_5587,N_5685);
nor U5777 (N_5777,N_5675,N_5662);
nor U5778 (N_5778,N_5571,N_5542);
or U5779 (N_5779,N_5596,N_5552);
nand U5780 (N_5780,N_5690,N_5623);
xor U5781 (N_5781,N_5541,N_5580);
nand U5782 (N_5782,N_5709,N_5594);
or U5783 (N_5783,N_5553,N_5591);
nand U5784 (N_5784,N_5523,N_5578);
and U5785 (N_5785,N_5527,N_5713);
nand U5786 (N_5786,N_5622,N_5585);
or U5787 (N_5787,N_5593,N_5506);
nor U5788 (N_5788,N_5723,N_5673);
or U5789 (N_5789,N_5515,N_5521);
xnor U5790 (N_5790,N_5530,N_5608);
or U5791 (N_5791,N_5659,N_5563);
and U5792 (N_5792,N_5631,N_5700);
nor U5793 (N_5793,N_5603,N_5566);
nor U5794 (N_5794,N_5516,N_5722);
xnor U5795 (N_5795,N_5555,N_5746);
xnor U5796 (N_5796,N_5724,N_5606);
or U5797 (N_5797,N_5688,N_5703);
and U5798 (N_5798,N_5522,N_5535);
and U5799 (N_5799,N_5588,N_5616);
nor U5800 (N_5800,N_5671,N_5680);
and U5801 (N_5801,N_5669,N_5733);
and U5802 (N_5802,N_5660,N_5501);
and U5803 (N_5803,N_5628,N_5513);
nand U5804 (N_5804,N_5702,N_5641);
and U5805 (N_5805,N_5554,N_5509);
and U5806 (N_5806,N_5511,N_5707);
nand U5807 (N_5807,N_5721,N_5518);
or U5808 (N_5808,N_5635,N_5570);
nor U5809 (N_5809,N_5584,N_5668);
nand U5810 (N_5810,N_5738,N_5576);
nand U5811 (N_5811,N_5670,N_5543);
and U5812 (N_5812,N_5633,N_5505);
or U5813 (N_5813,N_5708,N_5545);
or U5814 (N_5814,N_5621,N_5657);
nor U5815 (N_5815,N_5717,N_5637);
nand U5816 (N_5816,N_5529,N_5579);
xor U5817 (N_5817,N_5605,N_5575);
nor U5818 (N_5818,N_5533,N_5601);
and U5819 (N_5819,N_5589,N_5643);
xnor U5820 (N_5820,N_5534,N_5716);
nor U5821 (N_5821,N_5650,N_5731);
nand U5822 (N_5822,N_5682,N_5510);
nand U5823 (N_5823,N_5627,N_5677);
xnor U5824 (N_5824,N_5745,N_5725);
nand U5825 (N_5825,N_5697,N_5747);
nand U5826 (N_5826,N_5692,N_5514);
nor U5827 (N_5827,N_5726,N_5592);
and U5828 (N_5828,N_5611,N_5613);
or U5829 (N_5829,N_5667,N_5590);
or U5830 (N_5830,N_5678,N_5569);
nand U5831 (N_5831,N_5524,N_5609);
xnor U5832 (N_5832,N_5520,N_5681);
xnor U5833 (N_5833,N_5547,N_5730);
and U5834 (N_5834,N_5532,N_5674);
or U5835 (N_5835,N_5718,N_5536);
and U5836 (N_5836,N_5691,N_5630);
or U5837 (N_5837,N_5735,N_5581);
xnor U5838 (N_5838,N_5639,N_5720);
xor U5839 (N_5839,N_5651,N_5559);
nor U5840 (N_5840,N_5629,N_5619);
and U5841 (N_5841,N_5664,N_5558);
nor U5842 (N_5842,N_5634,N_5686);
xor U5843 (N_5843,N_5556,N_5704);
nand U5844 (N_5844,N_5715,N_5687);
nand U5845 (N_5845,N_5538,N_5645);
and U5846 (N_5846,N_5564,N_5739);
nand U5847 (N_5847,N_5672,N_5711);
or U5848 (N_5848,N_5658,N_5632);
and U5849 (N_5849,N_5698,N_5653);
nor U5850 (N_5850,N_5539,N_5519);
and U5851 (N_5851,N_5640,N_5595);
xnor U5852 (N_5852,N_5649,N_5740);
nand U5853 (N_5853,N_5600,N_5624);
nor U5854 (N_5854,N_5727,N_5607);
xnor U5855 (N_5855,N_5573,N_5665);
nor U5856 (N_5856,N_5684,N_5729);
or U5857 (N_5857,N_5550,N_5712);
xnor U5858 (N_5858,N_5537,N_5500);
xor U5859 (N_5859,N_5654,N_5551);
nor U5860 (N_5860,N_5748,N_5548);
nor U5861 (N_5861,N_5696,N_5744);
or U5862 (N_5862,N_5617,N_5597);
or U5863 (N_5863,N_5625,N_5656);
xnor U5864 (N_5864,N_5614,N_5572);
nand U5865 (N_5865,N_5517,N_5586);
and U5866 (N_5866,N_5689,N_5561);
nand U5867 (N_5867,N_5526,N_5693);
xor U5868 (N_5868,N_5737,N_5604);
and U5869 (N_5869,N_5504,N_5567);
or U5870 (N_5870,N_5714,N_5676);
and U5871 (N_5871,N_5683,N_5582);
xnor U5872 (N_5872,N_5612,N_5565);
nand U5873 (N_5873,N_5705,N_5701);
nor U5874 (N_5874,N_5560,N_5694);
nand U5875 (N_5875,N_5503,N_5545);
nand U5876 (N_5876,N_5604,N_5552);
xnor U5877 (N_5877,N_5570,N_5745);
and U5878 (N_5878,N_5663,N_5681);
nor U5879 (N_5879,N_5504,N_5695);
nor U5880 (N_5880,N_5565,N_5639);
nand U5881 (N_5881,N_5666,N_5654);
and U5882 (N_5882,N_5567,N_5706);
nor U5883 (N_5883,N_5604,N_5712);
xor U5884 (N_5884,N_5570,N_5577);
nor U5885 (N_5885,N_5675,N_5529);
xnor U5886 (N_5886,N_5604,N_5533);
or U5887 (N_5887,N_5629,N_5613);
nand U5888 (N_5888,N_5624,N_5704);
nand U5889 (N_5889,N_5634,N_5553);
nand U5890 (N_5890,N_5540,N_5579);
xnor U5891 (N_5891,N_5740,N_5633);
or U5892 (N_5892,N_5590,N_5506);
xnor U5893 (N_5893,N_5508,N_5605);
nand U5894 (N_5894,N_5703,N_5521);
and U5895 (N_5895,N_5569,N_5602);
xor U5896 (N_5896,N_5513,N_5519);
nor U5897 (N_5897,N_5609,N_5578);
nor U5898 (N_5898,N_5632,N_5602);
nor U5899 (N_5899,N_5527,N_5663);
nand U5900 (N_5900,N_5559,N_5562);
xnor U5901 (N_5901,N_5579,N_5628);
xor U5902 (N_5902,N_5534,N_5521);
and U5903 (N_5903,N_5655,N_5722);
and U5904 (N_5904,N_5727,N_5658);
xor U5905 (N_5905,N_5682,N_5512);
or U5906 (N_5906,N_5721,N_5717);
and U5907 (N_5907,N_5713,N_5744);
xnor U5908 (N_5908,N_5539,N_5588);
nand U5909 (N_5909,N_5629,N_5705);
and U5910 (N_5910,N_5710,N_5713);
and U5911 (N_5911,N_5541,N_5690);
nor U5912 (N_5912,N_5526,N_5586);
nor U5913 (N_5913,N_5662,N_5543);
nand U5914 (N_5914,N_5545,N_5532);
xnor U5915 (N_5915,N_5623,N_5660);
and U5916 (N_5916,N_5748,N_5640);
nor U5917 (N_5917,N_5704,N_5670);
xnor U5918 (N_5918,N_5520,N_5560);
nor U5919 (N_5919,N_5542,N_5651);
or U5920 (N_5920,N_5717,N_5515);
nand U5921 (N_5921,N_5698,N_5586);
and U5922 (N_5922,N_5604,N_5654);
xor U5923 (N_5923,N_5579,N_5523);
nand U5924 (N_5924,N_5545,N_5623);
and U5925 (N_5925,N_5505,N_5535);
or U5926 (N_5926,N_5573,N_5566);
xnor U5927 (N_5927,N_5641,N_5740);
and U5928 (N_5928,N_5644,N_5640);
xnor U5929 (N_5929,N_5677,N_5618);
nor U5930 (N_5930,N_5678,N_5630);
and U5931 (N_5931,N_5653,N_5691);
nor U5932 (N_5932,N_5626,N_5635);
nand U5933 (N_5933,N_5509,N_5689);
xor U5934 (N_5934,N_5600,N_5721);
or U5935 (N_5935,N_5579,N_5653);
nand U5936 (N_5936,N_5668,N_5616);
nand U5937 (N_5937,N_5591,N_5728);
and U5938 (N_5938,N_5661,N_5681);
and U5939 (N_5939,N_5682,N_5611);
nor U5940 (N_5940,N_5539,N_5569);
nand U5941 (N_5941,N_5533,N_5506);
xnor U5942 (N_5942,N_5641,N_5650);
nor U5943 (N_5943,N_5690,N_5589);
xnor U5944 (N_5944,N_5673,N_5590);
or U5945 (N_5945,N_5680,N_5577);
and U5946 (N_5946,N_5651,N_5630);
or U5947 (N_5947,N_5745,N_5621);
or U5948 (N_5948,N_5567,N_5623);
or U5949 (N_5949,N_5628,N_5562);
nand U5950 (N_5950,N_5523,N_5721);
nor U5951 (N_5951,N_5608,N_5697);
or U5952 (N_5952,N_5746,N_5717);
xor U5953 (N_5953,N_5687,N_5548);
nand U5954 (N_5954,N_5657,N_5640);
xnor U5955 (N_5955,N_5630,N_5524);
and U5956 (N_5956,N_5697,N_5694);
nand U5957 (N_5957,N_5534,N_5594);
nand U5958 (N_5958,N_5610,N_5614);
xnor U5959 (N_5959,N_5571,N_5562);
and U5960 (N_5960,N_5629,N_5722);
nor U5961 (N_5961,N_5610,N_5720);
and U5962 (N_5962,N_5502,N_5685);
nand U5963 (N_5963,N_5701,N_5598);
nand U5964 (N_5964,N_5647,N_5671);
or U5965 (N_5965,N_5643,N_5581);
or U5966 (N_5966,N_5666,N_5545);
xnor U5967 (N_5967,N_5699,N_5648);
or U5968 (N_5968,N_5682,N_5684);
xnor U5969 (N_5969,N_5630,N_5667);
nand U5970 (N_5970,N_5507,N_5543);
nor U5971 (N_5971,N_5694,N_5527);
xor U5972 (N_5972,N_5520,N_5571);
nor U5973 (N_5973,N_5713,N_5562);
nor U5974 (N_5974,N_5638,N_5705);
nand U5975 (N_5975,N_5577,N_5530);
nand U5976 (N_5976,N_5648,N_5566);
or U5977 (N_5977,N_5628,N_5665);
and U5978 (N_5978,N_5608,N_5694);
xor U5979 (N_5979,N_5542,N_5621);
nand U5980 (N_5980,N_5541,N_5589);
nand U5981 (N_5981,N_5738,N_5728);
or U5982 (N_5982,N_5691,N_5571);
and U5983 (N_5983,N_5677,N_5586);
xnor U5984 (N_5984,N_5714,N_5679);
or U5985 (N_5985,N_5705,N_5674);
xnor U5986 (N_5986,N_5673,N_5687);
and U5987 (N_5987,N_5571,N_5606);
and U5988 (N_5988,N_5640,N_5558);
or U5989 (N_5989,N_5595,N_5683);
nor U5990 (N_5990,N_5686,N_5687);
xor U5991 (N_5991,N_5749,N_5577);
or U5992 (N_5992,N_5568,N_5735);
or U5993 (N_5993,N_5566,N_5662);
or U5994 (N_5994,N_5521,N_5721);
or U5995 (N_5995,N_5680,N_5618);
or U5996 (N_5996,N_5675,N_5544);
xor U5997 (N_5997,N_5716,N_5734);
and U5998 (N_5998,N_5742,N_5587);
and U5999 (N_5999,N_5729,N_5604);
nor U6000 (N_6000,N_5783,N_5791);
xor U6001 (N_6001,N_5974,N_5830);
nand U6002 (N_6002,N_5819,N_5834);
and U6003 (N_6003,N_5848,N_5851);
and U6004 (N_6004,N_5939,N_5870);
xor U6005 (N_6005,N_5949,N_5998);
nand U6006 (N_6006,N_5868,N_5981);
nand U6007 (N_6007,N_5904,N_5840);
or U6008 (N_6008,N_5975,N_5962);
nor U6009 (N_6009,N_5751,N_5978);
or U6010 (N_6010,N_5766,N_5780);
xnor U6011 (N_6011,N_5935,N_5817);
or U6012 (N_6012,N_5992,N_5768);
or U6013 (N_6013,N_5794,N_5806);
or U6014 (N_6014,N_5779,N_5786);
and U6015 (N_6015,N_5883,N_5973);
and U6016 (N_6016,N_5857,N_5898);
nor U6017 (N_6017,N_5863,N_5968);
or U6018 (N_6018,N_5896,N_5999);
xor U6019 (N_6019,N_5946,N_5832);
or U6020 (N_6020,N_5777,N_5812);
and U6021 (N_6021,N_5754,N_5858);
and U6022 (N_6022,N_5790,N_5867);
or U6023 (N_6023,N_5861,N_5967);
xnor U6024 (N_6024,N_5818,N_5866);
xnor U6025 (N_6025,N_5924,N_5796);
and U6026 (N_6026,N_5805,N_5882);
or U6027 (N_6027,N_5825,N_5960);
nor U6028 (N_6028,N_5893,N_5774);
xnor U6029 (N_6029,N_5944,N_5782);
xnor U6030 (N_6030,N_5918,N_5936);
or U6031 (N_6031,N_5801,N_5993);
xnor U6032 (N_6032,N_5839,N_5810);
nand U6033 (N_6033,N_5837,N_5943);
xnor U6034 (N_6034,N_5894,N_5966);
nand U6035 (N_6035,N_5907,N_5873);
or U6036 (N_6036,N_5910,N_5776);
or U6037 (N_6037,N_5959,N_5831);
xnor U6038 (N_6038,N_5821,N_5976);
or U6039 (N_6039,N_5938,N_5787);
xor U6040 (N_6040,N_5778,N_5835);
xnor U6041 (N_6041,N_5878,N_5877);
or U6042 (N_6042,N_5916,N_5864);
xor U6043 (N_6043,N_5802,N_5970);
and U6044 (N_6044,N_5969,N_5755);
nand U6045 (N_6045,N_5881,N_5875);
nand U6046 (N_6046,N_5847,N_5876);
and U6047 (N_6047,N_5797,N_5862);
and U6048 (N_6048,N_5979,N_5888);
xnor U6049 (N_6049,N_5921,N_5899);
nand U6050 (N_6050,N_5892,N_5809);
nand U6051 (N_6051,N_5757,N_5905);
nand U6052 (N_6052,N_5849,N_5769);
or U6053 (N_6053,N_5972,N_5799);
or U6054 (N_6054,N_5761,N_5824);
nand U6055 (N_6055,N_5953,N_5872);
or U6056 (N_6056,N_5995,N_5767);
or U6057 (N_6057,N_5895,N_5901);
nand U6058 (N_6058,N_5990,N_5937);
nor U6059 (N_6059,N_5865,N_5854);
nand U6060 (N_6060,N_5833,N_5971);
xnor U6061 (N_6061,N_5900,N_5951);
xor U6062 (N_6062,N_5983,N_5765);
nand U6063 (N_6063,N_5930,N_5991);
nand U6064 (N_6064,N_5793,N_5869);
or U6065 (N_6065,N_5752,N_5795);
or U6066 (N_6066,N_5948,N_5917);
nor U6067 (N_6067,N_5813,N_5792);
and U6068 (N_6068,N_5989,N_5909);
nand U6069 (N_6069,N_5803,N_5852);
nand U6070 (N_6070,N_5773,N_5919);
nand U6071 (N_6071,N_5758,N_5997);
nand U6072 (N_6072,N_5996,N_5952);
or U6073 (N_6073,N_5926,N_5928);
and U6074 (N_6074,N_5955,N_5932);
and U6075 (N_6075,N_5855,N_5986);
xnor U6076 (N_6076,N_5826,N_5950);
nand U6077 (N_6077,N_5889,N_5923);
nor U6078 (N_6078,N_5816,N_5902);
nor U6079 (N_6079,N_5850,N_5763);
and U6080 (N_6080,N_5856,N_5775);
and U6081 (N_6081,N_5804,N_5942);
nand U6082 (N_6082,N_5756,N_5984);
or U6083 (N_6083,N_5982,N_5933);
nand U6084 (N_6084,N_5785,N_5827);
and U6085 (N_6085,N_5925,N_5843);
and U6086 (N_6086,N_5891,N_5800);
or U6087 (N_6087,N_5890,N_5945);
nor U6088 (N_6088,N_5771,N_5841);
or U6089 (N_6089,N_5903,N_5922);
and U6090 (N_6090,N_5823,N_5963);
or U6091 (N_6091,N_5822,N_5940);
and U6092 (N_6092,N_5836,N_5987);
and U6093 (N_6093,N_5815,N_5859);
and U6094 (N_6094,N_5964,N_5954);
or U6095 (N_6095,N_5762,N_5871);
and U6096 (N_6096,N_5912,N_5759);
nand U6097 (N_6097,N_5808,N_5811);
or U6098 (N_6098,N_5807,N_5844);
or U6099 (N_6099,N_5798,N_5887);
or U6100 (N_6100,N_5886,N_5956);
and U6101 (N_6101,N_5920,N_5906);
nand U6102 (N_6102,N_5879,N_5764);
xnor U6103 (N_6103,N_5829,N_5958);
xor U6104 (N_6104,N_5770,N_5884);
xor U6105 (N_6105,N_5941,N_5860);
and U6106 (N_6106,N_5988,N_5820);
or U6107 (N_6107,N_5760,N_5980);
nor U6108 (N_6108,N_5927,N_5885);
xnor U6109 (N_6109,N_5915,N_5985);
and U6110 (N_6110,N_5846,N_5853);
nor U6111 (N_6111,N_5880,N_5957);
or U6112 (N_6112,N_5842,N_5838);
and U6113 (N_6113,N_5845,N_5772);
and U6114 (N_6114,N_5914,N_5961);
xor U6115 (N_6115,N_5750,N_5977);
nand U6116 (N_6116,N_5934,N_5994);
and U6117 (N_6117,N_5789,N_5947);
nor U6118 (N_6118,N_5828,N_5931);
and U6119 (N_6119,N_5788,N_5908);
and U6120 (N_6120,N_5911,N_5897);
and U6121 (N_6121,N_5913,N_5929);
nand U6122 (N_6122,N_5814,N_5781);
and U6123 (N_6123,N_5784,N_5965);
or U6124 (N_6124,N_5874,N_5753);
or U6125 (N_6125,N_5902,N_5940);
xor U6126 (N_6126,N_5753,N_5945);
or U6127 (N_6127,N_5845,N_5792);
and U6128 (N_6128,N_5874,N_5821);
nand U6129 (N_6129,N_5907,N_5793);
and U6130 (N_6130,N_5953,N_5836);
or U6131 (N_6131,N_5867,N_5791);
nand U6132 (N_6132,N_5885,N_5766);
nand U6133 (N_6133,N_5970,N_5879);
nor U6134 (N_6134,N_5923,N_5969);
xnor U6135 (N_6135,N_5986,N_5898);
or U6136 (N_6136,N_5984,N_5871);
and U6137 (N_6137,N_5780,N_5831);
xor U6138 (N_6138,N_5938,N_5890);
nor U6139 (N_6139,N_5836,N_5766);
nand U6140 (N_6140,N_5913,N_5904);
nand U6141 (N_6141,N_5940,N_5859);
nand U6142 (N_6142,N_5971,N_5978);
and U6143 (N_6143,N_5797,N_5928);
nor U6144 (N_6144,N_5861,N_5948);
xnor U6145 (N_6145,N_5945,N_5840);
or U6146 (N_6146,N_5788,N_5947);
or U6147 (N_6147,N_5897,N_5872);
nor U6148 (N_6148,N_5947,N_5881);
xnor U6149 (N_6149,N_5866,N_5984);
xnor U6150 (N_6150,N_5775,N_5850);
and U6151 (N_6151,N_5911,N_5796);
nor U6152 (N_6152,N_5864,N_5874);
nand U6153 (N_6153,N_5985,N_5874);
and U6154 (N_6154,N_5780,N_5757);
or U6155 (N_6155,N_5759,N_5949);
xor U6156 (N_6156,N_5902,N_5936);
or U6157 (N_6157,N_5950,N_5762);
nand U6158 (N_6158,N_5855,N_5980);
nand U6159 (N_6159,N_5930,N_5931);
xnor U6160 (N_6160,N_5859,N_5834);
nand U6161 (N_6161,N_5880,N_5953);
and U6162 (N_6162,N_5898,N_5871);
and U6163 (N_6163,N_5867,N_5955);
nor U6164 (N_6164,N_5819,N_5909);
xor U6165 (N_6165,N_5842,N_5960);
and U6166 (N_6166,N_5832,N_5776);
xnor U6167 (N_6167,N_5906,N_5942);
and U6168 (N_6168,N_5991,N_5911);
nand U6169 (N_6169,N_5982,N_5751);
nor U6170 (N_6170,N_5883,N_5764);
nand U6171 (N_6171,N_5966,N_5895);
nor U6172 (N_6172,N_5992,N_5841);
and U6173 (N_6173,N_5815,N_5912);
nor U6174 (N_6174,N_5818,N_5858);
and U6175 (N_6175,N_5837,N_5903);
nand U6176 (N_6176,N_5953,N_5763);
xor U6177 (N_6177,N_5968,N_5936);
nand U6178 (N_6178,N_5860,N_5901);
nand U6179 (N_6179,N_5832,N_5904);
nor U6180 (N_6180,N_5864,N_5826);
and U6181 (N_6181,N_5876,N_5957);
nor U6182 (N_6182,N_5956,N_5970);
nor U6183 (N_6183,N_5973,N_5972);
or U6184 (N_6184,N_5818,N_5985);
or U6185 (N_6185,N_5892,N_5887);
or U6186 (N_6186,N_5817,N_5814);
xor U6187 (N_6187,N_5812,N_5957);
or U6188 (N_6188,N_5950,N_5812);
nand U6189 (N_6189,N_5831,N_5977);
xnor U6190 (N_6190,N_5947,N_5928);
nor U6191 (N_6191,N_5940,N_5773);
and U6192 (N_6192,N_5776,N_5807);
nor U6193 (N_6193,N_5936,N_5816);
xnor U6194 (N_6194,N_5893,N_5897);
and U6195 (N_6195,N_5801,N_5836);
xor U6196 (N_6196,N_5944,N_5959);
or U6197 (N_6197,N_5864,N_5920);
and U6198 (N_6198,N_5995,N_5821);
xnor U6199 (N_6199,N_5831,N_5783);
or U6200 (N_6200,N_5805,N_5939);
nor U6201 (N_6201,N_5970,N_5777);
and U6202 (N_6202,N_5784,N_5907);
xor U6203 (N_6203,N_5813,N_5846);
and U6204 (N_6204,N_5918,N_5985);
xor U6205 (N_6205,N_5944,N_5810);
nor U6206 (N_6206,N_5773,N_5905);
nor U6207 (N_6207,N_5809,N_5925);
xnor U6208 (N_6208,N_5757,N_5967);
and U6209 (N_6209,N_5753,N_5851);
or U6210 (N_6210,N_5869,N_5866);
or U6211 (N_6211,N_5806,N_5918);
or U6212 (N_6212,N_5794,N_5904);
nor U6213 (N_6213,N_5767,N_5764);
xnor U6214 (N_6214,N_5754,N_5934);
nand U6215 (N_6215,N_5860,N_5937);
and U6216 (N_6216,N_5966,N_5893);
and U6217 (N_6217,N_5879,N_5903);
xor U6218 (N_6218,N_5800,N_5892);
or U6219 (N_6219,N_5789,N_5896);
and U6220 (N_6220,N_5816,N_5884);
and U6221 (N_6221,N_5984,N_5905);
xor U6222 (N_6222,N_5917,N_5864);
nand U6223 (N_6223,N_5974,N_5786);
or U6224 (N_6224,N_5896,N_5776);
xor U6225 (N_6225,N_5920,N_5887);
nor U6226 (N_6226,N_5789,N_5908);
nor U6227 (N_6227,N_5822,N_5970);
nand U6228 (N_6228,N_5925,N_5759);
xnor U6229 (N_6229,N_5979,N_5806);
nor U6230 (N_6230,N_5874,N_5883);
xor U6231 (N_6231,N_5794,N_5907);
xor U6232 (N_6232,N_5849,N_5985);
xnor U6233 (N_6233,N_5985,N_5960);
or U6234 (N_6234,N_5979,N_5853);
and U6235 (N_6235,N_5956,N_5766);
nand U6236 (N_6236,N_5835,N_5819);
and U6237 (N_6237,N_5793,N_5868);
xnor U6238 (N_6238,N_5970,N_5856);
and U6239 (N_6239,N_5782,N_5899);
xor U6240 (N_6240,N_5918,N_5916);
xnor U6241 (N_6241,N_5772,N_5993);
nand U6242 (N_6242,N_5830,N_5851);
xor U6243 (N_6243,N_5959,N_5763);
or U6244 (N_6244,N_5826,N_5912);
or U6245 (N_6245,N_5987,N_5903);
xnor U6246 (N_6246,N_5762,N_5895);
xor U6247 (N_6247,N_5806,N_5773);
nand U6248 (N_6248,N_5894,N_5927);
nor U6249 (N_6249,N_5818,N_5871);
nand U6250 (N_6250,N_6110,N_6103);
xor U6251 (N_6251,N_6173,N_6165);
nand U6252 (N_6252,N_6037,N_6137);
nor U6253 (N_6253,N_6162,N_6062);
nor U6254 (N_6254,N_6152,N_6247);
xnor U6255 (N_6255,N_6028,N_6190);
nor U6256 (N_6256,N_6217,N_6083);
nand U6257 (N_6257,N_6229,N_6241);
nor U6258 (N_6258,N_6038,N_6199);
and U6259 (N_6259,N_6196,N_6139);
and U6260 (N_6260,N_6090,N_6091);
nand U6261 (N_6261,N_6182,N_6202);
nor U6262 (N_6262,N_6086,N_6054);
or U6263 (N_6263,N_6140,N_6027);
or U6264 (N_6264,N_6016,N_6188);
and U6265 (N_6265,N_6204,N_6058);
nor U6266 (N_6266,N_6120,N_6078);
nor U6267 (N_6267,N_6242,N_6208);
nand U6268 (N_6268,N_6019,N_6092);
and U6269 (N_6269,N_6003,N_6117);
or U6270 (N_6270,N_6187,N_6213);
or U6271 (N_6271,N_6100,N_6222);
and U6272 (N_6272,N_6101,N_6146);
nand U6273 (N_6273,N_6061,N_6015);
or U6274 (N_6274,N_6226,N_6025);
nand U6275 (N_6275,N_6144,N_6109);
or U6276 (N_6276,N_6115,N_6236);
and U6277 (N_6277,N_6148,N_6057);
xor U6278 (N_6278,N_6046,N_6104);
nor U6279 (N_6279,N_6067,N_6099);
and U6280 (N_6280,N_6200,N_6131);
nand U6281 (N_6281,N_6237,N_6158);
and U6282 (N_6282,N_6167,N_6020);
xnor U6283 (N_6283,N_6042,N_6193);
or U6284 (N_6284,N_6160,N_6141);
xnor U6285 (N_6285,N_6002,N_6218);
nand U6286 (N_6286,N_6001,N_6068);
nand U6287 (N_6287,N_6221,N_6201);
or U6288 (N_6288,N_6230,N_6189);
nor U6289 (N_6289,N_6047,N_6079);
or U6290 (N_6290,N_6235,N_6031);
or U6291 (N_6291,N_6000,N_6082);
nand U6292 (N_6292,N_6097,N_6178);
nand U6293 (N_6293,N_6024,N_6192);
nand U6294 (N_6294,N_6069,N_6014);
and U6295 (N_6295,N_6026,N_6071);
xor U6296 (N_6296,N_6053,N_6183);
or U6297 (N_6297,N_6040,N_6012);
nor U6298 (N_6298,N_6116,N_6070);
or U6299 (N_6299,N_6239,N_6179);
nand U6300 (N_6300,N_6170,N_6008);
and U6301 (N_6301,N_6154,N_6045);
xor U6302 (N_6302,N_6050,N_6007);
or U6303 (N_6303,N_6233,N_6246);
nand U6304 (N_6304,N_6072,N_6084);
nand U6305 (N_6305,N_6123,N_6171);
nor U6306 (N_6306,N_6075,N_6030);
xnor U6307 (N_6307,N_6074,N_6186);
nor U6308 (N_6308,N_6177,N_6168);
or U6309 (N_6309,N_6087,N_6238);
or U6310 (N_6310,N_6005,N_6094);
nor U6311 (N_6311,N_6107,N_6039);
nor U6312 (N_6312,N_6064,N_6106);
xor U6313 (N_6313,N_6081,N_6108);
nand U6314 (N_6314,N_6102,N_6210);
nor U6315 (N_6315,N_6049,N_6234);
and U6316 (N_6316,N_6125,N_6129);
and U6317 (N_6317,N_6011,N_6142);
nor U6318 (N_6318,N_6176,N_6051);
xnor U6319 (N_6319,N_6017,N_6029);
nor U6320 (N_6320,N_6052,N_6044);
nand U6321 (N_6321,N_6243,N_6043);
nor U6322 (N_6322,N_6164,N_6198);
nand U6323 (N_6323,N_6130,N_6076);
or U6324 (N_6324,N_6112,N_6227);
or U6325 (N_6325,N_6180,N_6157);
or U6326 (N_6326,N_6105,N_6095);
or U6327 (N_6327,N_6041,N_6004);
or U6328 (N_6328,N_6127,N_6207);
nand U6329 (N_6329,N_6018,N_6195);
or U6330 (N_6330,N_6184,N_6248);
or U6331 (N_6331,N_6118,N_6169);
nor U6332 (N_6332,N_6175,N_6132);
or U6333 (N_6333,N_6096,N_6205);
and U6334 (N_6334,N_6066,N_6077);
or U6335 (N_6335,N_6006,N_6151);
xor U6336 (N_6336,N_6224,N_6089);
nand U6337 (N_6337,N_6145,N_6048);
or U6338 (N_6338,N_6060,N_6035);
or U6339 (N_6339,N_6220,N_6065);
and U6340 (N_6340,N_6055,N_6216);
nand U6341 (N_6341,N_6240,N_6085);
xor U6342 (N_6342,N_6022,N_6033);
nor U6343 (N_6343,N_6172,N_6021);
xnor U6344 (N_6344,N_6155,N_6114);
nor U6345 (N_6345,N_6034,N_6009);
nor U6346 (N_6346,N_6244,N_6219);
or U6347 (N_6347,N_6163,N_6203);
or U6348 (N_6348,N_6249,N_6150);
nor U6349 (N_6349,N_6211,N_6093);
nand U6350 (N_6350,N_6161,N_6063);
nor U6351 (N_6351,N_6194,N_6225);
and U6352 (N_6352,N_6088,N_6159);
and U6353 (N_6353,N_6098,N_6128);
nor U6354 (N_6354,N_6138,N_6174);
nor U6355 (N_6355,N_6056,N_6080);
xor U6356 (N_6356,N_6124,N_6149);
xor U6357 (N_6357,N_6228,N_6136);
and U6358 (N_6358,N_6111,N_6166);
or U6359 (N_6359,N_6143,N_6119);
or U6360 (N_6360,N_6134,N_6232);
xnor U6361 (N_6361,N_6113,N_6059);
nand U6362 (N_6362,N_6036,N_6206);
nand U6363 (N_6363,N_6032,N_6013);
and U6364 (N_6364,N_6126,N_6122);
xor U6365 (N_6365,N_6073,N_6135);
or U6366 (N_6366,N_6147,N_6156);
nand U6367 (N_6367,N_6023,N_6181);
nor U6368 (N_6368,N_6245,N_6010);
and U6369 (N_6369,N_6133,N_6153);
or U6370 (N_6370,N_6191,N_6212);
nor U6371 (N_6371,N_6214,N_6185);
nor U6372 (N_6372,N_6223,N_6121);
and U6373 (N_6373,N_6215,N_6209);
nor U6374 (N_6374,N_6231,N_6197);
and U6375 (N_6375,N_6130,N_6121);
nand U6376 (N_6376,N_6027,N_6086);
nor U6377 (N_6377,N_6111,N_6070);
nor U6378 (N_6378,N_6012,N_6074);
nor U6379 (N_6379,N_6171,N_6155);
nor U6380 (N_6380,N_6118,N_6014);
or U6381 (N_6381,N_6036,N_6081);
xnor U6382 (N_6382,N_6043,N_6087);
nand U6383 (N_6383,N_6160,N_6071);
or U6384 (N_6384,N_6134,N_6123);
or U6385 (N_6385,N_6187,N_6212);
nor U6386 (N_6386,N_6014,N_6083);
and U6387 (N_6387,N_6042,N_6146);
and U6388 (N_6388,N_6137,N_6164);
nor U6389 (N_6389,N_6052,N_6160);
or U6390 (N_6390,N_6058,N_6139);
and U6391 (N_6391,N_6175,N_6198);
or U6392 (N_6392,N_6088,N_6152);
xnor U6393 (N_6393,N_6031,N_6075);
nor U6394 (N_6394,N_6085,N_6248);
xor U6395 (N_6395,N_6012,N_6127);
nand U6396 (N_6396,N_6162,N_6227);
or U6397 (N_6397,N_6247,N_6030);
xnor U6398 (N_6398,N_6049,N_6123);
or U6399 (N_6399,N_6203,N_6193);
nor U6400 (N_6400,N_6129,N_6131);
nand U6401 (N_6401,N_6048,N_6198);
xor U6402 (N_6402,N_6084,N_6193);
or U6403 (N_6403,N_6185,N_6211);
and U6404 (N_6404,N_6086,N_6058);
nand U6405 (N_6405,N_6171,N_6234);
xor U6406 (N_6406,N_6193,N_6064);
nand U6407 (N_6407,N_6009,N_6021);
and U6408 (N_6408,N_6058,N_6162);
nand U6409 (N_6409,N_6113,N_6241);
nor U6410 (N_6410,N_6184,N_6140);
nor U6411 (N_6411,N_6021,N_6174);
nor U6412 (N_6412,N_6248,N_6022);
xor U6413 (N_6413,N_6028,N_6206);
xor U6414 (N_6414,N_6202,N_6240);
nor U6415 (N_6415,N_6118,N_6238);
nand U6416 (N_6416,N_6200,N_6221);
or U6417 (N_6417,N_6164,N_6235);
and U6418 (N_6418,N_6203,N_6142);
or U6419 (N_6419,N_6240,N_6204);
and U6420 (N_6420,N_6028,N_6148);
nand U6421 (N_6421,N_6086,N_6064);
nor U6422 (N_6422,N_6221,N_6094);
or U6423 (N_6423,N_6125,N_6034);
xnor U6424 (N_6424,N_6072,N_6207);
and U6425 (N_6425,N_6136,N_6008);
nor U6426 (N_6426,N_6187,N_6085);
xor U6427 (N_6427,N_6105,N_6201);
or U6428 (N_6428,N_6171,N_6104);
nand U6429 (N_6429,N_6075,N_6003);
nand U6430 (N_6430,N_6031,N_6009);
or U6431 (N_6431,N_6139,N_6010);
and U6432 (N_6432,N_6003,N_6157);
and U6433 (N_6433,N_6052,N_6233);
nor U6434 (N_6434,N_6118,N_6153);
nor U6435 (N_6435,N_6012,N_6195);
and U6436 (N_6436,N_6144,N_6067);
nand U6437 (N_6437,N_6231,N_6243);
or U6438 (N_6438,N_6043,N_6026);
or U6439 (N_6439,N_6164,N_6196);
or U6440 (N_6440,N_6162,N_6198);
and U6441 (N_6441,N_6088,N_6229);
or U6442 (N_6442,N_6168,N_6238);
or U6443 (N_6443,N_6227,N_6215);
nand U6444 (N_6444,N_6165,N_6025);
and U6445 (N_6445,N_6078,N_6129);
nor U6446 (N_6446,N_6117,N_6103);
and U6447 (N_6447,N_6098,N_6001);
and U6448 (N_6448,N_6235,N_6161);
nand U6449 (N_6449,N_6013,N_6198);
or U6450 (N_6450,N_6242,N_6107);
and U6451 (N_6451,N_6187,N_6232);
nor U6452 (N_6452,N_6228,N_6139);
or U6453 (N_6453,N_6098,N_6123);
nor U6454 (N_6454,N_6176,N_6126);
nor U6455 (N_6455,N_6004,N_6037);
nand U6456 (N_6456,N_6011,N_6085);
nand U6457 (N_6457,N_6075,N_6167);
or U6458 (N_6458,N_6202,N_6020);
nor U6459 (N_6459,N_6141,N_6214);
and U6460 (N_6460,N_6016,N_6220);
and U6461 (N_6461,N_6164,N_6131);
nor U6462 (N_6462,N_6116,N_6203);
nand U6463 (N_6463,N_6193,N_6229);
xnor U6464 (N_6464,N_6006,N_6226);
xor U6465 (N_6465,N_6209,N_6022);
nor U6466 (N_6466,N_6056,N_6096);
and U6467 (N_6467,N_6215,N_6047);
or U6468 (N_6468,N_6222,N_6201);
nor U6469 (N_6469,N_6223,N_6173);
xor U6470 (N_6470,N_6077,N_6025);
and U6471 (N_6471,N_6128,N_6135);
and U6472 (N_6472,N_6148,N_6097);
nor U6473 (N_6473,N_6156,N_6054);
xor U6474 (N_6474,N_6200,N_6223);
or U6475 (N_6475,N_6121,N_6096);
nor U6476 (N_6476,N_6017,N_6000);
nor U6477 (N_6477,N_6218,N_6195);
or U6478 (N_6478,N_6111,N_6010);
nand U6479 (N_6479,N_6112,N_6048);
xor U6480 (N_6480,N_6184,N_6038);
nor U6481 (N_6481,N_6151,N_6045);
xor U6482 (N_6482,N_6200,N_6160);
or U6483 (N_6483,N_6137,N_6150);
or U6484 (N_6484,N_6036,N_6113);
and U6485 (N_6485,N_6232,N_6248);
nor U6486 (N_6486,N_6156,N_6135);
nor U6487 (N_6487,N_6171,N_6188);
nor U6488 (N_6488,N_6024,N_6199);
or U6489 (N_6489,N_6095,N_6184);
xor U6490 (N_6490,N_6191,N_6097);
nand U6491 (N_6491,N_6063,N_6206);
xnor U6492 (N_6492,N_6210,N_6154);
and U6493 (N_6493,N_6164,N_6108);
and U6494 (N_6494,N_6069,N_6170);
nor U6495 (N_6495,N_6193,N_6011);
nor U6496 (N_6496,N_6040,N_6232);
or U6497 (N_6497,N_6218,N_6246);
nand U6498 (N_6498,N_6120,N_6021);
or U6499 (N_6499,N_6195,N_6247);
xor U6500 (N_6500,N_6381,N_6427);
xor U6501 (N_6501,N_6287,N_6420);
nor U6502 (N_6502,N_6294,N_6293);
nand U6503 (N_6503,N_6378,N_6309);
or U6504 (N_6504,N_6360,N_6333);
or U6505 (N_6505,N_6313,N_6327);
and U6506 (N_6506,N_6410,N_6318);
and U6507 (N_6507,N_6397,N_6369);
and U6508 (N_6508,N_6489,N_6289);
nor U6509 (N_6509,N_6450,N_6371);
or U6510 (N_6510,N_6418,N_6492);
and U6511 (N_6511,N_6477,N_6292);
nor U6512 (N_6512,N_6376,N_6323);
and U6513 (N_6513,N_6373,N_6261);
or U6514 (N_6514,N_6411,N_6276);
nor U6515 (N_6515,N_6328,N_6298);
xor U6516 (N_6516,N_6312,N_6282);
nor U6517 (N_6517,N_6280,N_6403);
xnor U6518 (N_6518,N_6463,N_6361);
xor U6519 (N_6519,N_6429,N_6480);
nor U6520 (N_6520,N_6274,N_6315);
nand U6521 (N_6521,N_6324,N_6446);
nand U6522 (N_6522,N_6344,N_6299);
nor U6523 (N_6523,N_6445,N_6340);
or U6524 (N_6524,N_6406,N_6363);
and U6525 (N_6525,N_6488,N_6367);
and U6526 (N_6526,N_6329,N_6264);
xor U6527 (N_6527,N_6437,N_6354);
or U6528 (N_6528,N_6311,N_6314);
xor U6529 (N_6529,N_6356,N_6383);
and U6530 (N_6530,N_6382,N_6417);
xnor U6531 (N_6531,N_6422,N_6265);
or U6532 (N_6532,N_6468,N_6352);
xor U6533 (N_6533,N_6283,N_6442);
and U6534 (N_6534,N_6470,N_6370);
or U6535 (N_6535,N_6337,N_6375);
and U6536 (N_6536,N_6257,N_6472);
or U6537 (N_6537,N_6284,N_6320);
and U6538 (N_6538,N_6421,N_6399);
and U6539 (N_6539,N_6286,N_6485);
or U6540 (N_6540,N_6434,N_6270);
and U6541 (N_6541,N_6279,N_6338);
or U6542 (N_6542,N_6493,N_6304);
nand U6543 (N_6543,N_6347,N_6255);
and U6544 (N_6544,N_6390,N_6474);
xor U6545 (N_6545,N_6414,N_6362);
nand U6546 (N_6546,N_6321,N_6322);
xor U6547 (N_6547,N_6357,N_6343);
nand U6548 (N_6548,N_6325,N_6497);
nand U6549 (N_6549,N_6387,N_6316);
and U6550 (N_6550,N_6365,N_6425);
or U6551 (N_6551,N_6359,N_6345);
nor U6552 (N_6552,N_6465,N_6455);
nand U6553 (N_6553,N_6405,N_6481);
or U6554 (N_6554,N_6300,N_6394);
xnor U6555 (N_6555,N_6440,N_6393);
and U6556 (N_6556,N_6395,N_6400);
nor U6557 (N_6557,N_6402,N_6253);
nand U6558 (N_6558,N_6346,N_6288);
xnor U6559 (N_6559,N_6460,N_6368);
nand U6560 (N_6560,N_6491,N_6419);
and U6561 (N_6561,N_6487,N_6475);
or U6562 (N_6562,N_6262,N_6266);
nand U6563 (N_6563,N_6388,N_6430);
xnor U6564 (N_6564,N_6296,N_6484);
nand U6565 (N_6565,N_6486,N_6438);
and U6566 (N_6566,N_6290,N_6379);
xor U6567 (N_6567,N_6331,N_6307);
nand U6568 (N_6568,N_6407,N_6416);
and U6569 (N_6569,N_6413,N_6495);
xor U6570 (N_6570,N_6389,N_6391);
or U6571 (N_6571,N_6490,N_6332);
nor U6572 (N_6572,N_6386,N_6432);
xnor U6573 (N_6573,N_6341,N_6431);
nor U6574 (N_6574,N_6401,N_6366);
xnor U6575 (N_6575,N_6269,N_6334);
nor U6576 (N_6576,N_6482,N_6272);
nor U6577 (N_6577,N_6424,N_6297);
or U6578 (N_6578,N_6295,N_6342);
or U6579 (N_6579,N_6336,N_6443);
or U6580 (N_6580,N_6412,N_6404);
and U6581 (N_6581,N_6499,N_6308);
nand U6582 (N_6582,N_6436,N_6317);
and U6583 (N_6583,N_6392,N_6351);
or U6584 (N_6584,N_6348,N_6374);
nand U6585 (N_6585,N_6372,N_6476);
xnor U6586 (N_6586,N_6330,N_6350);
or U6587 (N_6587,N_6415,N_6250);
nand U6588 (N_6588,N_6433,N_6451);
nor U6589 (N_6589,N_6306,N_6285);
or U6590 (N_6590,N_6498,N_6483);
nand U6591 (N_6591,N_6467,N_6478);
or U6592 (N_6592,N_6471,N_6385);
or U6593 (N_6593,N_6268,N_6408);
nand U6594 (N_6594,N_6259,N_6358);
or U6595 (N_6595,N_6278,N_6380);
nand U6596 (N_6596,N_6252,N_6339);
or U6597 (N_6597,N_6251,N_6423);
or U6598 (N_6598,N_6310,N_6409);
nand U6599 (N_6599,N_6447,N_6258);
or U6600 (N_6600,N_6275,N_6454);
and U6601 (N_6601,N_6444,N_6301);
or U6602 (N_6602,N_6466,N_6494);
xnor U6603 (N_6603,N_6459,N_6441);
nor U6604 (N_6604,N_6353,N_6435);
or U6605 (N_6605,N_6398,N_6326);
or U6606 (N_6606,N_6267,N_6254);
or U6607 (N_6607,N_6469,N_6349);
and U6608 (N_6608,N_6384,N_6473);
or U6609 (N_6609,N_6462,N_6291);
xor U6610 (N_6610,N_6335,N_6457);
nand U6611 (N_6611,N_6426,N_6271);
xnor U6612 (N_6612,N_6260,N_6355);
and U6613 (N_6613,N_6303,N_6439);
xor U6614 (N_6614,N_6302,N_6319);
nand U6615 (N_6615,N_6305,N_6377);
nor U6616 (N_6616,N_6479,N_6456);
xnor U6617 (N_6617,N_6496,N_6453);
nor U6618 (N_6618,N_6364,N_6263);
and U6619 (N_6619,N_6449,N_6273);
nand U6620 (N_6620,N_6428,N_6277);
and U6621 (N_6621,N_6396,N_6256);
or U6622 (N_6622,N_6448,N_6458);
nor U6623 (N_6623,N_6281,N_6464);
or U6624 (N_6624,N_6452,N_6461);
nor U6625 (N_6625,N_6335,N_6444);
or U6626 (N_6626,N_6450,N_6428);
and U6627 (N_6627,N_6396,N_6266);
nand U6628 (N_6628,N_6383,N_6373);
or U6629 (N_6629,N_6460,N_6476);
or U6630 (N_6630,N_6492,N_6261);
nor U6631 (N_6631,N_6399,N_6251);
and U6632 (N_6632,N_6385,N_6451);
or U6633 (N_6633,N_6398,N_6289);
and U6634 (N_6634,N_6475,N_6363);
xor U6635 (N_6635,N_6436,N_6354);
and U6636 (N_6636,N_6318,N_6265);
nand U6637 (N_6637,N_6430,N_6263);
nor U6638 (N_6638,N_6450,N_6447);
or U6639 (N_6639,N_6371,N_6416);
nor U6640 (N_6640,N_6257,N_6297);
nor U6641 (N_6641,N_6342,N_6485);
or U6642 (N_6642,N_6453,N_6393);
xor U6643 (N_6643,N_6367,N_6408);
or U6644 (N_6644,N_6333,N_6303);
xor U6645 (N_6645,N_6267,N_6344);
and U6646 (N_6646,N_6302,N_6442);
nor U6647 (N_6647,N_6295,N_6291);
or U6648 (N_6648,N_6274,N_6472);
and U6649 (N_6649,N_6283,N_6259);
and U6650 (N_6650,N_6479,N_6289);
nor U6651 (N_6651,N_6430,N_6260);
or U6652 (N_6652,N_6420,N_6350);
xnor U6653 (N_6653,N_6285,N_6462);
nor U6654 (N_6654,N_6481,N_6407);
xnor U6655 (N_6655,N_6463,N_6467);
nor U6656 (N_6656,N_6270,N_6421);
nand U6657 (N_6657,N_6378,N_6252);
nand U6658 (N_6658,N_6473,N_6252);
or U6659 (N_6659,N_6489,N_6440);
nor U6660 (N_6660,N_6281,N_6361);
and U6661 (N_6661,N_6349,N_6389);
nand U6662 (N_6662,N_6373,N_6264);
nor U6663 (N_6663,N_6487,N_6451);
nor U6664 (N_6664,N_6380,N_6326);
nand U6665 (N_6665,N_6414,N_6377);
and U6666 (N_6666,N_6314,N_6386);
xnor U6667 (N_6667,N_6405,N_6415);
nor U6668 (N_6668,N_6353,N_6266);
or U6669 (N_6669,N_6336,N_6325);
or U6670 (N_6670,N_6437,N_6499);
nand U6671 (N_6671,N_6485,N_6361);
nand U6672 (N_6672,N_6297,N_6460);
xor U6673 (N_6673,N_6418,N_6471);
xor U6674 (N_6674,N_6261,N_6385);
and U6675 (N_6675,N_6445,N_6390);
xnor U6676 (N_6676,N_6315,N_6393);
nor U6677 (N_6677,N_6250,N_6431);
nand U6678 (N_6678,N_6372,N_6449);
or U6679 (N_6679,N_6356,N_6308);
and U6680 (N_6680,N_6477,N_6327);
or U6681 (N_6681,N_6455,N_6282);
or U6682 (N_6682,N_6483,N_6365);
or U6683 (N_6683,N_6453,N_6296);
and U6684 (N_6684,N_6269,N_6363);
and U6685 (N_6685,N_6287,N_6486);
xnor U6686 (N_6686,N_6266,N_6441);
or U6687 (N_6687,N_6457,N_6448);
nand U6688 (N_6688,N_6401,N_6411);
and U6689 (N_6689,N_6265,N_6335);
or U6690 (N_6690,N_6363,N_6337);
nor U6691 (N_6691,N_6296,N_6440);
nor U6692 (N_6692,N_6287,N_6475);
xor U6693 (N_6693,N_6399,N_6436);
nor U6694 (N_6694,N_6361,N_6367);
nor U6695 (N_6695,N_6419,N_6387);
and U6696 (N_6696,N_6335,N_6488);
or U6697 (N_6697,N_6456,N_6278);
or U6698 (N_6698,N_6342,N_6419);
and U6699 (N_6699,N_6310,N_6340);
or U6700 (N_6700,N_6422,N_6297);
or U6701 (N_6701,N_6410,N_6365);
xor U6702 (N_6702,N_6448,N_6347);
nor U6703 (N_6703,N_6424,N_6280);
nand U6704 (N_6704,N_6478,N_6396);
xor U6705 (N_6705,N_6378,N_6448);
and U6706 (N_6706,N_6332,N_6413);
or U6707 (N_6707,N_6457,N_6325);
nor U6708 (N_6708,N_6455,N_6275);
nand U6709 (N_6709,N_6393,N_6452);
nor U6710 (N_6710,N_6472,N_6292);
and U6711 (N_6711,N_6343,N_6391);
or U6712 (N_6712,N_6418,N_6304);
and U6713 (N_6713,N_6452,N_6289);
and U6714 (N_6714,N_6421,N_6309);
and U6715 (N_6715,N_6273,N_6488);
nor U6716 (N_6716,N_6275,N_6258);
and U6717 (N_6717,N_6479,N_6345);
xor U6718 (N_6718,N_6327,N_6445);
and U6719 (N_6719,N_6437,N_6458);
nand U6720 (N_6720,N_6423,N_6374);
or U6721 (N_6721,N_6274,N_6341);
and U6722 (N_6722,N_6484,N_6337);
and U6723 (N_6723,N_6414,N_6422);
and U6724 (N_6724,N_6454,N_6311);
nand U6725 (N_6725,N_6455,N_6437);
xor U6726 (N_6726,N_6404,N_6463);
and U6727 (N_6727,N_6396,N_6267);
xor U6728 (N_6728,N_6409,N_6330);
or U6729 (N_6729,N_6317,N_6397);
or U6730 (N_6730,N_6380,N_6448);
and U6731 (N_6731,N_6476,N_6485);
and U6732 (N_6732,N_6295,N_6424);
xnor U6733 (N_6733,N_6284,N_6396);
xnor U6734 (N_6734,N_6433,N_6350);
nor U6735 (N_6735,N_6454,N_6315);
or U6736 (N_6736,N_6455,N_6397);
nor U6737 (N_6737,N_6295,N_6254);
or U6738 (N_6738,N_6389,N_6403);
nor U6739 (N_6739,N_6253,N_6423);
and U6740 (N_6740,N_6326,N_6378);
nor U6741 (N_6741,N_6321,N_6251);
nor U6742 (N_6742,N_6267,N_6484);
or U6743 (N_6743,N_6357,N_6487);
nor U6744 (N_6744,N_6429,N_6323);
and U6745 (N_6745,N_6443,N_6426);
xnor U6746 (N_6746,N_6342,N_6297);
or U6747 (N_6747,N_6290,N_6309);
nor U6748 (N_6748,N_6412,N_6449);
or U6749 (N_6749,N_6284,N_6421);
or U6750 (N_6750,N_6602,N_6685);
nor U6751 (N_6751,N_6726,N_6744);
nor U6752 (N_6752,N_6672,N_6617);
nand U6753 (N_6753,N_6552,N_6700);
xnor U6754 (N_6754,N_6671,N_6631);
or U6755 (N_6755,N_6598,N_6544);
and U6756 (N_6756,N_6662,N_6718);
and U6757 (N_6757,N_6524,N_6574);
nand U6758 (N_6758,N_6500,N_6695);
or U6759 (N_6759,N_6710,N_6706);
and U6760 (N_6760,N_6721,N_6687);
nand U6761 (N_6761,N_6513,N_6593);
xnor U6762 (N_6762,N_6742,N_6656);
nand U6763 (N_6763,N_6545,N_6605);
nor U6764 (N_6764,N_6735,N_6741);
nor U6765 (N_6765,N_6573,N_6564);
nand U6766 (N_6766,N_6562,N_6578);
nor U6767 (N_6767,N_6746,N_6572);
nand U6768 (N_6768,N_6659,N_6576);
xor U6769 (N_6769,N_6575,N_6677);
xnor U6770 (N_6770,N_6546,N_6698);
nand U6771 (N_6771,N_6689,N_6679);
and U6772 (N_6772,N_6711,N_6604);
or U6773 (N_6773,N_6648,N_6702);
or U6774 (N_6774,N_6723,N_6673);
nand U6775 (N_6775,N_6590,N_6684);
nor U6776 (N_6776,N_6682,N_6503);
nand U6777 (N_6777,N_6534,N_6600);
or U6778 (N_6778,N_6589,N_6577);
nand U6779 (N_6779,N_6618,N_6733);
or U6780 (N_6780,N_6611,N_6712);
nand U6781 (N_6781,N_6643,N_6529);
and U6782 (N_6782,N_6620,N_6654);
xnor U6783 (N_6783,N_6606,N_6715);
or U6784 (N_6784,N_6616,N_6716);
and U6785 (N_6785,N_6555,N_6632);
and U6786 (N_6786,N_6699,N_6688);
xor U6787 (N_6787,N_6686,N_6506);
xor U6788 (N_6788,N_6514,N_6732);
or U6789 (N_6789,N_6502,N_6621);
or U6790 (N_6790,N_6515,N_6663);
or U6791 (N_6791,N_6557,N_6660);
nor U6792 (N_6792,N_6609,N_6717);
or U6793 (N_6793,N_6508,N_6597);
or U6794 (N_6794,N_6535,N_6638);
or U6795 (N_6795,N_6704,N_6678);
and U6796 (N_6796,N_6644,N_6667);
xor U6797 (N_6797,N_6640,N_6745);
and U6798 (N_6798,N_6665,N_6670);
nand U6799 (N_6799,N_6533,N_6691);
nor U6800 (N_6800,N_6683,N_6666);
or U6801 (N_6801,N_6720,N_6510);
xor U6802 (N_6802,N_6628,N_6520);
xor U6803 (N_6803,N_6626,N_6612);
nor U6804 (N_6804,N_6729,N_6675);
nand U6805 (N_6805,N_6650,N_6629);
nor U6806 (N_6806,N_6556,N_6630);
nor U6807 (N_6807,N_6610,N_6727);
nand U6808 (N_6808,N_6653,N_6748);
and U6809 (N_6809,N_6518,N_6747);
xnor U6810 (N_6810,N_6567,N_6669);
or U6811 (N_6811,N_6696,N_6581);
and U6812 (N_6812,N_6613,N_6724);
nand U6813 (N_6813,N_6505,N_6694);
and U6814 (N_6814,N_6588,N_6634);
nor U6815 (N_6815,N_6530,N_6594);
nor U6816 (N_6816,N_6693,N_6601);
or U6817 (N_6817,N_6708,N_6603);
xor U6818 (N_6818,N_6549,N_6587);
nor U6819 (N_6819,N_6658,N_6541);
nor U6820 (N_6820,N_6739,N_6560);
or U6821 (N_6821,N_6639,N_6730);
nor U6822 (N_6822,N_6615,N_6728);
and U6823 (N_6823,N_6550,N_6595);
xnor U6824 (N_6824,N_6501,N_6509);
or U6825 (N_6825,N_6516,N_6657);
or U6826 (N_6826,N_6540,N_6676);
xnor U6827 (N_6827,N_6583,N_6614);
nand U6828 (N_6828,N_6680,N_6517);
or U6829 (N_6829,N_6637,N_6553);
nand U6830 (N_6830,N_6649,N_6539);
nand U6831 (N_6831,N_6705,N_6543);
or U6832 (N_6832,N_6713,N_6625);
nand U6833 (N_6833,N_6738,N_6652);
xnor U6834 (N_6834,N_6547,N_6674);
and U6835 (N_6835,N_6647,N_6703);
and U6836 (N_6836,N_6627,N_6566);
xor U6837 (N_6837,N_6636,N_6664);
and U6838 (N_6838,N_6558,N_6707);
or U6839 (N_6839,N_6522,N_6641);
xor U6840 (N_6840,N_6519,N_6526);
nor U6841 (N_6841,N_6584,N_6661);
and U6842 (N_6842,N_6542,N_6525);
nand U6843 (N_6843,N_6697,N_6623);
nand U6844 (N_6844,N_6536,N_6521);
or U6845 (N_6845,N_6743,N_6528);
and U6846 (N_6846,N_6586,N_6511);
or U6847 (N_6847,N_6645,N_6563);
xor U6848 (N_6848,N_6531,N_6537);
and U6849 (N_6849,N_6635,N_6596);
nand U6850 (N_6850,N_6599,N_6668);
or U6851 (N_6851,N_6622,N_6607);
nand U6852 (N_6852,N_6538,N_6681);
xnor U6853 (N_6853,N_6619,N_6512);
and U6854 (N_6854,N_6507,N_6692);
nand U6855 (N_6855,N_6655,N_6570);
and U6856 (N_6856,N_6527,N_6737);
nor U6857 (N_6857,N_6701,N_6580);
and U6858 (N_6858,N_6719,N_6740);
or U6859 (N_6859,N_6709,N_6646);
and U6860 (N_6860,N_6736,N_6582);
xor U6861 (N_6861,N_6592,N_6633);
xor U6862 (N_6862,N_6714,N_6569);
nand U6863 (N_6863,N_6523,N_6749);
and U6864 (N_6864,N_6642,N_6725);
or U6865 (N_6865,N_6608,N_6551);
xnor U6866 (N_6866,N_6585,N_6734);
or U6867 (N_6867,N_6565,N_6731);
nor U6868 (N_6868,N_6624,N_6561);
or U6869 (N_6869,N_6690,N_6571);
or U6870 (N_6870,N_6554,N_6559);
xor U6871 (N_6871,N_6568,N_6651);
and U6872 (N_6872,N_6504,N_6591);
and U6873 (N_6873,N_6532,N_6548);
nor U6874 (N_6874,N_6579,N_6722);
xor U6875 (N_6875,N_6567,N_6708);
and U6876 (N_6876,N_6606,N_6595);
or U6877 (N_6877,N_6573,N_6555);
nor U6878 (N_6878,N_6561,N_6710);
xor U6879 (N_6879,N_6508,N_6577);
nand U6880 (N_6880,N_6725,N_6517);
xnor U6881 (N_6881,N_6597,N_6696);
and U6882 (N_6882,N_6619,N_6656);
nor U6883 (N_6883,N_6674,N_6609);
nor U6884 (N_6884,N_6729,N_6740);
nand U6885 (N_6885,N_6532,N_6666);
and U6886 (N_6886,N_6520,N_6644);
nand U6887 (N_6887,N_6511,N_6507);
xor U6888 (N_6888,N_6607,N_6588);
or U6889 (N_6889,N_6583,N_6561);
and U6890 (N_6890,N_6729,N_6529);
nand U6891 (N_6891,N_6564,N_6591);
and U6892 (N_6892,N_6615,N_6579);
nor U6893 (N_6893,N_6659,N_6667);
and U6894 (N_6894,N_6513,N_6551);
or U6895 (N_6895,N_6616,N_6737);
nand U6896 (N_6896,N_6685,N_6689);
nand U6897 (N_6897,N_6529,N_6646);
xor U6898 (N_6898,N_6743,N_6691);
or U6899 (N_6899,N_6593,N_6543);
and U6900 (N_6900,N_6651,N_6685);
nand U6901 (N_6901,N_6547,N_6725);
and U6902 (N_6902,N_6714,N_6533);
xnor U6903 (N_6903,N_6572,N_6655);
xnor U6904 (N_6904,N_6710,N_6679);
or U6905 (N_6905,N_6681,N_6545);
and U6906 (N_6906,N_6604,N_6542);
nor U6907 (N_6907,N_6646,N_6530);
or U6908 (N_6908,N_6519,N_6646);
or U6909 (N_6909,N_6691,N_6696);
xor U6910 (N_6910,N_6683,N_6576);
nand U6911 (N_6911,N_6523,N_6519);
and U6912 (N_6912,N_6569,N_6712);
nand U6913 (N_6913,N_6735,N_6686);
and U6914 (N_6914,N_6654,N_6594);
and U6915 (N_6915,N_6613,N_6572);
nor U6916 (N_6916,N_6702,N_6564);
and U6917 (N_6917,N_6513,N_6500);
or U6918 (N_6918,N_6577,N_6660);
xor U6919 (N_6919,N_6667,N_6617);
nor U6920 (N_6920,N_6667,N_6600);
xnor U6921 (N_6921,N_6630,N_6612);
or U6922 (N_6922,N_6731,N_6568);
and U6923 (N_6923,N_6537,N_6642);
nand U6924 (N_6924,N_6632,N_6668);
nor U6925 (N_6925,N_6520,N_6705);
nand U6926 (N_6926,N_6743,N_6537);
xnor U6927 (N_6927,N_6725,N_6743);
or U6928 (N_6928,N_6640,N_6672);
and U6929 (N_6929,N_6708,N_6523);
nor U6930 (N_6930,N_6524,N_6529);
nor U6931 (N_6931,N_6506,N_6584);
xnor U6932 (N_6932,N_6549,N_6703);
nor U6933 (N_6933,N_6584,N_6695);
or U6934 (N_6934,N_6668,N_6512);
xnor U6935 (N_6935,N_6722,N_6500);
and U6936 (N_6936,N_6629,N_6724);
nor U6937 (N_6937,N_6744,N_6677);
or U6938 (N_6938,N_6520,N_6560);
xnor U6939 (N_6939,N_6681,N_6610);
and U6940 (N_6940,N_6550,N_6649);
nor U6941 (N_6941,N_6604,N_6628);
xnor U6942 (N_6942,N_6510,N_6734);
xnor U6943 (N_6943,N_6726,N_6574);
and U6944 (N_6944,N_6688,N_6662);
or U6945 (N_6945,N_6621,N_6503);
nor U6946 (N_6946,N_6579,N_6660);
xnor U6947 (N_6947,N_6659,N_6542);
and U6948 (N_6948,N_6504,N_6737);
nor U6949 (N_6949,N_6616,N_6641);
or U6950 (N_6950,N_6565,N_6719);
nor U6951 (N_6951,N_6565,N_6597);
nor U6952 (N_6952,N_6567,N_6556);
or U6953 (N_6953,N_6537,N_6561);
nand U6954 (N_6954,N_6603,N_6700);
and U6955 (N_6955,N_6554,N_6546);
or U6956 (N_6956,N_6556,N_6687);
and U6957 (N_6957,N_6605,N_6509);
and U6958 (N_6958,N_6582,N_6502);
nand U6959 (N_6959,N_6714,N_6662);
nand U6960 (N_6960,N_6743,N_6731);
and U6961 (N_6961,N_6666,N_6628);
xor U6962 (N_6962,N_6634,N_6691);
and U6963 (N_6963,N_6583,N_6631);
xor U6964 (N_6964,N_6686,N_6647);
or U6965 (N_6965,N_6596,N_6653);
nor U6966 (N_6966,N_6552,N_6639);
and U6967 (N_6967,N_6555,N_6556);
nor U6968 (N_6968,N_6503,N_6623);
nand U6969 (N_6969,N_6644,N_6715);
or U6970 (N_6970,N_6579,N_6511);
xnor U6971 (N_6971,N_6701,N_6723);
xor U6972 (N_6972,N_6561,N_6687);
or U6973 (N_6973,N_6523,N_6718);
and U6974 (N_6974,N_6631,N_6593);
xor U6975 (N_6975,N_6543,N_6549);
nor U6976 (N_6976,N_6580,N_6542);
xnor U6977 (N_6977,N_6581,N_6653);
nor U6978 (N_6978,N_6527,N_6574);
nand U6979 (N_6979,N_6733,N_6648);
or U6980 (N_6980,N_6535,N_6692);
and U6981 (N_6981,N_6647,N_6639);
or U6982 (N_6982,N_6534,N_6660);
nor U6983 (N_6983,N_6621,N_6552);
and U6984 (N_6984,N_6552,N_6688);
or U6985 (N_6985,N_6618,N_6611);
nor U6986 (N_6986,N_6672,N_6634);
nor U6987 (N_6987,N_6530,N_6706);
and U6988 (N_6988,N_6612,N_6574);
xnor U6989 (N_6989,N_6714,N_6575);
or U6990 (N_6990,N_6546,N_6528);
xnor U6991 (N_6991,N_6723,N_6622);
or U6992 (N_6992,N_6616,N_6636);
or U6993 (N_6993,N_6692,N_6592);
and U6994 (N_6994,N_6656,N_6727);
xor U6995 (N_6995,N_6531,N_6570);
and U6996 (N_6996,N_6670,N_6632);
nor U6997 (N_6997,N_6619,N_6548);
nand U6998 (N_6998,N_6634,N_6579);
nand U6999 (N_6999,N_6577,N_6656);
xnor U7000 (N_7000,N_6766,N_6933);
xor U7001 (N_7001,N_6784,N_6946);
or U7002 (N_7002,N_6789,N_6776);
xor U7003 (N_7003,N_6992,N_6841);
nand U7004 (N_7004,N_6937,N_6932);
and U7005 (N_7005,N_6958,N_6983);
and U7006 (N_7006,N_6869,N_6904);
or U7007 (N_7007,N_6984,N_6837);
nor U7008 (N_7008,N_6876,N_6786);
nor U7009 (N_7009,N_6930,N_6763);
xor U7010 (N_7010,N_6927,N_6835);
nor U7011 (N_7011,N_6805,N_6795);
and U7012 (N_7012,N_6815,N_6808);
nor U7013 (N_7013,N_6890,N_6757);
xnor U7014 (N_7014,N_6911,N_6814);
xor U7015 (N_7015,N_6993,N_6909);
nor U7016 (N_7016,N_6793,N_6996);
nand U7017 (N_7017,N_6913,N_6752);
nand U7018 (N_7018,N_6981,N_6824);
nor U7019 (N_7019,N_6968,N_6885);
xor U7020 (N_7020,N_6751,N_6770);
nand U7021 (N_7021,N_6754,N_6920);
nor U7022 (N_7022,N_6926,N_6801);
or U7023 (N_7023,N_6857,N_6940);
nand U7024 (N_7024,N_6989,N_6846);
nor U7025 (N_7025,N_6887,N_6790);
xnor U7026 (N_7026,N_6922,N_6791);
and U7027 (N_7027,N_6759,N_6900);
and U7028 (N_7028,N_6907,N_6939);
xor U7029 (N_7029,N_6942,N_6921);
or U7030 (N_7030,N_6943,N_6768);
nand U7031 (N_7031,N_6951,N_6781);
or U7032 (N_7032,N_6800,N_6972);
nand U7033 (N_7033,N_6971,N_6832);
nor U7034 (N_7034,N_6892,N_6868);
or U7035 (N_7035,N_6818,N_6870);
nand U7036 (N_7036,N_6903,N_6894);
nor U7037 (N_7037,N_6965,N_6925);
or U7038 (N_7038,N_6947,N_6782);
xnor U7039 (N_7039,N_6838,N_6758);
nor U7040 (N_7040,N_6973,N_6901);
or U7041 (N_7041,N_6843,N_6998);
nand U7042 (N_7042,N_6982,N_6812);
and U7043 (N_7043,N_6883,N_6976);
xnor U7044 (N_7044,N_6941,N_6856);
and U7045 (N_7045,N_6773,N_6806);
or U7046 (N_7046,N_6803,N_6975);
nor U7047 (N_7047,N_6848,N_6986);
nor U7048 (N_7048,N_6798,N_6771);
or U7049 (N_7049,N_6817,N_6851);
nor U7050 (N_7050,N_6956,N_6961);
and U7051 (N_7051,N_6881,N_6915);
xnor U7052 (N_7052,N_6845,N_6750);
xor U7053 (N_7053,N_6767,N_6990);
or U7054 (N_7054,N_6966,N_6788);
and U7055 (N_7055,N_6978,N_6960);
or U7056 (N_7056,N_6809,N_6871);
xnor U7057 (N_7057,N_6955,N_6827);
nand U7058 (N_7058,N_6979,N_6760);
nor U7059 (N_7059,N_6830,N_6884);
or U7060 (N_7060,N_6948,N_6895);
nor U7061 (N_7061,N_6836,N_6755);
or U7062 (N_7062,N_6878,N_6874);
nor U7063 (N_7063,N_6792,N_6967);
xnor U7064 (N_7064,N_6822,N_6854);
xnor U7065 (N_7065,N_6852,N_6977);
and U7066 (N_7066,N_6834,N_6859);
xor U7067 (N_7067,N_6810,N_6825);
or U7068 (N_7068,N_6826,N_6844);
xnor U7069 (N_7069,N_6936,N_6811);
xnor U7070 (N_7070,N_6753,N_6823);
nor U7071 (N_7071,N_6945,N_6858);
xor U7072 (N_7072,N_6860,N_6863);
or U7073 (N_7073,N_6917,N_6774);
nand U7074 (N_7074,N_6797,N_6764);
or U7075 (N_7075,N_6756,N_6987);
nand U7076 (N_7076,N_6957,N_6866);
and U7077 (N_7077,N_6910,N_6783);
nor U7078 (N_7078,N_6928,N_6873);
or U7079 (N_7079,N_6938,N_6898);
nor U7080 (N_7080,N_6829,N_6761);
nand U7081 (N_7081,N_6912,N_6861);
and U7082 (N_7082,N_6799,N_6879);
or U7083 (N_7083,N_6902,N_6880);
nor U7084 (N_7084,N_6905,N_6980);
nor U7085 (N_7085,N_6850,N_6787);
nor U7086 (N_7086,N_6842,N_6923);
and U7087 (N_7087,N_6855,N_6916);
and U7088 (N_7088,N_6862,N_6991);
and U7089 (N_7089,N_6821,N_6819);
or U7090 (N_7090,N_6853,N_6962);
or U7091 (N_7091,N_6974,N_6995);
nand U7092 (N_7092,N_6908,N_6919);
nor U7093 (N_7093,N_6839,N_6796);
and U7094 (N_7094,N_6867,N_6899);
nand U7095 (N_7095,N_6999,N_6762);
and U7096 (N_7096,N_6875,N_6831);
nor U7097 (N_7097,N_6775,N_6804);
and U7098 (N_7098,N_6802,N_6954);
xnor U7099 (N_7099,N_6931,N_6849);
nand U7100 (N_7100,N_6944,N_6906);
nand U7101 (N_7101,N_6877,N_6865);
nand U7102 (N_7102,N_6780,N_6779);
nand U7103 (N_7103,N_6949,N_6772);
or U7104 (N_7104,N_6886,N_6769);
nand U7105 (N_7105,N_6813,N_6882);
xnor U7106 (N_7106,N_6970,N_6765);
nor U7107 (N_7107,N_6896,N_6816);
nand U7108 (N_7108,N_6988,N_6833);
or U7109 (N_7109,N_6914,N_6964);
xor U7110 (N_7110,N_6794,N_6847);
nor U7111 (N_7111,N_6994,N_6889);
nor U7112 (N_7112,N_6924,N_6820);
or U7113 (N_7113,N_6959,N_6935);
and U7114 (N_7114,N_6934,N_6985);
xor U7115 (N_7115,N_6963,N_6918);
nand U7116 (N_7116,N_6893,N_6777);
xor U7117 (N_7117,N_6840,N_6953);
or U7118 (N_7118,N_6888,N_6929);
nor U7119 (N_7119,N_6950,N_6997);
nand U7120 (N_7120,N_6891,N_6872);
or U7121 (N_7121,N_6785,N_6969);
and U7122 (N_7122,N_6778,N_6807);
nand U7123 (N_7123,N_6828,N_6897);
xor U7124 (N_7124,N_6952,N_6864);
or U7125 (N_7125,N_6955,N_6835);
or U7126 (N_7126,N_6754,N_6777);
xnor U7127 (N_7127,N_6934,N_6944);
nand U7128 (N_7128,N_6983,N_6896);
or U7129 (N_7129,N_6890,N_6826);
or U7130 (N_7130,N_6843,N_6993);
nand U7131 (N_7131,N_6950,N_6974);
nor U7132 (N_7132,N_6782,N_6975);
xnor U7133 (N_7133,N_6930,N_6953);
and U7134 (N_7134,N_6801,N_6800);
nor U7135 (N_7135,N_6832,N_6894);
nand U7136 (N_7136,N_6920,N_6936);
or U7137 (N_7137,N_6930,N_6802);
nor U7138 (N_7138,N_6828,N_6841);
or U7139 (N_7139,N_6790,N_6971);
nand U7140 (N_7140,N_6775,N_6876);
and U7141 (N_7141,N_6901,N_6778);
or U7142 (N_7142,N_6753,N_6765);
and U7143 (N_7143,N_6805,N_6784);
nand U7144 (N_7144,N_6891,N_6904);
nand U7145 (N_7145,N_6774,N_6902);
or U7146 (N_7146,N_6919,N_6871);
or U7147 (N_7147,N_6829,N_6780);
nor U7148 (N_7148,N_6996,N_6983);
xor U7149 (N_7149,N_6798,N_6896);
nand U7150 (N_7150,N_6814,N_6756);
nor U7151 (N_7151,N_6923,N_6799);
nand U7152 (N_7152,N_6985,N_6949);
nor U7153 (N_7153,N_6929,N_6753);
and U7154 (N_7154,N_6894,N_6841);
nand U7155 (N_7155,N_6876,N_6947);
xnor U7156 (N_7156,N_6790,N_6938);
or U7157 (N_7157,N_6786,N_6958);
or U7158 (N_7158,N_6853,N_6921);
nor U7159 (N_7159,N_6926,N_6920);
xor U7160 (N_7160,N_6909,N_6802);
and U7161 (N_7161,N_6808,N_6937);
and U7162 (N_7162,N_6973,N_6859);
nor U7163 (N_7163,N_6806,N_6780);
nand U7164 (N_7164,N_6765,N_6897);
nor U7165 (N_7165,N_6843,N_6852);
or U7166 (N_7166,N_6910,N_6942);
nand U7167 (N_7167,N_6773,N_6873);
or U7168 (N_7168,N_6789,N_6944);
nand U7169 (N_7169,N_6854,N_6980);
and U7170 (N_7170,N_6754,N_6994);
nand U7171 (N_7171,N_6878,N_6986);
nand U7172 (N_7172,N_6986,N_6812);
xnor U7173 (N_7173,N_6917,N_6929);
nor U7174 (N_7174,N_6925,N_6929);
nand U7175 (N_7175,N_6886,N_6877);
and U7176 (N_7176,N_6754,N_6846);
nand U7177 (N_7177,N_6874,N_6752);
nand U7178 (N_7178,N_6882,N_6852);
nand U7179 (N_7179,N_6786,N_6974);
or U7180 (N_7180,N_6790,N_6979);
or U7181 (N_7181,N_6831,N_6818);
and U7182 (N_7182,N_6932,N_6866);
or U7183 (N_7183,N_6997,N_6866);
or U7184 (N_7184,N_6768,N_6804);
nand U7185 (N_7185,N_6881,N_6963);
or U7186 (N_7186,N_6959,N_6967);
and U7187 (N_7187,N_6906,N_6957);
nand U7188 (N_7188,N_6919,N_6813);
xor U7189 (N_7189,N_6975,N_6907);
and U7190 (N_7190,N_6940,N_6844);
nor U7191 (N_7191,N_6815,N_6855);
and U7192 (N_7192,N_6913,N_6844);
or U7193 (N_7193,N_6966,N_6952);
nand U7194 (N_7194,N_6993,N_6937);
and U7195 (N_7195,N_6923,N_6926);
or U7196 (N_7196,N_6859,N_6928);
and U7197 (N_7197,N_6965,N_6828);
nor U7198 (N_7198,N_6884,N_6948);
xnor U7199 (N_7199,N_6821,N_6825);
and U7200 (N_7200,N_6945,N_6877);
nor U7201 (N_7201,N_6993,N_6964);
and U7202 (N_7202,N_6915,N_6832);
nor U7203 (N_7203,N_6830,N_6922);
xor U7204 (N_7204,N_6855,N_6989);
nor U7205 (N_7205,N_6790,N_6882);
xor U7206 (N_7206,N_6850,N_6840);
and U7207 (N_7207,N_6800,N_6765);
nand U7208 (N_7208,N_6942,N_6900);
nor U7209 (N_7209,N_6992,N_6973);
and U7210 (N_7210,N_6839,N_6852);
or U7211 (N_7211,N_6808,N_6977);
or U7212 (N_7212,N_6774,N_6956);
nor U7213 (N_7213,N_6757,N_6769);
or U7214 (N_7214,N_6873,N_6943);
nand U7215 (N_7215,N_6830,N_6991);
xnor U7216 (N_7216,N_6834,N_6825);
or U7217 (N_7217,N_6885,N_6776);
and U7218 (N_7218,N_6796,N_6928);
nor U7219 (N_7219,N_6874,N_6979);
and U7220 (N_7220,N_6772,N_6764);
and U7221 (N_7221,N_6788,N_6800);
nand U7222 (N_7222,N_6966,N_6789);
and U7223 (N_7223,N_6765,N_6987);
and U7224 (N_7224,N_6967,N_6762);
or U7225 (N_7225,N_6956,N_6928);
nand U7226 (N_7226,N_6838,N_6796);
nand U7227 (N_7227,N_6925,N_6776);
xor U7228 (N_7228,N_6943,N_6761);
and U7229 (N_7229,N_6853,N_6843);
nand U7230 (N_7230,N_6907,N_6851);
nand U7231 (N_7231,N_6982,N_6823);
or U7232 (N_7232,N_6774,N_6851);
nor U7233 (N_7233,N_6789,N_6869);
and U7234 (N_7234,N_6843,N_6807);
and U7235 (N_7235,N_6856,N_6921);
nor U7236 (N_7236,N_6771,N_6970);
or U7237 (N_7237,N_6878,N_6985);
and U7238 (N_7238,N_6985,N_6917);
or U7239 (N_7239,N_6756,N_6752);
or U7240 (N_7240,N_6908,N_6806);
nand U7241 (N_7241,N_6877,N_6833);
or U7242 (N_7242,N_6796,N_6871);
and U7243 (N_7243,N_6797,N_6855);
or U7244 (N_7244,N_6957,N_6832);
nand U7245 (N_7245,N_6938,N_6951);
or U7246 (N_7246,N_6844,N_6938);
or U7247 (N_7247,N_6808,N_6925);
or U7248 (N_7248,N_6836,N_6792);
nor U7249 (N_7249,N_6836,N_6868);
nor U7250 (N_7250,N_7049,N_7228);
nor U7251 (N_7251,N_7217,N_7074);
nor U7252 (N_7252,N_7161,N_7065);
nand U7253 (N_7253,N_7214,N_7023);
nand U7254 (N_7254,N_7156,N_7088);
or U7255 (N_7255,N_7116,N_7052);
nor U7256 (N_7256,N_7084,N_7095);
nor U7257 (N_7257,N_7097,N_7129);
or U7258 (N_7258,N_7075,N_7222);
nand U7259 (N_7259,N_7237,N_7041);
or U7260 (N_7260,N_7103,N_7062);
or U7261 (N_7261,N_7236,N_7037);
and U7262 (N_7262,N_7026,N_7066);
nor U7263 (N_7263,N_7039,N_7140);
and U7264 (N_7264,N_7051,N_7215);
nand U7265 (N_7265,N_7144,N_7061);
or U7266 (N_7266,N_7220,N_7107);
xor U7267 (N_7267,N_7212,N_7029);
nor U7268 (N_7268,N_7008,N_7243);
and U7269 (N_7269,N_7170,N_7001);
nor U7270 (N_7270,N_7046,N_7077);
and U7271 (N_7271,N_7213,N_7043);
nand U7272 (N_7272,N_7028,N_7106);
nand U7273 (N_7273,N_7171,N_7015);
or U7274 (N_7274,N_7021,N_7101);
nor U7275 (N_7275,N_7069,N_7120);
nor U7276 (N_7276,N_7132,N_7241);
nor U7277 (N_7277,N_7246,N_7179);
nand U7278 (N_7278,N_7035,N_7059);
or U7279 (N_7279,N_7188,N_7187);
xnor U7280 (N_7280,N_7112,N_7163);
or U7281 (N_7281,N_7100,N_7191);
nor U7282 (N_7282,N_7175,N_7031);
nand U7283 (N_7283,N_7134,N_7159);
and U7284 (N_7284,N_7180,N_7135);
or U7285 (N_7285,N_7048,N_7200);
nand U7286 (N_7286,N_7192,N_7042);
or U7287 (N_7287,N_7169,N_7231);
or U7288 (N_7288,N_7147,N_7121);
nand U7289 (N_7289,N_7010,N_7072);
and U7290 (N_7290,N_7151,N_7184);
and U7291 (N_7291,N_7076,N_7030);
and U7292 (N_7292,N_7011,N_7118);
nand U7293 (N_7293,N_7149,N_7128);
nand U7294 (N_7294,N_7110,N_7206);
xnor U7295 (N_7295,N_7125,N_7181);
or U7296 (N_7296,N_7024,N_7244);
nor U7297 (N_7297,N_7098,N_7119);
nand U7298 (N_7298,N_7033,N_7104);
or U7299 (N_7299,N_7248,N_7005);
xnor U7300 (N_7300,N_7201,N_7064);
nor U7301 (N_7301,N_7233,N_7017);
nor U7302 (N_7302,N_7056,N_7045);
or U7303 (N_7303,N_7019,N_7242);
nand U7304 (N_7304,N_7070,N_7238);
nor U7305 (N_7305,N_7225,N_7114);
nor U7306 (N_7306,N_7190,N_7032);
nand U7307 (N_7307,N_7167,N_7012);
or U7308 (N_7308,N_7089,N_7142);
or U7309 (N_7309,N_7050,N_7060);
and U7310 (N_7310,N_7210,N_7002);
nand U7311 (N_7311,N_7091,N_7000);
or U7312 (N_7312,N_7057,N_7115);
nor U7313 (N_7313,N_7153,N_7189);
and U7314 (N_7314,N_7224,N_7160);
and U7315 (N_7315,N_7124,N_7203);
nand U7316 (N_7316,N_7194,N_7036);
and U7317 (N_7317,N_7018,N_7109);
nand U7318 (N_7318,N_7131,N_7229);
or U7319 (N_7319,N_7207,N_7155);
and U7320 (N_7320,N_7234,N_7195);
and U7321 (N_7321,N_7227,N_7127);
xor U7322 (N_7322,N_7138,N_7247);
or U7323 (N_7323,N_7090,N_7216);
xor U7324 (N_7324,N_7232,N_7053);
and U7325 (N_7325,N_7136,N_7145);
and U7326 (N_7326,N_7117,N_7126);
xor U7327 (N_7327,N_7096,N_7063);
nor U7328 (N_7328,N_7087,N_7223);
xor U7329 (N_7329,N_7094,N_7158);
nand U7330 (N_7330,N_7082,N_7071);
and U7331 (N_7331,N_7113,N_7092);
or U7332 (N_7332,N_7073,N_7172);
nor U7333 (N_7333,N_7186,N_7085);
or U7334 (N_7334,N_7183,N_7157);
nor U7335 (N_7335,N_7235,N_7165);
and U7336 (N_7336,N_7006,N_7249);
nand U7337 (N_7337,N_7221,N_7141);
xor U7338 (N_7338,N_7014,N_7055);
or U7339 (N_7339,N_7130,N_7068);
xor U7340 (N_7340,N_7111,N_7208);
nor U7341 (N_7341,N_7081,N_7025);
or U7342 (N_7342,N_7185,N_7143);
or U7343 (N_7343,N_7197,N_7146);
or U7344 (N_7344,N_7086,N_7004);
nand U7345 (N_7345,N_7080,N_7168);
or U7346 (N_7346,N_7044,N_7016);
nand U7347 (N_7347,N_7102,N_7083);
xnor U7348 (N_7348,N_7047,N_7209);
xnor U7349 (N_7349,N_7245,N_7079);
or U7350 (N_7350,N_7105,N_7218);
or U7351 (N_7351,N_7020,N_7013);
or U7352 (N_7352,N_7162,N_7219);
nor U7353 (N_7353,N_7099,N_7230);
nor U7354 (N_7354,N_7108,N_7152);
and U7355 (N_7355,N_7240,N_7178);
or U7356 (N_7356,N_7196,N_7148);
xnor U7357 (N_7357,N_7007,N_7174);
or U7358 (N_7358,N_7040,N_7164);
or U7359 (N_7359,N_7054,N_7204);
nand U7360 (N_7360,N_7038,N_7226);
xnor U7361 (N_7361,N_7027,N_7173);
or U7362 (N_7362,N_7211,N_7123);
nand U7363 (N_7363,N_7058,N_7122);
nor U7364 (N_7364,N_7182,N_7239);
nor U7365 (N_7365,N_7193,N_7154);
and U7366 (N_7366,N_7176,N_7003);
nand U7367 (N_7367,N_7078,N_7177);
nor U7368 (N_7368,N_7009,N_7166);
nand U7369 (N_7369,N_7205,N_7150);
xor U7370 (N_7370,N_7198,N_7199);
or U7371 (N_7371,N_7133,N_7093);
xnor U7372 (N_7372,N_7137,N_7139);
nor U7373 (N_7373,N_7202,N_7022);
nand U7374 (N_7374,N_7034,N_7067);
nor U7375 (N_7375,N_7083,N_7165);
xor U7376 (N_7376,N_7149,N_7132);
or U7377 (N_7377,N_7036,N_7059);
nor U7378 (N_7378,N_7064,N_7138);
nand U7379 (N_7379,N_7228,N_7153);
or U7380 (N_7380,N_7129,N_7049);
and U7381 (N_7381,N_7116,N_7036);
and U7382 (N_7382,N_7163,N_7008);
nor U7383 (N_7383,N_7109,N_7057);
xnor U7384 (N_7384,N_7046,N_7013);
xor U7385 (N_7385,N_7072,N_7053);
or U7386 (N_7386,N_7102,N_7219);
and U7387 (N_7387,N_7033,N_7235);
xnor U7388 (N_7388,N_7055,N_7215);
xor U7389 (N_7389,N_7012,N_7236);
nor U7390 (N_7390,N_7115,N_7063);
or U7391 (N_7391,N_7142,N_7101);
and U7392 (N_7392,N_7019,N_7076);
or U7393 (N_7393,N_7051,N_7108);
nand U7394 (N_7394,N_7228,N_7208);
xor U7395 (N_7395,N_7183,N_7143);
or U7396 (N_7396,N_7216,N_7019);
or U7397 (N_7397,N_7171,N_7118);
xor U7398 (N_7398,N_7244,N_7173);
or U7399 (N_7399,N_7083,N_7186);
or U7400 (N_7400,N_7032,N_7153);
and U7401 (N_7401,N_7028,N_7185);
and U7402 (N_7402,N_7152,N_7247);
nor U7403 (N_7403,N_7133,N_7237);
nor U7404 (N_7404,N_7106,N_7168);
and U7405 (N_7405,N_7046,N_7219);
and U7406 (N_7406,N_7240,N_7164);
nand U7407 (N_7407,N_7189,N_7052);
nor U7408 (N_7408,N_7179,N_7247);
or U7409 (N_7409,N_7165,N_7181);
nand U7410 (N_7410,N_7247,N_7088);
xnor U7411 (N_7411,N_7146,N_7018);
nand U7412 (N_7412,N_7222,N_7148);
xor U7413 (N_7413,N_7139,N_7016);
and U7414 (N_7414,N_7146,N_7163);
and U7415 (N_7415,N_7244,N_7073);
nand U7416 (N_7416,N_7028,N_7196);
nand U7417 (N_7417,N_7078,N_7095);
xor U7418 (N_7418,N_7119,N_7057);
xnor U7419 (N_7419,N_7134,N_7111);
and U7420 (N_7420,N_7233,N_7203);
xnor U7421 (N_7421,N_7092,N_7184);
or U7422 (N_7422,N_7231,N_7154);
xor U7423 (N_7423,N_7223,N_7079);
or U7424 (N_7424,N_7185,N_7161);
nand U7425 (N_7425,N_7141,N_7005);
xnor U7426 (N_7426,N_7152,N_7102);
nand U7427 (N_7427,N_7081,N_7181);
xnor U7428 (N_7428,N_7233,N_7055);
and U7429 (N_7429,N_7072,N_7159);
nor U7430 (N_7430,N_7228,N_7086);
xor U7431 (N_7431,N_7096,N_7224);
or U7432 (N_7432,N_7058,N_7066);
nand U7433 (N_7433,N_7072,N_7192);
or U7434 (N_7434,N_7176,N_7092);
nor U7435 (N_7435,N_7052,N_7057);
xnor U7436 (N_7436,N_7140,N_7155);
xnor U7437 (N_7437,N_7118,N_7042);
or U7438 (N_7438,N_7146,N_7161);
nand U7439 (N_7439,N_7090,N_7044);
nand U7440 (N_7440,N_7163,N_7089);
nor U7441 (N_7441,N_7163,N_7173);
nor U7442 (N_7442,N_7003,N_7070);
and U7443 (N_7443,N_7087,N_7161);
or U7444 (N_7444,N_7203,N_7101);
xor U7445 (N_7445,N_7024,N_7089);
and U7446 (N_7446,N_7176,N_7134);
nand U7447 (N_7447,N_7153,N_7062);
or U7448 (N_7448,N_7216,N_7054);
xor U7449 (N_7449,N_7153,N_7236);
nor U7450 (N_7450,N_7036,N_7135);
xor U7451 (N_7451,N_7167,N_7067);
xnor U7452 (N_7452,N_7174,N_7013);
nand U7453 (N_7453,N_7181,N_7014);
xor U7454 (N_7454,N_7117,N_7022);
and U7455 (N_7455,N_7176,N_7096);
nand U7456 (N_7456,N_7131,N_7140);
and U7457 (N_7457,N_7244,N_7233);
xor U7458 (N_7458,N_7226,N_7055);
xor U7459 (N_7459,N_7176,N_7230);
and U7460 (N_7460,N_7029,N_7162);
nor U7461 (N_7461,N_7059,N_7029);
or U7462 (N_7462,N_7052,N_7050);
nor U7463 (N_7463,N_7120,N_7062);
xnor U7464 (N_7464,N_7076,N_7135);
and U7465 (N_7465,N_7164,N_7098);
xnor U7466 (N_7466,N_7195,N_7134);
nand U7467 (N_7467,N_7078,N_7000);
xnor U7468 (N_7468,N_7232,N_7044);
or U7469 (N_7469,N_7237,N_7178);
xnor U7470 (N_7470,N_7135,N_7072);
nor U7471 (N_7471,N_7126,N_7205);
and U7472 (N_7472,N_7037,N_7174);
xor U7473 (N_7473,N_7131,N_7024);
nand U7474 (N_7474,N_7248,N_7117);
or U7475 (N_7475,N_7230,N_7018);
xor U7476 (N_7476,N_7089,N_7058);
nand U7477 (N_7477,N_7137,N_7105);
and U7478 (N_7478,N_7193,N_7068);
xor U7479 (N_7479,N_7245,N_7175);
nor U7480 (N_7480,N_7116,N_7230);
nor U7481 (N_7481,N_7103,N_7108);
nand U7482 (N_7482,N_7066,N_7127);
and U7483 (N_7483,N_7221,N_7150);
nor U7484 (N_7484,N_7087,N_7077);
and U7485 (N_7485,N_7230,N_7111);
nand U7486 (N_7486,N_7055,N_7249);
or U7487 (N_7487,N_7019,N_7026);
xor U7488 (N_7488,N_7154,N_7241);
nand U7489 (N_7489,N_7043,N_7231);
or U7490 (N_7490,N_7029,N_7187);
or U7491 (N_7491,N_7016,N_7094);
xnor U7492 (N_7492,N_7243,N_7078);
nor U7493 (N_7493,N_7075,N_7152);
nand U7494 (N_7494,N_7083,N_7088);
and U7495 (N_7495,N_7154,N_7215);
and U7496 (N_7496,N_7019,N_7163);
or U7497 (N_7497,N_7041,N_7133);
or U7498 (N_7498,N_7122,N_7076);
nand U7499 (N_7499,N_7049,N_7086);
xor U7500 (N_7500,N_7312,N_7367);
and U7501 (N_7501,N_7438,N_7404);
nand U7502 (N_7502,N_7325,N_7497);
and U7503 (N_7503,N_7326,N_7432);
xor U7504 (N_7504,N_7381,N_7468);
nand U7505 (N_7505,N_7335,N_7282);
or U7506 (N_7506,N_7406,N_7331);
and U7507 (N_7507,N_7339,N_7320);
and U7508 (N_7508,N_7270,N_7334);
nand U7509 (N_7509,N_7358,N_7460);
nor U7510 (N_7510,N_7480,N_7471);
nor U7511 (N_7511,N_7494,N_7276);
xor U7512 (N_7512,N_7280,N_7436);
and U7513 (N_7513,N_7360,N_7274);
xor U7514 (N_7514,N_7369,N_7351);
nand U7515 (N_7515,N_7267,N_7366);
or U7516 (N_7516,N_7321,N_7344);
and U7517 (N_7517,N_7493,N_7250);
or U7518 (N_7518,N_7411,N_7472);
xor U7519 (N_7519,N_7286,N_7353);
nor U7520 (N_7520,N_7302,N_7253);
nor U7521 (N_7521,N_7435,N_7398);
nand U7522 (N_7522,N_7393,N_7455);
nand U7523 (N_7523,N_7347,N_7299);
xor U7524 (N_7524,N_7462,N_7285);
or U7525 (N_7525,N_7444,N_7394);
and U7526 (N_7526,N_7346,N_7456);
or U7527 (N_7527,N_7425,N_7419);
nand U7528 (N_7528,N_7473,N_7402);
and U7529 (N_7529,N_7341,N_7281);
nor U7530 (N_7530,N_7356,N_7409);
nor U7531 (N_7531,N_7475,N_7386);
nor U7532 (N_7532,N_7291,N_7319);
nor U7533 (N_7533,N_7445,N_7403);
nand U7534 (N_7534,N_7314,N_7466);
and U7535 (N_7535,N_7397,N_7449);
nand U7536 (N_7536,N_7375,N_7478);
or U7537 (N_7537,N_7417,N_7490);
nand U7538 (N_7538,N_7441,N_7450);
and U7539 (N_7539,N_7437,N_7328);
or U7540 (N_7540,N_7284,N_7476);
xor U7541 (N_7541,N_7295,N_7430);
nand U7542 (N_7542,N_7447,N_7296);
xor U7543 (N_7543,N_7443,N_7477);
and U7544 (N_7544,N_7348,N_7370);
nor U7545 (N_7545,N_7499,N_7421);
nand U7546 (N_7546,N_7297,N_7440);
and U7547 (N_7547,N_7498,N_7293);
xor U7548 (N_7548,N_7332,N_7254);
nor U7549 (N_7549,N_7371,N_7448);
nor U7550 (N_7550,N_7469,N_7266);
xnor U7551 (N_7551,N_7413,N_7337);
or U7552 (N_7552,N_7350,N_7272);
xor U7553 (N_7553,N_7365,N_7484);
or U7554 (N_7554,N_7357,N_7277);
or U7555 (N_7555,N_7340,N_7414);
and U7556 (N_7556,N_7491,N_7434);
nand U7557 (N_7557,N_7269,N_7345);
nor U7558 (N_7558,N_7483,N_7261);
nand U7559 (N_7559,N_7488,N_7316);
nor U7560 (N_7560,N_7385,N_7467);
or U7561 (N_7561,N_7265,N_7336);
or U7562 (N_7562,N_7359,N_7292);
xor U7563 (N_7563,N_7308,N_7259);
xor U7564 (N_7564,N_7401,N_7378);
nor U7565 (N_7565,N_7301,N_7306);
or U7566 (N_7566,N_7463,N_7288);
nor U7567 (N_7567,N_7395,N_7283);
nor U7568 (N_7568,N_7322,N_7362);
nor U7569 (N_7569,N_7492,N_7424);
xor U7570 (N_7570,N_7464,N_7279);
nand U7571 (N_7571,N_7256,N_7298);
xnor U7572 (N_7572,N_7383,N_7415);
nor U7573 (N_7573,N_7465,N_7278);
nand U7574 (N_7574,N_7433,N_7426);
and U7575 (N_7575,N_7376,N_7387);
nor U7576 (N_7576,N_7439,N_7373);
and U7577 (N_7577,N_7264,N_7429);
xnor U7578 (N_7578,N_7405,N_7271);
and U7579 (N_7579,N_7252,N_7262);
nor U7580 (N_7580,N_7470,N_7294);
nand U7581 (N_7581,N_7354,N_7489);
or U7582 (N_7582,N_7486,N_7311);
and U7583 (N_7583,N_7391,N_7352);
nand U7584 (N_7584,N_7303,N_7377);
nand U7585 (N_7585,N_7482,N_7310);
nor U7586 (N_7586,N_7452,N_7407);
nor U7587 (N_7587,N_7479,N_7368);
or U7588 (N_7588,N_7307,N_7379);
and U7589 (N_7589,N_7263,N_7446);
and U7590 (N_7590,N_7390,N_7380);
xor U7591 (N_7591,N_7324,N_7290);
nor U7592 (N_7592,N_7338,N_7323);
nand U7593 (N_7593,N_7453,N_7333);
or U7594 (N_7594,N_7487,N_7313);
nor U7595 (N_7595,N_7481,N_7372);
nand U7596 (N_7596,N_7343,N_7374);
nor U7597 (N_7597,N_7318,N_7361);
xor U7598 (N_7598,N_7396,N_7408);
nand U7599 (N_7599,N_7427,N_7289);
xnor U7600 (N_7600,N_7255,N_7416);
or U7601 (N_7601,N_7317,N_7251);
xnor U7602 (N_7602,N_7388,N_7454);
or U7603 (N_7603,N_7461,N_7420);
nor U7604 (N_7604,N_7458,N_7275);
xor U7605 (N_7605,N_7327,N_7412);
nor U7606 (N_7606,N_7329,N_7442);
or U7607 (N_7607,N_7257,N_7418);
or U7608 (N_7608,N_7459,N_7400);
or U7609 (N_7609,N_7423,N_7384);
xor U7610 (N_7610,N_7315,N_7273);
or U7611 (N_7611,N_7305,N_7268);
nand U7612 (N_7612,N_7304,N_7363);
xnor U7613 (N_7613,N_7287,N_7485);
and U7614 (N_7614,N_7474,N_7399);
nand U7615 (N_7615,N_7349,N_7260);
nand U7616 (N_7616,N_7258,N_7495);
xor U7617 (N_7617,N_7364,N_7389);
nor U7618 (N_7618,N_7300,N_7428);
nor U7619 (N_7619,N_7330,N_7309);
or U7620 (N_7620,N_7342,N_7410);
nand U7621 (N_7621,N_7422,N_7392);
xor U7622 (N_7622,N_7355,N_7431);
and U7623 (N_7623,N_7457,N_7496);
nand U7624 (N_7624,N_7451,N_7382);
nor U7625 (N_7625,N_7463,N_7364);
nor U7626 (N_7626,N_7295,N_7347);
xor U7627 (N_7627,N_7298,N_7414);
xnor U7628 (N_7628,N_7388,N_7277);
xnor U7629 (N_7629,N_7444,N_7339);
nand U7630 (N_7630,N_7468,N_7408);
xnor U7631 (N_7631,N_7324,N_7478);
and U7632 (N_7632,N_7394,N_7342);
xnor U7633 (N_7633,N_7264,N_7422);
xnor U7634 (N_7634,N_7360,N_7379);
nand U7635 (N_7635,N_7302,N_7266);
nor U7636 (N_7636,N_7310,N_7336);
nor U7637 (N_7637,N_7298,N_7405);
nor U7638 (N_7638,N_7351,N_7466);
xnor U7639 (N_7639,N_7365,N_7260);
nand U7640 (N_7640,N_7300,N_7435);
or U7641 (N_7641,N_7394,N_7354);
nand U7642 (N_7642,N_7280,N_7400);
xor U7643 (N_7643,N_7271,N_7372);
nor U7644 (N_7644,N_7344,N_7350);
and U7645 (N_7645,N_7377,N_7451);
or U7646 (N_7646,N_7335,N_7263);
and U7647 (N_7647,N_7459,N_7412);
and U7648 (N_7648,N_7487,N_7457);
nor U7649 (N_7649,N_7294,N_7406);
xnor U7650 (N_7650,N_7359,N_7385);
nor U7651 (N_7651,N_7310,N_7403);
and U7652 (N_7652,N_7371,N_7437);
xnor U7653 (N_7653,N_7387,N_7373);
or U7654 (N_7654,N_7274,N_7384);
nand U7655 (N_7655,N_7356,N_7302);
nand U7656 (N_7656,N_7301,N_7444);
nand U7657 (N_7657,N_7368,N_7354);
and U7658 (N_7658,N_7261,N_7428);
or U7659 (N_7659,N_7302,N_7284);
and U7660 (N_7660,N_7459,N_7448);
xor U7661 (N_7661,N_7264,N_7404);
xor U7662 (N_7662,N_7320,N_7393);
xnor U7663 (N_7663,N_7392,N_7385);
nor U7664 (N_7664,N_7474,N_7492);
nand U7665 (N_7665,N_7283,N_7303);
xor U7666 (N_7666,N_7283,N_7309);
or U7667 (N_7667,N_7379,N_7356);
and U7668 (N_7668,N_7485,N_7354);
xnor U7669 (N_7669,N_7308,N_7368);
or U7670 (N_7670,N_7359,N_7423);
and U7671 (N_7671,N_7471,N_7479);
and U7672 (N_7672,N_7372,N_7362);
nand U7673 (N_7673,N_7403,N_7414);
nand U7674 (N_7674,N_7330,N_7382);
nand U7675 (N_7675,N_7416,N_7331);
and U7676 (N_7676,N_7264,N_7316);
or U7677 (N_7677,N_7252,N_7487);
xnor U7678 (N_7678,N_7436,N_7415);
nand U7679 (N_7679,N_7391,N_7423);
nor U7680 (N_7680,N_7476,N_7384);
and U7681 (N_7681,N_7371,N_7403);
and U7682 (N_7682,N_7355,N_7262);
nand U7683 (N_7683,N_7328,N_7349);
nand U7684 (N_7684,N_7353,N_7345);
xor U7685 (N_7685,N_7287,N_7451);
xnor U7686 (N_7686,N_7465,N_7439);
nor U7687 (N_7687,N_7419,N_7409);
xnor U7688 (N_7688,N_7289,N_7426);
nand U7689 (N_7689,N_7454,N_7427);
xnor U7690 (N_7690,N_7290,N_7299);
and U7691 (N_7691,N_7268,N_7390);
and U7692 (N_7692,N_7410,N_7380);
nor U7693 (N_7693,N_7496,N_7322);
or U7694 (N_7694,N_7286,N_7348);
and U7695 (N_7695,N_7255,N_7265);
xnor U7696 (N_7696,N_7270,N_7273);
nand U7697 (N_7697,N_7485,N_7442);
xor U7698 (N_7698,N_7285,N_7436);
and U7699 (N_7699,N_7490,N_7472);
xor U7700 (N_7700,N_7362,N_7297);
or U7701 (N_7701,N_7302,N_7465);
nor U7702 (N_7702,N_7341,N_7306);
nand U7703 (N_7703,N_7486,N_7428);
or U7704 (N_7704,N_7417,N_7455);
nor U7705 (N_7705,N_7375,N_7497);
xor U7706 (N_7706,N_7403,N_7341);
nand U7707 (N_7707,N_7395,N_7280);
nor U7708 (N_7708,N_7400,N_7255);
nor U7709 (N_7709,N_7486,N_7341);
nand U7710 (N_7710,N_7493,N_7406);
nand U7711 (N_7711,N_7363,N_7264);
and U7712 (N_7712,N_7305,N_7425);
and U7713 (N_7713,N_7271,N_7380);
or U7714 (N_7714,N_7265,N_7424);
nand U7715 (N_7715,N_7398,N_7358);
and U7716 (N_7716,N_7336,N_7391);
nor U7717 (N_7717,N_7332,N_7464);
xnor U7718 (N_7718,N_7458,N_7258);
or U7719 (N_7719,N_7457,N_7357);
or U7720 (N_7720,N_7282,N_7340);
and U7721 (N_7721,N_7451,N_7374);
nand U7722 (N_7722,N_7330,N_7274);
xor U7723 (N_7723,N_7397,N_7369);
nor U7724 (N_7724,N_7459,N_7457);
nand U7725 (N_7725,N_7259,N_7362);
nor U7726 (N_7726,N_7428,N_7367);
nand U7727 (N_7727,N_7290,N_7291);
nand U7728 (N_7728,N_7345,N_7391);
and U7729 (N_7729,N_7305,N_7366);
nor U7730 (N_7730,N_7499,N_7300);
or U7731 (N_7731,N_7267,N_7336);
nand U7732 (N_7732,N_7351,N_7321);
nor U7733 (N_7733,N_7432,N_7473);
and U7734 (N_7734,N_7326,N_7336);
nand U7735 (N_7735,N_7373,N_7413);
xnor U7736 (N_7736,N_7282,N_7291);
or U7737 (N_7737,N_7450,N_7315);
nor U7738 (N_7738,N_7426,N_7376);
nor U7739 (N_7739,N_7444,N_7285);
nand U7740 (N_7740,N_7459,N_7450);
or U7741 (N_7741,N_7296,N_7472);
and U7742 (N_7742,N_7454,N_7438);
nor U7743 (N_7743,N_7265,N_7421);
nor U7744 (N_7744,N_7403,N_7400);
or U7745 (N_7745,N_7373,N_7384);
or U7746 (N_7746,N_7272,N_7263);
xor U7747 (N_7747,N_7292,N_7395);
and U7748 (N_7748,N_7463,N_7358);
nor U7749 (N_7749,N_7291,N_7408);
xnor U7750 (N_7750,N_7520,N_7619);
xor U7751 (N_7751,N_7686,N_7640);
or U7752 (N_7752,N_7638,N_7610);
nand U7753 (N_7753,N_7591,N_7564);
or U7754 (N_7754,N_7708,N_7733);
nand U7755 (N_7755,N_7651,N_7681);
and U7756 (N_7756,N_7687,N_7658);
nand U7757 (N_7757,N_7558,N_7728);
nand U7758 (N_7758,N_7677,N_7525);
xnor U7759 (N_7759,N_7675,N_7614);
nor U7760 (N_7760,N_7663,N_7706);
or U7761 (N_7761,N_7628,N_7569);
nor U7762 (N_7762,N_7669,N_7590);
and U7763 (N_7763,N_7512,N_7670);
or U7764 (N_7764,N_7534,N_7615);
xor U7765 (N_7765,N_7611,N_7514);
nand U7766 (N_7766,N_7637,N_7500);
and U7767 (N_7767,N_7504,N_7541);
nor U7768 (N_7768,N_7549,N_7722);
or U7769 (N_7769,N_7662,N_7603);
xor U7770 (N_7770,N_7597,N_7616);
xor U7771 (N_7771,N_7550,N_7711);
xor U7772 (N_7772,N_7606,N_7593);
and U7773 (N_7773,N_7680,N_7529);
or U7774 (N_7774,N_7579,N_7599);
nor U7775 (N_7775,N_7556,N_7505);
nor U7776 (N_7776,N_7609,N_7661);
or U7777 (N_7777,N_7655,N_7513);
nand U7778 (N_7778,N_7607,N_7538);
nand U7779 (N_7779,N_7527,N_7709);
nand U7780 (N_7780,N_7641,N_7678);
nand U7781 (N_7781,N_7725,N_7546);
xor U7782 (N_7782,N_7632,N_7705);
or U7783 (N_7783,N_7642,N_7713);
nand U7784 (N_7784,N_7712,N_7526);
and U7785 (N_7785,N_7622,N_7608);
or U7786 (N_7786,N_7543,N_7693);
and U7787 (N_7787,N_7745,N_7629);
nand U7788 (N_7788,N_7671,N_7739);
and U7789 (N_7789,N_7717,N_7578);
or U7790 (N_7790,N_7691,N_7519);
xor U7791 (N_7791,N_7692,N_7581);
xor U7792 (N_7792,N_7699,N_7555);
xor U7793 (N_7793,N_7589,N_7730);
nand U7794 (N_7794,N_7639,N_7666);
or U7795 (N_7795,N_7624,N_7653);
nor U7796 (N_7796,N_7649,N_7650);
xnor U7797 (N_7797,N_7732,N_7511);
xnor U7798 (N_7798,N_7565,N_7571);
nand U7799 (N_7799,N_7716,N_7747);
nor U7800 (N_7800,N_7690,N_7531);
nand U7801 (N_7801,N_7647,N_7635);
xnor U7802 (N_7802,N_7592,N_7723);
and U7803 (N_7803,N_7617,N_7654);
and U7804 (N_7804,N_7503,N_7673);
and U7805 (N_7805,N_7659,N_7553);
or U7806 (N_7806,N_7676,N_7714);
and U7807 (N_7807,N_7535,N_7645);
or U7808 (N_7808,N_7586,N_7742);
xor U7809 (N_7809,N_7643,N_7539);
and U7810 (N_7810,N_7510,N_7679);
nor U7811 (N_7811,N_7623,N_7580);
and U7812 (N_7812,N_7559,N_7567);
xor U7813 (N_7813,N_7502,N_7695);
xor U7814 (N_7814,N_7696,N_7583);
and U7815 (N_7815,N_7554,N_7704);
or U7816 (N_7816,N_7524,N_7521);
and U7817 (N_7817,N_7729,N_7741);
or U7818 (N_7818,N_7573,N_7618);
nand U7819 (N_7819,N_7584,N_7574);
or U7820 (N_7820,N_7646,N_7537);
or U7821 (N_7821,N_7726,N_7575);
and U7822 (N_7822,N_7707,N_7598);
xnor U7823 (N_7823,N_7698,N_7701);
and U7824 (N_7824,N_7507,N_7562);
nor U7825 (N_7825,N_7667,N_7631);
and U7826 (N_7826,N_7621,N_7737);
and U7827 (N_7827,N_7672,N_7545);
xnor U7828 (N_7828,N_7721,N_7548);
or U7829 (N_7829,N_7509,N_7633);
and U7830 (N_7830,N_7625,N_7738);
or U7831 (N_7831,N_7748,N_7736);
and U7832 (N_7832,N_7517,N_7508);
nand U7833 (N_7833,N_7594,N_7665);
or U7834 (N_7834,N_7577,N_7664);
nand U7835 (N_7835,N_7660,N_7694);
nor U7836 (N_7836,N_7604,N_7501);
or U7837 (N_7837,N_7601,N_7700);
nand U7838 (N_7838,N_7697,N_7746);
nand U7839 (N_7839,N_7600,N_7533);
and U7840 (N_7840,N_7561,N_7719);
xnor U7841 (N_7841,N_7582,N_7612);
or U7842 (N_7842,N_7689,N_7718);
and U7843 (N_7843,N_7551,N_7528);
and U7844 (N_7844,N_7735,N_7656);
xnor U7845 (N_7845,N_7540,N_7731);
nor U7846 (N_7846,N_7715,N_7668);
nand U7847 (N_7847,N_7605,N_7557);
or U7848 (N_7848,N_7749,N_7702);
nor U7849 (N_7849,N_7518,N_7596);
nand U7850 (N_7850,N_7522,N_7710);
xor U7851 (N_7851,N_7572,N_7724);
or U7852 (N_7852,N_7570,N_7542);
xnor U7853 (N_7853,N_7740,N_7506);
and U7854 (N_7854,N_7585,N_7627);
or U7855 (N_7855,N_7516,N_7587);
nand U7856 (N_7856,N_7682,N_7634);
nand U7857 (N_7857,N_7552,N_7734);
nor U7858 (N_7858,N_7743,N_7620);
and U7859 (N_7859,N_7720,N_7684);
or U7860 (N_7860,N_7588,N_7595);
and U7861 (N_7861,N_7568,N_7536);
and U7862 (N_7862,N_7532,N_7544);
xnor U7863 (N_7863,N_7602,N_7630);
nor U7864 (N_7864,N_7547,N_7576);
nand U7865 (N_7865,N_7560,N_7688);
xor U7866 (N_7866,N_7523,N_7563);
or U7867 (N_7867,N_7657,N_7613);
nor U7868 (N_7868,N_7644,N_7674);
nor U7869 (N_7869,N_7636,N_7652);
and U7870 (N_7870,N_7566,N_7703);
xnor U7871 (N_7871,N_7727,N_7744);
or U7872 (N_7872,N_7685,N_7683);
xnor U7873 (N_7873,N_7648,N_7626);
and U7874 (N_7874,N_7515,N_7530);
or U7875 (N_7875,N_7568,N_7683);
nand U7876 (N_7876,N_7552,N_7706);
xor U7877 (N_7877,N_7746,N_7508);
and U7878 (N_7878,N_7672,N_7504);
or U7879 (N_7879,N_7744,N_7546);
or U7880 (N_7880,N_7731,N_7505);
and U7881 (N_7881,N_7702,N_7529);
or U7882 (N_7882,N_7551,N_7589);
nand U7883 (N_7883,N_7711,N_7696);
and U7884 (N_7884,N_7697,N_7549);
nand U7885 (N_7885,N_7504,N_7580);
and U7886 (N_7886,N_7584,N_7598);
nand U7887 (N_7887,N_7639,N_7579);
and U7888 (N_7888,N_7702,N_7540);
and U7889 (N_7889,N_7512,N_7618);
nand U7890 (N_7890,N_7519,N_7603);
or U7891 (N_7891,N_7517,N_7706);
or U7892 (N_7892,N_7589,N_7631);
or U7893 (N_7893,N_7705,N_7511);
and U7894 (N_7894,N_7731,N_7631);
xnor U7895 (N_7895,N_7637,N_7715);
nand U7896 (N_7896,N_7640,N_7706);
and U7897 (N_7897,N_7609,N_7590);
and U7898 (N_7898,N_7555,N_7660);
nor U7899 (N_7899,N_7636,N_7579);
xnor U7900 (N_7900,N_7726,N_7581);
and U7901 (N_7901,N_7596,N_7504);
or U7902 (N_7902,N_7573,N_7565);
and U7903 (N_7903,N_7588,N_7513);
nand U7904 (N_7904,N_7614,N_7547);
nor U7905 (N_7905,N_7576,N_7683);
and U7906 (N_7906,N_7519,N_7686);
and U7907 (N_7907,N_7570,N_7708);
or U7908 (N_7908,N_7712,N_7595);
nor U7909 (N_7909,N_7551,N_7521);
and U7910 (N_7910,N_7608,N_7713);
nand U7911 (N_7911,N_7566,N_7616);
nand U7912 (N_7912,N_7743,N_7613);
or U7913 (N_7913,N_7678,N_7642);
or U7914 (N_7914,N_7516,N_7619);
and U7915 (N_7915,N_7737,N_7612);
xor U7916 (N_7916,N_7732,N_7513);
nor U7917 (N_7917,N_7569,N_7600);
and U7918 (N_7918,N_7642,N_7710);
and U7919 (N_7919,N_7710,N_7674);
and U7920 (N_7920,N_7576,N_7688);
xnor U7921 (N_7921,N_7581,N_7719);
nor U7922 (N_7922,N_7548,N_7684);
or U7923 (N_7923,N_7614,N_7590);
nor U7924 (N_7924,N_7577,N_7529);
xnor U7925 (N_7925,N_7559,N_7539);
nor U7926 (N_7926,N_7716,N_7644);
xor U7927 (N_7927,N_7577,N_7573);
or U7928 (N_7928,N_7539,N_7538);
or U7929 (N_7929,N_7613,N_7557);
nor U7930 (N_7930,N_7628,N_7620);
nand U7931 (N_7931,N_7692,N_7539);
nand U7932 (N_7932,N_7500,N_7667);
or U7933 (N_7933,N_7715,N_7517);
nor U7934 (N_7934,N_7682,N_7674);
nor U7935 (N_7935,N_7656,N_7746);
and U7936 (N_7936,N_7593,N_7576);
and U7937 (N_7937,N_7564,N_7733);
nand U7938 (N_7938,N_7501,N_7571);
or U7939 (N_7939,N_7618,N_7639);
and U7940 (N_7940,N_7725,N_7624);
and U7941 (N_7941,N_7510,N_7736);
or U7942 (N_7942,N_7535,N_7671);
xor U7943 (N_7943,N_7708,N_7690);
nor U7944 (N_7944,N_7554,N_7594);
or U7945 (N_7945,N_7533,N_7635);
nor U7946 (N_7946,N_7575,N_7723);
nand U7947 (N_7947,N_7742,N_7587);
and U7948 (N_7948,N_7584,N_7592);
nand U7949 (N_7949,N_7550,N_7596);
xnor U7950 (N_7950,N_7671,N_7609);
nor U7951 (N_7951,N_7713,N_7600);
xor U7952 (N_7952,N_7715,N_7706);
xnor U7953 (N_7953,N_7596,N_7744);
or U7954 (N_7954,N_7732,N_7706);
nor U7955 (N_7955,N_7698,N_7546);
nor U7956 (N_7956,N_7647,N_7633);
or U7957 (N_7957,N_7623,N_7582);
nand U7958 (N_7958,N_7584,N_7722);
nand U7959 (N_7959,N_7683,N_7642);
and U7960 (N_7960,N_7635,N_7662);
and U7961 (N_7961,N_7650,N_7652);
xor U7962 (N_7962,N_7509,N_7710);
xor U7963 (N_7963,N_7606,N_7513);
or U7964 (N_7964,N_7516,N_7660);
and U7965 (N_7965,N_7507,N_7529);
xnor U7966 (N_7966,N_7556,N_7609);
or U7967 (N_7967,N_7746,N_7559);
xnor U7968 (N_7968,N_7683,N_7646);
and U7969 (N_7969,N_7617,N_7622);
nor U7970 (N_7970,N_7562,N_7732);
or U7971 (N_7971,N_7698,N_7729);
and U7972 (N_7972,N_7607,N_7609);
xor U7973 (N_7973,N_7510,N_7553);
xnor U7974 (N_7974,N_7589,N_7702);
or U7975 (N_7975,N_7731,N_7702);
nor U7976 (N_7976,N_7541,N_7729);
or U7977 (N_7977,N_7558,N_7706);
nand U7978 (N_7978,N_7660,N_7717);
nor U7979 (N_7979,N_7586,N_7665);
or U7980 (N_7980,N_7530,N_7679);
nand U7981 (N_7981,N_7562,N_7683);
and U7982 (N_7982,N_7727,N_7627);
and U7983 (N_7983,N_7518,N_7601);
and U7984 (N_7984,N_7723,N_7726);
or U7985 (N_7985,N_7588,N_7542);
xnor U7986 (N_7986,N_7616,N_7526);
or U7987 (N_7987,N_7720,N_7692);
nor U7988 (N_7988,N_7558,N_7688);
and U7989 (N_7989,N_7643,N_7682);
or U7990 (N_7990,N_7524,N_7543);
and U7991 (N_7991,N_7506,N_7528);
xnor U7992 (N_7992,N_7740,N_7585);
nor U7993 (N_7993,N_7652,N_7729);
xnor U7994 (N_7994,N_7602,N_7747);
xor U7995 (N_7995,N_7510,N_7668);
xnor U7996 (N_7996,N_7545,N_7511);
nand U7997 (N_7997,N_7749,N_7509);
and U7998 (N_7998,N_7604,N_7739);
nor U7999 (N_7999,N_7670,N_7502);
nor U8000 (N_8000,N_7937,N_7777);
xnor U8001 (N_8001,N_7866,N_7904);
and U8002 (N_8002,N_7966,N_7855);
nand U8003 (N_8003,N_7827,N_7938);
xnor U8004 (N_8004,N_7876,N_7895);
nand U8005 (N_8005,N_7980,N_7981);
xnor U8006 (N_8006,N_7897,N_7756);
xnor U8007 (N_8007,N_7965,N_7944);
or U8008 (N_8008,N_7752,N_7901);
xor U8009 (N_8009,N_7975,N_7973);
nor U8010 (N_8010,N_7917,N_7772);
nand U8011 (N_8011,N_7935,N_7916);
or U8012 (N_8012,N_7905,N_7954);
and U8013 (N_8013,N_7779,N_7919);
or U8014 (N_8014,N_7896,N_7939);
and U8015 (N_8015,N_7891,N_7840);
and U8016 (N_8016,N_7970,N_7979);
xor U8017 (N_8017,N_7789,N_7851);
and U8018 (N_8018,N_7774,N_7910);
or U8019 (N_8019,N_7996,N_7961);
xor U8020 (N_8020,N_7800,N_7757);
nand U8021 (N_8021,N_7962,N_7931);
and U8022 (N_8022,N_7924,N_7869);
xor U8023 (N_8023,N_7786,N_7862);
nor U8024 (N_8024,N_7834,N_7788);
or U8025 (N_8025,N_7761,N_7948);
nor U8026 (N_8026,N_7835,N_7999);
nor U8027 (N_8027,N_7803,N_7923);
and U8028 (N_8028,N_7854,N_7775);
nor U8029 (N_8029,N_7816,N_7982);
or U8030 (N_8030,N_7860,N_7831);
and U8031 (N_8031,N_7837,N_7994);
and U8032 (N_8032,N_7806,N_7941);
nand U8033 (N_8033,N_7934,N_7972);
nor U8034 (N_8034,N_7952,N_7881);
and U8035 (N_8035,N_7811,N_7852);
xor U8036 (N_8036,N_7823,N_7785);
and U8037 (N_8037,N_7783,N_7971);
nor U8038 (N_8038,N_7805,N_7960);
nor U8039 (N_8039,N_7977,N_7873);
nand U8040 (N_8040,N_7802,N_7947);
and U8041 (N_8041,N_7875,N_7986);
nand U8042 (N_8042,N_7893,N_7997);
and U8043 (N_8043,N_7976,N_7892);
nand U8044 (N_8044,N_7959,N_7932);
nor U8045 (N_8045,N_7769,N_7794);
nor U8046 (N_8046,N_7763,N_7781);
nor U8047 (N_8047,N_7818,N_7838);
and U8048 (N_8048,N_7985,N_7922);
nor U8049 (N_8049,N_7753,N_7762);
nor U8050 (N_8050,N_7795,N_7861);
or U8051 (N_8051,N_7841,N_7877);
xnor U8052 (N_8052,N_7859,N_7846);
and U8053 (N_8053,N_7815,N_7819);
nor U8054 (N_8054,N_7771,N_7953);
xnor U8055 (N_8055,N_7902,N_7908);
or U8056 (N_8056,N_7950,N_7874);
or U8057 (N_8057,N_7940,N_7909);
xor U8058 (N_8058,N_7974,N_7995);
nor U8059 (N_8059,N_7864,N_7886);
nand U8060 (N_8060,N_7914,N_7998);
xor U8061 (N_8061,N_7764,N_7957);
xor U8062 (N_8062,N_7810,N_7949);
or U8063 (N_8063,N_7817,N_7857);
nor U8064 (N_8064,N_7820,N_7865);
nand U8065 (N_8065,N_7770,N_7798);
nor U8066 (N_8066,N_7899,N_7898);
or U8067 (N_8067,N_7946,N_7766);
nand U8068 (N_8068,N_7907,N_7787);
nor U8069 (N_8069,N_7936,N_7767);
xor U8070 (N_8070,N_7987,N_7822);
and U8071 (N_8071,N_7990,N_7821);
nor U8072 (N_8072,N_7760,N_7768);
nand U8073 (N_8073,N_7993,N_7913);
and U8074 (N_8074,N_7808,N_7958);
or U8075 (N_8075,N_7793,N_7903);
xor U8076 (N_8076,N_7967,N_7751);
and U8077 (N_8077,N_7983,N_7928);
and U8078 (N_8078,N_7890,N_7836);
xnor U8079 (N_8079,N_7858,N_7833);
xor U8080 (N_8080,N_7863,N_7792);
nor U8081 (N_8081,N_7889,N_7778);
nand U8082 (N_8082,N_7799,N_7839);
or U8083 (N_8083,N_7844,N_7918);
nor U8084 (N_8084,N_7871,N_7872);
or U8085 (N_8085,N_7921,N_7867);
nor U8086 (N_8086,N_7945,N_7870);
or U8087 (N_8087,N_7942,N_7930);
xnor U8088 (N_8088,N_7926,N_7978);
or U8089 (N_8089,N_7885,N_7813);
or U8090 (N_8090,N_7964,N_7887);
or U8091 (N_8091,N_7991,N_7847);
and U8092 (N_8092,N_7984,N_7754);
or U8093 (N_8093,N_7814,N_7782);
nand U8094 (N_8094,N_7920,N_7879);
and U8095 (N_8095,N_7929,N_7888);
nor U8096 (N_8096,N_7758,N_7915);
nand U8097 (N_8097,N_7848,N_7825);
or U8098 (N_8098,N_7828,N_7824);
nor U8099 (N_8099,N_7988,N_7884);
or U8100 (N_8100,N_7992,N_7925);
and U8101 (N_8101,N_7784,N_7943);
xnor U8102 (N_8102,N_7812,N_7791);
nand U8103 (N_8103,N_7850,N_7765);
nor U8104 (N_8104,N_7951,N_7956);
and U8105 (N_8105,N_7927,N_7829);
or U8106 (N_8106,N_7900,N_7790);
and U8107 (N_8107,N_7968,N_7856);
xnor U8108 (N_8108,N_7969,N_7989);
xor U8109 (N_8109,N_7809,N_7801);
or U8110 (N_8110,N_7882,N_7826);
xor U8111 (N_8111,N_7878,N_7759);
nand U8112 (N_8112,N_7755,N_7880);
xnor U8113 (N_8113,N_7807,N_7830);
nor U8114 (N_8114,N_7906,N_7804);
and U8115 (N_8115,N_7845,N_7796);
nor U8116 (N_8116,N_7894,N_7912);
xnor U8117 (N_8117,N_7750,N_7797);
xnor U8118 (N_8118,N_7776,N_7955);
and U8119 (N_8119,N_7843,N_7853);
nand U8120 (N_8120,N_7868,N_7773);
xor U8121 (N_8121,N_7849,N_7780);
xor U8122 (N_8122,N_7933,N_7963);
or U8123 (N_8123,N_7911,N_7832);
and U8124 (N_8124,N_7842,N_7883);
and U8125 (N_8125,N_7774,N_7851);
xnor U8126 (N_8126,N_7870,N_7940);
xor U8127 (N_8127,N_7894,N_7941);
nor U8128 (N_8128,N_7823,N_7864);
nor U8129 (N_8129,N_7847,N_7783);
or U8130 (N_8130,N_7830,N_7971);
or U8131 (N_8131,N_7969,N_7785);
and U8132 (N_8132,N_7840,N_7824);
or U8133 (N_8133,N_7988,N_7970);
or U8134 (N_8134,N_7854,N_7890);
or U8135 (N_8135,N_7807,N_7845);
or U8136 (N_8136,N_7883,N_7862);
xnor U8137 (N_8137,N_7816,N_7837);
xor U8138 (N_8138,N_7983,N_7917);
nor U8139 (N_8139,N_7990,N_7861);
and U8140 (N_8140,N_7802,N_7766);
and U8141 (N_8141,N_7847,N_7828);
nand U8142 (N_8142,N_7840,N_7864);
and U8143 (N_8143,N_7832,N_7940);
nand U8144 (N_8144,N_7835,N_7890);
nor U8145 (N_8145,N_7971,N_7969);
nor U8146 (N_8146,N_7841,N_7751);
and U8147 (N_8147,N_7805,N_7969);
nor U8148 (N_8148,N_7983,N_7956);
xor U8149 (N_8149,N_7981,N_7984);
or U8150 (N_8150,N_7978,N_7925);
and U8151 (N_8151,N_7768,N_7847);
and U8152 (N_8152,N_7955,N_7849);
and U8153 (N_8153,N_7833,N_7939);
and U8154 (N_8154,N_7945,N_7818);
nand U8155 (N_8155,N_7890,N_7773);
nand U8156 (N_8156,N_7781,N_7959);
nor U8157 (N_8157,N_7879,N_7924);
xor U8158 (N_8158,N_7771,N_7966);
or U8159 (N_8159,N_7757,N_7906);
and U8160 (N_8160,N_7992,N_7970);
or U8161 (N_8161,N_7998,N_7823);
and U8162 (N_8162,N_7860,N_7803);
xor U8163 (N_8163,N_7961,N_7926);
and U8164 (N_8164,N_7830,N_7774);
nor U8165 (N_8165,N_7824,N_7783);
nand U8166 (N_8166,N_7841,N_7903);
xnor U8167 (N_8167,N_7960,N_7933);
and U8168 (N_8168,N_7750,N_7767);
nand U8169 (N_8169,N_7980,N_7915);
nor U8170 (N_8170,N_7915,N_7981);
xor U8171 (N_8171,N_7975,N_7823);
and U8172 (N_8172,N_7874,N_7759);
nor U8173 (N_8173,N_7938,N_7921);
nand U8174 (N_8174,N_7798,N_7953);
or U8175 (N_8175,N_7829,N_7919);
or U8176 (N_8176,N_7972,N_7887);
nor U8177 (N_8177,N_7932,N_7792);
xor U8178 (N_8178,N_7959,N_7848);
or U8179 (N_8179,N_7893,N_7870);
and U8180 (N_8180,N_7854,N_7900);
nand U8181 (N_8181,N_7769,N_7890);
nand U8182 (N_8182,N_7912,N_7908);
nand U8183 (N_8183,N_7859,N_7977);
nand U8184 (N_8184,N_7837,N_7860);
nand U8185 (N_8185,N_7773,N_7936);
nor U8186 (N_8186,N_7958,N_7966);
nand U8187 (N_8187,N_7750,N_7813);
nand U8188 (N_8188,N_7890,N_7761);
xnor U8189 (N_8189,N_7870,N_7753);
or U8190 (N_8190,N_7877,N_7949);
nand U8191 (N_8191,N_7844,N_7959);
xor U8192 (N_8192,N_7939,N_7953);
nand U8193 (N_8193,N_7791,N_7763);
or U8194 (N_8194,N_7810,N_7913);
and U8195 (N_8195,N_7911,N_7990);
nor U8196 (N_8196,N_7984,N_7868);
nor U8197 (N_8197,N_7928,N_7816);
xnor U8198 (N_8198,N_7814,N_7788);
nand U8199 (N_8199,N_7915,N_7889);
or U8200 (N_8200,N_7882,N_7807);
nand U8201 (N_8201,N_7849,N_7882);
nand U8202 (N_8202,N_7969,N_7772);
xor U8203 (N_8203,N_7752,N_7917);
nand U8204 (N_8204,N_7754,N_7916);
nor U8205 (N_8205,N_7974,N_7805);
nand U8206 (N_8206,N_7910,N_7883);
nor U8207 (N_8207,N_7764,N_7917);
or U8208 (N_8208,N_7786,N_7787);
nor U8209 (N_8209,N_7916,N_7984);
or U8210 (N_8210,N_7906,N_7963);
xor U8211 (N_8211,N_7986,N_7930);
and U8212 (N_8212,N_7891,N_7924);
nor U8213 (N_8213,N_7866,N_7919);
nor U8214 (N_8214,N_7939,N_7956);
xnor U8215 (N_8215,N_7863,N_7946);
nor U8216 (N_8216,N_7755,N_7879);
nor U8217 (N_8217,N_7931,N_7961);
or U8218 (N_8218,N_7967,N_7787);
nand U8219 (N_8219,N_7802,N_7792);
nor U8220 (N_8220,N_7986,N_7983);
xor U8221 (N_8221,N_7842,N_7984);
xnor U8222 (N_8222,N_7753,N_7820);
or U8223 (N_8223,N_7832,N_7824);
and U8224 (N_8224,N_7995,N_7950);
nand U8225 (N_8225,N_7975,N_7852);
xor U8226 (N_8226,N_7894,N_7995);
nor U8227 (N_8227,N_7837,N_7829);
and U8228 (N_8228,N_7922,N_7996);
or U8229 (N_8229,N_7952,N_7977);
nor U8230 (N_8230,N_7965,N_7789);
xnor U8231 (N_8231,N_7978,N_7901);
or U8232 (N_8232,N_7842,N_7809);
and U8233 (N_8233,N_7756,N_7956);
and U8234 (N_8234,N_7920,N_7803);
xnor U8235 (N_8235,N_7903,N_7808);
or U8236 (N_8236,N_7879,N_7875);
or U8237 (N_8237,N_7926,N_7893);
nor U8238 (N_8238,N_7782,N_7972);
nand U8239 (N_8239,N_7967,N_7852);
nand U8240 (N_8240,N_7769,N_7977);
nor U8241 (N_8241,N_7982,N_7839);
and U8242 (N_8242,N_7972,N_7935);
and U8243 (N_8243,N_7805,N_7881);
and U8244 (N_8244,N_7912,N_7755);
nor U8245 (N_8245,N_7863,N_7794);
nand U8246 (N_8246,N_7935,N_7928);
or U8247 (N_8247,N_7999,N_7940);
or U8248 (N_8248,N_7963,N_7878);
or U8249 (N_8249,N_7860,N_7885);
nand U8250 (N_8250,N_8185,N_8062);
xor U8251 (N_8251,N_8091,N_8180);
xnor U8252 (N_8252,N_8023,N_8226);
or U8253 (N_8253,N_8043,N_8008);
nand U8254 (N_8254,N_8233,N_8065);
and U8255 (N_8255,N_8105,N_8031);
nand U8256 (N_8256,N_8005,N_8142);
and U8257 (N_8257,N_8203,N_8088);
nor U8258 (N_8258,N_8015,N_8093);
or U8259 (N_8259,N_8209,N_8044);
nand U8260 (N_8260,N_8011,N_8077);
or U8261 (N_8261,N_8136,N_8162);
nand U8262 (N_8262,N_8187,N_8198);
xor U8263 (N_8263,N_8217,N_8184);
nor U8264 (N_8264,N_8117,N_8205);
and U8265 (N_8265,N_8033,N_8219);
nor U8266 (N_8266,N_8041,N_8210);
and U8267 (N_8267,N_8102,N_8202);
or U8268 (N_8268,N_8097,N_8177);
nor U8269 (N_8269,N_8006,N_8140);
or U8270 (N_8270,N_8155,N_8207);
xnor U8271 (N_8271,N_8112,N_8249);
or U8272 (N_8272,N_8007,N_8159);
and U8273 (N_8273,N_8014,N_8020);
xor U8274 (N_8274,N_8199,N_8016);
nor U8275 (N_8275,N_8060,N_8188);
and U8276 (N_8276,N_8022,N_8017);
xor U8277 (N_8277,N_8146,N_8235);
or U8278 (N_8278,N_8206,N_8139);
xnor U8279 (N_8279,N_8059,N_8069);
xnor U8280 (N_8280,N_8190,N_8000);
nor U8281 (N_8281,N_8021,N_8029);
or U8282 (N_8282,N_8125,N_8248);
xor U8283 (N_8283,N_8072,N_8193);
nand U8284 (N_8284,N_8231,N_8138);
nand U8285 (N_8285,N_8213,N_8153);
xor U8286 (N_8286,N_8025,N_8237);
and U8287 (N_8287,N_8001,N_8009);
and U8288 (N_8288,N_8034,N_8042);
or U8289 (N_8289,N_8208,N_8081);
and U8290 (N_8290,N_8238,N_8221);
or U8291 (N_8291,N_8036,N_8243);
nand U8292 (N_8292,N_8149,N_8076);
and U8293 (N_8293,N_8167,N_8108);
nand U8294 (N_8294,N_8145,N_8071);
or U8295 (N_8295,N_8212,N_8051);
xnor U8296 (N_8296,N_8228,N_8030);
or U8297 (N_8297,N_8067,N_8144);
nand U8298 (N_8298,N_8224,N_8160);
nor U8299 (N_8299,N_8063,N_8054);
and U8300 (N_8300,N_8003,N_8133);
or U8301 (N_8301,N_8082,N_8090);
and U8302 (N_8302,N_8178,N_8242);
nor U8303 (N_8303,N_8247,N_8049);
or U8304 (N_8304,N_8245,N_8053);
nor U8305 (N_8305,N_8244,N_8018);
and U8306 (N_8306,N_8151,N_8218);
and U8307 (N_8307,N_8129,N_8152);
nand U8308 (N_8308,N_8137,N_8103);
nor U8309 (N_8309,N_8191,N_8118);
and U8310 (N_8310,N_8120,N_8115);
nand U8311 (N_8311,N_8122,N_8032);
xnor U8312 (N_8312,N_8079,N_8046);
xor U8313 (N_8313,N_8204,N_8229);
and U8314 (N_8314,N_8083,N_8215);
nor U8315 (N_8315,N_8058,N_8107);
or U8316 (N_8316,N_8239,N_8172);
xnor U8317 (N_8317,N_8052,N_8087);
nand U8318 (N_8318,N_8240,N_8220);
nand U8319 (N_8319,N_8236,N_8156);
xnor U8320 (N_8320,N_8075,N_8230);
xor U8321 (N_8321,N_8040,N_8078);
xor U8322 (N_8322,N_8168,N_8089);
or U8323 (N_8323,N_8126,N_8127);
and U8324 (N_8324,N_8197,N_8012);
and U8325 (N_8325,N_8154,N_8181);
nor U8326 (N_8326,N_8047,N_8195);
nand U8327 (N_8327,N_8057,N_8048);
xor U8328 (N_8328,N_8101,N_8134);
nor U8329 (N_8329,N_8124,N_8165);
or U8330 (N_8330,N_8116,N_8234);
xor U8331 (N_8331,N_8070,N_8182);
and U8332 (N_8332,N_8171,N_8131);
xnor U8333 (N_8333,N_8169,N_8128);
xor U8334 (N_8334,N_8158,N_8080);
and U8335 (N_8335,N_8123,N_8225);
xnor U8336 (N_8336,N_8183,N_8109);
nand U8337 (N_8337,N_8246,N_8161);
xnor U8338 (N_8338,N_8179,N_8232);
nor U8339 (N_8339,N_8010,N_8175);
nor U8340 (N_8340,N_8216,N_8106);
and U8341 (N_8341,N_8192,N_8119);
or U8342 (N_8342,N_8073,N_8002);
nand U8343 (N_8343,N_8099,N_8166);
or U8344 (N_8344,N_8096,N_8214);
xnor U8345 (N_8345,N_8196,N_8150);
xor U8346 (N_8346,N_8026,N_8227);
or U8347 (N_8347,N_8028,N_8147);
or U8348 (N_8348,N_8094,N_8113);
and U8349 (N_8349,N_8004,N_8039);
or U8350 (N_8350,N_8061,N_8130);
or U8351 (N_8351,N_8189,N_8186);
nand U8352 (N_8352,N_8035,N_8086);
nand U8353 (N_8353,N_8170,N_8050);
nor U8354 (N_8354,N_8066,N_8055);
and U8355 (N_8355,N_8013,N_8092);
nand U8356 (N_8356,N_8164,N_8148);
nor U8357 (N_8357,N_8174,N_8114);
xor U8358 (N_8358,N_8211,N_8241);
and U8359 (N_8359,N_8163,N_8111);
and U8360 (N_8360,N_8056,N_8084);
and U8361 (N_8361,N_8027,N_8194);
xor U8362 (N_8362,N_8104,N_8132);
nand U8363 (N_8363,N_8100,N_8200);
xnor U8364 (N_8364,N_8110,N_8064);
nand U8365 (N_8365,N_8037,N_8143);
or U8366 (N_8366,N_8222,N_8019);
and U8367 (N_8367,N_8038,N_8098);
nor U8368 (N_8368,N_8135,N_8173);
or U8369 (N_8369,N_8095,N_8141);
or U8370 (N_8370,N_8068,N_8085);
or U8371 (N_8371,N_8024,N_8176);
xor U8372 (N_8372,N_8201,N_8074);
nand U8373 (N_8373,N_8157,N_8121);
or U8374 (N_8374,N_8223,N_8045);
and U8375 (N_8375,N_8039,N_8140);
nand U8376 (N_8376,N_8100,N_8070);
and U8377 (N_8377,N_8174,N_8084);
or U8378 (N_8378,N_8193,N_8206);
nand U8379 (N_8379,N_8213,N_8180);
nand U8380 (N_8380,N_8015,N_8109);
nand U8381 (N_8381,N_8106,N_8070);
and U8382 (N_8382,N_8009,N_8105);
nor U8383 (N_8383,N_8045,N_8115);
nand U8384 (N_8384,N_8037,N_8170);
nand U8385 (N_8385,N_8023,N_8231);
nor U8386 (N_8386,N_8067,N_8085);
nand U8387 (N_8387,N_8014,N_8109);
nor U8388 (N_8388,N_8119,N_8157);
or U8389 (N_8389,N_8198,N_8040);
or U8390 (N_8390,N_8012,N_8193);
nor U8391 (N_8391,N_8197,N_8149);
and U8392 (N_8392,N_8041,N_8148);
nand U8393 (N_8393,N_8191,N_8086);
nor U8394 (N_8394,N_8225,N_8057);
or U8395 (N_8395,N_8231,N_8237);
and U8396 (N_8396,N_8153,N_8094);
nand U8397 (N_8397,N_8003,N_8241);
nor U8398 (N_8398,N_8183,N_8081);
and U8399 (N_8399,N_8022,N_8222);
nand U8400 (N_8400,N_8247,N_8082);
nand U8401 (N_8401,N_8151,N_8140);
and U8402 (N_8402,N_8074,N_8203);
xnor U8403 (N_8403,N_8209,N_8000);
nor U8404 (N_8404,N_8008,N_8230);
xor U8405 (N_8405,N_8221,N_8199);
nand U8406 (N_8406,N_8010,N_8095);
or U8407 (N_8407,N_8176,N_8144);
nand U8408 (N_8408,N_8161,N_8231);
and U8409 (N_8409,N_8051,N_8218);
xor U8410 (N_8410,N_8031,N_8051);
and U8411 (N_8411,N_8154,N_8161);
nor U8412 (N_8412,N_8084,N_8164);
nor U8413 (N_8413,N_8177,N_8242);
or U8414 (N_8414,N_8045,N_8075);
or U8415 (N_8415,N_8107,N_8204);
xnor U8416 (N_8416,N_8125,N_8097);
nand U8417 (N_8417,N_8061,N_8069);
and U8418 (N_8418,N_8172,N_8199);
nand U8419 (N_8419,N_8012,N_8210);
xor U8420 (N_8420,N_8010,N_8096);
xnor U8421 (N_8421,N_8040,N_8136);
nand U8422 (N_8422,N_8014,N_8119);
or U8423 (N_8423,N_8152,N_8046);
and U8424 (N_8424,N_8178,N_8055);
or U8425 (N_8425,N_8231,N_8179);
or U8426 (N_8426,N_8234,N_8113);
and U8427 (N_8427,N_8077,N_8052);
nor U8428 (N_8428,N_8060,N_8121);
and U8429 (N_8429,N_8088,N_8161);
or U8430 (N_8430,N_8032,N_8233);
nand U8431 (N_8431,N_8019,N_8062);
or U8432 (N_8432,N_8067,N_8145);
or U8433 (N_8433,N_8155,N_8102);
xnor U8434 (N_8434,N_8081,N_8219);
nand U8435 (N_8435,N_8146,N_8001);
or U8436 (N_8436,N_8149,N_8006);
xnor U8437 (N_8437,N_8025,N_8236);
nor U8438 (N_8438,N_8062,N_8247);
nor U8439 (N_8439,N_8171,N_8035);
xor U8440 (N_8440,N_8106,N_8098);
and U8441 (N_8441,N_8074,N_8211);
and U8442 (N_8442,N_8160,N_8135);
nor U8443 (N_8443,N_8172,N_8151);
nor U8444 (N_8444,N_8177,N_8100);
or U8445 (N_8445,N_8076,N_8111);
and U8446 (N_8446,N_8019,N_8074);
xnor U8447 (N_8447,N_8019,N_8046);
nand U8448 (N_8448,N_8033,N_8002);
or U8449 (N_8449,N_8099,N_8220);
or U8450 (N_8450,N_8227,N_8041);
and U8451 (N_8451,N_8072,N_8121);
or U8452 (N_8452,N_8147,N_8111);
nand U8453 (N_8453,N_8029,N_8081);
xnor U8454 (N_8454,N_8208,N_8179);
nand U8455 (N_8455,N_8130,N_8188);
xor U8456 (N_8456,N_8068,N_8117);
and U8457 (N_8457,N_8224,N_8010);
and U8458 (N_8458,N_8085,N_8093);
nand U8459 (N_8459,N_8162,N_8051);
xnor U8460 (N_8460,N_8183,N_8002);
nand U8461 (N_8461,N_8140,N_8247);
and U8462 (N_8462,N_8062,N_8207);
xnor U8463 (N_8463,N_8063,N_8127);
nor U8464 (N_8464,N_8189,N_8157);
xor U8465 (N_8465,N_8092,N_8170);
nand U8466 (N_8466,N_8239,N_8086);
xnor U8467 (N_8467,N_8147,N_8170);
xor U8468 (N_8468,N_8003,N_8112);
and U8469 (N_8469,N_8130,N_8186);
or U8470 (N_8470,N_8200,N_8063);
or U8471 (N_8471,N_8086,N_8217);
and U8472 (N_8472,N_8070,N_8167);
or U8473 (N_8473,N_8034,N_8021);
nor U8474 (N_8474,N_8079,N_8025);
nand U8475 (N_8475,N_8137,N_8223);
or U8476 (N_8476,N_8063,N_8016);
nor U8477 (N_8477,N_8010,N_8202);
xnor U8478 (N_8478,N_8025,N_8004);
and U8479 (N_8479,N_8175,N_8235);
and U8480 (N_8480,N_8080,N_8019);
nand U8481 (N_8481,N_8063,N_8201);
or U8482 (N_8482,N_8049,N_8160);
and U8483 (N_8483,N_8213,N_8151);
xnor U8484 (N_8484,N_8236,N_8132);
nor U8485 (N_8485,N_8106,N_8197);
xor U8486 (N_8486,N_8225,N_8077);
nor U8487 (N_8487,N_8239,N_8107);
nor U8488 (N_8488,N_8169,N_8134);
or U8489 (N_8489,N_8150,N_8227);
and U8490 (N_8490,N_8198,N_8131);
nor U8491 (N_8491,N_8103,N_8173);
and U8492 (N_8492,N_8029,N_8155);
nor U8493 (N_8493,N_8010,N_8077);
nor U8494 (N_8494,N_8223,N_8046);
or U8495 (N_8495,N_8162,N_8084);
nand U8496 (N_8496,N_8149,N_8021);
xor U8497 (N_8497,N_8114,N_8231);
and U8498 (N_8498,N_8102,N_8004);
or U8499 (N_8499,N_8111,N_8022);
nand U8500 (N_8500,N_8352,N_8396);
nor U8501 (N_8501,N_8429,N_8499);
nand U8502 (N_8502,N_8377,N_8400);
xnor U8503 (N_8503,N_8361,N_8363);
xnor U8504 (N_8504,N_8468,N_8258);
xnor U8505 (N_8505,N_8279,N_8473);
nand U8506 (N_8506,N_8333,N_8321);
or U8507 (N_8507,N_8327,N_8386);
or U8508 (N_8508,N_8308,N_8381);
nor U8509 (N_8509,N_8455,N_8476);
xnor U8510 (N_8510,N_8304,N_8357);
nand U8511 (N_8511,N_8434,N_8358);
or U8512 (N_8512,N_8413,N_8452);
xor U8513 (N_8513,N_8456,N_8348);
and U8514 (N_8514,N_8447,N_8360);
or U8515 (N_8515,N_8305,N_8376);
nand U8516 (N_8516,N_8469,N_8446);
nand U8517 (N_8517,N_8474,N_8415);
xnor U8518 (N_8518,N_8260,N_8323);
or U8519 (N_8519,N_8438,N_8265);
nor U8520 (N_8520,N_8314,N_8421);
nor U8521 (N_8521,N_8355,N_8387);
or U8522 (N_8522,N_8435,N_8481);
and U8523 (N_8523,N_8382,N_8384);
and U8524 (N_8524,N_8417,N_8310);
and U8525 (N_8525,N_8450,N_8431);
and U8526 (N_8526,N_8458,N_8419);
and U8527 (N_8527,N_8313,N_8418);
or U8528 (N_8528,N_8330,N_8471);
and U8529 (N_8529,N_8251,N_8370);
nand U8530 (N_8530,N_8485,N_8380);
and U8531 (N_8531,N_8273,N_8318);
nand U8532 (N_8532,N_8451,N_8395);
or U8533 (N_8533,N_8495,N_8325);
nor U8534 (N_8534,N_8408,N_8454);
xnor U8535 (N_8535,N_8426,N_8367);
xnor U8536 (N_8536,N_8414,N_8302);
nor U8537 (N_8537,N_8297,N_8269);
and U8538 (N_8538,N_8389,N_8441);
or U8539 (N_8539,N_8420,N_8298);
nor U8540 (N_8540,N_8388,N_8287);
and U8541 (N_8541,N_8393,N_8276);
nor U8542 (N_8542,N_8311,N_8428);
and U8543 (N_8543,N_8394,N_8479);
or U8544 (N_8544,N_8489,N_8339);
or U8545 (N_8545,N_8315,N_8398);
xnor U8546 (N_8546,N_8371,N_8328);
nand U8547 (N_8547,N_8422,N_8493);
xor U8548 (N_8548,N_8296,N_8462);
or U8549 (N_8549,N_8294,N_8404);
nand U8550 (N_8550,N_8280,N_8259);
nor U8551 (N_8551,N_8487,N_8402);
xor U8552 (N_8552,N_8340,N_8320);
nor U8553 (N_8553,N_8436,N_8437);
nor U8554 (N_8554,N_8282,N_8254);
nand U8555 (N_8555,N_8326,N_8263);
xor U8556 (N_8556,N_8406,N_8270);
nand U8557 (N_8557,N_8286,N_8477);
or U8558 (N_8558,N_8427,N_8300);
nor U8559 (N_8559,N_8329,N_8337);
nand U8560 (N_8560,N_8289,N_8264);
xnor U8561 (N_8561,N_8498,N_8409);
nor U8562 (N_8562,N_8262,N_8401);
nand U8563 (N_8563,N_8478,N_8375);
and U8564 (N_8564,N_8484,N_8482);
and U8565 (N_8565,N_8424,N_8342);
or U8566 (N_8566,N_8332,N_8372);
xnor U8567 (N_8567,N_8453,N_8488);
and U8568 (N_8568,N_8354,N_8324);
nor U8569 (N_8569,N_8465,N_8445);
and U8570 (N_8570,N_8459,N_8391);
or U8571 (N_8571,N_8369,N_8309);
nor U8572 (N_8572,N_8299,N_8353);
nand U8573 (N_8573,N_8266,N_8457);
xnor U8574 (N_8574,N_8261,N_8350);
nor U8575 (N_8575,N_8378,N_8356);
xor U8576 (N_8576,N_8442,N_8345);
nor U8577 (N_8577,N_8432,N_8288);
nand U8578 (N_8578,N_8322,N_8317);
xor U8579 (N_8579,N_8491,N_8397);
nor U8580 (N_8580,N_8492,N_8257);
and U8581 (N_8581,N_8433,N_8461);
xor U8582 (N_8582,N_8336,N_8341);
nand U8583 (N_8583,N_8359,N_8272);
nand U8584 (N_8584,N_8448,N_8368);
nor U8585 (N_8585,N_8464,N_8496);
nor U8586 (N_8586,N_8292,N_8365);
or U8587 (N_8587,N_8475,N_8274);
xor U8588 (N_8588,N_8440,N_8449);
and U8589 (N_8589,N_8390,N_8291);
and U8590 (N_8590,N_8307,N_8271);
and U8591 (N_8591,N_8423,N_8425);
xnor U8592 (N_8592,N_8466,N_8439);
and U8593 (N_8593,N_8374,N_8385);
xnor U8594 (N_8594,N_8351,N_8344);
nand U8595 (N_8595,N_8335,N_8347);
nand U8596 (N_8596,N_8331,N_8281);
and U8597 (N_8597,N_8416,N_8410);
or U8598 (N_8598,N_8301,N_8312);
xor U8599 (N_8599,N_8252,N_8366);
and U8600 (N_8600,N_8275,N_8497);
nor U8601 (N_8601,N_8303,N_8490);
nor U8602 (N_8602,N_8486,N_8349);
xor U8603 (N_8603,N_8403,N_8444);
and U8604 (N_8604,N_8306,N_8362);
nand U8605 (N_8605,N_8293,N_8407);
or U8606 (N_8606,N_8277,N_8460);
nand U8607 (N_8607,N_8430,N_8411);
or U8608 (N_8608,N_8284,N_8316);
and U8609 (N_8609,N_8338,N_8250);
nand U8610 (N_8610,N_8483,N_8379);
and U8611 (N_8611,N_8494,N_8373);
xnor U8612 (N_8612,N_8399,N_8405);
or U8613 (N_8613,N_8443,N_8364);
xnor U8614 (N_8614,N_8295,N_8472);
and U8615 (N_8615,N_8392,N_8283);
nand U8616 (N_8616,N_8346,N_8343);
xor U8617 (N_8617,N_8412,N_8470);
nand U8618 (N_8618,N_8319,N_8463);
xor U8619 (N_8619,N_8334,N_8253);
nand U8620 (N_8620,N_8267,N_8290);
nor U8621 (N_8621,N_8467,N_8255);
xor U8622 (N_8622,N_8278,N_8256);
xnor U8623 (N_8623,N_8285,N_8268);
xnor U8624 (N_8624,N_8383,N_8480);
nor U8625 (N_8625,N_8308,N_8422);
nand U8626 (N_8626,N_8265,N_8393);
xnor U8627 (N_8627,N_8341,N_8489);
nand U8628 (N_8628,N_8314,N_8398);
nand U8629 (N_8629,N_8371,N_8482);
and U8630 (N_8630,N_8255,N_8446);
or U8631 (N_8631,N_8445,N_8369);
nor U8632 (N_8632,N_8482,N_8385);
nor U8633 (N_8633,N_8375,N_8365);
or U8634 (N_8634,N_8494,N_8347);
nand U8635 (N_8635,N_8287,N_8365);
and U8636 (N_8636,N_8466,N_8429);
xnor U8637 (N_8637,N_8350,N_8485);
nand U8638 (N_8638,N_8409,N_8344);
nor U8639 (N_8639,N_8401,N_8493);
nand U8640 (N_8640,N_8462,N_8337);
and U8641 (N_8641,N_8373,N_8427);
nor U8642 (N_8642,N_8418,N_8448);
nor U8643 (N_8643,N_8429,N_8347);
nor U8644 (N_8644,N_8273,N_8393);
and U8645 (N_8645,N_8465,N_8338);
nor U8646 (N_8646,N_8434,N_8324);
and U8647 (N_8647,N_8443,N_8293);
or U8648 (N_8648,N_8300,N_8389);
xnor U8649 (N_8649,N_8387,N_8285);
nand U8650 (N_8650,N_8465,N_8401);
nor U8651 (N_8651,N_8400,N_8415);
xnor U8652 (N_8652,N_8313,N_8450);
and U8653 (N_8653,N_8301,N_8442);
nand U8654 (N_8654,N_8331,N_8461);
xnor U8655 (N_8655,N_8398,N_8473);
nor U8656 (N_8656,N_8482,N_8404);
nor U8657 (N_8657,N_8485,N_8442);
nor U8658 (N_8658,N_8477,N_8363);
or U8659 (N_8659,N_8488,N_8376);
or U8660 (N_8660,N_8388,N_8282);
xor U8661 (N_8661,N_8461,N_8428);
xnor U8662 (N_8662,N_8466,N_8411);
or U8663 (N_8663,N_8301,N_8292);
and U8664 (N_8664,N_8306,N_8386);
xor U8665 (N_8665,N_8458,N_8404);
or U8666 (N_8666,N_8338,N_8457);
or U8667 (N_8667,N_8348,N_8491);
or U8668 (N_8668,N_8296,N_8373);
xor U8669 (N_8669,N_8372,N_8300);
and U8670 (N_8670,N_8398,N_8328);
and U8671 (N_8671,N_8336,N_8264);
nand U8672 (N_8672,N_8412,N_8276);
nor U8673 (N_8673,N_8414,N_8308);
and U8674 (N_8674,N_8495,N_8394);
or U8675 (N_8675,N_8441,N_8291);
nand U8676 (N_8676,N_8309,N_8265);
xnor U8677 (N_8677,N_8270,N_8396);
nor U8678 (N_8678,N_8422,N_8413);
nor U8679 (N_8679,N_8282,N_8355);
or U8680 (N_8680,N_8447,N_8267);
or U8681 (N_8681,N_8345,N_8367);
nor U8682 (N_8682,N_8358,N_8471);
nor U8683 (N_8683,N_8461,N_8276);
xnor U8684 (N_8684,N_8250,N_8411);
xnor U8685 (N_8685,N_8259,N_8295);
nor U8686 (N_8686,N_8448,N_8267);
xnor U8687 (N_8687,N_8431,N_8326);
nand U8688 (N_8688,N_8449,N_8324);
nand U8689 (N_8689,N_8402,N_8328);
xor U8690 (N_8690,N_8382,N_8416);
nand U8691 (N_8691,N_8417,N_8306);
xnor U8692 (N_8692,N_8267,N_8446);
xnor U8693 (N_8693,N_8300,N_8465);
and U8694 (N_8694,N_8357,N_8423);
or U8695 (N_8695,N_8435,N_8463);
xor U8696 (N_8696,N_8443,N_8257);
or U8697 (N_8697,N_8412,N_8345);
nor U8698 (N_8698,N_8280,N_8459);
nor U8699 (N_8699,N_8262,N_8446);
or U8700 (N_8700,N_8381,N_8315);
xnor U8701 (N_8701,N_8493,N_8488);
nand U8702 (N_8702,N_8441,N_8296);
nor U8703 (N_8703,N_8465,N_8397);
and U8704 (N_8704,N_8269,N_8410);
nor U8705 (N_8705,N_8327,N_8266);
nor U8706 (N_8706,N_8346,N_8326);
or U8707 (N_8707,N_8498,N_8267);
nand U8708 (N_8708,N_8457,N_8466);
and U8709 (N_8709,N_8380,N_8397);
and U8710 (N_8710,N_8342,N_8343);
and U8711 (N_8711,N_8487,N_8471);
or U8712 (N_8712,N_8315,N_8494);
xor U8713 (N_8713,N_8470,N_8296);
or U8714 (N_8714,N_8371,N_8368);
nor U8715 (N_8715,N_8457,N_8303);
nor U8716 (N_8716,N_8277,N_8436);
or U8717 (N_8717,N_8348,N_8363);
xnor U8718 (N_8718,N_8319,N_8335);
xnor U8719 (N_8719,N_8262,N_8482);
xor U8720 (N_8720,N_8490,N_8293);
xor U8721 (N_8721,N_8328,N_8256);
or U8722 (N_8722,N_8451,N_8413);
nand U8723 (N_8723,N_8453,N_8421);
nor U8724 (N_8724,N_8347,N_8302);
and U8725 (N_8725,N_8485,N_8393);
nand U8726 (N_8726,N_8297,N_8460);
nand U8727 (N_8727,N_8312,N_8330);
nand U8728 (N_8728,N_8488,N_8394);
and U8729 (N_8729,N_8346,N_8364);
or U8730 (N_8730,N_8394,N_8450);
nor U8731 (N_8731,N_8427,N_8479);
and U8732 (N_8732,N_8419,N_8314);
and U8733 (N_8733,N_8436,N_8450);
nand U8734 (N_8734,N_8377,N_8313);
nor U8735 (N_8735,N_8398,N_8395);
or U8736 (N_8736,N_8431,N_8393);
and U8737 (N_8737,N_8280,N_8461);
xor U8738 (N_8738,N_8405,N_8430);
xor U8739 (N_8739,N_8294,N_8320);
and U8740 (N_8740,N_8268,N_8266);
nand U8741 (N_8741,N_8443,N_8406);
xor U8742 (N_8742,N_8251,N_8389);
xnor U8743 (N_8743,N_8448,N_8381);
or U8744 (N_8744,N_8493,N_8450);
and U8745 (N_8745,N_8364,N_8353);
nor U8746 (N_8746,N_8436,N_8365);
xnor U8747 (N_8747,N_8410,N_8296);
nand U8748 (N_8748,N_8447,N_8331);
and U8749 (N_8749,N_8350,N_8360);
and U8750 (N_8750,N_8636,N_8668);
and U8751 (N_8751,N_8658,N_8531);
and U8752 (N_8752,N_8656,N_8663);
xnor U8753 (N_8753,N_8506,N_8640);
nor U8754 (N_8754,N_8721,N_8715);
nand U8755 (N_8755,N_8562,N_8675);
nand U8756 (N_8756,N_8536,N_8699);
xnor U8757 (N_8757,N_8652,N_8690);
and U8758 (N_8758,N_8623,N_8530);
nand U8759 (N_8759,N_8559,N_8748);
or U8760 (N_8760,N_8581,N_8518);
xnor U8761 (N_8761,N_8547,N_8705);
nor U8762 (N_8762,N_8622,N_8621);
nand U8763 (N_8763,N_8510,N_8661);
xor U8764 (N_8764,N_8588,N_8679);
nor U8765 (N_8765,N_8599,N_8670);
or U8766 (N_8766,N_8578,N_8647);
or U8767 (N_8767,N_8589,N_8501);
nand U8768 (N_8768,N_8740,N_8685);
nand U8769 (N_8769,N_8565,N_8645);
and U8770 (N_8770,N_8520,N_8602);
nand U8771 (N_8771,N_8664,N_8720);
or U8772 (N_8772,N_8634,N_8724);
nand U8773 (N_8773,N_8537,N_8567);
or U8774 (N_8774,N_8655,N_8545);
or U8775 (N_8775,N_8666,N_8557);
nand U8776 (N_8776,N_8593,N_8564);
xor U8777 (N_8777,N_8500,N_8734);
nand U8778 (N_8778,N_8672,N_8612);
nand U8779 (N_8779,N_8566,N_8582);
nand U8780 (N_8780,N_8717,N_8569);
xor U8781 (N_8781,N_8563,N_8525);
nand U8782 (N_8782,N_8575,N_8597);
or U8783 (N_8783,N_8628,N_8613);
nor U8784 (N_8784,N_8702,N_8727);
xor U8785 (N_8785,N_8519,N_8718);
nor U8786 (N_8786,N_8529,N_8576);
xnor U8787 (N_8787,N_8744,N_8732);
nand U8788 (N_8788,N_8590,N_8541);
xnor U8789 (N_8789,N_8696,N_8741);
or U8790 (N_8790,N_8616,N_8714);
or U8791 (N_8791,N_8642,N_8708);
or U8792 (N_8792,N_8502,N_8669);
xnor U8793 (N_8793,N_8644,N_8643);
nand U8794 (N_8794,N_8538,N_8695);
xnor U8795 (N_8795,N_8604,N_8657);
or U8796 (N_8796,N_8677,N_8553);
nand U8797 (N_8797,N_8646,N_8585);
or U8798 (N_8798,N_8701,N_8710);
or U8799 (N_8799,N_8684,N_8624);
and U8800 (N_8800,N_8505,N_8517);
xnor U8801 (N_8801,N_8521,N_8507);
nor U8802 (N_8802,N_8596,N_8697);
nor U8803 (N_8803,N_8549,N_8735);
and U8804 (N_8804,N_8629,N_8554);
nor U8805 (N_8805,N_8625,N_8598);
nand U8806 (N_8806,N_8686,N_8560);
xor U8807 (N_8807,N_8676,N_8733);
or U8808 (N_8808,N_8546,N_8595);
xnor U8809 (N_8809,N_8706,N_8561);
nand U8810 (N_8810,N_8739,N_8527);
nor U8811 (N_8811,N_8609,N_8680);
nor U8812 (N_8812,N_8713,N_8522);
and U8813 (N_8813,N_8660,N_8535);
nor U8814 (N_8814,N_8511,N_8515);
nor U8815 (N_8815,N_8601,N_8618);
nor U8816 (N_8816,N_8540,N_8681);
and U8817 (N_8817,N_8722,N_8558);
and U8818 (N_8818,N_8700,N_8610);
nor U8819 (N_8819,N_8580,N_8725);
nand U8820 (N_8820,N_8620,N_8641);
and U8821 (N_8821,N_8552,N_8745);
nand U8822 (N_8822,N_8528,N_8539);
nor U8823 (N_8823,N_8627,N_8587);
or U8824 (N_8824,N_8551,N_8683);
xor U8825 (N_8825,N_8736,N_8572);
and U8826 (N_8826,N_8555,N_8550);
xor U8827 (N_8827,N_8606,N_8692);
nand U8828 (N_8828,N_8514,N_8543);
and U8829 (N_8829,N_8665,N_8548);
or U8830 (N_8830,N_8698,N_8503);
nand U8831 (N_8831,N_8586,N_8707);
nor U8832 (N_8832,N_8730,N_8654);
or U8833 (N_8833,N_8533,N_8594);
or U8834 (N_8834,N_8523,N_8703);
nand U8835 (N_8835,N_8607,N_8731);
or U8836 (N_8836,N_8632,N_8687);
and U8837 (N_8837,N_8704,N_8611);
and U8838 (N_8838,N_8556,N_8694);
nand U8839 (N_8839,N_8630,N_8746);
xnor U8840 (N_8840,N_8678,N_8508);
xnor U8841 (N_8841,N_8544,N_8579);
nand U8842 (N_8842,N_8693,N_8749);
or U8843 (N_8843,N_8526,N_8709);
nand U8844 (N_8844,N_8716,N_8738);
xnor U8845 (N_8845,N_8723,N_8592);
or U8846 (N_8846,N_8516,N_8649);
and U8847 (N_8847,N_8639,N_8637);
or U8848 (N_8848,N_8577,N_8673);
or U8849 (N_8849,N_8615,N_8534);
nand U8850 (N_8850,N_8743,N_8667);
nand U8851 (N_8851,N_8619,N_8568);
nor U8852 (N_8852,N_8728,N_8617);
nand U8853 (N_8853,N_8712,N_8726);
nor U8854 (N_8854,N_8729,N_8650);
xnor U8855 (N_8855,N_8513,N_8682);
xnor U8856 (N_8856,N_8653,N_8659);
and U8857 (N_8857,N_8689,N_8651);
or U8858 (N_8858,N_8691,N_8635);
xor U8859 (N_8859,N_8742,N_8737);
nand U8860 (N_8860,N_8570,N_8747);
nand U8861 (N_8861,N_8674,N_8608);
nor U8862 (N_8862,N_8671,N_8631);
nor U8863 (N_8863,N_8600,N_8583);
xnor U8864 (N_8864,N_8626,N_8584);
nor U8865 (N_8865,N_8648,N_8532);
or U8866 (N_8866,N_8638,N_8603);
xnor U8867 (N_8867,N_8711,N_8571);
nor U8868 (N_8868,N_8614,N_8662);
xor U8869 (N_8869,N_8509,N_8574);
nor U8870 (N_8870,N_8719,N_8524);
and U8871 (N_8871,N_8591,N_8688);
or U8872 (N_8872,N_8605,N_8633);
and U8873 (N_8873,N_8542,N_8512);
or U8874 (N_8874,N_8573,N_8504);
and U8875 (N_8875,N_8639,N_8710);
nand U8876 (N_8876,N_8602,N_8603);
nor U8877 (N_8877,N_8591,N_8656);
and U8878 (N_8878,N_8749,N_8526);
nor U8879 (N_8879,N_8525,N_8725);
and U8880 (N_8880,N_8698,N_8630);
xnor U8881 (N_8881,N_8609,N_8637);
xor U8882 (N_8882,N_8576,N_8615);
or U8883 (N_8883,N_8725,N_8656);
or U8884 (N_8884,N_8742,N_8570);
and U8885 (N_8885,N_8671,N_8741);
and U8886 (N_8886,N_8672,N_8550);
xnor U8887 (N_8887,N_8534,N_8670);
nor U8888 (N_8888,N_8559,N_8685);
nand U8889 (N_8889,N_8748,N_8669);
nand U8890 (N_8890,N_8510,N_8671);
nor U8891 (N_8891,N_8747,N_8519);
or U8892 (N_8892,N_8706,N_8617);
nor U8893 (N_8893,N_8536,N_8748);
and U8894 (N_8894,N_8618,N_8517);
xor U8895 (N_8895,N_8515,N_8625);
nor U8896 (N_8896,N_8700,N_8665);
nand U8897 (N_8897,N_8605,N_8532);
and U8898 (N_8898,N_8573,N_8664);
nor U8899 (N_8899,N_8656,N_8735);
or U8900 (N_8900,N_8728,N_8731);
and U8901 (N_8901,N_8547,N_8504);
xnor U8902 (N_8902,N_8640,N_8687);
or U8903 (N_8903,N_8600,N_8687);
nand U8904 (N_8904,N_8700,N_8663);
nor U8905 (N_8905,N_8737,N_8531);
xnor U8906 (N_8906,N_8713,N_8661);
xnor U8907 (N_8907,N_8742,N_8512);
and U8908 (N_8908,N_8689,N_8509);
nand U8909 (N_8909,N_8717,N_8567);
xnor U8910 (N_8910,N_8623,N_8520);
and U8911 (N_8911,N_8648,N_8530);
or U8912 (N_8912,N_8728,N_8749);
xnor U8913 (N_8913,N_8588,N_8713);
nor U8914 (N_8914,N_8556,N_8635);
xnor U8915 (N_8915,N_8714,N_8649);
xnor U8916 (N_8916,N_8591,N_8509);
and U8917 (N_8917,N_8549,N_8542);
or U8918 (N_8918,N_8567,N_8518);
xnor U8919 (N_8919,N_8603,N_8559);
nor U8920 (N_8920,N_8676,N_8625);
nor U8921 (N_8921,N_8601,N_8619);
nand U8922 (N_8922,N_8550,N_8737);
nor U8923 (N_8923,N_8622,N_8591);
or U8924 (N_8924,N_8707,N_8612);
and U8925 (N_8925,N_8558,N_8595);
xor U8926 (N_8926,N_8738,N_8575);
and U8927 (N_8927,N_8531,N_8565);
or U8928 (N_8928,N_8500,N_8636);
and U8929 (N_8929,N_8533,N_8680);
and U8930 (N_8930,N_8552,N_8574);
nand U8931 (N_8931,N_8500,N_8612);
nand U8932 (N_8932,N_8641,N_8522);
xor U8933 (N_8933,N_8672,N_8515);
nor U8934 (N_8934,N_8559,N_8615);
nand U8935 (N_8935,N_8646,N_8501);
and U8936 (N_8936,N_8530,N_8596);
or U8937 (N_8937,N_8710,N_8743);
or U8938 (N_8938,N_8744,N_8697);
nand U8939 (N_8939,N_8519,N_8545);
nand U8940 (N_8940,N_8634,N_8573);
nand U8941 (N_8941,N_8604,N_8610);
or U8942 (N_8942,N_8599,N_8595);
or U8943 (N_8943,N_8727,N_8675);
nor U8944 (N_8944,N_8539,N_8745);
nand U8945 (N_8945,N_8694,N_8614);
or U8946 (N_8946,N_8613,N_8736);
nand U8947 (N_8947,N_8504,N_8728);
nand U8948 (N_8948,N_8544,N_8721);
nor U8949 (N_8949,N_8673,N_8671);
and U8950 (N_8950,N_8535,N_8553);
and U8951 (N_8951,N_8617,N_8627);
or U8952 (N_8952,N_8534,N_8642);
nor U8953 (N_8953,N_8560,N_8621);
and U8954 (N_8954,N_8592,N_8703);
nor U8955 (N_8955,N_8557,N_8708);
and U8956 (N_8956,N_8743,N_8697);
and U8957 (N_8957,N_8727,N_8629);
xor U8958 (N_8958,N_8745,N_8652);
xor U8959 (N_8959,N_8624,N_8578);
nand U8960 (N_8960,N_8597,N_8578);
nor U8961 (N_8961,N_8625,N_8507);
nand U8962 (N_8962,N_8576,N_8611);
xor U8963 (N_8963,N_8527,N_8623);
nor U8964 (N_8964,N_8528,N_8565);
nor U8965 (N_8965,N_8701,N_8537);
nand U8966 (N_8966,N_8503,N_8507);
and U8967 (N_8967,N_8690,N_8521);
nor U8968 (N_8968,N_8615,N_8638);
and U8969 (N_8969,N_8523,N_8543);
and U8970 (N_8970,N_8586,N_8735);
xor U8971 (N_8971,N_8614,N_8585);
nand U8972 (N_8972,N_8695,N_8681);
and U8973 (N_8973,N_8686,N_8616);
xor U8974 (N_8974,N_8552,N_8747);
and U8975 (N_8975,N_8596,N_8718);
or U8976 (N_8976,N_8656,N_8731);
or U8977 (N_8977,N_8744,N_8509);
or U8978 (N_8978,N_8589,N_8534);
or U8979 (N_8979,N_8660,N_8740);
nor U8980 (N_8980,N_8587,N_8651);
or U8981 (N_8981,N_8594,N_8534);
or U8982 (N_8982,N_8680,N_8688);
and U8983 (N_8983,N_8607,N_8501);
and U8984 (N_8984,N_8578,N_8608);
nand U8985 (N_8985,N_8521,N_8660);
nand U8986 (N_8986,N_8711,N_8632);
xor U8987 (N_8987,N_8579,N_8542);
and U8988 (N_8988,N_8710,N_8542);
nor U8989 (N_8989,N_8526,N_8568);
xnor U8990 (N_8990,N_8536,N_8562);
and U8991 (N_8991,N_8729,N_8719);
xnor U8992 (N_8992,N_8529,N_8673);
and U8993 (N_8993,N_8542,N_8598);
nor U8994 (N_8994,N_8699,N_8701);
nor U8995 (N_8995,N_8600,N_8543);
nor U8996 (N_8996,N_8578,N_8717);
or U8997 (N_8997,N_8527,N_8573);
and U8998 (N_8998,N_8551,N_8610);
or U8999 (N_8999,N_8598,N_8666);
nand U9000 (N_9000,N_8883,N_8991);
or U9001 (N_9001,N_8844,N_8988);
and U9002 (N_9002,N_8816,N_8808);
or U9003 (N_9003,N_8912,N_8961);
xnor U9004 (N_9004,N_8923,N_8751);
nor U9005 (N_9005,N_8801,N_8983);
or U9006 (N_9006,N_8812,N_8900);
or U9007 (N_9007,N_8794,N_8953);
xor U9008 (N_9008,N_8821,N_8978);
or U9009 (N_9009,N_8885,N_8916);
nand U9010 (N_9010,N_8835,N_8798);
nor U9011 (N_9011,N_8946,N_8926);
and U9012 (N_9012,N_8990,N_8815);
and U9013 (N_9013,N_8898,N_8968);
and U9014 (N_9014,N_8967,N_8787);
or U9015 (N_9015,N_8992,N_8868);
nand U9016 (N_9016,N_8754,N_8833);
xor U9017 (N_9017,N_8939,N_8804);
xnor U9018 (N_9018,N_8929,N_8799);
xnor U9019 (N_9019,N_8826,N_8897);
or U9020 (N_9020,N_8889,N_8874);
xnor U9021 (N_9021,N_8764,N_8785);
nor U9022 (N_9022,N_8811,N_8981);
nand U9023 (N_9023,N_8843,N_8849);
and U9024 (N_9024,N_8913,N_8860);
and U9025 (N_9025,N_8925,N_8813);
nor U9026 (N_9026,N_8862,N_8959);
and U9027 (N_9027,N_8853,N_8822);
or U9028 (N_9028,N_8872,N_8841);
nor U9029 (N_9029,N_8884,N_8907);
and U9030 (N_9030,N_8784,N_8979);
or U9031 (N_9031,N_8899,N_8768);
nand U9032 (N_9032,N_8984,N_8788);
or U9033 (N_9033,N_8938,N_8765);
xnor U9034 (N_9034,N_8850,N_8996);
nor U9035 (N_9035,N_8937,N_8891);
and U9036 (N_9036,N_8973,N_8831);
xnor U9037 (N_9037,N_8987,N_8915);
nand U9038 (N_9038,N_8893,N_8917);
xor U9039 (N_9039,N_8886,N_8905);
nand U9040 (N_9040,N_8875,N_8969);
xnor U9041 (N_9041,N_8944,N_8920);
nand U9042 (N_9042,N_8772,N_8780);
nand U9043 (N_9043,N_8910,N_8753);
xnor U9044 (N_9044,N_8999,N_8796);
and U9045 (N_9045,N_8790,N_8773);
and U9046 (N_9046,N_8805,N_8976);
xor U9047 (N_9047,N_8792,N_8986);
nand U9048 (N_9048,N_8966,N_8834);
and U9049 (N_9049,N_8750,N_8774);
or U9050 (N_9050,N_8896,N_8894);
and U9051 (N_9051,N_8838,N_8881);
nand U9052 (N_9052,N_8880,N_8775);
nor U9053 (N_9053,N_8827,N_8975);
nor U9054 (N_9054,N_8857,N_8809);
nand U9055 (N_9055,N_8824,N_8895);
nor U9056 (N_9056,N_8779,N_8914);
or U9057 (N_9057,N_8947,N_8807);
or U9058 (N_9058,N_8935,N_8830);
or U9059 (N_9059,N_8758,N_8819);
xnor U9060 (N_9060,N_8771,N_8803);
nor U9061 (N_9061,N_8806,N_8814);
nor U9062 (N_9062,N_8823,N_8802);
or U9063 (N_9063,N_8980,N_8783);
and U9064 (N_9064,N_8972,N_8954);
nor U9065 (N_9065,N_8882,N_8852);
or U9066 (N_9066,N_8970,N_8951);
or U9067 (N_9067,N_8964,N_8859);
xor U9068 (N_9068,N_8836,N_8977);
xnor U9069 (N_9069,N_8791,N_8948);
nand U9070 (N_9070,N_8845,N_8778);
xor U9071 (N_9071,N_8861,N_8867);
or U9072 (N_9072,N_8847,N_8931);
xnor U9073 (N_9073,N_8865,N_8924);
or U9074 (N_9074,N_8878,N_8869);
nand U9075 (N_9075,N_8928,N_8846);
and U9076 (N_9076,N_8909,N_8763);
and U9077 (N_9077,N_8974,N_8797);
nor U9078 (N_9078,N_8837,N_8877);
xor U9079 (N_9079,N_8902,N_8820);
xor U9080 (N_9080,N_8871,N_8918);
or U9081 (N_9081,N_8933,N_8793);
nand U9082 (N_9082,N_8906,N_8858);
xor U9083 (N_9083,N_8864,N_8795);
or U9084 (N_9084,N_8776,N_8848);
nor U9085 (N_9085,N_8901,N_8777);
and U9086 (N_9086,N_8840,N_8766);
xnor U9087 (N_9087,N_8919,N_8839);
and U9088 (N_9088,N_8866,N_8940);
nor U9089 (N_9089,N_8958,N_8985);
or U9090 (N_9090,N_8943,N_8922);
xnor U9091 (N_9091,N_8876,N_8971);
nand U9092 (N_9092,N_8911,N_8769);
and U9093 (N_9093,N_8851,N_8952);
and U9094 (N_9094,N_8781,N_8760);
nand U9095 (N_9095,N_8927,N_8829);
nand U9096 (N_9096,N_8989,N_8892);
xor U9097 (N_9097,N_8908,N_8817);
nand U9098 (N_9098,N_8904,N_8782);
nor U9099 (N_9099,N_8761,N_8998);
xor U9100 (N_9100,N_8993,N_8887);
and U9101 (N_9101,N_8767,N_8879);
and U9102 (N_9102,N_8888,N_8962);
and U9103 (N_9103,N_8965,N_8936);
nor U9104 (N_9104,N_8873,N_8762);
nor U9105 (N_9105,N_8994,N_8800);
and U9106 (N_9106,N_8810,N_8995);
or U9107 (N_9107,N_8756,N_8832);
or U9108 (N_9108,N_8842,N_8942);
and U9109 (N_9109,N_8863,N_8997);
and U9110 (N_9110,N_8870,N_8960);
nor U9111 (N_9111,N_8855,N_8755);
nand U9112 (N_9112,N_8770,N_8890);
nand U9113 (N_9113,N_8955,N_8818);
nor U9114 (N_9114,N_8956,N_8945);
xnor U9115 (N_9115,N_8903,N_8934);
nor U9116 (N_9116,N_8982,N_8957);
nor U9117 (N_9117,N_8921,N_8825);
nand U9118 (N_9118,N_8757,N_8963);
xor U9119 (N_9119,N_8759,N_8856);
and U9120 (N_9120,N_8941,N_8949);
and U9121 (N_9121,N_8828,N_8786);
and U9122 (N_9122,N_8950,N_8789);
and U9123 (N_9123,N_8854,N_8930);
xnor U9124 (N_9124,N_8752,N_8932);
nor U9125 (N_9125,N_8775,N_8818);
nand U9126 (N_9126,N_8909,N_8948);
xor U9127 (N_9127,N_8842,N_8963);
and U9128 (N_9128,N_8943,N_8804);
or U9129 (N_9129,N_8966,N_8751);
xnor U9130 (N_9130,N_8850,N_8855);
nor U9131 (N_9131,N_8795,N_8848);
nand U9132 (N_9132,N_8797,N_8779);
and U9133 (N_9133,N_8889,N_8925);
nor U9134 (N_9134,N_8751,N_8847);
and U9135 (N_9135,N_8859,N_8771);
nand U9136 (N_9136,N_8869,N_8898);
xor U9137 (N_9137,N_8999,N_8898);
nor U9138 (N_9138,N_8855,N_8839);
nor U9139 (N_9139,N_8952,N_8765);
xor U9140 (N_9140,N_8757,N_8933);
xnor U9141 (N_9141,N_8821,N_8844);
nor U9142 (N_9142,N_8866,N_8919);
xor U9143 (N_9143,N_8949,N_8993);
xnor U9144 (N_9144,N_8938,N_8795);
or U9145 (N_9145,N_8800,N_8897);
nor U9146 (N_9146,N_8826,N_8819);
nand U9147 (N_9147,N_8996,N_8882);
nand U9148 (N_9148,N_8862,N_8914);
xnor U9149 (N_9149,N_8774,N_8807);
nor U9150 (N_9150,N_8891,N_8754);
and U9151 (N_9151,N_8946,N_8890);
or U9152 (N_9152,N_8864,N_8794);
xnor U9153 (N_9153,N_8790,N_8863);
and U9154 (N_9154,N_8803,N_8995);
nand U9155 (N_9155,N_8778,N_8903);
nand U9156 (N_9156,N_8920,N_8858);
xnor U9157 (N_9157,N_8967,N_8786);
nor U9158 (N_9158,N_8771,N_8921);
nor U9159 (N_9159,N_8955,N_8757);
xnor U9160 (N_9160,N_8958,N_8812);
nand U9161 (N_9161,N_8799,N_8926);
nand U9162 (N_9162,N_8899,N_8860);
nand U9163 (N_9163,N_8969,N_8894);
xor U9164 (N_9164,N_8929,N_8770);
nand U9165 (N_9165,N_8826,N_8813);
xnor U9166 (N_9166,N_8851,N_8797);
nor U9167 (N_9167,N_8833,N_8783);
or U9168 (N_9168,N_8936,N_8811);
and U9169 (N_9169,N_8817,N_8999);
nor U9170 (N_9170,N_8896,N_8912);
nand U9171 (N_9171,N_8953,N_8832);
and U9172 (N_9172,N_8904,N_8925);
and U9173 (N_9173,N_8814,N_8780);
xnor U9174 (N_9174,N_8945,N_8840);
and U9175 (N_9175,N_8830,N_8801);
xor U9176 (N_9176,N_8821,N_8916);
nor U9177 (N_9177,N_8927,N_8885);
nor U9178 (N_9178,N_8956,N_8794);
and U9179 (N_9179,N_8941,N_8769);
nor U9180 (N_9180,N_8941,N_8913);
nor U9181 (N_9181,N_8918,N_8819);
nor U9182 (N_9182,N_8921,N_8917);
or U9183 (N_9183,N_8768,N_8874);
xor U9184 (N_9184,N_8997,N_8756);
or U9185 (N_9185,N_8818,N_8778);
xor U9186 (N_9186,N_8862,N_8904);
or U9187 (N_9187,N_8936,N_8795);
nand U9188 (N_9188,N_8855,N_8929);
nor U9189 (N_9189,N_8804,N_8867);
and U9190 (N_9190,N_8757,N_8961);
and U9191 (N_9191,N_8807,N_8783);
xor U9192 (N_9192,N_8841,N_8882);
xnor U9193 (N_9193,N_8889,N_8956);
nand U9194 (N_9194,N_8847,N_8937);
or U9195 (N_9195,N_8853,N_8830);
nor U9196 (N_9196,N_8774,N_8789);
xnor U9197 (N_9197,N_8911,N_8783);
nand U9198 (N_9198,N_8809,N_8802);
nor U9199 (N_9199,N_8817,N_8945);
or U9200 (N_9200,N_8993,N_8792);
xor U9201 (N_9201,N_8853,N_8990);
nand U9202 (N_9202,N_8832,N_8840);
nand U9203 (N_9203,N_8826,N_8937);
nand U9204 (N_9204,N_8772,N_8995);
nor U9205 (N_9205,N_8820,N_8778);
nor U9206 (N_9206,N_8881,N_8953);
nor U9207 (N_9207,N_8796,N_8827);
xor U9208 (N_9208,N_8792,N_8777);
xnor U9209 (N_9209,N_8751,N_8860);
nor U9210 (N_9210,N_8798,N_8990);
and U9211 (N_9211,N_8794,N_8942);
xnor U9212 (N_9212,N_8844,N_8890);
xor U9213 (N_9213,N_8910,N_8976);
xor U9214 (N_9214,N_8790,N_8824);
nand U9215 (N_9215,N_8784,N_8942);
xnor U9216 (N_9216,N_8802,N_8853);
xnor U9217 (N_9217,N_8798,N_8979);
and U9218 (N_9218,N_8870,N_8792);
xnor U9219 (N_9219,N_8945,N_8950);
or U9220 (N_9220,N_8771,N_8991);
nand U9221 (N_9221,N_8912,N_8954);
and U9222 (N_9222,N_8856,N_8779);
nand U9223 (N_9223,N_8922,N_8954);
nand U9224 (N_9224,N_8869,N_8824);
nand U9225 (N_9225,N_8833,N_8929);
or U9226 (N_9226,N_8941,N_8918);
nor U9227 (N_9227,N_8942,N_8881);
nand U9228 (N_9228,N_8930,N_8898);
or U9229 (N_9229,N_8804,N_8881);
nor U9230 (N_9230,N_8953,N_8951);
or U9231 (N_9231,N_8971,N_8897);
xor U9232 (N_9232,N_8827,N_8795);
nand U9233 (N_9233,N_8918,N_8790);
nor U9234 (N_9234,N_8764,N_8816);
nand U9235 (N_9235,N_8758,N_8976);
nor U9236 (N_9236,N_8847,N_8790);
nor U9237 (N_9237,N_8974,N_8780);
nand U9238 (N_9238,N_8791,N_8860);
nor U9239 (N_9239,N_8896,N_8945);
xor U9240 (N_9240,N_8764,N_8938);
xor U9241 (N_9241,N_8799,N_8952);
xor U9242 (N_9242,N_8868,N_8996);
nand U9243 (N_9243,N_8866,N_8763);
nand U9244 (N_9244,N_8985,N_8800);
xor U9245 (N_9245,N_8895,N_8839);
and U9246 (N_9246,N_8991,N_8862);
or U9247 (N_9247,N_8786,N_8846);
or U9248 (N_9248,N_8902,N_8999);
nand U9249 (N_9249,N_8790,N_8905);
and U9250 (N_9250,N_9196,N_9142);
xnor U9251 (N_9251,N_9080,N_9189);
nor U9252 (N_9252,N_9211,N_9095);
or U9253 (N_9253,N_9069,N_9234);
nor U9254 (N_9254,N_9081,N_9088);
or U9255 (N_9255,N_9181,N_9191);
nor U9256 (N_9256,N_9216,N_9085);
nor U9257 (N_9257,N_9140,N_9035);
xnor U9258 (N_9258,N_9056,N_9032);
nor U9259 (N_9259,N_9029,N_9052);
nand U9260 (N_9260,N_9133,N_9022);
or U9261 (N_9261,N_9010,N_9223);
nor U9262 (N_9262,N_9147,N_9040);
and U9263 (N_9263,N_9113,N_9242);
and U9264 (N_9264,N_9114,N_9003);
and U9265 (N_9265,N_9120,N_9155);
xor U9266 (N_9266,N_9002,N_9007);
nor U9267 (N_9267,N_9031,N_9129);
and U9268 (N_9268,N_9078,N_9084);
nor U9269 (N_9269,N_9206,N_9004);
or U9270 (N_9270,N_9062,N_9188);
nor U9271 (N_9271,N_9187,N_9126);
nor U9272 (N_9272,N_9030,N_9121);
nor U9273 (N_9273,N_9238,N_9146);
nand U9274 (N_9274,N_9009,N_9170);
and U9275 (N_9275,N_9151,N_9186);
nand U9276 (N_9276,N_9145,N_9075);
or U9277 (N_9277,N_9054,N_9159);
or U9278 (N_9278,N_9177,N_9039);
nor U9279 (N_9279,N_9005,N_9101);
or U9280 (N_9280,N_9082,N_9086);
nor U9281 (N_9281,N_9135,N_9201);
xor U9282 (N_9282,N_9094,N_9046);
or U9283 (N_9283,N_9018,N_9106);
and U9284 (N_9284,N_9225,N_9090);
nand U9285 (N_9285,N_9228,N_9066);
nand U9286 (N_9286,N_9163,N_9027);
or U9287 (N_9287,N_9233,N_9100);
and U9288 (N_9288,N_9131,N_9092);
nor U9289 (N_9289,N_9011,N_9128);
nor U9290 (N_9290,N_9025,N_9174);
nand U9291 (N_9291,N_9134,N_9227);
xnor U9292 (N_9292,N_9093,N_9143);
xnor U9293 (N_9293,N_9105,N_9117);
nand U9294 (N_9294,N_9026,N_9068);
xor U9295 (N_9295,N_9023,N_9049);
nor U9296 (N_9296,N_9115,N_9184);
nor U9297 (N_9297,N_9214,N_9125);
or U9298 (N_9298,N_9110,N_9220);
xor U9299 (N_9299,N_9083,N_9226);
nand U9300 (N_9300,N_9042,N_9122);
xnor U9301 (N_9301,N_9195,N_9243);
xnor U9302 (N_9302,N_9169,N_9099);
or U9303 (N_9303,N_9192,N_9034);
and U9304 (N_9304,N_9141,N_9176);
xnor U9305 (N_9305,N_9229,N_9076);
nor U9306 (N_9306,N_9213,N_9036);
and U9307 (N_9307,N_9098,N_9240);
or U9308 (N_9308,N_9070,N_9179);
nor U9309 (N_9309,N_9212,N_9047);
or U9310 (N_9310,N_9059,N_9183);
and U9311 (N_9311,N_9118,N_9246);
or U9312 (N_9312,N_9157,N_9158);
nand U9313 (N_9313,N_9130,N_9116);
and U9314 (N_9314,N_9015,N_9087);
nor U9315 (N_9315,N_9019,N_9153);
xnor U9316 (N_9316,N_9139,N_9150);
or U9317 (N_9317,N_9205,N_9180);
and U9318 (N_9318,N_9199,N_9058);
and U9319 (N_9319,N_9245,N_9045);
or U9320 (N_9320,N_9171,N_9091);
nor U9321 (N_9321,N_9144,N_9063);
nor U9322 (N_9322,N_9020,N_9102);
xnor U9323 (N_9323,N_9111,N_9182);
xnor U9324 (N_9324,N_9152,N_9073);
xnor U9325 (N_9325,N_9221,N_9044);
or U9326 (N_9326,N_9048,N_9248);
or U9327 (N_9327,N_9024,N_9000);
and U9328 (N_9328,N_9190,N_9249);
xor U9329 (N_9329,N_9060,N_9200);
and U9330 (N_9330,N_9028,N_9198);
and U9331 (N_9331,N_9232,N_9108);
and U9332 (N_9332,N_9197,N_9097);
or U9333 (N_9333,N_9231,N_9241);
nor U9334 (N_9334,N_9137,N_9154);
nand U9335 (N_9335,N_9001,N_9017);
and U9336 (N_9336,N_9193,N_9104);
and U9337 (N_9337,N_9037,N_9168);
and U9338 (N_9338,N_9235,N_9178);
or U9339 (N_9339,N_9239,N_9209);
or U9340 (N_9340,N_9132,N_9013);
nor U9341 (N_9341,N_9172,N_9127);
nor U9342 (N_9342,N_9204,N_9096);
nor U9343 (N_9343,N_9203,N_9202);
nand U9344 (N_9344,N_9208,N_9247);
and U9345 (N_9345,N_9072,N_9112);
nor U9346 (N_9346,N_9149,N_9043);
xor U9347 (N_9347,N_9021,N_9016);
xor U9348 (N_9348,N_9038,N_9051);
nor U9349 (N_9349,N_9218,N_9207);
and U9350 (N_9350,N_9156,N_9064);
xnor U9351 (N_9351,N_9103,N_9077);
xnor U9352 (N_9352,N_9160,N_9175);
xnor U9353 (N_9353,N_9210,N_9053);
nor U9354 (N_9354,N_9014,N_9185);
xnor U9355 (N_9355,N_9161,N_9167);
nand U9356 (N_9356,N_9065,N_9074);
nand U9357 (N_9357,N_9119,N_9057);
and U9358 (N_9358,N_9164,N_9236);
nor U9359 (N_9359,N_9107,N_9244);
and U9360 (N_9360,N_9165,N_9162);
nand U9361 (N_9361,N_9215,N_9109);
or U9362 (N_9362,N_9061,N_9071);
nor U9363 (N_9363,N_9123,N_9230);
nand U9364 (N_9364,N_9148,N_9041);
nand U9365 (N_9365,N_9219,N_9166);
and U9366 (N_9366,N_9124,N_9012);
or U9367 (N_9367,N_9067,N_9224);
nand U9368 (N_9368,N_9050,N_9079);
nor U9369 (N_9369,N_9237,N_9089);
nand U9370 (N_9370,N_9136,N_9173);
nor U9371 (N_9371,N_9033,N_9222);
nor U9372 (N_9372,N_9138,N_9194);
nor U9373 (N_9373,N_9055,N_9217);
and U9374 (N_9374,N_9008,N_9006);
nand U9375 (N_9375,N_9001,N_9016);
xnor U9376 (N_9376,N_9172,N_9091);
or U9377 (N_9377,N_9175,N_9042);
xnor U9378 (N_9378,N_9008,N_9063);
and U9379 (N_9379,N_9051,N_9097);
nor U9380 (N_9380,N_9103,N_9070);
nand U9381 (N_9381,N_9082,N_9230);
and U9382 (N_9382,N_9192,N_9070);
and U9383 (N_9383,N_9202,N_9208);
nand U9384 (N_9384,N_9184,N_9225);
and U9385 (N_9385,N_9049,N_9141);
nand U9386 (N_9386,N_9081,N_9236);
or U9387 (N_9387,N_9045,N_9224);
and U9388 (N_9388,N_9120,N_9002);
and U9389 (N_9389,N_9215,N_9137);
nor U9390 (N_9390,N_9205,N_9234);
and U9391 (N_9391,N_9001,N_9003);
or U9392 (N_9392,N_9122,N_9058);
nand U9393 (N_9393,N_9186,N_9122);
and U9394 (N_9394,N_9151,N_9054);
nor U9395 (N_9395,N_9095,N_9187);
nor U9396 (N_9396,N_9089,N_9005);
and U9397 (N_9397,N_9173,N_9088);
nand U9398 (N_9398,N_9090,N_9184);
nand U9399 (N_9399,N_9166,N_9146);
or U9400 (N_9400,N_9047,N_9141);
and U9401 (N_9401,N_9081,N_9026);
nand U9402 (N_9402,N_9139,N_9001);
nand U9403 (N_9403,N_9175,N_9126);
and U9404 (N_9404,N_9204,N_9227);
xor U9405 (N_9405,N_9088,N_9177);
or U9406 (N_9406,N_9033,N_9233);
or U9407 (N_9407,N_9219,N_9097);
nor U9408 (N_9408,N_9131,N_9048);
xor U9409 (N_9409,N_9031,N_9123);
nand U9410 (N_9410,N_9172,N_9035);
and U9411 (N_9411,N_9134,N_9085);
or U9412 (N_9412,N_9034,N_9223);
nand U9413 (N_9413,N_9175,N_9142);
nand U9414 (N_9414,N_9095,N_9247);
nor U9415 (N_9415,N_9164,N_9128);
nor U9416 (N_9416,N_9050,N_9039);
nand U9417 (N_9417,N_9060,N_9070);
or U9418 (N_9418,N_9014,N_9237);
nor U9419 (N_9419,N_9068,N_9126);
nand U9420 (N_9420,N_9145,N_9244);
nor U9421 (N_9421,N_9154,N_9083);
or U9422 (N_9422,N_9233,N_9052);
and U9423 (N_9423,N_9061,N_9102);
xnor U9424 (N_9424,N_9015,N_9013);
nor U9425 (N_9425,N_9234,N_9134);
or U9426 (N_9426,N_9159,N_9244);
xor U9427 (N_9427,N_9057,N_9188);
or U9428 (N_9428,N_9076,N_9217);
nand U9429 (N_9429,N_9083,N_9131);
nor U9430 (N_9430,N_9032,N_9057);
and U9431 (N_9431,N_9156,N_9133);
or U9432 (N_9432,N_9170,N_9063);
xnor U9433 (N_9433,N_9112,N_9148);
or U9434 (N_9434,N_9159,N_9190);
nand U9435 (N_9435,N_9173,N_9114);
or U9436 (N_9436,N_9125,N_9118);
nand U9437 (N_9437,N_9006,N_9135);
or U9438 (N_9438,N_9113,N_9247);
nand U9439 (N_9439,N_9099,N_9098);
or U9440 (N_9440,N_9120,N_9071);
or U9441 (N_9441,N_9191,N_9053);
or U9442 (N_9442,N_9112,N_9175);
and U9443 (N_9443,N_9202,N_9077);
nor U9444 (N_9444,N_9206,N_9183);
and U9445 (N_9445,N_9038,N_9124);
or U9446 (N_9446,N_9050,N_9042);
or U9447 (N_9447,N_9161,N_9049);
or U9448 (N_9448,N_9216,N_9154);
nor U9449 (N_9449,N_9151,N_9208);
and U9450 (N_9450,N_9012,N_9073);
or U9451 (N_9451,N_9172,N_9023);
or U9452 (N_9452,N_9121,N_9240);
nand U9453 (N_9453,N_9050,N_9209);
nor U9454 (N_9454,N_9052,N_9058);
xor U9455 (N_9455,N_9166,N_9206);
xor U9456 (N_9456,N_9002,N_9043);
nor U9457 (N_9457,N_9153,N_9209);
or U9458 (N_9458,N_9029,N_9144);
and U9459 (N_9459,N_9106,N_9245);
nand U9460 (N_9460,N_9019,N_9199);
or U9461 (N_9461,N_9012,N_9235);
or U9462 (N_9462,N_9127,N_9169);
or U9463 (N_9463,N_9134,N_9209);
nand U9464 (N_9464,N_9223,N_9167);
xnor U9465 (N_9465,N_9228,N_9205);
xnor U9466 (N_9466,N_9085,N_9092);
nor U9467 (N_9467,N_9133,N_9224);
nor U9468 (N_9468,N_9038,N_9063);
xor U9469 (N_9469,N_9182,N_9026);
nor U9470 (N_9470,N_9231,N_9148);
or U9471 (N_9471,N_9159,N_9084);
nand U9472 (N_9472,N_9051,N_9146);
xnor U9473 (N_9473,N_9141,N_9244);
xnor U9474 (N_9474,N_9222,N_9139);
nor U9475 (N_9475,N_9077,N_9142);
or U9476 (N_9476,N_9047,N_9080);
nor U9477 (N_9477,N_9100,N_9161);
and U9478 (N_9478,N_9173,N_9201);
xnor U9479 (N_9479,N_9036,N_9233);
or U9480 (N_9480,N_9155,N_9094);
xor U9481 (N_9481,N_9169,N_9002);
and U9482 (N_9482,N_9032,N_9042);
xnor U9483 (N_9483,N_9095,N_9057);
xnor U9484 (N_9484,N_9177,N_9012);
or U9485 (N_9485,N_9001,N_9156);
xor U9486 (N_9486,N_9243,N_9110);
or U9487 (N_9487,N_9124,N_9180);
or U9488 (N_9488,N_9064,N_9118);
nand U9489 (N_9489,N_9070,N_9143);
xnor U9490 (N_9490,N_9002,N_9234);
and U9491 (N_9491,N_9171,N_9007);
or U9492 (N_9492,N_9042,N_9141);
xnor U9493 (N_9493,N_9020,N_9144);
nand U9494 (N_9494,N_9048,N_9026);
and U9495 (N_9495,N_9249,N_9094);
or U9496 (N_9496,N_9112,N_9200);
or U9497 (N_9497,N_9132,N_9057);
nand U9498 (N_9498,N_9005,N_9185);
and U9499 (N_9499,N_9070,N_9138);
and U9500 (N_9500,N_9343,N_9486);
nand U9501 (N_9501,N_9275,N_9311);
or U9502 (N_9502,N_9451,N_9359);
nor U9503 (N_9503,N_9378,N_9419);
and U9504 (N_9504,N_9409,N_9297);
nor U9505 (N_9505,N_9340,N_9338);
and U9506 (N_9506,N_9305,N_9326);
or U9507 (N_9507,N_9347,N_9283);
xnor U9508 (N_9508,N_9331,N_9334);
xnor U9509 (N_9509,N_9467,N_9389);
xnor U9510 (N_9510,N_9294,N_9487);
and U9511 (N_9511,N_9375,N_9418);
or U9512 (N_9512,N_9333,N_9397);
nor U9513 (N_9513,N_9479,N_9357);
or U9514 (N_9514,N_9439,N_9404);
and U9515 (N_9515,N_9355,N_9281);
nand U9516 (N_9516,N_9406,N_9282);
xnor U9517 (N_9517,N_9356,N_9427);
or U9518 (N_9518,N_9461,N_9327);
or U9519 (N_9519,N_9412,N_9319);
or U9520 (N_9520,N_9325,N_9335);
nand U9521 (N_9521,N_9434,N_9482);
nor U9522 (N_9522,N_9318,N_9269);
xnor U9523 (N_9523,N_9278,N_9387);
nand U9524 (N_9524,N_9483,N_9377);
or U9525 (N_9525,N_9413,N_9403);
nor U9526 (N_9526,N_9447,N_9370);
nor U9527 (N_9527,N_9432,N_9259);
xnor U9528 (N_9528,N_9456,N_9264);
and U9529 (N_9529,N_9438,N_9251);
nand U9530 (N_9530,N_9381,N_9273);
or U9531 (N_9531,N_9390,N_9298);
and U9532 (N_9532,N_9464,N_9498);
xor U9533 (N_9533,N_9323,N_9256);
nor U9534 (N_9534,N_9488,N_9499);
xor U9535 (N_9535,N_9497,N_9396);
xnor U9536 (N_9536,N_9384,N_9459);
or U9537 (N_9537,N_9443,N_9385);
nor U9538 (N_9538,N_9277,N_9368);
nor U9539 (N_9539,N_9321,N_9457);
nor U9540 (N_9540,N_9288,N_9460);
and U9541 (N_9541,N_9312,N_9324);
nand U9542 (N_9542,N_9369,N_9279);
nand U9543 (N_9543,N_9440,N_9431);
nand U9544 (N_9544,N_9257,N_9358);
nor U9545 (N_9545,N_9280,N_9348);
xor U9546 (N_9546,N_9490,N_9346);
nor U9547 (N_9547,N_9435,N_9437);
xor U9548 (N_9548,N_9265,N_9255);
nor U9549 (N_9549,N_9455,N_9252);
nand U9550 (N_9550,N_9469,N_9337);
nor U9551 (N_9551,N_9442,N_9401);
nor U9552 (N_9552,N_9322,N_9268);
nor U9553 (N_9553,N_9367,N_9405);
nand U9554 (N_9554,N_9393,N_9478);
and U9555 (N_9555,N_9466,N_9417);
xnor U9556 (N_9556,N_9446,N_9339);
or U9557 (N_9557,N_9362,N_9386);
and U9558 (N_9558,N_9448,N_9271);
xnor U9559 (N_9559,N_9481,N_9270);
and U9560 (N_9560,N_9313,N_9424);
nand U9561 (N_9561,N_9302,N_9263);
or U9562 (N_9562,N_9491,N_9329);
nand U9563 (N_9563,N_9472,N_9480);
nor U9564 (N_9564,N_9428,N_9473);
and U9565 (N_9565,N_9361,N_9300);
xor U9566 (N_9566,N_9299,N_9291);
nand U9567 (N_9567,N_9363,N_9304);
nand U9568 (N_9568,N_9272,N_9320);
xnor U9569 (N_9569,N_9344,N_9383);
xnor U9570 (N_9570,N_9414,N_9293);
xnor U9571 (N_9571,N_9258,N_9253);
xor U9572 (N_9572,N_9328,N_9398);
and U9573 (N_9573,N_9317,N_9365);
nor U9574 (N_9574,N_9352,N_9462);
nand U9575 (N_9575,N_9489,N_9426);
nor U9576 (N_9576,N_9441,N_9388);
xnor U9577 (N_9577,N_9394,N_9336);
nor U9578 (N_9578,N_9290,N_9422);
xnor U9579 (N_9579,N_9260,N_9276);
and U9580 (N_9580,N_9463,N_9341);
xnor U9581 (N_9581,N_9354,N_9289);
or U9582 (N_9582,N_9485,N_9250);
nor U9583 (N_9583,N_9303,N_9391);
or U9584 (N_9584,N_9254,N_9342);
nand U9585 (N_9585,N_9444,N_9453);
xor U9586 (N_9586,N_9316,N_9445);
xnor U9587 (N_9587,N_9430,N_9262);
xnor U9588 (N_9588,N_9274,N_9306);
nor U9589 (N_9589,N_9493,N_9425);
and U9590 (N_9590,N_9474,N_9374);
or U9591 (N_9591,N_9471,N_9416);
and U9592 (N_9592,N_9410,N_9392);
and U9593 (N_9593,N_9465,N_9454);
nand U9594 (N_9594,N_9286,N_9420);
and U9595 (N_9595,N_9309,N_9360);
xnor U9596 (N_9596,N_9314,N_9399);
xnor U9597 (N_9597,N_9400,N_9261);
nor U9598 (N_9598,N_9366,N_9433);
nor U9599 (N_9599,N_9468,N_9350);
or U9600 (N_9600,N_9415,N_9476);
nand U9601 (N_9601,N_9429,N_9373);
nand U9602 (N_9602,N_9296,N_9496);
nand U9603 (N_9603,N_9477,N_9411);
and U9604 (N_9604,N_9495,N_9266);
nor U9605 (N_9605,N_9492,N_9372);
or U9606 (N_9606,N_9407,N_9458);
nor U9607 (N_9607,N_9345,N_9452);
xnor U9608 (N_9608,N_9308,N_9287);
and U9609 (N_9609,N_9310,N_9295);
or U9610 (N_9610,N_9353,N_9484);
and U9611 (N_9611,N_9285,N_9267);
or U9612 (N_9612,N_9395,N_9307);
xnor U9613 (N_9613,N_9382,N_9379);
or U9614 (N_9614,N_9371,N_9330);
nand U9615 (N_9615,N_9301,N_9315);
nand U9616 (N_9616,N_9475,N_9364);
or U9617 (N_9617,N_9449,N_9408);
and U9618 (N_9618,N_9376,N_9423);
xnor U9619 (N_9619,N_9494,N_9450);
nor U9620 (N_9620,N_9470,N_9351);
and U9621 (N_9621,N_9436,N_9349);
or U9622 (N_9622,N_9402,N_9421);
nand U9623 (N_9623,N_9380,N_9284);
and U9624 (N_9624,N_9332,N_9292);
and U9625 (N_9625,N_9489,N_9298);
and U9626 (N_9626,N_9336,N_9418);
xnor U9627 (N_9627,N_9276,N_9370);
nand U9628 (N_9628,N_9406,N_9445);
xnor U9629 (N_9629,N_9404,N_9284);
and U9630 (N_9630,N_9365,N_9259);
or U9631 (N_9631,N_9451,N_9392);
nor U9632 (N_9632,N_9480,N_9372);
xor U9633 (N_9633,N_9346,N_9485);
and U9634 (N_9634,N_9275,N_9265);
nor U9635 (N_9635,N_9403,N_9398);
xnor U9636 (N_9636,N_9347,N_9305);
xor U9637 (N_9637,N_9263,N_9319);
nor U9638 (N_9638,N_9274,N_9295);
nand U9639 (N_9639,N_9278,N_9374);
xnor U9640 (N_9640,N_9478,N_9446);
xnor U9641 (N_9641,N_9494,N_9423);
and U9642 (N_9642,N_9302,N_9307);
or U9643 (N_9643,N_9462,N_9479);
and U9644 (N_9644,N_9417,N_9474);
or U9645 (N_9645,N_9349,N_9364);
nor U9646 (N_9646,N_9446,N_9494);
xnor U9647 (N_9647,N_9294,N_9286);
or U9648 (N_9648,N_9439,N_9330);
nor U9649 (N_9649,N_9331,N_9302);
nand U9650 (N_9650,N_9472,N_9336);
or U9651 (N_9651,N_9492,N_9381);
nor U9652 (N_9652,N_9491,N_9436);
or U9653 (N_9653,N_9396,N_9291);
and U9654 (N_9654,N_9473,N_9297);
and U9655 (N_9655,N_9303,N_9491);
nor U9656 (N_9656,N_9428,N_9271);
nand U9657 (N_9657,N_9298,N_9363);
nand U9658 (N_9658,N_9417,N_9253);
and U9659 (N_9659,N_9259,N_9354);
xnor U9660 (N_9660,N_9272,N_9333);
and U9661 (N_9661,N_9459,N_9412);
and U9662 (N_9662,N_9276,N_9445);
xor U9663 (N_9663,N_9339,N_9280);
nor U9664 (N_9664,N_9263,N_9486);
xor U9665 (N_9665,N_9327,N_9463);
xnor U9666 (N_9666,N_9397,N_9469);
and U9667 (N_9667,N_9315,N_9269);
nand U9668 (N_9668,N_9271,N_9282);
and U9669 (N_9669,N_9256,N_9346);
xnor U9670 (N_9670,N_9265,N_9464);
nand U9671 (N_9671,N_9310,N_9301);
nand U9672 (N_9672,N_9254,N_9414);
or U9673 (N_9673,N_9324,N_9436);
nor U9674 (N_9674,N_9453,N_9479);
or U9675 (N_9675,N_9255,N_9344);
or U9676 (N_9676,N_9423,N_9496);
nand U9677 (N_9677,N_9406,N_9455);
and U9678 (N_9678,N_9272,N_9271);
and U9679 (N_9679,N_9447,N_9492);
and U9680 (N_9680,N_9416,N_9469);
nand U9681 (N_9681,N_9399,N_9374);
nand U9682 (N_9682,N_9268,N_9455);
nand U9683 (N_9683,N_9380,N_9321);
nor U9684 (N_9684,N_9317,N_9298);
and U9685 (N_9685,N_9386,N_9342);
nand U9686 (N_9686,N_9486,N_9338);
nand U9687 (N_9687,N_9251,N_9402);
or U9688 (N_9688,N_9468,N_9357);
nor U9689 (N_9689,N_9463,N_9421);
or U9690 (N_9690,N_9336,N_9398);
nor U9691 (N_9691,N_9255,N_9399);
nand U9692 (N_9692,N_9456,N_9411);
xor U9693 (N_9693,N_9476,N_9441);
nor U9694 (N_9694,N_9494,N_9403);
nor U9695 (N_9695,N_9483,N_9440);
or U9696 (N_9696,N_9350,N_9451);
nor U9697 (N_9697,N_9496,N_9394);
and U9698 (N_9698,N_9433,N_9492);
xnor U9699 (N_9699,N_9401,N_9470);
nand U9700 (N_9700,N_9283,N_9481);
and U9701 (N_9701,N_9317,N_9457);
nor U9702 (N_9702,N_9363,N_9324);
and U9703 (N_9703,N_9376,N_9415);
nand U9704 (N_9704,N_9406,N_9402);
xor U9705 (N_9705,N_9251,N_9358);
xor U9706 (N_9706,N_9332,N_9372);
nor U9707 (N_9707,N_9453,N_9422);
or U9708 (N_9708,N_9432,N_9393);
and U9709 (N_9709,N_9441,N_9364);
or U9710 (N_9710,N_9288,N_9396);
or U9711 (N_9711,N_9276,N_9319);
or U9712 (N_9712,N_9474,N_9297);
nand U9713 (N_9713,N_9319,N_9444);
xnor U9714 (N_9714,N_9351,N_9344);
nor U9715 (N_9715,N_9496,N_9410);
nand U9716 (N_9716,N_9421,N_9411);
or U9717 (N_9717,N_9463,N_9367);
and U9718 (N_9718,N_9466,N_9344);
or U9719 (N_9719,N_9340,N_9415);
nand U9720 (N_9720,N_9418,N_9305);
nor U9721 (N_9721,N_9350,N_9341);
nand U9722 (N_9722,N_9488,N_9355);
nand U9723 (N_9723,N_9426,N_9355);
xnor U9724 (N_9724,N_9371,N_9276);
and U9725 (N_9725,N_9397,N_9398);
nor U9726 (N_9726,N_9389,N_9384);
or U9727 (N_9727,N_9259,N_9285);
nor U9728 (N_9728,N_9386,N_9280);
or U9729 (N_9729,N_9289,N_9395);
or U9730 (N_9730,N_9455,N_9320);
nand U9731 (N_9731,N_9370,N_9335);
nand U9732 (N_9732,N_9311,N_9374);
nand U9733 (N_9733,N_9317,N_9431);
or U9734 (N_9734,N_9275,N_9359);
and U9735 (N_9735,N_9276,N_9297);
nor U9736 (N_9736,N_9476,N_9289);
xor U9737 (N_9737,N_9480,N_9462);
or U9738 (N_9738,N_9281,N_9321);
nand U9739 (N_9739,N_9360,N_9434);
nor U9740 (N_9740,N_9422,N_9389);
or U9741 (N_9741,N_9311,N_9409);
xnor U9742 (N_9742,N_9400,N_9273);
nor U9743 (N_9743,N_9473,N_9484);
nand U9744 (N_9744,N_9441,N_9363);
and U9745 (N_9745,N_9325,N_9396);
xnor U9746 (N_9746,N_9357,N_9417);
or U9747 (N_9747,N_9463,N_9411);
nor U9748 (N_9748,N_9255,N_9290);
nand U9749 (N_9749,N_9298,N_9376);
xor U9750 (N_9750,N_9527,N_9583);
nand U9751 (N_9751,N_9544,N_9647);
xnor U9752 (N_9752,N_9520,N_9504);
or U9753 (N_9753,N_9600,N_9556);
or U9754 (N_9754,N_9575,N_9514);
nand U9755 (N_9755,N_9724,N_9743);
or U9756 (N_9756,N_9533,N_9648);
or U9757 (N_9757,N_9566,N_9727);
or U9758 (N_9758,N_9665,N_9693);
nor U9759 (N_9759,N_9578,N_9584);
xor U9760 (N_9760,N_9542,N_9680);
and U9761 (N_9761,N_9684,N_9740);
xor U9762 (N_9762,N_9617,N_9748);
xnor U9763 (N_9763,N_9598,N_9595);
xnor U9764 (N_9764,N_9722,N_9576);
nor U9765 (N_9765,N_9638,N_9601);
or U9766 (N_9766,N_9732,N_9741);
or U9767 (N_9767,N_9700,N_9521);
nor U9768 (N_9768,N_9609,N_9688);
and U9769 (N_9769,N_9505,N_9550);
or U9770 (N_9770,N_9611,N_9634);
xnor U9771 (N_9771,N_9579,N_9667);
and U9772 (N_9772,N_9678,N_9581);
nor U9773 (N_9773,N_9618,N_9517);
nand U9774 (N_9774,N_9559,N_9711);
nand U9775 (N_9775,N_9589,N_9610);
nand U9776 (N_9776,N_9552,N_9586);
nor U9777 (N_9777,N_9535,N_9644);
and U9778 (N_9778,N_9636,N_9744);
and U9779 (N_9779,N_9511,N_9738);
or U9780 (N_9780,N_9500,N_9572);
and U9781 (N_9781,N_9567,N_9608);
and U9782 (N_9782,N_9716,N_9574);
xor U9783 (N_9783,N_9673,N_9605);
and U9784 (N_9784,N_9614,N_9737);
xor U9785 (N_9785,N_9561,N_9540);
and U9786 (N_9786,N_9590,N_9626);
xnor U9787 (N_9787,N_9606,N_9512);
nor U9788 (N_9788,N_9645,N_9670);
nand U9789 (N_9789,N_9705,N_9747);
nand U9790 (N_9790,N_9591,N_9739);
xor U9791 (N_9791,N_9526,N_9503);
and U9792 (N_9792,N_9532,N_9646);
xnor U9793 (N_9793,N_9719,N_9546);
and U9794 (N_9794,N_9588,N_9686);
nor U9795 (N_9795,N_9523,N_9676);
nor U9796 (N_9796,N_9721,N_9694);
xor U9797 (N_9797,N_9674,N_9704);
nor U9798 (N_9798,N_9687,N_9742);
nand U9799 (N_9799,N_9663,N_9649);
or U9800 (N_9800,N_9720,N_9725);
xnor U9801 (N_9801,N_9616,N_9539);
or U9802 (N_9802,N_9513,N_9525);
or U9803 (N_9803,N_9713,N_9690);
or U9804 (N_9804,N_9675,N_9746);
or U9805 (N_9805,N_9615,N_9656);
nor U9806 (N_9806,N_9712,N_9660);
xnor U9807 (N_9807,N_9631,N_9554);
nor U9808 (N_9808,N_9730,N_9652);
and U9809 (N_9809,N_9695,N_9549);
nand U9810 (N_9810,N_9571,N_9507);
xor U9811 (N_9811,N_9502,N_9585);
nand U9812 (N_9812,N_9735,N_9710);
or U9813 (N_9813,N_9594,N_9662);
nor U9814 (N_9814,N_9717,N_9622);
nor U9815 (N_9815,N_9661,N_9592);
or U9816 (N_9816,N_9632,N_9613);
nand U9817 (N_9817,N_9515,N_9602);
nand U9818 (N_9818,N_9596,N_9733);
nor U9819 (N_9819,N_9570,N_9536);
nand U9820 (N_9820,N_9573,N_9545);
nor U9821 (N_9821,N_9708,N_9619);
nor U9822 (N_9822,N_9692,N_9519);
nand U9823 (N_9823,N_9541,N_9707);
xnor U9824 (N_9824,N_9577,N_9629);
or U9825 (N_9825,N_9709,N_9604);
xnor U9826 (N_9826,N_9553,N_9657);
nand U9827 (N_9827,N_9637,N_9564);
xor U9828 (N_9828,N_9557,N_9669);
nand U9829 (N_9829,N_9640,N_9518);
nand U9830 (N_9830,N_9558,N_9734);
nand U9831 (N_9831,N_9714,N_9728);
and U9832 (N_9832,N_9666,N_9551);
xnor U9833 (N_9833,N_9715,N_9718);
and U9834 (N_9834,N_9587,N_9563);
nand U9835 (N_9835,N_9677,N_9701);
nor U9836 (N_9836,N_9562,N_9508);
nand U9837 (N_9837,N_9664,N_9597);
or U9838 (N_9838,N_9582,N_9706);
and U9839 (N_9839,N_9547,N_9599);
nand U9840 (N_9840,N_9543,N_9703);
or U9841 (N_9841,N_9528,N_9555);
nand U9842 (N_9842,N_9623,N_9650);
and U9843 (N_9843,N_9659,N_9537);
nor U9844 (N_9844,N_9699,N_9723);
or U9845 (N_9845,N_9627,N_9625);
nor U9846 (N_9846,N_9509,N_9529);
nand U9847 (N_9847,N_9593,N_9522);
or U9848 (N_9848,N_9681,N_9569);
and U9849 (N_9849,N_9643,N_9538);
nand U9850 (N_9850,N_9603,N_9736);
or U9851 (N_9851,N_9726,N_9516);
and U9852 (N_9852,N_9531,N_9729);
or U9853 (N_9853,N_9696,N_9682);
and U9854 (N_9854,N_9691,N_9560);
nor U9855 (N_9855,N_9683,N_9565);
and U9856 (N_9856,N_9568,N_9658);
or U9857 (N_9857,N_9641,N_9628);
and U9858 (N_9858,N_9530,N_9689);
and U9859 (N_9859,N_9501,N_9697);
and U9860 (N_9860,N_9607,N_9653);
xnor U9861 (N_9861,N_9655,N_9642);
and U9862 (N_9862,N_9698,N_9668);
nor U9863 (N_9863,N_9749,N_9651);
nand U9864 (N_9864,N_9624,N_9534);
or U9865 (N_9865,N_9639,N_9524);
and U9866 (N_9866,N_9702,N_9672);
or U9867 (N_9867,N_9745,N_9612);
or U9868 (N_9868,N_9510,N_9685);
nor U9869 (N_9869,N_9633,N_9671);
xnor U9870 (N_9870,N_9621,N_9630);
nor U9871 (N_9871,N_9679,N_9580);
nor U9872 (N_9872,N_9635,N_9654);
nor U9873 (N_9873,N_9620,N_9506);
xnor U9874 (N_9874,N_9731,N_9548);
or U9875 (N_9875,N_9683,N_9625);
and U9876 (N_9876,N_9670,N_9727);
and U9877 (N_9877,N_9545,N_9547);
nor U9878 (N_9878,N_9504,N_9612);
nor U9879 (N_9879,N_9533,N_9643);
or U9880 (N_9880,N_9576,N_9643);
nand U9881 (N_9881,N_9624,N_9667);
nand U9882 (N_9882,N_9739,N_9743);
and U9883 (N_9883,N_9705,N_9635);
and U9884 (N_9884,N_9579,N_9586);
xor U9885 (N_9885,N_9739,N_9737);
xnor U9886 (N_9886,N_9747,N_9693);
xor U9887 (N_9887,N_9504,N_9666);
and U9888 (N_9888,N_9533,N_9507);
xnor U9889 (N_9889,N_9500,N_9734);
xor U9890 (N_9890,N_9551,N_9657);
nand U9891 (N_9891,N_9572,N_9581);
and U9892 (N_9892,N_9535,N_9627);
nor U9893 (N_9893,N_9668,N_9510);
or U9894 (N_9894,N_9514,N_9685);
and U9895 (N_9895,N_9520,N_9595);
nand U9896 (N_9896,N_9675,N_9726);
nor U9897 (N_9897,N_9619,N_9729);
nor U9898 (N_9898,N_9618,N_9690);
nand U9899 (N_9899,N_9555,N_9744);
or U9900 (N_9900,N_9721,N_9708);
or U9901 (N_9901,N_9570,N_9566);
or U9902 (N_9902,N_9655,N_9583);
nor U9903 (N_9903,N_9591,N_9634);
nand U9904 (N_9904,N_9640,N_9742);
or U9905 (N_9905,N_9549,N_9521);
and U9906 (N_9906,N_9607,N_9516);
xor U9907 (N_9907,N_9692,N_9605);
nand U9908 (N_9908,N_9657,N_9736);
or U9909 (N_9909,N_9629,N_9585);
and U9910 (N_9910,N_9630,N_9613);
nand U9911 (N_9911,N_9532,N_9642);
and U9912 (N_9912,N_9667,N_9730);
nand U9913 (N_9913,N_9522,N_9612);
xor U9914 (N_9914,N_9726,N_9534);
nand U9915 (N_9915,N_9667,N_9746);
and U9916 (N_9916,N_9690,N_9519);
or U9917 (N_9917,N_9659,N_9555);
nand U9918 (N_9918,N_9511,N_9621);
or U9919 (N_9919,N_9594,N_9681);
nand U9920 (N_9920,N_9704,N_9633);
or U9921 (N_9921,N_9671,N_9704);
and U9922 (N_9922,N_9680,N_9586);
nand U9923 (N_9923,N_9521,N_9627);
and U9924 (N_9924,N_9600,N_9641);
and U9925 (N_9925,N_9514,N_9601);
xor U9926 (N_9926,N_9546,N_9572);
or U9927 (N_9927,N_9521,N_9708);
xor U9928 (N_9928,N_9612,N_9556);
nor U9929 (N_9929,N_9699,N_9709);
and U9930 (N_9930,N_9590,N_9724);
and U9931 (N_9931,N_9619,N_9646);
or U9932 (N_9932,N_9591,N_9633);
and U9933 (N_9933,N_9685,N_9649);
and U9934 (N_9934,N_9671,N_9718);
nor U9935 (N_9935,N_9536,N_9648);
or U9936 (N_9936,N_9697,N_9564);
xnor U9937 (N_9937,N_9628,N_9724);
or U9938 (N_9938,N_9641,N_9726);
and U9939 (N_9939,N_9506,N_9539);
nand U9940 (N_9940,N_9660,N_9692);
or U9941 (N_9941,N_9525,N_9610);
and U9942 (N_9942,N_9586,N_9716);
and U9943 (N_9943,N_9570,N_9539);
or U9944 (N_9944,N_9613,N_9648);
and U9945 (N_9945,N_9563,N_9679);
nor U9946 (N_9946,N_9563,N_9662);
nor U9947 (N_9947,N_9720,N_9675);
and U9948 (N_9948,N_9580,N_9554);
or U9949 (N_9949,N_9706,N_9724);
xnor U9950 (N_9950,N_9665,N_9688);
and U9951 (N_9951,N_9729,N_9608);
xor U9952 (N_9952,N_9666,N_9512);
nor U9953 (N_9953,N_9741,N_9547);
or U9954 (N_9954,N_9664,N_9619);
xor U9955 (N_9955,N_9566,N_9651);
xor U9956 (N_9956,N_9589,N_9591);
nor U9957 (N_9957,N_9674,N_9550);
xnor U9958 (N_9958,N_9591,N_9644);
or U9959 (N_9959,N_9534,N_9685);
nand U9960 (N_9960,N_9587,N_9680);
nand U9961 (N_9961,N_9517,N_9599);
nand U9962 (N_9962,N_9628,N_9531);
or U9963 (N_9963,N_9703,N_9536);
and U9964 (N_9964,N_9652,N_9700);
nor U9965 (N_9965,N_9520,N_9635);
xor U9966 (N_9966,N_9678,N_9638);
or U9967 (N_9967,N_9695,N_9654);
or U9968 (N_9968,N_9682,N_9541);
nor U9969 (N_9969,N_9574,N_9689);
or U9970 (N_9970,N_9657,N_9731);
nor U9971 (N_9971,N_9513,N_9548);
and U9972 (N_9972,N_9745,N_9701);
and U9973 (N_9973,N_9572,N_9706);
nand U9974 (N_9974,N_9629,N_9723);
nor U9975 (N_9975,N_9727,N_9610);
xor U9976 (N_9976,N_9592,N_9707);
and U9977 (N_9977,N_9735,N_9670);
and U9978 (N_9978,N_9576,N_9618);
and U9979 (N_9979,N_9720,N_9577);
nor U9980 (N_9980,N_9576,N_9526);
xor U9981 (N_9981,N_9595,N_9732);
nor U9982 (N_9982,N_9537,N_9516);
nand U9983 (N_9983,N_9513,N_9538);
or U9984 (N_9984,N_9658,N_9738);
or U9985 (N_9985,N_9657,N_9584);
and U9986 (N_9986,N_9697,N_9694);
nand U9987 (N_9987,N_9701,N_9541);
nand U9988 (N_9988,N_9683,N_9736);
nand U9989 (N_9989,N_9671,N_9639);
nand U9990 (N_9990,N_9733,N_9529);
xnor U9991 (N_9991,N_9551,N_9685);
xnor U9992 (N_9992,N_9532,N_9565);
xor U9993 (N_9993,N_9520,N_9573);
nand U9994 (N_9994,N_9628,N_9529);
or U9995 (N_9995,N_9670,N_9597);
xnor U9996 (N_9996,N_9546,N_9700);
xnor U9997 (N_9997,N_9676,N_9703);
xnor U9998 (N_9998,N_9593,N_9544);
and U9999 (N_9999,N_9563,N_9617);
or U10000 (N_10000,N_9831,N_9975);
xor U10001 (N_10001,N_9867,N_9878);
or U10002 (N_10002,N_9846,N_9929);
nor U10003 (N_10003,N_9790,N_9838);
xnor U10004 (N_10004,N_9821,N_9999);
nand U10005 (N_10005,N_9912,N_9839);
or U10006 (N_10006,N_9882,N_9970);
nor U10007 (N_10007,N_9927,N_9766);
or U10008 (N_10008,N_9916,N_9818);
nor U10009 (N_10009,N_9907,N_9752);
xor U10010 (N_10010,N_9777,N_9813);
or U10011 (N_10011,N_9981,N_9926);
nand U10012 (N_10012,N_9875,N_9759);
and U10013 (N_10013,N_9978,N_9842);
and U10014 (N_10014,N_9967,N_9773);
nor U10015 (N_10015,N_9765,N_9778);
or U10016 (N_10016,N_9788,N_9898);
nor U10017 (N_10017,N_9872,N_9850);
xnor U10018 (N_10018,N_9866,N_9883);
and U10019 (N_10019,N_9841,N_9923);
xor U10020 (N_10020,N_9902,N_9990);
or U10021 (N_10021,N_9946,N_9901);
and U10022 (N_10022,N_9993,N_9801);
xnor U10023 (N_10023,N_9936,N_9855);
nand U10024 (N_10024,N_9822,N_9787);
and U10025 (N_10025,N_9824,N_9772);
nand U10026 (N_10026,N_9976,N_9940);
or U10027 (N_10027,N_9789,N_9931);
nand U10028 (N_10028,N_9953,N_9964);
or U10029 (N_10029,N_9886,N_9969);
and U10030 (N_10030,N_9819,N_9827);
nand U10031 (N_10031,N_9933,N_9844);
xnor U10032 (N_10032,N_9982,N_9817);
nand U10033 (N_10033,N_9753,N_9919);
or U10034 (N_10034,N_9979,N_9899);
or U10035 (N_10035,N_9816,N_9986);
xnor U10036 (N_10036,N_9770,N_9750);
or U10037 (N_10037,N_9767,N_9891);
and U10038 (N_10038,N_9915,N_9843);
and U10039 (N_10039,N_9998,N_9992);
xnor U10040 (N_10040,N_9961,N_9851);
nand U10041 (N_10041,N_9894,N_9892);
and U10042 (N_10042,N_9868,N_9852);
nand U10043 (N_10043,N_9779,N_9879);
and U10044 (N_10044,N_9974,N_9954);
nor U10045 (N_10045,N_9939,N_9870);
nor U10046 (N_10046,N_9896,N_9857);
nor U10047 (N_10047,N_9861,N_9823);
xnor U10048 (N_10048,N_9792,N_9871);
nand U10049 (N_10049,N_9905,N_9985);
and U10050 (N_10050,N_9854,N_9924);
nand U10051 (N_10051,N_9925,N_9786);
xor U10052 (N_10052,N_9781,N_9965);
and U10053 (N_10053,N_9888,N_9780);
or U10054 (N_10054,N_9890,N_9908);
or U10055 (N_10055,N_9906,N_9984);
and U10056 (N_10056,N_9805,N_9917);
nand U10057 (N_10057,N_9859,N_9795);
xnor U10058 (N_10058,N_9885,N_9847);
nor U10059 (N_10059,N_9904,N_9849);
nor U10060 (N_10060,N_9913,N_9944);
xnor U10061 (N_10061,N_9811,N_9865);
xor U10062 (N_10062,N_9881,N_9968);
and U10063 (N_10063,N_9793,N_9895);
and U10064 (N_10064,N_9810,N_9791);
nand U10065 (N_10065,N_9832,N_9803);
and U10066 (N_10066,N_9941,N_9966);
or U10067 (N_10067,N_9764,N_9932);
nor U10068 (N_10068,N_9799,N_9897);
nor U10069 (N_10069,N_9952,N_9948);
xnor U10070 (N_10070,N_9755,N_9834);
and U10071 (N_10071,N_9774,N_9930);
nand U10072 (N_10072,N_9880,N_9958);
and U10073 (N_10073,N_9971,N_9806);
nand U10074 (N_10074,N_9826,N_9949);
and U10075 (N_10075,N_9768,N_9874);
and U10076 (N_10076,N_9889,N_9771);
xnor U10077 (N_10077,N_9956,N_9783);
nand U10078 (N_10078,N_9876,N_9922);
or U10079 (N_10079,N_9973,N_9853);
nor U10080 (N_10080,N_9960,N_9836);
nand U10081 (N_10081,N_9942,N_9815);
nor U10082 (N_10082,N_9785,N_9959);
nand U10083 (N_10083,N_9950,N_9873);
nand U10084 (N_10084,N_9845,N_9807);
xnor U10085 (N_10085,N_9918,N_9921);
or U10086 (N_10086,N_9935,N_9928);
or U10087 (N_10087,N_9763,N_9760);
nor U10088 (N_10088,N_9962,N_9893);
nand U10089 (N_10089,N_9863,N_9911);
or U10090 (N_10090,N_9784,N_9754);
or U10091 (N_10091,N_9937,N_9947);
nand U10092 (N_10092,N_9812,N_9858);
xor U10093 (N_10093,N_9996,N_9989);
and U10094 (N_10094,N_9856,N_9814);
xnor U10095 (N_10095,N_9945,N_9980);
and U10096 (N_10096,N_9769,N_9910);
and U10097 (N_10097,N_9884,N_9914);
xor U10098 (N_10098,N_9994,N_9758);
xor U10099 (N_10099,N_9951,N_9782);
or U10100 (N_10100,N_9808,N_9820);
nand U10101 (N_10101,N_9751,N_9835);
or U10102 (N_10102,N_9848,N_9862);
xor U10103 (N_10103,N_9798,N_9830);
or U10104 (N_10104,N_9869,N_9900);
or U10105 (N_10105,N_9909,N_9833);
nor U10106 (N_10106,N_9762,N_9804);
xor U10107 (N_10107,N_9776,N_9938);
or U10108 (N_10108,N_9864,N_9987);
xor U10109 (N_10109,N_9756,N_9963);
and U10110 (N_10110,N_9797,N_9903);
nand U10111 (N_10111,N_9991,N_9934);
nand U10112 (N_10112,N_9995,N_9829);
or U10113 (N_10113,N_9825,N_9997);
and U10114 (N_10114,N_9757,N_9775);
or U10115 (N_10115,N_9860,N_9977);
nor U10116 (N_10116,N_9809,N_9943);
nand U10117 (N_10117,N_9840,N_9800);
nor U10118 (N_10118,N_9983,N_9802);
xor U10119 (N_10119,N_9955,N_9837);
nor U10120 (N_10120,N_9920,N_9761);
xor U10121 (N_10121,N_9887,N_9877);
nor U10122 (N_10122,N_9828,N_9957);
or U10123 (N_10123,N_9988,N_9794);
and U10124 (N_10124,N_9972,N_9796);
or U10125 (N_10125,N_9935,N_9797);
nand U10126 (N_10126,N_9918,N_9849);
or U10127 (N_10127,N_9844,N_9768);
nand U10128 (N_10128,N_9982,N_9804);
and U10129 (N_10129,N_9975,N_9794);
nor U10130 (N_10130,N_9857,N_9815);
nor U10131 (N_10131,N_9877,N_9905);
and U10132 (N_10132,N_9752,N_9998);
nand U10133 (N_10133,N_9858,N_9919);
nor U10134 (N_10134,N_9826,N_9924);
and U10135 (N_10135,N_9813,N_9920);
nor U10136 (N_10136,N_9751,N_9957);
nand U10137 (N_10137,N_9985,N_9920);
and U10138 (N_10138,N_9793,N_9854);
nand U10139 (N_10139,N_9907,N_9836);
xor U10140 (N_10140,N_9836,N_9942);
nand U10141 (N_10141,N_9796,N_9805);
or U10142 (N_10142,N_9757,N_9867);
and U10143 (N_10143,N_9971,N_9911);
and U10144 (N_10144,N_9826,N_9881);
or U10145 (N_10145,N_9853,N_9773);
nand U10146 (N_10146,N_9926,N_9956);
xnor U10147 (N_10147,N_9975,N_9962);
nor U10148 (N_10148,N_9810,N_9899);
xor U10149 (N_10149,N_9975,N_9988);
and U10150 (N_10150,N_9971,N_9932);
xnor U10151 (N_10151,N_9931,N_9968);
or U10152 (N_10152,N_9892,N_9923);
and U10153 (N_10153,N_9946,N_9829);
xor U10154 (N_10154,N_9957,N_9750);
nand U10155 (N_10155,N_9953,N_9877);
xnor U10156 (N_10156,N_9861,N_9778);
nor U10157 (N_10157,N_9796,N_9870);
nand U10158 (N_10158,N_9896,N_9916);
and U10159 (N_10159,N_9830,N_9819);
nand U10160 (N_10160,N_9872,N_9833);
nor U10161 (N_10161,N_9972,N_9752);
xnor U10162 (N_10162,N_9754,N_9952);
nand U10163 (N_10163,N_9750,N_9982);
and U10164 (N_10164,N_9818,N_9852);
nand U10165 (N_10165,N_9884,N_9890);
nor U10166 (N_10166,N_9889,N_9900);
xnor U10167 (N_10167,N_9756,N_9914);
nor U10168 (N_10168,N_9801,N_9936);
nor U10169 (N_10169,N_9952,N_9978);
nor U10170 (N_10170,N_9782,N_9750);
nand U10171 (N_10171,N_9818,N_9802);
xnor U10172 (N_10172,N_9765,N_9923);
xor U10173 (N_10173,N_9994,N_9862);
xor U10174 (N_10174,N_9951,N_9852);
nand U10175 (N_10175,N_9835,N_9929);
or U10176 (N_10176,N_9885,N_9835);
nor U10177 (N_10177,N_9770,N_9882);
or U10178 (N_10178,N_9819,N_9982);
nand U10179 (N_10179,N_9904,N_9913);
xor U10180 (N_10180,N_9873,N_9991);
or U10181 (N_10181,N_9914,N_9853);
or U10182 (N_10182,N_9776,N_9914);
xnor U10183 (N_10183,N_9812,N_9900);
nor U10184 (N_10184,N_9910,N_9974);
or U10185 (N_10185,N_9985,N_9799);
nor U10186 (N_10186,N_9869,N_9996);
and U10187 (N_10187,N_9965,N_9865);
nand U10188 (N_10188,N_9758,N_9971);
and U10189 (N_10189,N_9830,N_9791);
or U10190 (N_10190,N_9808,N_9869);
nand U10191 (N_10191,N_9795,N_9776);
or U10192 (N_10192,N_9860,N_9797);
nand U10193 (N_10193,N_9955,N_9927);
xnor U10194 (N_10194,N_9902,N_9872);
and U10195 (N_10195,N_9983,N_9957);
nand U10196 (N_10196,N_9775,N_9967);
xor U10197 (N_10197,N_9794,N_9770);
or U10198 (N_10198,N_9985,N_9756);
xnor U10199 (N_10199,N_9848,N_9918);
nor U10200 (N_10200,N_9755,N_9842);
nor U10201 (N_10201,N_9971,N_9819);
nand U10202 (N_10202,N_9940,N_9754);
or U10203 (N_10203,N_9798,N_9945);
or U10204 (N_10204,N_9912,N_9978);
xor U10205 (N_10205,N_9922,N_9837);
or U10206 (N_10206,N_9998,N_9990);
xor U10207 (N_10207,N_9781,N_9830);
nand U10208 (N_10208,N_9822,N_9988);
or U10209 (N_10209,N_9936,N_9784);
or U10210 (N_10210,N_9930,N_9992);
nor U10211 (N_10211,N_9818,N_9795);
xnor U10212 (N_10212,N_9813,N_9788);
nor U10213 (N_10213,N_9882,N_9991);
xnor U10214 (N_10214,N_9951,N_9776);
xnor U10215 (N_10215,N_9925,N_9754);
xnor U10216 (N_10216,N_9800,N_9896);
xnor U10217 (N_10217,N_9900,N_9930);
nor U10218 (N_10218,N_9954,N_9825);
nand U10219 (N_10219,N_9997,N_9911);
and U10220 (N_10220,N_9930,N_9805);
nor U10221 (N_10221,N_9885,N_9925);
nand U10222 (N_10222,N_9785,N_9881);
xnor U10223 (N_10223,N_9767,N_9988);
nor U10224 (N_10224,N_9926,N_9953);
nor U10225 (N_10225,N_9790,N_9788);
xor U10226 (N_10226,N_9809,N_9823);
nor U10227 (N_10227,N_9859,N_9929);
nor U10228 (N_10228,N_9838,N_9880);
or U10229 (N_10229,N_9987,N_9753);
or U10230 (N_10230,N_9852,N_9890);
and U10231 (N_10231,N_9797,N_9915);
or U10232 (N_10232,N_9759,N_9770);
nor U10233 (N_10233,N_9762,N_9944);
or U10234 (N_10234,N_9927,N_9846);
xor U10235 (N_10235,N_9766,N_9940);
or U10236 (N_10236,N_9919,N_9771);
xor U10237 (N_10237,N_9982,N_9910);
xor U10238 (N_10238,N_9959,N_9898);
and U10239 (N_10239,N_9917,N_9782);
or U10240 (N_10240,N_9800,N_9768);
xor U10241 (N_10241,N_9937,N_9806);
nor U10242 (N_10242,N_9820,N_9890);
xor U10243 (N_10243,N_9882,N_9795);
or U10244 (N_10244,N_9758,N_9841);
nor U10245 (N_10245,N_9987,N_9807);
nor U10246 (N_10246,N_9960,N_9892);
or U10247 (N_10247,N_9878,N_9950);
nand U10248 (N_10248,N_9929,N_9799);
nand U10249 (N_10249,N_9987,N_9940);
xor U10250 (N_10250,N_10131,N_10031);
nand U10251 (N_10251,N_10152,N_10042);
nor U10252 (N_10252,N_10230,N_10187);
xnor U10253 (N_10253,N_10147,N_10166);
nor U10254 (N_10254,N_10245,N_10008);
xnor U10255 (N_10255,N_10025,N_10141);
xnor U10256 (N_10256,N_10097,N_10045);
nor U10257 (N_10257,N_10027,N_10159);
xor U10258 (N_10258,N_10011,N_10148);
and U10259 (N_10259,N_10144,N_10209);
or U10260 (N_10260,N_10110,N_10091);
xnor U10261 (N_10261,N_10009,N_10063);
nand U10262 (N_10262,N_10158,N_10219);
nand U10263 (N_10263,N_10059,N_10107);
and U10264 (N_10264,N_10122,N_10016);
nor U10265 (N_10265,N_10015,N_10229);
or U10266 (N_10266,N_10129,N_10193);
or U10267 (N_10267,N_10167,N_10086);
nor U10268 (N_10268,N_10202,N_10056);
nor U10269 (N_10269,N_10084,N_10127);
and U10270 (N_10270,N_10010,N_10217);
or U10271 (N_10271,N_10249,N_10115);
or U10272 (N_10272,N_10154,N_10182);
nand U10273 (N_10273,N_10036,N_10197);
nand U10274 (N_10274,N_10043,N_10001);
nand U10275 (N_10275,N_10236,N_10006);
nor U10276 (N_10276,N_10005,N_10113);
and U10277 (N_10277,N_10248,N_10096);
xnor U10278 (N_10278,N_10116,N_10003);
nand U10279 (N_10279,N_10174,N_10157);
nand U10280 (N_10280,N_10239,N_10076);
xor U10281 (N_10281,N_10169,N_10026);
and U10282 (N_10282,N_10156,N_10223);
xor U10283 (N_10283,N_10083,N_10004);
or U10284 (N_10284,N_10028,N_10051);
xnor U10285 (N_10285,N_10205,N_10178);
and U10286 (N_10286,N_10067,N_10186);
or U10287 (N_10287,N_10049,N_10139);
or U10288 (N_10288,N_10188,N_10022);
and U10289 (N_10289,N_10071,N_10165);
nand U10290 (N_10290,N_10247,N_10093);
or U10291 (N_10291,N_10125,N_10023);
nor U10292 (N_10292,N_10055,N_10181);
or U10293 (N_10293,N_10094,N_10092);
or U10294 (N_10294,N_10200,N_10149);
or U10295 (N_10295,N_10037,N_10231);
xnor U10296 (N_10296,N_10198,N_10013);
xor U10297 (N_10297,N_10109,N_10073);
and U10298 (N_10298,N_10102,N_10064);
or U10299 (N_10299,N_10095,N_10044);
or U10300 (N_10300,N_10021,N_10069);
or U10301 (N_10301,N_10104,N_10201);
nand U10302 (N_10302,N_10054,N_10119);
or U10303 (N_10303,N_10007,N_10194);
nand U10304 (N_10304,N_10032,N_10243);
or U10305 (N_10305,N_10020,N_10216);
xnor U10306 (N_10306,N_10053,N_10244);
or U10307 (N_10307,N_10241,N_10087);
or U10308 (N_10308,N_10014,N_10208);
nand U10309 (N_10309,N_10121,N_10210);
nor U10310 (N_10310,N_10117,N_10111);
nand U10311 (N_10311,N_10101,N_10126);
or U10312 (N_10312,N_10046,N_10103);
and U10313 (N_10313,N_10146,N_10153);
nand U10314 (N_10314,N_10089,N_10114);
xor U10315 (N_10315,N_10047,N_10235);
and U10316 (N_10316,N_10143,N_10150);
or U10317 (N_10317,N_10177,N_10088);
nand U10318 (N_10318,N_10163,N_10124);
and U10319 (N_10319,N_10134,N_10228);
nand U10320 (N_10320,N_10171,N_10220);
or U10321 (N_10321,N_10048,N_10242);
xnor U10322 (N_10322,N_10078,N_10211);
or U10323 (N_10323,N_10214,N_10072);
nand U10324 (N_10324,N_10128,N_10140);
nand U10325 (N_10325,N_10176,N_10195);
nor U10326 (N_10326,N_10218,N_10075);
or U10327 (N_10327,N_10120,N_10070);
and U10328 (N_10328,N_10168,N_10038);
and U10329 (N_10329,N_10029,N_10246);
xnor U10330 (N_10330,N_10172,N_10196);
xnor U10331 (N_10331,N_10033,N_10002);
and U10332 (N_10332,N_10066,N_10137);
nor U10333 (N_10333,N_10138,N_10068);
nor U10334 (N_10334,N_10173,N_10155);
xnor U10335 (N_10335,N_10151,N_10175);
nand U10336 (N_10336,N_10082,N_10133);
and U10337 (N_10337,N_10238,N_10224);
xor U10338 (N_10338,N_10052,N_10040);
nor U10339 (N_10339,N_10012,N_10185);
or U10340 (N_10340,N_10061,N_10112);
and U10341 (N_10341,N_10203,N_10184);
and U10342 (N_10342,N_10034,N_10060);
xor U10343 (N_10343,N_10018,N_10019);
xnor U10344 (N_10344,N_10190,N_10135);
nand U10345 (N_10345,N_10118,N_10160);
nor U10346 (N_10346,N_10179,N_10130);
xor U10347 (N_10347,N_10183,N_10161);
nand U10348 (N_10348,N_10050,N_10199);
or U10349 (N_10349,N_10024,N_10080);
or U10350 (N_10350,N_10145,N_10212);
nor U10351 (N_10351,N_10105,N_10098);
xnor U10352 (N_10352,N_10221,N_10132);
nor U10353 (N_10353,N_10233,N_10108);
and U10354 (N_10354,N_10017,N_10035);
or U10355 (N_10355,N_10232,N_10227);
xor U10356 (N_10356,N_10237,N_10090);
nand U10357 (N_10357,N_10136,N_10062);
xnor U10358 (N_10358,N_10204,N_10081);
xnor U10359 (N_10359,N_10191,N_10039);
and U10360 (N_10360,N_10074,N_10041);
nand U10361 (N_10361,N_10085,N_10225);
xnor U10362 (N_10362,N_10030,N_10162);
xnor U10363 (N_10363,N_10058,N_10142);
nand U10364 (N_10364,N_10180,N_10240);
or U10365 (N_10365,N_10192,N_10079);
nand U10366 (N_10366,N_10222,N_10106);
or U10367 (N_10367,N_10123,N_10170);
nand U10368 (N_10368,N_10213,N_10057);
or U10369 (N_10369,N_10065,N_10077);
nor U10370 (N_10370,N_10000,N_10206);
nor U10371 (N_10371,N_10226,N_10099);
nand U10372 (N_10372,N_10164,N_10189);
and U10373 (N_10373,N_10207,N_10234);
nand U10374 (N_10374,N_10100,N_10215);
nor U10375 (N_10375,N_10053,N_10184);
nor U10376 (N_10376,N_10095,N_10058);
and U10377 (N_10377,N_10052,N_10229);
or U10378 (N_10378,N_10132,N_10196);
nand U10379 (N_10379,N_10128,N_10088);
xor U10380 (N_10380,N_10119,N_10039);
xnor U10381 (N_10381,N_10037,N_10221);
nand U10382 (N_10382,N_10235,N_10175);
nand U10383 (N_10383,N_10236,N_10024);
or U10384 (N_10384,N_10108,N_10137);
or U10385 (N_10385,N_10218,N_10186);
and U10386 (N_10386,N_10219,N_10040);
nand U10387 (N_10387,N_10182,N_10078);
nand U10388 (N_10388,N_10168,N_10036);
or U10389 (N_10389,N_10191,N_10073);
nor U10390 (N_10390,N_10209,N_10084);
and U10391 (N_10391,N_10107,N_10204);
nand U10392 (N_10392,N_10000,N_10234);
xnor U10393 (N_10393,N_10020,N_10078);
or U10394 (N_10394,N_10223,N_10021);
or U10395 (N_10395,N_10181,N_10173);
xor U10396 (N_10396,N_10143,N_10196);
or U10397 (N_10397,N_10042,N_10044);
or U10398 (N_10398,N_10158,N_10094);
and U10399 (N_10399,N_10123,N_10039);
nand U10400 (N_10400,N_10125,N_10205);
xnor U10401 (N_10401,N_10233,N_10044);
nor U10402 (N_10402,N_10133,N_10010);
or U10403 (N_10403,N_10158,N_10106);
nor U10404 (N_10404,N_10243,N_10079);
and U10405 (N_10405,N_10122,N_10039);
and U10406 (N_10406,N_10044,N_10049);
or U10407 (N_10407,N_10027,N_10152);
or U10408 (N_10408,N_10199,N_10033);
nor U10409 (N_10409,N_10139,N_10209);
nor U10410 (N_10410,N_10157,N_10219);
or U10411 (N_10411,N_10080,N_10167);
or U10412 (N_10412,N_10092,N_10139);
and U10413 (N_10413,N_10101,N_10231);
xnor U10414 (N_10414,N_10214,N_10048);
or U10415 (N_10415,N_10107,N_10033);
xnor U10416 (N_10416,N_10138,N_10150);
nand U10417 (N_10417,N_10226,N_10171);
and U10418 (N_10418,N_10207,N_10236);
nor U10419 (N_10419,N_10166,N_10070);
nand U10420 (N_10420,N_10076,N_10091);
xnor U10421 (N_10421,N_10159,N_10021);
nand U10422 (N_10422,N_10096,N_10053);
or U10423 (N_10423,N_10144,N_10152);
xor U10424 (N_10424,N_10229,N_10140);
xor U10425 (N_10425,N_10146,N_10178);
or U10426 (N_10426,N_10206,N_10096);
xnor U10427 (N_10427,N_10147,N_10182);
nor U10428 (N_10428,N_10050,N_10168);
xor U10429 (N_10429,N_10241,N_10063);
xnor U10430 (N_10430,N_10187,N_10025);
xnor U10431 (N_10431,N_10242,N_10212);
and U10432 (N_10432,N_10139,N_10046);
xnor U10433 (N_10433,N_10130,N_10239);
nand U10434 (N_10434,N_10159,N_10017);
or U10435 (N_10435,N_10011,N_10039);
and U10436 (N_10436,N_10107,N_10111);
nand U10437 (N_10437,N_10029,N_10123);
nor U10438 (N_10438,N_10130,N_10062);
or U10439 (N_10439,N_10213,N_10015);
nand U10440 (N_10440,N_10025,N_10195);
or U10441 (N_10441,N_10129,N_10004);
and U10442 (N_10442,N_10183,N_10019);
and U10443 (N_10443,N_10153,N_10088);
xor U10444 (N_10444,N_10058,N_10248);
and U10445 (N_10445,N_10114,N_10088);
or U10446 (N_10446,N_10072,N_10032);
or U10447 (N_10447,N_10022,N_10241);
or U10448 (N_10448,N_10061,N_10189);
xor U10449 (N_10449,N_10184,N_10063);
or U10450 (N_10450,N_10033,N_10046);
nand U10451 (N_10451,N_10231,N_10110);
or U10452 (N_10452,N_10150,N_10171);
nand U10453 (N_10453,N_10197,N_10195);
or U10454 (N_10454,N_10084,N_10158);
or U10455 (N_10455,N_10154,N_10195);
and U10456 (N_10456,N_10031,N_10206);
nand U10457 (N_10457,N_10192,N_10111);
and U10458 (N_10458,N_10081,N_10000);
nand U10459 (N_10459,N_10190,N_10114);
or U10460 (N_10460,N_10004,N_10135);
nand U10461 (N_10461,N_10012,N_10016);
and U10462 (N_10462,N_10026,N_10113);
nand U10463 (N_10463,N_10073,N_10118);
nand U10464 (N_10464,N_10206,N_10231);
xor U10465 (N_10465,N_10192,N_10183);
nor U10466 (N_10466,N_10156,N_10012);
nand U10467 (N_10467,N_10097,N_10109);
nor U10468 (N_10468,N_10083,N_10235);
nand U10469 (N_10469,N_10130,N_10070);
nor U10470 (N_10470,N_10163,N_10203);
and U10471 (N_10471,N_10205,N_10017);
or U10472 (N_10472,N_10178,N_10062);
and U10473 (N_10473,N_10111,N_10094);
or U10474 (N_10474,N_10209,N_10101);
nor U10475 (N_10475,N_10236,N_10043);
nand U10476 (N_10476,N_10068,N_10204);
nand U10477 (N_10477,N_10160,N_10019);
and U10478 (N_10478,N_10158,N_10100);
or U10479 (N_10479,N_10031,N_10109);
and U10480 (N_10480,N_10048,N_10079);
or U10481 (N_10481,N_10169,N_10249);
xor U10482 (N_10482,N_10058,N_10017);
xnor U10483 (N_10483,N_10033,N_10192);
nand U10484 (N_10484,N_10047,N_10199);
nor U10485 (N_10485,N_10095,N_10198);
nand U10486 (N_10486,N_10184,N_10133);
xor U10487 (N_10487,N_10056,N_10146);
nor U10488 (N_10488,N_10000,N_10155);
xnor U10489 (N_10489,N_10038,N_10060);
nor U10490 (N_10490,N_10086,N_10169);
nand U10491 (N_10491,N_10101,N_10240);
nor U10492 (N_10492,N_10092,N_10076);
and U10493 (N_10493,N_10085,N_10240);
or U10494 (N_10494,N_10141,N_10153);
and U10495 (N_10495,N_10101,N_10248);
xor U10496 (N_10496,N_10011,N_10009);
or U10497 (N_10497,N_10011,N_10208);
and U10498 (N_10498,N_10155,N_10103);
and U10499 (N_10499,N_10099,N_10073);
and U10500 (N_10500,N_10274,N_10329);
nand U10501 (N_10501,N_10396,N_10409);
and U10502 (N_10502,N_10452,N_10295);
xor U10503 (N_10503,N_10445,N_10321);
and U10504 (N_10504,N_10455,N_10281);
and U10505 (N_10505,N_10402,N_10314);
nor U10506 (N_10506,N_10359,N_10428);
nor U10507 (N_10507,N_10439,N_10414);
and U10508 (N_10508,N_10421,N_10497);
nand U10509 (N_10509,N_10398,N_10440);
nor U10510 (N_10510,N_10324,N_10433);
or U10511 (N_10511,N_10381,N_10385);
and U10512 (N_10512,N_10446,N_10363);
and U10513 (N_10513,N_10313,N_10411);
or U10514 (N_10514,N_10320,N_10420);
and U10515 (N_10515,N_10304,N_10372);
and U10516 (N_10516,N_10474,N_10494);
and U10517 (N_10517,N_10340,N_10294);
or U10518 (N_10518,N_10480,N_10312);
nand U10519 (N_10519,N_10356,N_10378);
xnor U10520 (N_10520,N_10271,N_10416);
and U10521 (N_10521,N_10283,N_10422);
and U10522 (N_10522,N_10460,N_10308);
xnor U10523 (N_10523,N_10397,N_10386);
xnor U10524 (N_10524,N_10256,N_10262);
xor U10525 (N_10525,N_10395,N_10290);
xnor U10526 (N_10526,N_10392,N_10326);
xnor U10527 (N_10527,N_10318,N_10344);
and U10528 (N_10528,N_10470,N_10465);
nor U10529 (N_10529,N_10337,N_10405);
nor U10530 (N_10530,N_10374,N_10403);
xnor U10531 (N_10531,N_10400,N_10268);
nand U10532 (N_10532,N_10331,N_10347);
nand U10533 (N_10533,N_10469,N_10406);
nor U10534 (N_10534,N_10490,N_10484);
nand U10535 (N_10535,N_10483,N_10430);
nand U10536 (N_10536,N_10479,N_10489);
xor U10537 (N_10537,N_10437,N_10390);
and U10538 (N_10538,N_10250,N_10487);
and U10539 (N_10539,N_10427,N_10473);
or U10540 (N_10540,N_10267,N_10302);
and U10541 (N_10541,N_10301,N_10298);
and U10542 (N_10542,N_10459,N_10441);
xor U10543 (N_10543,N_10463,N_10485);
nor U10544 (N_10544,N_10355,N_10462);
and U10545 (N_10545,N_10266,N_10444);
nand U10546 (N_10546,N_10252,N_10259);
nor U10547 (N_10547,N_10410,N_10388);
nor U10548 (N_10548,N_10453,N_10387);
nor U10549 (N_10549,N_10467,N_10350);
nor U10550 (N_10550,N_10289,N_10415);
and U10551 (N_10551,N_10286,N_10438);
and U10552 (N_10552,N_10419,N_10323);
and U10553 (N_10553,N_10457,N_10491);
xor U10554 (N_10554,N_10309,N_10496);
and U10555 (N_10555,N_10364,N_10270);
nor U10556 (N_10556,N_10448,N_10291);
xor U10557 (N_10557,N_10334,N_10303);
xnor U10558 (N_10558,N_10375,N_10328);
or U10559 (N_10559,N_10341,N_10342);
nand U10560 (N_10560,N_10288,N_10492);
or U10561 (N_10561,N_10273,N_10495);
xor U10562 (N_10562,N_10345,N_10424);
xnor U10563 (N_10563,N_10377,N_10429);
xnor U10564 (N_10564,N_10282,N_10257);
nor U10565 (N_10565,N_10349,N_10316);
nand U10566 (N_10566,N_10351,N_10434);
nand U10567 (N_10567,N_10373,N_10436);
and U10568 (N_10568,N_10454,N_10293);
or U10569 (N_10569,N_10482,N_10315);
or U10570 (N_10570,N_10339,N_10251);
or U10571 (N_10571,N_10263,N_10384);
nand U10572 (N_10572,N_10443,N_10412);
or U10573 (N_10573,N_10407,N_10435);
xnor U10574 (N_10574,N_10404,N_10285);
nand U10575 (N_10575,N_10253,N_10292);
nor U10576 (N_10576,N_10466,N_10338);
and U10577 (N_10577,N_10317,N_10376);
or U10578 (N_10578,N_10343,N_10305);
and U10579 (N_10579,N_10311,N_10335);
nand U10580 (N_10580,N_10475,N_10493);
nor U10581 (N_10581,N_10399,N_10468);
nor U10582 (N_10582,N_10472,N_10394);
and U10583 (N_10583,N_10417,N_10255);
or U10584 (N_10584,N_10279,N_10450);
and U10585 (N_10585,N_10383,N_10449);
or U10586 (N_10586,N_10319,N_10348);
or U10587 (N_10587,N_10481,N_10284);
or U10588 (N_10588,N_10365,N_10477);
and U10589 (N_10589,N_10379,N_10478);
or U10590 (N_10590,N_10307,N_10476);
nand U10591 (N_10591,N_10280,N_10336);
or U10592 (N_10592,N_10451,N_10425);
or U10593 (N_10593,N_10297,N_10471);
or U10594 (N_10594,N_10413,N_10498);
or U10595 (N_10595,N_10393,N_10360);
nand U10596 (N_10596,N_10464,N_10357);
xnor U10597 (N_10597,N_10299,N_10310);
xnor U10598 (N_10598,N_10423,N_10431);
nand U10599 (N_10599,N_10369,N_10277);
nor U10600 (N_10600,N_10380,N_10265);
and U10601 (N_10601,N_10296,N_10426);
nand U10602 (N_10602,N_10272,N_10269);
nor U10603 (N_10603,N_10287,N_10361);
or U10604 (N_10604,N_10300,N_10258);
or U10605 (N_10605,N_10401,N_10260);
xor U10606 (N_10606,N_10264,N_10261);
nor U10607 (N_10607,N_10346,N_10368);
and U10608 (N_10608,N_10382,N_10442);
xnor U10609 (N_10609,N_10254,N_10391);
or U10610 (N_10610,N_10352,N_10327);
xor U10611 (N_10611,N_10371,N_10332);
nand U10612 (N_10612,N_10354,N_10275);
and U10613 (N_10613,N_10408,N_10366);
nand U10614 (N_10614,N_10325,N_10358);
and U10615 (N_10615,N_10456,N_10333);
nor U10616 (N_10616,N_10486,N_10447);
nand U10617 (N_10617,N_10458,N_10488);
and U10618 (N_10618,N_10418,N_10370);
or U10619 (N_10619,N_10389,N_10432);
and U10620 (N_10620,N_10362,N_10306);
nor U10621 (N_10621,N_10276,N_10499);
xor U10622 (N_10622,N_10461,N_10367);
or U10623 (N_10623,N_10322,N_10353);
xnor U10624 (N_10624,N_10278,N_10330);
nand U10625 (N_10625,N_10406,N_10380);
nor U10626 (N_10626,N_10446,N_10260);
or U10627 (N_10627,N_10298,N_10387);
nor U10628 (N_10628,N_10290,N_10325);
xnor U10629 (N_10629,N_10495,N_10436);
nor U10630 (N_10630,N_10490,N_10300);
or U10631 (N_10631,N_10329,N_10285);
nor U10632 (N_10632,N_10387,N_10270);
nand U10633 (N_10633,N_10268,N_10257);
and U10634 (N_10634,N_10299,N_10376);
or U10635 (N_10635,N_10307,N_10467);
nor U10636 (N_10636,N_10371,N_10455);
and U10637 (N_10637,N_10380,N_10351);
nand U10638 (N_10638,N_10310,N_10473);
and U10639 (N_10639,N_10315,N_10405);
and U10640 (N_10640,N_10301,N_10449);
or U10641 (N_10641,N_10398,N_10341);
or U10642 (N_10642,N_10442,N_10415);
nand U10643 (N_10643,N_10445,N_10397);
and U10644 (N_10644,N_10489,N_10306);
or U10645 (N_10645,N_10264,N_10472);
xor U10646 (N_10646,N_10306,N_10285);
xor U10647 (N_10647,N_10358,N_10390);
or U10648 (N_10648,N_10413,N_10383);
or U10649 (N_10649,N_10428,N_10493);
nand U10650 (N_10650,N_10311,N_10481);
xor U10651 (N_10651,N_10462,N_10359);
xor U10652 (N_10652,N_10259,N_10352);
nand U10653 (N_10653,N_10474,N_10303);
or U10654 (N_10654,N_10278,N_10270);
or U10655 (N_10655,N_10279,N_10473);
and U10656 (N_10656,N_10407,N_10481);
and U10657 (N_10657,N_10411,N_10266);
and U10658 (N_10658,N_10306,N_10474);
or U10659 (N_10659,N_10450,N_10475);
xnor U10660 (N_10660,N_10429,N_10369);
xnor U10661 (N_10661,N_10330,N_10493);
nor U10662 (N_10662,N_10335,N_10303);
nand U10663 (N_10663,N_10275,N_10268);
or U10664 (N_10664,N_10469,N_10413);
nor U10665 (N_10665,N_10353,N_10399);
xor U10666 (N_10666,N_10462,N_10309);
nand U10667 (N_10667,N_10311,N_10280);
xnor U10668 (N_10668,N_10347,N_10289);
and U10669 (N_10669,N_10308,N_10436);
nor U10670 (N_10670,N_10298,N_10340);
nand U10671 (N_10671,N_10262,N_10321);
and U10672 (N_10672,N_10290,N_10438);
or U10673 (N_10673,N_10438,N_10302);
or U10674 (N_10674,N_10438,N_10306);
or U10675 (N_10675,N_10273,N_10441);
nand U10676 (N_10676,N_10450,N_10491);
and U10677 (N_10677,N_10467,N_10357);
and U10678 (N_10678,N_10281,N_10479);
xnor U10679 (N_10679,N_10413,N_10484);
nand U10680 (N_10680,N_10392,N_10255);
nand U10681 (N_10681,N_10260,N_10319);
and U10682 (N_10682,N_10271,N_10287);
and U10683 (N_10683,N_10438,N_10254);
and U10684 (N_10684,N_10448,N_10397);
or U10685 (N_10685,N_10434,N_10477);
or U10686 (N_10686,N_10330,N_10356);
xnor U10687 (N_10687,N_10435,N_10393);
or U10688 (N_10688,N_10325,N_10298);
nor U10689 (N_10689,N_10372,N_10335);
or U10690 (N_10690,N_10473,N_10482);
and U10691 (N_10691,N_10398,N_10355);
nor U10692 (N_10692,N_10386,N_10300);
or U10693 (N_10693,N_10435,N_10427);
or U10694 (N_10694,N_10260,N_10352);
xnor U10695 (N_10695,N_10432,N_10418);
and U10696 (N_10696,N_10356,N_10488);
and U10697 (N_10697,N_10467,N_10314);
nand U10698 (N_10698,N_10448,N_10431);
nor U10699 (N_10699,N_10329,N_10341);
and U10700 (N_10700,N_10453,N_10463);
xnor U10701 (N_10701,N_10425,N_10307);
nand U10702 (N_10702,N_10289,N_10250);
nand U10703 (N_10703,N_10362,N_10482);
nor U10704 (N_10704,N_10460,N_10355);
nand U10705 (N_10705,N_10447,N_10351);
or U10706 (N_10706,N_10268,N_10303);
nor U10707 (N_10707,N_10255,N_10289);
and U10708 (N_10708,N_10367,N_10327);
and U10709 (N_10709,N_10492,N_10444);
and U10710 (N_10710,N_10389,N_10360);
or U10711 (N_10711,N_10491,N_10305);
or U10712 (N_10712,N_10497,N_10304);
nor U10713 (N_10713,N_10388,N_10454);
nor U10714 (N_10714,N_10454,N_10335);
xor U10715 (N_10715,N_10409,N_10270);
or U10716 (N_10716,N_10464,N_10418);
nor U10717 (N_10717,N_10486,N_10326);
xnor U10718 (N_10718,N_10382,N_10319);
nand U10719 (N_10719,N_10318,N_10454);
or U10720 (N_10720,N_10445,N_10271);
xnor U10721 (N_10721,N_10294,N_10267);
xor U10722 (N_10722,N_10435,N_10420);
and U10723 (N_10723,N_10368,N_10344);
nand U10724 (N_10724,N_10400,N_10325);
or U10725 (N_10725,N_10310,N_10346);
nor U10726 (N_10726,N_10434,N_10337);
xnor U10727 (N_10727,N_10496,N_10406);
or U10728 (N_10728,N_10260,N_10268);
nor U10729 (N_10729,N_10395,N_10291);
nand U10730 (N_10730,N_10327,N_10329);
xnor U10731 (N_10731,N_10262,N_10399);
and U10732 (N_10732,N_10364,N_10386);
nand U10733 (N_10733,N_10330,N_10309);
or U10734 (N_10734,N_10288,N_10438);
or U10735 (N_10735,N_10275,N_10489);
nand U10736 (N_10736,N_10394,N_10366);
xor U10737 (N_10737,N_10372,N_10418);
nand U10738 (N_10738,N_10362,N_10376);
or U10739 (N_10739,N_10279,N_10493);
and U10740 (N_10740,N_10255,N_10290);
or U10741 (N_10741,N_10258,N_10330);
nand U10742 (N_10742,N_10310,N_10301);
nand U10743 (N_10743,N_10415,N_10471);
or U10744 (N_10744,N_10389,N_10427);
nand U10745 (N_10745,N_10470,N_10350);
nor U10746 (N_10746,N_10339,N_10375);
nand U10747 (N_10747,N_10320,N_10274);
nand U10748 (N_10748,N_10285,N_10326);
xor U10749 (N_10749,N_10492,N_10392);
and U10750 (N_10750,N_10657,N_10622);
or U10751 (N_10751,N_10713,N_10565);
xor U10752 (N_10752,N_10562,N_10735);
or U10753 (N_10753,N_10558,N_10568);
and U10754 (N_10754,N_10700,N_10736);
or U10755 (N_10755,N_10682,N_10672);
and U10756 (N_10756,N_10689,N_10704);
xnor U10757 (N_10757,N_10506,N_10570);
xor U10758 (N_10758,N_10712,N_10597);
nand U10759 (N_10759,N_10602,N_10635);
xnor U10760 (N_10760,N_10746,N_10652);
and U10761 (N_10761,N_10545,N_10518);
nand U10762 (N_10762,N_10728,N_10690);
xor U10763 (N_10763,N_10738,N_10503);
nor U10764 (N_10764,N_10705,N_10547);
or U10765 (N_10765,N_10594,N_10541);
nor U10766 (N_10766,N_10725,N_10701);
xor U10767 (N_10767,N_10715,N_10677);
and U10768 (N_10768,N_10663,N_10519);
xnor U10769 (N_10769,N_10645,N_10505);
or U10770 (N_10770,N_10706,N_10520);
or U10771 (N_10771,N_10563,N_10685);
nand U10772 (N_10772,N_10630,N_10721);
and U10773 (N_10773,N_10666,N_10532);
nor U10774 (N_10774,N_10687,N_10676);
nor U10775 (N_10775,N_10683,N_10620);
xnor U10776 (N_10776,N_10569,N_10743);
xor U10777 (N_10777,N_10637,N_10732);
or U10778 (N_10778,N_10688,N_10609);
and U10779 (N_10779,N_10729,N_10640);
xnor U10780 (N_10780,N_10703,N_10686);
nand U10781 (N_10781,N_10698,N_10525);
nor U10782 (N_10782,N_10572,N_10575);
or U10783 (N_10783,N_10508,N_10718);
or U10784 (N_10784,N_10650,N_10542);
and U10785 (N_10785,N_10539,N_10606);
nor U10786 (N_10786,N_10538,N_10692);
nand U10787 (N_10787,N_10591,N_10707);
nand U10788 (N_10788,N_10583,N_10509);
or U10789 (N_10789,N_10550,N_10739);
or U10790 (N_10790,N_10699,N_10643);
nand U10791 (N_10791,N_10719,N_10574);
nand U10792 (N_10792,N_10559,N_10566);
nor U10793 (N_10793,N_10593,N_10576);
nand U10794 (N_10794,N_10561,N_10530);
or U10795 (N_10795,N_10618,N_10596);
nor U10796 (N_10796,N_10610,N_10616);
and U10797 (N_10797,N_10534,N_10653);
and U10798 (N_10798,N_10533,N_10727);
nand U10799 (N_10799,N_10536,N_10709);
or U10800 (N_10800,N_10669,N_10678);
nand U10801 (N_10801,N_10749,N_10560);
xor U10802 (N_10802,N_10580,N_10555);
xor U10803 (N_10803,N_10543,N_10614);
xnor U10804 (N_10804,N_10649,N_10624);
or U10805 (N_10805,N_10540,N_10680);
nor U10806 (N_10806,N_10553,N_10512);
and U10807 (N_10807,N_10599,N_10537);
or U10808 (N_10808,N_10696,N_10517);
nand U10809 (N_10809,N_10548,N_10639);
nand U10810 (N_10810,N_10664,N_10582);
nor U10811 (N_10811,N_10651,N_10590);
and U10812 (N_10812,N_10507,N_10720);
or U10813 (N_10813,N_10510,N_10668);
and U10814 (N_10814,N_10638,N_10697);
xnor U10815 (N_10815,N_10629,N_10611);
or U10816 (N_10816,N_10551,N_10586);
nor U10817 (N_10817,N_10607,N_10601);
or U10818 (N_10818,N_10625,N_10722);
and U10819 (N_10819,N_10714,N_10675);
nand U10820 (N_10820,N_10628,N_10627);
and U10821 (N_10821,N_10577,N_10617);
nor U10822 (N_10822,N_10605,N_10587);
or U10823 (N_10823,N_10619,N_10531);
nor U10824 (N_10824,N_10702,N_10581);
xnor U10825 (N_10825,N_10571,N_10573);
and U10826 (N_10826,N_10513,N_10521);
nand U10827 (N_10827,N_10679,N_10578);
and U10828 (N_10828,N_10710,N_10684);
nand U10829 (N_10829,N_10589,N_10623);
and U10830 (N_10830,N_10667,N_10644);
or U10831 (N_10831,N_10671,N_10633);
xor U10832 (N_10832,N_10726,N_10552);
nor U10833 (N_10833,N_10724,N_10527);
and U10834 (N_10834,N_10656,N_10529);
nand U10835 (N_10835,N_10579,N_10544);
nand U10836 (N_10836,N_10654,N_10546);
nand U10837 (N_10837,N_10691,N_10695);
xnor U10838 (N_10838,N_10584,N_10501);
nor U10839 (N_10839,N_10693,N_10516);
xor U10840 (N_10840,N_10708,N_10740);
or U10841 (N_10841,N_10681,N_10603);
and U10842 (N_10842,N_10608,N_10535);
or U10843 (N_10843,N_10741,N_10665);
or U10844 (N_10844,N_10648,N_10647);
xor U10845 (N_10845,N_10658,N_10604);
nand U10846 (N_10846,N_10564,N_10747);
xor U10847 (N_10847,N_10661,N_10549);
or U10848 (N_10848,N_10673,N_10612);
nor U10849 (N_10849,N_10744,N_10557);
nand U10850 (N_10850,N_10659,N_10515);
or U10851 (N_10851,N_10621,N_10522);
xnor U10852 (N_10852,N_10567,N_10500);
xor U10853 (N_10853,N_10730,N_10626);
xor U10854 (N_10854,N_10655,N_10748);
nor U10855 (N_10855,N_10556,N_10528);
nand U10856 (N_10856,N_10731,N_10631);
or U10857 (N_10857,N_10588,N_10511);
nor U10858 (N_10858,N_10733,N_10592);
nor U10859 (N_10859,N_10634,N_10742);
nand U10860 (N_10860,N_10524,N_10504);
and U10861 (N_10861,N_10642,N_10615);
xor U10862 (N_10862,N_10660,N_10502);
nand U10863 (N_10863,N_10737,N_10600);
and U10864 (N_10864,N_10711,N_10723);
nor U10865 (N_10865,N_10716,N_10526);
or U10866 (N_10866,N_10717,N_10745);
xnor U10867 (N_10867,N_10523,N_10662);
nor U10868 (N_10868,N_10694,N_10595);
and U10869 (N_10869,N_10641,N_10554);
xnor U10870 (N_10870,N_10734,N_10674);
nor U10871 (N_10871,N_10646,N_10613);
or U10872 (N_10872,N_10632,N_10670);
or U10873 (N_10873,N_10598,N_10585);
and U10874 (N_10874,N_10636,N_10514);
nand U10875 (N_10875,N_10636,N_10533);
nand U10876 (N_10876,N_10700,N_10615);
xor U10877 (N_10877,N_10546,N_10624);
xnor U10878 (N_10878,N_10626,N_10537);
nor U10879 (N_10879,N_10713,N_10574);
or U10880 (N_10880,N_10715,N_10642);
or U10881 (N_10881,N_10511,N_10646);
and U10882 (N_10882,N_10539,N_10537);
nand U10883 (N_10883,N_10549,N_10504);
nor U10884 (N_10884,N_10547,N_10745);
nor U10885 (N_10885,N_10747,N_10502);
or U10886 (N_10886,N_10549,N_10555);
nand U10887 (N_10887,N_10735,N_10572);
xnor U10888 (N_10888,N_10658,N_10710);
nand U10889 (N_10889,N_10533,N_10696);
and U10890 (N_10890,N_10690,N_10656);
xor U10891 (N_10891,N_10511,N_10603);
and U10892 (N_10892,N_10565,N_10689);
and U10893 (N_10893,N_10652,N_10727);
nor U10894 (N_10894,N_10702,N_10739);
xor U10895 (N_10895,N_10621,N_10678);
and U10896 (N_10896,N_10714,N_10564);
nand U10897 (N_10897,N_10643,N_10648);
nand U10898 (N_10898,N_10550,N_10678);
xor U10899 (N_10899,N_10516,N_10691);
and U10900 (N_10900,N_10592,N_10562);
or U10901 (N_10901,N_10700,N_10606);
or U10902 (N_10902,N_10681,N_10561);
nand U10903 (N_10903,N_10645,N_10693);
and U10904 (N_10904,N_10710,N_10644);
nand U10905 (N_10905,N_10555,N_10572);
nor U10906 (N_10906,N_10747,N_10624);
nor U10907 (N_10907,N_10616,N_10743);
and U10908 (N_10908,N_10595,N_10679);
or U10909 (N_10909,N_10564,N_10638);
and U10910 (N_10910,N_10673,N_10526);
or U10911 (N_10911,N_10605,N_10596);
xnor U10912 (N_10912,N_10723,N_10513);
nor U10913 (N_10913,N_10553,N_10674);
nand U10914 (N_10914,N_10606,N_10720);
nand U10915 (N_10915,N_10671,N_10717);
nand U10916 (N_10916,N_10589,N_10666);
nor U10917 (N_10917,N_10742,N_10598);
and U10918 (N_10918,N_10575,N_10574);
xnor U10919 (N_10919,N_10537,N_10592);
and U10920 (N_10920,N_10522,N_10629);
xor U10921 (N_10921,N_10602,N_10571);
nand U10922 (N_10922,N_10593,N_10546);
and U10923 (N_10923,N_10663,N_10602);
and U10924 (N_10924,N_10621,N_10611);
nor U10925 (N_10925,N_10557,N_10620);
xnor U10926 (N_10926,N_10656,N_10749);
nor U10927 (N_10927,N_10646,N_10712);
nor U10928 (N_10928,N_10518,N_10636);
and U10929 (N_10929,N_10652,N_10736);
and U10930 (N_10930,N_10518,N_10649);
nor U10931 (N_10931,N_10711,N_10661);
nand U10932 (N_10932,N_10583,N_10515);
or U10933 (N_10933,N_10678,N_10717);
nor U10934 (N_10934,N_10615,N_10562);
nand U10935 (N_10935,N_10683,N_10629);
or U10936 (N_10936,N_10511,N_10614);
and U10937 (N_10937,N_10601,N_10651);
nand U10938 (N_10938,N_10633,N_10600);
or U10939 (N_10939,N_10595,N_10531);
nor U10940 (N_10940,N_10701,N_10573);
nand U10941 (N_10941,N_10551,N_10572);
or U10942 (N_10942,N_10603,N_10585);
xor U10943 (N_10943,N_10581,N_10688);
and U10944 (N_10944,N_10505,N_10641);
or U10945 (N_10945,N_10612,N_10572);
or U10946 (N_10946,N_10581,N_10655);
and U10947 (N_10947,N_10512,N_10545);
nor U10948 (N_10948,N_10721,N_10687);
nor U10949 (N_10949,N_10692,N_10547);
and U10950 (N_10950,N_10660,N_10534);
or U10951 (N_10951,N_10680,N_10740);
and U10952 (N_10952,N_10587,N_10685);
xor U10953 (N_10953,N_10556,N_10634);
nand U10954 (N_10954,N_10666,N_10682);
and U10955 (N_10955,N_10606,N_10638);
xnor U10956 (N_10956,N_10617,N_10687);
or U10957 (N_10957,N_10698,N_10711);
or U10958 (N_10958,N_10574,N_10727);
nand U10959 (N_10959,N_10742,N_10693);
nand U10960 (N_10960,N_10686,N_10521);
nand U10961 (N_10961,N_10702,N_10728);
nor U10962 (N_10962,N_10533,N_10500);
and U10963 (N_10963,N_10568,N_10677);
or U10964 (N_10964,N_10536,N_10531);
or U10965 (N_10965,N_10688,N_10676);
nor U10966 (N_10966,N_10569,N_10525);
or U10967 (N_10967,N_10703,N_10658);
xnor U10968 (N_10968,N_10724,N_10631);
xor U10969 (N_10969,N_10613,N_10578);
nand U10970 (N_10970,N_10561,N_10737);
nor U10971 (N_10971,N_10548,N_10743);
and U10972 (N_10972,N_10598,N_10650);
xnor U10973 (N_10973,N_10728,N_10709);
or U10974 (N_10974,N_10530,N_10577);
xor U10975 (N_10975,N_10715,N_10621);
nor U10976 (N_10976,N_10627,N_10655);
or U10977 (N_10977,N_10643,N_10607);
nor U10978 (N_10978,N_10730,N_10684);
xnor U10979 (N_10979,N_10719,N_10505);
xnor U10980 (N_10980,N_10624,N_10545);
nand U10981 (N_10981,N_10732,N_10720);
nand U10982 (N_10982,N_10588,N_10603);
xor U10983 (N_10983,N_10729,N_10676);
xnor U10984 (N_10984,N_10503,N_10678);
or U10985 (N_10985,N_10748,N_10725);
nand U10986 (N_10986,N_10649,N_10601);
nand U10987 (N_10987,N_10709,N_10652);
xnor U10988 (N_10988,N_10711,N_10674);
nor U10989 (N_10989,N_10714,N_10526);
xnor U10990 (N_10990,N_10717,N_10733);
and U10991 (N_10991,N_10637,N_10502);
and U10992 (N_10992,N_10511,N_10642);
xnor U10993 (N_10993,N_10748,N_10588);
xor U10994 (N_10994,N_10660,N_10526);
and U10995 (N_10995,N_10718,N_10621);
nor U10996 (N_10996,N_10562,N_10525);
or U10997 (N_10997,N_10684,N_10716);
xnor U10998 (N_10998,N_10553,N_10730);
nor U10999 (N_10999,N_10614,N_10656);
and U11000 (N_11000,N_10781,N_10904);
or U11001 (N_11001,N_10896,N_10816);
or U11002 (N_11002,N_10988,N_10960);
xor U11003 (N_11003,N_10795,N_10940);
or U11004 (N_11004,N_10894,N_10970);
nor U11005 (N_11005,N_10887,N_10989);
nand U11006 (N_11006,N_10953,N_10804);
and U11007 (N_11007,N_10885,N_10939);
and U11008 (N_11008,N_10875,N_10874);
nor U11009 (N_11009,N_10857,N_10907);
nor U11010 (N_11010,N_10780,N_10889);
nor U11011 (N_11011,N_10976,N_10846);
and U11012 (N_11012,N_10901,N_10829);
and U11013 (N_11013,N_10883,N_10784);
nor U11014 (N_11014,N_10937,N_10991);
nand U11015 (N_11015,N_10802,N_10975);
nor U11016 (N_11016,N_10929,N_10872);
and U11017 (N_11017,N_10933,N_10965);
xnor U11018 (N_11018,N_10941,N_10915);
and U11019 (N_11019,N_10899,N_10811);
xnor U11020 (N_11020,N_10777,N_10759);
and U11021 (N_11021,N_10834,N_10840);
and U11022 (N_11022,N_10832,N_10876);
nor U11023 (N_11023,N_10974,N_10779);
nand U11024 (N_11024,N_10958,N_10823);
or U11025 (N_11025,N_10870,N_10842);
xor U11026 (N_11026,N_10961,N_10789);
nand U11027 (N_11027,N_10805,N_10987);
xnor U11028 (N_11028,N_10930,N_10913);
xor U11029 (N_11029,N_10962,N_10757);
or U11030 (N_11030,N_10798,N_10931);
xor U11031 (N_11031,N_10888,N_10927);
nor U11032 (N_11032,N_10910,N_10853);
nor U11033 (N_11033,N_10905,N_10922);
nand U11034 (N_11034,N_10774,N_10864);
and U11035 (N_11035,N_10914,N_10812);
nand U11036 (N_11036,N_10978,N_10850);
xnor U11037 (N_11037,N_10835,N_10790);
nand U11038 (N_11038,N_10918,N_10977);
or U11039 (N_11039,N_10868,N_10766);
nor U11040 (N_11040,N_10856,N_10809);
nand U11041 (N_11041,N_10878,N_10803);
or U11042 (N_11042,N_10908,N_10843);
nor U11043 (N_11043,N_10955,N_10919);
nor U11044 (N_11044,N_10821,N_10928);
xnor U11045 (N_11045,N_10946,N_10860);
xor U11046 (N_11046,N_10817,N_10971);
and U11047 (N_11047,N_10851,N_10818);
nor U11048 (N_11048,N_10898,N_10964);
nand U11049 (N_11049,N_10943,N_10893);
and U11050 (N_11050,N_10813,N_10948);
xor U11051 (N_11051,N_10873,N_10782);
xnor U11052 (N_11052,N_10882,N_10830);
or U11053 (N_11053,N_10980,N_10932);
nand U11054 (N_11054,N_10753,N_10909);
xor U11055 (N_11055,N_10773,N_10886);
xor U11056 (N_11056,N_10819,N_10900);
nor U11057 (N_11057,N_10848,N_10847);
and U11058 (N_11058,N_10767,N_10996);
xnor U11059 (N_11059,N_10994,N_10778);
nor U11060 (N_11060,N_10892,N_10810);
xor U11061 (N_11061,N_10799,N_10825);
nand U11062 (N_11062,N_10783,N_10897);
or U11063 (N_11063,N_10787,N_10984);
nor U11064 (N_11064,N_10770,N_10979);
or U11065 (N_11065,N_10895,N_10827);
nor U11066 (N_11066,N_10833,N_10866);
nor U11067 (N_11067,N_10902,N_10890);
xnor U11068 (N_11068,N_10951,N_10761);
nor U11069 (N_11069,N_10754,N_10785);
nand U11070 (N_11070,N_10775,N_10763);
xnor U11071 (N_11071,N_10750,N_10966);
nand U11072 (N_11072,N_10983,N_10801);
xnor U11073 (N_11073,N_10815,N_10935);
and U11074 (N_11074,N_10982,N_10942);
nor U11075 (N_11075,N_10924,N_10891);
nor U11076 (N_11076,N_10758,N_10755);
and U11077 (N_11077,N_10800,N_10752);
nand U11078 (N_11078,N_10877,N_10852);
nor U11079 (N_11079,N_10995,N_10926);
xor U11080 (N_11080,N_10884,N_10865);
nand U11081 (N_11081,N_10957,N_10950);
nand U11082 (N_11082,N_10796,N_10776);
nand U11083 (N_11083,N_10792,N_10985);
nand U11084 (N_11084,N_10954,N_10938);
nor U11085 (N_11085,N_10997,N_10765);
and U11086 (N_11086,N_10786,N_10969);
nor U11087 (N_11087,N_10838,N_10855);
or U11088 (N_11088,N_10934,N_10925);
nor U11089 (N_11089,N_10764,N_10820);
nor U11090 (N_11090,N_10854,N_10945);
nand U11091 (N_11091,N_10963,N_10772);
and U11092 (N_11092,N_10871,N_10920);
nor U11093 (N_11093,N_10992,N_10822);
nand U11094 (N_11094,N_10956,N_10849);
and U11095 (N_11095,N_10807,N_10771);
nor U11096 (N_11096,N_10862,N_10993);
xnor U11097 (N_11097,N_10769,N_10867);
nand U11098 (N_11098,N_10916,N_10831);
nor U11099 (N_11099,N_10828,N_10797);
xor U11100 (N_11100,N_10949,N_10826);
nor U11101 (N_11101,N_10990,N_10912);
xor U11102 (N_11102,N_10788,N_10986);
or U11103 (N_11103,N_10808,N_10768);
xnor U11104 (N_11104,N_10858,N_10972);
and U11105 (N_11105,N_10814,N_10760);
and U11106 (N_11106,N_10998,N_10999);
nor U11107 (N_11107,N_10824,N_10844);
nand U11108 (N_11108,N_10880,N_10917);
or U11109 (N_11109,N_10881,N_10947);
xor U11110 (N_11110,N_10837,N_10903);
nand U11111 (N_11111,N_10762,N_10952);
or U11112 (N_11112,N_10859,N_10879);
xnor U11113 (N_11113,N_10973,N_10959);
or U11114 (N_11114,N_10968,N_10861);
and U11115 (N_11115,N_10836,N_10923);
xnor U11116 (N_11116,N_10793,N_10936);
xnor U11117 (N_11117,N_10863,N_10756);
or U11118 (N_11118,N_10906,N_10911);
or U11119 (N_11119,N_10967,N_10806);
xnor U11120 (N_11120,N_10921,N_10751);
xor U11121 (N_11121,N_10791,N_10845);
xnor U11122 (N_11122,N_10944,N_10839);
xnor U11123 (N_11123,N_10794,N_10841);
nor U11124 (N_11124,N_10981,N_10869);
nand U11125 (N_11125,N_10757,N_10873);
xor U11126 (N_11126,N_10772,N_10974);
and U11127 (N_11127,N_10815,N_10905);
or U11128 (N_11128,N_10779,N_10821);
nor U11129 (N_11129,N_10919,N_10808);
and U11130 (N_11130,N_10860,N_10957);
or U11131 (N_11131,N_10833,N_10993);
xor U11132 (N_11132,N_10758,N_10995);
nand U11133 (N_11133,N_10926,N_10966);
nor U11134 (N_11134,N_10778,N_10877);
or U11135 (N_11135,N_10850,N_10997);
or U11136 (N_11136,N_10927,N_10893);
or U11137 (N_11137,N_10862,N_10902);
and U11138 (N_11138,N_10824,N_10799);
or U11139 (N_11139,N_10907,N_10999);
and U11140 (N_11140,N_10975,N_10978);
or U11141 (N_11141,N_10877,N_10832);
and U11142 (N_11142,N_10814,N_10976);
nand U11143 (N_11143,N_10869,N_10983);
and U11144 (N_11144,N_10755,N_10813);
and U11145 (N_11145,N_10828,N_10896);
or U11146 (N_11146,N_10826,N_10757);
and U11147 (N_11147,N_10849,N_10893);
nand U11148 (N_11148,N_10849,N_10966);
or U11149 (N_11149,N_10931,N_10840);
nor U11150 (N_11150,N_10807,N_10981);
xnor U11151 (N_11151,N_10809,N_10866);
nand U11152 (N_11152,N_10909,N_10944);
and U11153 (N_11153,N_10878,N_10835);
nand U11154 (N_11154,N_10865,N_10763);
nand U11155 (N_11155,N_10916,N_10790);
nand U11156 (N_11156,N_10809,N_10767);
nand U11157 (N_11157,N_10921,N_10879);
nor U11158 (N_11158,N_10923,N_10986);
nor U11159 (N_11159,N_10976,N_10847);
xnor U11160 (N_11160,N_10940,N_10978);
nand U11161 (N_11161,N_10871,N_10970);
xor U11162 (N_11162,N_10919,N_10988);
nand U11163 (N_11163,N_10897,N_10908);
xnor U11164 (N_11164,N_10890,N_10868);
xor U11165 (N_11165,N_10946,N_10828);
nor U11166 (N_11166,N_10880,N_10954);
nor U11167 (N_11167,N_10912,N_10916);
nor U11168 (N_11168,N_10820,N_10894);
nand U11169 (N_11169,N_10884,N_10832);
or U11170 (N_11170,N_10895,N_10995);
or U11171 (N_11171,N_10771,N_10960);
xor U11172 (N_11172,N_10759,N_10853);
nor U11173 (N_11173,N_10927,N_10946);
nor U11174 (N_11174,N_10922,N_10787);
nor U11175 (N_11175,N_10851,N_10919);
or U11176 (N_11176,N_10830,N_10829);
or U11177 (N_11177,N_10950,N_10835);
xnor U11178 (N_11178,N_10753,N_10843);
or U11179 (N_11179,N_10811,N_10885);
and U11180 (N_11180,N_10856,N_10919);
or U11181 (N_11181,N_10816,N_10866);
nor U11182 (N_11182,N_10821,N_10932);
nand U11183 (N_11183,N_10931,N_10996);
or U11184 (N_11184,N_10980,N_10803);
and U11185 (N_11185,N_10869,N_10790);
nand U11186 (N_11186,N_10909,N_10844);
nand U11187 (N_11187,N_10797,N_10940);
and U11188 (N_11188,N_10888,N_10875);
and U11189 (N_11189,N_10906,N_10803);
and U11190 (N_11190,N_10959,N_10822);
and U11191 (N_11191,N_10755,N_10790);
or U11192 (N_11192,N_10803,N_10989);
nor U11193 (N_11193,N_10764,N_10752);
nor U11194 (N_11194,N_10980,N_10754);
nand U11195 (N_11195,N_10965,N_10951);
nand U11196 (N_11196,N_10804,N_10990);
nand U11197 (N_11197,N_10933,N_10890);
nand U11198 (N_11198,N_10826,N_10909);
or U11199 (N_11199,N_10827,N_10991);
xor U11200 (N_11200,N_10824,N_10873);
xor U11201 (N_11201,N_10929,N_10818);
or U11202 (N_11202,N_10759,N_10829);
xor U11203 (N_11203,N_10875,N_10821);
nor U11204 (N_11204,N_10852,N_10956);
and U11205 (N_11205,N_10883,N_10908);
nand U11206 (N_11206,N_10819,N_10889);
nor U11207 (N_11207,N_10979,N_10988);
nor U11208 (N_11208,N_10871,N_10849);
nor U11209 (N_11209,N_10965,N_10816);
nor U11210 (N_11210,N_10811,N_10775);
xor U11211 (N_11211,N_10939,N_10861);
nor U11212 (N_11212,N_10986,N_10965);
nand U11213 (N_11213,N_10853,N_10857);
nor U11214 (N_11214,N_10766,N_10769);
nor U11215 (N_11215,N_10917,N_10807);
xor U11216 (N_11216,N_10768,N_10782);
and U11217 (N_11217,N_10943,N_10927);
and U11218 (N_11218,N_10767,N_10942);
nor U11219 (N_11219,N_10850,N_10945);
nand U11220 (N_11220,N_10944,N_10780);
and U11221 (N_11221,N_10809,N_10950);
xnor U11222 (N_11222,N_10827,N_10924);
nor U11223 (N_11223,N_10928,N_10931);
or U11224 (N_11224,N_10959,N_10931);
xor U11225 (N_11225,N_10876,N_10752);
or U11226 (N_11226,N_10978,N_10864);
nor U11227 (N_11227,N_10861,N_10776);
nor U11228 (N_11228,N_10905,N_10777);
xor U11229 (N_11229,N_10958,N_10811);
xnor U11230 (N_11230,N_10990,N_10872);
and U11231 (N_11231,N_10924,N_10990);
xnor U11232 (N_11232,N_10794,N_10785);
nor U11233 (N_11233,N_10977,N_10996);
xnor U11234 (N_11234,N_10965,N_10802);
or U11235 (N_11235,N_10785,N_10915);
nand U11236 (N_11236,N_10765,N_10859);
nor U11237 (N_11237,N_10812,N_10891);
xor U11238 (N_11238,N_10784,N_10866);
nor U11239 (N_11239,N_10950,N_10754);
or U11240 (N_11240,N_10798,N_10911);
nand U11241 (N_11241,N_10967,N_10893);
nand U11242 (N_11242,N_10948,N_10925);
nor U11243 (N_11243,N_10801,N_10814);
nand U11244 (N_11244,N_10857,N_10768);
nor U11245 (N_11245,N_10901,N_10904);
xnor U11246 (N_11246,N_10950,N_10965);
nor U11247 (N_11247,N_10930,N_10946);
nor U11248 (N_11248,N_10920,N_10820);
nand U11249 (N_11249,N_10901,N_10827);
nand U11250 (N_11250,N_11148,N_11220);
xor U11251 (N_11251,N_11201,N_11244);
nor U11252 (N_11252,N_11014,N_11233);
and U11253 (N_11253,N_11139,N_11223);
nand U11254 (N_11254,N_11144,N_11023);
nand U11255 (N_11255,N_11130,N_11133);
or U11256 (N_11256,N_11041,N_11132);
nand U11257 (N_11257,N_11001,N_11020);
nor U11258 (N_11258,N_11157,N_11056);
xnor U11259 (N_11259,N_11111,N_11225);
nand U11260 (N_11260,N_11228,N_11007);
and U11261 (N_11261,N_11052,N_11069);
xnor U11262 (N_11262,N_11150,N_11018);
or U11263 (N_11263,N_11151,N_11175);
xor U11264 (N_11264,N_11013,N_11221);
or U11265 (N_11265,N_11190,N_11029);
nand U11266 (N_11266,N_11181,N_11247);
or U11267 (N_11267,N_11083,N_11009);
and U11268 (N_11268,N_11230,N_11167);
xor U11269 (N_11269,N_11224,N_11030);
nor U11270 (N_11270,N_11153,N_11174);
nand U11271 (N_11271,N_11027,N_11168);
and U11272 (N_11272,N_11155,N_11022);
or U11273 (N_11273,N_11047,N_11234);
xor U11274 (N_11274,N_11037,N_11015);
and U11275 (N_11275,N_11112,N_11060);
nor U11276 (N_11276,N_11193,N_11004);
and U11277 (N_11277,N_11248,N_11238);
or U11278 (N_11278,N_11140,N_11191);
nand U11279 (N_11279,N_11057,N_11072);
xnor U11280 (N_11280,N_11040,N_11078);
nor U11281 (N_11281,N_11184,N_11171);
xnor U11282 (N_11282,N_11128,N_11046);
xnor U11283 (N_11283,N_11203,N_11218);
nor U11284 (N_11284,N_11079,N_11158);
and U11285 (N_11285,N_11156,N_11085);
or U11286 (N_11286,N_11162,N_11241);
or U11287 (N_11287,N_11061,N_11011);
or U11288 (N_11288,N_11043,N_11063);
nand U11289 (N_11289,N_11169,N_11135);
or U11290 (N_11290,N_11208,N_11067);
xor U11291 (N_11291,N_11245,N_11141);
and U11292 (N_11292,N_11229,N_11149);
or U11293 (N_11293,N_11104,N_11075);
nand U11294 (N_11294,N_11076,N_11180);
xor U11295 (N_11295,N_11217,N_11045);
and U11296 (N_11296,N_11071,N_11161);
and U11297 (N_11297,N_11219,N_11206);
nand U11298 (N_11298,N_11235,N_11202);
xnor U11299 (N_11299,N_11215,N_11145);
nor U11300 (N_11300,N_11098,N_11124);
nor U11301 (N_11301,N_11138,N_11086);
or U11302 (N_11302,N_11088,N_11142);
xnor U11303 (N_11303,N_11147,N_11212);
or U11304 (N_11304,N_11077,N_11107);
nor U11305 (N_11305,N_11110,N_11105);
or U11306 (N_11306,N_11050,N_11249);
nand U11307 (N_11307,N_11242,N_11092);
and U11308 (N_11308,N_11048,N_11231);
or U11309 (N_11309,N_11134,N_11003);
nor U11310 (N_11310,N_11146,N_11097);
nor U11311 (N_11311,N_11000,N_11035);
nor U11312 (N_11312,N_11197,N_11089);
or U11313 (N_11313,N_11164,N_11044);
nor U11314 (N_11314,N_11154,N_11006);
nor U11315 (N_11315,N_11049,N_11096);
xnor U11316 (N_11316,N_11173,N_11166);
nand U11317 (N_11317,N_11002,N_11059);
xor U11318 (N_11318,N_11116,N_11207);
xnor U11319 (N_11319,N_11125,N_11042);
nor U11320 (N_11320,N_11131,N_11159);
nor U11321 (N_11321,N_11216,N_11120);
xnor U11322 (N_11322,N_11054,N_11080);
or U11323 (N_11323,N_11036,N_11198);
and U11324 (N_11324,N_11113,N_11055);
nand U11325 (N_11325,N_11199,N_11033);
and U11326 (N_11326,N_11081,N_11152);
or U11327 (N_11327,N_11091,N_11196);
or U11328 (N_11328,N_11211,N_11185);
xnor U11329 (N_11329,N_11090,N_11100);
or U11330 (N_11330,N_11237,N_11165);
nand U11331 (N_11331,N_11010,N_11160);
xnor U11332 (N_11332,N_11119,N_11017);
or U11333 (N_11333,N_11213,N_11176);
or U11334 (N_11334,N_11031,N_11205);
nand U11335 (N_11335,N_11227,N_11024);
and U11336 (N_11336,N_11222,N_11170);
nor U11337 (N_11337,N_11058,N_11129);
and U11338 (N_11338,N_11062,N_11019);
and U11339 (N_11339,N_11204,N_11115);
nand U11340 (N_11340,N_11200,N_11183);
and U11341 (N_11341,N_11095,N_11194);
or U11342 (N_11342,N_11070,N_11051);
xnor U11343 (N_11343,N_11122,N_11103);
nand U11344 (N_11344,N_11239,N_11082);
and U11345 (N_11345,N_11137,N_11240);
and U11346 (N_11346,N_11178,N_11232);
xor U11347 (N_11347,N_11118,N_11123);
nor U11348 (N_11348,N_11005,N_11093);
and U11349 (N_11349,N_11177,N_11008);
nor U11350 (N_11350,N_11064,N_11246);
and U11351 (N_11351,N_11074,N_11114);
or U11352 (N_11352,N_11143,N_11021);
or U11353 (N_11353,N_11121,N_11073);
or U11354 (N_11354,N_11109,N_11053);
nor U11355 (N_11355,N_11084,N_11195);
xor U11356 (N_11356,N_11187,N_11182);
xnor U11357 (N_11357,N_11065,N_11189);
nor U11358 (N_11358,N_11106,N_11032);
xor U11359 (N_11359,N_11243,N_11127);
or U11360 (N_11360,N_11087,N_11094);
nand U11361 (N_11361,N_11117,N_11126);
nor U11362 (N_11362,N_11172,N_11226);
xor U11363 (N_11363,N_11025,N_11136);
nor U11364 (N_11364,N_11034,N_11066);
or U11365 (N_11365,N_11026,N_11108);
and U11366 (N_11366,N_11039,N_11028);
or U11367 (N_11367,N_11186,N_11012);
and U11368 (N_11368,N_11099,N_11068);
xor U11369 (N_11369,N_11163,N_11188);
nand U11370 (N_11370,N_11016,N_11179);
and U11371 (N_11371,N_11209,N_11210);
xnor U11372 (N_11372,N_11101,N_11102);
xnor U11373 (N_11373,N_11214,N_11236);
nand U11374 (N_11374,N_11192,N_11038);
nand U11375 (N_11375,N_11189,N_11036);
and U11376 (N_11376,N_11172,N_11150);
and U11377 (N_11377,N_11012,N_11158);
or U11378 (N_11378,N_11222,N_11135);
xnor U11379 (N_11379,N_11045,N_11077);
and U11380 (N_11380,N_11191,N_11160);
xnor U11381 (N_11381,N_11247,N_11170);
and U11382 (N_11382,N_11111,N_11149);
and U11383 (N_11383,N_11220,N_11047);
and U11384 (N_11384,N_11181,N_11140);
xnor U11385 (N_11385,N_11144,N_11244);
nand U11386 (N_11386,N_11171,N_11193);
nand U11387 (N_11387,N_11125,N_11214);
or U11388 (N_11388,N_11219,N_11039);
xor U11389 (N_11389,N_11008,N_11229);
and U11390 (N_11390,N_11141,N_11228);
nor U11391 (N_11391,N_11008,N_11046);
and U11392 (N_11392,N_11094,N_11029);
nand U11393 (N_11393,N_11212,N_11068);
xor U11394 (N_11394,N_11148,N_11212);
and U11395 (N_11395,N_11072,N_11216);
nand U11396 (N_11396,N_11180,N_11093);
nand U11397 (N_11397,N_11095,N_11029);
nor U11398 (N_11398,N_11089,N_11237);
nand U11399 (N_11399,N_11233,N_11029);
xor U11400 (N_11400,N_11004,N_11053);
and U11401 (N_11401,N_11210,N_11131);
and U11402 (N_11402,N_11036,N_11108);
and U11403 (N_11403,N_11218,N_11223);
and U11404 (N_11404,N_11097,N_11187);
xnor U11405 (N_11405,N_11151,N_11169);
and U11406 (N_11406,N_11049,N_11013);
or U11407 (N_11407,N_11083,N_11108);
xnor U11408 (N_11408,N_11147,N_11214);
xnor U11409 (N_11409,N_11050,N_11016);
or U11410 (N_11410,N_11125,N_11022);
and U11411 (N_11411,N_11037,N_11029);
nand U11412 (N_11412,N_11167,N_11048);
xor U11413 (N_11413,N_11041,N_11113);
or U11414 (N_11414,N_11003,N_11181);
nand U11415 (N_11415,N_11178,N_11222);
nand U11416 (N_11416,N_11173,N_11131);
xor U11417 (N_11417,N_11151,N_11100);
nand U11418 (N_11418,N_11242,N_11238);
nand U11419 (N_11419,N_11010,N_11089);
and U11420 (N_11420,N_11179,N_11030);
or U11421 (N_11421,N_11218,N_11153);
or U11422 (N_11422,N_11085,N_11216);
nor U11423 (N_11423,N_11131,N_11241);
nor U11424 (N_11424,N_11234,N_11081);
nor U11425 (N_11425,N_11065,N_11130);
or U11426 (N_11426,N_11055,N_11098);
nand U11427 (N_11427,N_11078,N_11181);
nor U11428 (N_11428,N_11005,N_11103);
or U11429 (N_11429,N_11196,N_11141);
nand U11430 (N_11430,N_11166,N_11117);
nor U11431 (N_11431,N_11249,N_11015);
nor U11432 (N_11432,N_11181,N_11225);
or U11433 (N_11433,N_11092,N_11049);
nand U11434 (N_11434,N_11098,N_11057);
nand U11435 (N_11435,N_11086,N_11005);
nor U11436 (N_11436,N_11227,N_11117);
nand U11437 (N_11437,N_11013,N_11196);
and U11438 (N_11438,N_11046,N_11097);
nand U11439 (N_11439,N_11060,N_11021);
xor U11440 (N_11440,N_11072,N_11170);
nand U11441 (N_11441,N_11022,N_11159);
nor U11442 (N_11442,N_11161,N_11042);
and U11443 (N_11443,N_11054,N_11122);
nand U11444 (N_11444,N_11130,N_11221);
xor U11445 (N_11445,N_11105,N_11154);
or U11446 (N_11446,N_11096,N_11137);
or U11447 (N_11447,N_11148,N_11121);
or U11448 (N_11448,N_11133,N_11139);
and U11449 (N_11449,N_11176,N_11243);
nand U11450 (N_11450,N_11094,N_11020);
nor U11451 (N_11451,N_11042,N_11238);
and U11452 (N_11452,N_11176,N_11027);
or U11453 (N_11453,N_11144,N_11140);
nand U11454 (N_11454,N_11214,N_11022);
nor U11455 (N_11455,N_11244,N_11005);
nor U11456 (N_11456,N_11021,N_11044);
or U11457 (N_11457,N_11069,N_11019);
and U11458 (N_11458,N_11235,N_11151);
or U11459 (N_11459,N_11223,N_11000);
nand U11460 (N_11460,N_11003,N_11117);
or U11461 (N_11461,N_11072,N_11008);
nor U11462 (N_11462,N_11075,N_11226);
and U11463 (N_11463,N_11013,N_11168);
xnor U11464 (N_11464,N_11109,N_11102);
xnor U11465 (N_11465,N_11134,N_11136);
xnor U11466 (N_11466,N_11064,N_11043);
nand U11467 (N_11467,N_11104,N_11107);
nand U11468 (N_11468,N_11075,N_11052);
and U11469 (N_11469,N_11202,N_11019);
and U11470 (N_11470,N_11217,N_11171);
nand U11471 (N_11471,N_11105,N_11033);
nor U11472 (N_11472,N_11199,N_11035);
and U11473 (N_11473,N_11140,N_11220);
xor U11474 (N_11474,N_11159,N_11240);
and U11475 (N_11475,N_11087,N_11044);
and U11476 (N_11476,N_11125,N_11179);
or U11477 (N_11477,N_11131,N_11181);
xor U11478 (N_11478,N_11131,N_11011);
nor U11479 (N_11479,N_11034,N_11168);
nand U11480 (N_11480,N_11211,N_11184);
nor U11481 (N_11481,N_11041,N_11043);
nor U11482 (N_11482,N_11234,N_11051);
xor U11483 (N_11483,N_11069,N_11080);
nand U11484 (N_11484,N_11183,N_11055);
xnor U11485 (N_11485,N_11192,N_11052);
and U11486 (N_11486,N_11169,N_11099);
nor U11487 (N_11487,N_11230,N_11206);
nand U11488 (N_11488,N_11013,N_11116);
nor U11489 (N_11489,N_11038,N_11181);
or U11490 (N_11490,N_11141,N_11088);
nor U11491 (N_11491,N_11233,N_11182);
nand U11492 (N_11492,N_11032,N_11037);
nand U11493 (N_11493,N_11106,N_11044);
or U11494 (N_11494,N_11149,N_11171);
xnor U11495 (N_11495,N_11081,N_11090);
nand U11496 (N_11496,N_11060,N_11049);
nand U11497 (N_11497,N_11247,N_11217);
nand U11498 (N_11498,N_11201,N_11223);
nand U11499 (N_11499,N_11206,N_11089);
xor U11500 (N_11500,N_11327,N_11404);
nor U11501 (N_11501,N_11411,N_11345);
nor U11502 (N_11502,N_11479,N_11308);
and U11503 (N_11503,N_11390,N_11459);
and U11504 (N_11504,N_11273,N_11317);
nor U11505 (N_11505,N_11460,N_11357);
xor U11506 (N_11506,N_11360,N_11480);
or U11507 (N_11507,N_11320,N_11375);
nor U11508 (N_11508,N_11292,N_11484);
xor U11509 (N_11509,N_11420,N_11408);
or U11510 (N_11510,N_11286,N_11359);
and U11511 (N_11511,N_11306,N_11337);
nor U11512 (N_11512,N_11435,N_11425);
nand U11513 (N_11513,N_11302,N_11464);
xnor U11514 (N_11514,N_11407,N_11295);
or U11515 (N_11515,N_11467,N_11280);
nand U11516 (N_11516,N_11437,N_11453);
xnor U11517 (N_11517,N_11285,N_11356);
or U11518 (N_11518,N_11284,N_11419);
nand U11519 (N_11519,N_11254,N_11489);
and U11520 (N_11520,N_11454,N_11331);
nor U11521 (N_11521,N_11444,N_11499);
xnor U11522 (N_11522,N_11393,N_11324);
nor U11523 (N_11523,N_11279,N_11386);
xnor U11524 (N_11524,N_11450,N_11342);
nand U11525 (N_11525,N_11353,N_11270);
nor U11526 (N_11526,N_11255,N_11352);
nor U11527 (N_11527,N_11329,N_11333);
nand U11528 (N_11528,N_11322,N_11347);
and U11529 (N_11529,N_11442,N_11487);
xnor U11530 (N_11530,N_11478,N_11415);
nor U11531 (N_11531,N_11335,N_11341);
nor U11532 (N_11532,N_11281,N_11271);
and U11533 (N_11533,N_11349,N_11438);
nand U11534 (N_11534,N_11429,N_11446);
xor U11535 (N_11535,N_11447,N_11492);
and U11536 (N_11536,N_11339,N_11498);
and U11537 (N_11537,N_11410,N_11465);
nand U11538 (N_11538,N_11294,N_11448);
nor U11539 (N_11539,N_11326,N_11276);
xor U11540 (N_11540,N_11401,N_11430);
nor U11541 (N_11541,N_11323,N_11259);
or U11542 (N_11542,N_11421,N_11253);
or U11543 (N_11543,N_11431,N_11298);
or U11544 (N_11544,N_11458,N_11378);
xor U11545 (N_11545,N_11367,N_11383);
or U11546 (N_11546,N_11481,N_11427);
nand U11547 (N_11547,N_11348,N_11377);
xor U11548 (N_11548,N_11371,N_11256);
or U11549 (N_11549,N_11334,N_11261);
and U11550 (N_11550,N_11396,N_11391);
xnor U11551 (N_11551,N_11372,N_11440);
or U11552 (N_11552,N_11423,N_11387);
and U11553 (N_11553,N_11382,N_11290);
nand U11554 (N_11554,N_11397,N_11346);
or U11555 (N_11555,N_11486,N_11265);
nor U11556 (N_11556,N_11466,N_11417);
and U11557 (N_11557,N_11304,N_11332);
and U11558 (N_11558,N_11260,N_11385);
xor U11559 (N_11559,N_11409,N_11312);
and U11560 (N_11560,N_11328,N_11433);
nor U11561 (N_11561,N_11491,N_11314);
or U11562 (N_11562,N_11282,N_11267);
nand U11563 (N_11563,N_11451,N_11363);
and U11564 (N_11564,N_11403,N_11493);
nand U11565 (N_11565,N_11266,N_11405);
nor U11566 (N_11566,N_11288,N_11398);
nor U11567 (N_11567,N_11457,N_11496);
xor U11568 (N_11568,N_11384,N_11283);
or U11569 (N_11569,N_11272,N_11293);
nor U11570 (N_11570,N_11399,N_11380);
xor U11571 (N_11571,N_11354,N_11251);
xnor U11572 (N_11572,N_11316,N_11370);
and U11573 (N_11573,N_11414,N_11452);
nor U11574 (N_11574,N_11319,N_11264);
or U11575 (N_11575,N_11497,N_11469);
xor U11576 (N_11576,N_11389,N_11388);
and U11577 (N_11577,N_11488,N_11258);
xnor U11578 (N_11578,N_11418,N_11311);
nand U11579 (N_11579,N_11278,N_11340);
and U11580 (N_11580,N_11362,N_11351);
xor U11581 (N_11581,N_11369,N_11455);
nand U11582 (N_11582,N_11344,N_11374);
xnor U11583 (N_11583,N_11392,N_11318);
and U11584 (N_11584,N_11474,N_11468);
and U11585 (N_11585,N_11343,N_11263);
and U11586 (N_11586,N_11301,N_11313);
and U11587 (N_11587,N_11445,N_11355);
nor U11588 (N_11588,N_11424,N_11416);
nand U11589 (N_11589,N_11432,N_11422);
nand U11590 (N_11590,N_11366,N_11287);
nand U11591 (N_11591,N_11381,N_11321);
or U11592 (N_11592,N_11494,N_11461);
and U11593 (N_11593,N_11307,N_11483);
nor U11594 (N_11594,N_11330,N_11441);
nor U11595 (N_11595,N_11365,N_11413);
and U11596 (N_11596,N_11262,N_11275);
nand U11597 (N_11597,N_11305,N_11368);
xor U11598 (N_11598,N_11472,N_11268);
nor U11599 (N_11599,N_11379,N_11473);
xnor U11600 (N_11600,N_11361,N_11470);
and U11601 (N_11601,N_11364,N_11289);
nor U11602 (N_11602,N_11426,N_11297);
or U11603 (N_11603,N_11338,N_11475);
and U11604 (N_11604,N_11299,N_11257);
nor U11605 (N_11605,N_11309,N_11394);
nand U11606 (N_11606,N_11315,N_11310);
or U11607 (N_11607,N_11373,N_11428);
or U11608 (N_11608,N_11358,N_11456);
nor U11609 (N_11609,N_11436,N_11495);
or U11610 (N_11610,N_11274,N_11269);
nand U11611 (N_11611,N_11462,N_11477);
nor U11612 (N_11612,N_11250,N_11463);
nand U11613 (N_11613,N_11350,N_11412);
nand U11614 (N_11614,N_11395,N_11277);
nor U11615 (N_11615,N_11406,N_11402);
nor U11616 (N_11616,N_11336,N_11449);
xor U11617 (N_11617,N_11439,N_11485);
xor U11618 (N_11618,N_11476,N_11443);
nor U11619 (N_11619,N_11376,N_11291);
nor U11620 (N_11620,N_11252,N_11471);
nand U11621 (N_11621,N_11490,N_11296);
or U11622 (N_11622,N_11300,N_11434);
and U11623 (N_11623,N_11400,N_11482);
and U11624 (N_11624,N_11303,N_11325);
nor U11625 (N_11625,N_11460,N_11459);
or U11626 (N_11626,N_11420,N_11445);
and U11627 (N_11627,N_11397,N_11306);
xnor U11628 (N_11628,N_11354,N_11451);
and U11629 (N_11629,N_11260,N_11442);
xor U11630 (N_11630,N_11489,N_11438);
and U11631 (N_11631,N_11402,N_11395);
and U11632 (N_11632,N_11498,N_11349);
xnor U11633 (N_11633,N_11351,N_11475);
xor U11634 (N_11634,N_11402,N_11272);
xor U11635 (N_11635,N_11491,N_11262);
or U11636 (N_11636,N_11478,N_11349);
xor U11637 (N_11637,N_11316,N_11440);
nor U11638 (N_11638,N_11425,N_11291);
and U11639 (N_11639,N_11308,N_11257);
nor U11640 (N_11640,N_11412,N_11393);
nand U11641 (N_11641,N_11436,N_11472);
nand U11642 (N_11642,N_11288,N_11402);
nand U11643 (N_11643,N_11358,N_11407);
nand U11644 (N_11644,N_11391,N_11320);
nor U11645 (N_11645,N_11495,N_11322);
nand U11646 (N_11646,N_11427,N_11260);
or U11647 (N_11647,N_11254,N_11400);
xor U11648 (N_11648,N_11280,N_11383);
and U11649 (N_11649,N_11382,N_11373);
nor U11650 (N_11650,N_11332,N_11442);
nand U11651 (N_11651,N_11350,N_11447);
nand U11652 (N_11652,N_11445,N_11397);
nor U11653 (N_11653,N_11296,N_11381);
and U11654 (N_11654,N_11429,N_11447);
nor U11655 (N_11655,N_11468,N_11330);
nor U11656 (N_11656,N_11335,N_11291);
nor U11657 (N_11657,N_11363,N_11473);
nand U11658 (N_11658,N_11317,N_11487);
and U11659 (N_11659,N_11416,N_11327);
or U11660 (N_11660,N_11304,N_11416);
xor U11661 (N_11661,N_11336,N_11377);
nor U11662 (N_11662,N_11308,N_11301);
nor U11663 (N_11663,N_11423,N_11256);
nand U11664 (N_11664,N_11386,N_11447);
nand U11665 (N_11665,N_11341,N_11293);
xnor U11666 (N_11666,N_11485,N_11454);
nor U11667 (N_11667,N_11408,N_11256);
xnor U11668 (N_11668,N_11307,N_11487);
and U11669 (N_11669,N_11405,N_11363);
and U11670 (N_11670,N_11468,N_11302);
xnor U11671 (N_11671,N_11369,N_11335);
and U11672 (N_11672,N_11437,N_11406);
nor U11673 (N_11673,N_11449,N_11250);
nand U11674 (N_11674,N_11477,N_11408);
or U11675 (N_11675,N_11298,N_11327);
xor U11676 (N_11676,N_11267,N_11474);
or U11677 (N_11677,N_11250,N_11357);
and U11678 (N_11678,N_11362,N_11333);
nand U11679 (N_11679,N_11385,N_11380);
xnor U11680 (N_11680,N_11323,N_11295);
and U11681 (N_11681,N_11415,N_11432);
xor U11682 (N_11682,N_11358,N_11315);
or U11683 (N_11683,N_11345,N_11441);
xor U11684 (N_11684,N_11378,N_11322);
and U11685 (N_11685,N_11439,N_11440);
or U11686 (N_11686,N_11252,N_11349);
nor U11687 (N_11687,N_11479,N_11252);
nor U11688 (N_11688,N_11417,N_11436);
or U11689 (N_11689,N_11397,N_11470);
nand U11690 (N_11690,N_11471,N_11434);
nor U11691 (N_11691,N_11269,N_11287);
xor U11692 (N_11692,N_11446,N_11456);
xor U11693 (N_11693,N_11499,N_11295);
and U11694 (N_11694,N_11346,N_11427);
nand U11695 (N_11695,N_11311,N_11287);
nand U11696 (N_11696,N_11481,N_11448);
nand U11697 (N_11697,N_11281,N_11497);
or U11698 (N_11698,N_11366,N_11496);
or U11699 (N_11699,N_11420,N_11365);
xor U11700 (N_11700,N_11489,N_11295);
xnor U11701 (N_11701,N_11333,N_11454);
nand U11702 (N_11702,N_11446,N_11434);
or U11703 (N_11703,N_11318,N_11325);
and U11704 (N_11704,N_11322,N_11297);
nand U11705 (N_11705,N_11460,N_11329);
nor U11706 (N_11706,N_11396,N_11458);
nand U11707 (N_11707,N_11384,N_11275);
nand U11708 (N_11708,N_11394,N_11257);
xor U11709 (N_11709,N_11299,N_11432);
xor U11710 (N_11710,N_11271,N_11400);
and U11711 (N_11711,N_11260,N_11428);
nor U11712 (N_11712,N_11470,N_11274);
nor U11713 (N_11713,N_11272,N_11367);
xnor U11714 (N_11714,N_11407,N_11419);
and U11715 (N_11715,N_11426,N_11379);
nor U11716 (N_11716,N_11364,N_11471);
xnor U11717 (N_11717,N_11282,N_11452);
nor U11718 (N_11718,N_11473,N_11362);
nor U11719 (N_11719,N_11361,N_11374);
nor U11720 (N_11720,N_11317,N_11345);
nor U11721 (N_11721,N_11326,N_11353);
xnor U11722 (N_11722,N_11268,N_11482);
xor U11723 (N_11723,N_11464,N_11413);
nand U11724 (N_11724,N_11319,N_11453);
or U11725 (N_11725,N_11483,N_11271);
nand U11726 (N_11726,N_11311,N_11434);
xor U11727 (N_11727,N_11353,N_11424);
xor U11728 (N_11728,N_11461,N_11485);
and U11729 (N_11729,N_11364,N_11323);
and U11730 (N_11730,N_11311,N_11315);
and U11731 (N_11731,N_11496,N_11293);
nand U11732 (N_11732,N_11330,N_11440);
and U11733 (N_11733,N_11493,N_11266);
nand U11734 (N_11734,N_11499,N_11305);
or U11735 (N_11735,N_11347,N_11486);
and U11736 (N_11736,N_11319,N_11438);
and U11737 (N_11737,N_11451,N_11254);
xnor U11738 (N_11738,N_11349,N_11423);
nor U11739 (N_11739,N_11400,N_11383);
nand U11740 (N_11740,N_11322,N_11277);
nor U11741 (N_11741,N_11404,N_11316);
or U11742 (N_11742,N_11472,N_11467);
nor U11743 (N_11743,N_11357,N_11488);
and U11744 (N_11744,N_11481,N_11252);
xnor U11745 (N_11745,N_11484,N_11271);
xnor U11746 (N_11746,N_11389,N_11393);
xnor U11747 (N_11747,N_11438,N_11368);
nor U11748 (N_11748,N_11287,N_11270);
nor U11749 (N_11749,N_11403,N_11318);
nand U11750 (N_11750,N_11624,N_11641);
nand U11751 (N_11751,N_11568,N_11533);
or U11752 (N_11752,N_11721,N_11591);
and U11753 (N_11753,N_11714,N_11674);
nor U11754 (N_11754,N_11733,N_11740);
xnor U11755 (N_11755,N_11739,N_11571);
and U11756 (N_11756,N_11693,N_11622);
and U11757 (N_11757,N_11692,N_11700);
or U11758 (N_11758,N_11734,N_11630);
and U11759 (N_11759,N_11749,N_11648);
or U11760 (N_11760,N_11653,N_11594);
or U11761 (N_11761,N_11511,N_11500);
and U11762 (N_11762,N_11650,N_11603);
or U11763 (N_11763,N_11747,N_11689);
and U11764 (N_11764,N_11561,N_11703);
xnor U11765 (N_11765,N_11556,N_11608);
xor U11766 (N_11766,N_11679,N_11616);
nor U11767 (N_11767,N_11558,N_11553);
nor U11768 (N_11768,N_11644,N_11663);
nor U11769 (N_11769,N_11620,N_11623);
and U11770 (N_11770,N_11519,N_11720);
and U11771 (N_11771,N_11547,N_11612);
xnor U11772 (N_11772,N_11598,N_11711);
or U11773 (N_11773,N_11705,N_11557);
nor U11774 (N_11774,N_11523,N_11536);
or U11775 (N_11775,N_11617,N_11570);
and U11776 (N_11776,N_11567,N_11719);
or U11777 (N_11777,N_11508,N_11618);
xnor U11778 (N_11778,N_11701,N_11518);
or U11779 (N_11779,N_11673,N_11524);
nor U11780 (N_11780,N_11710,N_11666);
nand U11781 (N_11781,N_11602,N_11636);
xnor U11782 (N_11782,N_11527,N_11580);
or U11783 (N_11783,N_11549,N_11731);
nand U11784 (N_11784,N_11708,N_11681);
xor U11785 (N_11785,N_11569,N_11715);
nand U11786 (N_11786,N_11626,N_11716);
or U11787 (N_11787,N_11590,N_11610);
xor U11788 (N_11788,N_11619,N_11668);
nand U11789 (N_11789,N_11564,N_11707);
xnor U11790 (N_11790,N_11676,N_11577);
or U11791 (N_11791,N_11690,N_11722);
or U11792 (N_11792,N_11537,N_11584);
nand U11793 (N_11793,N_11607,N_11670);
or U11794 (N_11794,N_11504,N_11639);
nor U11795 (N_11795,N_11604,N_11545);
xnor U11796 (N_11796,N_11588,N_11565);
or U11797 (N_11797,N_11677,N_11509);
or U11798 (N_11798,N_11551,N_11534);
or U11799 (N_11799,N_11600,N_11736);
or U11800 (N_11800,N_11633,N_11709);
and U11801 (N_11801,N_11697,N_11682);
nand U11802 (N_11802,N_11548,N_11742);
nand U11803 (N_11803,N_11543,N_11559);
nor U11804 (N_11804,N_11506,N_11688);
xor U11805 (N_11805,N_11525,N_11593);
nor U11806 (N_11806,N_11660,N_11686);
nand U11807 (N_11807,N_11573,N_11625);
and U11808 (N_11808,N_11637,N_11729);
xor U11809 (N_11809,N_11513,N_11542);
xor U11810 (N_11810,N_11685,N_11541);
and U11811 (N_11811,N_11581,N_11582);
and U11812 (N_11812,N_11635,N_11520);
nand U11813 (N_11813,N_11638,N_11704);
and U11814 (N_11814,N_11535,N_11662);
and U11815 (N_11815,N_11694,N_11683);
or U11816 (N_11816,N_11579,N_11655);
or U11817 (N_11817,N_11611,N_11601);
nand U11818 (N_11818,N_11587,N_11727);
xnor U11819 (N_11819,N_11738,N_11669);
and U11820 (N_11820,N_11672,N_11578);
xor U11821 (N_11821,N_11628,N_11656);
and U11822 (N_11822,N_11671,N_11646);
and U11823 (N_11823,N_11664,N_11732);
or U11824 (N_11824,N_11661,N_11503);
and U11825 (N_11825,N_11631,N_11526);
xor U11826 (N_11826,N_11546,N_11658);
xor U11827 (N_11827,N_11657,N_11654);
xor U11828 (N_11828,N_11699,N_11691);
or U11829 (N_11829,N_11507,N_11675);
xor U11830 (N_11830,N_11552,N_11560);
or U11831 (N_11831,N_11634,N_11647);
or U11832 (N_11832,N_11632,N_11605);
nor U11833 (N_11833,N_11550,N_11576);
xor U11834 (N_11834,N_11665,N_11696);
or U11835 (N_11835,N_11589,N_11514);
xnor U11836 (N_11836,N_11725,N_11515);
nor U11837 (N_11837,N_11643,N_11599);
and U11838 (N_11838,N_11712,N_11609);
nand U11839 (N_11839,N_11528,N_11583);
nand U11840 (N_11840,N_11615,N_11717);
xor U11841 (N_11841,N_11743,N_11586);
or U11842 (N_11842,N_11574,N_11735);
or U11843 (N_11843,N_11516,N_11510);
or U11844 (N_11844,N_11563,N_11521);
nand U11845 (N_11845,N_11649,N_11585);
or U11846 (N_11846,N_11531,N_11695);
or U11847 (N_11847,N_11621,N_11572);
nand U11848 (N_11848,N_11726,N_11517);
nor U11849 (N_11849,N_11505,N_11746);
nor U11850 (N_11850,N_11554,N_11724);
nor U11851 (N_11851,N_11614,N_11566);
xor U11852 (N_11852,N_11713,N_11640);
nand U11853 (N_11853,N_11748,N_11737);
nand U11854 (N_11854,N_11741,N_11502);
nor U11855 (N_11855,N_11698,N_11744);
or U11856 (N_11856,N_11659,N_11540);
xor U11857 (N_11857,N_11522,N_11684);
or U11858 (N_11858,N_11629,N_11529);
xnor U11859 (N_11859,N_11530,N_11718);
and U11860 (N_11860,N_11613,N_11687);
nor U11861 (N_11861,N_11680,N_11651);
and U11862 (N_11862,N_11597,N_11595);
xor U11863 (N_11863,N_11596,N_11606);
or U11864 (N_11864,N_11575,N_11730);
nand U11865 (N_11865,N_11539,N_11652);
nand U11866 (N_11866,N_11501,N_11627);
and U11867 (N_11867,N_11706,N_11555);
and U11868 (N_11868,N_11702,N_11723);
and U11869 (N_11869,N_11544,N_11562);
or U11870 (N_11870,N_11728,N_11645);
xnor U11871 (N_11871,N_11592,N_11512);
or U11872 (N_11872,N_11667,N_11538);
or U11873 (N_11873,N_11745,N_11642);
or U11874 (N_11874,N_11532,N_11678);
or U11875 (N_11875,N_11736,N_11586);
xor U11876 (N_11876,N_11672,N_11656);
nor U11877 (N_11877,N_11676,N_11519);
nand U11878 (N_11878,N_11542,N_11713);
or U11879 (N_11879,N_11734,N_11532);
nor U11880 (N_11880,N_11515,N_11596);
and U11881 (N_11881,N_11721,N_11741);
nor U11882 (N_11882,N_11518,N_11616);
nand U11883 (N_11883,N_11629,N_11546);
or U11884 (N_11884,N_11560,N_11581);
nand U11885 (N_11885,N_11744,N_11643);
or U11886 (N_11886,N_11539,N_11605);
or U11887 (N_11887,N_11565,N_11637);
nand U11888 (N_11888,N_11658,N_11648);
and U11889 (N_11889,N_11510,N_11749);
nand U11890 (N_11890,N_11559,N_11655);
and U11891 (N_11891,N_11515,N_11699);
xor U11892 (N_11892,N_11663,N_11671);
or U11893 (N_11893,N_11748,N_11657);
nor U11894 (N_11894,N_11514,N_11663);
nor U11895 (N_11895,N_11717,N_11537);
and U11896 (N_11896,N_11694,N_11686);
and U11897 (N_11897,N_11588,N_11519);
xor U11898 (N_11898,N_11555,N_11700);
nand U11899 (N_11899,N_11736,N_11548);
nor U11900 (N_11900,N_11651,N_11712);
xor U11901 (N_11901,N_11581,N_11666);
and U11902 (N_11902,N_11561,N_11642);
nand U11903 (N_11903,N_11532,N_11565);
nor U11904 (N_11904,N_11681,N_11658);
and U11905 (N_11905,N_11663,N_11629);
and U11906 (N_11906,N_11623,N_11658);
xor U11907 (N_11907,N_11711,N_11543);
or U11908 (N_11908,N_11697,N_11599);
and U11909 (N_11909,N_11553,N_11578);
nand U11910 (N_11910,N_11734,N_11597);
or U11911 (N_11911,N_11641,N_11698);
and U11912 (N_11912,N_11668,N_11718);
nor U11913 (N_11913,N_11738,N_11634);
xnor U11914 (N_11914,N_11678,N_11697);
xor U11915 (N_11915,N_11639,N_11701);
and U11916 (N_11916,N_11696,N_11642);
xor U11917 (N_11917,N_11725,N_11561);
xor U11918 (N_11918,N_11535,N_11676);
or U11919 (N_11919,N_11626,N_11533);
or U11920 (N_11920,N_11608,N_11590);
xor U11921 (N_11921,N_11638,N_11727);
xnor U11922 (N_11922,N_11557,N_11679);
and U11923 (N_11923,N_11676,N_11629);
nand U11924 (N_11924,N_11713,N_11626);
nor U11925 (N_11925,N_11742,N_11625);
and U11926 (N_11926,N_11719,N_11548);
or U11927 (N_11927,N_11571,N_11572);
nand U11928 (N_11928,N_11508,N_11687);
and U11929 (N_11929,N_11600,N_11623);
and U11930 (N_11930,N_11720,N_11597);
and U11931 (N_11931,N_11670,N_11737);
nor U11932 (N_11932,N_11525,N_11647);
or U11933 (N_11933,N_11651,N_11613);
nand U11934 (N_11934,N_11599,N_11712);
xor U11935 (N_11935,N_11664,N_11724);
nor U11936 (N_11936,N_11729,N_11746);
nand U11937 (N_11937,N_11628,N_11654);
nand U11938 (N_11938,N_11594,N_11726);
or U11939 (N_11939,N_11596,N_11526);
nor U11940 (N_11940,N_11685,N_11506);
and U11941 (N_11941,N_11509,N_11664);
and U11942 (N_11942,N_11559,N_11577);
xnor U11943 (N_11943,N_11675,N_11648);
and U11944 (N_11944,N_11606,N_11745);
or U11945 (N_11945,N_11675,N_11692);
nor U11946 (N_11946,N_11626,N_11507);
nor U11947 (N_11947,N_11551,N_11597);
nand U11948 (N_11948,N_11717,N_11625);
or U11949 (N_11949,N_11552,N_11570);
nand U11950 (N_11950,N_11637,N_11591);
and U11951 (N_11951,N_11676,N_11575);
xnor U11952 (N_11952,N_11659,N_11646);
nand U11953 (N_11953,N_11550,N_11549);
nand U11954 (N_11954,N_11625,N_11737);
nand U11955 (N_11955,N_11725,N_11638);
and U11956 (N_11956,N_11529,N_11701);
nor U11957 (N_11957,N_11576,N_11557);
and U11958 (N_11958,N_11746,N_11583);
and U11959 (N_11959,N_11510,N_11716);
nand U11960 (N_11960,N_11683,N_11557);
or U11961 (N_11961,N_11709,N_11540);
or U11962 (N_11962,N_11612,N_11598);
nor U11963 (N_11963,N_11666,N_11588);
and U11964 (N_11964,N_11725,N_11548);
and U11965 (N_11965,N_11741,N_11700);
or U11966 (N_11966,N_11670,N_11727);
xnor U11967 (N_11967,N_11749,N_11624);
nand U11968 (N_11968,N_11555,N_11576);
nand U11969 (N_11969,N_11567,N_11606);
nand U11970 (N_11970,N_11581,N_11591);
xor U11971 (N_11971,N_11585,N_11689);
and U11972 (N_11972,N_11629,N_11559);
and U11973 (N_11973,N_11574,N_11601);
and U11974 (N_11974,N_11624,N_11518);
nor U11975 (N_11975,N_11712,N_11600);
xnor U11976 (N_11976,N_11720,N_11543);
xnor U11977 (N_11977,N_11635,N_11656);
nor U11978 (N_11978,N_11570,N_11688);
or U11979 (N_11979,N_11736,N_11530);
nand U11980 (N_11980,N_11594,N_11583);
nor U11981 (N_11981,N_11690,N_11749);
nand U11982 (N_11982,N_11639,N_11717);
xor U11983 (N_11983,N_11692,N_11505);
nand U11984 (N_11984,N_11506,N_11592);
nand U11985 (N_11985,N_11509,N_11528);
xnor U11986 (N_11986,N_11592,N_11500);
and U11987 (N_11987,N_11584,N_11691);
xor U11988 (N_11988,N_11693,N_11623);
xor U11989 (N_11989,N_11511,N_11543);
nand U11990 (N_11990,N_11704,N_11749);
nand U11991 (N_11991,N_11637,N_11579);
or U11992 (N_11992,N_11578,N_11734);
xnor U11993 (N_11993,N_11602,N_11536);
xor U11994 (N_11994,N_11581,N_11614);
xnor U11995 (N_11995,N_11684,N_11690);
or U11996 (N_11996,N_11632,N_11531);
or U11997 (N_11997,N_11640,N_11675);
nor U11998 (N_11998,N_11522,N_11592);
xnor U11999 (N_11999,N_11575,N_11526);
or U12000 (N_12000,N_11915,N_11772);
or U12001 (N_12001,N_11920,N_11836);
nor U12002 (N_12002,N_11906,N_11794);
or U12003 (N_12003,N_11857,N_11851);
and U12004 (N_12004,N_11888,N_11829);
and U12005 (N_12005,N_11973,N_11943);
nand U12006 (N_12006,N_11872,N_11776);
or U12007 (N_12007,N_11764,N_11948);
and U12008 (N_12008,N_11890,N_11899);
and U12009 (N_12009,N_11803,N_11775);
and U12010 (N_12010,N_11752,N_11821);
nor U12011 (N_12011,N_11918,N_11870);
nand U12012 (N_12012,N_11937,N_11986);
xor U12013 (N_12013,N_11841,N_11991);
or U12014 (N_12014,N_11863,N_11939);
nand U12015 (N_12015,N_11839,N_11827);
nand U12016 (N_12016,N_11987,N_11818);
nand U12017 (N_12017,N_11756,N_11981);
nand U12018 (N_12018,N_11842,N_11945);
nor U12019 (N_12019,N_11860,N_11902);
or U12020 (N_12020,N_11966,N_11784);
or U12021 (N_12021,N_11944,N_11799);
and U12022 (N_12022,N_11810,N_11858);
nand U12023 (N_12023,N_11961,N_11787);
xnor U12024 (N_12024,N_11903,N_11934);
nand U12025 (N_12025,N_11993,N_11876);
nor U12026 (N_12026,N_11874,N_11958);
nand U12027 (N_12027,N_11814,N_11909);
xor U12028 (N_12028,N_11845,N_11941);
or U12029 (N_12029,N_11761,N_11817);
xnor U12030 (N_12030,N_11954,N_11795);
xor U12031 (N_12031,N_11807,N_11826);
or U12032 (N_12032,N_11896,N_11780);
nand U12033 (N_12033,N_11820,N_11783);
nor U12034 (N_12034,N_11854,N_11975);
xnor U12035 (N_12035,N_11886,N_11869);
nand U12036 (N_12036,N_11805,N_11861);
nand U12037 (N_12037,N_11901,N_11751);
or U12038 (N_12038,N_11949,N_11788);
xnor U12039 (N_12039,N_11924,N_11999);
or U12040 (N_12040,N_11984,N_11925);
and U12041 (N_12041,N_11959,N_11878);
xnor U12042 (N_12042,N_11983,N_11773);
and U12043 (N_12043,N_11768,N_11913);
xnor U12044 (N_12044,N_11792,N_11955);
nand U12045 (N_12045,N_11992,N_11859);
nor U12046 (N_12046,N_11759,N_11850);
nand U12047 (N_12047,N_11911,N_11848);
or U12048 (N_12048,N_11804,N_11942);
and U12049 (N_12049,N_11813,N_11774);
nand U12050 (N_12050,N_11977,N_11840);
xor U12051 (N_12051,N_11905,N_11976);
xnor U12052 (N_12052,N_11957,N_11847);
or U12053 (N_12053,N_11968,N_11815);
xor U12054 (N_12054,N_11912,N_11762);
or U12055 (N_12055,N_11811,N_11835);
or U12056 (N_12056,N_11947,N_11871);
xor U12057 (N_12057,N_11929,N_11812);
and U12058 (N_12058,N_11793,N_11982);
nor U12059 (N_12059,N_11830,N_11960);
nand U12060 (N_12060,N_11769,N_11972);
or U12061 (N_12061,N_11940,N_11921);
nand U12062 (N_12062,N_11952,N_11823);
nand U12063 (N_12063,N_11922,N_11928);
xnor U12064 (N_12064,N_11825,N_11962);
xor U12065 (N_12065,N_11831,N_11882);
nand U12066 (N_12066,N_11953,N_11971);
nor U12067 (N_12067,N_11907,N_11765);
nand U12068 (N_12068,N_11758,N_11837);
nand U12069 (N_12069,N_11832,N_11927);
nor U12070 (N_12070,N_11856,N_11843);
or U12071 (N_12071,N_11766,N_11964);
nor U12072 (N_12072,N_11797,N_11763);
nor U12073 (N_12073,N_11767,N_11800);
or U12074 (N_12074,N_11979,N_11898);
and U12075 (N_12075,N_11760,N_11778);
and U12076 (N_12076,N_11853,N_11779);
and U12077 (N_12077,N_11798,N_11777);
or U12078 (N_12078,N_11938,N_11895);
nand U12079 (N_12079,N_11910,N_11781);
or U12080 (N_12080,N_11923,N_11950);
nand U12081 (N_12081,N_11790,N_11935);
nand U12082 (N_12082,N_11791,N_11916);
nor U12083 (N_12083,N_11785,N_11750);
and U12084 (N_12084,N_11806,N_11908);
nor U12085 (N_12085,N_11844,N_11951);
and U12086 (N_12086,N_11995,N_11933);
nor U12087 (N_12087,N_11757,N_11926);
nor U12088 (N_12088,N_11822,N_11900);
nand U12089 (N_12089,N_11828,N_11789);
nand U12090 (N_12090,N_11877,N_11978);
xor U12091 (N_12091,N_11771,N_11892);
nor U12092 (N_12092,N_11965,N_11932);
xor U12093 (N_12093,N_11914,N_11919);
or U12094 (N_12094,N_11834,N_11824);
or U12095 (N_12095,N_11884,N_11786);
and U12096 (N_12096,N_11770,N_11985);
and U12097 (N_12097,N_11967,N_11930);
nand U12098 (N_12098,N_11897,N_11855);
nand U12099 (N_12099,N_11980,N_11796);
nor U12100 (N_12100,N_11970,N_11782);
or U12101 (N_12101,N_11754,N_11904);
or U12102 (N_12102,N_11989,N_11956);
xor U12103 (N_12103,N_11808,N_11755);
nor U12104 (N_12104,N_11833,N_11879);
nand U12105 (N_12105,N_11819,N_11865);
nand U12106 (N_12106,N_11849,N_11852);
or U12107 (N_12107,N_11969,N_11889);
or U12108 (N_12108,N_11936,N_11881);
nor U12109 (N_12109,N_11997,N_11974);
and U12110 (N_12110,N_11887,N_11883);
nand U12111 (N_12111,N_11816,N_11862);
or U12112 (N_12112,N_11988,N_11809);
or U12113 (N_12113,N_11838,N_11994);
or U12114 (N_12114,N_11963,N_11875);
nor U12115 (N_12115,N_11864,N_11873);
and U12116 (N_12116,N_11880,N_11846);
or U12117 (N_12117,N_11802,N_11801);
or U12118 (N_12118,N_11753,N_11867);
xnor U12119 (N_12119,N_11946,N_11996);
and U12120 (N_12120,N_11891,N_11894);
nand U12121 (N_12121,N_11866,N_11917);
or U12122 (N_12122,N_11931,N_11990);
and U12123 (N_12123,N_11885,N_11998);
nand U12124 (N_12124,N_11868,N_11893);
xnor U12125 (N_12125,N_11812,N_11767);
nor U12126 (N_12126,N_11786,N_11782);
and U12127 (N_12127,N_11977,N_11897);
or U12128 (N_12128,N_11975,N_11993);
nand U12129 (N_12129,N_11830,N_11883);
nand U12130 (N_12130,N_11771,N_11850);
xnor U12131 (N_12131,N_11860,N_11858);
nand U12132 (N_12132,N_11771,N_11867);
or U12133 (N_12133,N_11983,N_11906);
nand U12134 (N_12134,N_11973,N_11998);
nand U12135 (N_12135,N_11964,N_11905);
nand U12136 (N_12136,N_11833,N_11816);
and U12137 (N_12137,N_11847,N_11804);
and U12138 (N_12138,N_11896,N_11914);
and U12139 (N_12139,N_11942,N_11891);
and U12140 (N_12140,N_11997,N_11767);
xnor U12141 (N_12141,N_11844,N_11776);
xnor U12142 (N_12142,N_11943,N_11775);
and U12143 (N_12143,N_11864,N_11971);
or U12144 (N_12144,N_11822,N_11968);
and U12145 (N_12145,N_11985,N_11987);
or U12146 (N_12146,N_11994,N_11853);
nor U12147 (N_12147,N_11799,N_11982);
nor U12148 (N_12148,N_11922,N_11976);
nor U12149 (N_12149,N_11962,N_11950);
and U12150 (N_12150,N_11759,N_11861);
nand U12151 (N_12151,N_11971,N_11813);
nand U12152 (N_12152,N_11830,N_11853);
nor U12153 (N_12153,N_11904,N_11806);
nor U12154 (N_12154,N_11864,N_11785);
xnor U12155 (N_12155,N_11900,N_11975);
or U12156 (N_12156,N_11795,N_11755);
or U12157 (N_12157,N_11848,N_11949);
nand U12158 (N_12158,N_11930,N_11806);
or U12159 (N_12159,N_11909,N_11852);
xnor U12160 (N_12160,N_11939,N_11883);
xor U12161 (N_12161,N_11991,N_11894);
nand U12162 (N_12162,N_11843,N_11996);
xnor U12163 (N_12163,N_11767,N_11904);
and U12164 (N_12164,N_11978,N_11916);
or U12165 (N_12165,N_11877,N_11972);
nor U12166 (N_12166,N_11984,N_11858);
nor U12167 (N_12167,N_11781,N_11767);
nand U12168 (N_12168,N_11801,N_11927);
xor U12169 (N_12169,N_11998,N_11917);
nor U12170 (N_12170,N_11825,N_11782);
xnor U12171 (N_12171,N_11950,N_11766);
xnor U12172 (N_12172,N_11973,N_11806);
or U12173 (N_12173,N_11841,N_11937);
xnor U12174 (N_12174,N_11985,N_11981);
nor U12175 (N_12175,N_11958,N_11804);
xor U12176 (N_12176,N_11968,N_11800);
or U12177 (N_12177,N_11891,N_11964);
xnor U12178 (N_12178,N_11794,N_11939);
xnor U12179 (N_12179,N_11773,N_11757);
nand U12180 (N_12180,N_11857,N_11862);
and U12181 (N_12181,N_11885,N_11798);
or U12182 (N_12182,N_11756,N_11862);
nor U12183 (N_12183,N_11858,N_11929);
and U12184 (N_12184,N_11934,N_11800);
or U12185 (N_12185,N_11915,N_11813);
nor U12186 (N_12186,N_11925,N_11763);
nand U12187 (N_12187,N_11931,N_11883);
or U12188 (N_12188,N_11850,N_11916);
xnor U12189 (N_12189,N_11837,N_11792);
and U12190 (N_12190,N_11830,N_11892);
xnor U12191 (N_12191,N_11922,N_11978);
and U12192 (N_12192,N_11790,N_11813);
and U12193 (N_12193,N_11888,N_11865);
nor U12194 (N_12194,N_11807,N_11793);
xor U12195 (N_12195,N_11826,N_11830);
or U12196 (N_12196,N_11981,N_11910);
nand U12197 (N_12197,N_11804,N_11914);
nor U12198 (N_12198,N_11883,N_11952);
or U12199 (N_12199,N_11874,N_11991);
nand U12200 (N_12200,N_11996,N_11776);
and U12201 (N_12201,N_11990,N_11876);
nand U12202 (N_12202,N_11794,N_11758);
nand U12203 (N_12203,N_11870,N_11872);
xor U12204 (N_12204,N_11813,N_11750);
or U12205 (N_12205,N_11822,N_11873);
nand U12206 (N_12206,N_11765,N_11849);
xor U12207 (N_12207,N_11836,N_11864);
xor U12208 (N_12208,N_11841,N_11842);
and U12209 (N_12209,N_11860,N_11842);
or U12210 (N_12210,N_11861,N_11752);
nand U12211 (N_12211,N_11877,N_11860);
or U12212 (N_12212,N_11969,N_11863);
and U12213 (N_12213,N_11790,N_11773);
nand U12214 (N_12214,N_11995,N_11977);
xor U12215 (N_12215,N_11887,N_11946);
xor U12216 (N_12216,N_11750,N_11884);
or U12217 (N_12217,N_11879,N_11889);
or U12218 (N_12218,N_11858,N_11934);
and U12219 (N_12219,N_11840,N_11807);
and U12220 (N_12220,N_11851,N_11897);
nor U12221 (N_12221,N_11762,N_11950);
and U12222 (N_12222,N_11954,N_11774);
nor U12223 (N_12223,N_11803,N_11876);
nor U12224 (N_12224,N_11789,N_11974);
nor U12225 (N_12225,N_11867,N_11986);
nand U12226 (N_12226,N_11983,N_11897);
nand U12227 (N_12227,N_11979,N_11874);
nor U12228 (N_12228,N_11817,N_11879);
xnor U12229 (N_12229,N_11942,N_11861);
nand U12230 (N_12230,N_11953,N_11822);
and U12231 (N_12231,N_11942,N_11806);
xnor U12232 (N_12232,N_11903,N_11876);
or U12233 (N_12233,N_11822,N_11898);
or U12234 (N_12234,N_11751,N_11930);
nor U12235 (N_12235,N_11944,N_11813);
xor U12236 (N_12236,N_11805,N_11819);
xor U12237 (N_12237,N_11963,N_11774);
nor U12238 (N_12238,N_11986,N_11899);
or U12239 (N_12239,N_11871,N_11880);
nor U12240 (N_12240,N_11787,N_11813);
or U12241 (N_12241,N_11805,N_11814);
or U12242 (N_12242,N_11783,N_11977);
nand U12243 (N_12243,N_11864,N_11936);
nor U12244 (N_12244,N_11983,N_11759);
xnor U12245 (N_12245,N_11883,N_11977);
and U12246 (N_12246,N_11851,N_11908);
and U12247 (N_12247,N_11756,N_11875);
nand U12248 (N_12248,N_11861,N_11823);
or U12249 (N_12249,N_11929,N_11938);
nand U12250 (N_12250,N_12002,N_12142);
or U12251 (N_12251,N_12017,N_12188);
nor U12252 (N_12252,N_12029,N_12092);
xnor U12253 (N_12253,N_12144,N_12052);
or U12254 (N_12254,N_12172,N_12143);
and U12255 (N_12255,N_12030,N_12196);
nor U12256 (N_12256,N_12060,N_12076);
or U12257 (N_12257,N_12074,N_12127);
and U12258 (N_12258,N_12079,N_12219);
or U12259 (N_12259,N_12013,N_12221);
nand U12260 (N_12260,N_12176,N_12215);
and U12261 (N_12261,N_12241,N_12012);
and U12262 (N_12262,N_12182,N_12028);
and U12263 (N_12263,N_12042,N_12171);
xnor U12264 (N_12264,N_12065,N_12032);
or U12265 (N_12265,N_12115,N_12035);
or U12266 (N_12266,N_12124,N_12061);
nor U12267 (N_12267,N_12062,N_12151);
and U12268 (N_12268,N_12208,N_12118);
or U12269 (N_12269,N_12108,N_12131);
nand U12270 (N_12270,N_12248,N_12132);
and U12271 (N_12271,N_12003,N_12077);
nand U12272 (N_12272,N_12187,N_12058);
nor U12273 (N_12273,N_12066,N_12016);
and U12274 (N_12274,N_12110,N_12243);
xnor U12275 (N_12275,N_12162,N_12008);
nor U12276 (N_12276,N_12034,N_12056);
or U12277 (N_12277,N_12129,N_12156);
and U12278 (N_12278,N_12211,N_12233);
nor U12279 (N_12279,N_12088,N_12015);
or U12280 (N_12280,N_12239,N_12206);
nor U12281 (N_12281,N_12199,N_12036);
and U12282 (N_12282,N_12152,N_12101);
or U12283 (N_12283,N_12126,N_12128);
nor U12284 (N_12284,N_12137,N_12078);
and U12285 (N_12285,N_12134,N_12240);
xor U12286 (N_12286,N_12022,N_12112);
and U12287 (N_12287,N_12155,N_12195);
or U12288 (N_12288,N_12067,N_12089);
nor U12289 (N_12289,N_12031,N_12054);
and U12290 (N_12290,N_12249,N_12020);
and U12291 (N_12291,N_12049,N_12235);
nand U12292 (N_12292,N_12202,N_12136);
and U12293 (N_12293,N_12197,N_12238);
xor U12294 (N_12294,N_12069,N_12198);
and U12295 (N_12295,N_12212,N_12138);
xor U12296 (N_12296,N_12107,N_12234);
nor U12297 (N_12297,N_12068,N_12141);
xnor U12298 (N_12298,N_12040,N_12057);
nand U12299 (N_12299,N_12210,N_12053);
xor U12300 (N_12300,N_12063,N_12217);
nor U12301 (N_12301,N_12231,N_12098);
and U12302 (N_12302,N_12072,N_12158);
nand U12303 (N_12303,N_12145,N_12184);
and U12304 (N_12304,N_12207,N_12095);
or U12305 (N_12305,N_12023,N_12175);
nor U12306 (N_12306,N_12099,N_12105);
xnor U12307 (N_12307,N_12139,N_12026);
and U12308 (N_12308,N_12045,N_12192);
xnor U12309 (N_12309,N_12037,N_12019);
xnor U12310 (N_12310,N_12181,N_12185);
xnor U12311 (N_12311,N_12117,N_12071);
xor U12312 (N_12312,N_12021,N_12203);
or U12313 (N_12313,N_12097,N_12087);
nor U12314 (N_12314,N_12227,N_12170);
or U12315 (N_12315,N_12167,N_12194);
nor U12316 (N_12316,N_12153,N_12247);
xnor U12317 (N_12317,N_12174,N_12006);
or U12318 (N_12318,N_12051,N_12193);
nor U12319 (N_12319,N_12205,N_12004);
or U12320 (N_12320,N_12044,N_12083);
xnor U12321 (N_12321,N_12223,N_12119);
nand U12322 (N_12322,N_12218,N_12059);
xnor U12323 (N_12323,N_12055,N_12220);
nand U12324 (N_12324,N_12080,N_12146);
or U12325 (N_12325,N_12135,N_12047);
nand U12326 (N_12326,N_12244,N_12041);
and U12327 (N_12327,N_12070,N_12140);
xor U12328 (N_12328,N_12073,N_12122);
xnor U12329 (N_12329,N_12213,N_12164);
nand U12330 (N_12330,N_12106,N_12024);
nor U12331 (N_12331,N_12100,N_12237);
nand U12332 (N_12332,N_12005,N_12165);
nor U12333 (N_12333,N_12200,N_12186);
or U12334 (N_12334,N_12091,N_12224);
or U12335 (N_12335,N_12190,N_12130);
xor U12336 (N_12336,N_12064,N_12096);
and U12337 (N_12337,N_12232,N_12007);
nor U12338 (N_12338,N_12093,N_12075);
and U12339 (N_12339,N_12111,N_12226);
xor U12340 (N_12340,N_12084,N_12046);
nand U12341 (N_12341,N_12082,N_12001);
nor U12342 (N_12342,N_12000,N_12180);
nor U12343 (N_12343,N_12114,N_12094);
nand U12344 (N_12344,N_12014,N_12113);
nor U12345 (N_12345,N_12033,N_12245);
and U12346 (N_12346,N_12120,N_12038);
xnor U12347 (N_12347,N_12173,N_12011);
xnor U12348 (N_12348,N_12009,N_12225);
and U12349 (N_12349,N_12242,N_12025);
or U12350 (N_12350,N_12216,N_12201);
xor U12351 (N_12351,N_12222,N_12043);
nor U12352 (N_12352,N_12086,N_12191);
or U12353 (N_12353,N_12168,N_12050);
or U12354 (N_12354,N_12189,N_12179);
and U12355 (N_12355,N_12090,N_12147);
and U12356 (N_12356,N_12163,N_12183);
nor U12357 (N_12357,N_12125,N_12228);
or U12358 (N_12358,N_12148,N_12150);
or U12359 (N_12359,N_12177,N_12102);
xor U12360 (N_12360,N_12209,N_12039);
and U12361 (N_12361,N_12154,N_12116);
xor U12362 (N_12362,N_12103,N_12048);
nor U12363 (N_12363,N_12229,N_12149);
and U12364 (N_12364,N_12157,N_12159);
or U12365 (N_12365,N_12178,N_12204);
xnor U12366 (N_12366,N_12081,N_12085);
xnor U12367 (N_12367,N_12230,N_12018);
and U12368 (N_12368,N_12160,N_12161);
xnor U12369 (N_12369,N_12166,N_12121);
and U12370 (N_12370,N_12104,N_12109);
nor U12371 (N_12371,N_12236,N_12027);
or U12372 (N_12372,N_12214,N_12246);
or U12373 (N_12373,N_12123,N_12169);
or U12374 (N_12374,N_12133,N_12010);
xor U12375 (N_12375,N_12239,N_12245);
or U12376 (N_12376,N_12130,N_12071);
nand U12377 (N_12377,N_12056,N_12148);
nor U12378 (N_12378,N_12055,N_12085);
nand U12379 (N_12379,N_12245,N_12080);
nand U12380 (N_12380,N_12057,N_12011);
xnor U12381 (N_12381,N_12195,N_12132);
or U12382 (N_12382,N_12243,N_12165);
and U12383 (N_12383,N_12065,N_12135);
nand U12384 (N_12384,N_12046,N_12039);
and U12385 (N_12385,N_12168,N_12026);
nor U12386 (N_12386,N_12217,N_12080);
or U12387 (N_12387,N_12185,N_12096);
nand U12388 (N_12388,N_12080,N_12158);
nor U12389 (N_12389,N_12131,N_12109);
or U12390 (N_12390,N_12117,N_12171);
or U12391 (N_12391,N_12054,N_12191);
and U12392 (N_12392,N_12091,N_12073);
nor U12393 (N_12393,N_12225,N_12216);
nand U12394 (N_12394,N_12226,N_12156);
and U12395 (N_12395,N_12193,N_12112);
nor U12396 (N_12396,N_12192,N_12237);
nor U12397 (N_12397,N_12005,N_12144);
and U12398 (N_12398,N_12000,N_12034);
and U12399 (N_12399,N_12003,N_12117);
nor U12400 (N_12400,N_12173,N_12007);
xnor U12401 (N_12401,N_12061,N_12188);
xnor U12402 (N_12402,N_12128,N_12041);
nand U12403 (N_12403,N_12020,N_12023);
and U12404 (N_12404,N_12184,N_12157);
or U12405 (N_12405,N_12038,N_12116);
or U12406 (N_12406,N_12139,N_12130);
and U12407 (N_12407,N_12246,N_12184);
and U12408 (N_12408,N_12136,N_12114);
nor U12409 (N_12409,N_12109,N_12051);
or U12410 (N_12410,N_12012,N_12158);
nor U12411 (N_12411,N_12126,N_12007);
nor U12412 (N_12412,N_12072,N_12172);
or U12413 (N_12413,N_12171,N_12180);
nor U12414 (N_12414,N_12094,N_12245);
xnor U12415 (N_12415,N_12065,N_12205);
nor U12416 (N_12416,N_12114,N_12089);
xnor U12417 (N_12417,N_12070,N_12231);
and U12418 (N_12418,N_12115,N_12142);
and U12419 (N_12419,N_12054,N_12134);
or U12420 (N_12420,N_12141,N_12123);
xor U12421 (N_12421,N_12054,N_12222);
or U12422 (N_12422,N_12195,N_12084);
and U12423 (N_12423,N_12079,N_12166);
nand U12424 (N_12424,N_12202,N_12077);
nand U12425 (N_12425,N_12187,N_12172);
or U12426 (N_12426,N_12021,N_12071);
xnor U12427 (N_12427,N_12056,N_12215);
nor U12428 (N_12428,N_12111,N_12081);
nor U12429 (N_12429,N_12027,N_12089);
nand U12430 (N_12430,N_12221,N_12237);
or U12431 (N_12431,N_12197,N_12156);
nand U12432 (N_12432,N_12131,N_12171);
nand U12433 (N_12433,N_12043,N_12246);
or U12434 (N_12434,N_12123,N_12209);
and U12435 (N_12435,N_12042,N_12109);
and U12436 (N_12436,N_12042,N_12046);
xor U12437 (N_12437,N_12120,N_12060);
and U12438 (N_12438,N_12224,N_12012);
and U12439 (N_12439,N_12181,N_12246);
or U12440 (N_12440,N_12101,N_12249);
nand U12441 (N_12441,N_12108,N_12162);
xnor U12442 (N_12442,N_12214,N_12221);
nand U12443 (N_12443,N_12043,N_12119);
nor U12444 (N_12444,N_12023,N_12097);
and U12445 (N_12445,N_12137,N_12084);
and U12446 (N_12446,N_12181,N_12123);
nand U12447 (N_12447,N_12088,N_12171);
or U12448 (N_12448,N_12121,N_12191);
and U12449 (N_12449,N_12097,N_12018);
or U12450 (N_12450,N_12181,N_12183);
xnor U12451 (N_12451,N_12056,N_12117);
nor U12452 (N_12452,N_12171,N_12090);
nand U12453 (N_12453,N_12025,N_12184);
xor U12454 (N_12454,N_12072,N_12230);
and U12455 (N_12455,N_12141,N_12131);
or U12456 (N_12456,N_12081,N_12184);
and U12457 (N_12457,N_12191,N_12219);
or U12458 (N_12458,N_12054,N_12060);
nor U12459 (N_12459,N_12087,N_12072);
xor U12460 (N_12460,N_12091,N_12020);
or U12461 (N_12461,N_12086,N_12231);
nor U12462 (N_12462,N_12200,N_12235);
and U12463 (N_12463,N_12133,N_12101);
nand U12464 (N_12464,N_12120,N_12244);
xor U12465 (N_12465,N_12152,N_12171);
or U12466 (N_12466,N_12144,N_12034);
nand U12467 (N_12467,N_12045,N_12196);
nand U12468 (N_12468,N_12046,N_12069);
xor U12469 (N_12469,N_12161,N_12071);
nand U12470 (N_12470,N_12020,N_12008);
and U12471 (N_12471,N_12074,N_12154);
nand U12472 (N_12472,N_12202,N_12219);
and U12473 (N_12473,N_12167,N_12056);
xor U12474 (N_12474,N_12066,N_12142);
xnor U12475 (N_12475,N_12035,N_12015);
nor U12476 (N_12476,N_12125,N_12008);
xor U12477 (N_12477,N_12019,N_12069);
xor U12478 (N_12478,N_12041,N_12187);
nand U12479 (N_12479,N_12164,N_12041);
or U12480 (N_12480,N_12237,N_12186);
and U12481 (N_12481,N_12117,N_12023);
nor U12482 (N_12482,N_12131,N_12128);
xnor U12483 (N_12483,N_12116,N_12212);
or U12484 (N_12484,N_12153,N_12135);
nor U12485 (N_12485,N_12008,N_12113);
xor U12486 (N_12486,N_12185,N_12213);
nor U12487 (N_12487,N_12220,N_12184);
nor U12488 (N_12488,N_12234,N_12018);
nor U12489 (N_12489,N_12203,N_12222);
nand U12490 (N_12490,N_12062,N_12175);
xor U12491 (N_12491,N_12099,N_12185);
nand U12492 (N_12492,N_12137,N_12182);
or U12493 (N_12493,N_12075,N_12101);
nor U12494 (N_12494,N_12040,N_12008);
or U12495 (N_12495,N_12085,N_12203);
xnor U12496 (N_12496,N_12104,N_12175);
nor U12497 (N_12497,N_12090,N_12056);
xor U12498 (N_12498,N_12057,N_12068);
nor U12499 (N_12499,N_12108,N_12153);
nand U12500 (N_12500,N_12307,N_12352);
and U12501 (N_12501,N_12395,N_12469);
and U12502 (N_12502,N_12455,N_12423);
and U12503 (N_12503,N_12499,N_12279);
nor U12504 (N_12504,N_12303,N_12453);
nand U12505 (N_12505,N_12321,N_12315);
nand U12506 (N_12506,N_12374,N_12465);
or U12507 (N_12507,N_12470,N_12413);
nand U12508 (N_12508,N_12342,N_12323);
nor U12509 (N_12509,N_12471,N_12353);
nand U12510 (N_12510,N_12280,N_12488);
nor U12511 (N_12511,N_12306,N_12466);
or U12512 (N_12512,N_12474,N_12350);
and U12513 (N_12513,N_12344,N_12447);
and U12514 (N_12514,N_12430,N_12347);
and U12515 (N_12515,N_12480,N_12327);
nand U12516 (N_12516,N_12359,N_12394);
and U12517 (N_12517,N_12376,N_12490);
nor U12518 (N_12518,N_12408,N_12265);
nand U12519 (N_12519,N_12497,N_12366);
xnor U12520 (N_12520,N_12457,N_12355);
nand U12521 (N_12521,N_12271,N_12485);
or U12522 (N_12522,N_12328,N_12392);
nor U12523 (N_12523,N_12496,N_12459);
xor U12524 (N_12524,N_12282,N_12334);
nand U12525 (N_12525,N_12288,N_12351);
nor U12526 (N_12526,N_12338,N_12448);
or U12527 (N_12527,N_12293,N_12358);
and U12528 (N_12528,N_12391,N_12377);
xor U12529 (N_12529,N_12285,N_12283);
xnor U12530 (N_12530,N_12380,N_12363);
nand U12531 (N_12531,N_12425,N_12481);
xor U12532 (N_12532,N_12415,N_12393);
nand U12533 (N_12533,N_12274,N_12446);
xnor U12534 (N_12534,N_12254,N_12368);
or U12535 (N_12535,N_12317,N_12487);
nand U12536 (N_12536,N_12440,N_12267);
nor U12537 (N_12537,N_12349,N_12291);
or U12538 (N_12538,N_12320,N_12275);
and U12539 (N_12539,N_12258,N_12403);
nand U12540 (N_12540,N_12322,N_12407);
xor U12541 (N_12541,N_12437,N_12435);
nor U12542 (N_12542,N_12445,N_12257);
nor U12543 (N_12543,N_12493,N_12489);
nor U12544 (N_12544,N_12364,N_12292);
and U12545 (N_12545,N_12467,N_12477);
nand U12546 (N_12546,N_12450,N_12373);
and U12547 (N_12547,N_12332,N_12313);
nand U12548 (N_12548,N_12397,N_12308);
nand U12549 (N_12549,N_12337,N_12464);
xor U12550 (N_12550,N_12482,N_12396);
nor U12551 (N_12551,N_12297,N_12284);
xnor U12552 (N_12552,N_12406,N_12433);
nor U12553 (N_12553,N_12411,N_12498);
and U12554 (N_12554,N_12398,N_12438);
or U12555 (N_12555,N_12314,N_12375);
nand U12556 (N_12556,N_12382,N_12354);
xnor U12557 (N_12557,N_12256,N_12277);
nand U12558 (N_12558,N_12473,N_12309);
nor U12559 (N_12559,N_12422,N_12386);
and U12560 (N_12560,N_12268,N_12319);
nor U12561 (N_12561,N_12259,N_12476);
and U12562 (N_12562,N_12443,N_12451);
or U12563 (N_12563,N_12272,N_12478);
xnor U12564 (N_12564,N_12266,N_12287);
or U12565 (N_12565,N_12281,N_12399);
xnor U12566 (N_12566,N_12318,N_12343);
xnor U12567 (N_12567,N_12360,N_12458);
nand U12568 (N_12568,N_12330,N_12372);
nor U12569 (N_12569,N_12356,N_12341);
and U12570 (N_12570,N_12405,N_12316);
or U12571 (N_12571,N_12427,N_12310);
nor U12572 (N_12572,N_12460,N_12252);
and U12573 (N_12573,N_12494,N_12357);
or U12574 (N_12574,N_12424,N_12312);
or U12575 (N_12575,N_12270,N_12461);
nor U12576 (N_12576,N_12388,N_12333);
or U12577 (N_12577,N_12441,N_12304);
or U12578 (N_12578,N_12421,N_12420);
or U12579 (N_12579,N_12409,N_12444);
nor U12580 (N_12580,N_12432,N_12326);
xor U12581 (N_12581,N_12381,N_12339);
xnor U12582 (N_12582,N_12429,N_12475);
or U12583 (N_12583,N_12289,N_12324);
xnor U12584 (N_12584,N_12462,N_12251);
nand U12585 (N_12585,N_12404,N_12491);
xnor U12586 (N_12586,N_12449,N_12463);
xnor U12587 (N_12587,N_12390,N_12296);
nor U12588 (N_12588,N_12298,N_12325);
nand U12589 (N_12589,N_12483,N_12486);
and U12590 (N_12590,N_12294,N_12336);
nor U12591 (N_12591,N_12348,N_12479);
and U12592 (N_12592,N_12442,N_12419);
nor U12593 (N_12593,N_12346,N_12495);
and U12594 (N_12594,N_12454,N_12367);
nand U12595 (N_12595,N_12278,N_12264);
nor U12596 (N_12596,N_12362,N_12389);
nor U12597 (N_12597,N_12414,N_12369);
and U12598 (N_12598,N_12387,N_12295);
or U12599 (N_12599,N_12261,N_12379);
nand U12600 (N_12600,N_12378,N_12302);
nor U12601 (N_12601,N_12468,N_12345);
or U12602 (N_12602,N_12371,N_12255);
and U12603 (N_12603,N_12436,N_12384);
nand U12604 (N_12604,N_12431,N_12401);
nand U12605 (N_12605,N_12370,N_12434);
or U12606 (N_12606,N_12340,N_12311);
and U12607 (N_12607,N_12361,N_12383);
nor U12608 (N_12608,N_12402,N_12335);
nand U12609 (N_12609,N_12492,N_12452);
and U12610 (N_12610,N_12276,N_12286);
nor U12611 (N_12611,N_12273,N_12417);
or U12612 (N_12612,N_12439,N_12428);
nor U12613 (N_12613,N_12300,N_12263);
nand U12614 (N_12614,N_12262,N_12426);
nor U12615 (N_12615,N_12416,N_12299);
or U12616 (N_12616,N_12250,N_12290);
nand U12617 (N_12617,N_12305,N_12365);
nor U12618 (N_12618,N_12301,N_12329);
and U12619 (N_12619,N_12412,N_12410);
and U12620 (N_12620,N_12331,N_12253);
xnor U12621 (N_12621,N_12456,N_12400);
nor U12622 (N_12622,N_12472,N_12418);
xor U12623 (N_12623,N_12269,N_12385);
and U12624 (N_12624,N_12484,N_12260);
or U12625 (N_12625,N_12432,N_12485);
nor U12626 (N_12626,N_12341,N_12420);
and U12627 (N_12627,N_12358,N_12479);
and U12628 (N_12628,N_12463,N_12296);
xnor U12629 (N_12629,N_12476,N_12325);
nand U12630 (N_12630,N_12481,N_12470);
xor U12631 (N_12631,N_12360,N_12391);
and U12632 (N_12632,N_12342,N_12367);
nor U12633 (N_12633,N_12260,N_12263);
and U12634 (N_12634,N_12458,N_12480);
or U12635 (N_12635,N_12357,N_12305);
nor U12636 (N_12636,N_12370,N_12281);
nor U12637 (N_12637,N_12337,N_12449);
nand U12638 (N_12638,N_12276,N_12466);
and U12639 (N_12639,N_12390,N_12437);
or U12640 (N_12640,N_12415,N_12440);
and U12641 (N_12641,N_12460,N_12471);
xnor U12642 (N_12642,N_12310,N_12357);
and U12643 (N_12643,N_12425,N_12381);
nor U12644 (N_12644,N_12328,N_12409);
and U12645 (N_12645,N_12287,N_12375);
nand U12646 (N_12646,N_12370,N_12298);
and U12647 (N_12647,N_12266,N_12382);
and U12648 (N_12648,N_12433,N_12415);
nor U12649 (N_12649,N_12486,N_12308);
xnor U12650 (N_12650,N_12427,N_12268);
nand U12651 (N_12651,N_12370,N_12354);
or U12652 (N_12652,N_12349,N_12477);
nor U12653 (N_12653,N_12252,N_12278);
xor U12654 (N_12654,N_12257,N_12385);
xnor U12655 (N_12655,N_12372,N_12480);
nor U12656 (N_12656,N_12391,N_12271);
nand U12657 (N_12657,N_12326,N_12273);
xnor U12658 (N_12658,N_12494,N_12342);
nor U12659 (N_12659,N_12414,N_12268);
or U12660 (N_12660,N_12422,N_12497);
nand U12661 (N_12661,N_12268,N_12410);
or U12662 (N_12662,N_12411,N_12381);
nand U12663 (N_12663,N_12398,N_12380);
and U12664 (N_12664,N_12480,N_12452);
xor U12665 (N_12665,N_12340,N_12291);
or U12666 (N_12666,N_12471,N_12451);
xnor U12667 (N_12667,N_12299,N_12336);
and U12668 (N_12668,N_12428,N_12322);
nor U12669 (N_12669,N_12469,N_12288);
nor U12670 (N_12670,N_12298,N_12374);
or U12671 (N_12671,N_12479,N_12251);
and U12672 (N_12672,N_12303,N_12354);
nand U12673 (N_12673,N_12307,N_12383);
and U12674 (N_12674,N_12366,N_12354);
xor U12675 (N_12675,N_12296,N_12308);
nor U12676 (N_12676,N_12487,N_12371);
nor U12677 (N_12677,N_12333,N_12394);
and U12678 (N_12678,N_12320,N_12330);
nand U12679 (N_12679,N_12435,N_12333);
nand U12680 (N_12680,N_12417,N_12441);
xor U12681 (N_12681,N_12348,N_12320);
xor U12682 (N_12682,N_12487,N_12289);
nand U12683 (N_12683,N_12275,N_12330);
and U12684 (N_12684,N_12341,N_12454);
nand U12685 (N_12685,N_12282,N_12429);
xor U12686 (N_12686,N_12445,N_12448);
and U12687 (N_12687,N_12455,N_12496);
xnor U12688 (N_12688,N_12423,N_12308);
or U12689 (N_12689,N_12257,N_12481);
xor U12690 (N_12690,N_12375,N_12264);
nand U12691 (N_12691,N_12319,N_12432);
nand U12692 (N_12692,N_12448,N_12412);
nand U12693 (N_12693,N_12393,N_12276);
or U12694 (N_12694,N_12314,N_12383);
or U12695 (N_12695,N_12407,N_12257);
and U12696 (N_12696,N_12387,N_12486);
nand U12697 (N_12697,N_12435,N_12298);
nand U12698 (N_12698,N_12373,N_12405);
xor U12699 (N_12699,N_12480,N_12323);
and U12700 (N_12700,N_12322,N_12492);
nand U12701 (N_12701,N_12441,N_12380);
or U12702 (N_12702,N_12348,N_12475);
xor U12703 (N_12703,N_12330,N_12321);
and U12704 (N_12704,N_12386,N_12424);
nor U12705 (N_12705,N_12351,N_12359);
or U12706 (N_12706,N_12353,N_12372);
and U12707 (N_12707,N_12412,N_12299);
or U12708 (N_12708,N_12348,N_12369);
or U12709 (N_12709,N_12254,N_12458);
xnor U12710 (N_12710,N_12368,N_12303);
or U12711 (N_12711,N_12428,N_12459);
or U12712 (N_12712,N_12279,N_12385);
xnor U12713 (N_12713,N_12494,N_12465);
nand U12714 (N_12714,N_12374,N_12437);
xor U12715 (N_12715,N_12288,N_12278);
nor U12716 (N_12716,N_12474,N_12322);
and U12717 (N_12717,N_12310,N_12489);
or U12718 (N_12718,N_12348,N_12439);
nor U12719 (N_12719,N_12493,N_12359);
nand U12720 (N_12720,N_12274,N_12457);
nor U12721 (N_12721,N_12434,N_12460);
nand U12722 (N_12722,N_12440,N_12424);
and U12723 (N_12723,N_12473,N_12360);
and U12724 (N_12724,N_12302,N_12359);
nor U12725 (N_12725,N_12252,N_12381);
or U12726 (N_12726,N_12437,N_12382);
nand U12727 (N_12727,N_12310,N_12494);
xnor U12728 (N_12728,N_12351,N_12406);
nand U12729 (N_12729,N_12491,N_12406);
or U12730 (N_12730,N_12261,N_12325);
nor U12731 (N_12731,N_12424,N_12439);
or U12732 (N_12732,N_12302,N_12292);
or U12733 (N_12733,N_12275,N_12496);
or U12734 (N_12734,N_12262,N_12413);
nand U12735 (N_12735,N_12463,N_12309);
or U12736 (N_12736,N_12295,N_12472);
xor U12737 (N_12737,N_12468,N_12383);
nor U12738 (N_12738,N_12253,N_12338);
xor U12739 (N_12739,N_12392,N_12439);
xnor U12740 (N_12740,N_12333,N_12325);
nand U12741 (N_12741,N_12327,N_12253);
or U12742 (N_12742,N_12291,N_12450);
xor U12743 (N_12743,N_12305,N_12353);
or U12744 (N_12744,N_12295,N_12452);
xor U12745 (N_12745,N_12413,N_12265);
xor U12746 (N_12746,N_12471,N_12464);
or U12747 (N_12747,N_12477,N_12388);
xor U12748 (N_12748,N_12253,N_12325);
xor U12749 (N_12749,N_12342,N_12444);
nand U12750 (N_12750,N_12600,N_12673);
nand U12751 (N_12751,N_12610,N_12729);
nand U12752 (N_12752,N_12583,N_12700);
and U12753 (N_12753,N_12508,N_12694);
nor U12754 (N_12754,N_12615,N_12545);
xnor U12755 (N_12755,N_12530,N_12690);
and U12756 (N_12756,N_12618,N_12547);
nand U12757 (N_12757,N_12704,N_12743);
nand U12758 (N_12758,N_12635,N_12601);
nand U12759 (N_12759,N_12726,N_12539);
nor U12760 (N_12760,N_12506,N_12513);
and U12761 (N_12761,N_12682,N_12685);
nand U12762 (N_12762,N_12703,N_12578);
nor U12763 (N_12763,N_12579,N_12723);
and U12764 (N_12764,N_12549,N_12533);
nor U12765 (N_12765,N_12681,N_12526);
xor U12766 (N_12766,N_12660,N_12701);
and U12767 (N_12767,N_12702,N_12632);
and U12768 (N_12768,N_12639,N_12689);
and U12769 (N_12769,N_12577,N_12551);
nand U12770 (N_12770,N_12634,N_12564);
xnor U12771 (N_12771,N_12705,N_12696);
xor U12772 (N_12772,N_12646,N_12567);
or U12773 (N_12773,N_12621,N_12569);
nand U12774 (N_12774,N_12736,N_12648);
or U12775 (N_12775,N_12565,N_12645);
nor U12776 (N_12776,N_12688,N_12663);
nand U12777 (N_12777,N_12586,N_12584);
or U12778 (N_12778,N_12517,N_12536);
or U12779 (N_12779,N_12607,N_12713);
nand U12780 (N_12780,N_12747,N_12570);
nor U12781 (N_12781,N_12587,N_12502);
nor U12782 (N_12782,N_12557,N_12515);
or U12783 (N_12783,N_12711,N_12715);
nor U12784 (N_12784,N_12738,N_12541);
xnor U12785 (N_12785,N_12653,N_12603);
nand U12786 (N_12786,N_12636,N_12650);
or U12787 (N_12787,N_12678,N_12592);
or U12788 (N_12788,N_12616,N_12611);
nand U12789 (N_12789,N_12649,N_12679);
xor U12790 (N_12790,N_12739,N_12529);
and U12791 (N_12791,N_12745,N_12698);
nor U12792 (N_12792,N_12631,N_12588);
and U12793 (N_12793,N_12582,N_12626);
nand U12794 (N_12794,N_12655,N_12590);
or U12795 (N_12795,N_12683,N_12581);
and U12796 (N_12796,N_12677,N_12624);
or U12797 (N_12797,N_12562,N_12593);
nor U12798 (N_12798,N_12730,N_12642);
or U12799 (N_12799,N_12604,N_12518);
and U12800 (N_12800,N_12623,N_12671);
xor U12801 (N_12801,N_12609,N_12612);
nand U12802 (N_12802,N_12658,N_12544);
xnor U12803 (N_12803,N_12641,N_12516);
nand U12804 (N_12804,N_12652,N_12534);
nor U12805 (N_12805,N_12602,N_12669);
nor U12806 (N_12806,N_12680,N_12695);
and U12807 (N_12807,N_12532,N_12691);
or U12808 (N_12808,N_12501,N_12563);
nand U12809 (N_12809,N_12596,N_12554);
nor U12810 (N_12810,N_12598,N_12628);
nor U12811 (N_12811,N_12523,N_12656);
nor U12812 (N_12812,N_12651,N_12748);
nand U12813 (N_12813,N_12620,N_12708);
and U12814 (N_12814,N_12540,N_12555);
and U12815 (N_12815,N_12566,N_12637);
nand U12816 (N_12816,N_12521,N_12640);
xor U12817 (N_12817,N_12672,N_12505);
and U12818 (N_12818,N_12737,N_12718);
or U12819 (N_12819,N_12556,N_12599);
nand U12820 (N_12820,N_12619,N_12527);
xor U12821 (N_12821,N_12659,N_12668);
and U12822 (N_12822,N_12714,N_12693);
or U12823 (N_12823,N_12722,N_12749);
xnor U12824 (N_12824,N_12727,N_12538);
or U12825 (N_12825,N_12724,N_12699);
nand U12826 (N_12826,N_12525,N_12697);
xor U12827 (N_12827,N_12720,N_12742);
nor U12828 (N_12828,N_12537,N_12524);
nand U12829 (N_12829,N_12509,N_12574);
or U12830 (N_12830,N_12512,N_12644);
nor U12831 (N_12831,N_12731,N_12511);
nor U12832 (N_12832,N_12528,N_12719);
xor U12833 (N_12833,N_12732,N_12675);
xor U12834 (N_12834,N_12520,N_12709);
nand U12835 (N_12835,N_12560,N_12510);
nand U12836 (N_12836,N_12674,N_12746);
or U12837 (N_12837,N_12622,N_12734);
or U12838 (N_12838,N_12507,N_12667);
nor U12839 (N_12839,N_12580,N_12591);
or U12840 (N_12840,N_12670,N_12744);
nor U12841 (N_12841,N_12617,N_12546);
and U12842 (N_12842,N_12614,N_12661);
nand U12843 (N_12843,N_12608,N_12741);
xor U12844 (N_12844,N_12687,N_12630);
or U12845 (N_12845,N_12647,N_12543);
nand U12846 (N_12846,N_12504,N_12500);
xor U12847 (N_12847,N_12735,N_12606);
and U12848 (N_12848,N_12633,N_12519);
xor U12849 (N_12849,N_12712,N_12638);
and U12850 (N_12850,N_12522,N_12721);
nor U12851 (N_12851,N_12589,N_12740);
and U12852 (N_12852,N_12725,N_12676);
and U12853 (N_12853,N_12552,N_12550);
nor U12854 (N_12854,N_12733,N_12728);
or U12855 (N_12855,N_12605,N_12657);
and U12856 (N_12856,N_12627,N_12559);
and U12857 (N_12857,N_12576,N_12706);
and U12858 (N_12858,N_12594,N_12561);
and U12859 (N_12859,N_12531,N_12572);
and U12860 (N_12860,N_12625,N_12666);
nor U12861 (N_12861,N_12548,N_12707);
nor U12862 (N_12862,N_12710,N_12568);
nand U12863 (N_12863,N_12542,N_12665);
nor U12864 (N_12864,N_12503,N_12571);
nand U12865 (N_12865,N_12654,N_12717);
nand U12866 (N_12866,N_12684,N_12573);
or U12867 (N_12867,N_12662,N_12613);
and U12868 (N_12868,N_12585,N_12535);
nor U12869 (N_12869,N_12514,N_12597);
and U12870 (N_12870,N_12558,N_12643);
nor U12871 (N_12871,N_12629,N_12595);
and U12872 (N_12872,N_12716,N_12664);
nand U12873 (N_12873,N_12575,N_12692);
or U12874 (N_12874,N_12553,N_12686);
nand U12875 (N_12875,N_12531,N_12568);
nand U12876 (N_12876,N_12520,N_12675);
or U12877 (N_12877,N_12720,N_12707);
nand U12878 (N_12878,N_12652,N_12699);
xor U12879 (N_12879,N_12528,N_12732);
or U12880 (N_12880,N_12694,N_12551);
nor U12881 (N_12881,N_12657,N_12540);
nand U12882 (N_12882,N_12627,N_12616);
nand U12883 (N_12883,N_12508,N_12505);
nand U12884 (N_12884,N_12726,N_12549);
nor U12885 (N_12885,N_12519,N_12527);
nor U12886 (N_12886,N_12745,N_12670);
and U12887 (N_12887,N_12597,N_12730);
nor U12888 (N_12888,N_12744,N_12535);
or U12889 (N_12889,N_12738,N_12510);
or U12890 (N_12890,N_12581,N_12663);
and U12891 (N_12891,N_12514,N_12561);
xor U12892 (N_12892,N_12538,N_12677);
nand U12893 (N_12893,N_12731,N_12734);
and U12894 (N_12894,N_12723,N_12725);
and U12895 (N_12895,N_12581,N_12719);
nor U12896 (N_12896,N_12569,N_12644);
nor U12897 (N_12897,N_12732,N_12604);
xor U12898 (N_12898,N_12532,N_12634);
or U12899 (N_12899,N_12721,N_12570);
xor U12900 (N_12900,N_12730,N_12671);
or U12901 (N_12901,N_12706,N_12546);
and U12902 (N_12902,N_12673,N_12692);
nor U12903 (N_12903,N_12727,N_12694);
or U12904 (N_12904,N_12673,N_12682);
nand U12905 (N_12905,N_12692,N_12655);
nor U12906 (N_12906,N_12673,N_12571);
nand U12907 (N_12907,N_12507,N_12631);
and U12908 (N_12908,N_12714,N_12501);
or U12909 (N_12909,N_12559,N_12587);
xor U12910 (N_12910,N_12720,N_12679);
nand U12911 (N_12911,N_12542,N_12518);
and U12912 (N_12912,N_12639,N_12693);
or U12913 (N_12913,N_12646,N_12530);
nor U12914 (N_12914,N_12678,N_12632);
or U12915 (N_12915,N_12582,N_12745);
nor U12916 (N_12916,N_12670,N_12566);
nor U12917 (N_12917,N_12749,N_12598);
nor U12918 (N_12918,N_12527,N_12679);
nand U12919 (N_12919,N_12568,N_12540);
or U12920 (N_12920,N_12684,N_12610);
nor U12921 (N_12921,N_12506,N_12674);
nor U12922 (N_12922,N_12646,N_12664);
and U12923 (N_12923,N_12675,N_12635);
or U12924 (N_12924,N_12749,N_12638);
nor U12925 (N_12925,N_12694,N_12696);
nand U12926 (N_12926,N_12589,N_12748);
xnor U12927 (N_12927,N_12509,N_12610);
nand U12928 (N_12928,N_12506,N_12587);
and U12929 (N_12929,N_12613,N_12740);
nand U12930 (N_12930,N_12716,N_12549);
xor U12931 (N_12931,N_12721,N_12661);
nor U12932 (N_12932,N_12737,N_12602);
and U12933 (N_12933,N_12507,N_12677);
xor U12934 (N_12934,N_12642,N_12527);
xnor U12935 (N_12935,N_12594,N_12644);
xor U12936 (N_12936,N_12554,N_12540);
or U12937 (N_12937,N_12738,N_12724);
nand U12938 (N_12938,N_12540,N_12698);
or U12939 (N_12939,N_12747,N_12660);
nor U12940 (N_12940,N_12544,N_12543);
nand U12941 (N_12941,N_12648,N_12705);
xnor U12942 (N_12942,N_12589,N_12540);
nand U12943 (N_12943,N_12684,N_12538);
xnor U12944 (N_12944,N_12718,N_12623);
or U12945 (N_12945,N_12520,N_12598);
xnor U12946 (N_12946,N_12699,N_12679);
or U12947 (N_12947,N_12630,N_12721);
xor U12948 (N_12948,N_12705,N_12651);
and U12949 (N_12949,N_12617,N_12680);
nand U12950 (N_12950,N_12661,N_12745);
xnor U12951 (N_12951,N_12670,N_12594);
or U12952 (N_12952,N_12749,N_12569);
xnor U12953 (N_12953,N_12627,N_12509);
xnor U12954 (N_12954,N_12662,N_12529);
and U12955 (N_12955,N_12728,N_12637);
nand U12956 (N_12956,N_12653,N_12645);
xnor U12957 (N_12957,N_12719,N_12715);
and U12958 (N_12958,N_12738,N_12665);
and U12959 (N_12959,N_12716,N_12517);
xor U12960 (N_12960,N_12515,N_12585);
xor U12961 (N_12961,N_12669,N_12739);
nor U12962 (N_12962,N_12693,N_12504);
and U12963 (N_12963,N_12681,N_12541);
xnor U12964 (N_12964,N_12546,N_12569);
or U12965 (N_12965,N_12641,N_12518);
nand U12966 (N_12966,N_12516,N_12656);
or U12967 (N_12967,N_12712,N_12565);
or U12968 (N_12968,N_12565,N_12638);
nand U12969 (N_12969,N_12558,N_12736);
or U12970 (N_12970,N_12637,N_12575);
nand U12971 (N_12971,N_12592,N_12655);
and U12972 (N_12972,N_12561,N_12740);
nor U12973 (N_12973,N_12743,N_12698);
or U12974 (N_12974,N_12508,N_12744);
nand U12975 (N_12975,N_12598,N_12514);
xnor U12976 (N_12976,N_12689,N_12610);
nor U12977 (N_12977,N_12565,N_12744);
nor U12978 (N_12978,N_12645,N_12678);
xnor U12979 (N_12979,N_12508,N_12540);
or U12980 (N_12980,N_12703,N_12572);
and U12981 (N_12981,N_12616,N_12592);
xnor U12982 (N_12982,N_12725,N_12600);
and U12983 (N_12983,N_12589,N_12591);
or U12984 (N_12984,N_12622,N_12525);
nand U12985 (N_12985,N_12570,N_12712);
nor U12986 (N_12986,N_12601,N_12557);
nand U12987 (N_12987,N_12694,N_12628);
or U12988 (N_12988,N_12609,N_12567);
nor U12989 (N_12989,N_12744,N_12593);
or U12990 (N_12990,N_12524,N_12698);
xor U12991 (N_12991,N_12501,N_12731);
nor U12992 (N_12992,N_12687,N_12736);
nor U12993 (N_12993,N_12695,N_12531);
xnor U12994 (N_12994,N_12670,N_12501);
nand U12995 (N_12995,N_12642,N_12709);
and U12996 (N_12996,N_12553,N_12744);
and U12997 (N_12997,N_12577,N_12664);
and U12998 (N_12998,N_12525,N_12500);
and U12999 (N_12999,N_12600,N_12685);
and U13000 (N_13000,N_12928,N_12951);
or U13001 (N_13001,N_12966,N_12841);
or U13002 (N_13002,N_12782,N_12906);
nor U13003 (N_13003,N_12919,N_12950);
or U13004 (N_13004,N_12880,N_12959);
or U13005 (N_13005,N_12971,N_12778);
xnor U13006 (N_13006,N_12922,N_12877);
nor U13007 (N_13007,N_12903,N_12752);
xnor U13008 (N_13008,N_12861,N_12767);
and U13009 (N_13009,N_12977,N_12917);
nand U13010 (N_13010,N_12982,N_12780);
nor U13011 (N_13011,N_12965,N_12945);
nand U13012 (N_13012,N_12825,N_12975);
nand U13013 (N_13013,N_12785,N_12762);
xor U13014 (N_13014,N_12800,N_12827);
and U13015 (N_13015,N_12949,N_12924);
xor U13016 (N_13016,N_12986,N_12957);
or U13017 (N_13017,N_12769,N_12952);
and U13018 (N_13018,N_12820,N_12777);
xor U13019 (N_13019,N_12878,N_12842);
or U13020 (N_13020,N_12974,N_12870);
nor U13021 (N_13021,N_12997,N_12864);
xnor U13022 (N_13022,N_12942,N_12940);
nor U13023 (N_13023,N_12858,N_12969);
or U13024 (N_13024,N_12930,N_12756);
xor U13025 (N_13025,N_12863,N_12988);
and U13026 (N_13026,N_12753,N_12933);
or U13027 (N_13027,N_12781,N_12879);
xnor U13028 (N_13028,N_12811,N_12958);
nand U13029 (N_13029,N_12758,N_12770);
nor U13030 (N_13030,N_12771,N_12768);
and U13031 (N_13031,N_12983,N_12794);
xnor U13032 (N_13032,N_12885,N_12775);
nand U13033 (N_13033,N_12833,N_12995);
nand U13034 (N_13034,N_12801,N_12984);
nor U13035 (N_13035,N_12844,N_12886);
and U13036 (N_13036,N_12943,N_12809);
or U13037 (N_13037,N_12978,N_12750);
nor U13038 (N_13038,N_12865,N_12876);
and U13039 (N_13039,N_12921,N_12896);
xor U13040 (N_13040,N_12979,N_12760);
nand U13041 (N_13041,N_12815,N_12916);
nor U13042 (N_13042,N_12790,N_12889);
nor U13043 (N_13043,N_12985,N_12776);
xor U13044 (N_13044,N_12754,N_12956);
xnor U13045 (N_13045,N_12828,N_12838);
nand U13046 (N_13046,N_12802,N_12935);
xnor U13047 (N_13047,N_12901,N_12970);
and U13048 (N_13048,N_12837,N_12929);
nor U13049 (N_13049,N_12783,N_12938);
and U13050 (N_13050,N_12867,N_12796);
nor U13051 (N_13051,N_12751,N_12766);
xor U13052 (N_13052,N_12994,N_12991);
nor U13053 (N_13053,N_12947,N_12926);
and U13054 (N_13054,N_12845,N_12850);
nor U13055 (N_13055,N_12772,N_12904);
or U13056 (N_13056,N_12869,N_12789);
nor U13057 (N_13057,N_12819,N_12999);
nand U13058 (N_13058,N_12773,N_12996);
xnor U13059 (N_13059,N_12774,N_12804);
and U13060 (N_13060,N_12787,N_12962);
or U13061 (N_13061,N_12854,N_12909);
nor U13062 (N_13062,N_12972,N_12927);
xnor U13063 (N_13063,N_12799,N_12963);
and U13064 (N_13064,N_12814,N_12873);
nand U13065 (N_13065,N_12797,N_12792);
nor U13066 (N_13066,N_12857,N_12791);
and U13067 (N_13067,N_12853,N_12846);
xnor U13068 (N_13068,N_12887,N_12973);
xor U13069 (N_13069,N_12918,N_12840);
or U13070 (N_13070,N_12891,N_12788);
nor U13071 (N_13071,N_12831,N_12807);
nand U13072 (N_13072,N_12968,N_12824);
xnor U13073 (N_13073,N_12875,N_12786);
nor U13074 (N_13074,N_12868,N_12843);
nor U13075 (N_13075,N_12907,N_12855);
and U13076 (N_13076,N_12905,N_12798);
or U13077 (N_13077,N_12884,N_12953);
xor U13078 (N_13078,N_12849,N_12939);
and U13079 (N_13079,N_12765,N_12893);
nand U13080 (N_13080,N_12960,N_12888);
and U13081 (N_13081,N_12941,N_12822);
and U13082 (N_13082,N_12912,N_12852);
xor U13083 (N_13083,N_12899,N_12881);
nand U13084 (N_13084,N_12818,N_12764);
nand U13085 (N_13085,N_12931,N_12755);
nand U13086 (N_13086,N_12761,N_12836);
or U13087 (N_13087,N_12910,N_12954);
nand U13088 (N_13088,N_12872,N_12859);
or U13089 (N_13089,N_12961,N_12976);
nand U13090 (N_13090,N_12900,N_12810);
xor U13091 (N_13091,N_12848,N_12812);
nor U13092 (N_13092,N_12808,N_12894);
and U13093 (N_13093,N_12993,N_12832);
or U13094 (N_13094,N_12882,N_12989);
and U13095 (N_13095,N_12817,N_12805);
and U13096 (N_13096,N_12937,N_12839);
nor U13097 (N_13097,N_12990,N_12793);
and U13098 (N_13098,N_12874,N_12829);
nand U13099 (N_13099,N_12914,N_12892);
xor U13100 (N_13100,N_12944,N_12923);
nand U13101 (N_13101,N_12898,N_12826);
nor U13102 (N_13102,N_12908,N_12823);
nand U13103 (N_13103,N_12757,N_12934);
nand U13104 (N_13104,N_12998,N_12948);
or U13105 (N_13105,N_12834,N_12890);
or U13106 (N_13106,N_12946,N_12911);
nor U13107 (N_13107,N_12806,N_12897);
or U13108 (N_13108,N_12795,N_12992);
or U13109 (N_13109,N_12830,N_12920);
nand U13110 (N_13110,N_12763,N_12835);
and U13111 (N_13111,N_12851,N_12980);
nand U13112 (N_13112,N_12821,N_12932);
nand U13113 (N_13113,N_12967,N_12803);
nand U13114 (N_13114,N_12871,N_12759);
and U13115 (N_13115,N_12866,N_12779);
nor U13116 (N_13116,N_12936,N_12987);
and U13117 (N_13117,N_12981,N_12964);
or U13118 (N_13118,N_12925,N_12915);
nor U13119 (N_13119,N_12883,N_12856);
or U13120 (N_13120,N_12895,N_12816);
xnor U13121 (N_13121,N_12913,N_12902);
nor U13122 (N_13122,N_12955,N_12860);
xnor U13123 (N_13123,N_12862,N_12784);
or U13124 (N_13124,N_12847,N_12813);
or U13125 (N_13125,N_12939,N_12756);
nor U13126 (N_13126,N_12950,N_12883);
or U13127 (N_13127,N_12882,N_12970);
and U13128 (N_13128,N_12853,N_12912);
and U13129 (N_13129,N_12869,N_12756);
or U13130 (N_13130,N_12911,N_12880);
xnor U13131 (N_13131,N_12994,N_12838);
xnor U13132 (N_13132,N_12916,N_12937);
and U13133 (N_13133,N_12756,N_12813);
or U13134 (N_13134,N_12910,N_12871);
or U13135 (N_13135,N_12855,N_12952);
or U13136 (N_13136,N_12851,N_12798);
or U13137 (N_13137,N_12825,N_12848);
and U13138 (N_13138,N_12972,N_12768);
and U13139 (N_13139,N_12986,N_12887);
nor U13140 (N_13140,N_12879,N_12753);
or U13141 (N_13141,N_12845,N_12907);
and U13142 (N_13142,N_12796,N_12864);
xnor U13143 (N_13143,N_12814,N_12898);
nand U13144 (N_13144,N_12759,N_12770);
or U13145 (N_13145,N_12787,N_12837);
and U13146 (N_13146,N_12793,N_12770);
or U13147 (N_13147,N_12964,N_12910);
or U13148 (N_13148,N_12777,N_12963);
nand U13149 (N_13149,N_12755,N_12995);
or U13150 (N_13150,N_12829,N_12826);
nand U13151 (N_13151,N_12761,N_12903);
or U13152 (N_13152,N_12885,N_12906);
nor U13153 (N_13153,N_12886,N_12869);
nand U13154 (N_13154,N_12851,N_12959);
or U13155 (N_13155,N_12950,N_12763);
xnor U13156 (N_13156,N_12985,N_12873);
or U13157 (N_13157,N_12968,N_12853);
xnor U13158 (N_13158,N_12903,N_12931);
nor U13159 (N_13159,N_12888,N_12994);
xnor U13160 (N_13160,N_12971,N_12875);
and U13161 (N_13161,N_12892,N_12916);
xor U13162 (N_13162,N_12771,N_12907);
xnor U13163 (N_13163,N_12893,N_12820);
and U13164 (N_13164,N_12757,N_12752);
or U13165 (N_13165,N_12988,N_12769);
and U13166 (N_13166,N_12998,N_12888);
or U13167 (N_13167,N_12900,N_12757);
xnor U13168 (N_13168,N_12770,N_12810);
nor U13169 (N_13169,N_12950,N_12847);
and U13170 (N_13170,N_12841,N_12845);
nor U13171 (N_13171,N_12823,N_12755);
xor U13172 (N_13172,N_12764,N_12750);
nor U13173 (N_13173,N_12803,N_12840);
nor U13174 (N_13174,N_12785,N_12812);
xor U13175 (N_13175,N_12854,N_12935);
or U13176 (N_13176,N_12878,N_12825);
xnor U13177 (N_13177,N_12927,N_12974);
nand U13178 (N_13178,N_12795,N_12962);
nand U13179 (N_13179,N_12872,N_12958);
nand U13180 (N_13180,N_12862,N_12975);
nand U13181 (N_13181,N_12838,N_12791);
nor U13182 (N_13182,N_12953,N_12771);
nand U13183 (N_13183,N_12980,N_12810);
nor U13184 (N_13184,N_12850,N_12989);
or U13185 (N_13185,N_12976,N_12883);
and U13186 (N_13186,N_12875,N_12856);
nor U13187 (N_13187,N_12782,N_12927);
or U13188 (N_13188,N_12874,N_12891);
nand U13189 (N_13189,N_12896,N_12970);
nand U13190 (N_13190,N_12800,N_12882);
nor U13191 (N_13191,N_12805,N_12781);
xnor U13192 (N_13192,N_12855,N_12850);
xnor U13193 (N_13193,N_12815,N_12937);
nor U13194 (N_13194,N_12780,N_12873);
or U13195 (N_13195,N_12883,N_12816);
xnor U13196 (N_13196,N_12827,N_12912);
xor U13197 (N_13197,N_12992,N_12800);
or U13198 (N_13198,N_12962,N_12797);
and U13199 (N_13199,N_12978,N_12752);
xnor U13200 (N_13200,N_12972,N_12825);
or U13201 (N_13201,N_12811,N_12893);
nand U13202 (N_13202,N_12905,N_12928);
and U13203 (N_13203,N_12783,N_12996);
nor U13204 (N_13204,N_12791,N_12758);
or U13205 (N_13205,N_12896,N_12890);
and U13206 (N_13206,N_12809,N_12975);
xnor U13207 (N_13207,N_12893,N_12943);
and U13208 (N_13208,N_12841,N_12946);
xnor U13209 (N_13209,N_12966,N_12927);
nand U13210 (N_13210,N_12803,N_12970);
nor U13211 (N_13211,N_12979,N_12837);
nor U13212 (N_13212,N_12883,N_12945);
or U13213 (N_13213,N_12958,N_12854);
or U13214 (N_13214,N_12826,N_12794);
nand U13215 (N_13215,N_12907,N_12999);
xor U13216 (N_13216,N_12801,N_12964);
or U13217 (N_13217,N_12979,N_12768);
and U13218 (N_13218,N_12848,N_12840);
xor U13219 (N_13219,N_12981,N_12983);
nor U13220 (N_13220,N_12819,N_12920);
and U13221 (N_13221,N_12846,N_12995);
nand U13222 (N_13222,N_12998,N_12874);
nor U13223 (N_13223,N_12886,N_12833);
xor U13224 (N_13224,N_12827,N_12768);
or U13225 (N_13225,N_12863,N_12762);
xor U13226 (N_13226,N_12941,N_12781);
xnor U13227 (N_13227,N_12978,N_12942);
or U13228 (N_13228,N_12808,N_12854);
nor U13229 (N_13229,N_12907,N_12863);
or U13230 (N_13230,N_12961,N_12865);
xor U13231 (N_13231,N_12870,N_12752);
or U13232 (N_13232,N_12969,N_12827);
nand U13233 (N_13233,N_12993,N_12972);
nor U13234 (N_13234,N_12750,N_12877);
nand U13235 (N_13235,N_12923,N_12956);
and U13236 (N_13236,N_12901,N_12960);
or U13237 (N_13237,N_12770,N_12813);
or U13238 (N_13238,N_12944,N_12852);
nor U13239 (N_13239,N_12825,N_12765);
or U13240 (N_13240,N_12935,N_12923);
or U13241 (N_13241,N_12876,N_12924);
or U13242 (N_13242,N_12921,N_12801);
and U13243 (N_13243,N_12758,N_12821);
xor U13244 (N_13244,N_12922,N_12884);
and U13245 (N_13245,N_12920,N_12926);
xor U13246 (N_13246,N_12848,N_12821);
nor U13247 (N_13247,N_12893,N_12870);
nor U13248 (N_13248,N_12755,N_12849);
and U13249 (N_13249,N_12887,N_12953);
or U13250 (N_13250,N_13000,N_13161);
xor U13251 (N_13251,N_13217,N_13205);
and U13252 (N_13252,N_13175,N_13153);
nor U13253 (N_13253,N_13186,N_13201);
and U13254 (N_13254,N_13192,N_13029);
and U13255 (N_13255,N_13227,N_13133);
nand U13256 (N_13256,N_13117,N_13076);
nand U13257 (N_13257,N_13132,N_13122);
and U13258 (N_13258,N_13164,N_13069);
nor U13259 (N_13259,N_13024,N_13221);
and U13260 (N_13260,N_13085,N_13072);
xnor U13261 (N_13261,N_13015,N_13182);
xnor U13262 (N_13262,N_13229,N_13242);
and U13263 (N_13263,N_13098,N_13054);
nor U13264 (N_13264,N_13237,N_13095);
nor U13265 (N_13265,N_13119,N_13078);
or U13266 (N_13266,N_13167,N_13235);
nor U13267 (N_13267,N_13239,N_13169);
or U13268 (N_13268,N_13156,N_13089);
nand U13269 (N_13269,N_13103,N_13041);
xnor U13270 (N_13270,N_13135,N_13003);
and U13271 (N_13271,N_13203,N_13143);
xnor U13272 (N_13272,N_13097,N_13086);
nor U13273 (N_13273,N_13151,N_13130);
nand U13274 (N_13274,N_13127,N_13001);
nor U13275 (N_13275,N_13033,N_13144);
and U13276 (N_13276,N_13048,N_13163);
and U13277 (N_13277,N_13213,N_13025);
xor U13278 (N_13278,N_13050,N_13154);
nand U13279 (N_13279,N_13110,N_13188);
nand U13280 (N_13280,N_13123,N_13108);
or U13281 (N_13281,N_13241,N_13038);
nor U13282 (N_13282,N_13172,N_13109);
or U13283 (N_13283,N_13063,N_13039);
xor U13284 (N_13284,N_13114,N_13100);
nand U13285 (N_13285,N_13030,N_13136);
or U13286 (N_13286,N_13062,N_13170);
nor U13287 (N_13287,N_13007,N_13096);
nor U13288 (N_13288,N_13183,N_13075);
and U13289 (N_13289,N_13101,N_13009);
xnor U13290 (N_13290,N_13008,N_13055);
or U13291 (N_13291,N_13190,N_13247);
xor U13292 (N_13292,N_13131,N_13042);
xnor U13293 (N_13293,N_13145,N_13088);
xor U13294 (N_13294,N_13178,N_13141);
or U13295 (N_13295,N_13160,N_13134);
nor U13296 (N_13296,N_13027,N_13020);
nand U13297 (N_13297,N_13005,N_13052);
nand U13298 (N_13298,N_13112,N_13056);
nor U13299 (N_13299,N_13064,N_13120);
nand U13300 (N_13300,N_13142,N_13197);
xor U13301 (N_13301,N_13231,N_13232);
or U13302 (N_13302,N_13012,N_13196);
nor U13303 (N_13303,N_13035,N_13121);
and U13304 (N_13304,N_13073,N_13193);
and U13305 (N_13305,N_13225,N_13185);
nor U13306 (N_13306,N_13106,N_13090);
and U13307 (N_13307,N_13070,N_13199);
and U13308 (N_13308,N_13140,N_13159);
or U13309 (N_13309,N_13194,N_13236);
or U13310 (N_13310,N_13014,N_13113);
nor U13311 (N_13311,N_13066,N_13053);
and U13312 (N_13312,N_13102,N_13243);
and U13313 (N_13313,N_13176,N_13079);
nor U13314 (N_13314,N_13222,N_13223);
or U13315 (N_13315,N_13105,N_13116);
and U13316 (N_13316,N_13220,N_13040);
nand U13317 (N_13317,N_13094,N_13207);
or U13318 (N_13318,N_13084,N_13111);
and U13319 (N_13319,N_13023,N_13002);
or U13320 (N_13320,N_13034,N_13058);
xor U13321 (N_13321,N_13028,N_13139);
nor U13322 (N_13322,N_13202,N_13244);
and U13323 (N_13323,N_13204,N_13026);
nor U13324 (N_13324,N_13031,N_13045);
xor U13325 (N_13325,N_13047,N_13091);
nor U13326 (N_13326,N_13087,N_13118);
or U13327 (N_13327,N_13171,N_13226);
and U13328 (N_13328,N_13230,N_13124);
or U13329 (N_13329,N_13174,N_13157);
xor U13330 (N_13330,N_13016,N_13173);
nand U13331 (N_13331,N_13228,N_13240);
xnor U13332 (N_13332,N_13208,N_13046);
or U13333 (N_13333,N_13061,N_13082);
or U13334 (N_13334,N_13215,N_13125);
nand U13335 (N_13335,N_13150,N_13137);
nand U13336 (N_13336,N_13224,N_13099);
nor U13337 (N_13337,N_13104,N_13195);
and U13338 (N_13338,N_13074,N_13006);
xnor U13339 (N_13339,N_13148,N_13147);
or U13340 (N_13340,N_13037,N_13234);
and U13341 (N_13341,N_13107,N_13092);
nor U13342 (N_13342,N_13180,N_13013);
xor U13343 (N_13343,N_13249,N_13200);
or U13344 (N_13344,N_13032,N_13210);
and U13345 (N_13345,N_13211,N_13206);
nor U13346 (N_13346,N_13246,N_13238);
xor U13347 (N_13347,N_13218,N_13081);
xnor U13348 (N_13348,N_13017,N_13189);
nand U13349 (N_13349,N_13216,N_13093);
xor U13350 (N_13350,N_13152,N_13146);
nand U13351 (N_13351,N_13067,N_13060);
nand U13352 (N_13352,N_13128,N_13004);
xnor U13353 (N_13353,N_13065,N_13179);
xor U13354 (N_13354,N_13115,N_13245);
nand U13355 (N_13355,N_13044,N_13233);
nand U13356 (N_13356,N_13051,N_13184);
nand U13357 (N_13357,N_13149,N_13010);
xnor U13358 (N_13358,N_13129,N_13162);
nor U13359 (N_13359,N_13021,N_13018);
nand U13360 (N_13360,N_13191,N_13049);
nor U13361 (N_13361,N_13059,N_13043);
nand U13362 (N_13362,N_13138,N_13181);
nor U13363 (N_13363,N_13198,N_13212);
nor U13364 (N_13364,N_13057,N_13187);
nor U13365 (N_13365,N_13077,N_13177);
and U13366 (N_13366,N_13083,N_13158);
xor U13367 (N_13367,N_13165,N_13071);
xnor U13368 (N_13368,N_13022,N_13219);
or U13369 (N_13369,N_13068,N_13214);
nand U13370 (N_13370,N_13036,N_13080);
xor U13371 (N_13371,N_13248,N_13155);
xnor U13372 (N_13372,N_13019,N_13126);
and U13373 (N_13373,N_13168,N_13209);
nand U13374 (N_13374,N_13166,N_13011);
or U13375 (N_13375,N_13102,N_13210);
and U13376 (N_13376,N_13004,N_13046);
and U13377 (N_13377,N_13153,N_13042);
and U13378 (N_13378,N_13127,N_13160);
xor U13379 (N_13379,N_13086,N_13189);
or U13380 (N_13380,N_13215,N_13236);
and U13381 (N_13381,N_13125,N_13131);
or U13382 (N_13382,N_13070,N_13047);
nand U13383 (N_13383,N_13130,N_13071);
xor U13384 (N_13384,N_13142,N_13244);
nor U13385 (N_13385,N_13141,N_13169);
nor U13386 (N_13386,N_13152,N_13110);
or U13387 (N_13387,N_13006,N_13024);
nand U13388 (N_13388,N_13087,N_13199);
nor U13389 (N_13389,N_13161,N_13076);
and U13390 (N_13390,N_13097,N_13028);
and U13391 (N_13391,N_13156,N_13202);
or U13392 (N_13392,N_13137,N_13058);
and U13393 (N_13393,N_13190,N_13147);
and U13394 (N_13394,N_13154,N_13058);
and U13395 (N_13395,N_13242,N_13134);
nor U13396 (N_13396,N_13093,N_13143);
nand U13397 (N_13397,N_13104,N_13159);
or U13398 (N_13398,N_13005,N_13118);
nand U13399 (N_13399,N_13184,N_13176);
xor U13400 (N_13400,N_13111,N_13237);
and U13401 (N_13401,N_13190,N_13074);
or U13402 (N_13402,N_13028,N_13069);
or U13403 (N_13403,N_13033,N_13061);
nor U13404 (N_13404,N_13159,N_13045);
xnor U13405 (N_13405,N_13092,N_13203);
xnor U13406 (N_13406,N_13026,N_13179);
or U13407 (N_13407,N_13047,N_13133);
xnor U13408 (N_13408,N_13060,N_13035);
nand U13409 (N_13409,N_13007,N_13202);
nor U13410 (N_13410,N_13192,N_13174);
nor U13411 (N_13411,N_13244,N_13039);
nand U13412 (N_13412,N_13148,N_13195);
and U13413 (N_13413,N_13241,N_13118);
nand U13414 (N_13414,N_13188,N_13032);
nor U13415 (N_13415,N_13038,N_13229);
xnor U13416 (N_13416,N_13056,N_13192);
xnor U13417 (N_13417,N_13009,N_13148);
nor U13418 (N_13418,N_13030,N_13204);
xor U13419 (N_13419,N_13226,N_13118);
nand U13420 (N_13420,N_13106,N_13104);
xnor U13421 (N_13421,N_13014,N_13190);
or U13422 (N_13422,N_13204,N_13242);
and U13423 (N_13423,N_13218,N_13100);
xnor U13424 (N_13424,N_13065,N_13206);
nor U13425 (N_13425,N_13100,N_13191);
nand U13426 (N_13426,N_13077,N_13116);
nand U13427 (N_13427,N_13118,N_13218);
nand U13428 (N_13428,N_13082,N_13174);
or U13429 (N_13429,N_13193,N_13029);
nand U13430 (N_13430,N_13099,N_13214);
xor U13431 (N_13431,N_13005,N_13150);
xor U13432 (N_13432,N_13217,N_13027);
and U13433 (N_13433,N_13048,N_13026);
and U13434 (N_13434,N_13149,N_13039);
or U13435 (N_13435,N_13239,N_13154);
nor U13436 (N_13436,N_13066,N_13178);
xnor U13437 (N_13437,N_13024,N_13178);
nor U13438 (N_13438,N_13223,N_13057);
or U13439 (N_13439,N_13168,N_13029);
and U13440 (N_13440,N_13064,N_13011);
xor U13441 (N_13441,N_13238,N_13120);
and U13442 (N_13442,N_13043,N_13079);
nand U13443 (N_13443,N_13182,N_13226);
nor U13444 (N_13444,N_13001,N_13122);
nand U13445 (N_13445,N_13195,N_13047);
and U13446 (N_13446,N_13080,N_13045);
xor U13447 (N_13447,N_13164,N_13201);
nor U13448 (N_13448,N_13175,N_13015);
and U13449 (N_13449,N_13068,N_13230);
xnor U13450 (N_13450,N_13173,N_13218);
nand U13451 (N_13451,N_13006,N_13203);
nor U13452 (N_13452,N_13096,N_13102);
nor U13453 (N_13453,N_13045,N_13203);
and U13454 (N_13454,N_13039,N_13003);
xnor U13455 (N_13455,N_13074,N_13185);
nor U13456 (N_13456,N_13025,N_13086);
or U13457 (N_13457,N_13211,N_13123);
xor U13458 (N_13458,N_13201,N_13057);
nand U13459 (N_13459,N_13115,N_13024);
nand U13460 (N_13460,N_13103,N_13063);
or U13461 (N_13461,N_13083,N_13150);
or U13462 (N_13462,N_13041,N_13164);
and U13463 (N_13463,N_13005,N_13241);
nor U13464 (N_13464,N_13050,N_13228);
nand U13465 (N_13465,N_13079,N_13141);
nor U13466 (N_13466,N_13240,N_13170);
nand U13467 (N_13467,N_13090,N_13111);
and U13468 (N_13468,N_13049,N_13133);
nand U13469 (N_13469,N_13164,N_13071);
nand U13470 (N_13470,N_13068,N_13039);
nor U13471 (N_13471,N_13009,N_13225);
nor U13472 (N_13472,N_13194,N_13158);
nand U13473 (N_13473,N_13004,N_13247);
or U13474 (N_13474,N_13204,N_13077);
nand U13475 (N_13475,N_13188,N_13091);
or U13476 (N_13476,N_13081,N_13133);
or U13477 (N_13477,N_13069,N_13011);
xor U13478 (N_13478,N_13225,N_13117);
or U13479 (N_13479,N_13190,N_13241);
and U13480 (N_13480,N_13147,N_13031);
nand U13481 (N_13481,N_13144,N_13041);
or U13482 (N_13482,N_13046,N_13144);
or U13483 (N_13483,N_13231,N_13021);
nor U13484 (N_13484,N_13038,N_13067);
nand U13485 (N_13485,N_13229,N_13149);
nand U13486 (N_13486,N_13168,N_13141);
xnor U13487 (N_13487,N_13065,N_13137);
or U13488 (N_13488,N_13112,N_13201);
or U13489 (N_13489,N_13032,N_13225);
nand U13490 (N_13490,N_13165,N_13164);
and U13491 (N_13491,N_13083,N_13192);
and U13492 (N_13492,N_13138,N_13199);
and U13493 (N_13493,N_13196,N_13209);
nand U13494 (N_13494,N_13080,N_13009);
and U13495 (N_13495,N_13187,N_13102);
nor U13496 (N_13496,N_13192,N_13181);
nor U13497 (N_13497,N_13115,N_13042);
or U13498 (N_13498,N_13201,N_13110);
or U13499 (N_13499,N_13200,N_13056);
xor U13500 (N_13500,N_13363,N_13418);
nand U13501 (N_13501,N_13285,N_13432);
or U13502 (N_13502,N_13499,N_13453);
xnor U13503 (N_13503,N_13483,N_13258);
nor U13504 (N_13504,N_13484,N_13352);
nand U13505 (N_13505,N_13402,N_13326);
nor U13506 (N_13506,N_13403,N_13423);
or U13507 (N_13507,N_13472,N_13496);
nor U13508 (N_13508,N_13276,N_13444);
xnor U13509 (N_13509,N_13489,N_13293);
xnor U13510 (N_13510,N_13350,N_13333);
or U13511 (N_13511,N_13473,N_13411);
and U13512 (N_13512,N_13306,N_13260);
nand U13513 (N_13513,N_13421,N_13440);
or U13514 (N_13514,N_13450,N_13365);
nand U13515 (N_13515,N_13284,N_13275);
or U13516 (N_13516,N_13349,N_13386);
xnor U13517 (N_13517,N_13491,N_13289);
nor U13518 (N_13518,N_13255,N_13351);
or U13519 (N_13519,N_13320,N_13266);
xnor U13520 (N_13520,N_13252,N_13474);
and U13521 (N_13521,N_13318,N_13341);
nor U13522 (N_13522,N_13441,N_13494);
nand U13523 (N_13523,N_13420,N_13455);
and U13524 (N_13524,N_13353,N_13267);
nor U13525 (N_13525,N_13378,N_13456);
nor U13526 (N_13526,N_13467,N_13437);
nand U13527 (N_13527,N_13407,N_13305);
nor U13528 (N_13528,N_13254,N_13303);
or U13529 (N_13529,N_13443,N_13395);
and U13530 (N_13530,N_13463,N_13417);
and U13531 (N_13531,N_13493,N_13292);
nand U13532 (N_13532,N_13488,N_13259);
or U13533 (N_13533,N_13355,N_13253);
or U13534 (N_13534,N_13464,N_13412);
xor U13535 (N_13535,N_13283,N_13358);
or U13536 (N_13536,N_13366,N_13497);
and U13537 (N_13537,N_13398,N_13448);
nand U13538 (N_13538,N_13416,N_13406);
or U13539 (N_13539,N_13310,N_13291);
xor U13540 (N_13540,N_13446,N_13466);
nand U13541 (N_13541,N_13277,N_13287);
nand U13542 (N_13542,N_13390,N_13449);
and U13543 (N_13543,N_13486,N_13377);
nand U13544 (N_13544,N_13382,N_13263);
xnor U13545 (N_13545,N_13317,N_13470);
nor U13546 (N_13546,N_13435,N_13313);
nor U13547 (N_13547,N_13451,N_13408);
xor U13548 (N_13548,N_13401,N_13279);
xnor U13549 (N_13549,N_13281,N_13389);
nor U13550 (N_13550,N_13273,N_13274);
nand U13551 (N_13551,N_13300,N_13307);
nor U13552 (N_13552,N_13354,N_13415);
and U13553 (N_13553,N_13337,N_13471);
xor U13554 (N_13554,N_13301,N_13459);
or U13555 (N_13555,N_13438,N_13309);
xor U13556 (N_13556,N_13469,N_13481);
xor U13557 (N_13557,N_13344,N_13297);
nor U13558 (N_13558,N_13330,N_13323);
xnor U13559 (N_13559,N_13314,N_13371);
xor U13560 (N_13560,N_13348,N_13397);
and U13561 (N_13561,N_13261,N_13328);
or U13562 (N_13562,N_13270,N_13422);
and U13563 (N_13563,N_13356,N_13280);
or U13564 (N_13564,N_13431,N_13278);
nand U13565 (N_13565,N_13321,N_13383);
xor U13566 (N_13566,N_13414,N_13370);
xor U13567 (N_13567,N_13476,N_13428);
or U13568 (N_13568,N_13394,N_13250);
or U13569 (N_13569,N_13294,N_13399);
xnor U13570 (N_13570,N_13327,N_13374);
nand U13571 (N_13571,N_13329,N_13480);
nor U13572 (N_13572,N_13485,N_13482);
xor U13573 (N_13573,N_13458,N_13282);
xnor U13574 (N_13574,N_13339,N_13434);
and U13575 (N_13575,N_13302,N_13460);
nand U13576 (N_13576,N_13495,N_13465);
and U13577 (N_13577,N_13332,N_13359);
nand U13578 (N_13578,N_13430,N_13338);
nand U13579 (N_13579,N_13436,N_13396);
and U13580 (N_13580,N_13319,N_13295);
or U13581 (N_13581,N_13375,N_13308);
xor U13582 (N_13582,N_13312,N_13268);
xor U13583 (N_13583,N_13311,N_13478);
and U13584 (N_13584,N_13296,N_13335);
nor U13585 (N_13585,N_13316,N_13269);
xor U13586 (N_13586,N_13424,N_13343);
and U13587 (N_13587,N_13299,N_13409);
nor U13588 (N_13588,N_13479,N_13257);
and U13589 (N_13589,N_13393,N_13360);
or U13590 (N_13590,N_13380,N_13388);
xnor U13591 (N_13591,N_13367,N_13404);
nand U13592 (N_13592,N_13454,N_13304);
nor U13593 (N_13593,N_13251,N_13410);
nor U13594 (N_13594,N_13419,N_13413);
nand U13595 (N_13595,N_13265,N_13357);
nor U13596 (N_13596,N_13264,N_13361);
xnor U13597 (N_13597,N_13271,N_13364);
nor U13598 (N_13598,N_13381,N_13315);
nand U13599 (N_13599,N_13468,N_13452);
nor U13600 (N_13600,N_13445,N_13256);
xnor U13601 (N_13601,N_13324,N_13325);
and U13602 (N_13602,N_13272,N_13447);
nand U13603 (N_13603,N_13345,N_13427);
or U13604 (N_13604,N_13368,N_13346);
nand U13605 (N_13605,N_13492,N_13405);
nand U13606 (N_13606,N_13334,N_13487);
or U13607 (N_13607,N_13387,N_13376);
or U13608 (N_13608,N_13462,N_13439);
nand U13609 (N_13609,N_13331,N_13372);
or U13610 (N_13610,N_13426,N_13457);
and U13611 (N_13611,N_13347,N_13392);
xnor U13612 (N_13612,N_13429,N_13433);
nor U13613 (N_13613,N_13340,N_13384);
xnor U13614 (N_13614,N_13400,N_13477);
or U13615 (N_13615,N_13391,N_13262);
nand U13616 (N_13616,N_13475,N_13362);
and U13617 (N_13617,N_13385,N_13342);
xnor U13618 (N_13618,N_13461,N_13286);
nand U13619 (N_13619,N_13425,N_13442);
and U13620 (N_13620,N_13379,N_13322);
nand U13621 (N_13621,N_13298,N_13336);
or U13622 (N_13622,N_13373,N_13490);
nand U13623 (N_13623,N_13498,N_13288);
nand U13624 (N_13624,N_13369,N_13290);
xor U13625 (N_13625,N_13434,N_13253);
nor U13626 (N_13626,N_13411,N_13361);
nor U13627 (N_13627,N_13477,N_13344);
and U13628 (N_13628,N_13303,N_13353);
and U13629 (N_13629,N_13434,N_13287);
nand U13630 (N_13630,N_13487,N_13308);
nand U13631 (N_13631,N_13415,N_13428);
nand U13632 (N_13632,N_13471,N_13498);
xor U13633 (N_13633,N_13407,N_13454);
xnor U13634 (N_13634,N_13335,N_13475);
nand U13635 (N_13635,N_13480,N_13398);
and U13636 (N_13636,N_13433,N_13397);
xor U13637 (N_13637,N_13490,N_13473);
or U13638 (N_13638,N_13377,N_13265);
nand U13639 (N_13639,N_13346,N_13479);
nor U13640 (N_13640,N_13448,N_13343);
or U13641 (N_13641,N_13311,N_13337);
nand U13642 (N_13642,N_13400,N_13436);
or U13643 (N_13643,N_13303,N_13374);
xor U13644 (N_13644,N_13492,N_13281);
xnor U13645 (N_13645,N_13391,N_13426);
or U13646 (N_13646,N_13461,N_13483);
and U13647 (N_13647,N_13426,N_13386);
xnor U13648 (N_13648,N_13487,N_13372);
nand U13649 (N_13649,N_13254,N_13409);
nand U13650 (N_13650,N_13458,N_13366);
nor U13651 (N_13651,N_13454,N_13270);
and U13652 (N_13652,N_13485,N_13407);
nor U13653 (N_13653,N_13386,N_13336);
or U13654 (N_13654,N_13309,N_13310);
xor U13655 (N_13655,N_13253,N_13358);
nor U13656 (N_13656,N_13425,N_13348);
and U13657 (N_13657,N_13289,N_13261);
xnor U13658 (N_13658,N_13348,N_13358);
xor U13659 (N_13659,N_13275,N_13303);
or U13660 (N_13660,N_13415,N_13265);
nor U13661 (N_13661,N_13359,N_13255);
nor U13662 (N_13662,N_13363,N_13448);
nand U13663 (N_13663,N_13370,N_13476);
and U13664 (N_13664,N_13370,N_13380);
nand U13665 (N_13665,N_13320,N_13439);
and U13666 (N_13666,N_13307,N_13444);
xor U13667 (N_13667,N_13460,N_13328);
or U13668 (N_13668,N_13265,N_13260);
xor U13669 (N_13669,N_13438,N_13319);
xor U13670 (N_13670,N_13476,N_13349);
nand U13671 (N_13671,N_13286,N_13492);
nand U13672 (N_13672,N_13401,N_13291);
nand U13673 (N_13673,N_13285,N_13476);
nand U13674 (N_13674,N_13271,N_13253);
xnor U13675 (N_13675,N_13334,N_13406);
or U13676 (N_13676,N_13475,N_13304);
xnor U13677 (N_13677,N_13396,N_13488);
nor U13678 (N_13678,N_13281,N_13480);
nor U13679 (N_13679,N_13298,N_13432);
nand U13680 (N_13680,N_13455,N_13260);
and U13681 (N_13681,N_13485,N_13278);
and U13682 (N_13682,N_13320,N_13387);
xnor U13683 (N_13683,N_13411,N_13352);
and U13684 (N_13684,N_13353,N_13488);
or U13685 (N_13685,N_13411,N_13333);
nor U13686 (N_13686,N_13311,N_13397);
xor U13687 (N_13687,N_13422,N_13341);
or U13688 (N_13688,N_13405,N_13452);
nand U13689 (N_13689,N_13454,N_13317);
and U13690 (N_13690,N_13344,N_13408);
nor U13691 (N_13691,N_13287,N_13305);
xnor U13692 (N_13692,N_13441,N_13348);
nand U13693 (N_13693,N_13269,N_13255);
or U13694 (N_13694,N_13348,N_13257);
or U13695 (N_13695,N_13459,N_13469);
and U13696 (N_13696,N_13274,N_13433);
nor U13697 (N_13697,N_13447,N_13264);
nand U13698 (N_13698,N_13287,N_13361);
nor U13699 (N_13699,N_13371,N_13445);
nand U13700 (N_13700,N_13481,N_13443);
nor U13701 (N_13701,N_13391,N_13361);
nand U13702 (N_13702,N_13362,N_13470);
xnor U13703 (N_13703,N_13449,N_13436);
nand U13704 (N_13704,N_13353,N_13367);
nor U13705 (N_13705,N_13406,N_13370);
nand U13706 (N_13706,N_13463,N_13441);
and U13707 (N_13707,N_13449,N_13464);
xnor U13708 (N_13708,N_13365,N_13346);
nor U13709 (N_13709,N_13262,N_13455);
nor U13710 (N_13710,N_13386,N_13422);
nor U13711 (N_13711,N_13369,N_13446);
nor U13712 (N_13712,N_13326,N_13322);
or U13713 (N_13713,N_13383,N_13363);
and U13714 (N_13714,N_13303,N_13468);
nor U13715 (N_13715,N_13499,N_13254);
nor U13716 (N_13716,N_13362,N_13363);
xnor U13717 (N_13717,N_13323,N_13386);
nor U13718 (N_13718,N_13284,N_13445);
nor U13719 (N_13719,N_13467,N_13341);
nand U13720 (N_13720,N_13465,N_13481);
nor U13721 (N_13721,N_13259,N_13420);
and U13722 (N_13722,N_13402,N_13412);
nor U13723 (N_13723,N_13444,N_13381);
nor U13724 (N_13724,N_13306,N_13359);
nor U13725 (N_13725,N_13365,N_13435);
and U13726 (N_13726,N_13348,N_13365);
nor U13727 (N_13727,N_13429,N_13254);
nand U13728 (N_13728,N_13329,N_13494);
nand U13729 (N_13729,N_13379,N_13456);
xnor U13730 (N_13730,N_13376,N_13250);
and U13731 (N_13731,N_13408,N_13411);
xnor U13732 (N_13732,N_13338,N_13388);
or U13733 (N_13733,N_13438,N_13408);
nor U13734 (N_13734,N_13399,N_13426);
nor U13735 (N_13735,N_13300,N_13385);
xnor U13736 (N_13736,N_13456,N_13418);
or U13737 (N_13737,N_13330,N_13259);
or U13738 (N_13738,N_13257,N_13419);
and U13739 (N_13739,N_13267,N_13452);
nor U13740 (N_13740,N_13360,N_13327);
xor U13741 (N_13741,N_13326,N_13293);
nand U13742 (N_13742,N_13300,N_13299);
xnor U13743 (N_13743,N_13455,N_13288);
or U13744 (N_13744,N_13434,N_13457);
xnor U13745 (N_13745,N_13290,N_13392);
and U13746 (N_13746,N_13402,N_13449);
or U13747 (N_13747,N_13297,N_13354);
nor U13748 (N_13748,N_13299,N_13292);
xnor U13749 (N_13749,N_13409,N_13317);
or U13750 (N_13750,N_13647,N_13628);
xor U13751 (N_13751,N_13717,N_13700);
nand U13752 (N_13752,N_13694,N_13731);
and U13753 (N_13753,N_13719,N_13609);
nand U13754 (N_13754,N_13570,N_13699);
and U13755 (N_13755,N_13621,N_13691);
nand U13756 (N_13756,N_13692,N_13655);
nor U13757 (N_13757,N_13744,N_13687);
xor U13758 (N_13758,N_13522,N_13681);
nor U13759 (N_13759,N_13510,N_13605);
or U13760 (N_13760,N_13579,N_13586);
and U13761 (N_13761,N_13512,N_13627);
or U13762 (N_13762,N_13593,N_13653);
nor U13763 (N_13763,N_13544,N_13583);
xor U13764 (N_13764,N_13508,N_13594);
xnor U13765 (N_13765,N_13503,N_13553);
or U13766 (N_13766,N_13645,N_13701);
xor U13767 (N_13767,N_13732,N_13529);
nor U13768 (N_13768,N_13702,N_13611);
and U13769 (N_13769,N_13730,N_13704);
or U13770 (N_13770,N_13695,N_13527);
nand U13771 (N_13771,N_13632,N_13707);
xnor U13772 (N_13772,N_13690,N_13577);
nor U13773 (N_13773,N_13595,N_13603);
nor U13774 (N_13774,N_13662,N_13580);
or U13775 (N_13775,N_13743,N_13604);
and U13776 (N_13776,N_13502,N_13693);
nand U13777 (N_13777,N_13539,N_13623);
and U13778 (N_13778,N_13741,N_13723);
xnor U13779 (N_13779,N_13726,N_13557);
nand U13780 (N_13780,N_13561,N_13716);
and U13781 (N_13781,N_13651,N_13598);
and U13782 (N_13782,N_13516,N_13549);
and U13783 (N_13783,N_13520,N_13616);
xnor U13784 (N_13784,N_13547,N_13633);
or U13785 (N_13785,N_13737,N_13740);
and U13786 (N_13786,N_13565,N_13559);
nand U13787 (N_13787,N_13518,N_13703);
and U13788 (N_13788,N_13688,N_13531);
nand U13789 (N_13789,N_13711,N_13713);
nand U13790 (N_13790,N_13663,N_13513);
nor U13791 (N_13791,N_13581,N_13708);
or U13792 (N_13792,N_13501,N_13601);
or U13793 (N_13793,N_13666,N_13721);
or U13794 (N_13794,N_13641,N_13536);
nor U13795 (N_13795,N_13685,N_13587);
xnor U13796 (N_13796,N_13667,N_13618);
and U13797 (N_13797,N_13550,N_13571);
and U13798 (N_13798,N_13673,N_13639);
nor U13799 (N_13799,N_13634,N_13626);
xnor U13800 (N_13800,N_13686,N_13665);
nor U13801 (N_13801,N_13541,N_13588);
xor U13802 (N_13802,N_13567,N_13675);
and U13803 (N_13803,N_13552,N_13555);
nor U13804 (N_13804,N_13505,N_13504);
nor U13805 (N_13805,N_13709,N_13537);
nand U13806 (N_13806,N_13568,N_13602);
and U13807 (N_13807,N_13696,N_13720);
nor U13808 (N_13808,N_13674,N_13620);
nor U13809 (N_13809,N_13680,N_13728);
nor U13810 (N_13810,N_13683,N_13551);
nand U13811 (N_13811,N_13671,N_13715);
nor U13812 (N_13812,N_13742,N_13644);
nand U13813 (N_13813,N_13507,N_13676);
or U13814 (N_13814,N_13535,N_13657);
xor U13815 (N_13815,N_13722,N_13625);
nand U13816 (N_13816,N_13534,N_13624);
nand U13817 (N_13817,N_13519,N_13573);
nor U13818 (N_13818,N_13714,N_13533);
xor U13819 (N_13819,N_13727,N_13562);
or U13820 (N_13820,N_13545,N_13643);
xnor U13821 (N_13821,N_13725,N_13649);
and U13822 (N_13822,N_13660,N_13556);
nand U13823 (N_13823,N_13566,N_13540);
xor U13824 (N_13824,N_13615,N_13614);
nand U13825 (N_13825,N_13637,N_13613);
or U13826 (N_13826,N_13622,N_13697);
and U13827 (N_13827,N_13659,N_13589);
nor U13828 (N_13828,N_13523,N_13747);
nor U13829 (N_13829,N_13650,N_13608);
xor U13830 (N_13830,N_13664,N_13739);
nand U13831 (N_13831,N_13724,N_13712);
and U13832 (N_13832,N_13576,N_13590);
nor U13833 (N_13833,N_13517,N_13546);
nor U13834 (N_13834,N_13642,N_13554);
xnor U13835 (N_13835,N_13705,N_13630);
nand U13836 (N_13836,N_13746,N_13738);
xnor U13837 (N_13837,N_13654,N_13569);
nor U13838 (N_13838,N_13733,N_13572);
or U13839 (N_13839,N_13631,N_13735);
xor U13840 (N_13840,N_13564,N_13668);
and U13841 (N_13841,N_13525,N_13682);
and U13842 (N_13842,N_13584,N_13689);
and U13843 (N_13843,N_13607,N_13524);
xor U13844 (N_13844,N_13652,N_13582);
nand U13845 (N_13845,N_13585,N_13619);
and U13846 (N_13846,N_13574,N_13748);
nand U13847 (N_13847,N_13543,N_13736);
and U13848 (N_13848,N_13526,N_13677);
xor U13849 (N_13849,N_13679,N_13538);
nand U13850 (N_13850,N_13597,N_13500);
nor U13851 (N_13851,N_13734,N_13656);
or U13852 (N_13852,N_13636,N_13710);
nor U13853 (N_13853,N_13646,N_13640);
and U13854 (N_13854,N_13617,N_13591);
or U13855 (N_13855,N_13606,N_13706);
xor U13856 (N_13856,N_13521,N_13729);
nand U13857 (N_13857,N_13575,N_13530);
xor U13858 (N_13858,N_13749,N_13684);
nor U13859 (N_13859,N_13648,N_13592);
and U13860 (N_13860,N_13599,N_13718);
nand U13861 (N_13861,N_13511,N_13672);
nand U13862 (N_13862,N_13745,N_13506);
xor U13863 (N_13863,N_13542,N_13638);
or U13864 (N_13864,N_13532,N_13669);
nand U13865 (N_13865,N_13610,N_13514);
nand U13866 (N_13866,N_13515,N_13629);
nor U13867 (N_13867,N_13528,N_13548);
or U13868 (N_13868,N_13596,N_13509);
nor U13869 (N_13869,N_13578,N_13661);
and U13870 (N_13870,N_13560,N_13678);
and U13871 (N_13871,N_13658,N_13600);
nor U13872 (N_13872,N_13698,N_13670);
nor U13873 (N_13873,N_13612,N_13563);
nand U13874 (N_13874,N_13635,N_13558);
nand U13875 (N_13875,N_13739,N_13717);
and U13876 (N_13876,N_13549,N_13669);
nand U13877 (N_13877,N_13569,N_13521);
nand U13878 (N_13878,N_13663,N_13525);
xor U13879 (N_13879,N_13649,N_13676);
xor U13880 (N_13880,N_13645,N_13511);
xor U13881 (N_13881,N_13569,N_13709);
xnor U13882 (N_13882,N_13510,N_13742);
nor U13883 (N_13883,N_13709,N_13583);
or U13884 (N_13884,N_13612,N_13562);
or U13885 (N_13885,N_13615,N_13503);
xor U13886 (N_13886,N_13582,N_13511);
nor U13887 (N_13887,N_13734,N_13537);
and U13888 (N_13888,N_13630,N_13681);
and U13889 (N_13889,N_13658,N_13615);
and U13890 (N_13890,N_13745,N_13737);
nor U13891 (N_13891,N_13719,N_13661);
xnor U13892 (N_13892,N_13635,N_13580);
or U13893 (N_13893,N_13551,N_13687);
and U13894 (N_13894,N_13728,N_13556);
nand U13895 (N_13895,N_13739,N_13707);
xor U13896 (N_13896,N_13523,N_13536);
and U13897 (N_13897,N_13508,N_13657);
and U13898 (N_13898,N_13609,N_13500);
and U13899 (N_13899,N_13677,N_13722);
and U13900 (N_13900,N_13748,N_13653);
or U13901 (N_13901,N_13728,N_13659);
nor U13902 (N_13902,N_13528,N_13723);
and U13903 (N_13903,N_13678,N_13721);
nand U13904 (N_13904,N_13632,N_13702);
xnor U13905 (N_13905,N_13742,N_13592);
or U13906 (N_13906,N_13610,N_13661);
nor U13907 (N_13907,N_13601,N_13542);
and U13908 (N_13908,N_13504,N_13548);
or U13909 (N_13909,N_13584,N_13673);
or U13910 (N_13910,N_13560,N_13650);
or U13911 (N_13911,N_13667,N_13555);
nor U13912 (N_13912,N_13554,N_13600);
xnor U13913 (N_13913,N_13689,N_13697);
nor U13914 (N_13914,N_13728,N_13713);
and U13915 (N_13915,N_13599,N_13738);
and U13916 (N_13916,N_13507,N_13663);
and U13917 (N_13917,N_13543,N_13643);
and U13918 (N_13918,N_13587,N_13749);
or U13919 (N_13919,N_13543,N_13717);
nand U13920 (N_13920,N_13569,N_13500);
xor U13921 (N_13921,N_13573,N_13694);
nand U13922 (N_13922,N_13595,N_13584);
nor U13923 (N_13923,N_13667,N_13743);
or U13924 (N_13924,N_13593,N_13701);
xor U13925 (N_13925,N_13688,N_13709);
and U13926 (N_13926,N_13604,N_13622);
xor U13927 (N_13927,N_13589,N_13699);
nor U13928 (N_13928,N_13615,N_13641);
and U13929 (N_13929,N_13578,N_13673);
nor U13930 (N_13930,N_13597,N_13681);
nand U13931 (N_13931,N_13540,N_13655);
xor U13932 (N_13932,N_13714,N_13710);
or U13933 (N_13933,N_13665,N_13667);
nand U13934 (N_13934,N_13580,N_13537);
xor U13935 (N_13935,N_13618,N_13538);
nor U13936 (N_13936,N_13564,N_13642);
xor U13937 (N_13937,N_13633,N_13715);
xnor U13938 (N_13938,N_13622,N_13693);
and U13939 (N_13939,N_13525,N_13658);
nand U13940 (N_13940,N_13589,N_13548);
and U13941 (N_13941,N_13566,N_13660);
nor U13942 (N_13942,N_13509,N_13611);
or U13943 (N_13943,N_13658,N_13597);
or U13944 (N_13944,N_13699,N_13689);
and U13945 (N_13945,N_13720,N_13563);
nand U13946 (N_13946,N_13685,N_13627);
nand U13947 (N_13947,N_13739,N_13701);
or U13948 (N_13948,N_13650,N_13545);
nor U13949 (N_13949,N_13618,N_13702);
or U13950 (N_13950,N_13727,N_13702);
xor U13951 (N_13951,N_13631,N_13557);
nand U13952 (N_13952,N_13520,N_13642);
nand U13953 (N_13953,N_13698,N_13652);
and U13954 (N_13954,N_13672,N_13670);
and U13955 (N_13955,N_13707,N_13706);
and U13956 (N_13956,N_13748,N_13515);
nor U13957 (N_13957,N_13566,N_13734);
and U13958 (N_13958,N_13590,N_13628);
and U13959 (N_13959,N_13695,N_13583);
nor U13960 (N_13960,N_13659,N_13525);
and U13961 (N_13961,N_13681,N_13544);
nand U13962 (N_13962,N_13687,N_13567);
and U13963 (N_13963,N_13607,N_13720);
xor U13964 (N_13964,N_13603,N_13693);
nor U13965 (N_13965,N_13581,N_13571);
nor U13966 (N_13966,N_13711,N_13572);
nand U13967 (N_13967,N_13567,N_13737);
nor U13968 (N_13968,N_13743,N_13725);
xor U13969 (N_13969,N_13718,N_13534);
and U13970 (N_13970,N_13554,N_13611);
nor U13971 (N_13971,N_13533,N_13518);
xnor U13972 (N_13972,N_13672,N_13714);
xor U13973 (N_13973,N_13692,N_13648);
and U13974 (N_13974,N_13591,N_13734);
xnor U13975 (N_13975,N_13653,N_13548);
or U13976 (N_13976,N_13530,N_13601);
nor U13977 (N_13977,N_13681,N_13701);
nand U13978 (N_13978,N_13690,N_13705);
xnor U13979 (N_13979,N_13687,N_13604);
nand U13980 (N_13980,N_13714,N_13590);
and U13981 (N_13981,N_13556,N_13518);
and U13982 (N_13982,N_13712,N_13501);
or U13983 (N_13983,N_13711,N_13587);
or U13984 (N_13984,N_13601,N_13650);
xor U13985 (N_13985,N_13517,N_13629);
xor U13986 (N_13986,N_13662,N_13537);
or U13987 (N_13987,N_13564,N_13734);
nand U13988 (N_13988,N_13677,N_13670);
or U13989 (N_13989,N_13515,N_13705);
and U13990 (N_13990,N_13598,N_13516);
or U13991 (N_13991,N_13543,N_13712);
or U13992 (N_13992,N_13588,N_13545);
nand U13993 (N_13993,N_13531,N_13585);
and U13994 (N_13994,N_13651,N_13621);
xor U13995 (N_13995,N_13547,N_13682);
and U13996 (N_13996,N_13662,N_13704);
nor U13997 (N_13997,N_13563,N_13583);
and U13998 (N_13998,N_13630,N_13532);
nand U13999 (N_13999,N_13593,N_13584);
or U14000 (N_14000,N_13828,N_13899);
nor U14001 (N_14001,N_13783,N_13854);
nand U14002 (N_14002,N_13755,N_13822);
nor U14003 (N_14003,N_13756,N_13971);
nand U14004 (N_14004,N_13928,N_13992);
xnor U14005 (N_14005,N_13752,N_13860);
xor U14006 (N_14006,N_13907,N_13885);
nor U14007 (N_14007,N_13897,N_13954);
or U14008 (N_14008,N_13938,N_13948);
and U14009 (N_14009,N_13989,N_13763);
or U14010 (N_14010,N_13811,N_13936);
xor U14011 (N_14011,N_13847,N_13891);
nand U14012 (N_14012,N_13888,N_13842);
or U14013 (N_14013,N_13840,N_13784);
or U14014 (N_14014,N_13799,N_13772);
or U14015 (N_14015,N_13970,N_13835);
xnor U14016 (N_14016,N_13868,N_13773);
nand U14017 (N_14017,N_13781,N_13946);
and U14018 (N_14018,N_13850,N_13941);
nor U14019 (N_14019,N_13913,N_13795);
xnor U14020 (N_14020,N_13979,N_13793);
and U14021 (N_14021,N_13757,N_13764);
and U14022 (N_14022,N_13942,N_13880);
and U14023 (N_14023,N_13873,N_13875);
nand U14024 (N_14024,N_13844,N_13762);
and U14025 (N_14025,N_13804,N_13945);
nor U14026 (N_14026,N_13914,N_13931);
nor U14027 (N_14027,N_13851,N_13751);
nand U14028 (N_14028,N_13883,N_13845);
nor U14029 (N_14029,N_13857,N_13933);
xor U14030 (N_14030,N_13944,N_13892);
and U14031 (N_14031,N_13770,N_13967);
nor U14032 (N_14032,N_13965,N_13821);
and U14033 (N_14033,N_13994,N_13940);
or U14034 (N_14034,N_13829,N_13947);
xnor U14035 (N_14035,N_13866,N_13919);
or U14036 (N_14036,N_13900,N_13916);
xor U14037 (N_14037,N_13864,N_13951);
and U14038 (N_14038,N_13797,N_13978);
xor U14039 (N_14039,N_13805,N_13846);
and U14040 (N_14040,N_13836,N_13813);
and U14041 (N_14041,N_13917,N_13780);
nand U14042 (N_14042,N_13923,N_13761);
or U14043 (N_14043,N_13801,N_13816);
and U14044 (N_14044,N_13796,N_13839);
and U14045 (N_14045,N_13779,N_13915);
nand U14046 (N_14046,N_13869,N_13910);
nand U14047 (N_14047,N_13800,N_13974);
xor U14048 (N_14048,N_13879,N_13802);
and U14049 (N_14049,N_13861,N_13814);
nor U14050 (N_14050,N_13980,N_13960);
nor U14051 (N_14051,N_13754,N_13922);
nor U14052 (N_14052,N_13912,N_13937);
xnor U14053 (N_14053,N_13849,N_13935);
and U14054 (N_14054,N_13750,N_13927);
nand U14055 (N_14055,N_13958,N_13853);
or U14056 (N_14056,N_13898,N_13848);
nand U14057 (N_14057,N_13939,N_13905);
xnor U14058 (N_14058,N_13830,N_13977);
xor U14059 (N_14059,N_13862,N_13920);
nand U14060 (N_14060,N_13906,N_13823);
xor U14061 (N_14061,N_13815,N_13966);
xnor U14062 (N_14062,N_13881,N_13981);
xor U14063 (N_14063,N_13985,N_13837);
xor U14064 (N_14064,N_13766,N_13874);
nor U14065 (N_14065,N_13918,N_13808);
nor U14066 (N_14066,N_13990,N_13925);
xor U14067 (N_14067,N_13833,N_13894);
and U14068 (N_14068,N_13759,N_13789);
or U14069 (N_14069,N_13794,N_13984);
xor U14070 (N_14070,N_13841,N_13818);
nor U14071 (N_14071,N_13953,N_13975);
or U14072 (N_14072,N_13791,N_13758);
nor U14073 (N_14073,N_13778,N_13972);
xnor U14074 (N_14074,N_13768,N_13999);
nand U14075 (N_14075,N_13950,N_13983);
or U14076 (N_14076,N_13786,N_13987);
xor U14077 (N_14077,N_13878,N_13788);
xor U14078 (N_14078,N_13902,N_13926);
and U14079 (N_14079,N_13998,N_13831);
or U14080 (N_14080,N_13996,N_13832);
nand U14081 (N_14081,N_13993,N_13803);
xor U14082 (N_14082,N_13997,N_13776);
nor U14083 (N_14083,N_13882,N_13968);
and U14084 (N_14084,N_13765,N_13790);
or U14085 (N_14085,N_13825,N_13810);
xnor U14086 (N_14086,N_13895,N_13787);
nor U14087 (N_14087,N_13884,N_13774);
nand U14088 (N_14088,N_13929,N_13976);
or U14089 (N_14089,N_13956,N_13964);
xor U14090 (N_14090,N_13932,N_13952);
nor U14091 (N_14091,N_13792,N_13855);
xnor U14092 (N_14092,N_13986,N_13871);
or U14093 (N_14093,N_13934,N_13930);
or U14094 (N_14094,N_13973,N_13896);
nor U14095 (N_14095,N_13760,N_13817);
or U14096 (N_14096,N_13807,N_13863);
xor U14097 (N_14097,N_13921,N_13812);
and U14098 (N_14098,N_13904,N_13798);
xnor U14099 (N_14099,N_13834,N_13991);
or U14100 (N_14100,N_13843,N_13911);
nand U14101 (N_14101,N_13893,N_13887);
nor U14102 (N_14102,N_13955,N_13867);
and U14103 (N_14103,N_13982,N_13753);
or U14104 (N_14104,N_13769,N_13809);
xor U14105 (N_14105,N_13819,N_13782);
xor U14106 (N_14106,N_13767,N_13943);
nor U14107 (N_14107,N_13949,N_13824);
and U14108 (N_14108,N_13872,N_13865);
xnor U14109 (N_14109,N_13771,N_13908);
nor U14110 (N_14110,N_13889,N_13959);
or U14111 (N_14111,N_13924,N_13870);
nor U14112 (N_14112,N_13826,N_13890);
and U14113 (N_14113,N_13877,N_13969);
nand U14114 (N_14114,N_13962,N_13858);
xor U14115 (N_14115,N_13909,N_13856);
or U14116 (N_14116,N_13785,N_13995);
and U14117 (N_14117,N_13852,N_13961);
nand U14118 (N_14118,N_13777,N_13859);
nand U14119 (N_14119,N_13957,N_13886);
xor U14120 (N_14120,N_13988,N_13806);
or U14121 (N_14121,N_13827,N_13775);
nor U14122 (N_14122,N_13963,N_13838);
nand U14123 (N_14123,N_13903,N_13901);
nand U14124 (N_14124,N_13876,N_13820);
and U14125 (N_14125,N_13850,N_13938);
or U14126 (N_14126,N_13790,N_13813);
nor U14127 (N_14127,N_13851,N_13901);
xnor U14128 (N_14128,N_13824,N_13940);
or U14129 (N_14129,N_13936,N_13821);
xnor U14130 (N_14130,N_13996,N_13758);
nor U14131 (N_14131,N_13953,N_13910);
nand U14132 (N_14132,N_13913,N_13783);
xnor U14133 (N_14133,N_13931,N_13972);
xor U14134 (N_14134,N_13948,N_13912);
nor U14135 (N_14135,N_13750,N_13856);
or U14136 (N_14136,N_13953,N_13962);
nor U14137 (N_14137,N_13866,N_13897);
and U14138 (N_14138,N_13993,N_13953);
and U14139 (N_14139,N_13812,N_13890);
and U14140 (N_14140,N_13815,N_13832);
nand U14141 (N_14141,N_13751,N_13779);
or U14142 (N_14142,N_13862,N_13823);
xnor U14143 (N_14143,N_13750,N_13990);
nand U14144 (N_14144,N_13807,N_13756);
and U14145 (N_14145,N_13898,N_13960);
and U14146 (N_14146,N_13769,N_13982);
nor U14147 (N_14147,N_13953,N_13760);
xnor U14148 (N_14148,N_13982,N_13938);
nand U14149 (N_14149,N_13819,N_13999);
nand U14150 (N_14150,N_13868,N_13834);
nor U14151 (N_14151,N_13932,N_13782);
and U14152 (N_14152,N_13806,N_13765);
and U14153 (N_14153,N_13891,N_13897);
nand U14154 (N_14154,N_13849,N_13797);
and U14155 (N_14155,N_13775,N_13975);
nor U14156 (N_14156,N_13803,N_13831);
or U14157 (N_14157,N_13966,N_13996);
xor U14158 (N_14158,N_13988,N_13899);
and U14159 (N_14159,N_13844,N_13956);
and U14160 (N_14160,N_13864,N_13794);
or U14161 (N_14161,N_13813,N_13763);
and U14162 (N_14162,N_13786,N_13830);
nor U14163 (N_14163,N_13815,N_13883);
nand U14164 (N_14164,N_13849,N_13961);
and U14165 (N_14165,N_13983,N_13864);
xor U14166 (N_14166,N_13832,N_13966);
nand U14167 (N_14167,N_13816,N_13924);
or U14168 (N_14168,N_13931,N_13901);
and U14169 (N_14169,N_13963,N_13937);
nand U14170 (N_14170,N_13906,N_13797);
xor U14171 (N_14171,N_13927,N_13816);
nor U14172 (N_14172,N_13970,N_13910);
or U14173 (N_14173,N_13898,N_13881);
nor U14174 (N_14174,N_13811,N_13771);
nand U14175 (N_14175,N_13872,N_13818);
nand U14176 (N_14176,N_13814,N_13759);
or U14177 (N_14177,N_13773,N_13900);
and U14178 (N_14178,N_13750,N_13821);
and U14179 (N_14179,N_13909,N_13911);
nor U14180 (N_14180,N_13991,N_13972);
xnor U14181 (N_14181,N_13779,N_13923);
and U14182 (N_14182,N_13978,N_13864);
or U14183 (N_14183,N_13878,N_13782);
xnor U14184 (N_14184,N_13799,N_13842);
or U14185 (N_14185,N_13803,N_13920);
xor U14186 (N_14186,N_13997,N_13795);
nor U14187 (N_14187,N_13816,N_13890);
xnor U14188 (N_14188,N_13894,N_13988);
xnor U14189 (N_14189,N_13994,N_13921);
nor U14190 (N_14190,N_13781,N_13772);
xor U14191 (N_14191,N_13930,N_13811);
xor U14192 (N_14192,N_13829,N_13800);
nor U14193 (N_14193,N_13808,N_13836);
or U14194 (N_14194,N_13972,N_13975);
or U14195 (N_14195,N_13969,N_13977);
nand U14196 (N_14196,N_13811,N_13971);
xor U14197 (N_14197,N_13886,N_13966);
and U14198 (N_14198,N_13860,N_13888);
or U14199 (N_14199,N_13994,N_13870);
nand U14200 (N_14200,N_13931,N_13937);
and U14201 (N_14201,N_13851,N_13754);
or U14202 (N_14202,N_13903,N_13948);
and U14203 (N_14203,N_13765,N_13877);
nor U14204 (N_14204,N_13937,N_13905);
or U14205 (N_14205,N_13808,N_13894);
xor U14206 (N_14206,N_13787,N_13772);
nor U14207 (N_14207,N_13853,N_13763);
or U14208 (N_14208,N_13953,N_13983);
nor U14209 (N_14209,N_13764,N_13849);
nor U14210 (N_14210,N_13928,N_13902);
xor U14211 (N_14211,N_13915,N_13857);
and U14212 (N_14212,N_13802,N_13906);
nor U14213 (N_14213,N_13915,N_13970);
or U14214 (N_14214,N_13763,N_13958);
or U14215 (N_14215,N_13910,N_13806);
and U14216 (N_14216,N_13777,N_13778);
or U14217 (N_14217,N_13840,N_13985);
xnor U14218 (N_14218,N_13772,N_13778);
and U14219 (N_14219,N_13864,N_13823);
nor U14220 (N_14220,N_13951,N_13866);
nand U14221 (N_14221,N_13918,N_13754);
and U14222 (N_14222,N_13891,N_13971);
nor U14223 (N_14223,N_13943,N_13899);
or U14224 (N_14224,N_13752,N_13857);
and U14225 (N_14225,N_13976,N_13969);
or U14226 (N_14226,N_13911,N_13983);
nor U14227 (N_14227,N_13875,N_13914);
and U14228 (N_14228,N_13782,N_13875);
or U14229 (N_14229,N_13807,N_13880);
nor U14230 (N_14230,N_13977,N_13874);
and U14231 (N_14231,N_13869,N_13994);
and U14232 (N_14232,N_13776,N_13952);
nor U14233 (N_14233,N_13838,N_13815);
and U14234 (N_14234,N_13863,N_13907);
nor U14235 (N_14235,N_13842,N_13795);
nand U14236 (N_14236,N_13788,N_13823);
nand U14237 (N_14237,N_13940,N_13877);
nand U14238 (N_14238,N_13875,N_13852);
nand U14239 (N_14239,N_13760,N_13946);
and U14240 (N_14240,N_13940,N_13915);
and U14241 (N_14241,N_13788,N_13753);
xnor U14242 (N_14242,N_13964,N_13867);
nand U14243 (N_14243,N_13780,N_13872);
xor U14244 (N_14244,N_13782,N_13986);
nor U14245 (N_14245,N_13853,N_13865);
or U14246 (N_14246,N_13872,N_13895);
nor U14247 (N_14247,N_13759,N_13965);
nand U14248 (N_14248,N_13769,N_13907);
and U14249 (N_14249,N_13814,N_13815);
nand U14250 (N_14250,N_14143,N_14103);
xnor U14251 (N_14251,N_14000,N_14188);
nand U14252 (N_14252,N_14136,N_14064);
nand U14253 (N_14253,N_14206,N_14031);
or U14254 (N_14254,N_14222,N_14137);
or U14255 (N_14255,N_14180,N_14027);
or U14256 (N_14256,N_14035,N_14091);
and U14257 (N_14257,N_14216,N_14032);
and U14258 (N_14258,N_14119,N_14076);
xnor U14259 (N_14259,N_14139,N_14132);
and U14260 (N_14260,N_14049,N_14108);
and U14261 (N_14261,N_14097,N_14060);
or U14262 (N_14262,N_14124,N_14195);
nand U14263 (N_14263,N_14149,N_14085);
xor U14264 (N_14264,N_14230,N_14192);
or U14265 (N_14265,N_14185,N_14219);
or U14266 (N_14266,N_14039,N_14008);
nor U14267 (N_14267,N_14156,N_14007);
xor U14268 (N_14268,N_14019,N_14067);
and U14269 (N_14269,N_14203,N_14172);
nand U14270 (N_14270,N_14109,N_14092);
nor U14271 (N_14271,N_14193,N_14022);
or U14272 (N_14272,N_14118,N_14056);
nor U14273 (N_14273,N_14051,N_14102);
nand U14274 (N_14274,N_14231,N_14248);
xnor U14275 (N_14275,N_14162,N_14227);
xor U14276 (N_14276,N_14228,N_14126);
or U14277 (N_14277,N_14199,N_14177);
or U14278 (N_14278,N_14160,N_14011);
nor U14279 (N_14279,N_14146,N_14048);
nand U14280 (N_14280,N_14190,N_14047);
xor U14281 (N_14281,N_14120,N_14043);
nor U14282 (N_14282,N_14165,N_14058);
xnor U14283 (N_14283,N_14080,N_14041);
nand U14284 (N_14284,N_14096,N_14072);
nand U14285 (N_14285,N_14038,N_14157);
nor U14286 (N_14286,N_14223,N_14063);
nor U14287 (N_14287,N_14001,N_14189);
nor U14288 (N_14288,N_14084,N_14054);
or U14289 (N_14289,N_14239,N_14212);
nor U14290 (N_14290,N_14243,N_14168);
xor U14291 (N_14291,N_14073,N_14036);
nand U14292 (N_14292,N_14020,N_14217);
nor U14293 (N_14293,N_14152,N_14059);
or U14294 (N_14294,N_14181,N_14083);
or U14295 (N_14295,N_14012,N_14202);
and U14296 (N_14296,N_14077,N_14196);
nor U14297 (N_14297,N_14025,N_14095);
nor U14298 (N_14298,N_14174,N_14034);
nand U14299 (N_14299,N_14209,N_14090);
nor U14300 (N_14300,N_14194,N_14086);
and U14301 (N_14301,N_14233,N_14232);
and U14302 (N_14302,N_14053,N_14171);
and U14303 (N_14303,N_14173,N_14237);
and U14304 (N_14304,N_14121,N_14046);
and U14305 (N_14305,N_14018,N_14105);
or U14306 (N_14306,N_14045,N_14161);
xor U14307 (N_14307,N_14029,N_14153);
or U14308 (N_14308,N_14204,N_14116);
or U14309 (N_14309,N_14099,N_14130);
xor U14310 (N_14310,N_14110,N_14024);
or U14311 (N_14311,N_14205,N_14107);
nand U14312 (N_14312,N_14208,N_14028);
xnor U14313 (N_14313,N_14114,N_14178);
nor U14314 (N_14314,N_14089,N_14150);
xnor U14315 (N_14315,N_14127,N_14057);
nand U14316 (N_14316,N_14221,N_14117);
nand U14317 (N_14317,N_14186,N_14241);
or U14318 (N_14318,N_14210,N_14131);
nand U14319 (N_14319,N_14078,N_14016);
nor U14320 (N_14320,N_14154,N_14141);
nor U14321 (N_14321,N_14055,N_14170);
or U14322 (N_14322,N_14010,N_14179);
nor U14323 (N_14323,N_14068,N_14229);
nand U14324 (N_14324,N_14133,N_14071);
or U14325 (N_14325,N_14234,N_14070);
or U14326 (N_14326,N_14187,N_14242);
or U14327 (N_14327,N_14040,N_14225);
nor U14328 (N_14328,N_14098,N_14037);
xnor U14329 (N_14329,N_14088,N_14004);
nor U14330 (N_14330,N_14220,N_14148);
and U14331 (N_14331,N_14014,N_14244);
nand U14332 (N_14332,N_14175,N_14066);
nor U14333 (N_14333,N_14094,N_14201);
or U14334 (N_14334,N_14235,N_14009);
nand U14335 (N_14335,N_14122,N_14017);
and U14336 (N_14336,N_14198,N_14166);
nor U14337 (N_14337,N_14169,N_14218);
or U14338 (N_14338,N_14003,N_14249);
nor U14339 (N_14339,N_14134,N_14191);
xnor U14340 (N_14340,N_14042,N_14214);
nor U14341 (N_14341,N_14062,N_14147);
xnor U14342 (N_14342,N_14006,N_14013);
or U14343 (N_14343,N_14079,N_14052);
or U14344 (N_14344,N_14111,N_14113);
xor U14345 (N_14345,N_14184,N_14135);
nor U14346 (N_14346,N_14224,N_14112);
and U14347 (N_14347,N_14128,N_14081);
nand U14348 (N_14348,N_14226,N_14087);
nor U14349 (N_14349,N_14167,N_14069);
and U14350 (N_14350,N_14033,N_14200);
and U14351 (N_14351,N_14082,N_14182);
and U14352 (N_14352,N_14236,N_14151);
nor U14353 (N_14353,N_14158,N_14093);
nor U14354 (N_14354,N_14144,N_14023);
xor U14355 (N_14355,N_14238,N_14164);
and U14356 (N_14356,N_14015,N_14125);
nor U14357 (N_14357,N_14101,N_14075);
xor U14358 (N_14358,N_14176,N_14240);
nor U14359 (N_14359,N_14145,N_14005);
xor U14360 (N_14360,N_14183,N_14074);
and U14361 (N_14361,N_14140,N_14207);
xnor U14362 (N_14362,N_14138,N_14021);
nand U14363 (N_14363,N_14104,N_14044);
or U14364 (N_14364,N_14065,N_14129);
or U14365 (N_14365,N_14246,N_14245);
nand U14366 (N_14366,N_14026,N_14061);
nor U14367 (N_14367,N_14050,N_14155);
nand U14368 (N_14368,N_14163,N_14215);
xor U14369 (N_14369,N_14002,N_14211);
and U14370 (N_14370,N_14030,N_14115);
nor U14371 (N_14371,N_14247,N_14197);
or U14372 (N_14372,N_14159,N_14213);
xor U14373 (N_14373,N_14142,N_14123);
xnor U14374 (N_14374,N_14106,N_14100);
xor U14375 (N_14375,N_14101,N_14176);
xor U14376 (N_14376,N_14032,N_14213);
xor U14377 (N_14377,N_14180,N_14224);
and U14378 (N_14378,N_14050,N_14214);
xor U14379 (N_14379,N_14201,N_14041);
nor U14380 (N_14380,N_14077,N_14205);
nor U14381 (N_14381,N_14085,N_14023);
and U14382 (N_14382,N_14203,N_14153);
and U14383 (N_14383,N_14105,N_14001);
or U14384 (N_14384,N_14019,N_14148);
nand U14385 (N_14385,N_14027,N_14226);
nand U14386 (N_14386,N_14085,N_14145);
nor U14387 (N_14387,N_14160,N_14117);
xor U14388 (N_14388,N_14179,N_14083);
nor U14389 (N_14389,N_14159,N_14218);
or U14390 (N_14390,N_14225,N_14084);
nor U14391 (N_14391,N_14118,N_14059);
and U14392 (N_14392,N_14241,N_14134);
nor U14393 (N_14393,N_14107,N_14110);
nor U14394 (N_14394,N_14048,N_14217);
xnor U14395 (N_14395,N_14103,N_14082);
nor U14396 (N_14396,N_14000,N_14206);
xor U14397 (N_14397,N_14072,N_14248);
and U14398 (N_14398,N_14076,N_14141);
nand U14399 (N_14399,N_14206,N_14246);
nor U14400 (N_14400,N_14120,N_14227);
nand U14401 (N_14401,N_14005,N_14169);
and U14402 (N_14402,N_14057,N_14004);
nor U14403 (N_14403,N_14090,N_14068);
or U14404 (N_14404,N_14146,N_14044);
nor U14405 (N_14405,N_14104,N_14114);
nand U14406 (N_14406,N_14007,N_14078);
nand U14407 (N_14407,N_14204,N_14183);
xor U14408 (N_14408,N_14070,N_14068);
nand U14409 (N_14409,N_14000,N_14114);
nand U14410 (N_14410,N_14023,N_14160);
or U14411 (N_14411,N_14218,N_14242);
nand U14412 (N_14412,N_14058,N_14131);
and U14413 (N_14413,N_14095,N_14003);
or U14414 (N_14414,N_14147,N_14037);
xnor U14415 (N_14415,N_14169,N_14113);
nor U14416 (N_14416,N_14214,N_14084);
and U14417 (N_14417,N_14041,N_14197);
and U14418 (N_14418,N_14004,N_14013);
and U14419 (N_14419,N_14221,N_14125);
xor U14420 (N_14420,N_14206,N_14156);
xnor U14421 (N_14421,N_14228,N_14087);
xnor U14422 (N_14422,N_14113,N_14187);
nor U14423 (N_14423,N_14242,N_14078);
nand U14424 (N_14424,N_14133,N_14018);
or U14425 (N_14425,N_14137,N_14162);
nand U14426 (N_14426,N_14222,N_14085);
or U14427 (N_14427,N_14150,N_14223);
and U14428 (N_14428,N_14170,N_14128);
and U14429 (N_14429,N_14241,N_14001);
and U14430 (N_14430,N_14231,N_14085);
nand U14431 (N_14431,N_14214,N_14070);
or U14432 (N_14432,N_14243,N_14217);
and U14433 (N_14433,N_14048,N_14185);
or U14434 (N_14434,N_14109,N_14047);
nand U14435 (N_14435,N_14237,N_14008);
xor U14436 (N_14436,N_14142,N_14063);
or U14437 (N_14437,N_14214,N_14213);
nor U14438 (N_14438,N_14012,N_14127);
nor U14439 (N_14439,N_14016,N_14224);
and U14440 (N_14440,N_14217,N_14249);
nor U14441 (N_14441,N_14112,N_14241);
nor U14442 (N_14442,N_14227,N_14182);
nand U14443 (N_14443,N_14125,N_14042);
and U14444 (N_14444,N_14162,N_14170);
xnor U14445 (N_14445,N_14176,N_14132);
nand U14446 (N_14446,N_14012,N_14244);
nand U14447 (N_14447,N_14231,N_14019);
or U14448 (N_14448,N_14097,N_14051);
nand U14449 (N_14449,N_14231,N_14168);
xnor U14450 (N_14450,N_14075,N_14185);
nand U14451 (N_14451,N_14071,N_14178);
or U14452 (N_14452,N_14084,N_14176);
nor U14453 (N_14453,N_14244,N_14003);
nor U14454 (N_14454,N_14213,N_14094);
xnor U14455 (N_14455,N_14162,N_14038);
and U14456 (N_14456,N_14104,N_14233);
nor U14457 (N_14457,N_14199,N_14062);
xor U14458 (N_14458,N_14005,N_14086);
nor U14459 (N_14459,N_14202,N_14098);
xnor U14460 (N_14460,N_14049,N_14039);
nand U14461 (N_14461,N_14141,N_14020);
nor U14462 (N_14462,N_14216,N_14171);
nand U14463 (N_14463,N_14043,N_14121);
xnor U14464 (N_14464,N_14054,N_14108);
or U14465 (N_14465,N_14106,N_14024);
nor U14466 (N_14466,N_14063,N_14055);
xnor U14467 (N_14467,N_14106,N_14095);
or U14468 (N_14468,N_14189,N_14200);
and U14469 (N_14469,N_14112,N_14011);
and U14470 (N_14470,N_14004,N_14066);
nand U14471 (N_14471,N_14098,N_14058);
nor U14472 (N_14472,N_14231,N_14209);
nand U14473 (N_14473,N_14243,N_14157);
and U14474 (N_14474,N_14037,N_14052);
or U14475 (N_14475,N_14109,N_14005);
or U14476 (N_14476,N_14049,N_14208);
xor U14477 (N_14477,N_14095,N_14040);
nand U14478 (N_14478,N_14163,N_14114);
xor U14479 (N_14479,N_14038,N_14160);
nand U14480 (N_14480,N_14110,N_14172);
and U14481 (N_14481,N_14125,N_14177);
xor U14482 (N_14482,N_14229,N_14066);
or U14483 (N_14483,N_14083,N_14240);
or U14484 (N_14484,N_14143,N_14155);
or U14485 (N_14485,N_14078,N_14153);
nand U14486 (N_14486,N_14093,N_14126);
or U14487 (N_14487,N_14194,N_14075);
nor U14488 (N_14488,N_14121,N_14009);
or U14489 (N_14489,N_14111,N_14107);
nor U14490 (N_14490,N_14054,N_14235);
or U14491 (N_14491,N_14242,N_14175);
nor U14492 (N_14492,N_14119,N_14197);
nand U14493 (N_14493,N_14099,N_14194);
nor U14494 (N_14494,N_14244,N_14055);
nor U14495 (N_14495,N_14140,N_14114);
and U14496 (N_14496,N_14068,N_14247);
nor U14497 (N_14497,N_14208,N_14218);
nand U14498 (N_14498,N_14145,N_14097);
or U14499 (N_14499,N_14192,N_14102);
and U14500 (N_14500,N_14380,N_14400);
nand U14501 (N_14501,N_14449,N_14396);
xnor U14502 (N_14502,N_14284,N_14410);
and U14503 (N_14503,N_14277,N_14432);
nor U14504 (N_14504,N_14407,N_14493);
nor U14505 (N_14505,N_14348,N_14383);
xnor U14506 (N_14506,N_14460,N_14358);
nor U14507 (N_14507,N_14393,N_14262);
and U14508 (N_14508,N_14336,N_14471);
xor U14509 (N_14509,N_14479,N_14427);
or U14510 (N_14510,N_14436,N_14435);
xor U14511 (N_14511,N_14331,N_14496);
nor U14512 (N_14512,N_14487,N_14329);
xor U14513 (N_14513,N_14312,N_14325);
or U14514 (N_14514,N_14405,N_14353);
nand U14515 (N_14515,N_14297,N_14430);
nor U14516 (N_14516,N_14468,N_14453);
or U14517 (N_14517,N_14317,N_14374);
or U14518 (N_14518,N_14328,N_14365);
or U14519 (N_14519,N_14316,N_14324);
and U14520 (N_14520,N_14499,N_14344);
nand U14521 (N_14521,N_14268,N_14433);
nor U14522 (N_14522,N_14442,N_14295);
nor U14523 (N_14523,N_14422,N_14477);
xnor U14524 (N_14524,N_14327,N_14434);
and U14525 (N_14525,N_14409,N_14254);
nor U14526 (N_14526,N_14481,N_14415);
xor U14527 (N_14527,N_14386,N_14253);
xnor U14528 (N_14528,N_14315,N_14347);
or U14529 (N_14529,N_14462,N_14360);
nor U14530 (N_14530,N_14337,N_14369);
or U14531 (N_14531,N_14446,N_14343);
nor U14532 (N_14532,N_14346,N_14425);
nand U14533 (N_14533,N_14388,N_14318);
and U14534 (N_14534,N_14431,N_14299);
nor U14535 (N_14535,N_14291,N_14488);
xor U14536 (N_14536,N_14308,N_14426);
xor U14537 (N_14537,N_14489,N_14390);
or U14538 (N_14538,N_14322,N_14279);
xnor U14539 (N_14539,N_14439,N_14490);
and U14540 (N_14540,N_14314,N_14445);
nand U14541 (N_14541,N_14258,N_14391);
nand U14542 (N_14542,N_14320,N_14421);
nand U14543 (N_14543,N_14271,N_14259);
nor U14544 (N_14544,N_14486,N_14355);
xnor U14545 (N_14545,N_14286,N_14470);
or U14546 (N_14546,N_14257,N_14349);
nand U14547 (N_14547,N_14250,N_14474);
xor U14548 (N_14548,N_14376,N_14363);
or U14549 (N_14549,N_14492,N_14283);
and U14550 (N_14550,N_14332,N_14361);
xor U14551 (N_14551,N_14303,N_14455);
and U14552 (N_14552,N_14264,N_14472);
and U14553 (N_14553,N_14354,N_14389);
nand U14554 (N_14554,N_14367,N_14408);
nand U14555 (N_14555,N_14384,N_14302);
and U14556 (N_14556,N_14368,N_14273);
nand U14557 (N_14557,N_14265,N_14281);
nand U14558 (N_14558,N_14404,N_14377);
nor U14559 (N_14559,N_14413,N_14483);
and U14560 (N_14560,N_14330,N_14473);
or U14561 (N_14561,N_14313,N_14270);
nand U14562 (N_14562,N_14424,N_14382);
nor U14563 (N_14563,N_14357,N_14263);
xnor U14564 (N_14564,N_14420,N_14366);
or U14565 (N_14565,N_14401,N_14484);
nor U14566 (N_14566,N_14406,N_14371);
xor U14567 (N_14567,N_14423,N_14466);
or U14568 (N_14568,N_14298,N_14285);
and U14569 (N_14569,N_14387,N_14397);
and U14570 (N_14570,N_14480,N_14288);
xor U14571 (N_14571,N_14447,N_14260);
xnor U14572 (N_14572,N_14494,N_14469);
and U14573 (N_14573,N_14342,N_14463);
nor U14574 (N_14574,N_14441,N_14456);
nand U14575 (N_14575,N_14414,N_14282);
and U14576 (N_14576,N_14351,N_14292);
xor U14577 (N_14577,N_14311,N_14381);
xor U14578 (N_14578,N_14465,N_14399);
and U14579 (N_14579,N_14498,N_14495);
xor U14580 (N_14580,N_14373,N_14319);
nand U14581 (N_14581,N_14385,N_14375);
and U14582 (N_14582,N_14443,N_14461);
nand U14583 (N_14583,N_14321,N_14294);
nor U14584 (N_14584,N_14429,N_14491);
nand U14585 (N_14585,N_14450,N_14339);
nand U14586 (N_14586,N_14398,N_14255);
or U14587 (N_14587,N_14497,N_14252);
xnor U14588 (N_14588,N_14458,N_14372);
xor U14589 (N_14589,N_14266,N_14394);
nor U14590 (N_14590,N_14392,N_14280);
nor U14591 (N_14591,N_14323,N_14459);
and U14592 (N_14592,N_14478,N_14440);
or U14593 (N_14593,N_14411,N_14300);
and U14594 (N_14594,N_14261,N_14310);
nor U14595 (N_14595,N_14437,N_14309);
nor U14596 (N_14596,N_14476,N_14301);
nor U14597 (N_14597,N_14448,N_14272);
nand U14598 (N_14598,N_14287,N_14326);
nand U14599 (N_14599,N_14402,N_14289);
or U14600 (N_14600,N_14403,N_14370);
nor U14601 (N_14601,N_14444,N_14464);
nand U14602 (N_14602,N_14416,N_14306);
nand U14603 (N_14603,N_14338,N_14362);
nor U14604 (N_14604,N_14485,N_14333);
nand U14605 (N_14605,N_14275,N_14352);
or U14606 (N_14606,N_14419,N_14256);
nand U14607 (N_14607,N_14451,N_14359);
or U14608 (N_14608,N_14378,N_14296);
nand U14609 (N_14609,N_14340,N_14293);
and U14610 (N_14610,N_14364,N_14290);
xor U14611 (N_14611,N_14304,N_14418);
nand U14612 (N_14612,N_14274,N_14276);
or U14613 (N_14613,N_14452,N_14356);
and U14614 (N_14614,N_14305,N_14395);
nor U14615 (N_14615,N_14428,N_14345);
and U14616 (N_14616,N_14267,N_14457);
nand U14617 (N_14617,N_14417,N_14454);
or U14618 (N_14618,N_14307,N_14251);
and U14619 (N_14619,N_14475,N_14278);
xnor U14620 (N_14620,N_14467,N_14350);
and U14621 (N_14621,N_14341,N_14412);
nor U14622 (N_14622,N_14438,N_14482);
xnor U14623 (N_14623,N_14379,N_14269);
and U14624 (N_14624,N_14335,N_14334);
nor U14625 (N_14625,N_14462,N_14304);
or U14626 (N_14626,N_14348,N_14357);
xor U14627 (N_14627,N_14386,N_14414);
or U14628 (N_14628,N_14295,N_14260);
nor U14629 (N_14629,N_14425,N_14331);
nand U14630 (N_14630,N_14398,N_14371);
or U14631 (N_14631,N_14427,N_14262);
and U14632 (N_14632,N_14499,N_14353);
nand U14633 (N_14633,N_14494,N_14414);
nor U14634 (N_14634,N_14306,N_14263);
or U14635 (N_14635,N_14353,N_14374);
or U14636 (N_14636,N_14420,N_14327);
nor U14637 (N_14637,N_14323,N_14384);
nor U14638 (N_14638,N_14386,N_14353);
nand U14639 (N_14639,N_14328,N_14498);
or U14640 (N_14640,N_14250,N_14315);
and U14641 (N_14641,N_14433,N_14392);
nand U14642 (N_14642,N_14374,N_14310);
or U14643 (N_14643,N_14285,N_14427);
xnor U14644 (N_14644,N_14493,N_14455);
nand U14645 (N_14645,N_14440,N_14468);
or U14646 (N_14646,N_14478,N_14352);
xor U14647 (N_14647,N_14408,N_14256);
and U14648 (N_14648,N_14295,N_14273);
or U14649 (N_14649,N_14371,N_14348);
and U14650 (N_14650,N_14380,N_14481);
nand U14651 (N_14651,N_14490,N_14423);
nand U14652 (N_14652,N_14395,N_14297);
nor U14653 (N_14653,N_14366,N_14267);
nand U14654 (N_14654,N_14318,N_14477);
xnor U14655 (N_14655,N_14395,N_14398);
or U14656 (N_14656,N_14449,N_14399);
xor U14657 (N_14657,N_14387,N_14300);
or U14658 (N_14658,N_14373,N_14449);
xor U14659 (N_14659,N_14358,N_14483);
xnor U14660 (N_14660,N_14478,N_14433);
nand U14661 (N_14661,N_14304,N_14372);
and U14662 (N_14662,N_14407,N_14291);
nand U14663 (N_14663,N_14275,N_14378);
and U14664 (N_14664,N_14491,N_14401);
and U14665 (N_14665,N_14435,N_14315);
or U14666 (N_14666,N_14321,N_14391);
xnor U14667 (N_14667,N_14441,N_14258);
and U14668 (N_14668,N_14357,N_14338);
nand U14669 (N_14669,N_14381,N_14279);
nand U14670 (N_14670,N_14368,N_14270);
nor U14671 (N_14671,N_14415,N_14268);
or U14672 (N_14672,N_14274,N_14445);
xor U14673 (N_14673,N_14420,N_14340);
nor U14674 (N_14674,N_14445,N_14385);
nor U14675 (N_14675,N_14266,N_14351);
nor U14676 (N_14676,N_14456,N_14397);
nand U14677 (N_14677,N_14452,N_14385);
xor U14678 (N_14678,N_14368,N_14337);
xnor U14679 (N_14679,N_14368,N_14369);
xnor U14680 (N_14680,N_14349,N_14273);
and U14681 (N_14681,N_14387,N_14456);
or U14682 (N_14682,N_14397,N_14268);
nor U14683 (N_14683,N_14261,N_14422);
or U14684 (N_14684,N_14345,N_14386);
and U14685 (N_14685,N_14324,N_14350);
nand U14686 (N_14686,N_14368,N_14307);
or U14687 (N_14687,N_14473,N_14436);
nand U14688 (N_14688,N_14262,N_14307);
xor U14689 (N_14689,N_14312,N_14432);
nor U14690 (N_14690,N_14409,N_14441);
nor U14691 (N_14691,N_14371,N_14302);
nor U14692 (N_14692,N_14485,N_14398);
nor U14693 (N_14693,N_14263,N_14476);
or U14694 (N_14694,N_14480,N_14280);
nand U14695 (N_14695,N_14264,N_14418);
xnor U14696 (N_14696,N_14497,N_14381);
xor U14697 (N_14697,N_14349,N_14434);
nand U14698 (N_14698,N_14309,N_14479);
and U14699 (N_14699,N_14283,N_14388);
and U14700 (N_14700,N_14292,N_14429);
xor U14701 (N_14701,N_14375,N_14471);
and U14702 (N_14702,N_14274,N_14441);
nor U14703 (N_14703,N_14481,N_14441);
or U14704 (N_14704,N_14421,N_14450);
nor U14705 (N_14705,N_14484,N_14464);
and U14706 (N_14706,N_14385,N_14439);
xor U14707 (N_14707,N_14258,N_14378);
xor U14708 (N_14708,N_14375,N_14355);
and U14709 (N_14709,N_14493,N_14342);
nand U14710 (N_14710,N_14357,N_14268);
and U14711 (N_14711,N_14280,N_14472);
nand U14712 (N_14712,N_14434,N_14260);
xnor U14713 (N_14713,N_14250,N_14422);
xor U14714 (N_14714,N_14390,N_14404);
or U14715 (N_14715,N_14445,N_14434);
and U14716 (N_14716,N_14318,N_14327);
nand U14717 (N_14717,N_14254,N_14344);
xor U14718 (N_14718,N_14294,N_14302);
or U14719 (N_14719,N_14408,N_14386);
and U14720 (N_14720,N_14465,N_14312);
and U14721 (N_14721,N_14463,N_14320);
or U14722 (N_14722,N_14256,N_14372);
nor U14723 (N_14723,N_14434,N_14330);
or U14724 (N_14724,N_14410,N_14369);
nand U14725 (N_14725,N_14391,N_14426);
nand U14726 (N_14726,N_14390,N_14396);
and U14727 (N_14727,N_14491,N_14371);
xnor U14728 (N_14728,N_14251,N_14373);
and U14729 (N_14729,N_14327,N_14367);
xor U14730 (N_14730,N_14320,N_14458);
nor U14731 (N_14731,N_14364,N_14409);
and U14732 (N_14732,N_14476,N_14490);
nand U14733 (N_14733,N_14391,N_14432);
xnor U14734 (N_14734,N_14416,N_14483);
or U14735 (N_14735,N_14331,N_14453);
or U14736 (N_14736,N_14475,N_14371);
xor U14737 (N_14737,N_14383,N_14274);
nand U14738 (N_14738,N_14406,N_14397);
xnor U14739 (N_14739,N_14263,N_14458);
xor U14740 (N_14740,N_14419,N_14306);
xor U14741 (N_14741,N_14306,N_14319);
nand U14742 (N_14742,N_14440,N_14377);
nand U14743 (N_14743,N_14440,N_14278);
nor U14744 (N_14744,N_14366,N_14297);
nor U14745 (N_14745,N_14447,N_14437);
nand U14746 (N_14746,N_14260,N_14392);
nor U14747 (N_14747,N_14352,N_14355);
nand U14748 (N_14748,N_14420,N_14407);
and U14749 (N_14749,N_14291,N_14357);
and U14750 (N_14750,N_14721,N_14705);
or U14751 (N_14751,N_14609,N_14619);
xor U14752 (N_14752,N_14706,N_14654);
nand U14753 (N_14753,N_14579,N_14633);
nor U14754 (N_14754,N_14527,N_14732);
xnor U14755 (N_14755,N_14691,N_14558);
xor U14756 (N_14756,N_14522,N_14617);
xnor U14757 (N_14757,N_14516,N_14572);
nor U14758 (N_14758,N_14550,N_14581);
xnor U14759 (N_14759,N_14710,N_14690);
nor U14760 (N_14760,N_14600,N_14675);
xor U14761 (N_14761,N_14593,N_14728);
xor U14762 (N_14762,N_14526,N_14612);
nand U14763 (N_14763,N_14692,N_14589);
nor U14764 (N_14764,N_14741,N_14616);
nand U14765 (N_14765,N_14714,N_14547);
xor U14766 (N_14766,N_14746,N_14711);
and U14767 (N_14767,N_14587,N_14537);
and U14768 (N_14768,N_14667,N_14519);
xnor U14769 (N_14769,N_14716,N_14606);
xnor U14770 (N_14770,N_14583,N_14686);
xnor U14771 (N_14771,N_14742,N_14730);
and U14772 (N_14772,N_14666,N_14590);
nand U14773 (N_14773,N_14515,N_14552);
xor U14774 (N_14774,N_14739,N_14545);
xor U14775 (N_14775,N_14698,N_14709);
nor U14776 (N_14776,N_14726,N_14635);
nor U14777 (N_14777,N_14649,N_14659);
nand U14778 (N_14778,N_14614,N_14615);
and U14779 (N_14779,N_14544,N_14529);
nor U14780 (N_14780,N_14669,N_14502);
nand U14781 (N_14781,N_14682,N_14580);
nand U14782 (N_14782,N_14604,N_14717);
nor U14783 (N_14783,N_14508,N_14627);
nor U14784 (N_14784,N_14573,N_14598);
or U14785 (N_14785,N_14655,N_14531);
xor U14786 (N_14786,N_14503,N_14673);
and U14787 (N_14787,N_14591,N_14628);
or U14788 (N_14788,N_14511,N_14533);
or U14789 (N_14789,N_14510,N_14651);
or U14790 (N_14790,N_14555,N_14724);
xor U14791 (N_14791,N_14566,N_14672);
and U14792 (N_14792,N_14622,N_14592);
nor U14793 (N_14793,N_14677,N_14722);
or U14794 (N_14794,N_14629,N_14549);
and U14795 (N_14795,N_14582,N_14638);
nor U14796 (N_14796,N_14689,N_14605);
or U14797 (N_14797,N_14625,N_14568);
or U14798 (N_14798,N_14500,N_14599);
nand U14799 (N_14799,N_14607,N_14743);
and U14800 (N_14800,N_14674,N_14624);
or U14801 (N_14801,N_14576,N_14696);
or U14802 (N_14802,N_14652,N_14695);
or U14803 (N_14803,N_14548,N_14744);
xnor U14804 (N_14804,N_14685,N_14749);
or U14805 (N_14805,N_14643,N_14661);
nand U14806 (N_14806,N_14697,N_14687);
or U14807 (N_14807,N_14729,N_14525);
and U14808 (N_14808,N_14642,N_14506);
or U14809 (N_14809,N_14658,N_14540);
xor U14810 (N_14810,N_14584,N_14534);
nand U14811 (N_14811,N_14588,N_14532);
nand U14812 (N_14812,N_14740,N_14610);
nand U14813 (N_14813,N_14559,N_14562);
and U14814 (N_14814,N_14707,N_14578);
and U14815 (N_14815,N_14539,N_14644);
nor U14816 (N_14816,N_14524,N_14738);
nand U14817 (N_14817,N_14543,N_14631);
nor U14818 (N_14818,N_14703,N_14664);
nor U14819 (N_14819,N_14538,N_14603);
nor U14820 (N_14820,N_14520,N_14720);
nor U14821 (N_14821,N_14597,N_14679);
nand U14822 (N_14822,N_14554,N_14586);
xor U14823 (N_14823,N_14641,N_14648);
xor U14824 (N_14824,N_14736,N_14733);
xor U14825 (N_14825,N_14670,N_14735);
xor U14826 (N_14826,N_14645,N_14713);
and U14827 (N_14827,N_14715,N_14700);
nand U14828 (N_14828,N_14683,N_14618);
xor U14829 (N_14829,N_14608,N_14639);
xnor U14830 (N_14830,N_14694,N_14535);
xor U14831 (N_14831,N_14596,N_14708);
or U14832 (N_14832,N_14509,N_14719);
nor U14833 (N_14833,N_14681,N_14517);
and U14834 (N_14834,N_14632,N_14561);
nor U14835 (N_14835,N_14699,N_14727);
nand U14836 (N_14836,N_14536,N_14613);
nor U14837 (N_14837,N_14636,N_14571);
xnor U14838 (N_14838,N_14560,N_14553);
xnor U14839 (N_14839,N_14671,N_14542);
nand U14840 (N_14840,N_14702,N_14680);
nor U14841 (N_14841,N_14594,N_14676);
and U14842 (N_14842,N_14712,N_14701);
xor U14843 (N_14843,N_14541,N_14595);
and U14844 (N_14844,N_14505,N_14684);
nor U14845 (N_14845,N_14565,N_14564);
or U14846 (N_14846,N_14637,N_14567);
and U14847 (N_14847,N_14512,N_14725);
and U14848 (N_14848,N_14748,N_14662);
nor U14849 (N_14849,N_14747,N_14507);
nor U14850 (N_14850,N_14530,N_14620);
nor U14851 (N_14851,N_14563,N_14546);
nor U14852 (N_14852,N_14634,N_14660);
and U14853 (N_14853,N_14718,N_14621);
nor U14854 (N_14854,N_14657,N_14663);
nor U14855 (N_14855,N_14504,N_14668);
and U14856 (N_14856,N_14650,N_14678);
nor U14857 (N_14857,N_14745,N_14646);
and U14858 (N_14858,N_14656,N_14570);
nor U14859 (N_14859,N_14665,N_14623);
nand U14860 (N_14860,N_14574,N_14513);
and U14861 (N_14861,N_14647,N_14640);
and U14862 (N_14862,N_14556,N_14577);
nand U14863 (N_14863,N_14523,N_14585);
and U14864 (N_14864,N_14575,N_14602);
nor U14865 (N_14865,N_14551,N_14501);
or U14866 (N_14866,N_14704,N_14731);
nand U14867 (N_14867,N_14557,N_14601);
nor U14868 (N_14868,N_14569,N_14688);
nor U14869 (N_14869,N_14734,N_14693);
or U14870 (N_14870,N_14723,N_14528);
and U14871 (N_14871,N_14521,N_14737);
xor U14872 (N_14872,N_14518,N_14653);
nand U14873 (N_14873,N_14630,N_14514);
nor U14874 (N_14874,N_14626,N_14611);
nand U14875 (N_14875,N_14517,N_14732);
or U14876 (N_14876,N_14666,N_14565);
or U14877 (N_14877,N_14533,N_14728);
nand U14878 (N_14878,N_14666,N_14513);
xnor U14879 (N_14879,N_14591,N_14597);
xnor U14880 (N_14880,N_14687,N_14641);
or U14881 (N_14881,N_14630,N_14638);
nand U14882 (N_14882,N_14731,N_14736);
and U14883 (N_14883,N_14517,N_14510);
nand U14884 (N_14884,N_14718,N_14648);
nand U14885 (N_14885,N_14508,N_14736);
xor U14886 (N_14886,N_14636,N_14643);
nor U14887 (N_14887,N_14563,N_14625);
xnor U14888 (N_14888,N_14609,N_14691);
nand U14889 (N_14889,N_14714,N_14713);
nand U14890 (N_14890,N_14717,N_14531);
nand U14891 (N_14891,N_14563,N_14540);
nor U14892 (N_14892,N_14736,N_14744);
and U14893 (N_14893,N_14634,N_14723);
and U14894 (N_14894,N_14667,N_14609);
xnor U14895 (N_14895,N_14587,N_14717);
and U14896 (N_14896,N_14674,N_14584);
or U14897 (N_14897,N_14610,N_14587);
nand U14898 (N_14898,N_14707,N_14712);
and U14899 (N_14899,N_14633,N_14640);
nor U14900 (N_14900,N_14606,N_14732);
nor U14901 (N_14901,N_14545,N_14616);
nand U14902 (N_14902,N_14637,N_14669);
xor U14903 (N_14903,N_14537,N_14557);
and U14904 (N_14904,N_14628,N_14529);
nand U14905 (N_14905,N_14573,N_14712);
and U14906 (N_14906,N_14659,N_14697);
and U14907 (N_14907,N_14724,N_14731);
nand U14908 (N_14908,N_14575,N_14703);
xnor U14909 (N_14909,N_14741,N_14569);
nor U14910 (N_14910,N_14634,N_14717);
and U14911 (N_14911,N_14515,N_14517);
and U14912 (N_14912,N_14695,N_14610);
and U14913 (N_14913,N_14611,N_14731);
xor U14914 (N_14914,N_14549,N_14632);
nor U14915 (N_14915,N_14650,N_14625);
xor U14916 (N_14916,N_14505,N_14708);
nand U14917 (N_14917,N_14597,N_14705);
xnor U14918 (N_14918,N_14609,N_14611);
and U14919 (N_14919,N_14561,N_14702);
xor U14920 (N_14920,N_14580,N_14631);
or U14921 (N_14921,N_14680,N_14553);
nand U14922 (N_14922,N_14669,N_14517);
or U14923 (N_14923,N_14702,N_14645);
and U14924 (N_14924,N_14741,N_14684);
nor U14925 (N_14925,N_14514,N_14648);
nor U14926 (N_14926,N_14739,N_14622);
and U14927 (N_14927,N_14548,N_14735);
nand U14928 (N_14928,N_14604,N_14715);
nor U14929 (N_14929,N_14715,N_14568);
or U14930 (N_14930,N_14612,N_14644);
or U14931 (N_14931,N_14670,N_14678);
nand U14932 (N_14932,N_14541,N_14589);
nand U14933 (N_14933,N_14557,N_14737);
nor U14934 (N_14934,N_14539,N_14686);
xor U14935 (N_14935,N_14682,N_14545);
xor U14936 (N_14936,N_14695,N_14682);
nor U14937 (N_14937,N_14513,N_14660);
nand U14938 (N_14938,N_14547,N_14685);
nor U14939 (N_14939,N_14631,N_14740);
nor U14940 (N_14940,N_14502,N_14615);
xnor U14941 (N_14941,N_14650,N_14588);
nand U14942 (N_14942,N_14694,N_14516);
or U14943 (N_14943,N_14547,N_14528);
or U14944 (N_14944,N_14654,N_14746);
or U14945 (N_14945,N_14728,N_14621);
nand U14946 (N_14946,N_14637,N_14645);
and U14947 (N_14947,N_14686,N_14544);
nand U14948 (N_14948,N_14611,N_14711);
and U14949 (N_14949,N_14544,N_14534);
or U14950 (N_14950,N_14539,N_14729);
nand U14951 (N_14951,N_14742,N_14655);
nor U14952 (N_14952,N_14738,N_14540);
nand U14953 (N_14953,N_14512,N_14534);
nand U14954 (N_14954,N_14657,N_14664);
nand U14955 (N_14955,N_14671,N_14567);
nand U14956 (N_14956,N_14739,N_14720);
xnor U14957 (N_14957,N_14746,N_14579);
nor U14958 (N_14958,N_14702,N_14719);
nand U14959 (N_14959,N_14740,N_14647);
nand U14960 (N_14960,N_14682,N_14746);
or U14961 (N_14961,N_14740,N_14618);
or U14962 (N_14962,N_14643,N_14656);
xor U14963 (N_14963,N_14605,N_14673);
or U14964 (N_14964,N_14635,N_14542);
nor U14965 (N_14965,N_14557,N_14590);
xor U14966 (N_14966,N_14572,N_14734);
nor U14967 (N_14967,N_14599,N_14580);
xor U14968 (N_14968,N_14584,N_14549);
xor U14969 (N_14969,N_14588,N_14735);
nand U14970 (N_14970,N_14621,N_14599);
nand U14971 (N_14971,N_14583,N_14704);
or U14972 (N_14972,N_14562,N_14620);
nand U14973 (N_14973,N_14556,N_14530);
xor U14974 (N_14974,N_14612,N_14550);
xor U14975 (N_14975,N_14550,N_14566);
and U14976 (N_14976,N_14600,N_14715);
xor U14977 (N_14977,N_14546,N_14674);
and U14978 (N_14978,N_14545,N_14572);
and U14979 (N_14979,N_14626,N_14567);
or U14980 (N_14980,N_14562,N_14725);
or U14981 (N_14981,N_14563,N_14705);
or U14982 (N_14982,N_14718,N_14599);
xor U14983 (N_14983,N_14590,N_14540);
xor U14984 (N_14984,N_14508,N_14539);
and U14985 (N_14985,N_14516,N_14546);
xnor U14986 (N_14986,N_14551,N_14599);
xnor U14987 (N_14987,N_14632,N_14515);
nor U14988 (N_14988,N_14739,N_14511);
xor U14989 (N_14989,N_14734,N_14687);
or U14990 (N_14990,N_14673,N_14734);
or U14991 (N_14991,N_14618,N_14593);
or U14992 (N_14992,N_14669,N_14521);
xor U14993 (N_14993,N_14502,N_14718);
nor U14994 (N_14994,N_14610,N_14516);
nor U14995 (N_14995,N_14702,N_14638);
or U14996 (N_14996,N_14598,N_14682);
nand U14997 (N_14997,N_14522,N_14637);
or U14998 (N_14998,N_14608,N_14738);
xor U14999 (N_14999,N_14743,N_14630);
and U15000 (N_15000,N_14994,N_14759);
xnor U15001 (N_15001,N_14773,N_14959);
nand U15002 (N_15002,N_14795,N_14853);
and U15003 (N_15003,N_14999,N_14785);
xnor U15004 (N_15004,N_14920,N_14791);
xnor U15005 (N_15005,N_14937,N_14881);
nor U15006 (N_15006,N_14958,N_14888);
xnor U15007 (N_15007,N_14927,N_14776);
nand U15008 (N_15008,N_14950,N_14817);
or U15009 (N_15009,N_14799,N_14790);
nor U15010 (N_15010,N_14840,N_14839);
nand U15011 (N_15011,N_14873,N_14932);
nand U15012 (N_15012,N_14957,N_14893);
and U15013 (N_15013,N_14859,N_14879);
or U15014 (N_15014,N_14903,N_14783);
nor U15015 (N_15015,N_14789,N_14919);
nand U15016 (N_15016,N_14989,N_14844);
nand U15017 (N_15017,N_14915,N_14872);
or U15018 (N_15018,N_14857,N_14983);
nand U15019 (N_15019,N_14921,N_14856);
nand U15020 (N_15020,N_14751,N_14996);
nor U15021 (N_15021,N_14901,N_14981);
or U15022 (N_15022,N_14754,N_14855);
nor U15023 (N_15023,N_14916,N_14765);
nand U15024 (N_15024,N_14926,N_14990);
nor U15025 (N_15025,N_14818,N_14775);
and U15026 (N_15026,N_14833,N_14771);
or U15027 (N_15027,N_14966,N_14761);
and U15028 (N_15028,N_14805,N_14756);
xor U15029 (N_15029,N_14952,N_14870);
nor U15030 (N_15030,N_14768,N_14836);
nand U15031 (N_15031,N_14918,N_14894);
nand U15032 (N_15032,N_14930,N_14934);
nand U15033 (N_15033,N_14871,N_14831);
and U15034 (N_15034,N_14904,N_14963);
and U15035 (N_15035,N_14794,N_14887);
or U15036 (N_15036,N_14845,N_14955);
nor U15037 (N_15037,N_14917,N_14863);
nor U15038 (N_15038,N_14835,N_14792);
nor U15039 (N_15039,N_14925,N_14793);
and U15040 (N_15040,N_14995,N_14924);
or U15041 (N_15041,N_14956,N_14820);
or U15042 (N_15042,N_14854,N_14788);
xor U15043 (N_15043,N_14774,N_14987);
and U15044 (N_15044,N_14967,N_14882);
nor U15045 (N_15045,N_14997,N_14784);
xor U15046 (N_15046,N_14808,N_14874);
nor U15047 (N_15047,N_14822,N_14898);
nand U15048 (N_15048,N_14837,N_14778);
or U15049 (N_15049,N_14762,N_14798);
and U15050 (N_15050,N_14940,N_14852);
nand U15051 (N_15051,N_14905,N_14803);
xnor U15052 (N_15052,N_14953,N_14868);
nand U15053 (N_15053,N_14912,N_14896);
xor U15054 (N_15054,N_14886,N_14962);
nor U15055 (N_15055,N_14929,N_14968);
nor U15056 (N_15056,N_14975,N_14923);
or U15057 (N_15057,N_14787,N_14867);
or U15058 (N_15058,N_14908,N_14985);
xor U15059 (N_15059,N_14801,N_14781);
nor U15060 (N_15060,N_14939,N_14976);
nor U15061 (N_15061,N_14786,N_14851);
nor U15062 (N_15062,N_14988,N_14909);
or U15063 (N_15063,N_14815,N_14782);
xor U15064 (N_15064,N_14875,N_14910);
or U15065 (N_15065,N_14861,N_14802);
and U15066 (N_15066,N_14977,N_14758);
nand U15067 (N_15067,N_14780,N_14753);
nor U15068 (N_15068,N_14797,N_14906);
nor U15069 (N_15069,N_14755,N_14865);
xnor U15070 (N_15070,N_14843,N_14942);
nor U15071 (N_15071,N_14948,N_14769);
nor U15072 (N_15072,N_14984,N_14841);
nand U15073 (N_15073,N_14827,N_14913);
nand U15074 (N_15074,N_14825,N_14877);
xnor U15075 (N_15075,N_14878,N_14949);
xor U15076 (N_15076,N_14800,N_14998);
or U15077 (N_15077,N_14848,N_14970);
nor U15078 (N_15078,N_14850,N_14809);
xor U15079 (N_15079,N_14960,N_14770);
and U15080 (N_15080,N_14806,N_14902);
nand U15081 (N_15081,N_14973,N_14796);
or U15082 (N_15082,N_14847,N_14838);
nand U15083 (N_15083,N_14933,N_14779);
or U15084 (N_15084,N_14941,N_14757);
nand U15085 (N_15085,N_14750,N_14824);
nor U15086 (N_15086,N_14971,N_14928);
xor U15087 (N_15087,N_14980,N_14829);
or U15088 (N_15088,N_14811,N_14810);
nand U15089 (N_15089,N_14821,N_14830);
xnor U15090 (N_15090,N_14954,N_14883);
xnor U15091 (N_15091,N_14931,N_14826);
xor U15092 (N_15092,N_14846,N_14935);
nand U15093 (N_15093,N_14862,N_14876);
and U15094 (N_15094,N_14764,N_14816);
nor U15095 (N_15095,N_14936,N_14858);
and U15096 (N_15096,N_14772,N_14812);
or U15097 (N_15097,N_14889,N_14993);
nand U15098 (N_15098,N_14979,N_14938);
nand U15099 (N_15099,N_14965,N_14804);
and U15100 (N_15100,N_14899,N_14914);
nand U15101 (N_15101,N_14895,N_14978);
nor U15102 (N_15102,N_14907,N_14944);
nor U15103 (N_15103,N_14884,N_14992);
nor U15104 (N_15104,N_14991,N_14763);
nand U15105 (N_15105,N_14760,N_14880);
and U15106 (N_15106,N_14767,N_14892);
and U15107 (N_15107,N_14864,N_14982);
xnor U15108 (N_15108,N_14819,N_14946);
xnor U15109 (N_15109,N_14766,N_14849);
xor U15110 (N_15110,N_14969,N_14974);
nand U15111 (N_15111,N_14814,N_14869);
nand U15112 (N_15112,N_14945,N_14897);
or U15113 (N_15113,N_14900,N_14828);
and U15114 (N_15114,N_14885,N_14911);
nand U15115 (N_15115,N_14842,N_14834);
or U15116 (N_15116,N_14866,N_14891);
xor U15117 (N_15117,N_14823,N_14860);
or U15118 (N_15118,N_14964,N_14951);
nand U15119 (N_15119,N_14986,N_14961);
and U15120 (N_15120,N_14832,N_14972);
xor U15121 (N_15121,N_14777,N_14947);
nor U15122 (N_15122,N_14813,N_14807);
or U15123 (N_15123,N_14890,N_14752);
nor U15124 (N_15124,N_14943,N_14922);
nor U15125 (N_15125,N_14870,N_14831);
or U15126 (N_15126,N_14921,N_14959);
nor U15127 (N_15127,N_14766,N_14956);
or U15128 (N_15128,N_14750,N_14859);
nand U15129 (N_15129,N_14885,N_14824);
nand U15130 (N_15130,N_14976,N_14873);
and U15131 (N_15131,N_14944,N_14852);
and U15132 (N_15132,N_14967,N_14772);
nand U15133 (N_15133,N_14857,N_14969);
nand U15134 (N_15134,N_14930,N_14927);
nor U15135 (N_15135,N_14990,N_14955);
xnor U15136 (N_15136,N_14815,N_14905);
xor U15137 (N_15137,N_14876,N_14969);
or U15138 (N_15138,N_14756,N_14998);
or U15139 (N_15139,N_14857,N_14838);
or U15140 (N_15140,N_14761,N_14750);
or U15141 (N_15141,N_14763,N_14834);
nand U15142 (N_15142,N_14845,N_14952);
or U15143 (N_15143,N_14767,N_14905);
or U15144 (N_15144,N_14953,N_14966);
nand U15145 (N_15145,N_14908,N_14972);
xor U15146 (N_15146,N_14767,N_14893);
nor U15147 (N_15147,N_14962,N_14896);
nor U15148 (N_15148,N_14806,N_14970);
nand U15149 (N_15149,N_14950,N_14896);
nand U15150 (N_15150,N_14938,N_14906);
nor U15151 (N_15151,N_14962,N_14793);
or U15152 (N_15152,N_14842,N_14960);
xor U15153 (N_15153,N_14874,N_14807);
xnor U15154 (N_15154,N_14896,N_14898);
xnor U15155 (N_15155,N_14964,N_14987);
and U15156 (N_15156,N_14883,N_14824);
nand U15157 (N_15157,N_14991,N_14975);
nand U15158 (N_15158,N_14795,N_14938);
and U15159 (N_15159,N_14970,N_14850);
xnor U15160 (N_15160,N_14920,N_14945);
and U15161 (N_15161,N_14970,N_14982);
and U15162 (N_15162,N_14999,N_14926);
xnor U15163 (N_15163,N_14909,N_14769);
xnor U15164 (N_15164,N_14783,N_14949);
and U15165 (N_15165,N_14763,N_14979);
or U15166 (N_15166,N_14985,N_14921);
and U15167 (N_15167,N_14763,N_14797);
nand U15168 (N_15168,N_14865,N_14855);
xor U15169 (N_15169,N_14932,N_14917);
and U15170 (N_15170,N_14894,N_14933);
xor U15171 (N_15171,N_14907,N_14763);
nor U15172 (N_15172,N_14789,N_14855);
nor U15173 (N_15173,N_14989,N_14901);
nand U15174 (N_15174,N_14758,N_14897);
and U15175 (N_15175,N_14888,N_14985);
xnor U15176 (N_15176,N_14848,N_14800);
and U15177 (N_15177,N_14854,N_14986);
and U15178 (N_15178,N_14773,N_14943);
and U15179 (N_15179,N_14867,N_14750);
nor U15180 (N_15180,N_14818,N_14957);
or U15181 (N_15181,N_14811,N_14771);
nand U15182 (N_15182,N_14900,N_14861);
or U15183 (N_15183,N_14902,N_14867);
nor U15184 (N_15184,N_14881,N_14919);
or U15185 (N_15185,N_14909,N_14871);
and U15186 (N_15186,N_14766,N_14975);
and U15187 (N_15187,N_14821,N_14794);
xor U15188 (N_15188,N_14849,N_14900);
and U15189 (N_15189,N_14881,N_14974);
and U15190 (N_15190,N_14857,N_14918);
or U15191 (N_15191,N_14771,N_14936);
nor U15192 (N_15192,N_14917,N_14850);
or U15193 (N_15193,N_14832,N_14771);
xnor U15194 (N_15194,N_14934,N_14758);
xor U15195 (N_15195,N_14916,N_14999);
nand U15196 (N_15196,N_14819,N_14774);
xor U15197 (N_15197,N_14772,N_14889);
xor U15198 (N_15198,N_14833,N_14867);
and U15199 (N_15199,N_14825,N_14823);
xor U15200 (N_15200,N_14957,N_14854);
nor U15201 (N_15201,N_14816,N_14866);
or U15202 (N_15202,N_14801,N_14755);
nand U15203 (N_15203,N_14862,N_14817);
xnor U15204 (N_15204,N_14833,N_14796);
or U15205 (N_15205,N_14786,N_14969);
and U15206 (N_15206,N_14779,N_14757);
nand U15207 (N_15207,N_14927,N_14816);
and U15208 (N_15208,N_14798,N_14803);
and U15209 (N_15209,N_14788,N_14968);
nor U15210 (N_15210,N_14855,N_14856);
nor U15211 (N_15211,N_14816,N_14778);
nor U15212 (N_15212,N_14785,N_14942);
nand U15213 (N_15213,N_14873,N_14871);
nand U15214 (N_15214,N_14929,N_14859);
or U15215 (N_15215,N_14882,N_14994);
nor U15216 (N_15216,N_14842,N_14855);
nor U15217 (N_15217,N_14975,N_14941);
nand U15218 (N_15218,N_14821,N_14884);
or U15219 (N_15219,N_14934,N_14947);
nand U15220 (N_15220,N_14898,N_14816);
or U15221 (N_15221,N_14784,N_14852);
or U15222 (N_15222,N_14974,N_14993);
nand U15223 (N_15223,N_14851,N_14761);
and U15224 (N_15224,N_14872,N_14843);
xor U15225 (N_15225,N_14827,N_14819);
nor U15226 (N_15226,N_14887,N_14868);
nand U15227 (N_15227,N_14908,N_14924);
xnor U15228 (N_15228,N_14908,N_14856);
xor U15229 (N_15229,N_14981,N_14850);
xnor U15230 (N_15230,N_14754,N_14866);
and U15231 (N_15231,N_14988,N_14765);
and U15232 (N_15232,N_14801,N_14766);
and U15233 (N_15233,N_14814,N_14809);
nor U15234 (N_15234,N_14761,N_14839);
nand U15235 (N_15235,N_14900,N_14931);
or U15236 (N_15236,N_14821,N_14818);
nor U15237 (N_15237,N_14943,N_14899);
nand U15238 (N_15238,N_14913,N_14826);
xnor U15239 (N_15239,N_14770,N_14766);
xnor U15240 (N_15240,N_14952,N_14937);
and U15241 (N_15241,N_14802,N_14766);
and U15242 (N_15242,N_14972,N_14789);
and U15243 (N_15243,N_14817,N_14816);
and U15244 (N_15244,N_14994,N_14807);
nand U15245 (N_15245,N_14877,N_14931);
nor U15246 (N_15246,N_14771,N_14917);
xnor U15247 (N_15247,N_14895,N_14983);
xnor U15248 (N_15248,N_14978,N_14768);
nor U15249 (N_15249,N_14882,N_14843);
nand U15250 (N_15250,N_15140,N_15003);
and U15251 (N_15251,N_15022,N_15034);
or U15252 (N_15252,N_15045,N_15060);
nand U15253 (N_15253,N_15101,N_15051);
xnor U15254 (N_15254,N_15063,N_15235);
nand U15255 (N_15255,N_15199,N_15104);
nand U15256 (N_15256,N_15075,N_15027);
nor U15257 (N_15257,N_15130,N_15085);
xnor U15258 (N_15258,N_15097,N_15114);
and U15259 (N_15259,N_15217,N_15090);
nand U15260 (N_15260,N_15044,N_15058);
or U15261 (N_15261,N_15166,N_15126);
or U15262 (N_15262,N_15247,N_15216);
nand U15263 (N_15263,N_15198,N_15206);
xnor U15264 (N_15264,N_15156,N_15076);
nor U15265 (N_15265,N_15147,N_15221);
or U15266 (N_15266,N_15132,N_15088);
nand U15267 (N_15267,N_15139,N_15202);
nand U15268 (N_15268,N_15236,N_15239);
nand U15269 (N_15269,N_15006,N_15215);
or U15270 (N_15270,N_15201,N_15127);
nor U15271 (N_15271,N_15054,N_15231);
nor U15272 (N_15272,N_15129,N_15057);
or U15273 (N_15273,N_15228,N_15071);
or U15274 (N_15274,N_15077,N_15009);
nor U15275 (N_15275,N_15030,N_15041);
nor U15276 (N_15276,N_15070,N_15010);
xnor U15277 (N_15277,N_15011,N_15190);
xnor U15278 (N_15278,N_15210,N_15117);
xor U15279 (N_15279,N_15066,N_15102);
nor U15280 (N_15280,N_15227,N_15226);
or U15281 (N_15281,N_15040,N_15175);
nor U15282 (N_15282,N_15042,N_15138);
and U15283 (N_15283,N_15246,N_15179);
xnor U15284 (N_15284,N_15092,N_15020);
nand U15285 (N_15285,N_15038,N_15214);
and U15286 (N_15286,N_15200,N_15141);
and U15287 (N_15287,N_15035,N_15144);
nand U15288 (N_15288,N_15193,N_15116);
nor U15289 (N_15289,N_15048,N_15120);
xor U15290 (N_15290,N_15103,N_15123);
nand U15291 (N_15291,N_15079,N_15136);
nor U15292 (N_15292,N_15165,N_15183);
nor U15293 (N_15293,N_15204,N_15052);
xor U15294 (N_15294,N_15238,N_15154);
nand U15295 (N_15295,N_15000,N_15118);
or U15296 (N_15296,N_15167,N_15065);
nor U15297 (N_15297,N_15068,N_15184);
nand U15298 (N_15298,N_15112,N_15033);
nand U15299 (N_15299,N_15153,N_15053);
xnor U15300 (N_15300,N_15146,N_15242);
nand U15301 (N_15301,N_15072,N_15028);
nand U15302 (N_15302,N_15212,N_15232);
and U15303 (N_15303,N_15089,N_15161);
and U15304 (N_15304,N_15149,N_15121);
xnor U15305 (N_15305,N_15111,N_15182);
nor U15306 (N_15306,N_15218,N_15082);
nor U15307 (N_15307,N_15050,N_15158);
or U15308 (N_15308,N_15081,N_15189);
nand U15309 (N_15309,N_15015,N_15135);
nor U15310 (N_15310,N_15219,N_15115);
and U15311 (N_15311,N_15017,N_15207);
and U15312 (N_15312,N_15086,N_15025);
nor U15313 (N_15313,N_15078,N_15032);
and U15314 (N_15314,N_15180,N_15014);
nand U15315 (N_15315,N_15163,N_15105);
xnor U15316 (N_15316,N_15155,N_15098);
nor U15317 (N_15317,N_15224,N_15181);
and U15318 (N_15318,N_15091,N_15145);
or U15319 (N_15319,N_15056,N_15107);
and U15320 (N_15320,N_15191,N_15241);
and U15321 (N_15321,N_15205,N_15095);
or U15322 (N_15322,N_15037,N_15229);
xor U15323 (N_15323,N_15249,N_15187);
or U15324 (N_15324,N_15016,N_15248);
and U15325 (N_15325,N_15074,N_15222);
and U15326 (N_15326,N_15099,N_15142);
nor U15327 (N_15327,N_15192,N_15172);
xor U15328 (N_15328,N_15049,N_15233);
nor U15329 (N_15329,N_15240,N_15196);
nand U15330 (N_15330,N_15237,N_15005);
or U15331 (N_15331,N_15096,N_15209);
or U15332 (N_15332,N_15084,N_15178);
or U15333 (N_15333,N_15143,N_15039);
nand U15334 (N_15334,N_15152,N_15110);
xor U15335 (N_15335,N_15245,N_15137);
xnor U15336 (N_15336,N_15124,N_15108);
or U15337 (N_15337,N_15220,N_15186);
or U15338 (N_15338,N_15160,N_15168);
xor U15339 (N_15339,N_15026,N_15159);
xor U15340 (N_15340,N_15173,N_15113);
and U15341 (N_15341,N_15083,N_15019);
nor U15342 (N_15342,N_15185,N_15195);
nand U15343 (N_15343,N_15157,N_15174);
or U15344 (N_15344,N_15094,N_15021);
xnor U15345 (N_15345,N_15059,N_15067);
nor U15346 (N_15346,N_15170,N_15064);
or U15347 (N_15347,N_15046,N_15008);
nand U15348 (N_15348,N_15002,N_15073);
nand U15349 (N_15349,N_15243,N_15119);
nor U15350 (N_15350,N_15024,N_15029);
nor U15351 (N_15351,N_15208,N_15069);
and U15352 (N_15352,N_15244,N_15131);
and U15353 (N_15353,N_15213,N_15043);
and U15354 (N_15354,N_15055,N_15177);
and U15355 (N_15355,N_15109,N_15001);
xnor U15356 (N_15356,N_15087,N_15203);
and U15357 (N_15357,N_15225,N_15047);
or U15358 (N_15358,N_15031,N_15004);
nor U15359 (N_15359,N_15007,N_15230);
or U15360 (N_15360,N_15128,N_15223);
xnor U15361 (N_15361,N_15122,N_15197);
and U15362 (N_15362,N_15061,N_15169);
or U15363 (N_15363,N_15164,N_15125);
nor U15364 (N_15364,N_15148,N_15106);
nor U15365 (N_15365,N_15012,N_15018);
nor U15366 (N_15366,N_15133,N_15134);
and U15367 (N_15367,N_15194,N_15211);
xnor U15368 (N_15368,N_15036,N_15188);
or U15369 (N_15369,N_15234,N_15023);
or U15370 (N_15370,N_15013,N_15093);
and U15371 (N_15371,N_15150,N_15162);
or U15372 (N_15372,N_15080,N_15176);
xnor U15373 (N_15373,N_15151,N_15171);
nand U15374 (N_15374,N_15100,N_15062);
or U15375 (N_15375,N_15201,N_15173);
and U15376 (N_15376,N_15221,N_15019);
nand U15377 (N_15377,N_15188,N_15032);
and U15378 (N_15378,N_15232,N_15108);
and U15379 (N_15379,N_15016,N_15148);
and U15380 (N_15380,N_15005,N_15065);
nand U15381 (N_15381,N_15239,N_15012);
xor U15382 (N_15382,N_15089,N_15126);
nor U15383 (N_15383,N_15097,N_15065);
nand U15384 (N_15384,N_15039,N_15146);
and U15385 (N_15385,N_15181,N_15149);
and U15386 (N_15386,N_15137,N_15068);
or U15387 (N_15387,N_15020,N_15226);
and U15388 (N_15388,N_15110,N_15212);
or U15389 (N_15389,N_15201,N_15194);
xnor U15390 (N_15390,N_15071,N_15118);
nor U15391 (N_15391,N_15088,N_15106);
and U15392 (N_15392,N_15138,N_15022);
or U15393 (N_15393,N_15006,N_15116);
nor U15394 (N_15394,N_15058,N_15062);
xnor U15395 (N_15395,N_15012,N_15163);
and U15396 (N_15396,N_15220,N_15229);
nand U15397 (N_15397,N_15217,N_15009);
xor U15398 (N_15398,N_15155,N_15144);
xnor U15399 (N_15399,N_15149,N_15179);
xnor U15400 (N_15400,N_15155,N_15055);
and U15401 (N_15401,N_15040,N_15045);
xor U15402 (N_15402,N_15176,N_15108);
and U15403 (N_15403,N_15179,N_15211);
or U15404 (N_15404,N_15085,N_15039);
or U15405 (N_15405,N_15070,N_15222);
nor U15406 (N_15406,N_15160,N_15039);
nor U15407 (N_15407,N_15210,N_15049);
or U15408 (N_15408,N_15055,N_15145);
nand U15409 (N_15409,N_15219,N_15211);
or U15410 (N_15410,N_15003,N_15076);
xor U15411 (N_15411,N_15236,N_15067);
nand U15412 (N_15412,N_15046,N_15029);
nor U15413 (N_15413,N_15216,N_15007);
and U15414 (N_15414,N_15079,N_15032);
nor U15415 (N_15415,N_15236,N_15230);
nand U15416 (N_15416,N_15028,N_15225);
nand U15417 (N_15417,N_15151,N_15073);
and U15418 (N_15418,N_15074,N_15159);
or U15419 (N_15419,N_15204,N_15177);
or U15420 (N_15420,N_15142,N_15169);
or U15421 (N_15421,N_15137,N_15142);
or U15422 (N_15422,N_15084,N_15073);
xnor U15423 (N_15423,N_15181,N_15104);
nand U15424 (N_15424,N_15170,N_15091);
nor U15425 (N_15425,N_15201,N_15007);
xor U15426 (N_15426,N_15170,N_15234);
xnor U15427 (N_15427,N_15240,N_15006);
or U15428 (N_15428,N_15075,N_15031);
xor U15429 (N_15429,N_15245,N_15097);
and U15430 (N_15430,N_15074,N_15209);
nor U15431 (N_15431,N_15180,N_15161);
nor U15432 (N_15432,N_15113,N_15046);
xor U15433 (N_15433,N_15102,N_15012);
nand U15434 (N_15434,N_15219,N_15230);
or U15435 (N_15435,N_15034,N_15127);
nor U15436 (N_15436,N_15181,N_15007);
or U15437 (N_15437,N_15158,N_15098);
xor U15438 (N_15438,N_15146,N_15040);
nor U15439 (N_15439,N_15017,N_15170);
nand U15440 (N_15440,N_15067,N_15088);
and U15441 (N_15441,N_15190,N_15218);
nand U15442 (N_15442,N_15060,N_15157);
and U15443 (N_15443,N_15223,N_15099);
and U15444 (N_15444,N_15122,N_15003);
nand U15445 (N_15445,N_15061,N_15230);
nand U15446 (N_15446,N_15116,N_15213);
nor U15447 (N_15447,N_15245,N_15017);
and U15448 (N_15448,N_15129,N_15037);
or U15449 (N_15449,N_15145,N_15088);
xnor U15450 (N_15450,N_15059,N_15021);
or U15451 (N_15451,N_15085,N_15159);
nand U15452 (N_15452,N_15101,N_15176);
and U15453 (N_15453,N_15163,N_15166);
or U15454 (N_15454,N_15036,N_15222);
xnor U15455 (N_15455,N_15176,N_15239);
nor U15456 (N_15456,N_15078,N_15102);
nor U15457 (N_15457,N_15071,N_15089);
xor U15458 (N_15458,N_15210,N_15032);
and U15459 (N_15459,N_15210,N_15092);
nand U15460 (N_15460,N_15168,N_15008);
or U15461 (N_15461,N_15049,N_15165);
or U15462 (N_15462,N_15222,N_15200);
nor U15463 (N_15463,N_15176,N_15102);
or U15464 (N_15464,N_15108,N_15007);
or U15465 (N_15465,N_15216,N_15113);
nor U15466 (N_15466,N_15028,N_15201);
and U15467 (N_15467,N_15201,N_15236);
nand U15468 (N_15468,N_15093,N_15095);
and U15469 (N_15469,N_15045,N_15011);
or U15470 (N_15470,N_15238,N_15145);
nand U15471 (N_15471,N_15242,N_15162);
nand U15472 (N_15472,N_15072,N_15022);
nand U15473 (N_15473,N_15196,N_15083);
nand U15474 (N_15474,N_15062,N_15106);
xor U15475 (N_15475,N_15229,N_15052);
or U15476 (N_15476,N_15007,N_15248);
nand U15477 (N_15477,N_15019,N_15087);
xor U15478 (N_15478,N_15111,N_15158);
nor U15479 (N_15479,N_15121,N_15231);
nand U15480 (N_15480,N_15186,N_15202);
and U15481 (N_15481,N_15113,N_15098);
or U15482 (N_15482,N_15120,N_15090);
nor U15483 (N_15483,N_15032,N_15018);
xor U15484 (N_15484,N_15129,N_15119);
nor U15485 (N_15485,N_15202,N_15109);
xnor U15486 (N_15486,N_15068,N_15113);
nand U15487 (N_15487,N_15203,N_15175);
or U15488 (N_15488,N_15170,N_15185);
and U15489 (N_15489,N_15187,N_15110);
nor U15490 (N_15490,N_15028,N_15093);
and U15491 (N_15491,N_15164,N_15037);
or U15492 (N_15492,N_15205,N_15165);
or U15493 (N_15493,N_15059,N_15132);
nand U15494 (N_15494,N_15203,N_15167);
xnor U15495 (N_15495,N_15172,N_15153);
nand U15496 (N_15496,N_15081,N_15147);
or U15497 (N_15497,N_15022,N_15210);
and U15498 (N_15498,N_15184,N_15117);
or U15499 (N_15499,N_15003,N_15127);
xnor U15500 (N_15500,N_15362,N_15368);
nand U15501 (N_15501,N_15267,N_15397);
or U15502 (N_15502,N_15319,N_15474);
xor U15503 (N_15503,N_15352,N_15327);
xnor U15504 (N_15504,N_15308,N_15350);
xnor U15505 (N_15505,N_15439,N_15253);
nor U15506 (N_15506,N_15365,N_15422);
xnor U15507 (N_15507,N_15460,N_15446);
or U15508 (N_15508,N_15269,N_15453);
xor U15509 (N_15509,N_15465,N_15383);
or U15510 (N_15510,N_15372,N_15386);
nor U15511 (N_15511,N_15444,N_15356);
nand U15512 (N_15512,N_15336,N_15332);
xnor U15513 (N_15513,N_15314,N_15285);
nand U15514 (N_15514,N_15326,N_15398);
xnor U15515 (N_15515,N_15447,N_15413);
or U15516 (N_15516,N_15382,N_15270);
xor U15517 (N_15517,N_15361,N_15456);
nor U15518 (N_15518,N_15400,N_15256);
and U15519 (N_15519,N_15310,N_15313);
and U15520 (N_15520,N_15379,N_15497);
and U15521 (N_15521,N_15359,N_15323);
or U15522 (N_15522,N_15292,N_15293);
nor U15523 (N_15523,N_15409,N_15298);
xnor U15524 (N_15524,N_15405,N_15481);
and U15525 (N_15525,N_15311,N_15354);
and U15526 (N_15526,N_15425,N_15433);
nor U15527 (N_15527,N_15315,N_15454);
nand U15528 (N_15528,N_15341,N_15376);
xor U15529 (N_15529,N_15324,N_15282);
xnor U15530 (N_15530,N_15363,N_15305);
or U15531 (N_15531,N_15258,N_15499);
xor U15532 (N_15532,N_15389,N_15477);
and U15533 (N_15533,N_15448,N_15492);
nor U15534 (N_15534,N_15273,N_15255);
xor U15535 (N_15535,N_15366,N_15343);
or U15536 (N_15536,N_15457,N_15264);
and U15537 (N_15537,N_15261,N_15275);
xnor U15538 (N_15538,N_15377,N_15381);
xnor U15539 (N_15539,N_15297,N_15344);
nand U15540 (N_15540,N_15334,N_15325);
nor U15541 (N_15541,N_15289,N_15342);
nand U15542 (N_15542,N_15420,N_15340);
or U15543 (N_15543,N_15452,N_15288);
xnor U15544 (N_15544,N_15318,N_15300);
and U15545 (N_15545,N_15496,N_15494);
xnor U15546 (N_15546,N_15467,N_15345);
nor U15547 (N_15547,N_15274,N_15370);
and U15548 (N_15548,N_15412,N_15445);
nand U15549 (N_15549,N_15432,N_15331);
and U15550 (N_15550,N_15329,N_15455);
nand U15551 (N_15551,N_15309,N_15280);
nor U15552 (N_15552,N_15419,N_15435);
nand U15553 (N_15553,N_15487,N_15403);
nand U15554 (N_15554,N_15428,N_15387);
xor U15555 (N_15555,N_15304,N_15424);
or U15556 (N_15556,N_15493,N_15468);
nand U15557 (N_15557,N_15283,N_15259);
nand U15558 (N_15558,N_15385,N_15260);
or U15559 (N_15559,N_15482,N_15296);
or U15560 (N_15560,N_15351,N_15367);
nand U15561 (N_15561,N_15357,N_15450);
xnor U15562 (N_15562,N_15407,N_15478);
or U15563 (N_15563,N_15265,N_15429);
and U15564 (N_15564,N_15252,N_15414);
and U15565 (N_15565,N_15479,N_15491);
nor U15566 (N_15566,N_15306,N_15371);
or U15567 (N_15567,N_15411,N_15438);
or U15568 (N_15568,N_15437,N_15312);
nand U15569 (N_15569,N_15378,N_15473);
nor U15570 (N_15570,N_15348,N_15427);
nor U15571 (N_15571,N_15401,N_15333);
xnor U15572 (N_15572,N_15287,N_15278);
nor U15573 (N_15573,N_15294,N_15335);
nand U15574 (N_15574,N_15399,N_15459);
and U15575 (N_15575,N_15408,N_15423);
and U15576 (N_15576,N_15263,N_15321);
nand U15577 (N_15577,N_15286,N_15466);
xor U15578 (N_15578,N_15488,N_15418);
nor U15579 (N_15579,N_15355,N_15347);
and U15580 (N_15580,N_15390,N_15463);
or U15581 (N_15581,N_15375,N_15251);
xnor U15582 (N_15582,N_15290,N_15328);
nand U15583 (N_15583,N_15410,N_15291);
and U15584 (N_15584,N_15281,N_15404);
xnor U15585 (N_15585,N_15489,N_15358);
nor U15586 (N_15586,N_15303,N_15380);
or U15587 (N_15587,N_15388,N_15486);
nand U15588 (N_15588,N_15475,N_15402);
nand U15589 (N_15589,N_15484,N_15373);
nor U15590 (N_15590,N_15430,N_15320);
and U15591 (N_15591,N_15470,N_15495);
nand U15592 (N_15592,N_15349,N_15472);
nor U15593 (N_15593,N_15417,N_15277);
or U15594 (N_15594,N_15346,N_15384);
xnor U15595 (N_15595,N_15483,N_15431);
xnor U15596 (N_15596,N_15369,N_15434);
nand U15597 (N_15597,N_15272,N_15421);
or U15598 (N_15598,N_15480,N_15451);
xor U15599 (N_15599,N_15442,N_15393);
xor U15600 (N_15600,N_15396,N_15449);
and U15601 (N_15601,N_15316,N_15301);
and U15602 (N_15602,N_15469,N_15307);
or U15603 (N_15603,N_15353,N_15257);
xor U15604 (N_15604,N_15317,N_15276);
nand U15605 (N_15605,N_15266,N_15471);
xnor U15606 (N_15606,N_15443,N_15406);
nor U15607 (N_15607,N_15392,N_15426);
xnor U15608 (N_15608,N_15415,N_15458);
xnor U15609 (N_15609,N_15284,N_15498);
xor U15610 (N_15610,N_15250,N_15374);
and U15611 (N_15611,N_15339,N_15360);
nor U15612 (N_15612,N_15462,N_15338);
and U15613 (N_15613,N_15440,N_15302);
xor U15614 (N_15614,N_15299,N_15337);
xor U15615 (N_15615,N_15441,N_15262);
nor U15616 (N_15616,N_15395,N_15476);
xor U15617 (N_15617,N_15436,N_15490);
nand U15618 (N_15618,N_15330,N_15391);
or U15619 (N_15619,N_15461,N_15271);
nor U15620 (N_15620,N_15322,N_15268);
xnor U15621 (N_15621,N_15464,N_15394);
or U15622 (N_15622,N_15279,N_15295);
or U15623 (N_15623,N_15254,N_15485);
nor U15624 (N_15624,N_15364,N_15416);
and U15625 (N_15625,N_15481,N_15284);
xnor U15626 (N_15626,N_15376,N_15412);
nand U15627 (N_15627,N_15289,N_15304);
nor U15628 (N_15628,N_15418,N_15467);
and U15629 (N_15629,N_15469,N_15382);
nand U15630 (N_15630,N_15285,N_15489);
xor U15631 (N_15631,N_15424,N_15260);
nand U15632 (N_15632,N_15460,N_15289);
nand U15633 (N_15633,N_15445,N_15368);
and U15634 (N_15634,N_15251,N_15447);
nor U15635 (N_15635,N_15425,N_15400);
nor U15636 (N_15636,N_15362,N_15383);
or U15637 (N_15637,N_15355,N_15270);
nand U15638 (N_15638,N_15468,N_15499);
nor U15639 (N_15639,N_15400,N_15405);
xnor U15640 (N_15640,N_15330,N_15420);
nor U15641 (N_15641,N_15457,N_15357);
nor U15642 (N_15642,N_15396,N_15344);
or U15643 (N_15643,N_15309,N_15430);
xor U15644 (N_15644,N_15348,N_15377);
xnor U15645 (N_15645,N_15330,N_15259);
nand U15646 (N_15646,N_15280,N_15312);
or U15647 (N_15647,N_15427,N_15381);
xnor U15648 (N_15648,N_15275,N_15423);
and U15649 (N_15649,N_15308,N_15346);
nand U15650 (N_15650,N_15362,N_15413);
nand U15651 (N_15651,N_15335,N_15283);
nor U15652 (N_15652,N_15498,N_15288);
nor U15653 (N_15653,N_15431,N_15403);
nand U15654 (N_15654,N_15481,N_15466);
or U15655 (N_15655,N_15440,N_15346);
nor U15656 (N_15656,N_15281,N_15297);
nand U15657 (N_15657,N_15285,N_15438);
and U15658 (N_15658,N_15390,N_15314);
and U15659 (N_15659,N_15491,N_15495);
or U15660 (N_15660,N_15416,N_15435);
or U15661 (N_15661,N_15364,N_15291);
and U15662 (N_15662,N_15463,N_15451);
nand U15663 (N_15663,N_15464,N_15485);
or U15664 (N_15664,N_15301,N_15383);
and U15665 (N_15665,N_15265,N_15287);
and U15666 (N_15666,N_15260,N_15297);
and U15667 (N_15667,N_15359,N_15298);
or U15668 (N_15668,N_15283,N_15255);
xnor U15669 (N_15669,N_15418,N_15444);
nand U15670 (N_15670,N_15381,N_15400);
xor U15671 (N_15671,N_15473,N_15486);
and U15672 (N_15672,N_15473,N_15294);
xnor U15673 (N_15673,N_15393,N_15254);
nand U15674 (N_15674,N_15266,N_15367);
xnor U15675 (N_15675,N_15418,N_15285);
and U15676 (N_15676,N_15307,N_15374);
nand U15677 (N_15677,N_15328,N_15378);
and U15678 (N_15678,N_15376,N_15262);
or U15679 (N_15679,N_15392,N_15256);
nor U15680 (N_15680,N_15489,N_15493);
nor U15681 (N_15681,N_15280,N_15362);
and U15682 (N_15682,N_15418,N_15257);
xor U15683 (N_15683,N_15326,N_15381);
nand U15684 (N_15684,N_15403,N_15379);
nor U15685 (N_15685,N_15387,N_15430);
nand U15686 (N_15686,N_15318,N_15380);
nor U15687 (N_15687,N_15417,N_15397);
xor U15688 (N_15688,N_15296,N_15288);
or U15689 (N_15689,N_15276,N_15371);
nor U15690 (N_15690,N_15499,N_15281);
nand U15691 (N_15691,N_15320,N_15327);
xor U15692 (N_15692,N_15420,N_15275);
or U15693 (N_15693,N_15485,N_15384);
or U15694 (N_15694,N_15327,N_15460);
nor U15695 (N_15695,N_15261,N_15291);
or U15696 (N_15696,N_15355,N_15297);
nand U15697 (N_15697,N_15390,N_15298);
xnor U15698 (N_15698,N_15277,N_15453);
nand U15699 (N_15699,N_15297,N_15310);
xnor U15700 (N_15700,N_15444,N_15481);
or U15701 (N_15701,N_15267,N_15259);
nand U15702 (N_15702,N_15422,N_15380);
or U15703 (N_15703,N_15302,N_15391);
and U15704 (N_15704,N_15409,N_15424);
nand U15705 (N_15705,N_15356,N_15315);
nor U15706 (N_15706,N_15375,N_15373);
or U15707 (N_15707,N_15420,N_15284);
nand U15708 (N_15708,N_15345,N_15361);
nand U15709 (N_15709,N_15350,N_15306);
and U15710 (N_15710,N_15394,N_15358);
nand U15711 (N_15711,N_15309,N_15300);
or U15712 (N_15712,N_15434,N_15282);
nor U15713 (N_15713,N_15307,N_15448);
nand U15714 (N_15714,N_15340,N_15489);
nor U15715 (N_15715,N_15351,N_15346);
nand U15716 (N_15716,N_15427,N_15470);
nor U15717 (N_15717,N_15283,N_15287);
nand U15718 (N_15718,N_15357,N_15292);
nand U15719 (N_15719,N_15381,N_15463);
xor U15720 (N_15720,N_15305,N_15273);
xnor U15721 (N_15721,N_15268,N_15360);
and U15722 (N_15722,N_15290,N_15292);
and U15723 (N_15723,N_15341,N_15349);
or U15724 (N_15724,N_15347,N_15495);
and U15725 (N_15725,N_15295,N_15326);
nand U15726 (N_15726,N_15253,N_15349);
xnor U15727 (N_15727,N_15273,N_15319);
xor U15728 (N_15728,N_15317,N_15345);
xor U15729 (N_15729,N_15440,N_15463);
xnor U15730 (N_15730,N_15383,N_15495);
and U15731 (N_15731,N_15404,N_15385);
xor U15732 (N_15732,N_15456,N_15422);
and U15733 (N_15733,N_15365,N_15259);
and U15734 (N_15734,N_15301,N_15288);
and U15735 (N_15735,N_15338,N_15472);
nand U15736 (N_15736,N_15282,N_15387);
xnor U15737 (N_15737,N_15378,N_15274);
xor U15738 (N_15738,N_15441,N_15404);
or U15739 (N_15739,N_15330,N_15352);
and U15740 (N_15740,N_15297,N_15425);
and U15741 (N_15741,N_15394,N_15440);
nand U15742 (N_15742,N_15378,N_15393);
xor U15743 (N_15743,N_15445,N_15320);
nand U15744 (N_15744,N_15470,N_15494);
and U15745 (N_15745,N_15428,N_15331);
nand U15746 (N_15746,N_15463,N_15269);
xnor U15747 (N_15747,N_15398,N_15390);
xor U15748 (N_15748,N_15300,N_15430);
or U15749 (N_15749,N_15495,N_15477);
and U15750 (N_15750,N_15670,N_15649);
and U15751 (N_15751,N_15584,N_15641);
nor U15752 (N_15752,N_15608,N_15738);
and U15753 (N_15753,N_15697,N_15744);
xnor U15754 (N_15754,N_15685,N_15524);
nand U15755 (N_15755,N_15633,N_15729);
xnor U15756 (N_15756,N_15538,N_15630);
xnor U15757 (N_15757,N_15740,N_15725);
and U15758 (N_15758,N_15735,N_15518);
and U15759 (N_15759,N_15508,N_15691);
or U15760 (N_15760,N_15620,N_15663);
nor U15761 (N_15761,N_15515,N_15673);
nor U15762 (N_15762,N_15732,N_15650);
and U15763 (N_15763,N_15568,N_15619);
nand U15764 (N_15764,N_15644,N_15696);
nor U15765 (N_15765,N_15601,N_15539);
or U15766 (N_15766,N_15571,N_15566);
nor U15767 (N_15767,N_15546,N_15593);
and U15768 (N_15768,N_15737,N_15733);
nand U15769 (N_15769,N_15526,N_15639);
and U15770 (N_15770,N_15537,N_15646);
xnor U15771 (N_15771,N_15569,N_15509);
nand U15772 (N_15772,N_15564,N_15627);
nand U15773 (N_15773,N_15731,N_15565);
xnor U15774 (N_15774,N_15596,N_15623);
xor U15775 (N_15775,N_15578,N_15614);
nor U15776 (N_15776,N_15712,N_15617);
nor U15777 (N_15777,N_15552,N_15561);
xor U15778 (N_15778,N_15511,N_15698);
xor U15779 (N_15779,N_15536,N_15654);
nand U15780 (N_15780,N_15616,N_15553);
nor U15781 (N_15781,N_15651,N_15675);
or U15782 (N_15782,N_15545,N_15555);
or U15783 (N_15783,N_15661,N_15704);
nand U15784 (N_15784,N_15688,N_15559);
xnor U15785 (N_15785,N_15530,N_15551);
or U15786 (N_15786,N_15581,N_15507);
xnor U15787 (N_15787,N_15629,N_15582);
and U15788 (N_15788,N_15741,N_15557);
nand U15789 (N_15789,N_15607,N_15513);
xor U15790 (N_15790,N_15525,N_15647);
nor U15791 (N_15791,N_15631,N_15703);
xor U15792 (N_15792,N_15637,N_15626);
xnor U15793 (N_15793,N_15501,N_15597);
nor U15794 (N_15794,N_15594,N_15664);
nand U15795 (N_15795,N_15628,N_15726);
nor U15796 (N_15796,N_15622,N_15715);
and U15797 (N_15797,N_15684,N_15589);
and U15798 (N_15798,N_15745,N_15656);
and U15799 (N_15799,N_15632,N_15672);
nor U15800 (N_15800,N_15611,N_15541);
or U15801 (N_15801,N_15747,N_15516);
or U15802 (N_15802,N_15723,N_15610);
xnor U15803 (N_15803,N_15587,N_15682);
nor U15804 (N_15804,N_15570,N_15638);
or U15805 (N_15805,N_15576,N_15668);
or U15806 (N_15806,N_15573,N_15603);
or U15807 (N_15807,N_15567,N_15636);
or U15808 (N_15808,N_15572,N_15544);
xor U15809 (N_15809,N_15677,N_15635);
nor U15810 (N_15810,N_15739,N_15599);
nor U15811 (N_15811,N_15542,N_15579);
nor U15812 (N_15812,N_15709,N_15583);
nand U15813 (N_15813,N_15728,N_15692);
nand U15814 (N_15814,N_15681,N_15727);
or U15815 (N_15815,N_15535,N_15621);
or U15816 (N_15816,N_15618,N_15529);
and U15817 (N_15817,N_15592,N_15547);
or U15818 (N_15818,N_15543,N_15674);
nor U15819 (N_15819,N_15743,N_15716);
xor U15820 (N_15820,N_15522,N_15520);
and U15821 (N_15821,N_15640,N_15687);
nand U15822 (N_15822,N_15720,N_15724);
and U15823 (N_15823,N_15734,N_15708);
nand U15824 (N_15824,N_15604,N_15658);
and U15825 (N_15825,N_15690,N_15588);
xor U15826 (N_15826,N_15707,N_15503);
or U15827 (N_15827,N_15694,N_15642);
nor U15828 (N_15828,N_15502,N_15563);
nand U15829 (N_15829,N_15676,N_15742);
xnor U15830 (N_15830,N_15577,N_15580);
or U15831 (N_15831,N_15605,N_15648);
or U15832 (N_15832,N_15714,N_15519);
or U15833 (N_15833,N_15711,N_15686);
xnor U15834 (N_15834,N_15506,N_15510);
and U15835 (N_15835,N_15527,N_15562);
or U15836 (N_15836,N_15534,N_15625);
and U15837 (N_15837,N_15730,N_15615);
nor U15838 (N_15838,N_15624,N_15595);
xnor U15839 (N_15839,N_15693,N_15598);
or U15840 (N_15840,N_15655,N_15667);
xor U15841 (N_15841,N_15512,N_15533);
or U15842 (N_15842,N_15585,N_15556);
and U15843 (N_15843,N_15689,N_15531);
nor U15844 (N_15844,N_15700,N_15575);
xnor U15845 (N_15845,N_15748,N_15721);
nand U15846 (N_15846,N_15722,N_15736);
xnor U15847 (N_15847,N_15710,N_15548);
and U15848 (N_15848,N_15634,N_15532);
nand U15849 (N_15849,N_15591,N_15528);
xnor U15850 (N_15850,N_15662,N_15659);
nand U15851 (N_15851,N_15521,N_15657);
and U15852 (N_15852,N_15549,N_15701);
xor U15853 (N_15853,N_15713,N_15590);
nor U15854 (N_15854,N_15678,N_15560);
nand U15855 (N_15855,N_15613,N_15602);
nand U15856 (N_15856,N_15669,N_15660);
nor U15857 (N_15857,N_15717,N_15705);
nand U15858 (N_15858,N_15702,N_15523);
and U15859 (N_15859,N_15550,N_15665);
nor U15860 (N_15860,N_15666,N_15719);
nand U15861 (N_15861,N_15653,N_15517);
xnor U15862 (N_15862,N_15558,N_15612);
and U15863 (N_15863,N_15746,N_15574);
or U15864 (N_15864,N_15683,N_15680);
xor U15865 (N_15865,N_15679,N_15606);
and U15866 (N_15866,N_15695,N_15671);
or U15867 (N_15867,N_15706,N_15600);
nand U15868 (N_15868,N_15540,N_15554);
xnor U15869 (N_15869,N_15699,N_15586);
nor U15870 (N_15870,N_15609,N_15749);
and U15871 (N_15871,N_15505,N_15504);
xnor U15872 (N_15872,N_15645,N_15652);
nand U15873 (N_15873,N_15643,N_15514);
or U15874 (N_15874,N_15718,N_15500);
nor U15875 (N_15875,N_15601,N_15606);
nand U15876 (N_15876,N_15689,N_15643);
nand U15877 (N_15877,N_15651,N_15556);
and U15878 (N_15878,N_15540,N_15603);
nand U15879 (N_15879,N_15598,N_15624);
and U15880 (N_15880,N_15606,N_15670);
xor U15881 (N_15881,N_15583,N_15505);
or U15882 (N_15882,N_15504,N_15701);
and U15883 (N_15883,N_15548,N_15503);
nor U15884 (N_15884,N_15572,N_15639);
and U15885 (N_15885,N_15657,N_15501);
and U15886 (N_15886,N_15644,N_15667);
and U15887 (N_15887,N_15652,N_15684);
or U15888 (N_15888,N_15601,N_15744);
nor U15889 (N_15889,N_15609,N_15716);
xnor U15890 (N_15890,N_15500,N_15692);
and U15891 (N_15891,N_15554,N_15524);
nor U15892 (N_15892,N_15550,N_15604);
and U15893 (N_15893,N_15705,N_15617);
nor U15894 (N_15894,N_15580,N_15606);
nor U15895 (N_15895,N_15554,N_15574);
nor U15896 (N_15896,N_15645,N_15710);
and U15897 (N_15897,N_15581,N_15688);
nor U15898 (N_15898,N_15575,N_15602);
or U15899 (N_15899,N_15536,N_15533);
xor U15900 (N_15900,N_15580,N_15640);
or U15901 (N_15901,N_15689,N_15715);
nor U15902 (N_15902,N_15656,N_15584);
xnor U15903 (N_15903,N_15606,N_15687);
nor U15904 (N_15904,N_15573,N_15684);
and U15905 (N_15905,N_15576,N_15524);
xnor U15906 (N_15906,N_15632,N_15721);
nor U15907 (N_15907,N_15723,N_15524);
xor U15908 (N_15908,N_15675,N_15629);
or U15909 (N_15909,N_15666,N_15623);
or U15910 (N_15910,N_15708,N_15698);
xnor U15911 (N_15911,N_15672,N_15522);
nand U15912 (N_15912,N_15565,N_15548);
or U15913 (N_15913,N_15510,N_15615);
nor U15914 (N_15914,N_15664,N_15694);
and U15915 (N_15915,N_15681,N_15675);
xor U15916 (N_15916,N_15655,N_15685);
nand U15917 (N_15917,N_15543,N_15545);
nand U15918 (N_15918,N_15628,N_15584);
nand U15919 (N_15919,N_15589,N_15641);
or U15920 (N_15920,N_15611,N_15533);
or U15921 (N_15921,N_15692,N_15633);
nor U15922 (N_15922,N_15542,N_15531);
or U15923 (N_15923,N_15589,N_15501);
or U15924 (N_15924,N_15654,N_15574);
and U15925 (N_15925,N_15700,N_15708);
nor U15926 (N_15926,N_15631,N_15570);
or U15927 (N_15927,N_15685,N_15520);
and U15928 (N_15928,N_15560,N_15602);
and U15929 (N_15929,N_15526,N_15704);
or U15930 (N_15930,N_15702,N_15605);
and U15931 (N_15931,N_15727,N_15703);
and U15932 (N_15932,N_15613,N_15723);
xnor U15933 (N_15933,N_15629,N_15564);
nand U15934 (N_15934,N_15730,N_15715);
nor U15935 (N_15935,N_15566,N_15716);
xor U15936 (N_15936,N_15508,N_15703);
and U15937 (N_15937,N_15678,N_15723);
xor U15938 (N_15938,N_15528,N_15714);
nor U15939 (N_15939,N_15589,N_15653);
xnor U15940 (N_15940,N_15740,N_15535);
xor U15941 (N_15941,N_15525,N_15739);
and U15942 (N_15942,N_15576,N_15530);
or U15943 (N_15943,N_15679,N_15726);
nand U15944 (N_15944,N_15720,N_15696);
or U15945 (N_15945,N_15550,N_15614);
xnor U15946 (N_15946,N_15500,N_15573);
and U15947 (N_15947,N_15715,N_15691);
nand U15948 (N_15948,N_15671,N_15595);
xor U15949 (N_15949,N_15746,N_15591);
nand U15950 (N_15950,N_15584,N_15504);
xor U15951 (N_15951,N_15639,N_15603);
or U15952 (N_15952,N_15598,N_15716);
and U15953 (N_15953,N_15570,N_15746);
xor U15954 (N_15954,N_15718,N_15679);
and U15955 (N_15955,N_15593,N_15691);
or U15956 (N_15956,N_15584,N_15519);
nor U15957 (N_15957,N_15739,N_15523);
and U15958 (N_15958,N_15531,N_15559);
nor U15959 (N_15959,N_15675,N_15505);
xnor U15960 (N_15960,N_15686,N_15541);
nor U15961 (N_15961,N_15721,N_15621);
nand U15962 (N_15962,N_15507,N_15599);
nand U15963 (N_15963,N_15731,N_15508);
xnor U15964 (N_15964,N_15681,N_15679);
nand U15965 (N_15965,N_15696,N_15501);
or U15966 (N_15966,N_15514,N_15678);
nor U15967 (N_15967,N_15610,N_15628);
nor U15968 (N_15968,N_15672,N_15574);
or U15969 (N_15969,N_15562,N_15566);
xor U15970 (N_15970,N_15652,N_15743);
or U15971 (N_15971,N_15608,N_15677);
or U15972 (N_15972,N_15544,N_15694);
or U15973 (N_15973,N_15515,N_15631);
xnor U15974 (N_15974,N_15543,N_15743);
xnor U15975 (N_15975,N_15618,N_15737);
xnor U15976 (N_15976,N_15578,N_15725);
or U15977 (N_15977,N_15529,N_15547);
nor U15978 (N_15978,N_15708,N_15670);
xor U15979 (N_15979,N_15741,N_15529);
nand U15980 (N_15980,N_15640,N_15674);
or U15981 (N_15981,N_15579,N_15716);
xnor U15982 (N_15982,N_15739,N_15655);
or U15983 (N_15983,N_15566,N_15549);
or U15984 (N_15984,N_15523,N_15509);
xnor U15985 (N_15985,N_15533,N_15684);
and U15986 (N_15986,N_15640,N_15501);
nor U15987 (N_15987,N_15722,N_15659);
nand U15988 (N_15988,N_15504,N_15642);
nor U15989 (N_15989,N_15663,N_15666);
nand U15990 (N_15990,N_15527,N_15725);
or U15991 (N_15991,N_15725,N_15517);
and U15992 (N_15992,N_15724,N_15737);
and U15993 (N_15993,N_15727,N_15540);
and U15994 (N_15994,N_15559,N_15548);
and U15995 (N_15995,N_15734,N_15509);
nand U15996 (N_15996,N_15535,N_15726);
or U15997 (N_15997,N_15660,N_15564);
and U15998 (N_15998,N_15708,N_15689);
or U15999 (N_15999,N_15733,N_15508);
nand U16000 (N_16000,N_15917,N_15815);
nor U16001 (N_16001,N_15993,N_15903);
and U16002 (N_16002,N_15851,N_15850);
nand U16003 (N_16003,N_15871,N_15929);
and U16004 (N_16004,N_15803,N_15829);
xor U16005 (N_16005,N_15797,N_15808);
nand U16006 (N_16006,N_15837,N_15763);
nor U16007 (N_16007,N_15793,N_15933);
nor U16008 (N_16008,N_15774,N_15858);
or U16009 (N_16009,N_15819,N_15839);
or U16010 (N_16010,N_15824,N_15985);
or U16011 (N_16011,N_15990,N_15776);
and U16012 (N_16012,N_15771,N_15884);
or U16013 (N_16013,N_15977,N_15897);
xnor U16014 (N_16014,N_15923,N_15843);
xnor U16015 (N_16015,N_15809,N_15992);
nand U16016 (N_16016,N_15865,N_15930);
nor U16017 (N_16017,N_15986,N_15826);
xor U16018 (N_16018,N_15787,N_15972);
nor U16019 (N_16019,N_15994,N_15874);
or U16020 (N_16020,N_15879,N_15791);
and U16021 (N_16021,N_15991,N_15764);
nor U16022 (N_16022,N_15881,N_15833);
nor U16023 (N_16023,N_15947,N_15875);
or U16024 (N_16024,N_15788,N_15877);
nor U16025 (N_16025,N_15867,N_15913);
nand U16026 (N_16026,N_15946,N_15887);
or U16027 (N_16027,N_15810,N_15880);
nand U16028 (N_16028,N_15860,N_15770);
and U16029 (N_16029,N_15785,N_15959);
and U16030 (N_16030,N_15854,N_15998);
and U16031 (N_16031,N_15928,N_15900);
nor U16032 (N_16032,N_15934,N_15910);
nor U16033 (N_16033,N_15957,N_15869);
nor U16034 (N_16034,N_15790,N_15940);
or U16035 (N_16035,N_15795,N_15907);
nand U16036 (N_16036,N_15984,N_15909);
or U16037 (N_16037,N_15766,N_15817);
xnor U16038 (N_16038,N_15813,N_15948);
xnor U16039 (N_16039,N_15779,N_15757);
nand U16040 (N_16040,N_15845,N_15896);
nor U16041 (N_16041,N_15894,N_15944);
or U16042 (N_16042,N_15796,N_15921);
nand U16043 (N_16043,N_15798,N_15836);
nor U16044 (N_16044,N_15827,N_15772);
or U16045 (N_16045,N_15830,N_15769);
or U16046 (N_16046,N_15925,N_15814);
and U16047 (N_16047,N_15898,N_15762);
and U16048 (N_16048,N_15767,N_15890);
nor U16049 (N_16049,N_15778,N_15859);
nor U16050 (N_16050,N_15806,N_15954);
or U16051 (N_16051,N_15939,N_15799);
or U16052 (N_16052,N_15752,N_15842);
nor U16053 (N_16053,N_15783,N_15982);
xnor U16054 (N_16054,N_15932,N_15963);
xor U16055 (N_16055,N_15773,N_15807);
or U16056 (N_16056,N_15960,N_15840);
xnor U16057 (N_16057,N_15918,N_15951);
or U16058 (N_16058,N_15758,N_15961);
and U16059 (N_16059,N_15885,N_15983);
nor U16060 (N_16060,N_15943,N_15822);
and U16061 (N_16061,N_15996,N_15846);
xnor U16062 (N_16062,N_15852,N_15765);
xor U16063 (N_16063,N_15811,N_15883);
xor U16064 (N_16064,N_15886,N_15755);
and U16065 (N_16065,N_15892,N_15831);
nand U16066 (N_16066,N_15756,N_15927);
xnor U16067 (N_16067,N_15812,N_15849);
nand U16068 (N_16068,N_15878,N_15981);
nor U16069 (N_16069,N_15834,N_15955);
and U16070 (N_16070,N_15792,N_15856);
and U16071 (N_16071,N_15864,N_15825);
nor U16072 (N_16072,N_15821,N_15926);
or U16073 (N_16073,N_15978,N_15848);
nor U16074 (N_16074,N_15802,N_15781);
nand U16075 (N_16075,N_15924,N_15823);
nand U16076 (N_16076,N_15868,N_15901);
nor U16077 (N_16077,N_15820,N_15968);
nand U16078 (N_16078,N_15838,N_15979);
nand U16079 (N_16079,N_15976,N_15751);
xor U16080 (N_16080,N_15876,N_15780);
or U16081 (N_16081,N_15953,N_15789);
or U16082 (N_16082,N_15966,N_15862);
nor U16083 (N_16083,N_15818,N_15899);
or U16084 (N_16084,N_15967,N_15841);
xnor U16085 (N_16085,N_15935,N_15942);
or U16086 (N_16086,N_15888,N_15902);
or U16087 (N_16087,N_15989,N_15904);
nor U16088 (N_16088,N_15750,N_15988);
nand U16089 (N_16089,N_15995,N_15987);
or U16090 (N_16090,N_15949,N_15853);
and U16091 (N_16091,N_15753,N_15777);
or U16092 (N_16092,N_15801,N_15941);
and U16093 (N_16093,N_15919,N_15794);
xnor U16094 (N_16094,N_15945,N_15754);
and U16095 (N_16095,N_15759,N_15805);
xor U16096 (N_16096,N_15958,N_15970);
or U16097 (N_16097,N_15962,N_15975);
xor U16098 (N_16098,N_15956,N_15905);
and U16099 (N_16099,N_15964,N_15916);
nor U16100 (N_16100,N_15950,N_15893);
nor U16101 (N_16101,N_15873,N_15855);
and U16102 (N_16102,N_15914,N_15782);
xor U16103 (N_16103,N_15863,N_15908);
xor U16104 (N_16104,N_15784,N_15931);
and U16105 (N_16105,N_15816,N_15889);
nand U16106 (N_16106,N_15997,N_15761);
nand U16107 (N_16107,N_15915,N_15895);
nand U16108 (N_16108,N_15912,N_15911);
nand U16109 (N_16109,N_15832,N_15969);
or U16110 (N_16110,N_15866,N_15760);
nor U16111 (N_16111,N_15882,N_15775);
and U16112 (N_16112,N_15870,N_15906);
or U16113 (N_16113,N_15973,N_15872);
nand U16114 (N_16114,N_15800,N_15980);
nor U16115 (N_16115,N_15835,N_15847);
xnor U16116 (N_16116,N_15938,N_15965);
or U16117 (N_16117,N_15857,N_15999);
and U16118 (N_16118,N_15937,N_15922);
nand U16119 (N_16119,N_15786,N_15971);
or U16120 (N_16120,N_15861,N_15920);
and U16121 (N_16121,N_15768,N_15891);
xor U16122 (N_16122,N_15936,N_15974);
xor U16123 (N_16123,N_15952,N_15844);
xor U16124 (N_16124,N_15804,N_15828);
or U16125 (N_16125,N_15790,N_15795);
nand U16126 (N_16126,N_15771,N_15899);
nor U16127 (N_16127,N_15906,N_15802);
or U16128 (N_16128,N_15877,N_15752);
and U16129 (N_16129,N_15861,N_15809);
or U16130 (N_16130,N_15814,N_15792);
or U16131 (N_16131,N_15779,N_15768);
and U16132 (N_16132,N_15954,N_15888);
nand U16133 (N_16133,N_15818,N_15873);
nand U16134 (N_16134,N_15948,N_15877);
xnor U16135 (N_16135,N_15865,N_15829);
or U16136 (N_16136,N_15800,N_15916);
and U16137 (N_16137,N_15916,N_15945);
xnor U16138 (N_16138,N_15844,N_15981);
nor U16139 (N_16139,N_15909,N_15787);
nor U16140 (N_16140,N_15820,N_15838);
xor U16141 (N_16141,N_15996,N_15930);
xnor U16142 (N_16142,N_15809,N_15873);
or U16143 (N_16143,N_15831,N_15845);
nor U16144 (N_16144,N_15988,N_15757);
and U16145 (N_16145,N_15956,N_15840);
xor U16146 (N_16146,N_15862,N_15777);
and U16147 (N_16147,N_15900,N_15898);
xnor U16148 (N_16148,N_15916,N_15773);
and U16149 (N_16149,N_15959,N_15800);
nand U16150 (N_16150,N_15776,N_15958);
or U16151 (N_16151,N_15930,N_15892);
nand U16152 (N_16152,N_15943,N_15906);
nand U16153 (N_16153,N_15781,N_15988);
and U16154 (N_16154,N_15753,N_15887);
nor U16155 (N_16155,N_15903,N_15927);
and U16156 (N_16156,N_15820,N_15879);
and U16157 (N_16157,N_15986,N_15772);
and U16158 (N_16158,N_15808,N_15836);
nand U16159 (N_16159,N_15901,N_15946);
xnor U16160 (N_16160,N_15901,N_15859);
xor U16161 (N_16161,N_15934,N_15974);
and U16162 (N_16162,N_15853,N_15754);
and U16163 (N_16163,N_15933,N_15974);
nand U16164 (N_16164,N_15968,N_15920);
or U16165 (N_16165,N_15818,N_15980);
and U16166 (N_16166,N_15935,N_15762);
nand U16167 (N_16167,N_15917,N_15986);
or U16168 (N_16168,N_15875,N_15852);
xor U16169 (N_16169,N_15800,N_15870);
and U16170 (N_16170,N_15991,N_15913);
and U16171 (N_16171,N_15950,N_15855);
and U16172 (N_16172,N_15997,N_15891);
and U16173 (N_16173,N_15884,N_15869);
and U16174 (N_16174,N_15751,N_15750);
and U16175 (N_16175,N_15830,N_15932);
xor U16176 (N_16176,N_15913,N_15944);
nand U16177 (N_16177,N_15900,N_15850);
and U16178 (N_16178,N_15774,N_15862);
or U16179 (N_16179,N_15908,N_15813);
nand U16180 (N_16180,N_15899,N_15844);
and U16181 (N_16181,N_15993,N_15851);
nand U16182 (N_16182,N_15996,N_15927);
nor U16183 (N_16183,N_15840,N_15818);
and U16184 (N_16184,N_15910,N_15773);
nand U16185 (N_16185,N_15923,N_15789);
nor U16186 (N_16186,N_15884,N_15901);
nand U16187 (N_16187,N_15904,N_15887);
nand U16188 (N_16188,N_15928,N_15862);
nor U16189 (N_16189,N_15750,N_15844);
nand U16190 (N_16190,N_15887,N_15757);
xnor U16191 (N_16191,N_15781,N_15968);
and U16192 (N_16192,N_15885,N_15783);
nor U16193 (N_16193,N_15902,N_15821);
and U16194 (N_16194,N_15973,N_15997);
nand U16195 (N_16195,N_15815,N_15899);
nor U16196 (N_16196,N_15858,N_15951);
nor U16197 (N_16197,N_15839,N_15788);
nor U16198 (N_16198,N_15953,N_15763);
and U16199 (N_16199,N_15808,N_15776);
nor U16200 (N_16200,N_15857,N_15834);
nand U16201 (N_16201,N_15952,N_15852);
nor U16202 (N_16202,N_15874,N_15950);
or U16203 (N_16203,N_15799,N_15870);
or U16204 (N_16204,N_15954,N_15830);
xor U16205 (N_16205,N_15810,N_15830);
and U16206 (N_16206,N_15778,N_15917);
nor U16207 (N_16207,N_15990,N_15918);
nand U16208 (N_16208,N_15866,N_15849);
xnor U16209 (N_16209,N_15963,N_15810);
and U16210 (N_16210,N_15880,N_15894);
and U16211 (N_16211,N_15861,N_15956);
nand U16212 (N_16212,N_15757,N_15771);
or U16213 (N_16213,N_15829,N_15878);
or U16214 (N_16214,N_15950,N_15766);
and U16215 (N_16215,N_15923,N_15834);
or U16216 (N_16216,N_15814,N_15999);
and U16217 (N_16217,N_15874,N_15958);
or U16218 (N_16218,N_15842,N_15910);
or U16219 (N_16219,N_15846,N_15763);
or U16220 (N_16220,N_15977,N_15776);
or U16221 (N_16221,N_15781,N_15835);
or U16222 (N_16222,N_15831,N_15846);
or U16223 (N_16223,N_15888,N_15851);
xnor U16224 (N_16224,N_15767,N_15772);
nand U16225 (N_16225,N_15829,N_15949);
xor U16226 (N_16226,N_15847,N_15958);
nor U16227 (N_16227,N_15856,N_15752);
nor U16228 (N_16228,N_15822,N_15961);
xnor U16229 (N_16229,N_15814,N_15785);
xnor U16230 (N_16230,N_15930,N_15888);
nand U16231 (N_16231,N_15782,N_15898);
nor U16232 (N_16232,N_15755,N_15847);
nand U16233 (N_16233,N_15827,N_15835);
and U16234 (N_16234,N_15781,N_15928);
or U16235 (N_16235,N_15773,N_15867);
xor U16236 (N_16236,N_15923,N_15962);
and U16237 (N_16237,N_15927,N_15965);
xnor U16238 (N_16238,N_15974,N_15875);
nand U16239 (N_16239,N_15921,N_15759);
xor U16240 (N_16240,N_15802,N_15785);
and U16241 (N_16241,N_15996,N_15755);
xor U16242 (N_16242,N_15855,N_15996);
nand U16243 (N_16243,N_15895,N_15854);
nand U16244 (N_16244,N_15910,N_15800);
or U16245 (N_16245,N_15814,N_15984);
xor U16246 (N_16246,N_15905,N_15884);
nand U16247 (N_16247,N_15830,N_15991);
nor U16248 (N_16248,N_15846,N_15887);
xor U16249 (N_16249,N_15852,N_15861);
nand U16250 (N_16250,N_16123,N_16003);
nand U16251 (N_16251,N_16243,N_16033);
xnor U16252 (N_16252,N_16107,N_16129);
and U16253 (N_16253,N_16011,N_16166);
nand U16254 (N_16254,N_16085,N_16108);
nand U16255 (N_16255,N_16002,N_16088);
xor U16256 (N_16256,N_16144,N_16241);
nor U16257 (N_16257,N_16074,N_16201);
or U16258 (N_16258,N_16006,N_16235);
xor U16259 (N_16259,N_16190,N_16245);
or U16260 (N_16260,N_16221,N_16032);
nand U16261 (N_16261,N_16207,N_16179);
xnor U16262 (N_16262,N_16117,N_16073);
nor U16263 (N_16263,N_16130,N_16185);
nor U16264 (N_16264,N_16008,N_16023);
nand U16265 (N_16265,N_16173,N_16214);
and U16266 (N_16266,N_16019,N_16169);
or U16267 (N_16267,N_16204,N_16180);
nor U16268 (N_16268,N_16212,N_16047);
and U16269 (N_16269,N_16194,N_16138);
and U16270 (N_16270,N_16048,N_16225);
nand U16271 (N_16271,N_16058,N_16043);
nor U16272 (N_16272,N_16065,N_16103);
or U16273 (N_16273,N_16086,N_16186);
nor U16274 (N_16274,N_16104,N_16210);
nand U16275 (N_16275,N_16059,N_16247);
nand U16276 (N_16276,N_16052,N_16215);
xnor U16277 (N_16277,N_16010,N_16066);
nor U16278 (N_16278,N_16157,N_16229);
nand U16279 (N_16279,N_16249,N_16097);
nand U16280 (N_16280,N_16139,N_16147);
xnor U16281 (N_16281,N_16203,N_16209);
nand U16282 (N_16282,N_16146,N_16191);
nand U16283 (N_16283,N_16051,N_16055);
and U16284 (N_16284,N_16087,N_16044);
nor U16285 (N_16285,N_16234,N_16145);
or U16286 (N_16286,N_16135,N_16198);
nor U16287 (N_16287,N_16216,N_16132);
nand U16288 (N_16288,N_16165,N_16184);
nand U16289 (N_16289,N_16125,N_16140);
or U16290 (N_16290,N_16031,N_16178);
nor U16291 (N_16291,N_16056,N_16028);
and U16292 (N_16292,N_16098,N_16197);
nand U16293 (N_16293,N_16057,N_16054);
nor U16294 (N_16294,N_16038,N_16025);
and U16295 (N_16295,N_16187,N_16168);
and U16296 (N_16296,N_16183,N_16211);
nor U16297 (N_16297,N_16072,N_16005);
and U16298 (N_16298,N_16127,N_16174);
and U16299 (N_16299,N_16000,N_16099);
xnor U16300 (N_16300,N_16136,N_16120);
and U16301 (N_16301,N_16239,N_16017);
nor U16302 (N_16302,N_16218,N_16142);
xnor U16303 (N_16303,N_16071,N_16004);
xor U16304 (N_16304,N_16100,N_16018);
and U16305 (N_16305,N_16077,N_16222);
and U16306 (N_16306,N_16062,N_16037);
nor U16307 (N_16307,N_16200,N_16206);
nor U16308 (N_16308,N_16030,N_16115);
and U16309 (N_16309,N_16102,N_16213);
xnor U16310 (N_16310,N_16164,N_16172);
and U16311 (N_16311,N_16228,N_16192);
xnor U16312 (N_16312,N_16069,N_16177);
xnor U16313 (N_16313,N_16248,N_16149);
and U16314 (N_16314,N_16068,N_16022);
xnor U16315 (N_16315,N_16237,N_16095);
or U16316 (N_16316,N_16193,N_16230);
nor U16317 (N_16317,N_16133,N_16067);
nor U16318 (N_16318,N_16199,N_16233);
and U16319 (N_16319,N_16009,N_16153);
nor U16320 (N_16320,N_16171,N_16111);
nand U16321 (N_16321,N_16126,N_16015);
xor U16322 (N_16322,N_16134,N_16106);
and U16323 (N_16323,N_16114,N_16001);
xnor U16324 (N_16324,N_16110,N_16195);
xor U16325 (N_16325,N_16161,N_16188);
and U16326 (N_16326,N_16090,N_16202);
nor U16327 (N_16327,N_16049,N_16079);
and U16328 (N_16328,N_16205,N_16232);
xnor U16329 (N_16329,N_16013,N_16040);
nor U16330 (N_16330,N_16121,N_16116);
xnor U16331 (N_16331,N_16094,N_16113);
or U16332 (N_16332,N_16039,N_16167);
xnor U16333 (N_16333,N_16151,N_16101);
xnor U16334 (N_16334,N_16109,N_16093);
and U16335 (N_16335,N_16159,N_16208);
nand U16336 (N_16336,N_16224,N_16124);
nand U16337 (N_16337,N_16170,N_16020);
or U16338 (N_16338,N_16176,N_16112);
and U16339 (N_16339,N_16089,N_16105);
or U16340 (N_16340,N_16246,N_16143);
or U16341 (N_16341,N_16220,N_16026);
xor U16342 (N_16342,N_16118,N_16155);
or U16343 (N_16343,N_16091,N_16189);
xor U16344 (N_16344,N_16046,N_16227);
nor U16345 (N_16345,N_16223,N_16137);
xnor U16346 (N_16346,N_16182,N_16148);
nor U16347 (N_16347,N_16084,N_16240);
or U16348 (N_16348,N_16150,N_16141);
nor U16349 (N_16349,N_16175,N_16119);
nor U16350 (N_16350,N_16029,N_16236);
nand U16351 (N_16351,N_16082,N_16050);
xor U16352 (N_16352,N_16219,N_16080);
nor U16353 (N_16353,N_16092,N_16162);
or U16354 (N_16354,N_16007,N_16231);
nand U16355 (N_16355,N_16045,N_16128);
nor U16356 (N_16356,N_16163,N_16060);
nand U16357 (N_16357,N_16063,N_16061);
nand U16358 (N_16358,N_16036,N_16226);
nor U16359 (N_16359,N_16242,N_16027);
nand U16360 (N_16360,N_16083,N_16064);
xor U16361 (N_16361,N_16041,N_16053);
nand U16362 (N_16362,N_16244,N_16152);
or U16363 (N_16363,N_16160,N_16076);
xor U16364 (N_16364,N_16131,N_16075);
or U16365 (N_16365,N_16024,N_16035);
xor U16366 (N_16366,N_16016,N_16181);
nor U16367 (N_16367,N_16081,N_16070);
nand U16368 (N_16368,N_16034,N_16217);
nor U16369 (N_16369,N_16021,N_16238);
nand U16370 (N_16370,N_16096,N_16122);
or U16371 (N_16371,N_16196,N_16012);
nor U16372 (N_16372,N_16042,N_16078);
or U16373 (N_16373,N_16154,N_16014);
xnor U16374 (N_16374,N_16156,N_16158);
xnor U16375 (N_16375,N_16040,N_16016);
nand U16376 (N_16376,N_16230,N_16240);
xnor U16377 (N_16377,N_16029,N_16088);
nor U16378 (N_16378,N_16151,N_16242);
or U16379 (N_16379,N_16010,N_16205);
xor U16380 (N_16380,N_16105,N_16202);
nand U16381 (N_16381,N_16117,N_16235);
nor U16382 (N_16382,N_16218,N_16059);
nand U16383 (N_16383,N_16065,N_16145);
nor U16384 (N_16384,N_16202,N_16125);
nor U16385 (N_16385,N_16201,N_16219);
nor U16386 (N_16386,N_16072,N_16235);
nor U16387 (N_16387,N_16008,N_16099);
and U16388 (N_16388,N_16204,N_16118);
or U16389 (N_16389,N_16034,N_16047);
xnor U16390 (N_16390,N_16212,N_16087);
and U16391 (N_16391,N_16178,N_16187);
or U16392 (N_16392,N_16203,N_16010);
and U16393 (N_16393,N_16033,N_16131);
and U16394 (N_16394,N_16115,N_16086);
or U16395 (N_16395,N_16220,N_16226);
nor U16396 (N_16396,N_16245,N_16023);
xor U16397 (N_16397,N_16011,N_16000);
nand U16398 (N_16398,N_16224,N_16174);
or U16399 (N_16399,N_16152,N_16030);
or U16400 (N_16400,N_16206,N_16043);
or U16401 (N_16401,N_16070,N_16047);
and U16402 (N_16402,N_16210,N_16183);
nand U16403 (N_16403,N_16110,N_16200);
nand U16404 (N_16404,N_16035,N_16221);
nor U16405 (N_16405,N_16195,N_16025);
nor U16406 (N_16406,N_16200,N_16236);
nand U16407 (N_16407,N_16155,N_16124);
and U16408 (N_16408,N_16042,N_16020);
nor U16409 (N_16409,N_16082,N_16107);
and U16410 (N_16410,N_16162,N_16035);
xor U16411 (N_16411,N_16072,N_16126);
xor U16412 (N_16412,N_16123,N_16069);
or U16413 (N_16413,N_16229,N_16130);
nor U16414 (N_16414,N_16199,N_16060);
nor U16415 (N_16415,N_16162,N_16120);
xor U16416 (N_16416,N_16235,N_16183);
xor U16417 (N_16417,N_16242,N_16238);
or U16418 (N_16418,N_16093,N_16240);
nand U16419 (N_16419,N_16021,N_16176);
nand U16420 (N_16420,N_16186,N_16239);
and U16421 (N_16421,N_16016,N_16052);
nor U16422 (N_16422,N_16202,N_16058);
xnor U16423 (N_16423,N_16147,N_16095);
and U16424 (N_16424,N_16001,N_16078);
and U16425 (N_16425,N_16031,N_16126);
and U16426 (N_16426,N_16049,N_16065);
or U16427 (N_16427,N_16043,N_16222);
nor U16428 (N_16428,N_16240,N_16012);
and U16429 (N_16429,N_16103,N_16091);
nand U16430 (N_16430,N_16045,N_16231);
xnor U16431 (N_16431,N_16068,N_16221);
xnor U16432 (N_16432,N_16117,N_16234);
or U16433 (N_16433,N_16153,N_16133);
and U16434 (N_16434,N_16061,N_16222);
or U16435 (N_16435,N_16082,N_16108);
or U16436 (N_16436,N_16074,N_16230);
or U16437 (N_16437,N_16147,N_16069);
and U16438 (N_16438,N_16088,N_16077);
xor U16439 (N_16439,N_16011,N_16236);
xnor U16440 (N_16440,N_16069,N_16063);
nand U16441 (N_16441,N_16246,N_16004);
nor U16442 (N_16442,N_16236,N_16167);
nand U16443 (N_16443,N_16185,N_16201);
nand U16444 (N_16444,N_16065,N_16114);
and U16445 (N_16445,N_16217,N_16149);
and U16446 (N_16446,N_16117,N_16155);
and U16447 (N_16447,N_16237,N_16078);
xor U16448 (N_16448,N_16122,N_16165);
xnor U16449 (N_16449,N_16135,N_16095);
nand U16450 (N_16450,N_16141,N_16149);
nor U16451 (N_16451,N_16053,N_16131);
nand U16452 (N_16452,N_16026,N_16178);
nand U16453 (N_16453,N_16197,N_16028);
nand U16454 (N_16454,N_16239,N_16045);
or U16455 (N_16455,N_16195,N_16058);
xor U16456 (N_16456,N_16068,N_16015);
and U16457 (N_16457,N_16233,N_16065);
xnor U16458 (N_16458,N_16180,N_16048);
and U16459 (N_16459,N_16186,N_16243);
nor U16460 (N_16460,N_16201,N_16038);
or U16461 (N_16461,N_16172,N_16003);
nand U16462 (N_16462,N_16072,N_16160);
nor U16463 (N_16463,N_16084,N_16147);
nor U16464 (N_16464,N_16079,N_16077);
nor U16465 (N_16465,N_16155,N_16205);
nor U16466 (N_16466,N_16150,N_16011);
xnor U16467 (N_16467,N_16009,N_16006);
xor U16468 (N_16468,N_16193,N_16007);
nand U16469 (N_16469,N_16142,N_16195);
nor U16470 (N_16470,N_16022,N_16146);
nor U16471 (N_16471,N_16020,N_16126);
or U16472 (N_16472,N_16240,N_16008);
xor U16473 (N_16473,N_16131,N_16211);
and U16474 (N_16474,N_16044,N_16208);
nor U16475 (N_16475,N_16199,N_16118);
and U16476 (N_16476,N_16053,N_16180);
and U16477 (N_16477,N_16013,N_16128);
and U16478 (N_16478,N_16198,N_16126);
or U16479 (N_16479,N_16042,N_16094);
xnor U16480 (N_16480,N_16136,N_16194);
or U16481 (N_16481,N_16027,N_16129);
and U16482 (N_16482,N_16176,N_16125);
or U16483 (N_16483,N_16189,N_16174);
xor U16484 (N_16484,N_16191,N_16010);
nand U16485 (N_16485,N_16008,N_16161);
xnor U16486 (N_16486,N_16202,N_16161);
nor U16487 (N_16487,N_16139,N_16035);
xor U16488 (N_16488,N_16143,N_16004);
nor U16489 (N_16489,N_16012,N_16245);
and U16490 (N_16490,N_16117,N_16167);
nor U16491 (N_16491,N_16212,N_16007);
and U16492 (N_16492,N_16128,N_16034);
xor U16493 (N_16493,N_16127,N_16007);
nor U16494 (N_16494,N_16240,N_16149);
nand U16495 (N_16495,N_16002,N_16095);
or U16496 (N_16496,N_16093,N_16135);
and U16497 (N_16497,N_16224,N_16094);
nor U16498 (N_16498,N_16002,N_16224);
xnor U16499 (N_16499,N_16219,N_16120);
and U16500 (N_16500,N_16349,N_16355);
xor U16501 (N_16501,N_16340,N_16401);
or U16502 (N_16502,N_16296,N_16478);
xor U16503 (N_16503,N_16266,N_16325);
xnor U16504 (N_16504,N_16333,N_16301);
or U16505 (N_16505,N_16458,N_16286);
nor U16506 (N_16506,N_16343,N_16384);
or U16507 (N_16507,N_16405,N_16308);
xnor U16508 (N_16508,N_16294,N_16251);
nor U16509 (N_16509,N_16411,N_16434);
xnor U16510 (N_16510,N_16475,N_16331);
nand U16511 (N_16511,N_16389,N_16435);
and U16512 (N_16512,N_16302,N_16408);
nor U16513 (N_16513,N_16276,N_16469);
nand U16514 (N_16514,N_16414,N_16412);
nor U16515 (N_16515,N_16299,N_16400);
xor U16516 (N_16516,N_16317,N_16256);
nand U16517 (N_16517,N_16413,N_16375);
or U16518 (N_16518,N_16278,N_16318);
or U16519 (N_16519,N_16374,N_16303);
nor U16520 (N_16520,N_16494,N_16270);
xor U16521 (N_16521,N_16330,N_16338);
nor U16522 (N_16522,N_16269,N_16427);
nand U16523 (N_16523,N_16298,N_16311);
xor U16524 (N_16524,N_16394,N_16432);
and U16525 (N_16525,N_16257,N_16277);
or U16526 (N_16526,N_16390,N_16290);
nand U16527 (N_16527,N_16329,N_16463);
xnor U16528 (N_16528,N_16357,N_16382);
nor U16529 (N_16529,N_16319,N_16387);
or U16530 (N_16530,N_16467,N_16391);
nor U16531 (N_16531,N_16441,N_16309);
nand U16532 (N_16532,N_16466,N_16352);
or U16533 (N_16533,N_16465,N_16313);
or U16534 (N_16534,N_16315,N_16356);
xnor U16535 (N_16535,N_16380,N_16446);
and U16536 (N_16536,N_16392,N_16407);
xor U16537 (N_16537,N_16457,N_16451);
xnor U16538 (N_16538,N_16292,N_16496);
or U16539 (N_16539,N_16273,N_16284);
nor U16540 (N_16540,N_16481,N_16404);
or U16541 (N_16541,N_16271,N_16422);
nand U16542 (N_16542,N_16450,N_16279);
nor U16543 (N_16543,N_16474,N_16351);
or U16544 (N_16544,N_16342,N_16486);
nand U16545 (N_16545,N_16366,N_16485);
or U16546 (N_16546,N_16267,N_16250);
or U16547 (N_16547,N_16425,N_16498);
nor U16548 (N_16548,N_16370,N_16321);
and U16549 (N_16549,N_16473,N_16454);
nor U16550 (N_16550,N_16281,N_16310);
nor U16551 (N_16551,N_16381,N_16259);
and U16552 (N_16552,N_16283,N_16472);
nand U16553 (N_16553,N_16344,N_16499);
nor U16554 (N_16554,N_16448,N_16345);
nor U16555 (N_16555,N_16376,N_16272);
and U16556 (N_16556,N_16490,N_16263);
or U16557 (N_16557,N_16341,N_16488);
xor U16558 (N_16558,N_16287,N_16265);
nand U16559 (N_16559,N_16462,N_16395);
xor U16560 (N_16560,N_16452,N_16274);
or U16561 (N_16561,N_16449,N_16420);
nand U16562 (N_16562,N_16445,N_16360);
nor U16563 (N_16563,N_16346,N_16388);
nor U16564 (N_16564,N_16397,N_16428);
nor U16565 (N_16565,N_16305,N_16323);
or U16566 (N_16566,N_16406,N_16489);
or U16567 (N_16567,N_16368,N_16455);
nand U16568 (N_16568,N_16484,N_16495);
and U16569 (N_16569,N_16470,N_16419);
xor U16570 (N_16570,N_16453,N_16437);
and U16571 (N_16571,N_16433,N_16476);
xor U16572 (N_16572,N_16385,N_16430);
nor U16573 (N_16573,N_16289,N_16254);
nor U16574 (N_16574,N_16261,N_16324);
xnor U16575 (N_16575,N_16275,N_16363);
xnor U16576 (N_16576,N_16365,N_16328);
nor U16577 (N_16577,N_16264,N_16399);
xor U16578 (N_16578,N_16334,N_16402);
xnor U16579 (N_16579,N_16300,N_16461);
and U16580 (N_16580,N_16378,N_16326);
nor U16581 (N_16581,N_16436,N_16447);
or U16582 (N_16582,N_16354,N_16493);
and U16583 (N_16583,N_16285,N_16373);
nor U16584 (N_16584,N_16314,N_16280);
and U16585 (N_16585,N_16253,N_16492);
xnor U16586 (N_16586,N_16255,N_16336);
nand U16587 (N_16587,N_16377,N_16398);
nor U16588 (N_16588,N_16379,N_16480);
nor U16589 (N_16589,N_16293,N_16297);
or U16590 (N_16590,N_16393,N_16369);
xor U16591 (N_16591,N_16483,N_16347);
xor U16592 (N_16592,N_16282,N_16464);
nor U16593 (N_16593,N_16403,N_16304);
xor U16594 (N_16594,N_16337,N_16295);
or U16595 (N_16595,N_16383,N_16396);
or U16596 (N_16596,N_16440,N_16262);
nor U16597 (N_16597,N_16335,N_16418);
nand U16598 (N_16598,N_16339,N_16438);
xnor U16599 (N_16599,N_16471,N_16362);
and U16600 (N_16600,N_16477,N_16386);
and U16601 (N_16601,N_16364,N_16367);
nor U16602 (N_16602,N_16415,N_16306);
and U16603 (N_16603,N_16361,N_16497);
xor U16604 (N_16604,N_16459,N_16348);
or U16605 (N_16605,N_16487,N_16258);
and U16606 (N_16606,N_16431,N_16409);
nand U16607 (N_16607,N_16332,N_16316);
nor U16608 (N_16608,N_16312,N_16353);
nand U16609 (N_16609,N_16307,N_16288);
and U16610 (N_16610,N_16291,N_16350);
or U16611 (N_16611,N_16443,N_16442);
nor U16612 (N_16612,N_16460,N_16327);
or U16613 (N_16613,N_16456,N_16358);
xnor U16614 (N_16614,N_16320,N_16423);
nor U16615 (N_16615,N_16417,N_16372);
xnor U16616 (N_16616,N_16482,N_16439);
or U16617 (N_16617,N_16426,N_16424);
xor U16618 (N_16618,N_16359,N_16468);
or U16619 (N_16619,N_16491,N_16322);
nor U16620 (N_16620,N_16479,N_16444);
nand U16621 (N_16621,N_16268,N_16371);
nor U16622 (N_16622,N_16260,N_16421);
xor U16623 (N_16623,N_16252,N_16416);
nand U16624 (N_16624,N_16410,N_16429);
nand U16625 (N_16625,N_16471,N_16370);
or U16626 (N_16626,N_16304,N_16337);
and U16627 (N_16627,N_16446,N_16475);
nor U16628 (N_16628,N_16426,N_16299);
or U16629 (N_16629,N_16405,N_16266);
or U16630 (N_16630,N_16316,N_16487);
nor U16631 (N_16631,N_16463,N_16455);
nor U16632 (N_16632,N_16406,N_16424);
nor U16633 (N_16633,N_16383,N_16329);
nand U16634 (N_16634,N_16439,N_16348);
and U16635 (N_16635,N_16397,N_16392);
nor U16636 (N_16636,N_16418,N_16410);
nand U16637 (N_16637,N_16253,N_16311);
and U16638 (N_16638,N_16284,N_16260);
nor U16639 (N_16639,N_16404,N_16329);
xor U16640 (N_16640,N_16354,N_16478);
or U16641 (N_16641,N_16253,N_16413);
xor U16642 (N_16642,N_16431,N_16396);
or U16643 (N_16643,N_16320,N_16323);
nand U16644 (N_16644,N_16320,N_16273);
and U16645 (N_16645,N_16302,N_16414);
nor U16646 (N_16646,N_16409,N_16256);
nand U16647 (N_16647,N_16443,N_16251);
xnor U16648 (N_16648,N_16263,N_16409);
nand U16649 (N_16649,N_16457,N_16276);
nor U16650 (N_16650,N_16388,N_16347);
or U16651 (N_16651,N_16398,N_16333);
nand U16652 (N_16652,N_16326,N_16256);
and U16653 (N_16653,N_16464,N_16439);
or U16654 (N_16654,N_16492,N_16411);
and U16655 (N_16655,N_16396,N_16439);
nand U16656 (N_16656,N_16416,N_16250);
and U16657 (N_16657,N_16454,N_16334);
nor U16658 (N_16658,N_16489,N_16363);
and U16659 (N_16659,N_16378,N_16332);
xor U16660 (N_16660,N_16328,N_16493);
nor U16661 (N_16661,N_16476,N_16412);
nor U16662 (N_16662,N_16316,N_16448);
xor U16663 (N_16663,N_16449,N_16288);
nand U16664 (N_16664,N_16356,N_16499);
and U16665 (N_16665,N_16316,N_16329);
nor U16666 (N_16666,N_16496,N_16449);
nand U16667 (N_16667,N_16367,N_16332);
and U16668 (N_16668,N_16389,N_16366);
or U16669 (N_16669,N_16418,N_16298);
and U16670 (N_16670,N_16255,N_16314);
and U16671 (N_16671,N_16451,N_16443);
xor U16672 (N_16672,N_16280,N_16302);
xnor U16673 (N_16673,N_16389,N_16318);
nor U16674 (N_16674,N_16364,N_16304);
nand U16675 (N_16675,N_16283,N_16473);
nand U16676 (N_16676,N_16268,N_16441);
or U16677 (N_16677,N_16330,N_16334);
nor U16678 (N_16678,N_16372,N_16334);
or U16679 (N_16679,N_16434,N_16327);
or U16680 (N_16680,N_16398,N_16314);
and U16681 (N_16681,N_16365,N_16268);
and U16682 (N_16682,N_16485,N_16395);
nor U16683 (N_16683,N_16333,N_16277);
nand U16684 (N_16684,N_16403,N_16371);
xnor U16685 (N_16685,N_16316,N_16291);
or U16686 (N_16686,N_16462,N_16481);
nor U16687 (N_16687,N_16436,N_16455);
xor U16688 (N_16688,N_16258,N_16260);
or U16689 (N_16689,N_16334,N_16489);
or U16690 (N_16690,N_16380,N_16343);
nand U16691 (N_16691,N_16421,N_16250);
xor U16692 (N_16692,N_16476,N_16486);
xnor U16693 (N_16693,N_16488,N_16347);
or U16694 (N_16694,N_16473,N_16265);
nor U16695 (N_16695,N_16279,N_16251);
xor U16696 (N_16696,N_16476,N_16302);
and U16697 (N_16697,N_16460,N_16421);
nand U16698 (N_16698,N_16263,N_16332);
xor U16699 (N_16699,N_16397,N_16422);
nand U16700 (N_16700,N_16437,N_16341);
xnor U16701 (N_16701,N_16469,N_16303);
or U16702 (N_16702,N_16299,N_16286);
and U16703 (N_16703,N_16436,N_16429);
xnor U16704 (N_16704,N_16365,N_16302);
nand U16705 (N_16705,N_16492,N_16439);
and U16706 (N_16706,N_16458,N_16424);
or U16707 (N_16707,N_16490,N_16436);
nand U16708 (N_16708,N_16295,N_16340);
or U16709 (N_16709,N_16385,N_16446);
or U16710 (N_16710,N_16427,N_16374);
nand U16711 (N_16711,N_16416,N_16395);
nor U16712 (N_16712,N_16451,N_16370);
xnor U16713 (N_16713,N_16448,N_16466);
xor U16714 (N_16714,N_16361,N_16400);
nor U16715 (N_16715,N_16341,N_16261);
nand U16716 (N_16716,N_16282,N_16258);
nand U16717 (N_16717,N_16478,N_16415);
and U16718 (N_16718,N_16436,N_16337);
nor U16719 (N_16719,N_16471,N_16482);
and U16720 (N_16720,N_16307,N_16497);
nand U16721 (N_16721,N_16330,N_16496);
or U16722 (N_16722,N_16342,N_16351);
xnor U16723 (N_16723,N_16478,N_16338);
xnor U16724 (N_16724,N_16463,N_16433);
nand U16725 (N_16725,N_16349,N_16459);
and U16726 (N_16726,N_16288,N_16358);
or U16727 (N_16727,N_16412,N_16374);
or U16728 (N_16728,N_16315,N_16496);
nor U16729 (N_16729,N_16320,N_16364);
and U16730 (N_16730,N_16363,N_16343);
xor U16731 (N_16731,N_16252,N_16449);
xnor U16732 (N_16732,N_16311,N_16373);
xnor U16733 (N_16733,N_16254,N_16463);
xor U16734 (N_16734,N_16395,N_16402);
and U16735 (N_16735,N_16327,N_16310);
nor U16736 (N_16736,N_16363,N_16369);
nand U16737 (N_16737,N_16363,N_16472);
nand U16738 (N_16738,N_16281,N_16458);
and U16739 (N_16739,N_16436,N_16274);
nand U16740 (N_16740,N_16476,N_16447);
and U16741 (N_16741,N_16474,N_16283);
xnor U16742 (N_16742,N_16377,N_16404);
and U16743 (N_16743,N_16266,N_16487);
xor U16744 (N_16744,N_16346,N_16385);
nand U16745 (N_16745,N_16361,N_16336);
nor U16746 (N_16746,N_16299,N_16387);
nor U16747 (N_16747,N_16453,N_16446);
nand U16748 (N_16748,N_16484,N_16464);
and U16749 (N_16749,N_16460,N_16431);
nor U16750 (N_16750,N_16705,N_16703);
xnor U16751 (N_16751,N_16584,N_16716);
and U16752 (N_16752,N_16637,N_16537);
nand U16753 (N_16753,N_16598,N_16518);
nor U16754 (N_16754,N_16531,N_16694);
nor U16755 (N_16755,N_16513,N_16578);
xor U16756 (N_16756,N_16670,N_16674);
or U16757 (N_16757,N_16546,N_16742);
or U16758 (N_16758,N_16579,N_16559);
or U16759 (N_16759,N_16693,N_16515);
and U16760 (N_16760,N_16718,N_16627);
and U16761 (N_16761,N_16534,N_16591);
nor U16762 (N_16762,N_16508,N_16565);
nand U16763 (N_16763,N_16672,N_16741);
xor U16764 (N_16764,N_16553,N_16687);
nand U16765 (N_16765,N_16618,N_16509);
nor U16766 (N_16766,N_16695,N_16569);
and U16767 (N_16767,N_16549,N_16572);
xnor U16768 (N_16768,N_16512,N_16628);
nand U16769 (N_16769,N_16738,N_16630);
or U16770 (N_16770,N_16570,N_16737);
or U16771 (N_16771,N_16558,N_16673);
nand U16772 (N_16772,N_16679,N_16600);
nor U16773 (N_16773,N_16526,N_16568);
or U16774 (N_16774,N_16676,N_16721);
and U16775 (N_16775,N_16587,N_16582);
nor U16776 (N_16776,N_16659,N_16711);
nor U16777 (N_16777,N_16664,N_16543);
or U16778 (N_16778,N_16624,N_16617);
and U16779 (N_16779,N_16655,N_16644);
xor U16780 (N_16780,N_16744,N_16654);
or U16781 (N_16781,N_16653,N_16682);
nor U16782 (N_16782,N_16723,N_16639);
and U16783 (N_16783,N_16564,N_16666);
nor U16784 (N_16784,N_16671,N_16532);
or U16785 (N_16785,N_16593,N_16510);
nor U16786 (N_16786,N_16697,N_16590);
xnor U16787 (N_16787,N_16580,N_16658);
xnor U16788 (N_16788,N_16541,N_16610);
or U16789 (N_16789,N_16503,N_16739);
and U16790 (N_16790,N_16522,N_16749);
or U16791 (N_16791,N_16520,N_16605);
nand U16792 (N_16792,N_16606,N_16634);
or U16793 (N_16793,N_16609,N_16608);
and U16794 (N_16794,N_16714,N_16715);
nand U16795 (N_16795,N_16523,N_16560);
nor U16796 (N_16796,N_16648,N_16640);
and U16797 (N_16797,N_16542,N_16677);
nand U16798 (N_16798,N_16733,N_16571);
nor U16799 (N_16799,N_16688,N_16575);
nor U16800 (N_16800,N_16625,N_16528);
and U16801 (N_16801,N_16726,N_16743);
xor U16802 (N_16802,N_16650,N_16686);
and U16803 (N_16803,N_16588,N_16597);
nand U16804 (N_16804,N_16651,N_16663);
or U16805 (N_16805,N_16599,N_16595);
nand U16806 (N_16806,N_16667,N_16616);
and U16807 (N_16807,N_16709,N_16636);
and U16808 (N_16808,N_16533,N_16689);
xnor U16809 (N_16809,N_16529,N_16561);
nor U16810 (N_16810,N_16535,N_16736);
nand U16811 (N_16811,N_16719,N_16727);
and U16812 (N_16812,N_16585,N_16538);
nor U16813 (N_16813,N_16621,N_16657);
xnor U16814 (N_16814,N_16581,N_16620);
and U16815 (N_16815,N_16698,N_16574);
xnor U16816 (N_16816,N_16551,N_16554);
nand U16817 (N_16817,N_16746,N_16517);
xor U16818 (N_16818,N_16725,N_16665);
nand U16819 (N_16819,N_16652,N_16740);
nand U16820 (N_16820,N_16619,N_16586);
nand U16821 (N_16821,N_16681,N_16516);
nor U16822 (N_16822,N_16615,N_16557);
or U16823 (N_16823,N_16638,N_16603);
and U16824 (N_16824,N_16685,N_16507);
or U16825 (N_16825,N_16552,N_16730);
and U16826 (N_16826,N_16647,N_16556);
or U16827 (N_16827,N_16562,N_16717);
nor U16828 (N_16828,N_16734,N_16583);
nand U16829 (N_16829,N_16661,N_16708);
and U16830 (N_16830,N_16521,N_16645);
or U16831 (N_16831,N_16530,N_16635);
nor U16832 (N_16832,N_16505,N_16712);
nand U16833 (N_16833,N_16613,N_16700);
nor U16834 (N_16834,N_16643,N_16612);
or U16835 (N_16835,N_16631,N_16641);
and U16836 (N_16836,N_16544,N_16539);
nand U16837 (N_16837,N_16504,N_16622);
or U16838 (N_16838,N_16500,N_16547);
xnor U16839 (N_16839,N_16576,N_16669);
and U16840 (N_16840,N_16735,N_16592);
or U16841 (N_16841,N_16601,N_16745);
nor U16842 (N_16842,N_16626,N_16524);
nor U16843 (N_16843,N_16511,N_16589);
xor U16844 (N_16844,N_16713,N_16614);
and U16845 (N_16845,N_16692,N_16649);
nand U16846 (N_16846,N_16602,N_16690);
xnor U16847 (N_16847,N_16633,N_16567);
nor U16848 (N_16848,N_16632,N_16550);
and U16849 (N_16849,N_16660,N_16604);
nor U16850 (N_16850,N_16548,N_16696);
and U16851 (N_16851,N_16701,N_16707);
and U16852 (N_16852,N_16536,N_16678);
nor U16853 (N_16853,N_16720,N_16577);
xnor U16854 (N_16854,N_16566,N_16748);
nand U16855 (N_16855,N_16680,N_16747);
nand U16856 (N_16856,N_16729,N_16668);
and U16857 (N_16857,N_16540,N_16646);
xnor U16858 (N_16858,N_16656,N_16611);
and U16859 (N_16859,N_16691,N_16642);
or U16860 (N_16860,N_16728,N_16594);
and U16861 (N_16861,N_16684,N_16662);
nand U16862 (N_16862,N_16501,N_16596);
and U16863 (N_16863,N_16629,N_16699);
nand U16864 (N_16864,N_16527,N_16545);
xnor U16865 (N_16865,N_16519,N_16710);
nor U16866 (N_16866,N_16514,N_16731);
and U16867 (N_16867,N_16607,N_16573);
nor U16868 (N_16868,N_16525,N_16704);
or U16869 (N_16869,N_16506,N_16683);
nor U16870 (N_16870,N_16623,N_16675);
nand U16871 (N_16871,N_16706,N_16702);
and U16872 (N_16872,N_16722,N_16502);
nand U16873 (N_16873,N_16724,N_16563);
or U16874 (N_16874,N_16732,N_16555);
nor U16875 (N_16875,N_16629,N_16669);
nor U16876 (N_16876,N_16689,N_16591);
and U16877 (N_16877,N_16732,N_16520);
or U16878 (N_16878,N_16654,N_16593);
xor U16879 (N_16879,N_16539,N_16536);
and U16880 (N_16880,N_16744,N_16573);
or U16881 (N_16881,N_16606,N_16726);
nor U16882 (N_16882,N_16572,N_16744);
xnor U16883 (N_16883,N_16572,N_16745);
xor U16884 (N_16884,N_16630,N_16656);
and U16885 (N_16885,N_16659,N_16563);
xnor U16886 (N_16886,N_16512,N_16723);
and U16887 (N_16887,N_16731,N_16712);
xnor U16888 (N_16888,N_16637,N_16627);
or U16889 (N_16889,N_16552,N_16598);
and U16890 (N_16890,N_16736,N_16727);
nand U16891 (N_16891,N_16511,N_16502);
nand U16892 (N_16892,N_16527,N_16646);
nand U16893 (N_16893,N_16564,N_16579);
xor U16894 (N_16894,N_16672,N_16639);
and U16895 (N_16895,N_16675,N_16653);
nor U16896 (N_16896,N_16634,N_16715);
xnor U16897 (N_16897,N_16694,N_16522);
and U16898 (N_16898,N_16605,N_16574);
or U16899 (N_16899,N_16511,N_16572);
nor U16900 (N_16900,N_16533,N_16519);
nand U16901 (N_16901,N_16516,N_16693);
nand U16902 (N_16902,N_16531,N_16659);
xnor U16903 (N_16903,N_16544,N_16601);
xor U16904 (N_16904,N_16710,N_16504);
or U16905 (N_16905,N_16714,N_16664);
xnor U16906 (N_16906,N_16610,N_16510);
or U16907 (N_16907,N_16505,N_16537);
nand U16908 (N_16908,N_16658,N_16566);
or U16909 (N_16909,N_16688,N_16580);
xor U16910 (N_16910,N_16549,N_16519);
and U16911 (N_16911,N_16603,N_16563);
nand U16912 (N_16912,N_16603,N_16618);
xnor U16913 (N_16913,N_16658,N_16608);
xor U16914 (N_16914,N_16602,N_16607);
or U16915 (N_16915,N_16689,N_16707);
nand U16916 (N_16916,N_16666,N_16552);
and U16917 (N_16917,N_16624,N_16566);
or U16918 (N_16918,N_16689,N_16535);
nor U16919 (N_16919,N_16680,N_16723);
nor U16920 (N_16920,N_16695,N_16536);
nor U16921 (N_16921,N_16620,N_16642);
or U16922 (N_16922,N_16655,N_16598);
nor U16923 (N_16923,N_16718,N_16552);
xor U16924 (N_16924,N_16577,N_16526);
nor U16925 (N_16925,N_16527,N_16721);
nand U16926 (N_16926,N_16726,N_16516);
xor U16927 (N_16927,N_16526,N_16733);
nand U16928 (N_16928,N_16621,N_16581);
nand U16929 (N_16929,N_16648,N_16736);
nor U16930 (N_16930,N_16578,N_16745);
or U16931 (N_16931,N_16500,N_16530);
xnor U16932 (N_16932,N_16595,N_16727);
nor U16933 (N_16933,N_16716,N_16553);
and U16934 (N_16934,N_16747,N_16543);
nor U16935 (N_16935,N_16640,N_16572);
nand U16936 (N_16936,N_16690,N_16565);
and U16937 (N_16937,N_16717,N_16666);
nand U16938 (N_16938,N_16571,N_16562);
nor U16939 (N_16939,N_16546,N_16536);
and U16940 (N_16940,N_16505,N_16736);
nand U16941 (N_16941,N_16507,N_16584);
nor U16942 (N_16942,N_16646,N_16719);
xor U16943 (N_16943,N_16602,N_16631);
and U16944 (N_16944,N_16672,N_16546);
or U16945 (N_16945,N_16652,N_16580);
nor U16946 (N_16946,N_16637,N_16635);
nor U16947 (N_16947,N_16727,N_16594);
and U16948 (N_16948,N_16677,N_16602);
nand U16949 (N_16949,N_16566,N_16669);
xnor U16950 (N_16950,N_16675,N_16521);
or U16951 (N_16951,N_16723,N_16673);
xnor U16952 (N_16952,N_16605,N_16519);
and U16953 (N_16953,N_16605,N_16716);
or U16954 (N_16954,N_16736,N_16595);
and U16955 (N_16955,N_16545,N_16618);
xor U16956 (N_16956,N_16534,N_16601);
xnor U16957 (N_16957,N_16695,N_16736);
nor U16958 (N_16958,N_16571,N_16719);
and U16959 (N_16959,N_16689,N_16699);
nand U16960 (N_16960,N_16680,N_16659);
or U16961 (N_16961,N_16518,N_16686);
or U16962 (N_16962,N_16667,N_16585);
xnor U16963 (N_16963,N_16672,N_16631);
nor U16964 (N_16964,N_16720,N_16651);
nand U16965 (N_16965,N_16601,N_16549);
xor U16966 (N_16966,N_16581,N_16634);
xor U16967 (N_16967,N_16541,N_16676);
and U16968 (N_16968,N_16581,N_16741);
or U16969 (N_16969,N_16591,N_16530);
or U16970 (N_16970,N_16587,N_16560);
nor U16971 (N_16971,N_16545,N_16512);
or U16972 (N_16972,N_16666,N_16636);
and U16973 (N_16973,N_16559,N_16628);
or U16974 (N_16974,N_16656,N_16742);
nand U16975 (N_16975,N_16510,N_16522);
and U16976 (N_16976,N_16737,N_16564);
nor U16977 (N_16977,N_16660,N_16531);
or U16978 (N_16978,N_16645,N_16510);
and U16979 (N_16979,N_16519,N_16586);
xor U16980 (N_16980,N_16526,N_16713);
and U16981 (N_16981,N_16661,N_16748);
nand U16982 (N_16982,N_16604,N_16625);
and U16983 (N_16983,N_16712,N_16675);
or U16984 (N_16984,N_16543,N_16643);
nor U16985 (N_16985,N_16746,N_16687);
xor U16986 (N_16986,N_16592,N_16670);
and U16987 (N_16987,N_16675,N_16670);
xor U16988 (N_16988,N_16545,N_16678);
nor U16989 (N_16989,N_16522,N_16703);
or U16990 (N_16990,N_16550,N_16563);
xnor U16991 (N_16991,N_16568,N_16697);
xor U16992 (N_16992,N_16521,N_16632);
and U16993 (N_16993,N_16726,N_16549);
nand U16994 (N_16994,N_16625,N_16739);
nor U16995 (N_16995,N_16738,N_16694);
nand U16996 (N_16996,N_16627,N_16721);
nor U16997 (N_16997,N_16743,N_16623);
xnor U16998 (N_16998,N_16513,N_16731);
or U16999 (N_16999,N_16553,N_16513);
and U17000 (N_17000,N_16997,N_16994);
nor U17001 (N_17001,N_16782,N_16796);
xor U17002 (N_17002,N_16902,N_16855);
xor U17003 (N_17003,N_16768,N_16950);
nor U17004 (N_17004,N_16888,N_16995);
nor U17005 (N_17005,N_16928,N_16833);
and U17006 (N_17006,N_16805,N_16750);
and U17007 (N_17007,N_16887,N_16926);
or U17008 (N_17008,N_16906,N_16927);
xor U17009 (N_17009,N_16869,N_16815);
and U17010 (N_17010,N_16765,N_16785);
nor U17011 (N_17011,N_16908,N_16821);
and U17012 (N_17012,N_16968,N_16916);
or U17013 (N_17013,N_16914,N_16947);
xor U17014 (N_17014,N_16996,N_16766);
xor U17015 (N_17015,N_16757,N_16848);
nand U17016 (N_17016,N_16857,N_16783);
nor U17017 (N_17017,N_16779,N_16961);
xor U17018 (N_17018,N_16828,N_16763);
and U17019 (N_17019,N_16784,N_16965);
and U17020 (N_17020,N_16915,N_16764);
or U17021 (N_17021,N_16903,N_16778);
or U17022 (N_17022,N_16963,N_16879);
and U17023 (N_17023,N_16835,N_16889);
and U17024 (N_17024,N_16806,N_16864);
xor U17025 (N_17025,N_16954,N_16880);
and U17026 (N_17026,N_16948,N_16966);
nor U17027 (N_17027,N_16956,N_16911);
nor U17028 (N_17028,N_16972,N_16901);
or U17029 (N_17029,N_16999,N_16890);
and U17030 (N_17030,N_16813,N_16987);
nor U17031 (N_17031,N_16886,N_16992);
nor U17032 (N_17032,N_16893,N_16892);
xnor U17033 (N_17033,N_16852,N_16773);
and U17034 (N_17034,N_16876,N_16851);
xnor U17035 (N_17035,N_16867,N_16881);
or U17036 (N_17036,N_16812,N_16883);
or U17037 (N_17037,N_16817,N_16752);
nand U17038 (N_17038,N_16825,N_16858);
nand U17039 (N_17039,N_16925,N_16967);
nand U17040 (N_17040,N_16811,N_16781);
nor U17041 (N_17041,N_16826,N_16870);
nor U17042 (N_17042,N_16907,N_16933);
xor U17043 (N_17043,N_16841,N_16775);
xnor U17044 (N_17044,N_16866,N_16899);
or U17045 (N_17045,N_16885,N_16850);
or U17046 (N_17046,N_16830,N_16875);
xnor U17047 (N_17047,N_16993,N_16840);
nor U17048 (N_17048,N_16955,N_16756);
or U17049 (N_17049,N_16797,N_16774);
or U17050 (N_17050,N_16860,N_16922);
xor U17051 (N_17051,N_16871,N_16807);
nand U17052 (N_17052,N_16802,N_16753);
nand U17053 (N_17053,N_16896,N_16924);
nand U17054 (N_17054,N_16831,N_16854);
nand U17055 (N_17055,N_16957,N_16787);
and U17056 (N_17056,N_16863,N_16980);
nand U17057 (N_17057,N_16761,N_16904);
nand U17058 (N_17058,N_16873,N_16820);
xnor U17059 (N_17059,N_16845,N_16913);
nand U17060 (N_17060,N_16790,N_16844);
and U17061 (N_17061,N_16794,N_16912);
nand U17062 (N_17062,N_16982,N_16920);
nand U17063 (N_17063,N_16804,N_16829);
xor U17064 (N_17064,N_16984,N_16872);
or U17065 (N_17065,N_16874,N_16940);
or U17066 (N_17066,N_16791,N_16941);
nor U17067 (N_17067,N_16932,N_16960);
and U17068 (N_17068,N_16938,N_16792);
and U17069 (N_17069,N_16979,N_16990);
xnor U17070 (N_17070,N_16777,N_16989);
nand U17071 (N_17071,N_16921,N_16762);
and U17072 (N_17072,N_16978,N_16816);
xnor U17073 (N_17073,N_16898,N_16931);
nor U17074 (N_17074,N_16930,N_16962);
or U17075 (N_17075,N_16843,N_16793);
and U17076 (N_17076,N_16905,N_16918);
nor U17077 (N_17077,N_16936,N_16865);
or U17078 (N_17078,N_16808,N_16949);
nor U17079 (N_17079,N_16975,N_16900);
or U17080 (N_17080,N_16861,N_16929);
xor U17081 (N_17081,N_16799,N_16788);
or U17082 (N_17082,N_16970,N_16877);
xor U17083 (N_17083,N_16770,N_16859);
xnor U17084 (N_17084,N_16942,N_16946);
and U17085 (N_17085,N_16837,N_16827);
xor U17086 (N_17086,N_16758,N_16754);
xor U17087 (N_17087,N_16751,N_16919);
nand U17088 (N_17088,N_16952,N_16839);
or U17089 (N_17089,N_16823,N_16818);
xnor U17090 (N_17090,N_16958,N_16836);
xnor U17091 (N_17091,N_16849,N_16803);
nor U17092 (N_17092,N_16894,N_16944);
xnor U17093 (N_17093,N_16798,N_16973);
xnor U17094 (N_17094,N_16810,N_16759);
nor U17095 (N_17095,N_16834,N_16856);
xnor U17096 (N_17096,N_16800,N_16822);
xor U17097 (N_17097,N_16953,N_16939);
nand U17098 (N_17098,N_16786,N_16769);
and U17099 (N_17099,N_16985,N_16976);
nor U17100 (N_17100,N_16842,N_16923);
and U17101 (N_17101,N_16878,N_16934);
and U17102 (N_17102,N_16772,N_16824);
or U17103 (N_17103,N_16884,N_16776);
xor U17104 (N_17104,N_16838,N_16998);
or U17105 (N_17105,N_16974,N_16951);
or U17106 (N_17106,N_16819,N_16891);
xnor U17107 (N_17107,N_16988,N_16767);
or U17108 (N_17108,N_16977,N_16882);
nor U17109 (N_17109,N_16862,N_16895);
nand U17110 (N_17110,N_16789,N_16943);
nor U17111 (N_17111,N_16780,N_16771);
nand U17112 (N_17112,N_16832,N_16969);
nand U17113 (N_17113,N_16945,N_16986);
nand U17114 (N_17114,N_16809,N_16937);
xnor U17115 (N_17115,N_16935,N_16917);
nand U17116 (N_17116,N_16964,N_16910);
nand U17117 (N_17117,N_16760,N_16983);
nand U17118 (N_17118,N_16868,N_16846);
xor U17119 (N_17119,N_16853,N_16795);
nand U17120 (N_17120,N_16801,N_16909);
and U17121 (N_17121,N_16897,N_16847);
or U17122 (N_17122,N_16959,N_16981);
and U17123 (N_17123,N_16991,N_16971);
and U17124 (N_17124,N_16755,N_16814);
and U17125 (N_17125,N_16981,N_16926);
nor U17126 (N_17126,N_16821,N_16864);
nor U17127 (N_17127,N_16793,N_16831);
nor U17128 (N_17128,N_16789,N_16802);
nor U17129 (N_17129,N_16999,N_16903);
xor U17130 (N_17130,N_16788,N_16867);
and U17131 (N_17131,N_16843,N_16979);
xor U17132 (N_17132,N_16812,N_16942);
and U17133 (N_17133,N_16850,N_16882);
xor U17134 (N_17134,N_16928,N_16785);
or U17135 (N_17135,N_16959,N_16910);
xnor U17136 (N_17136,N_16840,N_16762);
nand U17137 (N_17137,N_16923,N_16954);
and U17138 (N_17138,N_16966,N_16818);
nor U17139 (N_17139,N_16954,N_16876);
and U17140 (N_17140,N_16837,N_16999);
or U17141 (N_17141,N_16752,N_16902);
and U17142 (N_17142,N_16893,N_16771);
xor U17143 (N_17143,N_16855,N_16786);
nor U17144 (N_17144,N_16917,N_16842);
xor U17145 (N_17145,N_16932,N_16855);
xnor U17146 (N_17146,N_16886,N_16760);
nand U17147 (N_17147,N_16901,N_16985);
xnor U17148 (N_17148,N_16884,N_16990);
and U17149 (N_17149,N_16956,N_16883);
xnor U17150 (N_17150,N_16756,N_16762);
and U17151 (N_17151,N_16840,N_16916);
nand U17152 (N_17152,N_16921,N_16816);
or U17153 (N_17153,N_16917,N_16998);
nand U17154 (N_17154,N_16842,N_16763);
nand U17155 (N_17155,N_16938,N_16861);
nand U17156 (N_17156,N_16912,N_16773);
xnor U17157 (N_17157,N_16760,N_16880);
and U17158 (N_17158,N_16905,N_16770);
xor U17159 (N_17159,N_16908,N_16939);
xor U17160 (N_17160,N_16759,N_16807);
and U17161 (N_17161,N_16987,N_16943);
xor U17162 (N_17162,N_16871,N_16979);
nor U17163 (N_17163,N_16787,N_16842);
xor U17164 (N_17164,N_16877,N_16752);
or U17165 (N_17165,N_16946,N_16920);
nor U17166 (N_17166,N_16909,N_16777);
xor U17167 (N_17167,N_16803,N_16867);
nand U17168 (N_17168,N_16989,N_16940);
or U17169 (N_17169,N_16779,N_16967);
or U17170 (N_17170,N_16965,N_16786);
nor U17171 (N_17171,N_16933,N_16889);
or U17172 (N_17172,N_16787,N_16840);
or U17173 (N_17173,N_16770,N_16901);
nand U17174 (N_17174,N_16863,N_16835);
xnor U17175 (N_17175,N_16800,N_16924);
nand U17176 (N_17176,N_16852,N_16938);
and U17177 (N_17177,N_16911,N_16855);
xnor U17178 (N_17178,N_16984,N_16839);
and U17179 (N_17179,N_16954,N_16798);
nand U17180 (N_17180,N_16912,N_16925);
nor U17181 (N_17181,N_16805,N_16936);
and U17182 (N_17182,N_16979,N_16766);
xnor U17183 (N_17183,N_16941,N_16954);
or U17184 (N_17184,N_16772,N_16874);
xnor U17185 (N_17185,N_16969,N_16956);
nand U17186 (N_17186,N_16896,N_16849);
and U17187 (N_17187,N_16969,N_16978);
nand U17188 (N_17188,N_16850,N_16840);
or U17189 (N_17189,N_16866,N_16928);
xnor U17190 (N_17190,N_16954,N_16875);
and U17191 (N_17191,N_16923,N_16913);
nand U17192 (N_17192,N_16894,N_16941);
or U17193 (N_17193,N_16972,N_16877);
or U17194 (N_17194,N_16982,N_16833);
nand U17195 (N_17195,N_16984,N_16865);
xnor U17196 (N_17196,N_16791,N_16956);
nor U17197 (N_17197,N_16790,N_16845);
xnor U17198 (N_17198,N_16794,N_16890);
or U17199 (N_17199,N_16835,N_16966);
nand U17200 (N_17200,N_16770,N_16896);
or U17201 (N_17201,N_16879,N_16997);
or U17202 (N_17202,N_16869,N_16791);
xnor U17203 (N_17203,N_16939,N_16994);
xor U17204 (N_17204,N_16755,N_16895);
or U17205 (N_17205,N_16812,N_16916);
and U17206 (N_17206,N_16896,N_16871);
xnor U17207 (N_17207,N_16953,N_16840);
or U17208 (N_17208,N_16775,N_16876);
or U17209 (N_17209,N_16914,N_16788);
and U17210 (N_17210,N_16786,N_16903);
xor U17211 (N_17211,N_16760,N_16917);
nor U17212 (N_17212,N_16976,N_16873);
xnor U17213 (N_17213,N_16874,N_16925);
xnor U17214 (N_17214,N_16835,N_16796);
or U17215 (N_17215,N_16932,N_16831);
xor U17216 (N_17216,N_16961,N_16757);
xor U17217 (N_17217,N_16870,N_16771);
nor U17218 (N_17218,N_16822,N_16767);
nor U17219 (N_17219,N_16957,N_16808);
or U17220 (N_17220,N_16806,N_16943);
or U17221 (N_17221,N_16798,N_16947);
nand U17222 (N_17222,N_16778,N_16961);
nand U17223 (N_17223,N_16991,N_16900);
xor U17224 (N_17224,N_16840,N_16930);
nor U17225 (N_17225,N_16863,N_16805);
xor U17226 (N_17226,N_16860,N_16792);
nor U17227 (N_17227,N_16752,N_16782);
nand U17228 (N_17228,N_16871,N_16771);
xnor U17229 (N_17229,N_16979,N_16840);
xnor U17230 (N_17230,N_16786,N_16986);
nor U17231 (N_17231,N_16910,N_16756);
xor U17232 (N_17232,N_16943,N_16876);
or U17233 (N_17233,N_16875,N_16750);
or U17234 (N_17234,N_16912,N_16795);
nor U17235 (N_17235,N_16958,N_16760);
xnor U17236 (N_17236,N_16852,N_16984);
and U17237 (N_17237,N_16886,N_16834);
xnor U17238 (N_17238,N_16792,N_16884);
or U17239 (N_17239,N_16780,N_16914);
and U17240 (N_17240,N_16821,N_16800);
nor U17241 (N_17241,N_16782,N_16975);
nor U17242 (N_17242,N_16813,N_16848);
and U17243 (N_17243,N_16824,N_16842);
xor U17244 (N_17244,N_16874,N_16973);
or U17245 (N_17245,N_16813,N_16881);
and U17246 (N_17246,N_16859,N_16943);
xor U17247 (N_17247,N_16926,N_16753);
nand U17248 (N_17248,N_16773,N_16969);
xnor U17249 (N_17249,N_16752,N_16987);
and U17250 (N_17250,N_17128,N_17146);
and U17251 (N_17251,N_17107,N_17061);
nand U17252 (N_17252,N_17007,N_17054);
nand U17253 (N_17253,N_17248,N_17129);
or U17254 (N_17254,N_17177,N_17203);
nand U17255 (N_17255,N_17210,N_17130);
and U17256 (N_17256,N_17197,N_17194);
and U17257 (N_17257,N_17149,N_17168);
nand U17258 (N_17258,N_17069,N_17243);
and U17259 (N_17259,N_17090,N_17086);
or U17260 (N_17260,N_17000,N_17133);
xor U17261 (N_17261,N_17077,N_17124);
xor U17262 (N_17262,N_17122,N_17208);
nor U17263 (N_17263,N_17010,N_17192);
or U17264 (N_17264,N_17118,N_17240);
xor U17265 (N_17265,N_17098,N_17155);
nand U17266 (N_17266,N_17110,N_17187);
or U17267 (N_17267,N_17137,N_17154);
nor U17268 (N_17268,N_17218,N_17042);
or U17269 (N_17269,N_17043,N_17055);
xor U17270 (N_17270,N_17163,N_17142);
or U17271 (N_17271,N_17034,N_17206);
xor U17272 (N_17272,N_17117,N_17028);
xnor U17273 (N_17273,N_17079,N_17231);
xnor U17274 (N_17274,N_17005,N_17171);
and U17275 (N_17275,N_17073,N_17037);
xor U17276 (N_17276,N_17169,N_17032);
nor U17277 (N_17277,N_17062,N_17121);
and U17278 (N_17278,N_17113,N_17224);
and U17279 (N_17279,N_17093,N_17120);
xor U17280 (N_17280,N_17150,N_17023);
nand U17281 (N_17281,N_17068,N_17239);
and U17282 (N_17282,N_17067,N_17012);
nand U17283 (N_17283,N_17095,N_17025);
xor U17284 (N_17284,N_17001,N_17220);
and U17285 (N_17285,N_17108,N_17085);
xor U17286 (N_17286,N_17176,N_17053);
nand U17287 (N_17287,N_17141,N_17204);
or U17288 (N_17288,N_17080,N_17157);
nand U17289 (N_17289,N_17195,N_17213);
and U17290 (N_17290,N_17145,N_17196);
and U17291 (N_17291,N_17106,N_17099);
xor U17292 (N_17292,N_17101,N_17234);
nor U17293 (N_17293,N_17065,N_17139);
xor U17294 (N_17294,N_17017,N_17103);
nand U17295 (N_17295,N_17189,N_17111);
and U17296 (N_17296,N_17071,N_17161);
nand U17297 (N_17297,N_17127,N_17217);
nor U17298 (N_17298,N_17242,N_17215);
nor U17299 (N_17299,N_17074,N_17066);
nor U17300 (N_17300,N_17035,N_17135);
nand U17301 (N_17301,N_17087,N_17207);
nor U17302 (N_17302,N_17094,N_17119);
xnor U17303 (N_17303,N_17013,N_17225);
and U17304 (N_17304,N_17116,N_17249);
nand U17305 (N_17305,N_17076,N_17190);
nor U17306 (N_17306,N_17165,N_17198);
and U17307 (N_17307,N_17202,N_17088);
nand U17308 (N_17308,N_17097,N_17082);
and U17309 (N_17309,N_17112,N_17022);
or U17310 (N_17310,N_17180,N_17148);
and U17311 (N_17311,N_17147,N_17031);
nand U17312 (N_17312,N_17184,N_17235);
xor U17313 (N_17313,N_17200,N_17226);
nor U17314 (N_17314,N_17221,N_17125);
nor U17315 (N_17315,N_17123,N_17051);
xnor U17316 (N_17316,N_17075,N_17105);
xnor U17317 (N_17317,N_17236,N_17030);
xnor U17318 (N_17318,N_17029,N_17078);
or U17319 (N_17319,N_17188,N_17152);
and U17320 (N_17320,N_17050,N_17064);
xor U17321 (N_17321,N_17175,N_17011);
and U17322 (N_17322,N_17179,N_17102);
xor U17323 (N_17323,N_17173,N_17070);
nand U17324 (N_17324,N_17191,N_17167);
nand U17325 (N_17325,N_17092,N_17109);
nand U17326 (N_17326,N_17057,N_17143);
xnor U17327 (N_17327,N_17229,N_17246);
or U17328 (N_17328,N_17199,N_17205);
xnor U17329 (N_17329,N_17056,N_17049);
nand U17330 (N_17330,N_17045,N_17016);
xor U17331 (N_17331,N_17230,N_17084);
nor U17332 (N_17332,N_17212,N_17136);
and U17333 (N_17333,N_17026,N_17048);
nor U17334 (N_17334,N_17044,N_17182);
or U17335 (N_17335,N_17241,N_17027);
and U17336 (N_17336,N_17039,N_17209);
and U17337 (N_17337,N_17134,N_17222);
and U17338 (N_17338,N_17186,N_17052);
and U17339 (N_17339,N_17060,N_17140);
or U17340 (N_17340,N_17096,N_17232);
and U17341 (N_17341,N_17100,N_17104);
or U17342 (N_17342,N_17002,N_17162);
xor U17343 (N_17343,N_17041,N_17009);
or U17344 (N_17344,N_17015,N_17153);
and U17345 (N_17345,N_17201,N_17156);
or U17346 (N_17346,N_17244,N_17238);
nor U17347 (N_17347,N_17083,N_17006);
or U17348 (N_17348,N_17223,N_17247);
and U17349 (N_17349,N_17144,N_17151);
nor U17350 (N_17350,N_17219,N_17164);
xor U17351 (N_17351,N_17183,N_17170);
xor U17352 (N_17352,N_17019,N_17072);
nand U17353 (N_17353,N_17126,N_17214);
and U17354 (N_17354,N_17004,N_17020);
xnor U17355 (N_17355,N_17166,N_17174);
xor U17356 (N_17356,N_17081,N_17193);
or U17357 (N_17357,N_17233,N_17227);
nand U17358 (N_17358,N_17046,N_17058);
nor U17359 (N_17359,N_17040,N_17228);
nand U17360 (N_17360,N_17211,N_17021);
and U17361 (N_17361,N_17138,N_17216);
or U17362 (N_17362,N_17014,N_17158);
nand U17363 (N_17363,N_17018,N_17178);
nor U17364 (N_17364,N_17114,N_17047);
nand U17365 (N_17365,N_17063,N_17185);
and U17366 (N_17366,N_17160,N_17003);
or U17367 (N_17367,N_17089,N_17033);
or U17368 (N_17368,N_17091,N_17131);
nor U17369 (N_17369,N_17008,N_17036);
nor U17370 (N_17370,N_17181,N_17172);
nand U17371 (N_17371,N_17024,N_17237);
nand U17372 (N_17372,N_17132,N_17245);
nand U17373 (N_17373,N_17159,N_17115);
and U17374 (N_17374,N_17059,N_17038);
nor U17375 (N_17375,N_17017,N_17032);
nand U17376 (N_17376,N_17177,N_17078);
nor U17377 (N_17377,N_17034,N_17224);
nand U17378 (N_17378,N_17151,N_17051);
xor U17379 (N_17379,N_17102,N_17220);
xnor U17380 (N_17380,N_17225,N_17157);
xor U17381 (N_17381,N_17144,N_17060);
or U17382 (N_17382,N_17036,N_17230);
xnor U17383 (N_17383,N_17059,N_17236);
and U17384 (N_17384,N_17031,N_17238);
xor U17385 (N_17385,N_17058,N_17031);
and U17386 (N_17386,N_17033,N_17001);
xor U17387 (N_17387,N_17200,N_17047);
xnor U17388 (N_17388,N_17165,N_17095);
and U17389 (N_17389,N_17229,N_17227);
nand U17390 (N_17390,N_17125,N_17178);
nor U17391 (N_17391,N_17215,N_17007);
nor U17392 (N_17392,N_17031,N_17000);
and U17393 (N_17393,N_17207,N_17108);
nand U17394 (N_17394,N_17091,N_17148);
or U17395 (N_17395,N_17044,N_17029);
nand U17396 (N_17396,N_17027,N_17227);
xnor U17397 (N_17397,N_17071,N_17140);
and U17398 (N_17398,N_17106,N_17179);
xor U17399 (N_17399,N_17141,N_17066);
nand U17400 (N_17400,N_17190,N_17179);
nand U17401 (N_17401,N_17026,N_17028);
and U17402 (N_17402,N_17049,N_17109);
nand U17403 (N_17403,N_17153,N_17000);
xnor U17404 (N_17404,N_17070,N_17234);
nor U17405 (N_17405,N_17236,N_17035);
and U17406 (N_17406,N_17159,N_17092);
or U17407 (N_17407,N_17054,N_17031);
and U17408 (N_17408,N_17036,N_17066);
nor U17409 (N_17409,N_17093,N_17075);
nand U17410 (N_17410,N_17093,N_17218);
xor U17411 (N_17411,N_17100,N_17112);
and U17412 (N_17412,N_17241,N_17053);
nand U17413 (N_17413,N_17233,N_17038);
nor U17414 (N_17414,N_17068,N_17083);
and U17415 (N_17415,N_17248,N_17166);
or U17416 (N_17416,N_17200,N_17243);
and U17417 (N_17417,N_17070,N_17036);
nor U17418 (N_17418,N_17057,N_17232);
xnor U17419 (N_17419,N_17188,N_17076);
nand U17420 (N_17420,N_17106,N_17192);
xor U17421 (N_17421,N_17087,N_17082);
xor U17422 (N_17422,N_17083,N_17162);
nor U17423 (N_17423,N_17065,N_17076);
and U17424 (N_17424,N_17093,N_17182);
nand U17425 (N_17425,N_17044,N_17059);
nand U17426 (N_17426,N_17167,N_17247);
and U17427 (N_17427,N_17051,N_17137);
nand U17428 (N_17428,N_17135,N_17066);
nand U17429 (N_17429,N_17075,N_17036);
nand U17430 (N_17430,N_17083,N_17078);
or U17431 (N_17431,N_17050,N_17043);
and U17432 (N_17432,N_17034,N_17099);
nor U17433 (N_17433,N_17150,N_17230);
or U17434 (N_17434,N_17115,N_17066);
nor U17435 (N_17435,N_17035,N_17013);
or U17436 (N_17436,N_17153,N_17175);
or U17437 (N_17437,N_17226,N_17001);
or U17438 (N_17438,N_17144,N_17103);
nand U17439 (N_17439,N_17223,N_17000);
and U17440 (N_17440,N_17148,N_17010);
or U17441 (N_17441,N_17106,N_17162);
xnor U17442 (N_17442,N_17114,N_17142);
and U17443 (N_17443,N_17017,N_17085);
or U17444 (N_17444,N_17170,N_17080);
nand U17445 (N_17445,N_17050,N_17203);
xnor U17446 (N_17446,N_17096,N_17105);
and U17447 (N_17447,N_17194,N_17202);
xnor U17448 (N_17448,N_17215,N_17061);
or U17449 (N_17449,N_17237,N_17218);
xor U17450 (N_17450,N_17184,N_17244);
or U17451 (N_17451,N_17121,N_17036);
and U17452 (N_17452,N_17207,N_17073);
or U17453 (N_17453,N_17221,N_17150);
xnor U17454 (N_17454,N_17011,N_17010);
or U17455 (N_17455,N_17178,N_17052);
nand U17456 (N_17456,N_17229,N_17163);
xnor U17457 (N_17457,N_17037,N_17139);
nand U17458 (N_17458,N_17056,N_17060);
or U17459 (N_17459,N_17201,N_17195);
or U17460 (N_17460,N_17121,N_17238);
and U17461 (N_17461,N_17084,N_17078);
or U17462 (N_17462,N_17166,N_17164);
nand U17463 (N_17463,N_17155,N_17033);
or U17464 (N_17464,N_17185,N_17183);
nand U17465 (N_17465,N_17230,N_17239);
nand U17466 (N_17466,N_17012,N_17153);
nand U17467 (N_17467,N_17240,N_17208);
nand U17468 (N_17468,N_17073,N_17192);
xnor U17469 (N_17469,N_17033,N_17096);
nand U17470 (N_17470,N_17191,N_17020);
nand U17471 (N_17471,N_17077,N_17185);
or U17472 (N_17472,N_17091,N_17157);
nand U17473 (N_17473,N_17136,N_17233);
and U17474 (N_17474,N_17192,N_17117);
nand U17475 (N_17475,N_17019,N_17132);
or U17476 (N_17476,N_17202,N_17074);
and U17477 (N_17477,N_17206,N_17211);
or U17478 (N_17478,N_17203,N_17163);
nor U17479 (N_17479,N_17122,N_17197);
nor U17480 (N_17480,N_17232,N_17173);
xnor U17481 (N_17481,N_17180,N_17113);
nand U17482 (N_17482,N_17103,N_17114);
nand U17483 (N_17483,N_17121,N_17095);
xnor U17484 (N_17484,N_17057,N_17094);
or U17485 (N_17485,N_17171,N_17002);
nand U17486 (N_17486,N_17237,N_17244);
nand U17487 (N_17487,N_17161,N_17085);
and U17488 (N_17488,N_17227,N_17098);
nand U17489 (N_17489,N_17151,N_17145);
and U17490 (N_17490,N_17243,N_17083);
xor U17491 (N_17491,N_17067,N_17126);
or U17492 (N_17492,N_17012,N_17106);
and U17493 (N_17493,N_17030,N_17055);
nor U17494 (N_17494,N_17138,N_17126);
or U17495 (N_17495,N_17061,N_17040);
and U17496 (N_17496,N_17127,N_17132);
xor U17497 (N_17497,N_17133,N_17079);
xor U17498 (N_17498,N_17238,N_17237);
and U17499 (N_17499,N_17100,N_17065);
or U17500 (N_17500,N_17302,N_17389);
or U17501 (N_17501,N_17305,N_17372);
xor U17502 (N_17502,N_17299,N_17361);
and U17503 (N_17503,N_17491,N_17337);
nand U17504 (N_17504,N_17394,N_17366);
xor U17505 (N_17505,N_17396,N_17453);
nand U17506 (N_17506,N_17317,N_17298);
xnor U17507 (N_17507,N_17340,N_17465);
xor U17508 (N_17508,N_17379,N_17376);
xor U17509 (N_17509,N_17280,N_17362);
and U17510 (N_17510,N_17464,N_17275);
or U17511 (N_17511,N_17477,N_17312);
and U17512 (N_17512,N_17296,N_17441);
nand U17513 (N_17513,N_17456,N_17256);
nand U17514 (N_17514,N_17314,N_17463);
xnor U17515 (N_17515,N_17404,N_17494);
or U17516 (N_17516,N_17390,N_17349);
nor U17517 (N_17517,N_17383,N_17402);
or U17518 (N_17518,N_17481,N_17270);
and U17519 (N_17519,N_17455,N_17281);
and U17520 (N_17520,N_17253,N_17313);
nand U17521 (N_17521,N_17346,N_17496);
nand U17522 (N_17522,N_17410,N_17310);
nor U17523 (N_17523,N_17415,N_17287);
and U17524 (N_17524,N_17333,N_17328);
or U17525 (N_17525,N_17325,N_17495);
and U17526 (N_17526,N_17445,N_17487);
xnor U17527 (N_17527,N_17433,N_17454);
nand U17528 (N_17528,N_17263,N_17265);
xnor U17529 (N_17529,N_17493,N_17427);
or U17530 (N_17530,N_17303,N_17420);
and U17531 (N_17531,N_17474,N_17286);
nor U17532 (N_17532,N_17426,N_17371);
nor U17533 (N_17533,N_17315,N_17397);
and U17534 (N_17534,N_17355,N_17339);
and U17535 (N_17535,N_17387,N_17484);
nor U17536 (N_17536,N_17447,N_17452);
nor U17537 (N_17537,N_17352,N_17438);
xnor U17538 (N_17538,N_17407,N_17442);
or U17539 (N_17539,N_17358,N_17262);
xnor U17540 (N_17540,N_17332,N_17359);
nand U17541 (N_17541,N_17272,N_17274);
or U17542 (N_17542,N_17408,N_17327);
or U17543 (N_17543,N_17271,N_17486);
xor U17544 (N_17544,N_17306,N_17468);
and U17545 (N_17545,N_17357,N_17334);
nor U17546 (N_17546,N_17326,N_17444);
nand U17547 (N_17547,N_17472,N_17460);
nor U17548 (N_17548,N_17418,N_17282);
nor U17549 (N_17549,N_17440,N_17375);
nor U17550 (N_17550,N_17335,N_17309);
or U17551 (N_17551,N_17250,N_17266);
or U17552 (N_17552,N_17419,N_17264);
and U17553 (N_17553,N_17300,N_17367);
nand U17554 (N_17554,N_17330,N_17391);
and U17555 (N_17555,N_17351,N_17320);
nand U17556 (N_17556,N_17329,N_17368);
nor U17557 (N_17557,N_17476,N_17319);
nor U17558 (N_17558,N_17382,N_17431);
or U17559 (N_17559,N_17421,N_17437);
xor U17560 (N_17560,N_17388,N_17260);
nor U17561 (N_17561,N_17276,N_17488);
nand U17562 (N_17562,N_17251,N_17373);
and U17563 (N_17563,N_17395,N_17492);
nor U17564 (N_17564,N_17331,N_17428);
or U17565 (N_17565,N_17462,N_17473);
or U17566 (N_17566,N_17301,N_17446);
nand U17567 (N_17567,N_17258,N_17277);
or U17568 (N_17568,N_17273,N_17365);
xor U17569 (N_17569,N_17448,N_17497);
nand U17570 (N_17570,N_17294,N_17451);
and U17571 (N_17571,N_17480,N_17422);
nor U17572 (N_17572,N_17400,N_17405);
xnor U17573 (N_17573,N_17345,N_17307);
nor U17574 (N_17574,N_17416,N_17435);
or U17575 (N_17575,N_17293,N_17254);
or U17576 (N_17576,N_17384,N_17283);
and U17577 (N_17577,N_17342,N_17436);
and U17578 (N_17578,N_17459,N_17311);
and U17579 (N_17579,N_17412,N_17385);
nand U17580 (N_17580,N_17429,N_17316);
and U17581 (N_17581,N_17269,N_17257);
nand U17582 (N_17582,N_17490,N_17353);
xor U17583 (N_17583,N_17469,N_17291);
or U17584 (N_17584,N_17483,N_17414);
or U17585 (N_17585,N_17259,N_17295);
and U17586 (N_17586,N_17409,N_17268);
nand U17587 (N_17587,N_17292,N_17489);
nand U17588 (N_17588,N_17386,N_17439);
xnor U17589 (N_17589,N_17434,N_17369);
nand U17590 (N_17590,N_17343,N_17399);
and U17591 (N_17591,N_17344,N_17354);
and U17592 (N_17592,N_17279,N_17479);
nor U17593 (N_17593,N_17443,N_17261);
nand U17594 (N_17594,N_17363,N_17338);
nand U17595 (N_17595,N_17423,N_17252);
nand U17596 (N_17596,N_17285,N_17392);
xnor U17597 (N_17597,N_17457,N_17485);
and U17598 (N_17598,N_17290,N_17364);
and U17599 (N_17599,N_17466,N_17471);
nor U17600 (N_17600,N_17498,N_17321);
and U17601 (N_17601,N_17360,N_17378);
nor U17602 (N_17602,N_17424,N_17348);
and U17603 (N_17603,N_17380,N_17406);
xor U17604 (N_17604,N_17255,N_17398);
xnor U17605 (N_17605,N_17377,N_17417);
or U17606 (N_17606,N_17336,N_17432);
nand U17607 (N_17607,N_17267,N_17467);
nor U17608 (N_17608,N_17393,N_17323);
or U17609 (N_17609,N_17425,N_17350);
xor U17610 (N_17610,N_17482,N_17430);
or U17611 (N_17611,N_17381,N_17478);
and U17612 (N_17612,N_17413,N_17289);
nor U17613 (N_17613,N_17304,N_17401);
nor U17614 (N_17614,N_17278,N_17318);
nor U17615 (N_17615,N_17324,N_17475);
nand U17616 (N_17616,N_17356,N_17449);
nand U17617 (N_17617,N_17297,N_17461);
xor U17618 (N_17618,N_17284,N_17450);
nand U17619 (N_17619,N_17470,N_17308);
nor U17620 (N_17620,N_17499,N_17288);
or U17621 (N_17621,N_17341,N_17347);
and U17622 (N_17622,N_17374,N_17322);
and U17623 (N_17623,N_17411,N_17403);
and U17624 (N_17624,N_17458,N_17370);
nor U17625 (N_17625,N_17356,N_17305);
nor U17626 (N_17626,N_17315,N_17493);
and U17627 (N_17627,N_17455,N_17261);
or U17628 (N_17628,N_17465,N_17395);
or U17629 (N_17629,N_17460,N_17440);
or U17630 (N_17630,N_17453,N_17487);
or U17631 (N_17631,N_17420,N_17270);
and U17632 (N_17632,N_17301,N_17260);
or U17633 (N_17633,N_17335,N_17261);
or U17634 (N_17634,N_17351,N_17457);
and U17635 (N_17635,N_17277,N_17381);
or U17636 (N_17636,N_17365,N_17386);
and U17637 (N_17637,N_17282,N_17391);
nor U17638 (N_17638,N_17390,N_17418);
nand U17639 (N_17639,N_17458,N_17334);
xor U17640 (N_17640,N_17330,N_17309);
nor U17641 (N_17641,N_17360,N_17475);
and U17642 (N_17642,N_17492,N_17454);
or U17643 (N_17643,N_17469,N_17281);
nand U17644 (N_17644,N_17483,N_17306);
nor U17645 (N_17645,N_17372,N_17367);
nand U17646 (N_17646,N_17432,N_17395);
xnor U17647 (N_17647,N_17493,N_17415);
and U17648 (N_17648,N_17355,N_17396);
nand U17649 (N_17649,N_17271,N_17262);
nand U17650 (N_17650,N_17399,N_17396);
or U17651 (N_17651,N_17408,N_17412);
and U17652 (N_17652,N_17264,N_17346);
nor U17653 (N_17653,N_17419,N_17341);
and U17654 (N_17654,N_17455,N_17429);
and U17655 (N_17655,N_17277,N_17431);
xor U17656 (N_17656,N_17279,N_17366);
xor U17657 (N_17657,N_17477,N_17474);
nand U17658 (N_17658,N_17364,N_17453);
and U17659 (N_17659,N_17445,N_17279);
or U17660 (N_17660,N_17390,N_17338);
nor U17661 (N_17661,N_17372,N_17309);
nor U17662 (N_17662,N_17308,N_17294);
and U17663 (N_17663,N_17478,N_17267);
nor U17664 (N_17664,N_17289,N_17395);
nor U17665 (N_17665,N_17429,N_17344);
and U17666 (N_17666,N_17280,N_17411);
or U17667 (N_17667,N_17447,N_17422);
nand U17668 (N_17668,N_17295,N_17465);
nor U17669 (N_17669,N_17484,N_17400);
xnor U17670 (N_17670,N_17264,N_17460);
nand U17671 (N_17671,N_17437,N_17347);
or U17672 (N_17672,N_17419,N_17403);
xor U17673 (N_17673,N_17275,N_17476);
xor U17674 (N_17674,N_17437,N_17287);
or U17675 (N_17675,N_17334,N_17385);
or U17676 (N_17676,N_17395,N_17490);
xnor U17677 (N_17677,N_17329,N_17423);
nor U17678 (N_17678,N_17493,N_17495);
xnor U17679 (N_17679,N_17357,N_17295);
nand U17680 (N_17680,N_17410,N_17287);
xor U17681 (N_17681,N_17302,N_17285);
or U17682 (N_17682,N_17493,N_17405);
and U17683 (N_17683,N_17436,N_17279);
nand U17684 (N_17684,N_17428,N_17364);
nand U17685 (N_17685,N_17424,N_17318);
xor U17686 (N_17686,N_17393,N_17349);
or U17687 (N_17687,N_17328,N_17338);
and U17688 (N_17688,N_17492,N_17427);
or U17689 (N_17689,N_17491,N_17343);
nor U17690 (N_17690,N_17342,N_17399);
nor U17691 (N_17691,N_17308,N_17495);
nor U17692 (N_17692,N_17358,N_17263);
nand U17693 (N_17693,N_17423,N_17285);
and U17694 (N_17694,N_17472,N_17367);
nand U17695 (N_17695,N_17250,N_17365);
nor U17696 (N_17696,N_17466,N_17439);
nand U17697 (N_17697,N_17443,N_17393);
nor U17698 (N_17698,N_17434,N_17477);
xnor U17699 (N_17699,N_17479,N_17390);
nor U17700 (N_17700,N_17312,N_17369);
and U17701 (N_17701,N_17333,N_17472);
nor U17702 (N_17702,N_17352,N_17334);
xnor U17703 (N_17703,N_17344,N_17473);
and U17704 (N_17704,N_17359,N_17478);
or U17705 (N_17705,N_17379,N_17260);
and U17706 (N_17706,N_17488,N_17345);
or U17707 (N_17707,N_17334,N_17324);
and U17708 (N_17708,N_17297,N_17439);
xor U17709 (N_17709,N_17361,N_17335);
and U17710 (N_17710,N_17477,N_17472);
and U17711 (N_17711,N_17462,N_17254);
or U17712 (N_17712,N_17330,N_17361);
nand U17713 (N_17713,N_17353,N_17448);
nor U17714 (N_17714,N_17270,N_17289);
xnor U17715 (N_17715,N_17488,N_17400);
nand U17716 (N_17716,N_17380,N_17476);
or U17717 (N_17717,N_17372,N_17311);
nor U17718 (N_17718,N_17370,N_17253);
xnor U17719 (N_17719,N_17362,N_17255);
or U17720 (N_17720,N_17483,N_17492);
nor U17721 (N_17721,N_17420,N_17479);
xnor U17722 (N_17722,N_17479,N_17316);
nand U17723 (N_17723,N_17255,N_17471);
nor U17724 (N_17724,N_17273,N_17408);
and U17725 (N_17725,N_17360,N_17496);
xnor U17726 (N_17726,N_17472,N_17361);
nand U17727 (N_17727,N_17477,N_17429);
nor U17728 (N_17728,N_17370,N_17492);
nor U17729 (N_17729,N_17484,N_17398);
or U17730 (N_17730,N_17414,N_17400);
or U17731 (N_17731,N_17357,N_17358);
or U17732 (N_17732,N_17471,N_17483);
and U17733 (N_17733,N_17458,N_17321);
or U17734 (N_17734,N_17365,N_17372);
or U17735 (N_17735,N_17254,N_17332);
nand U17736 (N_17736,N_17311,N_17265);
nor U17737 (N_17737,N_17447,N_17330);
and U17738 (N_17738,N_17423,N_17409);
xor U17739 (N_17739,N_17354,N_17380);
or U17740 (N_17740,N_17295,N_17269);
nor U17741 (N_17741,N_17353,N_17340);
or U17742 (N_17742,N_17280,N_17346);
or U17743 (N_17743,N_17317,N_17274);
nor U17744 (N_17744,N_17378,N_17390);
nand U17745 (N_17745,N_17300,N_17459);
nor U17746 (N_17746,N_17253,N_17382);
or U17747 (N_17747,N_17388,N_17366);
and U17748 (N_17748,N_17396,N_17409);
nor U17749 (N_17749,N_17383,N_17371);
or U17750 (N_17750,N_17539,N_17629);
or U17751 (N_17751,N_17604,N_17668);
xnor U17752 (N_17752,N_17608,N_17601);
xor U17753 (N_17753,N_17639,N_17677);
xor U17754 (N_17754,N_17503,N_17655);
and U17755 (N_17755,N_17674,N_17598);
and U17756 (N_17756,N_17571,N_17660);
and U17757 (N_17757,N_17715,N_17501);
nand U17758 (N_17758,N_17575,N_17510);
and U17759 (N_17759,N_17665,N_17541);
nor U17760 (N_17760,N_17648,N_17726);
nor U17761 (N_17761,N_17675,N_17702);
and U17762 (N_17762,N_17561,N_17500);
and U17763 (N_17763,N_17744,N_17673);
nor U17764 (N_17764,N_17507,N_17512);
nor U17765 (N_17765,N_17664,N_17689);
nor U17766 (N_17766,N_17530,N_17574);
and U17767 (N_17767,N_17667,N_17693);
nor U17768 (N_17768,N_17617,N_17672);
nand U17769 (N_17769,N_17662,N_17526);
nor U17770 (N_17770,N_17505,N_17635);
xor U17771 (N_17771,N_17699,N_17565);
nand U17772 (N_17772,N_17701,N_17698);
nor U17773 (N_17773,N_17594,N_17713);
xor U17774 (N_17774,N_17559,N_17663);
and U17775 (N_17775,N_17552,N_17725);
nand U17776 (N_17776,N_17728,N_17696);
and U17777 (N_17777,N_17700,N_17651);
or U17778 (N_17778,N_17543,N_17716);
xor U17779 (N_17779,N_17599,N_17633);
xor U17780 (N_17780,N_17516,N_17557);
nand U17781 (N_17781,N_17533,N_17636);
or U17782 (N_17782,N_17627,N_17618);
nor U17783 (N_17783,N_17523,N_17641);
and U17784 (N_17784,N_17741,N_17509);
xnor U17785 (N_17785,N_17707,N_17583);
or U17786 (N_17786,N_17563,N_17682);
or U17787 (N_17787,N_17595,N_17647);
xor U17788 (N_17788,N_17580,N_17592);
or U17789 (N_17789,N_17546,N_17721);
nor U17790 (N_17790,N_17537,N_17593);
nand U17791 (N_17791,N_17568,N_17531);
nor U17792 (N_17792,N_17714,N_17517);
and U17793 (N_17793,N_17643,N_17709);
and U17794 (N_17794,N_17745,N_17638);
nand U17795 (N_17795,N_17587,N_17658);
or U17796 (N_17796,N_17558,N_17749);
xnor U17797 (N_17797,N_17661,N_17630);
or U17798 (N_17798,N_17717,N_17506);
nand U17799 (N_17799,N_17562,N_17706);
xnor U17800 (N_17800,N_17632,N_17545);
and U17801 (N_17801,N_17591,N_17746);
nand U17802 (N_17802,N_17534,N_17579);
xnor U17803 (N_17803,N_17740,N_17642);
nand U17804 (N_17804,N_17613,N_17532);
nand U17805 (N_17805,N_17614,N_17600);
xnor U17806 (N_17806,N_17695,N_17504);
nor U17807 (N_17807,N_17747,N_17688);
nand U17808 (N_17808,N_17723,N_17649);
xor U17809 (N_17809,N_17684,N_17722);
or U17810 (N_17810,N_17602,N_17519);
nand U17811 (N_17811,N_17690,N_17739);
xor U17812 (N_17812,N_17584,N_17686);
nand U17813 (N_17813,N_17529,N_17513);
or U17814 (N_17814,N_17590,N_17724);
nor U17815 (N_17815,N_17720,N_17625);
xor U17816 (N_17816,N_17727,N_17634);
and U17817 (N_17817,N_17666,N_17650);
or U17818 (N_17818,N_17524,N_17680);
xor U17819 (N_17819,N_17527,N_17540);
or U17820 (N_17820,N_17576,N_17653);
xor U17821 (N_17821,N_17554,N_17742);
or U17822 (N_17822,N_17581,N_17656);
or U17823 (N_17823,N_17560,N_17681);
and U17824 (N_17824,N_17538,N_17611);
nand U17825 (N_17825,N_17549,N_17678);
nor U17826 (N_17826,N_17588,N_17619);
or U17827 (N_17827,N_17731,N_17697);
and U17828 (N_17828,N_17572,N_17712);
or U17829 (N_17829,N_17573,N_17603);
nand U17830 (N_17830,N_17631,N_17521);
nand U17831 (N_17831,N_17628,N_17518);
xor U17832 (N_17832,N_17582,N_17551);
nand U17833 (N_17833,N_17544,N_17585);
nand U17834 (N_17834,N_17620,N_17743);
nand U17835 (N_17835,N_17586,N_17708);
nor U17836 (N_17836,N_17646,N_17514);
or U17837 (N_17837,N_17606,N_17710);
nand U17838 (N_17838,N_17730,N_17654);
nand U17839 (N_17839,N_17652,N_17624);
nand U17840 (N_17840,N_17567,N_17703);
nand U17841 (N_17841,N_17569,N_17704);
nand U17842 (N_17842,N_17566,N_17548);
xnor U17843 (N_17843,N_17737,N_17685);
xor U17844 (N_17844,N_17607,N_17502);
xor U17845 (N_17845,N_17640,N_17748);
xor U17846 (N_17846,N_17609,N_17615);
xnor U17847 (N_17847,N_17623,N_17637);
nor U17848 (N_17848,N_17657,N_17691);
nor U17849 (N_17849,N_17645,N_17550);
xor U17850 (N_17850,N_17729,N_17616);
nor U17851 (N_17851,N_17553,N_17535);
nand U17852 (N_17852,N_17621,N_17589);
and U17853 (N_17853,N_17671,N_17687);
nand U17854 (N_17854,N_17705,N_17711);
and U17855 (N_17855,N_17556,N_17515);
nor U17856 (N_17856,N_17676,N_17733);
nor U17857 (N_17857,N_17669,N_17732);
and U17858 (N_17858,N_17577,N_17578);
and U17859 (N_17859,N_17570,N_17508);
nand U17860 (N_17860,N_17542,N_17536);
and U17861 (N_17861,N_17547,N_17564);
or U17862 (N_17862,N_17596,N_17735);
nor U17863 (N_17863,N_17520,N_17659);
or U17864 (N_17864,N_17511,N_17683);
and U17865 (N_17865,N_17626,N_17694);
nor U17866 (N_17866,N_17528,N_17605);
nand U17867 (N_17867,N_17734,N_17718);
xor U17868 (N_17868,N_17610,N_17738);
xor U17869 (N_17869,N_17597,N_17670);
and U17870 (N_17870,N_17622,N_17555);
nor U17871 (N_17871,N_17736,N_17612);
nor U17872 (N_17872,N_17692,N_17525);
and U17873 (N_17873,N_17522,N_17679);
or U17874 (N_17874,N_17644,N_17719);
or U17875 (N_17875,N_17612,N_17662);
or U17876 (N_17876,N_17637,N_17609);
or U17877 (N_17877,N_17585,N_17504);
and U17878 (N_17878,N_17631,N_17658);
nor U17879 (N_17879,N_17528,N_17554);
xnor U17880 (N_17880,N_17615,N_17581);
xnor U17881 (N_17881,N_17727,N_17657);
or U17882 (N_17882,N_17603,N_17692);
or U17883 (N_17883,N_17618,N_17664);
nand U17884 (N_17884,N_17612,N_17711);
and U17885 (N_17885,N_17620,N_17584);
nor U17886 (N_17886,N_17734,N_17724);
and U17887 (N_17887,N_17692,N_17517);
and U17888 (N_17888,N_17646,N_17544);
and U17889 (N_17889,N_17640,N_17505);
nor U17890 (N_17890,N_17530,N_17605);
nand U17891 (N_17891,N_17572,N_17552);
nor U17892 (N_17892,N_17545,N_17539);
or U17893 (N_17893,N_17522,N_17716);
nor U17894 (N_17894,N_17536,N_17535);
xor U17895 (N_17895,N_17645,N_17678);
xor U17896 (N_17896,N_17518,N_17684);
nand U17897 (N_17897,N_17718,N_17540);
nand U17898 (N_17898,N_17718,N_17714);
nor U17899 (N_17899,N_17613,N_17554);
nand U17900 (N_17900,N_17725,N_17683);
xor U17901 (N_17901,N_17614,N_17574);
or U17902 (N_17902,N_17730,N_17562);
or U17903 (N_17903,N_17518,N_17560);
or U17904 (N_17904,N_17539,N_17540);
xor U17905 (N_17905,N_17736,N_17662);
nand U17906 (N_17906,N_17716,N_17748);
and U17907 (N_17907,N_17729,N_17694);
nand U17908 (N_17908,N_17658,N_17740);
nor U17909 (N_17909,N_17739,N_17657);
xnor U17910 (N_17910,N_17589,N_17609);
or U17911 (N_17911,N_17657,N_17627);
xor U17912 (N_17912,N_17708,N_17706);
and U17913 (N_17913,N_17571,N_17645);
nand U17914 (N_17914,N_17619,N_17744);
or U17915 (N_17915,N_17663,N_17642);
nor U17916 (N_17916,N_17637,N_17669);
nand U17917 (N_17917,N_17534,N_17740);
or U17918 (N_17918,N_17743,N_17591);
and U17919 (N_17919,N_17510,N_17720);
nand U17920 (N_17920,N_17673,N_17644);
xor U17921 (N_17921,N_17714,N_17544);
nor U17922 (N_17922,N_17745,N_17703);
nand U17923 (N_17923,N_17675,N_17521);
or U17924 (N_17924,N_17697,N_17706);
nand U17925 (N_17925,N_17743,N_17581);
nand U17926 (N_17926,N_17686,N_17673);
and U17927 (N_17927,N_17745,N_17544);
or U17928 (N_17928,N_17581,N_17510);
and U17929 (N_17929,N_17706,N_17634);
nor U17930 (N_17930,N_17643,N_17591);
nor U17931 (N_17931,N_17506,N_17629);
nand U17932 (N_17932,N_17619,N_17675);
and U17933 (N_17933,N_17543,N_17672);
or U17934 (N_17934,N_17580,N_17609);
nand U17935 (N_17935,N_17696,N_17545);
or U17936 (N_17936,N_17573,N_17586);
nand U17937 (N_17937,N_17675,N_17641);
and U17938 (N_17938,N_17685,N_17518);
nor U17939 (N_17939,N_17736,N_17651);
or U17940 (N_17940,N_17529,N_17510);
nand U17941 (N_17941,N_17664,N_17625);
xnor U17942 (N_17942,N_17511,N_17659);
nor U17943 (N_17943,N_17530,N_17599);
nand U17944 (N_17944,N_17747,N_17534);
xnor U17945 (N_17945,N_17673,N_17608);
xor U17946 (N_17946,N_17505,N_17628);
nor U17947 (N_17947,N_17694,N_17543);
and U17948 (N_17948,N_17524,N_17516);
xnor U17949 (N_17949,N_17574,N_17737);
and U17950 (N_17950,N_17622,N_17668);
and U17951 (N_17951,N_17518,N_17584);
or U17952 (N_17952,N_17637,N_17746);
nor U17953 (N_17953,N_17547,N_17673);
or U17954 (N_17954,N_17720,N_17661);
or U17955 (N_17955,N_17529,N_17709);
or U17956 (N_17956,N_17610,N_17508);
nor U17957 (N_17957,N_17715,N_17679);
or U17958 (N_17958,N_17564,N_17590);
nor U17959 (N_17959,N_17635,N_17708);
nor U17960 (N_17960,N_17668,N_17679);
nor U17961 (N_17961,N_17732,N_17690);
and U17962 (N_17962,N_17521,N_17564);
nand U17963 (N_17963,N_17700,N_17717);
xor U17964 (N_17964,N_17705,N_17683);
nor U17965 (N_17965,N_17518,N_17619);
nor U17966 (N_17966,N_17533,N_17558);
xor U17967 (N_17967,N_17564,N_17660);
and U17968 (N_17968,N_17621,N_17659);
xnor U17969 (N_17969,N_17716,N_17541);
nand U17970 (N_17970,N_17576,N_17616);
and U17971 (N_17971,N_17722,N_17547);
and U17972 (N_17972,N_17529,N_17693);
xnor U17973 (N_17973,N_17554,N_17515);
xor U17974 (N_17974,N_17552,N_17637);
nand U17975 (N_17975,N_17608,N_17605);
or U17976 (N_17976,N_17587,N_17586);
and U17977 (N_17977,N_17614,N_17737);
and U17978 (N_17978,N_17638,N_17646);
nand U17979 (N_17979,N_17563,N_17734);
nor U17980 (N_17980,N_17526,N_17610);
nand U17981 (N_17981,N_17510,N_17676);
nand U17982 (N_17982,N_17674,N_17629);
nand U17983 (N_17983,N_17634,N_17542);
nor U17984 (N_17984,N_17606,N_17692);
nand U17985 (N_17985,N_17555,N_17700);
nor U17986 (N_17986,N_17684,N_17620);
nor U17987 (N_17987,N_17658,N_17532);
nand U17988 (N_17988,N_17716,N_17562);
xnor U17989 (N_17989,N_17590,N_17742);
or U17990 (N_17990,N_17690,N_17623);
and U17991 (N_17991,N_17546,N_17511);
nor U17992 (N_17992,N_17507,N_17574);
and U17993 (N_17993,N_17562,N_17666);
xor U17994 (N_17994,N_17610,N_17574);
and U17995 (N_17995,N_17727,N_17596);
nand U17996 (N_17996,N_17680,N_17507);
xor U17997 (N_17997,N_17506,N_17708);
xnor U17998 (N_17998,N_17598,N_17581);
nor U17999 (N_17999,N_17578,N_17736);
and U18000 (N_18000,N_17756,N_17813);
nor U18001 (N_18001,N_17934,N_17942);
or U18002 (N_18002,N_17783,N_17818);
and U18003 (N_18003,N_17795,N_17950);
xnor U18004 (N_18004,N_17765,N_17963);
xnor U18005 (N_18005,N_17954,N_17949);
nor U18006 (N_18006,N_17951,N_17830);
nand U18007 (N_18007,N_17993,N_17973);
and U18008 (N_18008,N_17866,N_17788);
nor U18009 (N_18009,N_17930,N_17971);
xnor U18010 (N_18010,N_17764,N_17856);
or U18011 (N_18011,N_17956,N_17944);
and U18012 (N_18012,N_17986,N_17787);
nor U18013 (N_18013,N_17881,N_17769);
and U18014 (N_18014,N_17924,N_17885);
or U18015 (N_18015,N_17774,N_17964);
or U18016 (N_18016,N_17758,N_17903);
xnor U18017 (N_18017,N_17894,N_17911);
xnor U18018 (N_18018,N_17821,N_17947);
nor U18019 (N_18019,N_17895,N_17864);
nor U18020 (N_18020,N_17886,N_17915);
and U18021 (N_18021,N_17896,N_17862);
nor U18022 (N_18022,N_17920,N_17926);
or U18023 (N_18023,N_17958,N_17803);
and U18024 (N_18024,N_17848,N_17790);
nor U18025 (N_18025,N_17806,N_17962);
or U18026 (N_18026,N_17922,N_17876);
nor U18027 (N_18027,N_17857,N_17804);
or U18028 (N_18028,N_17763,N_17939);
xor U18029 (N_18029,N_17861,N_17770);
or U18030 (N_18030,N_17840,N_17796);
or U18031 (N_18031,N_17843,N_17981);
nor U18032 (N_18032,N_17967,N_17780);
and U18033 (N_18033,N_17900,N_17837);
and U18034 (N_18034,N_17997,N_17928);
or U18035 (N_18035,N_17781,N_17753);
xnor U18036 (N_18036,N_17898,N_17937);
nor U18037 (N_18037,N_17999,N_17952);
xor U18038 (N_18038,N_17878,N_17799);
xnor U18039 (N_18039,N_17815,N_17771);
nand U18040 (N_18040,N_17792,N_17853);
nor U18041 (N_18041,N_17912,N_17929);
and U18042 (N_18042,N_17890,N_17871);
and U18043 (N_18043,N_17811,N_17814);
nand U18044 (N_18044,N_17976,N_17849);
and U18045 (N_18045,N_17933,N_17851);
or U18046 (N_18046,N_17831,N_17940);
and U18047 (N_18047,N_17972,N_17945);
nor U18048 (N_18048,N_17984,N_17836);
and U18049 (N_18049,N_17784,N_17782);
nand U18050 (N_18050,N_17902,N_17936);
or U18051 (N_18051,N_17983,N_17957);
xor U18052 (N_18052,N_17778,N_17880);
and U18053 (N_18053,N_17819,N_17916);
and U18054 (N_18054,N_17935,N_17845);
or U18055 (N_18055,N_17988,N_17991);
nor U18056 (N_18056,N_17833,N_17948);
or U18057 (N_18057,N_17752,N_17820);
xnor U18058 (N_18058,N_17875,N_17827);
xor U18059 (N_18059,N_17750,N_17828);
xnor U18060 (N_18060,N_17918,N_17809);
or U18061 (N_18061,N_17860,N_17858);
nand U18062 (N_18062,N_17882,N_17767);
nor U18063 (N_18063,N_17893,N_17901);
or U18064 (N_18064,N_17990,N_17887);
nand U18065 (N_18065,N_17970,N_17965);
nand U18066 (N_18066,N_17982,N_17798);
xor U18067 (N_18067,N_17992,N_17874);
xor U18068 (N_18068,N_17977,N_17995);
xnor U18069 (N_18069,N_17805,N_17969);
xor U18070 (N_18070,N_17888,N_17835);
xnor U18071 (N_18071,N_17966,N_17847);
nor U18072 (N_18072,N_17816,N_17850);
or U18073 (N_18073,N_17834,N_17807);
xnor U18074 (N_18074,N_17877,N_17914);
nor U18075 (N_18075,N_17846,N_17777);
or U18076 (N_18076,N_17960,N_17927);
and U18077 (N_18077,N_17953,N_17852);
xor U18078 (N_18078,N_17824,N_17772);
and U18079 (N_18079,N_17842,N_17791);
nand U18080 (N_18080,N_17823,N_17909);
nand U18081 (N_18081,N_17808,N_17946);
nor U18082 (N_18082,N_17844,N_17923);
nor U18083 (N_18083,N_17863,N_17921);
or U18084 (N_18084,N_17961,N_17906);
nor U18085 (N_18085,N_17959,N_17768);
or U18086 (N_18086,N_17829,N_17755);
nand U18087 (N_18087,N_17872,N_17985);
or U18088 (N_18088,N_17838,N_17802);
or U18089 (N_18089,N_17955,N_17817);
nor U18090 (N_18090,N_17757,N_17913);
nor U18091 (N_18091,N_17800,N_17996);
nand U18092 (N_18092,N_17868,N_17975);
nand U18093 (N_18093,N_17883,N_17775);
or U18094 (N_18094,N_17812,N_17907);
xor U18095 (N_18095,N_17841,N_17785);
or U18096 (N_18096,N_17839,N_17978);
nand U18097 (N_18097,N_17751,N_17826);
xnor U18098 (N_18098,N_17794,N_17797);
and U18099 (N_18099,N_17980,N_17889);
nor U18100 (N_18100,N_17766,N_17899);
nand U18101 (N_18101,N_17793,N_17989);
nand U18102 (N_18102,N_17905,N_17832);
nand U18103 (N_18103,N_17859,N_17910);
and U18104 (N_18104,N_17987,N_17867);
xnor U18105 (N_18105,N_17760,N_17779);
nor U18106 (N_18106,N_17925,N_17759);
nand U18107 (N_18107,N_17801,N_17776);
nor U18108 (N_18108,N_17979,N_17968);
nand U18109 (N_18109,N_17938,N_17891);
xor U18110 (N_18110,N_17897,N_17789);
and U18111 (N_18111,N_17998,N_17932);
nor U18112 (N_18112,N_17941,N_17908);
and U18113 (N_18113,N_17919,N_17854);
and U18114 (N_18114,N_17754,N_17822);
nand U18115 (N_18115,N_17879,N_17892);
xnor U18116 (N_18116,N_17884,N_17869);
xor U18117 (N_18117,N_17773,N_17904);
nand U18118 (N_18118,N_17786,N_17917);
nor U18119 (N_18119,N_17855,N_17974);
or U18120 (N_18120,N_17762,N_17865);
nor U18121 (N_18121,N_17810,N_17825);
and U18122 (N_18122,N_17994,N_17873);
nor U18123 (N_18123,N_17943,N_17931);
nor U18124 (N_18124,N_17761,N_17870);
nand U18125 (N_18125,N_17764,N_17754);
nand U18126 (N_18126,N_17926,N_17931);
xnor U18127 (N_18127,N_17752,N_17958);
nor U18128 (N_18128,N_17758,N_17980);
nor U18129 (N_18129,N_17916,N_17781);
and U18130 (N_18130,N_17769,N_17898);
or U18131 (N_18131,N_17886,N_17899);
or U18132 (N_18132,N_17798,N_17796);
nor U18133 (N_18133,N_17954,N_17806);
nand U18134 (N_18134,N_17955,N_17755);
nor U18135 (N_18135,N_17779,N_17950);
or U18136 (N_18136,N_17754,N_17882);
nor U18137 (N_18137,N_17936,N_17756);
xnor U18138 (N_18138,N_17849,N_17887);
nor U18139 (N_18139,N_17988,N_17753);
and U18140 (N_18140,N_17889,N_17814);
nor U18141 (N_18141,N_17869,N_17753);
nand U18142 (N_18142,N_17864,N_17946);
xnor U18143 (N_18143,N_17924,N_17825);
xnor U18144 (N_18144,N_17755,N_17882);
nand U18145 (N_18145,N_17980,N_17893);
nand U18146 (N_18146,N_17816,N_17751);
and U18147 (N_18147,N_17999,N_17757);
nand U18148 (N_18148,N_17861,N_17989);
or U18149 (N_18149,N_17921,N_17857);
nand U18150 (N_18150,N_17894,N_17902);
and U18151 (N_18151,N_17807,N_17775);
xor U18152 (N_18152,N_17932,N_17777);
or U18153 (N_18153,N_17904,N_17866);
xor U18154 (N_18154,N_17787,N_17940);
xor U18155 (N_18155,N_17867,N_17784);
xor U18156 (N_18156,N_17863,N_17798);
nand U18157 (N_18157,N_17948,N_17983);
and U18158 (N_18158,N_17796,N_17948);
or U18159 (N_18159,N_17877,N_17860);
xor U18160 (N_18160,N_17792,N_17867);
nor U18161 (N_18161,N_17772,N_17947);
xor U18162 (N_18162,N_17911,N_17758);
or U18163 (N_18163,N_17887,N_17932);
xnor U18164 (N_18164,N_17957,N_17962);
nor U18165 (N_18165,N_17903,N_17948);
nand U18166 (N_18166,N_17813,N_17854);
nand U18167 (N_18167,N_17880,N_17970);
nor U18168 (N_18168,N_17839,N_17921);
xnor U18169 (N_18169,N_17847,N_17995);
xnor U18170 (N_18170,N_17998,N_17965);
or U18171 (N_18171,N_17891,N_17960);
nand U18172 (N_18172,N_17772,N_17781);
nor U18173 (N_18173,N_17760,N_17781);
nand U18174 (N_18174,N_17757,N_17796);
nor U18175 (N_18175,N_17923,N_17895);
nand U18176 (N_18176,N_17752,N_17888);
or U18177 (N_18177,N_17844,N_17800);
nand U18178 (N_18178,N_17757,N_17968);
nand U18179 (N_18179,N_17943,N_17887);
and U18180 (N_18180,N_17807,N_17808);
or U18181 (N_18181,N_17754,N_17770);
or U18182 (N_18182,N_17956,N_17990);
nor U18183 (N_18183,N_17838,N_17971);
nor U18184 (N_18184,N_17892,N_17826);
or U18185 (N_18185,N_17885,N_17803);
and U18186 (N_18186,N_17938,N_17777);
or U18187 (N_18187,N_17840,N_17916);
xor U18188 (N_18188,N_17777,N_17982);
or U18189 (N_18189,N_17832,N_17862);
and U18190 (N_18190,N_17892,N_17847);
xnor U18191 (N_18191,N_17820,N_17960);
nor U18192 (N_18192,N_17945,N_17953);
nand U18193 (N_18193,N_17819,N_17758);
nor U18194 (N_18194,N_17898,N_17968);
nor U18195 (N_18195,N_17971,N_17804);
xor U18196 (N_18196,N_17795,N_17943);
nor U18197 (N_18197,N_17852,N_17888);
nand U18198 (N_18198,N_17789,N_17800);
xnor U18199 (N_18199,N_17999,N_17941);
nand U18200 (N_18200,N_17752,N_17886);
xor U18201 (N_18201,N_17852,N_17797);
xor U18202 (N_18202,N_17818,N_17985);
nand U18203 (N_18203,N_17757,N_17961);
xor U18204 (N_18204,N_17937,N_17835);
nor U18205 (N_18205,N_17767,N_17890);
nand U18206 (N_18206,N_17971,N_17954);
and U18207 (N_18207,N_17796,N_17993);
nor U18208 (N_18208,N_17996,N_17892);
nand U18209 (N_18209,N_17998,N_17979);
or U18210 (N_18210,N_17925,N_17999);
and U18211 (N_18211,N_17823,N_17953);
xnor U18212 (N_18212,N_17810,N_17968);
nand U18213 (N_18213,N_17804,N_17979);
nand U18214 (N_18214,N_17772,N_17786);
xnor U18215 (N_18215,N_17875,N_17866);
nor U18216 (N_18216,N_17980,N_17858);
nand U18217 (N_18217,N_17768,N_17802);
nand U18218 (N_18218,N_17753,N_17862);
xor U18219 (N_18219,N_17839,N_17946);
or U18220 (N_18220,N_17935,N_17966);
xor U18221 (N_18221,N_17939,N_17827);
xnor U18222 (N_18222,N_17968,N_17750);
xnor U18223 (N_18223,N_17759,N_17889);
xor U18224 (N_18224,N_17811,N_17930);
xnor U18225 (N_18225,N_17794,N_17944);
or U18226 (N_18226,N_17847,N_17777);
nor U18227 (N_18227,N_17992,N_17941);
nand U18228 (N_18228,N_17861,N_17755);
or U18229 (N_18229,N_17868,N_17793);
nand U18230 (N_18230,N_17818,N_17943);
or U18231 (N_18231,N_17968,N_17792);
nand U18232 (N_18232,N_17813,N_17871);
nor U18233 (N_18233,N_17789,N_17862);
nand U18234 (N_18234,N_17868,N_17781);
nor U18235 (N_18235,N_17831,N_17776);
nand U18236 (N_18236,N_17950,N_17926);
xor U18237 (N_18237,N_17970,N_17848);
and U18238 (N_18238,N_17998,N_17783);
nor U18239 (N_18239,N_17811,N_17962);
and U18240 (N_18240,N_17927,N_17989);
and U18241 (N_18241,N_17794,N_17996);
nand U18242 (N_18242,N_17879,N_17931);
nor U18243 (N_18243,N_17826,N_17797);
and U18244 (N_18244,N_17764,N_17767);
and U18245 (N_18245,N_17811,N_17792);
nor U18246 (N_18246,N_17837,N_17854);
or U18247 (N_18247,N_17880,N_17753);
or U18248 (N_18248,N_17809,N_17995);
xnor U18249 (N_18249,N_17958,N_17956);
xnor U18250 (N_18250,N_18132,N_18182);
xor U18251 (N_18251,N_18143,N_18010);
nor U18252 (N_18252,N_18111,N_18229);
xor U18253 (N_18253,N_18030,N_18233);
nor U18254 (N_18254,N_18057,N_18139);
or U18255 (N_18255,N_18045,N_18065);
or U18256 (N_18256,N_18008,N_18246);
nor U18257 (N_18257,N_18091,N_18096);
nor U18258 (N_18258,N_18101,N_18079);
xor U18259 (N_18259,N_18037,N_18009);
or U18260 (N_18260,N_18038,N_18196);
nand U18261 (N_18261,N_18136,N_18003);
nor U18262 (N_18262,N_18085,N_18201);
xnor U18263 (N_18263,N_18095,N_18186);
or U18264 (N_18264,N_18148,N_18142);
nand U18265 (N_18265,N_18108,N_18115);
xnor U18266 (N_18266,N_18058,N_18248);
xor U18267 (N_18267,N_18200,N_18176);
nor U18268 (N_18268,N_18192,N_18018);
xor U18269 (N_18269,N_18056,N_18088);
nand U18270 (N_18270,N_18226,N_18247);
and U18271 (N_18271,N_18110,N_18249);
xnor U18272 (N_18272,N_18118,N_18125);
and U18273 (N_18273,N_18100,N_18144);
nor U18274 (N_18274,N_18087,N_18166);
nor U18275 (N_18275,N_18209,N_18205);
and U18276 (N_18276,N_18178,N_18163);
or U18277 (N_18277,N_18202,N_18235);
or U18278 (N_18278,N_18214,N_18075);
xor U18279 (N_18279,N_18134,N_18116);
nand U18280 (N_18280,N_18208,N_18083);
xnor U18281 (N_18281,N_18044,N_18011);
xor U18282 (N_18282,N_18150,N_18103);
nand U18283 (N_18283,N_18033,N_18160);
xnor U18284 (N_18284,N_18162,N_18106);
nor U18285 (N_18285,N_18099,N_18220);
nand U18286 (N_18286,N_18180,N_18019);
nor U18287 (N_18287,N_18123,N_18028);
and U18288 (N_18288,N_18133,N_18051);
nor U18289 (N_18289,N_18173,N_18197);
xnor U18290 (N_18290,N_18046,N_18135);
nand U18291 (N_18291,N_18047,N_18076);
xnor U18292 (N_18292,N_18232,N_18187);
nor U18293 (N_18293,N_18069,N_18219);
nand U18294 (N_18294,N_18024,N_18241);
nand U18295 (N_18295,N_18114,N_18107);
nor U18296 (N_18296,N_18161,N_18002);
nand U18297 (N_18297,N_18199,N_18021);
nand U18298 (N_18298,N_18090,N_18014);
nor U18299 (N_18299,N_18013,N_18244);
xnor U18300 (N_18300,N_18032,N_18195);
and U18301 (N_18301,N_18126,N_18112);
and U18302 (N_18302,N_18077,N_18155);
nand U18303 (N_18303,N_18181,N_18210);
xnor U18304 (N_18304,N_18080,N_18198);
nand U18305 (N_18305,N_18119,N_18140);
nand U18306 (N_18306,N_18170,N_18104);
or U18307 (N_18307,N_18221,N_18015);
nor U18308 (N_18308,N_18147,N_18122);
nand U18309 (N_18309,N_18225,N_18190);
and U18310 (N_18310,N_18042,N_18102);
nand U18311 (N_18311,N_18053,N_18179);
xor U18312 (N_18312,N_18152,N_18184);
and U18313 (N_18313,N_18059,N_18218);
or U18314 (N_18314,N_18191,N_18138);
or U18315 (N_18315,N_18245,N_18060);
or U18316 (N_18316,N_18070,N_18129);
nor U18317 (N_18317,N_18213,N_18041);
nor U18318 (N_18318,N_18092,N_18023);
nor U18319 (N_18319,N_18215,N_18239);
nand U18320 (N_18320,N_18223,N_18063);
nand U18321 (N_18321,N_18212,N_18005);
nor U18322 (N_18322,N_18066,N_18216);
or U18323 (N_18323,N_18081,N_18130);
nor U18324 (N_18324,N_18031,N_18149);
and U18325 (N_18325,N_18206,N_18204);
or U18326 (N_18326,N_18211,N_18203);
nor U18327 (N_18327,N_18049,N_18084);
xnor U18328 (N_18328,N_18078,N_18169);
nor U18329 (N_18329,N_18194,N_18228);
xor U18330 (N_18330,N_18012,N_18240);
or U18331 (N_18331,N_18074,N_18141);
and U18332 (N_18332,N_18124,N_18109);
xnor U18333 (N_18333,N_18000,N_18004);
nor U18334 (N_18334,N_18222,N_18230);
xnor U18335 (N_18335,N_18036,N_18167);
or U18336 (N_18336,N_18043,N_18153);
and U18337 (N_18337,N_18025,N_18029);
and U18338 (N_18338,N_18097,N_18050);
xnor U18339 (N_18339,N_18175,N_18017);
and U18340 (N_18340,N_18242,N_18188);
nor U18341 (N_18341,N_18237,N_18128);
nor U18342 (N_18342,N_18082,N_18022);
and U18343 (N_18343,N_18131,N_18243);
xor U18344 (N_18344,N_18027,N_18062);
xor U18345 (N_18345,N_18193,N_18064);
or U18346 (N_18346,N_18052,N_18113);
xnor U18347 (N_18347,N_18217,N_18156);
nand U18348 (N_18348,N_18183,N_18068);
nand U18349 (N_18349,N_18054,N_18236);
and U18350 (N_18350,N_18157,N_18067);
xor U18351 (N_18351,N_18174,N_18185);
or U18352 (N_18352,N_18145,N_18146);
and U18353 (N_18353,N_18073,N_18168);
nand U18354 (N_18354,N_18089,N_18120);
nor U18355 (N_18355,N_18159,N_18171);
nor U18356 (N_18356,N_18035,N_18117);
or U18357 (N_18357,N_18039,N_18151);
nand U18358 (N_18358,N_18224,N_18098);
nand U18359 (N_18359,N_18172,N_18238);
and U18360 (N_18360,N_18105,N_18207);
nand U18361 (N_18361,N_18061,N_18137);
nor U18362 (N_18362,N_18086,N_18154);
nand U18363 (N_18363,N_18164,N_18016);
or U18364 (N_18364,N_18072,N_18094);
xnor U18365 (N_18365,N_18234,N_18231);
nand U18366 (N_18366,N_18006,N_18026);
xor U18367 (N_18367,N_18127,N_18121);
or U18368 (N_18368,N_18020,N_18227);
nand U18369 (N_18369,N_18189,N_18040);
nand U18370 (N_18370,N_18007,N_18055);
nor U18371 (N_18371,N_18165,N_18034);
or U18372 (N_18372,N_18048,N_18001);
xor U18373 (N_18373,N_18071,N_18158);
nand U18374 (N_18374,N_18177,N_18093);
or U18375 (N_18375,N_18177,N_18112);
nor U18376 (N_18376,N_18091,N_18158);
and U18377 (N_18377,N_18096,N_18085);
nor U18378 (N_18378,N_18246,N_18103);
nor U18379 (N_18379,N_18142,N_18067);
xnor U18380 (N_18380,N_18249,N_18173);
and U18381 (N_18381,N_18218,N_18190);
and U18382 (N_18382,N_18000,N_18192);
nor U18383 (N_18383,N_18205,N_18218);
nand U18384 (N_18384,N_18139,N_18105);
and U18385 (N_18385,N_18016,N_18202);
and U18386 (N_18386,N_18219,N_18222);
xor U18387 (N_18387,N_18077,N_18202);
xor U18388 (N_18388,N_18036,N_18198);
nand U18389 (N_18389,N_18243,N_18177);
nor U18390 (N_18390,N_18041,N_18177);
nor U18391 (N_18391,N_18016,N_18220);
or U18392 (N_18392,N_18057,N_18026);
and U18393 (N_18393,N_18170,N_18160);
nand U18394 (N_18394,N_18156,N_18141);
or U18395 (N_18395,N_18037,N_18050);
nand U18396 (N_18396,N_18184,N_18113);
nand U18397 (N_18397,N_18110,N_18150);
nand U18398 (N_18398,N_18075,N_18016);
nor U18399 (N_18399,N_18099,N_18182);
xor U18400 (N_18400,N_18178,N_18025);
xnor U18401 (N_18401,N_18058,N_18187);
and U18402 (N_18402,N_18212,N_18229);
or U18403 (N_18403,N_18013,N_18084);
xnor U18404 (N_18404,N_18153,N_18242);
xor U18405 (N_18405,N_18097,N_18153);
xor U18406 (N_18406,N_18182,N_18086);
xor U18407 (N_18407,N_18003,N_18208);
and U18408 (N_18408,N_18094,N_18116);
nand U18409 (N_18409,N_18012,N_18079);
or U18410 (N_18410,N_18166,N_18019);
xor U18411 (N_18411,N_18032,N_18140);
and U18412 (N_18412,N_18066,N_18085);
xor U18413 (N_18413,N_18132,N_18019);
nor U18414 (N_18414,N_18116,N_18101);
or U18415 (N_18415,N_18082,N_18120);
xnor U18416 (N_18416,N_18248,N_18005);
xnor U18417 (N_18417,N_18189,N_18216);
nand U18418 (N_18418,N_18238,N_18041);
nand U18419 (N_18419,N_18178,N_18071);
and U18420 (N_18420,N_18171,N_18055);
xnor U18421 (N_18421,N_18175,N_18004);
or U18422 (N_18422,N_18245,N_18106);
nor U18423 (N_18423,N_18238,N_18054);
nand U18424 (N_18424,N_18210,N_18071);
and U18425 (N_18425,N_18041,N_18131);
nor U18426 (N_18426,N_18213,N_18150);
and U18427 (N_18427,N_18147,N_18243);
xnor U18428 (N_18428,N_18021,N_18085);
nor U18429 (N_18429,N_18099,N_18168);
nor U18430 (N_18430,N_18134,N_18050);
or U18431 (N_18431,N_18029,N_18057);
xnor U18432 (N_18432,N_18195,N_18213);
xnor U18433 (N_18433,N_18181,N_18162);
xor U18434 (N_18434,N_18129,N_18198);
or U18435 (N_18435,N_18073,N_18139);
and U18436 (N_18436,N_18165,N_18010);
xor U18437 (N_18437,N_18153,N_18205);
nor U18438 (N_18438,N_18202,N_18080);
nor U18439 (N_18439,N_18234,N_18246);
nor U18440 (N_18440,N_18210,N_18152);
or U18441 (N_18441,N_18044,N_18049);
nor U18442 (N_18442,N_18049,N_18087);
and U18443 (N_18443,N_18189,N_18211);
and U18444 (N_18444,N_18123,N_18131);
or U18445 (N_18445,N_18174,N_18151);
nor U18446 (N_18446,N_18017,N_18173);
nand U18447 (N_18447,N_18204,N_18070);
nand U18448 (N_18448,N_18207,N_18004);
and U18449 (N_18449,N_18075,N_18027);
xnor U18450 (N_18450,N_18046,N_18197);
nand U18451 (N_18451,N_18009,N_18181);
nand U18452 (N_18452,N_18188,N_18130);
xor U18453 (N_18453,N_18123,N_18055);
nor U18454 (N_18454,N_18150,N_18012);
nor U18455 (N_18455,N_18210,N_18078);
and U18456 (N_18456,N_18014,N_18221);
or U18457 (N_18457,N_18020,N_18052);
or U18458 (N_18458,N_18087,N_18085);
xnor U18459 (N_18459,N_18051,N_18240);
nand U18460 (N_18460,N_18217,N_18051);
nand U18461 (N_18461,N_18171,N_18033);
or U18462 (N_18462,N_18207,N_18058);
nand U18463 (N_18463,N_18120,N_18008);
nor U18464 (N_18464,N_18034,N_18000);
and U18465 (N_18465,N_18103,N_18181);
xnor U18466 (N_18466,N_18098,N_18206);
nor U18467 (N_18467,N_18078,N_18244);
nor U18468 (N_18468,N_18183,N_18222);
xnor U18469 (N_18469,N_18043,N_18034);
or U18470 (N_18470,N_18026,N_18089);
nand U18471 (N_18471,N_18013,N_18193);
and U18472 (N_18472,N_18084,N_18032);
nor U18473 (N_18473,N_18129,N_18017);
nand U18474 (N_18474,N_18120,N_18019);
nand U18475 (N_18475,N_18188,N_18038);
xor U18476 (N_18476,N_18184,N_18234);
nor U18477 (N_18477,N_18058,N_18090);
xnor U18478 (N_18478,N_18154,N_18142);
or U18479 (N_18479,N_18167,N_18054);
and U18480 (N_18480,N_18101,N_18210);
nand U18481 (N_18481,N_18180,N_18002);
or U18482 (N_18482,N_18122,N_18096);
nand U18483 (N_18483,N_18067,N_18217);
or U18484 (N_18484,N_18174,N_18197);
and U18485 (N_18485,N_18246,N_18230);
xnor U18486 (N_18486,N_18117,N_18119);
and U18487 (N_18487,N_18096,N_18056);
or U18488 (N_18488,N_18173,N_18111);
nor U18489 (N_18489,N_18017,N_18169);
xor U18490 (N_18490,N_18071,N_18057);
or U18491 (N_18491,N_18232,N_18194);
or U18492 (N_18492,N_18240,N_18122);
and U18493 (N_18493,N_18063,N_18159);
or U18494 (N_18494,N_18181,N_18106);
nor U18495 (N_18495,N_18053,N_18069);
nor U18496 (N_18496,N_18022,N_18184);
xnor U18497 (N_18497,N_18124,N_18095);
or U18498 (N_18498,N_18049,N_18037);
nor U18499 (N_18499,N_18100,N_18152);
or U18500 (N_18500,N_18460,N_18433);
and U18501 (N_18501,N_18275,N_18288);
xnor U18502 (N_18502,N_18421,N_18337);
nand U18503 (N_18503,N_18308,N_18292);
or U18504 (N_18504,N_18360,N_18314);
and U18505 (N_18505,N_18443,N_18283);
xor U18506 (N_18506,N_18255,N_18355);
xnor U18507 (N_18507,N_18260,N_18340);
nand U18508 (N_18508,N_18434,N_18351);
nor U18509 (N_18509,N_18406,N_18285);
nor U18510 (N_18510,N_18386,N_18378);
or U18511 (N_18511,N_18322,N_18469);
nand U18512 (N_18512,N_18427,N_18279);
nand U18513 (N_18513,N_18422,N_18455);
nand U18514 (N_18514,N_18363,N_18484);
nand U18515 (N_18515,N_18332,N_18440);
or U18516 (N_18516,N_18416,N_18426);
xor U18517 (N_18517,N_18350,N_18453);
or U18518 (N_18518,N_18271,N_18284);
and U18519 (N_18519,N_18399,N_18376);
xor U18520 (N_18520,N_18382,N_18331);
xnor U18521 (N_18521,N_18429,N_18371);
and U18522 (N_18522,N_18449,N_18280);
and U18523 (N_18523,N_18297,N_18454);
nand U18524 (N_18524,N_18373,N_18298);
or U18525 (N_18525,N_18407,N_18320);
nand U18526 (N_18526,N_18310,N_18345);
or U18527 (N_18527,N_18306,N_18390);
nor U18528 (N_18528,N_18420,N_18383);
xor U18529 (N_18529,N_18388,N_18348);
and U18530 (N_18530,N_18341,N_18356);
or U18531 (N_18531,N_18274,N_18273);
nand U18532 (N_18532,N_18483,N_18364);
or U18533 (N_18533,N_18471,N_18423);
nor U18534 (N_18534,N_18456,N_18436);
and U18535 (N_18535,N_18267,N_18482);
nor U18536 (N_18536,N_18408,N_18485);
nand U18537 (N_18537,N_18374,N_18318);
and U18538 (N_18538,N_18492,N_18411);
xnor U18539 (N_18539,N_18402,N_18425);
xor U18540 (N_18540,N_18431,N_18493);
or U18541 (N_18541,N_18344,N_18415);
nor U18542 (N_18542,N_18354,N_18405);
nor U18543 (N_18543,N_18296,N_18282);
xnor U18544 (N_18544,N_18352,N_18265);
nor U18545 (N_18545,N_18457,N_18398);
xnor U18546 (N_18546,N_18389,N_18313);
nand U18547 (N_18547,N_18428,N_18257);
nand U18548 (N_18548,N_18384,N_18358);
xor U18549 (N_18549,N_18252,N_18424);
and U18550 (N_18550,N_18476,N_18262);
nand U18551 (N_18551,N_18495,N_18301);
xnor U18552 (N_18552,N_18319,N_18324);
nor U18553 (N_18553,N_18281,N_18317);
xor U18554 (N_18554,N_18487,N_18307);
or U18555 (N_18555,N_18393,N_18291);
xnor U18556 (N_18556,N_18451,N_18412);
xnor U18557 (N_18557,N_18387,N_18418);
nand U18558 (N_18558,N_18435,N_18299);
nor U18559 (N_18559,N_18253,N_18385);
or U18560 (N_18560,N_18413,N_18343);
or U18561 (N_18561,N_18349,N_18270);
xnor U18562 (N_18562,N_18269,N_18321);
nand U18563 (N_18563,N_18475,N_18309);
nand U18564 (N_18564,N_18368,N_18325);
nor U18565 (N_18565,N_18417,N_18338);
nor U18566 (N_18566,N_18414,N_18300);
xor U18567 (N_18567,N_18468,N_18369);
nor U18568 (N_18568,N_18254,N_18432);
nor U18569 (N_18569,N_18446,N_18347);
nor U18570 (N_18570,N_18463,N_18342);
nand U18571 (N_18571,N_18323,N_18334);
and U18572 (N_18572,N_18489,N_18251);
and U18573 (N_18573,N_18339,N_18330);
nand U18574 (N_18574,N_18365,N_18370);
nand U18575 (N_18575,N_18258,N_18496);
nor U18576 (N_18576,N_18333,N_18250);
or U18577 (N_18577,N_18277,N_18256);
and U18578 (N_18578,N_18261,N_18362);
and U18579 (N_18579,N_18391,N_18259);
nand U18580 (N_18580,N_18444,N_18400);
and U18581 (N_18581,N_18448,N_18381);
nand U18582 (N_18582,N_18294,N_18486);
nor U18583 (N_18583,N_18458,N_18295);
nor U18584 (N_18584,N_18395,N_18490);
xnor U18585 (N_18585,N_18336,N_18410);
xor U18586 (N_18586,N_18450,N_18272);
nor U18587 (N_18587,N_18419,N_18287);
nor U18588 (N_18588,N_18329,N_18477);
or U18589 (N_18589,N_18473,N_18396);
nor U18590 (N_18590,N_18498,N_18461);
nand U18591 (N_18591,N_18499,N_18380);
and U18592 (N_18592,N_18480,N_18401);
nor U18593 (N_18593,N_18442,N_18377);
or U18594 (N_18594,N_18311,N_18403);
nand U18595 (N_18595,N_18459,N_18276);
or U18596 (N_18596,N_18466,N_18379);
and U18597 (N_18597,N_18394,N_18327);
or U18598 (N_18598,N_18264,N_18409);
xnor U18599 (N_18599,N_18438,N_18302);
or U18600 (N_18600,N_18335,N_18346);
and U18601 (N_18601,N_18361,N_18316);
nor U18602 (N_18602,N_18289,N_18293);
or U18603 (N_18603,N_18312,N_18491);
and U18604 (N_18604,N_18478,N_18278);
and U18605 (N_18605,N_18268,N_18392);
nand U18606 (N_18606,N_18488,N_18470);
xor U18607 (N_18607,N_18367,N_18445);
xor U18608 (N_18608,N_18303,N_18439);
nand U18609 (N_18609,N_18430,N_18447);
xor U18610 (N_18610,N_18328,N_18353);
nor U18611 (N_18611,N_18315,N_18465);
xnor U18612 (N_18612,N_18479,N_18494);
or U18613 (N_18613,N_18357,N_18441);
xor U18614 (N_18614,N_18326,N_18290);
xor U18615 (N_18615,N_18437,N_18286);
xnor U18616 (N_18616,N_18366,N_18263);
nor U18617 (N_18617,N_18305,N_18372);
nor U18618 (N_18618,N_18304,N_18462);
or U18619 (N_18619,N_18404,N_18472);
nor U18620 (N_18620,N_18474,N_18266);
and U18621 (N_18621,N_18497,N_18359);
nor U18622 (N_18622,N_18452,N_18467);
and U18623 (N_18623,N_18375,N_18464);
nor U18624 (N_18624,N_18397,N_18481);
and U18625 (N_18625,N_18481,N_18387);
or U18626 (N_18626,N_18252,N_18374);
nand U18627 (N_18627,N_18258,N_18278);
or U18628 (N_18628,N_18347,N_18394);
and U18629 (N_18629,N_18289,N_18437);
or U18630 (N_18630,N_18286,N_18355);
xor U18631 (N_18631,N_18406,N_18271);
nand U18632 (N_18632,N_18341,N_18339);
and U18633 (N_18633,N_18394,N_18422);
and U18634 (N_18634,N_18319,N_18457);
xnor U18635 (N_18635,N_18368,N_18297);
xor U18636 (N_18636,N_18445,N_18251);
or U18637 (N_18637,N_18419,N_18317);
or U18638 (N_18638,N_18372,N_18267);
nor U18639 (N_18639,N_18321,N_18472);
xnor U18640 (N_18640,N_18312,N_18467);
nor U18641 (N_18641,N_18436,N_18299);
nand U18642 (N_18642,N_18333,N_18385);
xnor U18643 (N_18643,N_18410,N_18287);
nor U18644 (N_18644,N_18441,N_18424);
xnor U18645 (N_18645,N_18410,N_18463);
nand U18646 (N_18646,N_18373,N_18351);
or U18647 (N_18647,N_18454,N_18442);
or U18648 (N_18648,N_18285,N_18306);
nor U18649 (N_18649,N_18329,N_18366);
and U18650 (N_18650,N_18376,N_18496);
nand U18651 (N_18651,N_18291,N_18443);
nand U18652 (N_18652,N_18488,N_18271);
nor U18653 (N_18653,N_18397,N_18352);
nor U18654 (N_18654,N_18482,N_18287);
nor U18655 (N_18655,N_18255,N_18444);
nand U18656 (N_18656,N_18399,N_18266);
nor U18657 (N_18657,N_18332,N_18496);
nand U18658 (N_18658,N_18406,N_18447);
nor U18659 (N_18659,N_18440,N_18361);
or U18660 (N_18660,N_18453,N_18295);
nand U18661 (N_18661,N_18451,N_18359);
nand U18662 (N_18662,N_18266,N_18443);
and U18663 (N_18663,N_18353,N_18350);
and U18664 (N_18664,N_18486,N_18259);
nand U18665 (N_18665,N_18271,N_18373);
or U18666 (N_18666,N_18394,N_18393);
and U18667 (N_18667,N_18325,N_18310);
or U18668 (N_18668,N_18284,N_18467);
xor U18669 (N_18669,N_18288,N_18300);
nand U18670 (N_18670,N_18465,N_18495);
or U18671 (N_18671,N_18251,N_18275);
or U18672 (N_18672,N_18274,N_18298);
nor U18673 (N_18673,N_18490,N_18343);
nand U18674 (N_18674,N_18459,N_18306);
and U18675 (N_18675,N_18391,N_18403);
and U18676 (N_18676,N_18441,N_18282);
nand U18677 (N_18677,N_18447,N_18331);
or U18678 (N_18678,N_18265,N_18260);
and U18679 (N_18679,N_18388,N_18296);
nand U18680 (N_18680,N_18435,N_18476);
or U18681 (N_18681,N_18353,N_18481);
xor U18682 (N_18682,N_18294,N_18379);
xor U18683 (N_18683,N_18401,N_18354);
and U18684 (N_18684,N_18373,N_18418);
xor U18685 (N_18685,N_18388,N_18479);
and U18686 (N_18686,N_18254,N_18290);
and U18687 (N_18687,N_18355,N_18263);
or U18688 (N_18688,N_18398,N_18338);
nor U18689 (N_18689,N_18283,N_18489);
and U18690 (N_18690,N_18260,N_18452);
nand U18691 (N_18691,N_18430,N_18265);
or U18692 (N_18692,N_18264,N_18450);
or U18693 (N_18693,N_18438,N_18335);
xnor U18694 (N_18694,N_18376,N_18329);
nor U18695 (N_18695,N_18390,N_18430);
or U18696 (N_18696,N_18385,N_18470);
nand U18697 (N_18697,N_18357,N_18263);
or U18698 (N_18698,N_18260,N_18347);
and U18699 (N_18699,N_18399,N_18442);
nand U18700 (N_18700,N_18458,N_18350);
nand U18701 (N_18701,N_18251,N_18322);
or U18702 (N_18702,N_18353,N_18451);
and U18703 (N_18703,N_18360,N_18262);
and U18704 (N_18704,N_18429,N_18273);
nor U18705 (N_18705,N_18490,N_18366);
and U18706 (N_18706,N_18342,N_18259);
nand U18707 (N_18707,N_18250,N_18266);
xnor U18708 (N_18708,N_18327,N_18274);
xnor U18709 (N_18709,N_18295,N_18452);
and U18710 (N_18710,N_18338,N_18459);
and U18711 (N_18711,N_18353,N_18370);
and U18712 (N_18712,N_18253,N_18378);
nand U18713 (N_18713,N_18315,N_18397);
nand U18714 (N_18714,N_18412,N_18278);
and U18715 (N_18715,N_18499,N_18339);
or U18716 (N_18716,N_18295,N_18343);
nor U18717 (N_18717,N_18354,N_18455);
nand U18718 (N_18718,N_18299,N_18285);
nor U18719 (N_18719,N_18340,N_18381);
and U18720 (N_18720,N_18327,N_18279);
and U18721 (N_18721,N_18286,N_18333);
nor U18722 (N_18722,N_18261,N_18330);
nor U18723 (N_18723,N_18391,N_18254);
or U18724 (N_18724,N_18266,N_18451);
or U18725 (N_18725,N_18435,N_18389);
or U18726 (N_18726,N_18427,N_18499);
and U18727 (N_18727,N_18272,N_18335);
or U18728 (N_18728,N_18497,N_18378);
xor U18729 (N_18729,N_18272,N_18351);
nor U18730 (N_18730,N_18435,N_18462);
xnor U18731 (N_18731,N_18443,N_18375);
xor U18732 (N_18732,N_18497,N_18398);
xnor U18733 (N_18733,N_18484,N_18299);
xor U18734 (N_18734,N_18262,N_18398);
nor U18735 (N_18735,N_18462,N_18440);
xnor U18736 (N_18736,N_18440,N_18444);
nor U18737 (N_18737,N_18280,N_18329);
xor U18738 (N_18738,N_18285,N_18411);
xor U18739 (N_18739,N_18482,N_18363);
and U18740 (N_18740,N_18455,N_18491);
xor U18741 (N_18741,N_18378,N_18393);
xnor U18742 (N_18742,N_18471,N_18444);
nand U18743 (N_18743,N_18273,N_18496);
xnor U18744 (N_18744,N_18309,N_18492);
and U18745 (N_18745,N_18385,N_18287);
xnor U18746 (N_18746,N_18318,N_18344);
and U18747 (N_18747,N_18362,N_18339);
nand U18748 (N_18748,N_18472,N_18384);
xnor U18749 (N_18749,N_18274,N_18287);
or U18750 (N_18750,N_18668,N_18711);
nand U18751 (N_18751,N_18709,N_18721);
xnor U18752 (N_18752,N_18653,N_18730);
or U18753 (N_18753,N_18715,N_18518);
nor U18754 (N_18754,N_18595,N_18570);
and U18755 (N_18755,N_18725,N_18639);
nor U18756 (N_18756,N_18645,N_18511);
or U18757 (N_18757,N_18654,N_18661);
or U18758 (N_18758,N_18694,N_18734);
xor U18759 (N_18759,N_18744,N_18665);
nand U18760 (N_18760,N_18666,N_18615);
or U18761 (N_18761,N_18568,N_18728);
and U18762 (N_18762,N_18651,N_18524);
and U18763 (N_18763,N_18713,N_18735);
and U18764 (N_18764,N_18520,N_18591);
or U18765 (N_18765,N_18684,N_18526);
nand U18766 (N_18766,N_18634,N_18510);
nor U18767 (N_18767,N_18696,N_18545);
nand U18768 (N_18768,N_18572,N_18596);
nor U18769 (N_18769,N_18574,N_18675);
nand U18770 (N_18770,N_18682,N_18567);
or U18771 (N_18771,N_18600,N_18731);
nor U18772 (N_18772,N_18611,N_18602);
nor U18773 (N_18773,N_18680,N_18652);
nand U18774 (N_18774,N_18512,N_18544);
xnor U18775 (N_18775,N_18561,N_18739);
and U18776 (N_18776,N_18726,N_18560);
nor U18777 (N_18777,N_18610,N_18552);
nor U18778 (N_18778,N_18742,N_18573);
or U18779 (N_18779,N_18614,N_18535);
xnor U18780 (N_18780,N_18607,N_18530);
nand U18781 (N_18781,N_18692,N_18714);
nand U18782 (N_18782,N_18604,N_18577);
nor U18783 (N_18783,N_18631,N_18729);
and U18784 (N_18784,N_18699,N_18521);
nor U18785 (N_18785,N_18702,N_18594);
and U18786 (N_18786,N_18747,N_18674);
nor U18787 (N_18787,N_18718,N_18579);
nor U18788 (N_18788,N_18618,N_18647);
or U18789 (N_18789,N_18605,N_18622);
nor U18790 (N_18790,N_18550,N_18644);
nor U18791 (N_18791,N_18662,N_18632);
xnor U18792 (N_18792,N_18703,N_18529);
xnor U18793 (N_18793,N_18519,N_18543);
or U18794 (N_18794,N_18501,N_18708);
xor U18795 (N_18795,N_18664,N_18743);
nand U18796 (N_18796,N_18597,N_18583);
nor U18797 (N_18797,N_18569,N_18630);
xnor U18798 (N_18798,N_18626,N_18695);
and U18799 (N_18799,N_18504,N_18556);
nor U18800 (N_18800,N_18658,N_18599);
xnor U18801 (N_18801,N_18660,N_18612);
nor U18802 (N_18802,N_18677,N_18722);
nand U18803 (N_18803,N_18508,N_18659);
nor U18804 (N_18804,N_18513,N_18523);
or U18805 (N_18805,N_18749,N_18541);
or U18806 (N_18806,N_18723,N_18719);
nor U18807 (N_18807,N_18700,N_18720);
or U18808 (N_18808,N_18528,N_18689);
and U18809 (N_18809,N_18522,N_18687);
xnor U18810 (N_18810,N_18534,N_18635);
and U18811 (N_18811,N_18667,N_18643);
nor U18812 (N_18812,N_18616,N_18678);
nor U18813 (N_18813,N_18566,N_18738);
nand U18814 (N_18814,N_18514,N_18636);
xnor U18815 (N_18815,N_18539,N_18669);
nor U18816 (N_18816,N_18638,N_18542);
nand U18817 (N_18817,N_18681,N_18533);
and U18818 (N_18818,N_18690,N_18555);
and U18819 (N_18819,N_18717,N_18531);
nor U18820 (N_18820,N_18502,N_18564);
and U18821 (N_18821,N_18563,N_18624);
nor U18822 (N_18822,N_18628,N_18732);
and U18823 (N_18823,N_18633,N_18565);
nand U18824 (N_18824,N_18617,N_18698);
xor U18825 (N_18825,N_18705,N_18707);
xor U18826 (N_18826,N_18736,N_18503);
and U18827 (N_18827,N_18554,N_18562);
nor U18828 (N_18828,N_18685,N_18546);
nor U18829 (N_18829,N_18640,N_18507);
xor U18830 (N_18830,N_18549,N_18655);
nor U18831 (N_18831,N_18670,N_18724);
and U18832 (N_18832,N_18500,N_18525);
or U18833 (N_18833,N_18538,N_18505);
nor U18834 (N_18834,N_18532,N_18537);
or U18835 (N_18835,N_18515,N_18740);
nor U18836 (N_18836,N_18587,N_18540);
or U18837 (N_18837,N_18701,N_18716);
and U18838 (N_18838,N_18683,N_18578);
nor U18839 (N_18839,N_18619,N_18646);
nand U18840 (N_18840,N_18623,N_18727);
nor U18841 (N_18841,N_18745,N_18584);
xnor U18842 (N_18842,N_18517,N_18509);
nor U18843 (N_18843,N_18641,N_18582);
xor U18844 (N_18844,N_18558,N_18676);
and U18845 (N_18845,N_18613,N_18516);
nand U18846 (N_18846,N_18656,N_18592);
nand U18847 (N_18847,N_18637,N_18575);
and U18848 (N_18848,N_18671,N_18598);
and U18849 (N_18849,N_18649,N_18548);
or U18850 (N_18850,N_18733,N_18527);
nand U18851 (N_18851,N_18648,N_18559);
and U18852 (N_18852,N_18629,N_18551);
or U18853 (N_18853,N_18547,N_18741);
xor U18854 (N_18854,N_18580,N_18686);
or U18855 (N_18855,N_18589,N_18693);
nor U18856 (N_18856,N_18691,N_18608);
and U18857 (N_18857,N_18506,N_18601);
nand U18858 (N_18858,N_18581,N_18712);
nand U18859 (N_18859,N_18679,N_18688);
xor U18860 (N_18860,N_18748,N_18557);
and U18861 (N_18861,N_18650,N_18672);
nor U18862 (N_18862,N_18663,N_18706);
nor U18863 (N_18863,N_18536,N_18657);
nor U18864 (N_18864,N_18586,N_18609);
and U18865 (N_18865,N_18673,N_18625);
nand U18866 (N_18866,N_18606,N_18576);
and U18867 (N_18867,N_18588,N_18621);
xnor U18868 (N_18868,N_18737,N_18620);
nand U18869 (N_18869,N_18697,N_18710);
nor U18870 (N_18870,N_18593,N_18585);
or U18871 (N_18871,N_18590,N_18704);
and U18872 (N_18872,N_18553,N_18746);
xor U18873 (N_18873,N_18627,N_18603);
and U18874 (N_18874,N_18642,N_18571);
or U18875 (N_18875,N_18615,N_18677);
nand U18876 (N_18876,N_18537,N_18500);
xor U18877 (N_18877,N_18549,N_18504);
and U18878 (N_18878,N_18621,N_18741);
nor U18879 (N_18879,N_18525,N_18654);
or U18880 (N_18880,N_18539,N_18651);
or U18881 (N_18881,N_18744,N_18586);
and U18882 (N_18882,N_18556,N_18577);
and U18883 (N_18883,N_18558,N_18711);
or U18884 (N_18884,N_18613,N_18736);
and U18885 (N_18885,N_18727,N_18748);
or U18886 (N_18886,N_18716,N_18618);
and U18887 (N_18887,N_18515,N_18655);
and U18888 (N_18888,N_18660,N_18747);
and U18889 (N_18889,N_18519,N_18605);
or U18890 (N_18890,N_18531,N_18551);
and U18891 (N_18891,N_18544,N_18533);
xnor U18892 (N_18892,N_18715,N_18569);
nor U18893 (N_18893,N_18521,N_18580);
xnor U18894 (N_18894,N_18706,N_18732);
nor U18895 (N_18895,N_18559,N_18528);
or U18896 (N_18896,N_18535,N_18669);
or U18897 (N_18897,N_18636,N_18587);
or U18898 (N_18898,N_18693,N_18658);
and U18899 (N_18899,N_18658,N_18716);
xnor U18900 (N_18900,N_18690,N_18665);
and U18901 (N_18901,N_18683,N_18660);
xnor U18902 (N_18902,N_18623,N_18644);
xor U18903 (N_18903,N_18653,N_18719);
nand U18904 (N_18904,N_18566,N_18623);
xnor U18905 (N_18905,N_18699,N_18729);
nor U18906 (N_18906,N_18711,N_18543);
xnor U18907 (N_18907,N_18630,N_18573);
nand U18908 (N_18908,N_18648,N_18582);
or U18909 (N_18909,N_18746,N_18715);
or U18910 (N_18910,N_18704,N_18697);
nor U18911 (N_18911,N_18680,N_18633);
nand U18912 (N_18912,N_18618,N_18639);
and U18913 (N_18913,N_18572,N_18741);
or U18914 (N_18914,N_18607,N_18534);
nand U18915 (N_18915,N_18634,N_18529);
xnor U18916 (N_18916,N_18583,N_18563);
and U18917 (N_18917,N_18628,N_18721);
nand U18918 (N_18918,N_18619,N_18573);
or U18919 (N_18919,N_18686,N_18611);
nor U18920 (N_18920,N_18629,N_18628);
or U18921 (N_18921,N_18575,N_18538);
nand U18922 (N_18922,N_18585,N_18621);
xor U18923 (N_18923,N_18519,N_18712);
xnor U18924 (N_18924,N_18613,N_18733);
xor U18925 (N_18925,N_18670,N_18593);
and U18926 (N_18926,N_18539,N_18714);
nand U18927 (N_18927,N_18710,N_18534);
nor U18928 (N_18928,N_18736,N_18562);
xor U18929 (N_18929,N_18551,N_18721);
nor U18930 (N_18930,N_18595,N_18722);
nor U18931 (N_18931,N_18739,N_18578);
nand U18932 (N_18932,N_18582,N_18616);
xnor U18933 (N_18933,N_18550,N_18605);
nor U18934 (N_18934,N_18708,N_18720);
xor U18935 (N_18935,N_18637,N_18722);
nor U18936 (N_18936,N_18668,N_18692);
or U18937 (N_18937,N_18681,N_18647);
xor U18938 (N_18938,N_18735,N_18651);
or U18939 (N_18939,N_18709,N_18720);
xor U18940 (N_18940,N_18516,N_18691);
nand U18941 (N_18941,N_18535,N_18683);
xor U18942 (N_18942,N_18561,N_18669);
or U18943 (N_18943,N_18666,N_18508);
and U18944 (N_18944,N_18568,N_18592);
and U18945 (N_18945,N_18556,N_18521);
nor U18946 (N_18946,N_18587,N_18749);
xnor U18947 (N_18947,N_18502,N_18651);
xor U18948 (N_18948,N_18665,N_18669);
or U18949 (N_18949,N_18632,N_18681);
and U18950 (N_18950,N_18706,N_18610);
or U18951 (N_18951,N_18500,N_18688);
xor U18952 (N_18952,N_18616,N_18608);
nor U18953 (N_18953,N_18678,N_18634);
and U18954 (N_18954,N_18748,N_18543);
or U18955 (N_18955,N_18699,N_18600);
nand U18956 (N_18956,N_18663,N_18578);
and U18957 (N_18957,N_18692,N_18598);
nor U18958 (N_18958,N_18733,N_18603);
xnor U18959 (N_18959,N_18576,N_18670);
or U18960 (N_18960,N_18653,N_18541);
xor U18961 (N_18961,N_18513,N_18555);
nor U18962 (N_18962,N_18517,N_18731);
and U18963 (N_18963,N_18590,N_18525);
xor U18964 (N_18964,N_18743,N_18541);
xnor U18965 (N_18965,N_18631,N_18539);
xor U18966 (N_18966,N_18697,N_18718);
nor U18967 (N_18967,N_18525,N_18502);
nor U18968 (N_18968,N_18528,N_18524);
or U18969 (N_18969,N_18645,N_18635);
and U18970 (N_18970,N_18658,N_18728);
xor U18971 (N_18971,N_18684,N_18685);
nand U18972 (N_18972,N_18730,N_18663);
xor U18973 (N_18973,N_18701,N_18602);
or U18974 (N_18974,N_18670,N_18567);
or U18975 (N_18975,N_18724,N_18643);
nand U18976 (N_18976,N_18708,N_18594);
and U18977 (N_18977,N_18715,N_18693);
nand U18978 (N_18978,N_18572,N_18749);
or U18979 (N_18979,N_18579,N_18666);
and U18980 (N_18980,N_18665,N_18549);
and U18981 (N_18981,N_18701,N_18542);
or U18982 (N_18982,N_18561,N_18674);
and U18983 (N_18983,N_18747,N_18610);
nand U18984 (N_18984,N_18701,N_18512);
nor U18985 (N_18985,N_18716,N_18699);
and U18986 (N_18986,N_18726,N_18562);
nor U18987 (N_18987,N_18526,N_18653);
xnor U18988 (N_18988,N_18661,N_18547);
xor U18989 (N_18989,N_18728,N_18708);
and U18990 (N_18990,N_18500,N_18703);
nand U18991 (N_18991,N_18637,N_18672);
and U18992 (N_18992,N_18671,N_18576);
and U18993 (N_18993,N_18665,N_18671);
or U18994 (N_18994,N_18733,N_18606);
or U18995 (N_18995,N_18553,N_18727);
nand U18996 (N_18996,N_18732,N_18671);
nand U18997 (N_18997,N_18500,N_18510);
or U18998 (N_18998,N_18548,N_18553);
xnor U18999 (N_18999,N_18695,N_18599);
or U19000 (N_19000,N_18785,N_18781);
or U19001 (N_19001,N_18956,N_18971);
or U19002 (N_19002,N_18862,N_18866);
xnor U19003 (N_19003,N_18803,N_18821);
and U19004 (N_19004,N_18851,N_18874);
nor U19005 (N_19005,N_18825,N_18940);
xnor U19006 (N_19006,N_18761,N_18883);
xor U19007 (N_19007,N_18869,N_18770);
nor U19008 (N_19008,N_18878,N_18783);
xor U19009 (N_19009,N_18934,N_18918);
nor U19010 (N_19010,N_18993,N_18964);
nand U19011 (N_19011,N_18778,N_18840);
nand U19012 (N_19012,N_18750,N_18890);
nor U19013 (N_19013,N_18786,N_18978);
or U19014 (N_19014,N_18805,N_18804);
and U19015 (N_19015,N_18903,N_18856);
and U19016 (N_19016,N_18962,N_18985);
and U19017 (N_19017,N_18932,N_18996);
nor U19018 (N_19018,N_18974,N_18854);
nor U19019 (N_19019,N_18769,N_18759);
or U19020 (N_19020,N_18948,N_18842);
and U19021 (N_19021,N_18773,N_18975);
nor U19022 (N_19022,N_18861,N_18920);
nor U19023 (N_19023,N_18913,N_18855);
nand U19024 (N_19024,N_18958,N_18826);
and U19025 (N_19025,N_18789,N_18941);
nand U19026 (N_19026,N_18827,N_18968);
xnor U19027 (N_19027,N_18905,N_18991);
xnor U19028 (N_19028,N_18927,N_18972);
and U19029 (N_19029,N_18779,N_18796);
nor U19030 (N_19030,N_18983,N_18907);
and U19031 (N_19031,N_18908,N_18839);
and U19032 (N_19032,N_18800,N_18818);
and U19033 (N_19033,N_18950,N_18755);
xor U19034 (N_19034,N_18955,N_18867);
and U19035 (N_19035,N_18836,N_18772);
nand U19036 (N_19036,N_18868,N_18898);
and U19037 (N_19037,N_18838,N_18774);
nor U19038 (N_19038,N_18797,N_18888);
nor U19039 (N_19039,N_18792,N_18776);
xor U19040 (N_19040,N_18926,N_18909);
or U19041 (N_19041,N_18989,N_18764);
nand U19042 (N_19042,N_18756,N_18945);
xor U19043 (N_19043,N_18843,N_18794);
nand U19044 (N_19044,N_18911,N_18901);
or U19045 (N_19045,N_18849,N_18850);
nand U19046 (N_19046,N_18767,N_18837);
and U19047 (N_19047,N_18939,N_18963);
nor U19048 (N_19048,N_18885,N_18808);
or U19049 (N_19049,N_18981,N_18917);
or U19050 (N_19050,N_18806,N_18844);
and U19051 (N_19051,N_18896,N_18810);
nand U19052 (N_19052,N_18775,N_18899);
xnor U19053 (N_19053,N_18995,N_18858);
nand U19054 (N_19054,N_18892,N_18947);
and U19055 (N_19055,N_18997,N_18906);
xnor U19056 (N_19056,N_18863,N_18987);
xor U19057 (N_19057,N_18999,N_18782);
nor U19058 (N_19058,N_18807,N_18829);
and U19059 (N_19059,N_18799,N_18768);
nor U19060 (N_19060,N_18752,N_18816);
and U19061 (N_19061,N_18998,N_18910);
nand U19062 (N_19062,N_18845,N_18887);
nand U19063 (N_19063,N_18875,N_18884);
or U19064 (N_19064,N_18852,N_18787);
nand U19065 (N_19065,N_18790,N_18977);
xor U19066 (N_19066,N_18943,N_18865);
xor U19067 (N_19067,N_18988,N_18886);
and U19068 (N_19068,N_18793,N_18966);
nor U19069 (N_19069,N_18933,N_18814);
nor U19070 (N_19070,N_18915,N_18946);
nand U19071 (N_19071,N_18760,N_18980);
xnor U19072 (N_19072,N_18833,N_18965);
nor U19073 (N_19073,N_18949,N_18802);
nor U19074 (N_19074,N_18812,N_18938);
and U19075 (N_19075,N_18848,N_18990);
or U19076 (N_19076,N_18986,N_18900);
and U19077 (N_19077,N_18811,N_18766);
nor U19078 (N_19078,N_18824,N_18984);
xnor U19079 (N_19079,N_18753,N_18864);
nand U19080 (N_19080,N_18809,N_18820);
and U19081 (N_19081,N_18795,N_18817);
nor U19082 (N_19082,N_18944,N_18951);
or U19083 (N_19083,N_18872,N_18902);
and U19084 (N_19084,N_18813,N_18882);
or U19085 (N_19085,N_18819,N_18919);
or U19086 (N_19086,N_18930,N_18841);
and U19087 (N_19087,N_18967,N_18780);
xnor U19088 (N_19088,N_18823,N_18982);
or U19089 (N_19089,N_18784,N_18834);
xnor U19090 (N_19090,N_18889,N_18828);
xnor U19091 (N_19091,N_18970,N_18928);
and U19092 (N_19092,N_18931,N_18912);
or U19093 (N_19093,N_18959,N_18922);
xor U19094 (N_19094,N_18873,N_18914);
nand U19095 (N_19095,N_18871,N_18857);
nand U19096 (N_19096,N_18788,N_18937);
and U19097 (N_19097,N_18879,N_18954);
nand U19098 (N_19098,N_18757,N_18835);
nor U19099 (N_19099,N_18935,N_18870);
and U19100 (N_19100,N_18957,N_18846);
nand U19101 (N_19101,N_18895,N_18751);
and U19102 (N_19102,N_18880,N_18894);
and U19103 (N_19103,N_18801,N_18765);
and U19104 (N_19104,N_18777,N_18953);
nand U19105 (N_19105,N_18936,N_18762);
xor U19106 (N_19106,N_18952,N_18771);
nor U19107 (N_19107,N_18923,N_18754);
xor U19108 (N_19108,N_18859,N_18847);
or U19109 (N_19109,N_18853,N_18960);
and U19110 (N_19110,N_18830,N_18992);
or U19111 (N_19111,N_18976,N_18798);
xor U19112 (N_19112,N_18994,N_18893);
or U19113 (N_19113,N_18791,N_18904);
and U19114 (N_19114,N_18961,N_18973);
nor U19115 (N_19115,N_18891,N_18881);
or U19116 (N_19116,N_18876,N_18832);
nor U19117 (N_19117,N_18763,N_18860);
nor U19118 (N_19118,N_18921,N_18758);
and U19119 (N_19119,N_18979,N_18815);
nand U19120 (N_19120,N_18916,N_18969);
and U19121 (N_19121,N_18925,N_18831);
nor U19122 (N_19122,N_18877,N_18822);
xor U19123 (N_19123,N_18897,N_18929);
nor U19124 (N_19124,N_18942,N_18924);
and U19125 (N_19125,N_18855,N_18795);
or U19126 (N_19126,N_18928,N_18799);
nor U19127 (N_19127,N_18904,N_18942);
nor U19128 (N_19128,N_18974,N_18911);
nor U19129 (N_19129,N_18915,N_18816);
and U19130 (N_19130,N_18959,N_18813);
nor U19131 (N_19131,N_18993,N_18972);
nor U19132 (N_19132,N_18964,N_18823);
nor U19133 (N_19133,N_18882,N_18837);
nand U19134 (N_19134,N_18813,N_18942);
xor U19135 (N_19135,N_18902,N_18915);
nor U19136 (N_19136,N_18879,N_18870);
xor U19137 (N_19137,N_18840,N_18862);
or U19138 (N_19138,N_18827,N_18815);
and U19139 (N_19139,N_18751,N_18890);
xor U19140 (N_19140,N_18854,N_18976);
or U19141 (N_19141,N_18979,N_18789);
or U19142 (N_19142,N_18848,N_18821);
and U19143 (N_19143,N_18781,N_18754);
nand U19144 (N_19144,N_18764,N_18768);
or U19145 (N_19145,N_18999,N_18828);
nor U19146 (N_19146,N_18859,N_18864);
nand U19147 (N_19147,N_18872,N_18827);
xnor U19148 (N_19148,N_18986,N_18994);
or U19149 (N_19149,N_18874,N_18980);
and U19150 (N_19150,N_18785,N_18897);
or U19151 (N_19151,N_18939,N_18905);
and U19152 (N_19152,N_18950,N_18754);
xnor U19153 (N_19153,N_18811,N_18759);
nand U19154 (N_19154,N_18769,N_18819);
and U19155 (N_19155,N_18962,N_18995);
nand U19156 (N_19156,N_18789,N_18761);
nand U19157 (N_19157,N_18918,N_18814);
and U19158 (N_19158,N_18854,N_18960);
xor U19159 (N_19159,N_18936,N_18929);
or U19160 (N_19160,N_18933,N_18858);
and U19161 (N_19161,N_18875,N_18927);
xor U19162 (N_19162,N_18876,N_18946);
nand U19163 (N_19163,N_18867,N_18903);
nand U19164 (N_19164,N_18912,N_18822);
or U19165 (N_19165,N_18968,N_18960);
nand U19166 (N_19166,N_18847,N_18865);
nor U19167 (N_19167,N_18758,N_18796);
nor U19168 (N_19168,N_18934,N_18757);
or U19169 (N_19169,N_18975,N_18793);
nor U19170 (N_19170,N_18814,N_18856);
xor U19171 (N_19171,N_18752,N_18996);
nor U19172 (N_19172,N_18920,N_18979);
or U19173 (N_19173,N_18766,N_18924);
nand U19174 (N_19174,N_18835,N_18825);
and U19175 (N_19175,N_18869,N_18871);
or U19176 (N_19176,N_18968,N_18880);
xor U19177 (N_19177,N_18767,N_18937);
or U19178 (N_19178,N_18833,N_18891);
and U19179 (N_19179,N_18786,N_18826);
and U19180 (N_19180,N_18929,N_18860);
nor U19181 (N_19181,N_18778,N_18836);
nand U19182 (N_19182,N_18961,N_18865);
or U19183 (N_19183,N_18945,N_18903);
and U19184 (N_19184,N_18751,N_18777);
and U19185 (N_19185,N_18781,N_18983);
nand U19186 (N_19186,N_18766,N_18875);
nand U19187 (N_19187,N_18768,N_18757);
nand U19188 (N_19188,N_18984,N_18955);
and U19189 (N_19189,N_18896,N_18983);
nor U19190 (N_19190,N_18935,N_18827);
nand U19191 (N_19191,N_18945,N_18771);
or U19192 (N_19192,N_18967,N_18980);
nor U19193 (N_19193,N_18750,N_18901);
nor U19194 (N_19194,N_18835,N_18942);
nand U19195 (N_19195,N_18792,N_18999);
nand U19196 (N_19196,N_18851,N_18848);
or U19197 (N_19197,N_18794,N_18793);
or U19198 (N_19198,N_18800,N_18850);
or U19199 (N_19199,N_18956,N_18768);
xnor U19200 (N_19200,N_18890,N_18847);
xnor U19201 (N_19201,N_18868,N_18949);
nand U19202 (N_19202,N_18807,N_18956);
nor U19203 (N_19203,N_18950,N_18961);
or U19204 (N_19204,N_18874,N_18985);
nor U19205 (N_19205,N_18884,N_18830);
nor U19206 (N_19206,N_18997,N_18799);
nand U19207 (N_19207,N_18909,N_18875);
nor U19208 (N_19208,N_18841,N_18886);
nand U19209 (N_19209,N_18942,N_18906);
and U19210 (N_19210,N_18848,N_18825);
nand U19211 (N_19211,N_18878,N_18958);
nor U19212 (N_19212,N_18971,N_18754);
xor U19213 (N_19213,N_18799,N_18931);
nand U19214 (N_19214,N_18863,N_18750);
and U19215 (N_19215,N_18858,N_18817);
nand U19216 (N_19216,N_18992,N_18850);
nand U19217 (N_19217,N_18784,N_18815);
nor U19218 (N_19218,N_18859,N_18790);
nor U19219 (N_19219,N_18980,N_18783);
and U19220 (N_19220,N_18977,N_18919);
nand U19221 (N_19221,N_18994,N_18751);
and U19222 (N_19222,N_18918,N_18906);
nor U19223 (N_19223,N_18998,N_18839);
nor U19224 (N_19224,N_18936,N_18799);
nand U19225 (N_19225,N_18936,N_18772);
nand U19226 (N_19226,N_18824,N_18912);
xor U19227 (N_19227,N_18772,N_18899);
xor U19228 (N_19228,N_18825,N_18910);
nor U19229 (N_19229,N_18782,N_18792);
or U19230 (N_19230,N_18755,N_18973);
nand U19231 (N_19231,N_18796,N_18880);
and U19232 (N_19232,N_18911,N_18930);
xnor U19233 (N_19233,N_18756,N_18981);
and U19234 (N_19234,N_18955,N_18831);
nor U19235 (N_19235,N_18894,N_18951);
nor U19236 (N_19236,N_18968,N_18854);
or U19237 (N_19237,N_18784,N_18796);
and U19238 (N_19238,N_18871,N_18856);
or U19239 (N_19239,N_18984,N_18958);
and U19240 (N_19240,N_18854,N_18927);
and U19241 (N_19241,N_18908,N_18988);
nand U19242 (N_19242,N_18820,N_18956);
nand U19243 (N_19243,N_18925,N_18970);
nor U19244 (N_19244,N_18793,N_18778);
nand U19245 (N_19245,N_18989,N_18792);
nand U19246 (N_19246,N_18769,N_18862);
nor U19247 (N_19247,N_18915,N_18983);
or U19248 (N_19248,N_18889,N_18774);
and U19249 (N_19249,N_18943,N_18893);
or U19250 (N_19250,N_19147,N_19006);
nor U19251 (N_19251,N_19027,N_19129);
nor U19252 (N_19252,N_19068,N_19053);
and U19253 (N_19253,N_19047,N_19054);
nand U19254 (N_19254,N_19114,N_19151);
nor U19255 (N_19255,N_19049,N_19201);
and U19256 (N_19256,N_19168,N_19178);
or U19257 (N_19257,N_19005,N_19166);
or U19258 (N_19258,N_19187,N_19155);
or U19259 (N_19259,N_19014,N_19035);
or U19260 (N_19260,N_19222,N_19139);
xor U19261 (N_19261,N_19095,N_19110);
nor U19262 (N_19262,N_19193,N_19174);
and U19263 (N_19263,N_19196,N_19182);
nor U19264 (N_19264,N_19138,N_19244);
nand U19265 (N_19265,N_19144,N_19093);
or U19266 (N_19266,N_19055,N_19072);
xnor U19267 (N_19267,N_19013,N_19059);
and U19268 (N_19268,N_19097,N_19152);
or U19269 (N_19269,N_19123,N_19164);
or U19270 (N_19270,N_19061,N_19010);
or U19271 (N_19271,N_19169,N_19045);
nor U19272 (N_19272,N_19091,N_19162);
nand U19273 (N_19273,N_19238,N_19119);
or U19274 (N_19274,N_19028,N_19020);
and U19275 (N_19275,N_19009,N_19143);
xor U19276 (N_19276,N_19088,N_19221);
and U19277 (N_19277,N_19070,N_19094);
and U19278 (N_19278,N_19234,N_19112);
and U19279 (N_19279,N_19237,N_19180);
nor U19280 (N_19280,N_19242,N_19023);
xnor U19281 (N_19281,N_19213,N_19186);
or U19282 (N_19282,N_19086,N_19031);
xnor U19283 (N_19283,N_19248,N_19016);
nand U19284 (N_19284,N_19131,N_19230);
xnor U19285 (N_19285,N_19030,N_19024);
nor U19286 (N_19286,N_19223,N_19083);
nor U19287 (N_19287,N_19003,N_19165);
or U19288 (N_19288,N_19007,N_19203);
or U19289 (N_19289,N_19153,N_19000);
nor U19290 (N_19290,N_19171,N_19043);
xor U19291 (N_19291,N_19078,N_19179);
nor U19292 (N_19292,N_19046,N_19198);
nor U19293 (N_19293,N_19160,N_19041);
and U19294 (N_19294,N_19226,N_19181);
nor U19295 (N_19295,N_19154,N_19124);
or U19296 (N_19296,N_19133,N_19033);
or U19297 (N_19297,N_19177,N_19087);
or U19298 (N_19298,N_19192,N_19002);
nor U19299 (N_19299,N_19074,N_19206);
or U19300 (N_19300,N_19113,N_19116);
xor U19301 (N_19301,N_19018,N_19163);
nor U19302 (N_19302,N_19048,N_19077);
or U19303 (N_19303,N_19232,N_19079);
or U19304 (N_19304,N_19224,N_19036);
nand U19305 (N_19305,N_19202,N_19066);
nand U19306 (N_19306,N_19057,N_19246);
nand U19307 (N_19307,N_19157,N_19240);
nand U19308 (N_19308,N_19076,N_19195);
and U19309 (N_19309,N_19120,N_19044);
nor U19310 (N_19310,N_19051,N_19148);
or U19311 (N_19311,N_19249,N_19117);
nand U19312 (N_19312,N_19145,N_19073);
nand U19313 (N_19313,N_19245,N_19106);
xor U19314 (N_19314,N_19128,N_19012);
xnor U19315 (N_19315,N_19205,N_19214);
or U19316 (N_19316,N_19211,N_19040);
nor U19317 (N_19317,N_19219,N_19241);
xnor U19318 (N_19318,N_19137,N_19215);
nand U19319 (N_19319,N_19064,N_19141);
and U19320 (N_19320,N_19140,N_19111);
nand U19321 (N_19321,N_19052,N_19239);
and U19322 (N_19322,N_19204,N_19228);
or U19323 (N_19323,N_19185,N_19058);
nor U19324 (N_19324,N_19021,N_19008);
or U19325 (N_19325,N_19134,N_19015);
nor U19326 (N_19326,N_19183,N_19067);
xor U19327 (N_19327,N_19210,N_19243);
nor U19328 (N_19328,N_19081,N_19135);
nor U19329 (N_19329,N_19109,N_19208);
xor U19330 (N_19330,N_19170,N_19220);
or U19331 (N_19331,N_19056,N_19146);
xor U19332 (N_19332,N_19217,N_19167);
xor U19333 (N_19333,N_19105,N_19038);
nor U19334 (N_19334,N_19218,N_19103);
xor U19335 (N_19335,N_19071,N_19122);
or U19336 (N_19336,N_19184,N_19159);
nor U19337 (N_19337,N_19096,N_19089);
and U19338 (N_19338,N_19001,N_19026);
or U19339 (N_19339,N_19125,N_19063);
and U19340 (N_19340,N_19019,N_19050);
and U19341 (N_19341,N_19209,N_19084);
xnor U19342 (N_19342,N_19188,N_19069);
and U19343 (N_19343,N_19235,N_19212);
xnor U19344 (N_19344,N_19102,N_19101);
nor U19345 (N_19345,N_19216,N_19022);
or U19346 (N_19346,N_19231,N_19229);
or U19347 (N_19347,N_19104,N_19189);
nor U19348 (N_19348,N_19004,N_19197);
nor U19349 (N_19349,N_19130,N_19075);
nand U19350 (N_19350,N_19227,N_19200);
nand U19351 (N_19351,N_19099,N_19121);
or U19352 (N_19352,N_19080,N_19017);
and U19353 (N_19353,N_19107,N_19142);
nor U19354 (N_19354,N_19150,N_19161);
nand U19355 (N_19355,N_19034,N_19029);
or U19356 (N_19356,N_19085,N_19247);
and U19357 (N_19357,N_19172,N_19098);
nand U19358 (N_19358,N_19062,N_19090);
and U19359 (N_19359,N_19136,N_19176);
nand U19360 (N_19360,N_19199,N_19191);
xnor U19361 (N_19361,N_19115,N_19132);
or U19362 (N_19362,N_19082,N_19194);
or U19363 (N_19363,N_19127,N_19118);
nand U19364 (N_19364,N_19156,N_19092);
nor U19365 (N_19365,N_19065,N_19233);
nand U19366 (N_19366,N_19190,N_19011);
and U19367 (N_19367,N_19158,N_19207);
nor U19368 (N_19368,N_19032,N_19225);
or U19369 (N_19369,N_19100,N_19037);
and U19370 (N_19370,N_19042,N_19126);
nor U19371 (N_19371,N_19236,N_19175);
nand U19372 (N_19372,N_19149,N_19039);
nor U19373 (N_19373,N_19108,N_19173);
nand U19374 (N_19374,N_19060,N_19025);
or U19375 (N_19375,N_19046,N_19178);
and U19376 (N_19376,N_19048,N_19051);
nor U19377 (N_19377,N_19022,N_19030);
xnor U19378 (N_19378,N_19154,N_19206);
nor U19379 (N_19379,N_19100,N_19112);
and U19380 (N_19380,N_19146,N_19155);
or U19381 (N_19381,N_19141,N_19015);
or U19382 (N_19382,N_19144,N_19230);
nor U19383 (N_19383,N_19246,N_19171);
xnor U19384 (N_19384,N_19078,N_19083);
nor U19385 (N_19385,N_19130,N_19210);
nor U19386 (N_19386,N_19062,N_19172);
xor U19387 (N_19387,N_19033,N_19210);
nand U19388 (N_19388,N_19037,N_19125);
or U19389 (N_19389,N_19208,N_19165);
and U19390 (N_19390,N_19028,N_19162);
nand U19391 (N_19391,N_19095,N_19242);
and U19392 (N_19392,N_19232,N_19213);
nand U19393 (N_19393,N_19117,N_19226);
nand U19394 (N_19394,N_19226,N_19084);
nor U19395 (N_19395,N_19063,N_19208);
xnor U19396 (N_19396,N_19057,N_19144);
nand U19397 (N_19397,N_19034,N_19155);
xor U19398 (N_19398,N_19079,N_19121);
nand U19399 (N_19399,N_19041,N_19170);
xnor U19400 (N_19400,N_19030,N_19123);
and U19401 (N_19401,N_19109,N_19114);
or U19402 (N_19402,N_19197,N_19057);
and U19403 (N_19403,N_19023,N_19148);
nand U19404 (N_19404,N_19022,N_19159);
xnor U19405 (N_19405,N_19224,N_19067);
nor U19406 (N_19406,N_19072,N_19060);
or U19407 (N_19407,N_19132,N_19162);
or U19408 (N_19408,N_19185,N_19020);
and U19409 (N_19409,N_19164,N_19195);
nor U19410 (N_19410,N_19070,N_19218);
and U19411 (N_19411,N_19019,N_19197);
nand U19412 (N_19412,N_19078,N_19242);
xnor U19413 (N_19413,N_19029,N_19150);
or U19414 (N_19414,N_19246,N_19179);
nand U19415 (N_19415,N_19153,N_19070);
and U19416 (N_19416,N_19053,N_19126);
and U19417 (N_19417,N_19215,N_19087);
nor U19418 (N_19418,N_19148,N_19146);
or U19419 (N_19419,N_19112,N_19130);
or U19420 (N_19420,N_19097,N_19078);
or U19421 (N_19421,N_19221,N_19068);
xnor U19422 (N_19422,N_19096,N_19057);
or U19423 (N_19423,N_19087,N_19203);
nand U19424 (N_19424,N_19157,N_19211);
and U19425 (N_19425,N_19080,N_19245);
nand U19426 (N_19426,N_19193,N_19015);
and U19427 (N_19427,N_19117,N_19071);
and U19428 (N_19428,N_19036,N_19027);
nor U19429 (N_19429,N_19011,N_19188);
nand U19430 (N_19430,N_19059,N_19045);
and U19431 (N_19431,N_19106,N_19025);
xor U19432 (N_19432,N_19207,N_19155);
xor U19433 (N_19433,N_19208,N_19149);
and U19434 (N_19434,N_19103,N_19243);
nor U19435 (N_19435,N_19016,N_19212);
nor U19436 (N_19436,N_19028,N_19165);
and U19437 (N_19437,N_19219,N_19145);
nor U19438 (N_19438,N_19083,N_19059);
xor U19439 (N_19439,N_19234,N_19020);
nand U19440 (N_19440,N_19152,N_19087);
nor U19441 (N_19441,N_19135,N_19150);
and U19442 (N_19442,N_19094,N_19019);
xor U19443 (N_19443,N_19137,N_19101);
xnor U19444 (N_19444,N_19048,N_19094);
xnor U19445 (N_19445,N_19173,N_19209);
xnor U19446 (N_19446,N_19044,N_19040);
and U19447 (N_19447,N_19042,N_19142);
xor U19448 (N_19448,N_19145,N_19034);
and U19449 (N_19449,N_19073,N_19217);
nand U19450 (N_19450,N_19146,N_19202);
xor U19451 (N_19451,N_19077,N_19141);
xnor U19452 (N_19452,N_19099,N_19085);
and U19453 (N_19453,N_19156,N_19243);
nand U19454 (N_19454,N_19178,N_19029);
and U19455 (N_19455,N_19211,N_19102);
nor U19456 (N_19456,N_19179,N_19029);
xor U19457 (N_19457,N_19007,N_19002);
nand U19458 (N_19458,N_19035,N_19196);
nand U19459 (N_19459,N_19028,N_19110);
or U19460 (N_19460,N_19175,N_19176);
nand U19461 (N_19461,N_19137,N_19208);
xor U19462 (N_19462,N_19218,N_19112);
and U19463 (N_19463,N_19162,N_19149);
nand U19464 (N_19464,N_19008,N_19140);
or U19465 (N_19465,N_19159,N_19057);
xor U19466 (N_19466,N_19147,N_19152);
nand U19467 (N_19467,N_19177,N_19091);
and U19468 (N_19468,N_19192,N_19147);
xor U19469 (N_19469,N_19018,N_19042);
and U19470 (N_19470,N_19248,N_19113);
and U19471 (N_19471,N_19116,N_19176);
and U19472 (N_19472,N_19202,N_19087);
nor U19473 (N_19473,N_19209,N_19218);
nand U19474 (N_19474,N_19069,N_19138);
and U19475 (N_19475,N_19050,N_19000);
nand U19476 (N_19476,N_19217,N_19152);
nand U19477 (N_19477,N_19098,N_19033);
or U19478 (N_19478,N_19030,N_19097);
or U19479 (N_19479,N_19212,N_19027);
and U19480 (N_19480,N_19035,N_19088);
nor U19481 (N_19481,N_19191,N_19056);
nand U19482 (N_19482,N_19090,N_19061);
nand U19483 (N_19483,N_19149,N_19138);
or U19484 (N_19484,N_19022,N_19014);
xnor U19485 (N_19485,N_19073,N_19023);
nand U19486 (N_19486,N_19238,N_19026);
or U19487 (N_19487,N_19200,N_19046);
nor U19488 (N_19488,N_19116,N_19002);
nand U19489 (N_19489,N_19033,N_19218);
or U19490 (N_19490,N_19046,N_19235);
nand U19491 (N_19491,N_19031,N_19028);
nor U19492 (N_19492,N_19064,N_19232);
nand U19493 (N_19493,N_19067,N_19165);
or U19494 (N_19494,N_19148,N_19048);
xnor U19495 (N_19495,N_19233,N_19083);
nor U19496 (N_19496,N_19029,N_19073);
or U19497 (N_19497,N_19029,N_19114);
nand U19498 (N_19498,N_19157,N_19036);
or U19499 (N_19499,N_19213,N_19145);
xor U19500 (N_19500,N_19478,N_19393);
and U19501 (N_19501,N_19336,N_19413);
and U19502 (N_19502,N_19343,N_19483);
and U19503 (N_19503,N_19354,N_19275);
nand U19504 (N_19504,N_19280,N_19279);
nor U19505 (N_19505,N_19463,N_19287);
or U19506 (N_19506,N_19266,N_19370);
xnor U19507 (N_19507,N_19338,N_19314);
or U19508 (N_19508,N_19486,N_19305);
xnor U19509 (N_19509,N_19391,N_19258);
and U19510 (N_19510,N_19272,N_19284);
xor U19511 (N_19511,N_19481,N_19489);
or U19512 (N_19512,N_19307,N_19352);
or U19513 (N_19513,N_19276,N_19360);
or U19514 (N_19514,N_19376,N_19437);
or U19515 (N_19515,N_19265,N_19496);
and U19516 (N_19516,N_19297,N_19322);
nor U19517 (N_19517,N_19323,N_19440);
and U19518 (N_19518,N_19274,N_19432);
nor U19519 (N_19519,N_19395,N_19409);
xor U19520 (N_19520,N_19414,N_19306);
and U19521 (N_19521,N_19339,N_19282);
nor U19522 (N_19522,N_19400,N_19436);
nor U19523 (N_19523,N_19263,N_19383);
or U19524 (N_19524,N_19443,N_19388);
and U19525 (N_19525,N_19465,N_19427);
and U19526 (N_19526,N_19459,N_19498);
or U19527 (N_19527,N_19329,N_19411);
or U19528 (N_19528,N_19390,N_19325);
xnor U19529 (N_19529,N_19475,N_19277);
xnor U19530 (N_19530,N_19464,N_19317);
or U19531 (N_19531,N_19349,N_19319);
nand U19532 (N_19532,N_19273,N_19357);
and U19533 (N_19533,N_19442,N_19373);
xnor U19534 (N_19534,N_19353,N_19281);
xnor U19535 (N_19535,N_19366,N_19402);
nor U19536 (N_19536,N_19271,N_19454);
nor U19537 (N_19537,N_19374,N_19270);
and U19538 (N_19538,N_19342,N_19385);
or U19539 (N_19539,N_19394,N_19392);
or U19540 (N_19540,N_19455,N_19453);
and U19541 (N_19541,N_19415,N_19467);
nand U19542 (N_19542,N_19431,N_19365);
xnor U19543 (N_19543,N_19369,N_19350);
and U19544 (N_19544,N_19472,N_19253);
and U19545 (N_19545,N_19401,N_19396);
or U19546 (N_19546,N_19405,N_19381);
nand U19547 (N_19547,N_19468,N_19482);
or U19548 (N_19548,N_19303,N_19285);
nand U19549 (N_19549,N_19315,N_19439);
or U19550 (N_19550,N_19456,N_19458);
nand U19551 (N_19551,N_19452,N_19444);
or U19552 (N_19552,N_19286,N_19267);
nand U19553 (N_19553,N_19477,N_19435);
xor U19554 (N_19554,N_19426,N_19326);
nand U19555 (N_19555,N_19425,N_19497);
nor U19556 (N_19556,N_19490,N_19399);
xnor U19557 (N_19557,N_19371,N_19294);
or U19558 (N_19558,N_19480,N_19368);
xor U19559 (N_19559,N_19335,N_19330);
xnor U19560 (N_19560,N_19340,N_19257);
or U19561 (N_19561,N_19320,N_19445);
nor U19562 (N_19562,N_19324,N_19449);
nor U19563 (N_19563,N_19450,N_19422);
nor U19564 (N_19564,N_19261,N_19389);
or U19565 (N_19565,N_19304,N_19293);
nand U19566 (N_19566,N_19471,N_19355);
or U19567 (N_19567,N_19316,N_19462);
or U19568 (N_19568,N_19384,N_19466);
nand U19569 (N_19569,N_19416,N_19499);
nor U19570 (N_19570,N_19300,N_19312);
nor U19571 (N_19571,N_19259,N_19309);
nand U19572 (N_19572,N_19377,N_19457);
or U19573 (N_19573,N_19408,N_19491);
xnor U19574 (N_19574,N_19447,N_19397);
nand U19575 (N_19575,N_19251,N_19362);
xnor U19576 (N_19576,N_19255,N_19433);
nand U19577 (N_19577,N_19291,N_19260);
xor U19578 (N_19578,N_19407,N_19347);
xnor U19579 (N_19579,N_19327,N_19469);
and U19580 (N_19580,N_19460,N_19488);
or U19581 (N_19581,N_19479,N_19308);
or U19582 (N_19582,N_19250,N_19268);
and U19583 (N_19583,N_19341,N_19359);
nor U19584 (N_19584,N_19387,N_19412);
and U19585 (N_19585,N_19331,N_19404);
nor U19586 (N_19586,N_19429,N_19375);
and U19587 (N_19587,N_19283,N_19430);
nand U19588 (N_19588,N_19333,N_19348);
nand U19589 (N_19589,N_19321,N_19313);
and U19590 (N_19590,N_19364,N_19410);
nand U19591 (N_19591,N_19441,N_19474);
or U19592 (N_19592,N_19406,N_19344);
or U19593 (N_19593,N_19386,N_19337);
nand U19594 (N_19594,N_19351,N_19494);
xnor U19595 (N_19595,N_19424,N_19290);
xor U19596 (N_19596,N_19345,N_19301);
and U19597 (N_19597,N_19252,N_19302);
nand U19598 (N_19598,N_19418,N_19298);
and U19599 (N_19599,N_19332,N_19256);
or U19600 (N_19600,N_19473,N_19403);
and U19601 (N_19601,N_19380,N_19476);
xnor U19602 (N_19602,N_19278,N_19417);
and U19603 (N_19603,N_19428,N_19423);
nor U19604 (N_19604,N_19295,N_19363);
nor U19605 (N_19605,N_19379,N_19492);
xor U19606 (N_19606,N_19484,N_19361);
or U19607 (N_19607,N_19382,N_19378);
xor U19608 (N_19608,N_19269,N_19420);
xnor U19609 (N_19609,N_19311,N_19470);
and U19610 (N_19610,N_19451,N_19292);
xor U19611 (N_19611,N_19296,N_19446);
nand U19612 (N_19612,N_19398,N_19461);
nand U19613 (N_19613,N_19485,N_19356);
or U19614 (N_19614,N_19299,N_19421);
xor U19615 (N_19615,N_19288,N_19328);
xor U19616 (N_19616,N_19372,N_19262);
and U19617 (N_19617,N_19493,N_19318);
xor U19618 (N_19618,N_19419,N_19358);
or U19619 (N_19619,N_19438,N_19448);
or U19620 (N_19620,N_19434,N_19254);
or U19621 (N_19621,N_19310,N_19289);
nand U19622 (N_19622,N_19487,N_19346);
nor U19623 (N_19623,N_19367,N_19495);
nand U19624 (N_19624,N_19334,N_19264);
xor U19625 (N_19625,N_19313,N_19396);
or U19626 (N_19626,N_19334,N_19436);
xor U19627 (N_19627,N_19276,N_19370);
and U19628 (N_19628,N_19255,N_19486);
or U19629 (N_19629,N_19301,N_19253);
and U19630 (N_19630,N_19316,N_19426);
nor U19631 (N_19631,N_19437,N_19415);
xnor U19632 (N_19632,N_19471,N_19423);
nand U19633 (N_19633,N_19316,N_19322);
nor U19634 (N_19634,N_19476,N_19271);
nor U19635 (N_19635,N_19293,N_19463);
and U19636 (N_19636,N_19381,N_19462);
nor U19637 (N_19637,N_19365,N_19420);
xor U19638 (N_19638,N_19424,N_19322);
nor U19639 (N_19639,N_19281,N_19453);
and U19640 (N_19640,N_19392,N_19419);
nor U19641 (N_19641,N_19328,N_19385);
nor U19642 (N_19642,N_19366,N_19391);
or U19643 (N_19643,N_19387,N_19269);
or U19644 (N_19644,N_19455,N_19373);
xor U19645 (N_19645,N_19371,N_19413);
or U19646 (N_19646,N_19404,N_19301);
xor U19647 (N_19647,N_19365,N_19430);
xnor U19648 (N_19648,N_19426,N_19385);
xnor U19649 (N_19649,N_19344,N_19346);
nand U19650 (N_19650,N_19296,N_19337);
and U19651 (N_19651,N_19337,N_19305);
xnor U19652 (N_19652,N_19369,N_19437);
and U19653 (N_19653,N_19414,N_19277);
nor U19654 (N_19654,N_19432,N_19433);
or U19655 (N_19655,N_19297,N_19434);
and U19656 (N_19656,N_19427,N_19268);
nor U19657 (N_19657,N_19438,N_19399);
or U19658 (N_19658,N_19287,N_19291);
nand U19659 (N_19659,N_19469,N_19444);
xnor U19660 (N_19660,N_19261,N_19362);
and U19661 (N_19661,N_19358,N_19317);
and U19662 (N_19662,N_19400,N_19370);
and U19663 (N_19663,N_19479,N_19250);
xor U19664 (N_19664,N_19268,N_19413);
nand U19665 (N_19665,N_19482,N_19392);
nor U19666 (N_19666,N_19499,N_19456);
or U19667 (N_19667,N_19307,N_19359);
or U19668 (N_19668,N_19421,N_19499);
nand U19669 (N_19669,N_19311,N_19459);
xnor U19670 (N_19670,N_19418,N_19379);
xor U19671 (N_19671,N_19386,N_19358);
nor U19672 (N_19672,N_19414,N_19263);
nor U19673 (N_19673,N_19495,N_19286);
and U19674 (N_19674,N_19398,N_19375);
xnor U19675 (N_19675,N_19376,N_19468);
nor U19676 (N_19676,N_19286,N_19277);
nand U19677 (N_19677,N_19383,N_19320);
nor U19678 (N_19678,N_19291,N_19357);
nand U19679 (N_19679,N_19339,N_19411);
nand U19680 (N_19680,N_19328,N_19327);
or U19681 (N_19681,N_19476,N_19336);
and U19682 (N_19682,N_19488,N_19466);
or U19683 (N_19683,N_19357,N_19255);
xnor U19684 (N_19684,N_19422,N_19366);
xor U19685 (N_19685,N_19395,N_19403);
xor U19686 (N_19686,N_19328,N_19382);
and U19687 (N_19687,N_19499,N_19449);
xor U19688 (N_19688,N_19418,N_19320);
nor U19689 (N_19689,N_19484,N_19325);
or U19690 (N_19690,N_19330,N_19332);
nand U19691 (N_19691,N_19319,N_19401);
or U19692 (N_19692,N_19421,N_19425);
or U19693 (N_19693,N_19380,N_19361);
nand U19694 (N_19694,N_19414,N_19337);
nand U19695 (N_19695,N_19282,N_19272);
nor U19696 (N_19696,N_19335,N_19265);
nor U19697 (N_19697,N_19279,N_19434);
nand U19698 (N_19698,N_19332,N_19267);
nor U19699 (N_19699,N_19387,N_19304);
and U19700 (N_19700,N_19456,N_19264);
xor U19701 (N_19701,N_19432,N_19463);
or U19702 (N_19702,N_19383,N_19266);
nor U19703 (N_19703,N_19307,N_19330);
or U19704 (N_19704,N_19446,N_19429);
xnor U19705 (N_19705,N_19409,N_19471);
nor U19706 (N_19706,N_19371,N_19320);
and U19707 (N_19707,N_19431,N_19342);
xnor U19708 (N_19708,N_19343,N_19291);
and U19709 (N_19709,N_19315,N_19347);
xor U19710 (N_19710,N_19372,N_19253);
nand U19711 (N_19711,N_19477,N_19415);
xor U19712 (N_19712,N_19278,N_19494);
xor U19713 (N_19713,N_19479,N_19290);
xnor U19714 (N_19714,N_19363,N_19372);
and U19715 (N_19715,N_19496,N_19286);
and U19716 (N_19716,N_19403,N_19397);
nor U19717 (N_19717,N_19450,N_19250);
or U19718 (N_19718,N_19270,N_19449);
or U19719 (N_19719,N_19464,N_19397);
or U19720 (N_19720,N_19453,N_19382);
xor U19721 (N_19721,N_19441,N_19481);
or U19722 (N_19722,N_19490,N_19454);
or U19723 (N_19723,N_19386,N_19396);
nand U19724 (N_19724,N_19271,N_19260);
nor U19725 (N_19725,N_19333,N_19490);
or U19726 (N_19726,N_19335,N_19498);
nor U19727 (N_19727,N_19347,N_19287);
and U19728 (N_19728,N_19284,N_19433);
or U19729 (N_19729,N_19345,N_19419);
or U19730 (N_19730,N_19426,N_19263);
or U19731 (N_19731,N_19418,N_19399);
nand U19732 (N_19732,N_19293,N_19435);
nand U19733 (N_19733,N_19310,N_19484);
or U19734 (N_19734,N_19287,N_19316);
xor U19735 (N_19735,N_19391,N_19496);
xnor U19736 (N_19736,N_19473,N_19319);
or U19737 (N_19737,N_19314,N_19426);
nor U19738 (N_19738,N_19375,N_19458);
nand U19739 (N_19739,N_19327,N_19421);
xnor U19740 (N_19740,N_19388,N_19409);
and U19741 (N_19741,N_19291,N_19281);
xor U19742 (N_19742,N_19389,N_19375);
xor U19743 (N_19743,N_19271,N_19279);
nand U19744 (N_19744,N_19470,N_19429);
or U19745 (N_19745,N_19269,N_19260);
or U19746 (N_19746,N_19294,N_19402);
nand U19747 (N_19747,N_19366,N_19365);
nor U19748 (N_19748,N_19329,N_19327);
xnor U19749 (N_19749,N_19262,N_19417);
xor U19750 (N_19750,N_19512,N_19686);
or U19751 (N_19751,N_19554,N_19685);
xnor U19752 (N_19752,N_19507,N_19618);
nand U19753 (N_19753,N_19729,N_19639);
xor U19754 (N_19754,N_19516,N_19626);
and U19755 (N_19755,N_19657,N_19720);
or U19756 (N_19756,N_19744,N_19531);
nand U19757 (N_19757,N_19541,N_19612);
nand U19758 (N_19758,N_19680,N_19630);
and U19759 (N_19759,N_19544,N_19610);
xor U19760 (N_19760,N_19600,N_19688);
nor U19761 (N_19761,N_19687,N_19713);
nand U19762 (N_19762,N_19695,N_19517);
or U19763 (N_19763,N_19614,N_19673);
and U19764 (N_19764,N_19563,N_19712);
and U19765 (N_19765,N_19519,N_19530);
nand U19766 (N_19766,N_19606,N_19642);
or U19767 (N_19767,N_19522,N_19534);
xor U19768 (N_19768,N_19679,N_19550);
nor U19769 (N_19769,N_19631,N_19699);
and U19770 (N_19770,N_19553,N_19681);
and U19771 (N_19771,N_19638,N_19537);
and U19772 (N_19772,N_19640,N_19738);
and U19773 (N_19773,N_19532,N_19645);
xnor U19774 (N_19774,N_19654,N_19565);
and U19775 (N_19775,N_19545,N_19667);
and U19776 (N_19776,N_19671,N_19571);
xnor U19777 (N_19777,N_19653,N_19742);
nor U19778 (N_19778,N_19743,N_19584);
or U19779 (N_19779,N_19567,N_19514);
nor U19780 (N_19780,N_19697,N_19595);
or U19781 (N_19781,N_19566,N_19704);
or U19782 (N_19782,N_19669,N_19627);
nand U19783 (N_19783,N_19672,N_19585);
xnor U19784 (N_19784,N_19580,N_19573);
and U19785 (N_19785,N_19579,N_19561);
nand U19786 (N_19786,N_19726,N_19513);
nand U19787 (N_19787,N_19707,N_19528);
nand U19788 (N_19788,N_19521,N_19548);
nor U19789 (N_19789,N_19683,N_19505);
xnor U19790 (N_19790,N_19710,N_19502);
and U19791 (N_19791,N_19508,N_19737);
xnor U19792 (N_19792,N_19594,N_19529);
and U19793 (N_19793,N_19509,N_19655);
nor U19794 (N_19794,N_19598,N_19735);
and U19795 (N_19795,N_19564,N_19637);
nor U19796 (N_19796,N_19547,N_19702);
nor U19797 (N_19797,N_19504,N_19609);
nor U19798 (N_19798,N_19559,N_19734);
nor U19799 (N_19799,N_19590,N_19647);
nor U19800 (N_19800,N_19731,N_19656);
and U19801 (N_19801,N_19725,N_19506);
and U19802 (N_19802,N_19523,N_19659);
nor U19803 (N_19803,N_19730,N_19668);
or U19804 (N_19804,N_19555,N_19501);
xor U19805 (N_19805,N_19616,N_19660);
or U19806 (N_19806,N_19535,N_19719);
and U19807 (N_19807,N_19691,N_19629);
and U19808 (N_19808,N_19611,N_19745);
nor U19809 (N_19809,N_19515,N_19510);
nand U19810 (N_19810,N_19575,N_19677);
and U19811 (N_19811,N_19714,N_19665);
or U19812 (N_19812,N_19727,N_19634);
and U19813 (N_19813,N_19661,N_19666);
nor U19814 (N_19814,N_19636,N_19711);
nor U19815 (N_19815,N_19746,N_19525);
or U19816 (N_19816,N_19601,N_19641);
or U19817 (N_19817,N_19581,N_19748);
nand U19818 (N_19818,N_19582,N_19619);
or U19819 (N_19819,N_19538,N_19692);
nand U19820 (N_19820,N_19705,N_19607);
xnor U19821 (N_19821,N_19694,N_19568);
or U19822 (N_19822,N_19524,N_19676);
nor U19823 (N_19823,N_19662,N_19698);
nand U19824 (N_19824,N_19542,N_19608);
or U19825 (N_19825,N_19703,N_19664);
xor U19826 (N_19826,N_19526,N_19518);
xor U19827 (N_19827,N_19557,N_19520);
and U19828 (N_19828,N_19576,N_19635);
nor U19829 (N_19829,N_19722,N_19622);
nor U19830 (N_19830,N_19625,N_19570);
nand U19831 (N_19831,N_19588,N_19603);
and U19832 (N_19832,N_19690,N_19675);
and U19833 (N_19833,N_19706,N_19723);
or U19834 (N_19834,N_19546,N_19732);
or U19835 (N_19835,N_19733,N_19556);
and U19836 (N_19836,N_19560,N_19684);
and U19837 (N_19837,N_19717,N_19543);
nor U19838 (N_19838,N_19689,N_19511);
nor U19839 (N_19839,N_19740,N_19617);
xor U19840 (N_19840,N_19678,N_19551);
or U19841 (N_19841,N_19670,N_19597);
xnor U19842 (N_19842,N_19583,N_19592);
nand U19843 (N_19843,N_19574,N_19593);
or U19844 (N_19844,N_19682,N_19503);
or U19845 (N_19845,N_19527,N_19728);
xnor U19846 (N_19846,N_19533,N_19596);
nor U19847 (N_19847,N_19701,N_19628);
nand U19848 (N_19848,N_19623,N_19500);
xnor U19849 (N_19849,N_19589,N_19736);
nor U19850 (N_19850,N_19646,N_19715);
or U19851 (N_19851,N_19650,N_19747);
xor U19852 (N_19852,N_19591,N_19577);
nor U19853 (N_19853,N_19602,N_19700);
nor U19854 (N_19854,N_19562,N_19649);
xor U19855 (N_19855,N_19693,N_19539);
or U19856 (N_19856,N_19663,N_19615);
and U19857 (N_19857,N_19604,N_19718);
or U19858 (N_19858,N_19572,N_19708);
xnor U19859 (N_19859,N_19644,N_19549);
or U19860 (N_19860,N_19633,N_19605);
nor U19861 (N_19861,N_19586,N_19578);
or U19862 (N_19862,N_19724,N_19613);
xor U19863 (N_19863,N_19621,N_19624);
and U19864 (N_19864,N_19599,N_19632);
nor U19865 (N_19865,N_19648,N_19540);
nand U19866 (N_19866,N_19749,N_19739);
xor U19867 (N_19867,N_19569,N_19587);
nand U19868 (N_19868,N_19721,N_19674);
nor U19869 (N_19869,N_19741,N_19536);
xnor U19870 (N_19870,N_19716,N_19558);
nand U19871 (N_19871,N_19709,N_19552);
xnor U19872 (N_19872,N_19643,N_19658);
nand U19873 (N_19873,N_19620,N_19651);
xor U19874 (N_19874,N_19696,N_19652);
and U19875 (N_19875,N_19526,N_19537);
nand U19876 (N_19876,N_19594,N_19738);
or U19877 (N_19877,N_19641,N_19707);
and U19878 (N_19878,N_19581,N_19529);
and U19879 (N_19879,N_19682,N_19511);
xor U19880 (N_19880,N_19619,N_19738);
xor U19881 (N_19881,N_19580,N_19586);
nand U19882 (N_19882,N_19654,N_19712);
or U19883 (N_19883,N_19697,N_19503);
nand U19884 (N_19884,N_19728,N_19669);
nand U19885 (N_19885,N_19620,N_19577);
xor U19886 (N_19886,N_19593,N_19556);
xor U19887 (N_19887,N_19720,N_19602);
xor U19888 (N_19888,N_19507,N_19717);
nor U19889 (N_19889,N_19508,N_19590);
and U19890 (N_19890,N_19717,N_19619);
and U19891 (N_19891,N_19744,N_19740);
nor U19892 (N_19892,N_19628,N_19536);
or U19893 (N_19893,N_19589,N_19710);
nand U19894 (N_19894,N_19687,N_19716);
nand U19895 (N_19895,N_19704,N_19565);
nand U19896 (N_19896,N_19585,N_19712);
or U19897 (N_19897,N_19606,N_19591);
and U19898 (N_19898,N_19528,N_19554);
nand U19899 (N_19899,N_19590,N_19746);
nand U19900 (N_19900,N_19644,N_19616);
and U19901 (N_19901,N_19574,N_19615);
xor U19902 (N_19902,N_19688,N_19642);
nor U19903 (N_19903,N_19606,N_19705);
or U19904 (N_19904,N_19693,N_19562);
nor U19905 (N_19905,N_19541,N_19512);
xor U19906 (N_19906,N_19697,N_19536);
xor U19907 (N_19907,N_19729,N_19733);
xnor U19908 (N_19908,N_19648,N_19533);
and U19909 (N_19909,N_19573,N_19618);
and U19910 (N_19910,N_19627,N_19703);
and U19911 (N_19911,N_19523,N_19604);
xor U19912 (N_19912,N_19627,N_19588);
nand U19913 (N_19913,N_19616,N_19570);
or U19914 (N_19914,N_19730,N_19578);
xor U19915 (N_19915,N_19711,N_19712);
xnor U19916 (N_19916,N_19516,N_19735);
or U19917 (N_19917,N_19651,N_19716);
or U19918 (N_19918,N_19692,N_19597);
nand U19919 (N_19919,N_19654,N_19593);
or U19920 (N_19920,N_19749,N_19512);
or U19921 (N_19921,N_19562,N_19567);
nor U19922 (N_19922,N_19651,N_19652);
nor U19923 (N_19923,N_19649,N_19547);
and U19924 (N_19924,N_19610,N_19648);
and U19925 (N_19925,N_19706,N_19514);
or U19926 (N_19926,N_19520,N_19634);
and U19927 (N_19927,N_19724,N_19646);
and U19928 (N_19928,N_19503,N_19723);
xnor U19929 (N_19929,N_19503,N_19587);
xnor U19930 (N_19930,N_19518,N_19606);
nor U19931 (N_19931,N_19621,N_19531);
and U19932 (N_19932,N_19507,N_19737);
nor U19933 (N_19933,N_19630,N_19592);
xor U19934 (N_19934,N_19713,N_19541);
xor U19935 (N_19935,N_19566,N_19568);
nor U19936 (N_19936,N_19619,N_19639);
nor U19937 (N_19937,N_19743,N_19687);
nor U19938 (N_19938,N_19656,N_19651);
or U19939 (N_19939,N_19652,N_19640);
xnor U19940 (N_19940,N_19749,N_19546);
and U19941 (N_19941,N_19670,N_19731);
nand U19942 (N_19942,N_19597,N_19575);
xor U19943 (N_19943,N_19638,N_19585);
and U19944 (N_19944,N_19519,N_19523);
nor U19945 (N_19945,N_19618,N_19601);
or U19946 (N_19946,N_19716,N_19738);
nor U19947 (N_19947,N_19702,N_19565);
or U19948 (N_19948,N_19727,N_19701);
nand U19949 (N_19949,N_19686,N_19662);
or U19950 (N_19950,N_19632,N_19705);
nor U19951 (N_19951,N_19652,N_19608);
xor U19952 (N_19952,N_19709,N_19554);
nand U19953 (N_19953,N_19624,N_19614);
or U19954 (N_19954,N_19554,N_19690);
nand U19955 (N_19955,N_19733,N_19531);
nand U19956 (N_19956,N_19685,N_19546);
and U19957 (N_19957,N_19609,N_19742);
or U19958 (N_19958,N_19501,N_19719);
nand U19959 (N_19959,N_19511,N_19731);
xor U19960 (N_19960,N_19622,N_19634);
or U19961 (N_19961,N_19693,N_19524);
or U19962 (N_19962,N_19749,N_19632);
nor U19963 (N_19963,N_19500,N_19610);
xnor U19964 (N_19964,N_19694,N_19620);
nand U19965 (N_19965,N_19619,N_19681);
and U19966 (N_19966,N_19640,N_19584);
nor U19967 (N_19967,N_19536,N_19728);
xor U19968 (N_19968,N_19664,N_19680);
nand U19969 (N_19969,N_19589,N_19566);
or U19970 (N_19970,N_19593,N_19749);
or U19971 (N_19971,N_19587,N_19697);
and U19972 (N_19972,N_19669,N_19541);
nand U19973 (N_19973,N_19602,N_19674);
nand U19974 (N_19974,N_19657,N_19671);
xor U19975 (N_19975,N_19650,N_19694);
or U19976 (N_19976,N_19616,N_19711);
and U19977 (N_19977,N_19574,N_19657);
nand U19978 (N_19978,N_19553,N_19546);
xnor U19979 (N_19979,N_19701,N_19749);
or U19980 (N_19980,N_19690,N_19505);
xor U19981 (N_19981,N_19720,N_19654);
xnor U19982 (N_19982,N_19507,N_19703);
xor U19983 (N_19983,N_19701,N_19606);
or U19984 (N_19984,N_19629,N_19602);
nand U19985 (N_19985,N_19665,N_19643);
nand U19986 (N_19986,N_19672,N_19687);
or U19987 (N_19987,N_19655,N_19548);
nor U19988 (N_19988,N_19506,N_19568);
xnor U19989 (N_19989,N_19575,N_19559);
and U19990 (N_19990,N_19568,N_19581);
xor U19991 (N_19991,N_19712,N_19653);
and U19992 (N_19992,N_19528,N_19643);
xnor U19993 (N_19993,N_19586,N_19613);
and U19994 (N_19994,N_19648,N_19681);
or U19995 (N_19995,N_19712,N_19512);
xnor U19996 (N_19996,N_19523,N_19633);
or U19997 (N_19997,N_19667,N_19679);
nor U19998 (N_19998,N_19530,N_19655);
nand U19999 (N_19999,N_19517,N_19733);
nor U20000 (N_20000,N_19913,N_19956);
xor U20001 (N_20001,N_19943,N_19901);
xnor U20002 (N_20002,N_19835,N_19949);
nand U20003 (N_20003,N_19841,N_19850);
nand U20004 (N_20004,N_19767,N_19814);
nor U20005 (N_20005,N_19889,N_19908);
and U20006 (N_20006,N_19959,N_19880);
and U20007 (N_20007,N_19924,N_19948);
nand U20008 (N_20008,N_19992,N_19786);
and U20009 (N_20009,N_19967,N_19994);
xor U20010 (N_20010,N_19849,N_19754);
xor U20011 (N_20011,N_19751,N_19885);
nor U20012 (N_20012,N_19761,N_19920);
xor U20013 (N_20013,N_19810,N_19971);
or U20014 (N_20014,N_19927,N_19960);
or U20015 (N_20015,N_19921,N_19929);
nand U20016 (N_20016,N_19827,N_19890);
nor U20017 (N_20017,N_19842,N_19799);
nand U20018 (N_20018,N_19881,N_19978);
or U20019 (N_20019,N_19918,N_19750);
or U20020 (N_20020,N_19912,N_19982);
and U20021 (N_20021,N_19937,N_19891);
and U20022 (N_20022,N_19990,N_19866);
or U20023 (N_20023,N_19800,N_19764);
or U20024 (N_20024,N_19807,N_19878);
nand U20025 (N_20025,N_19855,N_19968);
nor U20026 (N_20026,N_19771,N_19780);
or U20027 (N_20027,N_19832,N_19875);
nand U20028 (N_20028,N_19934,N_19864);
or U20029 (N_20029,N_19820,N_19765);
and U20030 (N_20030,N_19945,N_19847);
xor U20031 (N_20031,N_19833,N_19887);
nor U20032 (N_20032,N_19942,N_19839);
or U20033 (N_20033,N_19845,N_19953);
or U20034 (N_20034,N_19843,N_19970);
nand U20035 (N_20035,N_19860,N_19798);
xor U20036 (N_20036,N_19870,N_19914);
xnor U20037 (N_20037,N_19922,N_19760);
nor U20038 (N_20038,N_19919,N_19974);
xnor U20039 (N_20039,N_19854,N_19972);
nor U20040 (N_20040,N_19784,N_19862);
xor U20041 (N_20041,N_19886,N_19865);
or U20042 (N_20042,N_19774,N_19828);
nor U20043 (N_20043,N_19838,N_19877);
or U20044 (N_20044,N_19902,N_19907);
or U20045 (N_20045,N_19925,N_19980);
nor U20046 (N_20046,N_19769,N_19926);
nor U20047 (N_20047,N_19822,N_19973);
nor U20048 (N_20048,N_19884,N_19808);
or U20049 (N_20049,N_19778,N_19869);
nor U20050 (N_20050,N_19876,N_19755);
nor U20051 (N_20051,N_19773,N_19836);
xor U20052 (N_20052,N_19830,N_19991);
nand U20053 (N_20053,N_19962,N_19928);
xor U20054 (N_20054,N_19763,N_19868);
nand U20055 (N_20055,N_19904,N_19947);
nand U20056 (N_20056,N_19939,N_19759);
nor U20057 (N_20057,N_19858,N_19861);
nor U20058 (N_20058,N_19995,N_19752);
nor U20059 (N_20059,N_19976,N_19882);
nand U20060 (N_20060,N_19906,N_19824);
nor U20061 (N_20061,N_19898,N_19793);
and U20062 (N_20062,N_19916,N_19900);
xnor U20063 (N_20063,N_19987,N_19903);
xor U20064 (N_20064,N_19909,N_19796);
or U20065 (N_20065,N_19917,N_19977);
xor U20066 (N_20066,N_19895,N_19811);
nor U20067 (N_20067,N_19941,N_19821);
and U20068 (N_20068,N_19753,N_19965);
and U20069 (N_20069,N_19950,N_19879);
nor U20070 (N_20070,N_19979,N_19857);
xnor U20071 (N_20071,N_19938,N_19844);
nand U20072 (N_20072,N_19911,N_19999);
or U20073 (N_20073,N_19923,N_19788);
or U20074 (N_20074,N_19888,N_19961);
nor U20075 (N_20075,N_19964,N_19766);
nand U20076 (N_20076,N_19932,N_19770);
or U20077 (N_20077,N_19874,N_19791);
or U20078 (N_20078,N_19789,N_19983);
or U20079 (N_20079,N_19993,N_19944);
xnor U20080 (N_20080,N_19803,N_19856);
or U20081 (N_20081,N_19989,N_19883);
and U20082 (N_20082,N_19825,N_19984);
nor U20083 (N_20083,N_19815,N_19829);
nand U20084 (N_20084,N_19863,N_19872);
nand U20085 (N_20085,N_19893,N_19936);
nand U20086 (N_20086,N_19975,N_19782);
and U20087 (N_20087,N_19951,N_19899);
and U20088 (N_20088,N_19958,N_19823);
nor U20089 (N_20089,N_19867,N_19757);
nand U20090 (N_20090,N_19802,N_19848);
and U20091 (N_20091,N_19834,N_19910);
or U20092 (N_20092,N_19846,N_19933);
nor U20093 (N_20093,N_19871,N_19783);
or U20094 (N_20094,N_19969,N_19897);
nand U20095 (N_20095,N_19840,N_19806);
nor U20096 (N_20096,N_19954,N_19986);
nand U20097 (N_20097,N_19805,N_19966);
nand U20098 (N_20098,N_19797,N_19859);
and U20099 (N_20099,N_19804,N_19896);
nand U20100 (N_20100,N_19787,N_19957);
nor U20101 (N_20101,N_19963,N_19985);
nand U20102 (N_20102,N_19779,N_19940);
or U20103 (N_20103,N_19768,N_19758);
xor U20104 (N_20104,N_19792,N_19818);
nand U20105 (N_20105,N_19781,N_19952);
xnor U20106 (N_20106,N_19930,N_19997);
and U20107 (N_20107,N_19996,N_19955);
nor U20108 (N_20108,N_19790,N_19826);
and U20109 (N_20109,N_19831,N_19988);
nand U20110 (N_20110,N_19812,N_19915);
xor U20111 (N_20111,N_19946,N_19873);
xnor U20112 (N_20112,N_19785,N_19935);
and U20113 (N_20113,N_19795,N_19892);
or U20114 (N_20114,N_19777,N_19852);
or U20115 (N_20115,N_19809,N_19905);
nand U20116 (N_20116,N_19837,N_19853);
nand U20117 (N_20117,N_19998,N_19851);
xor U20118 (N_20118,N_19981,N_19931);
nor U20119 (N_20119,N_19762,N_19801);
and U20120 (N_20120,N_19819,N_19817);
xnor U20121 (N_20121,N_19772,N_19813);
xnor U20122 (N_20122,N_19776,N_19816);
or U20123 (N_20123,N_19775,N_19756);
nor U20124 (N_20124,N_19894,N_19794);
nor U20125 (N_20125,N_19936,N_19975);
nor U20126 (N_20126,N_19787,N_19859);
nor U20127 (N_20127,N_19964,N_19935);
or U20128 (N_20128,N_19859,N_19807);
xor U20129 (N_20129,N_19907,N_19990);
nor U20130 (N_20130,N_19961,N_19752);
xnor U20131 (N_20131,N_19915,N_19966);
nand U20132 (N_20132,N_19821,N_19789);
nor U20133 (N_20133,N_19778,N_19839);
xor U20134 (N_20134,N_19833,N_19766);
xor U20135 (N_20135,N_19782,N_19788);
nor U20136 (N_20136,N_19915,N_19873);
nand U20137 (N_20137,N_19962,N_19838);
nor U20138 (N_20138,N_19928,N_19791);
xnor U20139 (N_20139,N_19810,N_19829);
and U20140 (N_20140,N_19892,N_19946);
or U20141 (N_20141,N_19959,N_19881);
or U20142 (N_20142,N_19941,N_19795);
xnor U20143 (N_20143,N_19800,N_19932);
or U20144 (N_20144,N_19795,N_19769);
nor U20145 (N_20145,N_19986,N_19845);
and U20146 (N_20146,N_19824,N_19858);
nand U20147 (N_20147,N_19794,N_19882);
nand U20148 (N_20148,N_19958,N_19947);
nand U20149 (N_20149,N_19910,N_19780);
and U20150 (N_20150,N_19986,N_19938);
xor U20151 (N_20151,N_19923,N_19882);
or U20152 (N_20152,N_19916,N_19955);
and U20153 (N_20153,N_19931,N_19810);
or U20154 (N_20154,N_19901,N_19771);
and U20155 (N_20155,N_19904,N_19869);
xnor U20156 (N_20156,N_19806,N_19872);
and U20157 (N_20157,N_19800,N_19914);
nor U20158 (N_20158,N_19811,N_19931);
xnor U20159 (N_20159,N_19838,N_19869);
nand U20160 (N_20160,N_19856,N_19876);
and U20161 (N_20161,N_19759,N_19966);
nor U20162 (N_20162,N_19954,N_19867);
and U20163 (N_20163,N_19785,N_19854);
or U20164 (N_20164,N_19828,N_19771);
and U20165 (N_20165,N_19834,N_19856);
nor U20166 (N_20166,N_19987,N_19833);
and U20167 (N_20167,N_19979,N_19968);
nor U20168 (N_20168,N_19998,N_19844);
nor U20169 (N_20169,N_19926,N_19822);
nor U20170 (N_20170,N_19893,N_19864);
xnor U20171 (N_20171,N_19879,N_19973);
nand U20172 (N_20172,N_19836,N_19770);
xnor U20173 (N_20173,N_19878,N_19931);
and U20174 (N_20174,N_19889,N_19936);
nor U20175 (N_20175,N_19851,N_19752);
and U20176 (N_20176,N_19975,N_19958);
or U20177 (N_20177,N_19984,N_19859);
nand U20178 (N_20178,N_19836,N_19787);
nor U20179 (N_20179,N_19796,N_19882);
and U20180 (N_20180,N_19889,N_19918);
and U20181 (N_20181,N_19872,N_19927);
and U20182 (N_20182,N_19949,N_19756);
xnor U20183 (N_20183,N_19862,N_19934);
nor U20184 (N_20184,N_19941,N_19770);
xnor U20185 (N_20185,N_19900,N_19982);
nor U20186 (N_20186,N_19882,N_19837);
xnor U20187 (N_20187,N_19909,N_19762);
xnor U20188 (N_20188,N_19817,N_19906);
nor U20189 (N_20189,N_19901,N_19864);
or U20190 (N_20190,N_19859,N_19973);
nor U20191 (N_20191,N_19995,N_19910);
nand U20192 (N_20192,N_19858,N_19759);
nor U20193 (N_20193,N_19998,N_19761);
or U20194 (N_20194,N_19913,N_19814);
xnor U20195 (N_20195,N_19942,N_19978);
xor U20196 (N_20196,N_19843,N_19963);
nand U20197 (N_20197,N_19901,N_19998);
xor U20198 (N_20198,N_19950,N_19777);
xor U20199 (N_20199,N_19832,N_19812);
or U20200 (N_20200,N_19824,N_19789);
nand U20201 (N_20201,N_19802,N_19796);
nor U20202 (N_20202,N_19854,N_19884);
nor U20203 (N_20203,N_19864,N_19854);
and U20204 (N_20204,N_19887,N_19982);
nor U20205 (N_20205,N_19960,N_19890);
nor U20206 (N_20206,N_19984,N_19994);
and U20207 (N_20207,N_19892,N_19783);
and U20208 (N_20208,N_19877,N_19869);
nor U20209 (N_20209,N_19860,N_19910);
and U20210 (N_20210,N_19997,N_19896);
xnor U20211 (N_20211,N_19872,N_19945);
or U20212 (N_20212,N_19794,N_19834);
or U20213 (N_20213,N_19995,N_19868);
nor U20214 (N_20214,N_19985,N_19994);
xnor U20215 (N_20215,N_19878,N_19907);
xnor U20216 (N_20216,N_19827,N_19779);
xnor U20217 (N_20217,N_19967,N_19872);
nand U20218 (N_20218,N_19975,N_19950);
xnor U20219 (N_20219,N_19794,N_19792);
and U20220 (N_20220,N_19796,N_19858);
nor U20221 (N_20221,N_19953,N_19848);
and U20222 (N_20222,N_19780,N_19945);
and U20223 (N_20223,N_19837,N_19852);
nor U20224 (N_20224,N_19943,N_19788);
nor U20225 (N_20225,N_19917,N_19993);
or U20226 (N_20226,N_19781,N_19974);
and U20227 (N_20227,N_19757,N_19995);
and U20228 (N_20228,N_19979,N_19934);
nor U20229 (N_20229,N_19908,N_19989);
or U20230 (N_20230,N_19805,N_19943);
xor U20231 (N_20231,N_19889,N_19888);
or U20232 (N_20232,N_19782,N_19884);
nand U20233 (N_20233,N_19952,N_19910);
nor U20234 (N_20234,N_19888,N_19887);
xnor U20235 (N_20235,N_19756,N_19991);
and U20236 (N_20236,N_19754,N_19800);
nor U20237 (N_20237,N_19769,N_19934);
and U20238 (N_20238,N_19955,N_19920);
xnor U20239 (N_20239,N_19903,N_19918);
nand U20240 (N_20240,N_19780,N_19873);
xor U20241 (N_20241,N_19808,N_19962);
nor U20242 (N_20242,N_19825,N_19775);
xnor U20243 (N_20243,N_19922,N_19775);
nand U20244 (N_20244,N_19811,N_19767);
and U20245 (N_20245,N_19931,N_19801);
or U20246 (N_20246,N_19886,N_19928);
xnor U20247 (N_20247,N_19853,N_19859);
or U20248 (N_20248,N_19815,N_19770);
nand U20249 (N_20249,N_19778,N_19823);
xor U20250 (N_20250,N_20128,N_20131);
xor U20251 (N_20251,N_20162,N_20170);
and U20252 (N_20252,N_20025,N_20217);
xnor U20253 (N_20253,N_20068,N_20235);
nor U20254 (N_20254,N_20148,N_20090);
and U20255 (N_20255,N_20231,N_20006);
and U20256 (N_20256,N_20163,N_20151);
nor U20257 (N_20257,N_20175,N_20165);
xor U20258 (N_20258,N_20112,N_20042);
nand U20259 (N_20259,N_20249,N_20184);
or U20260 (N_20260,N_20176,N_20041);
nand U20261 (N_20261,N_20153,N_20071);
nor U20262 (N_20262,N_20152,N_20023);
nor U20263 (N_20263,N_20186,N_20208);
or U20264 (N_20264,N_20237,N_20204);
xnor U20265 (N_20265,N_20066,N_20030);
or U20266 (N_20266,N_20027,N_20138);
nand U20267 (N_20267,N_20196,N_20088);
and U20268 (N_20268,N_20024,N_20069);
nand U20269 (N_20269,N_20084,N_20062);
nand U20270 (N_20270,N_20244,N_20040);
xnor U20271 (N_20271,N_20100,N_20218);
or U20272 (N_20272,N_20082,N_20233);
xor U20273 (N_20273,N_20242,N_20117);
nor U20274 (N_20274,N_20192,N_20081);
and U20275 (N_20275,N_20166,N_20180);
nor U20276 (N_20276,N_20094,N_20076);
nor U20277 (N_20277,N_20188,N_20241);
nor U20278 (N_20278,N_20055,N_20164);
nand U20279 (N_20279,N_20190,N_20087);
nor U20280 (N_20280,N_20109,N_20183);
or U20281 (N_20281,N_20048,N_20239);
nand U20282 (N_20282,N_20209,N_20141);
or U20283 (N_20283,N_20020,N_20009);
or U20284 (N_20284,N_20095,N_20168);
nor U20285 (N_20285,N_20125,N_20135);
or U20286 (N_20286,N_20116,N_20223);
or U20287 (N_20287,N_20245,N_20072);
xnor U20288 (N_20288,N_20182,N_20104);
nand U20289 (N_20289,N_20248,N_20043);
and U20290 (N_20290,N_20015,N_20139);
or U20291 (N_20291,N_20010,N_20086);
and U20292 (N_20292,N_20220,N_20181);
nand U20293 (N_20293,N_20002,N_20097);
nor U20294 (N_20294,N_20103,N_20063);
or U20295 (N_20295,N_20017,N_20227);
xnor U20296 (N_20296,N_20101,N_20222);
or U20297 (N_20297,N_20124,N_20083);
nor U20298 (N_20298,N_20193,N_20021);
or U20299 (N_20299,N_20102,N_20078);
nor U20300 (N_20300,N_20026,N_20126);
and U20301 (N_20301,N_20107,N_20234);
nor U20302 (N_20302,N_20130,N_20098);
or U20303 (N_20303,N_20140,N_20001);
xor U20304 (N_20304,N_20212,N_20099);
nand U20305 (N_20305,N_20174,N_20127);
or U20306 (N_20306,N_20045,N_20047);
or U20307 (N_20307,N_20123,N_20214);
xor U20308 (N_20308,N_20079,N_20177);
and U20309 (N_20309,N_20089,N_20169);
nor U20310 (N_20310,N_20018,N_20207);
or U20311 (N_20311,N_20160,N_20122);
nor U20312 (N_20312,N_20014,N_20247);
nand U20313 (N_20313,N_20199,N_20167);
and U20314 (N_20314,N_20155,N_20016);
and U20315 (N_20315,N_20110,N_20051);
xor U20316 (N_20316,N_20120,N_20039);
nand U20317 (N_20317,N_20011,N_20229);
and U20318 (N_20318,N_20058,N_20203);
nor U20319 (N_20319,N_20065,N_20156);
nand U20320 (N_20320,N_20022,N_20114);
and U20321 (N_20321,N_20224,N_20201);
nand U20322 (N_20322,N_20050,N_20035);
nand U20323 (N_20323,N_20154,N_20119);
nor U20324 (N_20324,N_20205,N_20198);
and U20325 (N_20325,N_20173,N_20061);
and U20326 (N_20326,N_20206,N_20004);
or U20327 (N_20327,N_20032,N_20054);
nand U20328 (N_20328,N_20129,N_20056);
nor U20329 (N_20329,N_20044,N_20092);
or U20330 (N_20330,N_20115,N_20143);
and U20331 (N_20331,N_20106,N_20142);
nor U20332 (N_20332,N_20105,N_20019);
nand U20333 (N_20333,N_20093,N_20091);
xor U20334 (N_20334,N_20221,N_20028);
or U20335 (N_20335,N_20064,N_20194);
nor U20336 (N_20336,N_20159,N_20074);
xnor U20337 (N_20337,N_20226,N_20200);
xnor U20338 (N_20338,N_20232,N_20236);
xor U20339 (N_20339,N_20118,N_20243);
nor U20340 (N_20340,N_20073,N_20185);
nor U20341 (N_20341,N_20070,N_20178);
nand U20342 (N_20342,N_20003,N_20172);
xnor U20343 (N_20343,N_20219,N_20147);
nand U20344 (N_20344,N_20033,N_20060);
nand U20345 (N_20345,N_20228,N_20034);
or U20346 (N_20346,N_20080,N_20057);
xor U20347 (N_20347,N_20195,N_20007);
nor U20348 (N_20348,N_20049,N_20132);
nand U20349 (N_20349,N_20171,N_20150);
and U20350 (N_20350,N_20113,N_20246);
nand U20351 (N_20351,N_20053,N_20036);
or U20352 (N_20352,N_20213,N_20029);
or U20353 (N_20353,N_20075,N_20096);
nand U20354 (N_20354,N_20077,N_20038);
xor U20355 (N_20355,N_20179,N_20157);
and U20356 (N_20356,N_20216,N_20189);
nor U20357 (N_20357,N_20013,N_20210);
and U20358 (N_20358,N_20134,N_20225);
or U20359 (N_20359,N_20145,N_20085);
nor U20360 (N_20360,N_20144,N_20052);
nand U20361 (N_20361,N_20108,N_20067);
xnor U20362 (N_20362,N_20037,N_20000);
nor U20363 (N_20363,N_20137,N_20046);
nor U20364 (N_20364,N_20158,N_20211);
xnor U20365 (N_20365,N_20059,N_20187);
nor U20366 (N_20366,N_20111,N_20191);
nor U20367 (N_20367,N_20197,N_20136);
and U20368 (N_20368,N_20240,N_20005);
nand U20369 (N_20369,N_20146,N_20121);
nor U20370 (N_20370,N_20230,N_20202);
or U20371 (N_20371,N_20215,N_20238);
and U20372 (N_20372,N_20161,N_20031);
nor U20373 (N_20373,N_20008,N_20133);
nor U20374 (N_20374,N_20012,N_20149);
and U20375 (N_20375,N_20033,N_20164);
or U20376 (N_20376,N_20229,N_20228);
nand U20377 (N_20377,N_20202,N_20078);
nand U20378 (N_20378,N_20182,N_20016);
nand U20379 (N_20379,N_20206,N_20061);
nand U20380 (N_20380,N_20051,N_20118);
xnor U20381 (N_20381,N_20109,N_20002);
nand U20382 (N_20382,N_20180,N_20104);
or U20383 (N_20383,N_20113,N_20221);
nor U20384 (N_20384,N_20159,N_20061);
xor U20385 (N_20385,N_20053,N_20108);
and U20386 (N_20386,N_20106,N_20040);
or U20387 (N_20387,N_20221,N_20204);
and U20388 (N_20388,N_20117,N_20194);
and U20389 (N_20389,N_20136,N_20161);
nand U20390 (N_20390,N_20105,N_20215);
xnor U20391 (N_20391,N_20137,N_20051);
and U20392 (N_20392,N_20051,N_20045);
or U20393 (N_20393,N_20039,N_20089);
and U20394 (N_20394,N_20033,N_20027);
and U20395 (N_20395,N_20119,N_20093);
nand U20396 (N_20396,N_20211,N_20249);
nand U20397 (N_20397,N_20179,N_20232);
nand U20398 (N_20398,N_20210,N_20178);
nor U20399 (N_20399,N_20050,N_20058);
nand U20400 (N_20400,N_20177,N_20163);
xnor U20401 (N_20401,N_20072,N_20057);
and U20402 (N_20402,N_20105,N_20091);
xor U20403 (N_20403,N_20246,N_20082);
xor U20404 (N_20404,N_20055,N_20113);
nor U20405 (N_20405,N_20168,N_20197);
or U20406 (N_20406,N_20172,N_20229);
and U20407 (N_20407,N_20101,N_20147);
and U20408 (N_20408,N_20051,N_20203);
and U20409 (N_20409,N_20238,N_20065);
and U20410 (N_20410,N_20136,N_20220);
xor U20411 (N_20411,N_20219,N_20188);
nor U20412 (N_20412,N_20223,N_20164);
nand U20413 (N_20413,N_20117,N_20207);
xor U20414 (N_20414,N_20244,N_20107);
nand U20415 (N_20415,N_20166,N_20200);
or U20416 (N_20416,N_20129,N_20221);
nor U20417 (N_20417,N_20082,N_20224);
or U20418 (N_20418,N_20149,N_20016);
xnor U20419 (N_20419,N_20136,N_20229);
and U20420 (N_20420,N_20018,N_20209);
xnor U20421 (N_20421,N_20140,N_20240);
xnor U20422 (N_20422,N_20248,N_20168);
xor U20423 (N_20423,N_20101,N_20148);
nand U20424 (N_20424,N_20007,N_20231);
or U20425 (N_20425,N_20184,N_20035);
or U20426 (N_20426,N_20020,N_20210);
nor U20427 (N_20427,N_20055,N_20019);
or U20428 (N_20428,N_20155,N_20160);
nor U20429 (N_20429,N_20035,N_20067);
nor U20430 (N_20430,N_20247,N_20057);
nand U20431 (N_20431,N_20086,N_20023);
and U20432 (N_20432,N_20026,N_20177);
xor U20433 (N_20433,N_20108,N_20145);
or U20434 (N_20434,N_20047,N_20033);
and U20435 (N_20435,N_20057,N_20032);
or U20436 (N_20436,N_20090,N_20062);
xnor U20437 (N_20437,N_20066,N_20195);
or U20438 (N_20438,N_20085,N_20137);
nand U20439 (N_20439,N_20069,N_20154);
and U20440 (N_20440,N_20184,N_20089);
or U20441 (N_20441,N_20066,N_20060);
nor U20442 (N_20442,N_20133,N_20196);
or U20443 (N_20443,N_20077,N_20123);
nand U20444 (N_20444,N_20199,N_20149);
nor U20445 (N_20445,N_20142,N_20030);
nand U20446 (N_20446,N_20129,N_20009);
xnor U20447 (N_20447,N_20194,N_20172);
xor U20448 (N_20448,N_20083,N_20160);
nor U20449 (N_20449,N_20147,N_20141);
xnor U20450 (N_20450,N_20111,N_20016);
nand U20451 (N_20451,N_20009,N_20194);
and U20452 (N_20452,N_20116,N_20195);
or U20453 (N_20453,N_20063,N_20231);
or U20454 (N_20454,N_20113,N_20179);
nand U20455 (N_20455,N_20156,N_20138);
or U20456 (N_20456,N_20235,N_20012);
nor U20457 (N_20457,N_20183,N_20075);
nor U20458 (N_20458,N_20120,N_20203);
and U20459 (N_20459,N_20035,N_20039);
xor U20460 (N_20460,N_20235,N_20159);
nor U20461 (N_20461,N_20194,N_20170);
or U20462 (N_20462,N_20245,N_20052);
or U20463 (N_20463,N_20198,N_20094);
nand U20464 (N_20464,N_20004,N_20105);
nand U20465 (N_20465,N_20202,N_20040);
xnor U20466 (N_20466,N_20189,N_20051);
and U20467 (N_20467,N_20094,N_20058);
nand U20468 (N_20468,N_20115,N_20011);
xnor U20469 (N_20469,N_20080,N_20202);
xnor U20470 (N_20470,N_20001,N_20061);
nand U20471 (N_20471,N_20183,N_20135);
xnor U20472 (N_20472,N_20196,N_20229);
nor U20473 (N_20473,N_20071,N_20075);
and U20474 (N_20474,N_20183,N_20066);
nor U20475 (N_20475,N_20233,N_20130);
xnor U20476 (N_20476,N_20101,N_20004);
nand U20477 (N_20477,N_20144,N_20126);
nor U20478 (N_20478,N_20017,N_20059);
xor U20479 (N_20479,N_20138,N_20043);
nand U20480 (N_20480,N_20041,N_20214);
and U20481 (N_20481,N_20070,N_20087);
or U20482 (N_20482,N_20074,N_20020);
nor U20483 (N_20483,N_20161,N_20192);
or U20484 (N_20484,N_20189,N_20026);
nand U20485 (N_20485,N_20117,N_20132);
xnor U20486 (N_20486,N_20246,N_20017);
and U20487 (N_20487,N_20039,N_20101);
xnor U20488 (N_20488,N_20215,N_20081);
nor U20489 (N_20489,N_20161,N_20169);
nor U20490 (N_20490,N_20124,N_20120);
or U20491 (N_20491,N_20242,N_20075);
nand U20492 (N_20492,N_20079,N_20119);
xor U20493 (N_20493,N_20206,N_20005);
or U20494 (N_20494,N_20208,N_20054);
or U20495 (N_20495,N_20066,N_20096);
nand U20496 (N_20496,N_20062,N_20076);
nand U20497 (N_20497,N_20025,N_20006);
nand U20498 (N_20498,N_20062,N_20068);
nor U20499 (N_20499,N_20062,N_20031);
and U20500 (N_20500,N_20315,N_20471);
and U20501 (N_20501,N_20383,N_20438);
and U20502 (N_20502,N_20370,N_20489);
xor U20503 (N_20503,N_20340,N_20285);
nor U20504 (N_20504,N_20412,N_20354);
xor U20505 (N_20505,N_20333,N_20452);
nand U20506 (N_20506,N_20373,N_20433);
xor U20507 (N_20507,N_20422,N_20280);
xor U20508 (N_20508,N_20446,N_20368);
and U20509 (N_20509,N_20402,N_20345);
or U20510 (N_20510,N_20485,N_20481);
nand U20511 (N_20511,N_20398,N_20392);
xor U20512 (N_20512,N_20273,N_20427);
and U20513 (N_20513,N_20428,N_20288);
or U20514 (N_20514,N_20305,N_20444);
or U20515 (N_20515,N_20498,N_20302);
and U20516 (N_20516,N_20282,N_20351);
nand U20517 (N_20517,N_20419,N_20350);
nand U20518 (N_20518,N_20355,N_20366);
nand U20519 (N_20519,N_20358,N_20429);
nor U20520 (N_20520,N_20272,N_20296);
nand U20521 (N_20521,N_20294,N_20318);
nor U20522 (N_20522,N_20352,N_20304);
nor U20523 (N_20523,N_20455,N_20321);
nand U20524 (N_20524,N_20406,N_20307);
nor U20525 (N_20525,N_20382,N_20411);
nor U20526 (N_20526,N_20258,N_20363);
and U20527 (N_20527,N_20461,N_20330);
nand U20528 (N_20528,N_20401,N_20483);
xor U20529 (N_20529,N_20391,N_20484);
xor U20530 (N_20530,N_20448,N_20323);
or U20531 (N_20531,N_20450,N_20343);
and U20532 (N_20532,N_20314,N_20408);
nand U20533 (N_20533,N_20460,N_20442);
nand U20534 (N_20534,N_20393,N_20454);
nand U20535 (N_20535,N_20365,N_20329);
and U20536 (N_20536,N_20413,N_20265);
nor U20537 (N_20537,N_20387,N_20259);
or U20538 (N_20538,N_20492,N_20451);
and U20539 (N_20539,N_20468,N_20381);
xor U20540 (N_20540,N_20263,N_20289);
xor U20541 (N_20541,N_20431,N_20415);
nor U20542 (N_20542,N_20439,N_20332);
nor U20543 (N_20543,N_20339,N_20430);
or U20544 (N_20544,N_20371,N_20287);
nand U20545 (N_20545,N_20399,N_20449);
nor U20546 (N_20546,N_20486,N_20416);
nor U20547 (N_20547,N_20327,N_20286);
nand U20548 (N_20548,N_20317,N_20361);
nor U20549 (N_20549,N_20303,N_20478);
and U20550 (N_20550,N_20487,N_20293);
or U20551 (N_20551,N_20308,N_20414);
and U20552 (N_20552,N_20338,N_20322);
and U20553 (N_20553,N_20277,N_20300);
and U20554 (N_20554,N_20497,N_20270);
or U20555 (N_20555,N_20385,N_20341);
and U20556 (N_20556,N_20326,N_20477);
nor U20557 (N_20557,N_20281,N_20283);
xor U20558 (N_20558,N_20337,N_20466);
nor U20559 (N_20559,N_20336,N_20469);
nand U20560 (N_20560,N_20292,N_20476);
nor U20561 (N_20561,N_20475,N_20377);
and U20562 (N_20562,N_20331,N_20251);
nand U20563 (N_20563,N_20395,N_20284);
xnor U20564 (N_20564,N_20253,N_20491);
nand U20565 (N_20565,N_20276,N_20313);
nand U20566 (N_20566,N_20353,N_20496);
and U20567 (N_20567,N_20495,N_20325);
xnor U20568 (N_20568,N_20360,N_20260);
nor U20569 (N_20569,N_20311,N_20403);
xnor U20570 (N_20570,N_20278,N_20410);
and U20571 (N_20571,N_20424,N_20290);
nor U20572 (N_20572,N_20378,N_20320);
nor U20573 (N_20573,N_20407,N_20390);
and U20574 (N_20574,N_20261,N_20254);
nand U20575 (N_20575,N_20369,N_20324);
and U20576 (N_20576,N_20462,N_20264);
nand U20577 (N_20577,N_20342,N_20372);
and U20578 (N_20578,N_20375,N_20463);
or U20579 (N_20579,N_20490,N_20295);
nand U20580 (N_20580,N_20328,N_20376);
or U20581 (N_20581,N_20423,N_20473);
and U20582 (N_20582,N_20275,N_20405);
and U20583 (N_20583,N_20456,N_20291);
or U20584 (N_20584,N_20386,N_20379);
and U20585 (N_20585,N_20384,N_20432);
or U20586 (N_20586,N_20364,N_20397);
nand U20587 (N_20587,N_20488,N_20359);
or U20588 (N_20588,N_20362,N_20297);
nand U20589 (N_20589,N_20301,N_20479);
nor U20590 (N_20590,N_20480,N_20396);
or U20591 (N_20591,N_20453,N_20348);
and U20592 (N_20592,N_20316,N_20306);
and U20593 (N_20593,N_20472,N_20404);
nor U20594 (N_20594,N_20458,N_20445);
or U20595 (N_20595,N_20389,N_20310);
xor U20596 (N_20596,N_20279,N_20426);
or U20597 (N_20597,N_20447,N_20349);
nand U20598 (N_20598,N_20367,N_20257);
xnor U20599 (N_20599,N_20356,N_20465);
or U20600 (N_20600,N_20299,N_20274);
or U20601 (N_20601,N_20464,N_20418);
nand U20602 (N_20602,N_20417,N_20437);
or U20603 (N_20603,N_20268,N_20319);
or U20604 (N_20604,N_20436,N_20309);
nand U20605 (N_20605,N_20443,N_20357);
nand U20606 (N_20606,N_20420,N_20425);
nand U20607 (N_20607,N_20346,N_20380);
nor U20608 (N_20608,N_20334,N_20344);
nor U20609 (N_20609,N_20266,N_20482);
nor U20610 (N_20610,N_20298,N_20493);
nand U20611 (N_20611,N_20250,N_20269);
or U20612 (N_20612,N_20494,N_20347);
and U20613 (N_20613,N_20374,N_20267);
or U20614 (N_20614,N_20335,N_20474);
and U20615 (N_20615,N_20388,N_20400);
nor U20616 (N_20616,N_20262,N_20421);
nor U20617 (N_20617,N_20409,N_20499);
nor U20618 (N_20618,N_20434,N_20467);
nand U20619 (N_20619,N_20394,N_20457);
nor U20620 (N_20620,N_20271,N_20435);
and U20621 (N_20621,N_20459,N_20312);
nor U20622 (N_20622,N_20256,N_20440);
xnor U20623 (N_20623,N_20441,N_20252);
nor U20624 (N_20624,N_20470,N_20255);
xor U20625 (N_20625,N_20258,N_20413);
nand U20626 (N_20626,N_20358,N_20455);
xor U20627 (N_20627,N_20424,N_20450);
xor U20628 (N_20628,N_20468,N_20409);
or U20629 (N_20629,N_20357,N_20450);
nand U20630 (N_20630,N_20459,N_20261);
and U20631 (N_20631,N_20313,N_20251);
xor U20632 (N_20632,N_20445,N_20333);
or U20633 (N_20633,N_20411,N_20488);
xor U20634 (N_20634,N_20323,N_20280);
xor U20635 (N_20635,N_20423,N_20277);
xor U20636 (N_20636,N_20462,N_20355);
nor U20637 (N_20637,N_20308,N_20302);
nor U20638 (N_20638,N_20474,N_20458);
nand U20639 (N_20639,N_20296,N_20465);
nor U20640 (N_20640,N_20497,N_20410);
nor U20641 (N_20641,N_20480,N_20331);
nor U20642 (N_20642,N_20499,N_20443);
and U20643 (N_20643,N_20444,N_20419);
nand U20644 (N_20644,N_20260,N_20406);
and U20645 (N_20645,N_20344,N_20349);
nor U20646 (N_20646,N_20485,N_20390);
xor U20647 (N_20647,N_20290,N_20473);
xnor U20648 (N_20648,N_20409,N_20394);
nor U20649 (N_20649,N_20443,N_20347);
xor U20650 (N_20650,N_20440,N_20273);
nand U20651 (N_20651,N_20398,N_20285);
nand U20652 (N_20652,N_20485,N_20300);
nand U20653 (N_20653,N_20298,N_20404);
and U20654 (N_20654,N_20424,N_20390);
nand U20655 (N_20655,N_20471,N_20257);
nor U20656 (N_20656,N_20372,N_20263);
xnor U20657 (N_20657,N_20318,N_20390);
nor U20658 (N_20658,N_20475,N_20434);
nor U20659 (N_20659,N_20359,N_20276);
or U20660 (N_20660,N_20351,N_20403);
and U20661 (N_20661,N_20428,N_20449);
nand U20662 (N_20662,N_20401,N_20315);
nand U20663 (N_20663,N_20251,N_20365);
nor U20664 (N_20664,N_20301,N_20414);
and U20665 (N_20665,N_20429,N_20323);
and U20666 (N_20666,N_20307,N_20453);
xor U20667 (N_20667,N_20434,N_20288);
nand U20668 (N_20668,N_20324,N_20430);
nor U20669 (N_20669,N_20470,N_20254);
and U20670 (N_20670,N_20256,N_20296);
and U20671 (N_20671,N_20367,N_20354);
and U20672 (N_20672,N_20461,N_20417);
or U20673 (N_20673,N_20354,N_20379);
nor U20674 (N_20674,N_20422,N_20411);
xnor U20675 (N_20675,N_20444,N_20353);
or U20676 (N_20676,N_20252,N_20254);
nor U20677 (N_20677,N_20383,N_20445);
and U20678 (N_20678,N_20476,N_20475);
nand U20679 (N_20679,N_20442,N_20392);
and U20680 (N_20680,N_20456,N_20252);
and U20681 (N_20681,N_20328,N_20304);
xor U20682 (N_20682,N_20351,N_20425);
and U20683 (N_20683,N_20314,N_20456);
or U20684 (N_20684,N_20406,N_20379);
nor U20685 (N_20685,N_20467,N_20256);
xor U20686 (N_20686,N_20426,N_20479);
nand U20687 (N_20687,N_20470,N_20276);
and U20688 (N_20688,N_20441,N_20271);
nor U20689 (N_20689,N_20442,N_20323);
nand U20690 (N_20690,N_20396,N_20392);
xnor U20691 (N_20691,N_20322,N_20370);
nor U20692 (N_20692,N_20482,N_20488);
nand U20693 (N_20693,N_20372,N_20468);
nor U20694 (N_20694,N_20448,N_20256);
nor U20695 (N_20695,N_20267,N_20472);
nand U20696 (N_20696,N_20486,N_20384);
nor U20697 (N_20697,N_20377,N_20431);
and U20698 (N_20698,N_20425,N_20343);
xnor U20699 (N_20699,N_20377,N_20282);
nand U20700 (N_20700,N_20295,N_20383);
or U20701 (N_20701,N_20437,N_20422);
and U20702 (N_20702,N_20366,N_20276);
nor U20703 (N_20703,N_20314,N_20281);
xor U20704 (N_20704,N_20321,N_20328);
nand U20705 (N_20705,N_20267,N_20355);
nor U20706 (N_20706,N_20487,N_20305);
nand U20707 (N_20707,N_20328,N_20340);
or U20708 (N_20708,N_20332,N_20351);
or U20709 (N_20709,N_20497,N_20475);
and U20710 (N_20710,N_20488,N_20407);
nor U20711 (N_20711,N_20298,N_20358);
xor U20712 (N_20712,N_20412,N_20443);
and U20713 (N_20713,N_20497,N_20499);
or U20714 (N_20714,N_20430,N_20361);
nor U20715 (N_20715,N_20328,N_20369);
and U20716 (N_20716,N_20464,N_20491);
or U20717 (N_20717,N_20454,N_20451);
nor U20718 (N_20718,N_20439,N_20409);
nand U20719 (N_20719,N_20359,N_20432);
nand U20720 (N_20720,N_20279,N_20380);
nand U20721 (N_20721,N_20365,N_20294);
and U20722 (N_20722,N_20270,N_20408);
nor U20723 (N_20723,N_20471,N_20287);
and U20724 (N_20724,N_20273,N_20296);
xnor U20725 (N_20725,N_20414,N_20378);
xor U20726 (N_20726,N_20306,N_20357);
nor U20727 (N_20727,N_20455,N_20275);
nor U20728 (N_20728,N_20451,N_20441);
and U20729 (N_20729,N_20314,N_20322);
nand U20730 (N_20730,N_20377,N_20427);
nand U20731 (N_20731,N_20263,N_20408);
xor U20732 (N_20732,N_20341,N_20297);
xnor U20733 (N_20733,N_20322,N_20451);
or U20734 (N_20734,N_20349,N_20413);
xnor U20735 (N_20735,N_20370,N_20499);
nor U20736 (N_20736,N_20467,N_20306);
nand U20737 (N_20737,N_20281,N_20300);
nand U20738 (N_20738,N_20411,N_20369);
and U20739 (N_20739,N_20295,N_20311);
nand U20740 (N_20740,N_20451,N_20468);
nand U20741 (N_20741,N_20251,N_20416);
or U20742 (N_20742,N_20373,N_20435);
xor U20743 (N_20743,N_20372,N_20472);
nand U20744 (N_20744,N_20292,N_20390);
xnor U20745 (N_20745,N_20460,N_20455);
nand U20746 (N_20746,N_20287,N_20273);
and U20747 (N_20747,N_20401,N_20419);
xor U20748 (N_20748,N_20455,N_20429);
xnor U20749 (N_20749,N_20275,N_20422);
nand U20750 (N_20750,N_20525,N_20631);
nor U20751 (N_20751,N_20502,N_20619);
nand U20752 (N_20752,N_20574,N_20583);
nor U20753 (N_20753,N_20522,N_20616);
or U20754 (N_20754,N_20708,N_20711);
xor U20755 (N_20755,N_20729,N_20604);
or U20756 (N_20756,N_20591,N_20548);
xnor U20757 (N_20757,N_20564,N_20713);
or U20758 (N_20758,N_20576,N_20733);
and U20759 (N_20759,N_20689,N_20568);
xor U20760 (N_20760,N_20683,N_20608);
xor U20761 (N_20761,N_20677,N_20510);
xor U20762 (N_20762,N_20722,N_20728);
nand U20763 (N_20763,N_20518,N_20503);
and U20764 (N_20764,N_20575,N_20546);
and U20765 (N_20765,N_20731,N_20526);
nand U20766 (N_20766,N_20530,N_20514);
nor U20767 (N_20767,N_20629,N_20587);
xnor U20768 (N_20768,N_20572,N_20664);
xor U20769 (N_20769,N_20688,N_20625);
and U20770 (N_20770,N_20584,N_20632);
xnor U20771 (N_20771,N_20519,N_20669);
nand U20772 (N_20772,N_20567,N_20709);
or U20773 (N_20773,N_20508,N_20638);
nor U20774 (N_20774,N_20714,N_20656);
and U20775 (N_20775,N_20734,N_20700);
nand U20776 (N_20776,N_20578,N_20727);
or U20777 (N_20777,N_20600,N_20555);
and U20778 (N_20778,N_20720,N_20529);
xnor U20779 (N_20779,N_20612,N_20739);
or U20780 (N_20780,N_20747,N_20630);
nand U20781 (N_20781,N_20624,N_20682);
or U20782 (N_20782,N_20540,N_20665);
nor U20783 (N_20783,N_20657,N_20699);
nor U20784 (N_20784,N_20618,N_20675);
and U20785 (N_20785,N_20660,N_20633);
nand U20786 (N_20786,N_20571,N_20609);
or U20787 (N_20787,N_20653,N_20539);
nand U20788 (N_20788,N_20563,N_20511);
nand U20789 (N_20789,N_20640,N_20698);
or U20790 (N_20790,N_20570,N_20593);
nand U20791 (N_20791,N_20556,N_20687);
or U20792 (N_20792,N_20562,N_20533);
nor U20793 (N_20793,N_20644,N_20706);
nor U20794 (N_20794,N_20697,N_20643);
xnor U20795 (N_20795,N_20686,N_20520);
nand U20796 (N_20796,N_20691,N_20500);
nand U20797 (N_20797,N_20627,N_20634);
nor U20798 (N_20798,N_20521,N_20719);
or U20799 (N_20799,N_20703,N_20573);
nand U20800 (N_20800,N_20726,N_20534);
xor U20801 (N_20801,N_20599,N_20553);
nor U20802 (N_20802,N_20702,N_20647);
and U20803 (N_20803,N_20628,N_20531);
nor U20804 (N_20804,N_20552,N_20679);
and U20805 (N_20805,N_20580,N_20651);
xnor U20806 (N_20806,N_20749,N_20527);
nand U20807 (N_20807,N_20672,N_20725);
xor U20808 (N_20808,N_20549,N_20673);
nand U20809 (N_20809,N_20622,N_20695);
or U20810 (N_20810,N_20742,N_20565);
nor U20811 (N_20811,N_20605,N_20545);
or U20812 (N_20812,N_20586,N_20501);
or U20813 (N_20813,N_20732,N_20707);
and U20814 (N_20814,N_20559,N_20504);
nor U20815 (N_20815,N_20694,N_20717);
nand U20816 (N_20816,N_20715,N_20606);
or U20817 (N_20817,N_20512,N_20537);
and U20818 (N_20818,N_20551,N_20577);
nand U20819 (N_20819,N_20560,N_20692);
nor U20820 (N_20820,N_20614,N_20582);
nor U20821 (N_20821,N_20536,N_20646);
nand U20822 (N_20822,N_20649,N_20636);
or U20823 (N_20823,N_20507,N_20671);
nor U20824 (N_20824,N_20650,N_20718);
xnor U20825 (N_20825,N_20685,N_20613);
nor U20826 (N_20826,N_20566,N_20513);
nor U20827 (N_20827,N_20524,N_20641);
xnor U20828 (N_20828,N_20617,N_20595);
or U20829 (N_20829,N_20710,N_20743);
or U20830 (N_20830,N_20645,N_20741);
or U20831 (N_20831,N_20542,N_20561);
nor U20832 (N_20832,N_20547,N_20523);
nor U20833 (N_20833,N_20544,N_20611);
nand U20834 (N_20834,N_20541,N_20598);
xor U20835 (N_20835,N_20745,N_20658);
nor U20836 (N_20836,N_20670,N_20588);
and U20837 (N_20837,N_20648,N_20661);
nor U20838 (N_20838,N_20602,N_20610);
xnor U20839 (N_20839,N_20626,N_20620);
nand U20840 (N_20840,N_20737,N_20678);
xor U20841 (N_20841,N_20736,N_20723);
nand U20842 (N_20842,N_20659,N_20738);
xnor U20843 (N_20843,N_20676,N_20596);
or U20844 (N_20844,N_20594,N_20538);
and U20845 (N_20845,N_20554,N_20696);
xnor U20846 (N_20846,N_20607,N_20693);
and U20847 (N_20847,N_20704,N_20581);
nor U20848 (N_20848,N_20667,N_20558);
xnor U20849 (N_20849,N_20516,N_20623);
and U20850 (N_20850,N_20666,N_20579);
xnor U20851 (N_20851,N_20505,N_20642);
or U20852 (N_20852,N_20712,N_20615);
xor U20853 (N_20853,N_20601,N_20621);
nor U20854 (N_20854,N_20674,N_20730);
xor U20855 (N_20855,N_20663,N_20681);
and U20856 (N_20856,N_20744,N_20690);
nand U20857 (N_20857,N_20535,N_20517);
and U20858 (N_20858,N_20635,N_20637);
nand U20859 (N_20859,N_20662,N_20589);
xor U20860 (N_20860,N_20701,N_20532);
nor U20861 (N_20861,N_20569,N_20585);
or U20862 (N_20862,N_20705,N_20740);
and U20863 (N_20863,N_20724,N_20509);
xnor U20864 (N_20864,N_20654,N_20515);
and U20865 (N_20865,N_20735,N_20655);
or U20866 (N_20866,N_20592,N_20639);
or U20867 (N_20867,N_20716,N_20597);
xnor U20868 (N_20868,N_20550,N_20590);
nand U20869 (N_20869,N_20528,N_20746);
nor U20870 (N_20870,N_20721,N_20684);
or U20871 (N_20871,N_20748,N_20603);
or U20872 (N_20872,N_20668,N_20506);
nand U20873 (N_20873,N_20652,N_20680);
or U20874 (N_20874,N_20543,N_20557);
and U20875 (N_20875,N_20571,N_20649);
nand U20876 (N_20876,N_20730,N_20680);
or U20877 (N_20877,N_20609,N_20585);
nor U20878 (N_20878,N_20507,N_20589);
and U20879 (N_20879,N_20648,N_20512);
nor U20880 (N_20880,N_20713,N_20718);
or U20881 (N_20881,N_20680,N_20553);
nor U20882 (N_20882,N_20558,N_20503);
or U20883 (N_20883,N_20705,N_20742);
or U20884 (N_20884,N_20504,N_20669);
nor U20885 (N_20885,N_20628,N_20614);
or U20886 (N_20886,N_20665,N_20527);
or U20887 (N_20887,N_20703,N_20665);
nand U20888 (N_20888,N_20679,N_20519);
and U20889 (N_20889,N_20688,N_20540);
nand U20890 (N_20890,N_20583,N_20501);
nor U20891 (N_20891,N_20501,N_20743);
xor U20892 (N_20892,N_20576,N_20621);
nor U20893 (N_20893,N_20608,N_20517);
or U20894 (N_20894,N_20625,N_20504);
or U20895 (N_20895,N_20693,N_20547);
xor U20896 (N_20896,N_20545,N_20589);
nand U20897 (N_20897,N_20749,N_20551);
or U20898 (N_20898,N_20701,N_20565);
and U20899 (N_20899,N_20685,N_20616);
and U20900 (N_20900,N_20536,N_20709);
or U20901 (N_20901,N_20504,N_20566);
and U20902 (N_20902,N_20630,N_20599);
nand U20903 (N_20903,N_20692,N_20666);
xnor U20904 (N_20904,N_20734,N_20720);
and U20905 (N_20905,N_20581,N_20728);
nand U20906 (N_20906,N_20533,N_20699);
xnor U20907 (N_20907,N_20748,N_20584);
and U20908 (N_20908,N_20577,N_20649);
xnor U20909 (N_20909,N_20735,N_20683);
and U20910 (N_20910,N_20650,N_20658);
nor U20911 (N_20911,N_20601,N_20638);
nand U20912 (N_20912,N_20689,N_20744);
or U20913 (N_20913,N_20530,N_20596);
xnor U20914 (N_20914,N_20596,N_20621);
xor U20915 (N_20915,N_20582,N_20747);
xor U20916 (N_20916,N_20701,N_20633);
nand U20917 (N_20917,N_20712,N_20634);
nor U20918 (N_20918,N_20557,N_20598);
nand U20919 (N_20919,N_20647,N_20678);
nor U20920 (N_20920,N_20688,N_20549);
or U20921 (N_20921,N_20568,N_20642);
and U20922 (N_20922,N_20738,N_20663);
or U20923 (N_20923,N_20622,N_20556);
and U20924 (N_20924,N_20710,N_20634);
or U20925 (N_20925,N_20672,N_20588);
or U20926 (N_20926,N_20512,N_20735);
xnor U20927 (N_20927,N_20669,N_20700);
nor U20928 (N_20928,N_20577,N_20678);
nor U20929 (N_20929,N_20626,N_20629);
and U20930 (N_20930,N_20589,N_20639);
xor U20931 (N_20931,N_20673,N_20718);
nor U20932 (N_20932,N_20574,N_20611);
xnor U20933 (N_20933,N_20592,N_20667);
nand U20934 (N_20934,N_20536,N_20610);
nand U20935 (N_20935,N_20516,N_20584);
xor U20936 (N_20936,N_20591,N_20651);
and U20937 (N_20937,N_20686,N_20552);
nand U20938 (N_20938,N_20695,N_20578);
and U20939 (N_20939,N_20663,N_20615);
and U20940 (N_20940,N_20531,N_20625);
or U20941 (N_20941,N_20648,N_20645);
and U20942 (N_20942,N_20526,N_20654);
nor U20943 (N_20943,N_20648,N_20520);
or U20944 (N_20944,N_20621,N_20554);
or U20945 (N_20945,N_20731,N_20523);
nor U20946 (N_20946,N_20522,N_20637);
and U20947 (N_20947,N_20742,N_20616);
nor U20948 (N_20948,N_20526,N_20637);
nand U20949 (N_20949,N_20539,N_20585);
nor U20950 (N_20950,N_20598,N_20683);
xnor U20951 (N_20951,N_20553,N_20712);
nor U20952 (N_20952,N_20723,N_20634);
or U20953 (N_20953,N_20575,N_20667);
and U20954 (N_20954,N_20637,N_20669);
xor U20955 (N_20955,N_20694,N_20655);
and U20956 (N_20956,N_20560,N_20659);
or U20957 (N_20957,N_20545,N_20501);
nor U20958 (N_20958,N_20555,N_20645);
or U20959 (N_20959,N_20601,N_20555);
nand U20960 (N_20960,N_20634,N_20653);
or U20961 (N_20961,N_20636,N_20525);
nor U20962 (N_20962,N_20592,N_20532);
nand U20963 (N_20963,N_20688,N_20652);
or U20964 (N_20964,N_20673,N_20511);
xnor U20965 (N_20965,N_20715,N_20562);
nand U20966 (N_20966,N_20537,N_20543);
or U20967 (N_20967,N_20673,N_20748);
and U20968 (N_20968,N_20647,N_20641);
and U20969 (N_20969,N_20613,N_20569);
nor U20970 (N_20970,N_20501,N_20707);
nor U20971 (N_20971,N_20648,N_20545);
xnor U20972 (N_20972,N_20613,N_20712);
and U20973 (N_20973,N_20684,N_20572);
xnor U20974 (N_20974,N_20618,N_20636);
or U20975 (N_20975,N_20675,N_20629);
or U20976 (N_20976,N_20522,N_20604);
nor U20977 (N_20977,N_20695,N_20523);
and U20978 (N_20978,N_20563,N_20504);
nand U20979 (N_20979,N_20544,N_20614);
nor U20980 (N_20980,N_20512,N_20631);
nor U20981 (N_20981,N_20660,N_20631);
or U20982 (N_20982,N_20597,N_20543);
and U20983 (N_20983,N_20597,N_20590);
nor U20984 (N_20984,N_20602,N_20701);
nand U20985 (N_20985,N_20682,N_20508);
nor U20986 (N_20986,N_20613,N_20555);
xor U20987 (N_20987,N_20510,N_20507);
or U20988 (N_20988,N_20506,N_20674);
nand U20989 (N_20989,N_20738,N_20649);
nand U20990 (N_20990,N_20616,N_20677);
or U20991 (N_20991,N_20655,N_20558);
xnor U20992 (N_20992,N_20696,N_20730);
and U20993 (N_20993,N_20699,N_20706);
xor U20994 (N_20994,N_20691,N_20724);
nand U20995 (N_20995,N_20598,N_20700);
nand U20996 (N_20996,N_20667,N_20521);
or U20997 (N_20997,N_20630,N_20594);
and U20998 (N_20998,N_20732,N_20552);
nand U20999 (N_20999,N_20501,N_20515);
or U21000 (N_21000,N_20920,N_20826);
or U21001 (N_21001,N_20782,N_20815);
nor U21002 (N_21002,N_20936,N_20896);
xnor U21003 (N_21003,N_20950,N_20867);
and U21004 (N_21004,N_20821,N_20797);
and U21005 (N_21005,N_20956,N_20981);
or U21006 (N_21006,N_20959,N_20984);
and U21007 (N_21007,N_20757,N_20752);
and U21008 (N_21008,N_20758,N_20760);
nor U21009 (N_21009,N_20799,N_20775);
xor U21010 (N_21010,N_20913,N_20883);
nand U21011 (N_21011,N_20862,N_20873);
and U21012 (N_21012,N_20898,N_20790);
nor U21013 (N_21013,N_20804,N_20979);
and U21014 (N_21014,N_20992,N_20791);
or U21015 (N_21015,N_20814,N_20893);
nor U21016 (N_21016,N_20876,N_20845);
xor U21017 (N_21017,N_20940,N_20947);
nor U21018 (N_21018,N_20923,N_20832);
nand U21019 (N_21019,N_20864,N_20915);
and U21020 (N_21020,N_20994,N_20833);
and U21021 (N_21021,N_20967,N_20878);
and U21022 (N_21022,N_20753,N_20870);
and U21023 (N_21023,N_20925,N_20930);
and U21024 (N_21024,N_20769,N_20822);
and U21025 (N_21025,N_20991,N_20808);
and U21026 (N_21026,N_20951,N_20837);
or U21027 (N_21027,N_20813,N_20774);
xnor U21028 (N_21028,N_20820,N_20768);
or U21029 (N_21029,N_20839,N_20772);
nand U21030 (N_21030,N_20776,N_20996);
or U21031 (N_21031,N_20946,N_20969);
and U21032 (N_21032,N_20886,N_20773);
xor U21033 (N_21033,N_20871,N_20770);
and U21034 (N_21034,N_20942,N_20789);
nand U21035 (N_21035,N_20971,N_20835);
nand U21036 (N_21036,N_20840,N_20931);
nand U21037 (N_21037,N_20927,N_20847);
and U21038 (N_21038,N_20784,N_20918);
xnor U21039 (N_21039,N_20879,N_20882);
or U21040 (N_21040,N_20811,N_20787);
or U21041 (N_21041,N_20795,N_20766);
nand U21042 (N_21042,N_20894,N_20903);
and U21043 (N_21043,N_20812,N_20976);
nor U21044 (N_21044,N_20962,N_20911);
and U21045 (N_21045,N_20957,N_20777);
and U21046 (N_21046,N_20819,N_20954);
or U21047 (N_21047,N_20972,N_20924);
or U21048 (N_21048,N_20817,N_20858);
or U21049 (N_21049,N_20834,N_20836);
nor U21050 (N_21050,N_20934,N_20937);
xnor U21051 (N_21051,N_20868,N_20977);
or U21052 (N_21052,N_20852,N_20865);
and U21053 (N_21053,N_20751,N_20779);
and U21054 (N_21054,N_20892,N_20884);
and U21055 (N_21055,N_20881,N_20853);
and U21056 (N_21056,N_20802,N_20765);
xor U21057 (N_21057,N_20805,N_20974);
nand U21058 (N_21058,N_20831,N_20785);
xnor U21059 (N_21059,N_20818,N_20860);
xor U21060 (N_21060,N_20952,N_20889);
and U21061 (N_21061,N_20933,N_20935);
xor U21062 (N_21062,N_20857,N_20914);
nand U21063 (N_21063,N_20995,N_20961);
nand U21064 (N_21064,N_20960,N_20964);
or U21065 (N_21065,N_20949,N_20816);
or U21066 (N_21066,N_20999,N_20885);
or U21067 (N_21067,N_20978,N_20855);
xnor U21068 (N_21068,N_20922,N_20750);
nand U21069 (N_21069,N_20987,N_20910);
or U21070 (N_21070,N_20771,N_20803);
and U21071 (N_21071,N_20869,N_20921);
and U21072 (N_21072,N_20842,N_20912);
nor U21073 (N_21073,N_20943,N_20998);
xor U21074 (N_21074,N_20850,N_20788);
xnor U21075 (N_21075,N_20756,N_20783);
xnor U21076 (N_21076,N_20906,N_20989);
or U21077 (N_21077,N_20973,N_20899);
nor U21078 (N_21078,N_20926,N_20905);
and U21079 (N_21079,N_20843,N_20901);
and U21080 (N_21080,N_20844,N_20767);
nand U21081 (N_21081,N_20919,N_20908);
nand U21082 (N_21082,N_20948,N_20986);
nor U21083 (N_21083,N_20928,N_20807);
and U21084 (N_21084,N_20975,N_20966);
xor U21085 (N_21085,N_20970,N_20849);
xor U21086 (N_21086,N_20997,N_20793);
and U21087 (N_21087,N_20778,N_20988);
xnor U21088 (N_21088,N_20965,N_20780);
or U21089 (N_21089,N_20801,N_20982);
or U21090 (N_21090,N_20880,N_20866);
nor U21091 (N_21091,N_20755,N_20872);
and U21092 (N_21092,N_20848,N_20891);
nor U21093 (N_21093,N_20754,N_20929);
nor U21094 (N_21094,N_20796,N_20846);
nor U21095 (N_21095,N_20993,N_20904);
nor U21096 (N_21096,N_20888,N_20968);
and U21097 (N_21097,N_20897,N_20875);
xnor U21098 (N_21098,N_20762,N_20916);
and U21099 (N_21099,N_20945,N_20764);
and U21100 (N_21100,N_20809,N_20902);
nand U21101 (N_21101,N_20877,N_20786);
xor U21102 (N_21102,N_20985,N_20953);
nand U21103 (N_21103,N_20955,N_20941);
nand U21104 (N_21104,N_20823,N_20863);
nand U21105 (N_21105,N_20829,N_20990);
and U21106 (N_21106,N_20938,N_20854);
xor U21107 (N_21107,N_20830,N_20900);
xnor U21108 (N_21108,N_20824,N_20851);
xor U21109 (N_21109,N_20810,N_20963);
nor U21110 (N_21110,N_20794,N_20759);
nor U21111 (N_21111,N_20944,N_20983);
xor U21112 (N_21112,N_20874,N_20841);
nand U21113 (N_21113,N_20887,N_20798);
nand U21114 (N_21114,N_20907,N_20825);
xor U21115 (N_21115,N_20890,N_20761);
nor U21116 (N_21116,N_20932,N_20856);
or U21117 (N_21117,N_20895,N_20939);
xnor U21118 (N_21118,N_20838,N_20806);
xor U21119 (N_21119,N_20917,N_20859);
and U21120 (N_21120,N_20792,N_20763);
nor U21121 (N_21121,N_20800,N_20781);
or U21122 (N_21122,N_20828,N_20861);
xor U21123 (N_21123,N_20958,N_20909);
xor U21124 (N_21124,N_20980,N_20827);
and U21125 (N_21125,N_20777,N_20995);
xnor U21126 (N_21126,N_20975,N_20977);
nand U21127 (N_21127,N_20760,N_20926);
and U21128 (N_21128,N_20952,N_20929);
nand U21129 (N_21129,N_20976,N_20959);
xor U21130 (N_21130,N_20886,N_20842);
xor U21131 (N_21131,N_20846,N_20852);
or U21132 (N_21132,N_20765,N_20753);
and U21133 (N_21133,N_20829,N_20833);
xnor U21134 (N_21134,N_20874,N_20866);
or U21135 (N_21135,N_20880,N_20771);
nand U21136 (N_21136,N_20782,N_20970);
or U21137 (N_21137,N_20822,N_20772);
nand U21138 (N_21138,N_20971,N_20930);
or U21139 (N_21139,N_20787,N_20856);
or U21140 (N_21140,N_20849,N_20765);
xnor U21141 (N_21141,N_20964,N_20877);
and U21142 (N_21142,N_20976,N_20971);
nand U21143 (N_21143,N_20985,N_20810);
nand U21144 (N_21144,N_20967,N_20995);
nor U21145 (N_21145,N_20763,N_20769);
xor U21146 (N_21146,N_20936,N_20954);
and U21147 (N_21147,N_20964,N_20847);
xor U21148 (N_21148,N_20918,N_20945);
xnor U21149 (N_21149,N_20760,N_20985);
nor U21150 (N_21150,N_20828,N_20878);
nor U21151 (N_21151,N_20833,N_20818);
nor U21152 (N_21152,N_20797,N_20791);
nor U21153 (N_21153,N_20834,N_20900);
nand U21154 (N_21154,N_20892,N_20754);
or U21155 (N_21155,N_20838,N_20864);
or U21156 (N_21156,N_20862,N_20905);
nand U21157 (N_21157,N_20936,N_20803);
or U21158 (N_21158,N_20772,N_20939);
xor U21159 (N_21159,N_20857,N_20902);
or U21160 (N_21160,N_20823,N_20833);
or U21161 (N_21161,N_20917,N_20815);
nor U21162 (N_21162,N_20829,N_20864);
or U21163 (N_21163,N_20944,N_20938);
xor U21164 (N_21164,N_20784,N_20785);
xor U21165 (N_21165,N_20961,N_20814);
nor U21166 (N_21166,N_20754,N_20778);
nand U21167 (N_21167,N_20892,N_20966);
and U21168 (N_21168,N_20984,N_20808);
and U21169 (N_21169,N_20830,N_20813);
nand U21170 (N_21170,N_20790,N_20956);
or U21171 (N_21171,N_20844,N_20843);
xor U21172 (N_21172,N_20960,N_20906);
and U21173 (N_21173,N_20918,N_20973);
nand U21174 (N_21174,N_20907,N_20830);
nand U21175 (N_21175,N_20858,N_20828);
and U21176 (N_21176,N_20811,N_20800);
xor U21177 (N_21177,N_20769,N_20994);
xnor U21178 (N_21178,N_20960,N_20866);
or U21179 (N_21179,N_20883,N_20843);
xnor U21180 (N_21180,N_20875,N_20872);
and U21181 (N_21181,N_20752,N_20900);
nor U21182 (N_21182,N_20936,N_20915);
xor U21183 (N_21183,N_20828,N_20763);
and U21184 (N_21184,N_20971,N_20771);
nor U21185 (N_21185,N_20810,N_20750);
nor U21186 (N_21186,N_20910,N_20826);
nor U21187 (N_21187,N_20788,N_20761);
and U21188 (N_21188,N_20783,N_20981);
and U21189 (N_21189,N_20844,N_20896);
nor U21190 (N_21190,N_20806,N_20902);
nor U21191 (N_21191,N_20862,N_20808);
xor U21192 (N_21192,N_20896,N_20842);
nand U21193 (N_21193,N_20854,N_20999);
nand U21194 (N_21194,N_20893,N_20828);
nand U21195 (N_21195,N_20754,N_20840);
xnor U21196 (N_21196,N_20811,N_20937);
nor U21197 (N_21197,N_20750,N_20936);
xnor U21198 (N_21198,N_20883,N_20899);
and U21199 (N_21199,N_20945,N_20854);
nand U21200 (N_21200,N_20884,N_20957);
or U21201 (N_21201,N_20759,N_20892);
and U21202 (N_21202,N_20763,N_20864);
nor U21203 (N_21203,N_20751,N_20859);
xor U21204 (N_21204,N_20994,N_20921);
or U21205 (N_21205,N_20838,N_20891);
or U21206 (N_21206,N_20888,N_20949);
nor U21207 (N_21207,N_20887,N_20964);
and U21208 (N_21208,N_20985,N_20848);
or U21209 (N_21209,N_20872,N_20783);
and U21210 (N_21210,N_20770,N_20760);
nor U21211 (N_21211,N_20836,N_20919);
nor U21212 (N_21212,N_20969,N_20935);
or U21213 (N_21213,N_20934,N_20904);
nor U21214 (N_21214,N_20997,N_20990);
and U21215 (N_21215,N_20903,N_20772);
and U21216 (N_21216,N_20910,N_20915);
nand U21217 (N_21217,N_20994,N_20900);
nand U21218 (N_21218,N_20775,N_20925);
or U21219 (N_21219,N_20762,N_20807);
nor U21220 (N_21220,N_20900,N_20803);
nand U21221 (N_21221,N_20806,N_20932);
and U21222 (N_21222,N_20993,N_20903);
nand U21223 (N_21223,N_20992,N_20839);
nor U21224 (N_21224,N_20990,N_20888);
and U21225 (N_21225,N_20908,N_20962);
xor U21226 (N_21226,N_20875,N_20888);
and U21227 (N_21227,N_20971,N_20888);
nand U21228 (N_21228,N_20783,N_20806);
nand U21229 (N_21229,N_20808,N_20815);
xor U21230 (N_21230,N_20791,N_20854);
xor U21231 (N_21231,N_20979,N_20937);
or U21232 (N_21232,N_20900,N_20767);
xor U21233 (N_21233,N_20929,N_20810);
xnor U21234 (N_21234,N_20845,N_20871);
nor U21235 (N_21235,N_20840,N_20853);
nor U21236 (N_21236,N_20757,N_20813);
and U21237 (N_21237,N_20808,N_20774);
or U21238 (N_21238,N_20770,N_20945);
and U21239 (N_21239,N_20992,N_20987);
nor U21240 (N_21240,N_20959,N_20840);
or U21241 (N_21241,N_20912,N_20816);
nand U21242 (N_21242,N_20846,N_20898);
or U21243 (N_21243,N_20801,N_20825);
nor U21244 (N_21244,N_20847,N_20996);
or U21245 (N_21245,N_20863,N_20982);
xor U21246 (N_21246,N_20756,N_20938);
nand U21247 (N_21247,N_20876,N_20942);
and U21248 (N_21248,N_20753,N_20989);
nor U21249 (N_21249,N_20987,N_20820);
nor U21250 (N_21250,N_21115,N_21069);
and U21251 (N_21251,N_21232,N_21180);
xnor U21252 (N_21252,N_21167,N_21042);
xor U21253 (N_21253,N_21229,N_21124);
and U21254 (N_21254,N_21247,N_21012);
nor U21255 (N_21255,N_21198,N_21159);
and U21256 (N_21256,N_21108,N_21082);
nor U21257 (N_21257,N_21106,N_21191);
or U21258 (N_21258,N_21164,N_21013);
xnor U21259 (N_21259,N_21096,N_21181);
xnor U21260 (N_21260,N_21016,N_21213);
or U21261 (N_21261,N_21178,N_21199);
nand U21262 (N_21262,N_21222,N_21128);
xnor U21263 (N_21263,N_21221,N_21084);
and U21264 (N_21264,N_21102,N_21205);
or U21265 (N_21265,N_21033,N_21158);
nor U21266 (N_21266,N_21119,N_21067);
xor U21267 (N_21267,N_21104,N_21000);
or U21268 (N_21268,N_21236,N_21014);
nand U21269 (N_21269,N_21246,N_21116);
or U21270 (N_21270,N_21061,N_21209);
xnor U21271 (N_21271,N_21126,N_21017);
nor U21272 (N_21272,N_21211,N_21056);
nor U21273 (N_21273,N_21154,N_21215);
nor U21274 (N_21274,N_21023,N_21078);
nor U21275 (N_21275,N_21018,N_21197);
nand U21276 (N_21276,N_21006,N_21185);
or U21277 (N_21277,N_21114,N_21010);
nor U21278 (N_21278,N_21117,N_21110);
nor U21279 (N_21279,N_21129,N_21040);
xnor U21280 (N_21280,N_21008,N_21171);
xor U21281 (N_21281,N_21193,N_21174);
or U21282 (N_21282,N_21065,N_21169);
and U21283 (N_21283,N_21044,N_21123);
nand U21284 (N_21284,N_21026,N_21064);
xor U21285 (N_21285,N_21046,N_21068);
xor U21286 (N_21286,N_21004,N_21245);
nand U21287 (N_21287,N_21240,N_21217);
nand U21288 (N_21288,N_21085,N_21184);
xor U21289 (N_21289,N_21091,N_21179);
xor U21290 (N_21290,N_21107,N_21045);
nor U21291 (N_21291,N_21070,N_21095);
or U21292 (N_21292,N_21021,N_21168);
and U21293 (N_21293,N_21192,N_21005);
or U21294 (N_21294,N_21182,N_21242);
nand U21295 (N_21295,N_21233,N_21138);
and U21296 (N_21296,N_21075,N_21218);
and U21297 (N_21297,N_21146,N_21077);
nand U21298 (N_21298,N_21022,N_21132);
nor U21299 (N_21299,N_21208,N_21157);
xor U21300 (N_21300,N_21212,N_21002);
or U21301 (N_21301,N_21032,N_21139);
xor U21302 (N_21302,N_21210,N_21223);
nor U21303 (N_21303,N_21059,N_21173);
or U21304 (N_21304,N_21113,N_21142);
nand U21305 (N_21305,N_21225,N_21235);
nor U21306 (N_21306,N_21172,N_21152);
nor U21307 (N_21307,N_21066,N_21060);
nor U21308 (N_21308,N_21140,N_21196);
nor U21309 (N_21309,N_21072,N_21080);
nor U21310 (N_21310,N_21137,N_21216);
xor U21311 (N_21311,N_21219,N_21133);
nor U21312 (N_21312,N_21189,N_21086);
xor U21313 (N_21313,N_21001,N_21083);
xor U21314 (N_21314,N_21220,N_21099);
xor U21315 (N_21315,N_21048,N_21019);
and U21316 (N_21316,N_21074,N_21248);
nor U21317 (N_21317,N_21063,N_21009);
xor U21318 (N_21318,N_21226,N_21024);
nor U21319 (N_21319,N_21043,N_21030);
nor U21320 (N_21320,N_21122,N_21062);
xor U21321 (N_21321,N_21161,N_21094);
nand U21322 (N_21322,N_21151,N_21194);
or U21323 (N_21323,N_21155,N_21076);
or U21324 (N_21324,N_21111,N_21163);
nor U21325 (N_21325,N_21041,N_21090);
xnor U21326 (N_21326,N_21103,N_21055);
and U21327 (N_21327,N_21131,N_21097);
xor U21328 (N_21328,N_21204,N_21202);
nand U21329 (N_21329,N_21249,N_21071);
xnor U21330 (N_21330,N_21047,N_21098);
and U21331 (N_21331,N_21144,N_21244);
xnor U21332 (N_21332,N_21195,N_21058);
nor U21333 (N_21333,N_21214,N_21127);
nand U21334 (N_21334,N_21141,N_21175);
nor U21335 (N_21335,N_21201,N_21148);
and U21336 (N_21336,N_21037,N_21206);
nor U21337 (N_21337,N_21230,N_21120);
nor U21338 (N_21338,N_21176,N_21130);
and U21339 (N_21339,N_21136,N_21190);
nand U21340 (N_21340,N_21200,N_21011);
or U21341 (N_21341,N_21027,N_21092);
nand U21342 (N_21342,N_21147,N_21007);
nor U21343 (N_21343,N_21081,N_21112);
nand U21344 (N_21344,N_21227,N_21101);
or U21345 (N_21345,N_21088,N_21057);
nor U21346 (N_21346,N_21020,N_21228);
or U21347 (N_21347,N_21203,N_21207);
or U21348 (N_21348,N_21187,N_21105);
nor U21349 (N_21349,N_21170,N_21109);
xnor U21350 (N_21350,N_21162,N_21052);
xor U21351 (N_21351,N_21243,N_21025);
or U21352 (N_21352,N_21186,N_21239);
xnor U21353 (N_21353,N_21237,N_21031);
nor U21354 (N_21354,N_21053,N_21153);
xnor U21355 (N_21355,N_21079,N_21143);
or U21356 (N_21356,N_21087,N_21035);
and U21357 (N_21357,N_21038,N_21036);
xnor U21358 (N_21358,N_21093,N_21234);
nand U21359 (N_21359,N_21050,N_21145);
nor U21360 (N_21360,N_21166,N_21125);
and U21361 (N_21361,N_21049,N_21029);
and U21362 (N_21362,N_21183,N_21134);
nor U21363 (N_21363,N_21224,N_21165);
nand U21364 (N_21364,N_21015,N_21156);
nand U21365 (N_21365,N_21089,N_21238);
or U21366 (N_21366,N_21003,N_21177);
nor U21367 (N_21367,N_21073,N_21051);
xnor U21368 (N_21368,N_21150,N_21241);
xnor U21369 (N_21369,N_21039,N_21121);
and U21370 (N_21370,N_21034,N_21149);
xnor U21371 (N_21371,N_21028,N_21188);
nand U21372 (N_21372,N_21118,N_21160);
nand U21373 (N_21373,N_21231,N_21100);
and U21374 (N_21374,N_21135,N_21054);
nor U21375 (N_21375,N_21087,N_21186);
and U21376 (N_21376,N_21213,N_21044);
xor U21377 (N_21377,N_21062,N_21235);
or U21378 (N_21378,N_21053,N_21114);
or U21379 (N_21379,N_21009,N_21168);
xnor U21380 (N_21380,N_21247,N_21130);
nor U21381 (N_21381,N_21244,N_21070);
nand U21382 (N_21382,N_21038,N_21050);
xnor U21383 (N_21383,N_21030,N_21067);
or U21384 (N_21384,N_21120,N_21163);
nand U21385 (N_21385,N_21144,N_21029);
nand U21386 (N_21386,N_21248,N_21200);
nor U21387 (N_21387,N_21009,N_21184);
nor U21388 (N_21388,N_21104,N_21232);
nor U21389 (N_21389,N_21064,N_21137);
nor U21390 (N_21390,N_21177,N_21137);
or U21391 (N_21391,N_21171,N_21045);
and U21392 (N_21392,N_21152,N_21053);
and U21393 (N_21393,N_21149,N_21150);
or U21394 (N_21394,N_21114,N_21201);
nor U21395 (N_21395,N_21200,N_21015);
nand U21396 (N_21396,N_21004,N_21076);
and U21397 (N_21397,N_21234,N_21110);
xor U21398 (N_21398,N_21067,N_21083);
or U21399 (N_21399,N_21004,N_21141);
nand U21400 (N_21400,N_21096,N_21082);
nor U21401 (N_21401,N_21063,N_21056);
nand U21402 (N_21402,N_21243,N_21188);
or U21403 (N_21403,N_21189,N_21061);
nand U21404 (N_21404,N_21048,N_21172);
nor U21405 (N_21405,N_21208,N_21005);
xor U21406 (N_21406,N_21042,N_21083);
and U21407 (N_21407,N_21157,N_21172);
nor U21408 (N_21408,N_21143,N_21090);
nand U21409 (N_21409,N_21045,N_21063);
or U21410 (N_21410,N_21246,N_21022);
or U21411 (N_21411,N_21075,N_21150);
nand U21412 (N_21412,N_21238,N_21217);
and U21413 (N_21413,N_21047,N_21240);
or U21414 (N_21414,N_21214,N_21162);
and U21415 (N_21415,N_21080,N_21151);
nor U21416 (N_21416,N_21004,N_21090);
nor U21417 (N_21417,N_21207,N_21110);
nand U21418 (N_21418,N_21018,N_21174);
xnor U21419 (N_21419,N_21244,N_21054);
nand U21420 (N_21420,N_21136,N_21064);
nand U21421 (N_21421,N_21202,N_21096);
nor U21422 (N_21422,N_21156,N_21036);
and U21423 (N_21423,N_21062,N_21195);
nor U21424 (N_21424,N_21195,N_21139);
nor U21425 (N_21425,N_21217,N_21220);
nand U21426 (N_21426,N_21082,N_21195);
nor U21427 (N_21427,N_21164,N_21101);
xnor U21428 (N_21428,N_21037,N_21119);
or U21429 (N_21429,N_21111,N_21182);
or U21430 (N_21430,N_21112,N_21153);
xnor U21431 (N_21431,N_21035,N_21180);
and U21432 (N_21432,N_21210,N_21229);
or U21433 (N_21433,N_21061,N_21043);
xnor U21434 (N_21434,N_21081,N_21218);
xnor U21435 (N_21435,N_21126,N_21239);
nand U21436 (N_21436,N_21035,N_21032);
or U21437 (N_21437,N_21029,N_21058);
and U21438 (N_21438,N_21081,N_21132);
nor U21439 (N_21439,N_21232,N_21010);
and U21440 (N_21440,N_21107,N_21147);
and U21441 (N_21441,N_21057,N_21228);
nor U21442 (N_21442,N_21184,N_21174);
or U21443 (N_21443,N_21136,N_21199);
nor U21444 (N_21444,N_21229,N_21115);
and U21445 (N_21445,N_21236,N_21063);
and U21446 (N_21446,N_21093,N_21217);
and U21447 (N_21447,N_21041,N_21082);
nand U21448 (N_21448,N_21092,N_21167);
or U21449 (N_21449,N_21140,N_21097);
nor U21450 (N_21450,N_21118,N_21051);
xor U21451 (N_21451,N_21182,N_21239);
or U21452 (N_21452,N_21129,N_21143);
or U21453 (N_21453,N_21013,N_21017);
nor U21454 (N_21454,N_21108,N_21019);
and U21455 (N_21455,N_21199,N_21225);
xor U21456 (N_21456,N_21058,N_21197);
and U21457 (N_21457,N_21053,N_21049);
nor U21458 (N_21458,N_21007,N_21195);
or U21459 (N_21459,N_21136,N_21001);
or U21460 (N_21460,N_21222,N_21219);
nor U21461 (N_21461,N_21128,N_21030);
or U21462 (N_21462,N_21060,N_21051);
or U21463 (N_21463,N_21182,N_21035);
nor U21464 (N_21464,N_21162,N_21147);
nand U21465 (N_21465,N_21013,N_21178);
and U21466 (N_21466,N_21200,N_21231);
nor U21467 (N_21467,N_21163,N_21203);
xor U21468 (N_21468,N_21078,N_21199);
nor U21469 (N_21469,N_21185,N_21203);
xnor U21470 (N_21470,N_21021,N_21051);
xor U21471 (N_21471,N_21101,N_21091);
and U21472 (N_21472,N_21247,N_21115);
and U21473 (N_21473,N_21210,N_21116);
or U21474 (N_21474,N_21076,N_21018);
or U21475 (N_21475,N_21149,N_21002);
nand U21476 (N_21476,N_21185,N_21202);
nor U21477 (N_21477,N_21137,N_21168);
or U21478 (N_21478,N_21133,N_21131);
and U21479 (N_21479,N_21117,N_21179);
and U21480 (N_21480,N_21206,N_21012);
nand U21481 (N_21481,N_21065,N_21180);
nand U21482 (N_21482,N_21189,N_21172);
nand U21483 (N_21483,N_21042,N_21206);
xnor U21484 (N_21484,N_21206,N_21181);
or U21485 (N_21485,N_21058,N_21132);
xnor U21486 (N_21486,N_21115,N_21235);
or U21487 (N_21487,N_21173,N_21217);
or U21488 (N_21488,N_21170,N_21034);
nor U21489 (N_21489,N_21018,N_21219);
or U21490 (N_21490,N_21182,N_21227);
and U21491 (N_21491,N_21108,N_21141);
and U21492 (N_21492,N_21140,N_21005);
xnor U21493 (N_21493,N_21025,N_21176);
nand U21494 (N_21494,N_21191,N_21078);
xor U21495 (N_21495,N_21243,N_21240);
or U21496 (N_21496,N_21216,N_21015);
nand U21497 (N_21497,N_21151,N_21179);
xor U21498 (N_21498,N_21179,N_21185);
nor U21499 (N_21499,N_21228,N_21075);
and U21500 (N_21500,N_21415,N_21322);
or U21501 (N_21501,N_21428,N_21370);
xnor U21502 (N_21502,N_21290,N_21444);
xnor U21503 (N_21503,N_21297,N_21286);
nand U21504 (N_21504,N_21406,N_21295);
xor U21505 (N_21505,N_21300,N_21414);
and U21506 (N_21506,N_21425,N_21293);
xnor U21507 (N_21507,N_21356,N_21326);
and U21508 (N_21508,N_21296,N_21294);
nor U21509 (N_21509,N_21391,N_21487);
nor U21510 (N_21510,N_21320,N_21256);
nor U21511 (N_21511,N_21364,N_21366);
xor U21512 (N_21512,N_21258,N_21386);
nand U21513 (N_21513,N_21291,N_21439);
or U21514 (N_21514,N_21448,N_21408);
xnor U21515 (N_21515,N_21251,N_21335);
xnor U21516 (N_21516,N_21298,N_21309);
or U21517 (N_21517,N_21261,N_21469);
xnor U21518 (N_21518,N_21314,N_21306);
and U21519 (N_21519,N_21289,N_21421);
xnor U21520 (N_21520,N_21404,N_21476);
or U21521 (N_21521,N_21253,N_21467);
nand U21522 (N_21522,N_21280,N_21429);
xnor U21523 (N_21523,N_21316,N_21343);
nand U21524 (N_21524,N_21260,N_21311);
nor U21525 (N_21525,N_21460,N_21478);
or U21526 (N_21526,N_21492,N_21303);
nor U21527 (N_21527,N_21266,N_21488);
nand U21528 (N_21528,N_21250,N_21495);
nor U21529 (N_21529,N_21401,N_21349);
xor U21530 (N_21530,N_21327,N_21259);
nand U21531 (N_21531,N_21485,N_21416);
nor U21532 (N_21532,N_21325,N_21497);
or U21533 (N_21533,N_21486,N_21365);
or U21534 (N_21534,N_21292,N_21449);
or U21535 (N_21535,N_21400,N_21452);
xor U21536 (N_21536,N_21436,N_21465);
nor U21537 (N_21537,N_21323,N_21264);
nand U21538 (N_21538,N_21281,N_21466);
xor U21539 (N_21539,N_21282,N_21474);
or U21540 (N_21540,N_21257,N_21288);
nand U21541 (N_21541,N_21403,N_21389);
or U21542 (N_21542,N_21437,N_21441);
and U21543 (N_21543,N_21407,N_21350);
nor U21544 (N_21544,N_21273,N_21346);
and U21545 (N_21545,N_21344,N_21479);
nand U21546 (N_21546,N_21284,N_21371);
nor U21547 (N_21547,N_21456,N_21412);
nand U21548 (N_21548,N_21464,N_21475);
nand U21549 (N_21549,N_21384,N_21328);
nand U21550 (N_21550,N_21397,N_21454);
nor U21551 (N_21551,N_21431,N_21376);
or U21552 (N_21552,N_21418,N_21269);
nand U21553 (N_21553,N_21402,N_21305);
xnor U21554 (N_21554,N_21361,N_21447);
and U21555 (N_21555,N_21473,N_21489);
nor U21556 (N_21556,N_21347,N_21274);
nand U21557 (N_21557,N_21304,N_21494);
and U21558 (N_21558,N_21276,N_21337);
xnor U21559 (N_21559,N_21424,N_21443);
and U21560 (N_21560,N_21332,N_21321);
nand U21561 (N_21561,N_21267,N_21278);
and U21562 (N_21562,N_21360,N_21413);
xor U21563 (N_21563,N_21468,N_21279);
nor U21564 (N_21564,N_21362,N_21382);
nor U21565 (N_21565,N_21383,N_21462);
nand U21566 (N_21566,N_21399,N_21324);
nand U21567 (N_21567,N_21345,N_21351);
nor U21568 (N_21568,N_21378,N_21355);
xor U21569 (N_21569,N_21419,N_21338);
xnor U21570 (N_21570,N_21353,N_21398);
and U21571 (N_21571,N_21265,N_21254);
or U21572 (N_21572,N_21333,N_21255);
and U21573 (N_21573,N_21363,N_21285);
nand U21574 (N_21574,N_21268,N_21329);
nor U21575 (N_21575,N_21302,N_21334);
and U21576 (N_21576,N_21381,N_21379);
and U21577 (N_21577,N_21368,N_21310);
xnor U21578 (N_21578,N_21433,N_21481);
nand U21579 (N_21579,N_21272,N_21480);
nor U21580 (N_21580,N_21318,N_21390);
nor U21581 (N_21581,N_21423,N_21499);
or U21582 (N_21582,N_21319,N_21312);
xnor U21583 (N_21583,N_21336,N_21417);
nor U21584 (N_21584,N_21341,N_21377);
or U21585 (N_21585,N_21409,N_21463);
nor U21586 (N_21586,N_21430,N_21446);
or U21587 (N_21587,N_21471,N_21358);
or U21588 (N_21588,N_21308,N_21369);
and U21589 (N_21589,N_21373,N_21270);
xor U21590 (N_21590,N_21275,N_21422);
or U21591 (N_21591,N_21375,N_21385);
or U21592 (N_21592,N_21396,N_21459);
xnor U21593 (N_21593,N_21339,N_21442);
nand U21594 (N_21594,N_21331,N_21445);
nor U21595 (N_21595,N_21359,N_21393);
nor U21596 (N_21596,N_21432,N_21461);
xor U21597 (N_21597,N_21287,N_21427);
and U21598 (N_21598,N_21411,N_21271);
or U21599 (N_21599,N_21301,N_21317);
or U21600 (N_21600,N_21405,N_21262);
nor U21601 (N_21601,N_21354,N_21434);
xor U21602 (N_21602,N_21496,N_21420);
nor U21603 (N_21603,N_21348,N_21490);
or U21604 (N_21604,N_21313,N_21392);
nand U21605 (N_21605,N_21435,N_21483);
xor U21606 (N_21606,N_21482,N_21455);
and U21607 (N_21607,N_21263,N_21440);
and U21608 (N_21608,N_21395,N_21457);
xnor U21609 (N_21609,N_21484,N_21477);
nand U21610 (N_21610,N_21498,N_21394);
nor U21611 (N_21611,N_21352,N_21451);
nand U21612 (N_21612,N_21340,N_21277);
or U21613 (N_21613,N_21367,N_21374);
xnor U21614 (N_21614,N_21387,N_21438);
or U21615 (N_21615,N_21342,N_21315);
nor U21616 (N_21616,N_21380,N_21493);
or U21617 (N_21617,N_21307,N_21357);
xnor U21618 (N_21618,N_21299,N_21388);
or U21619 (N_21619,N_21283,N_21330);
xor U21620 (N_21620,N_21426,N_21472);
xor U21621 (N_21621,N_21450,N_21470);
nand U21622 (N_21622,N_21252,N_21410);
xor U21623 (N_21623,N_21372,N_21458);
xor U21624 (N_21624,N_21453,N_21491);
xor U21625 (N_21625,N_21288,N_21364);
and U21626 (N_21626,N_21287,N_21331);
or U21627 (N_21627,N_21335,N_21301);
nor U21628 (N_21628,N_21264,N_21465);
nor U21629 (N_21629,N_21431,N_21330);
xnor U21630 (N_21630,N_21411,N_21448);
or U21631 (N_21631,N_21477,N_21385);
or U21632 (N_21632,N_21453,N_21479);
nor U21633 (N_21633,N_21470,N_21420);
nand U21634 (N_21634,N_21440,N_21364);
nand U21635 (N_21635,N_21353,N_21420);
nor U21636 (N_21636,N_21266,N_21472);
or U21637 (N_21637,N_21305,N_21284);
nand U21638 (N_21638,N_21472,N_21263);
and U21639 (N_21639,N_21399,N_21451);
and U21640 (N_21640,N_21296,N_21297);
or U21641 (N_21641,N_21286,N_21406);
and U21642 (N_21642,N_21265,N_21474);
xnor U21643 (N_21643,N_21476,N_21276);
nor U21644 (N_21644,N_21452,N_21385);
nand U21645 (N_21645,N_21354,N_21301);
xor U21646 (N_21646,N_21451,N_21306);
nand U21647 (N_21647,N_21353,N_21496);
or U21648 (N_21648,N_21277,N_21474);
nand U21649 (N_21649,N_21336,N_21272);
and U21650 (N_21650,N_21495,N_21360);
nand U21651 (N_21651,N_21318,N_21459);
and U21652 (N_21652,N_21333,N_21475);
nor U21653 (N_21653,N_21399,N_21257);
xnor U21654 (N_21654,N_21299,N_21263);
nand U21655 (N_21655,N_21467,N_21297);
nor U21656 (N_21656,N_21258,N_21266);
nor U21657 (N_21657,N_21309,N_21397);
and U21658 (N_21658,N_21460,N_21398);
or U21659 (N_21659,N_21469,N_21429);
or U21660 (N_21660,N_21398,N_21299);
nor U21661 (N_21661,N_21403,N_21287);
nor U21662 (N_21662,N_21337,N_21485);
nand U21663 (N_21663,N_21402,N_21281);
nor U21664 (N_21664,N_21372,N_21477);
or U21665 (N_21665,N_21432,N_21405);
and U21666 (N_21666,N_21330,N_21340);
nor U21667 (N_21667,N_21425,N_21427);
nor U21668 (N_21668,N_21261,N_21271);
nand U21669 (N_21669,N_21264,N_21306);
and U21670 (N_21670,N_21449,N_21430);
nor U21671 (N_21671,N_21454,N_21411);
and U21672 (N_21672,N_21338,N_21253);
nand U21673 (N_21673,N_21374,N_21368);
nand U21674 (N_21674,N_21279,N_21451);
nor U21675 (N_21675,N_21451,N_21417);
nand U21676 (N_21676,N_21488,N_21275);
or U21677 (N_21677,N_21456,N_21489);
nor U21678 (N_21678,N_21330,N_21400);
xor U21679 (N_21679,N_21388,N_21438);
nand U21680 (N_21680,N_21478,N_21345);
nor U21681 (N_21681,N_21333,N_21373);
nand U21682 (N_21682,N_21310,N_21442);
and U21683 (N_21683,N_21419,N_21411);
nor U21684 (N_21684,N_21414,N_21259);
or U21685 (N_21685,N_21406,N_21489);
and U21686 (N_21686,N_21288,N_21441);
nand U21687 (N_21687,N_21321,N_21293);
or U21688 (N_21688,N_21368,N_21358);
xnor U21689 (N_21689,N_21296,N_21257);
xnor U21690 (N_21690,N_21407,N_21275);
nand U21691 (N_21691,N_21427,N_21417);
and U21692 (N_21692,N_21402,N_21352);
xnor U21693 (N_21693,N_21373,N_21430);
nor U21694 (N_21694,N_21391,N_21332);
nor U21695 (N_21695,N_21403,N_21392);
nor U21696 (N_21696,N_21448,N_21414);
and U21697 (N_21697,N_21407,N_21309);
xor U21698 (N_21698,N_21351,N_21322);
and U21699 (N_21699,N_21378,N_21371);
nor U21700 (N_21700,N_21488,N_21310);
nand U21701 (N_21701,N_21360,N_21496);
or U21702 (N_21702,N_21495,N_21309);
xor U21703 (N_21703,N_21493,N_21323);
nor U21704 (N_21704,N_21302,N_21296);
xor U21705 (N_21705,N_21355,N_21361);
nor U21706 (N_21706,N_21264,N_21296);
xor U21707 (N_21707,N_21321,N_21394);
nor U21708 (N_21708,N_21369,N_21374);
and U21709 (N_21709,N_21419,N_21481);
and U21710 (N_21710,N_21482,N_21488);
nand U21711 (N_21711,N_21279,N_21473);
nand U21712 (N_21712,N_21488,N_21446);
xor U21713 (N_21713,N_21301,N_21363);
or U21714 (N_21714,N_21366,N_21375);
xnor U21715 (N_21715,N_21436,N_21329);
and U21716 (N_21716,N_21358,N_21290);
nand U21717 (N_21717,N_21335,N_21452);
nor U21718 (N_21718,N_21299,N_21498);
or U21719 (N_21719,N_21345,N_21385);
and U21720 (N_21720,N_21340,N_21486);
or U21721 (N_21721,N_21274,N_21296);
xor U21722 (N_21722,N_21361,N_21386);
or U21723 (N_21723,N_21262,N_21322);
or U21724 (N_21724,N_21259,N_21290);
or U21725 (N_21725,N_21353,N_21477);
or U21726 (N_21726,N_21268,N_21416);
xnor U21727 (N_21727,N_21494,N_21451);
or U21728 (N_21728,N_21325,N_21367);
or U21729 (N_21729,N_21309,N_21437);
nand U21730 (N_21730,N_21452,N_21451);
xnor U21731 (N_21731,N_21498,N_21472);
and U21732 (N_21732,N_21382,N_21376);
xnor U21733 (N_21733,N_21382,N_21495);
and U21734 (N_21734,N_21341,N_21257);
xnor U21735 (N_21735,N_21434,N_21419);
nand U21736 (N_21736,N_21313,N_21291);
nor U21737 (N_21737,N_21454,N_21314);
xor U21738 (N_21738,N_21480,N_21286);
and U21739 (N_21739,N_21448,N_21481);
or U21740 (N_21740,N_21351,N_21468);
xnor U21741 (N_21741,N_21413,N_21257);
and U21742 (N_21742,N_21431,N_21329);
or U21743 (N_21743,N_21327,N_21415);
xnor U21744 (N_21744,N_21434,N_21493);
or U21745 (N_21745,N_21359,N_21368);
and U21746 (N_21746,N_21296,N_21459);
nand U21747 (N_21747,N_21352,N_21416);
and U21748 (N_21748,N_21485,N_21404);
or U21749 (N_21749,N_21417,N_21278);
nor U21750 (N_21750,N_21535,N_21732);
nand U21751 (N_21751,N_21630,N_21571);
nor U21752 (N_21752,N_21632,N_21730);
nor U21753 (N_21753,N_21739,N_21504);
or U21754 (N_21754,N_21537,N_21547);
nor U21755 (N_21755,N_21714,N_21720);
and U21756 (N_21756,N_21601,N_21650);
nand U21757 (N_21757,N_21579,N_21511);
xnor U21758 (N_21758,N_21531,N_21690);
or U21759 (N_21759,N_21523,N_21611);
and U21760 (N_21760,N_21738,N_21530);
and U21761 (N_21761,N_21731,N_21681);
or U21762 (N_21762,N_21736,N_21508);
nor U21763 (N_21763,N_21599,N_21705);
and U21764 (N_21764,N_21696,N_21604);
xor U21765 (N_21765,N_21574,N_21592);
and U21766 (N_21766,N_21608,N_21694);
xor U21767 (N_21767,N_21578,N_21674);
and U21768 (N_21768,N_21622,N_21595);
nor U21769 (N_21769,N_21713,N_21518);
nand U21770 (N_21770,N_21575,N_21631);
nor U21771 (N_21771,N_21613,N_21671);
nand U21772 (N_21772,N_21610,N_21512);
nor U21773 (N_21773,N_21554,N_21698);
or U21774 (N_21774,N_21552,N_21729);
nand U21775 (N_21775,N_21623,N_21708);
xnor U21776 (N_21776,N_21600,N_21514);
xnor U21777 (N_21777,N_21524,N_21581);
and U21778 (N_21778,N_21706,N_21548);
and U21779 (N_21779,N_21702,N_21679);
nor U21780 (N_21780,N_21648,N_21593);
nor U21781 (N_21781,N_21687,N_21555);
xor U21782 (N_21782,N_21634,N_21689);
and U21783 (N_21783,N_21625,N_21586);
nand U21784 (N_21784,N_21543,N_21549);
or U21785 (N_21785,N_21527,N_21519);
xor U21786 (N_21786,N_21576,N_21737);
and U21787 (N_21787,N_21685,N_21725);
xor U21788 (N_21788,N_21636,N_21562);
or U21789 (N_21789,N_21747,N_21664);
xor U21790 (N_21790,N_21672,N_21724);
xor U21791 (N_21791,N_21528,N_21609);
nor U21792 (N_21792,N_21680,N_21645);
nor U21793 (N_21793,N_21564,N_21605);
and U21794 (N_21794,N_21651,N_21734);
nand U21795 (N_21795,N_21626,N_21550);
nor U21796 (N_21796,N_21726,N_21569);
nor U21797 (N_21797,N_21585,N_21742);
and U21798 (N_21798,N_21667,N_21642);
or U21799 (N_21799,N_21587,N_21612);
and U21800 (N_21800,N_21712,N_21596);
nand U21801 (N_21801,N_21715,N_21746);
nor U21802 (N_21802,N_21627,N_21529);
or U21803 (N_21803,N_21691,N_21614);
and U21804 (N_21804,N_21591,N_21561);
xor U21805 (N_21805,N_21516,N_21682);
and U21806 (N_21806,N_21520,N_21704);
or U21807 (N_21807,N_21649,N_21656);
xnor U21808 (N_21808,N_21540,N_21666);
or U21809 (N_21809,N_21657,N_21639);
and U21810 (N_21810,N_21616,N_21733);
and U21811 (N_21811,N_21545,N_21635);
nor U21812 (N_21812,N_21647,N_21534);
nor U21813 (N_21813,N_21583,N_21669);
and U21814 (N_21814,N_21655,N_21602);
xor U21815 (N_21815,N_21644,N_21629);
nand U21816 (N_21816,N_21638,N_21517);
and U21817 (N_21817,N_21515,N_21748);
and U21818 (N_21818,N_21503,N_21653);
nor U21819 (N_21819,N_21589,N_21701);
xor U21820 (N_21820,N_21743,N_21624);
and U21821 (N_21821,N_21709,N_21567);
or U21822 (N_21822,N_21711,N_21525);
or U21823 (N_21823,N_21594,N_21686);
nor U21824 (N_21824,N_21532,N_21526);
nand U21825 (N_21825,N_21665,N_21584);
and U21826 (N_21826,N_21717,N_21615);
and U21827 (N_21827,N_21501,N_21675);
or U21828 (N_21828,N_21621,N_21536);
and U21829 (N_21829,N_21546,N_21658);
or U21830 (N_21830,N_21640,N_21670);
or U21831 (N_21831,N_21618,N_21727);
nand U21832 (N_21832,N_21607,N_21707);
xnor U21833 (N_21833,N_21728,N_21565);
nor U21834 (N_21834,N_21570,N_21556);
nor U21835 (N_21835,N_21541,N_21577);
xnor U21836 (N_21836,N_21646,N_21533);
and U21837 (N_21837,N_21695,N_21673);
or U21838 (N_21838,N_21509,N_21603);
xor U21839 (N_21839,N_21722,N_21542);
nor U21840 (N_21840,N_21572,N_21740);
or U21841 (N_21841,N_21597,N_21505);
nor U21842 (N_21842,N_21684,N_21551);
xor U21843 (N_21843,N_21566,N_21582);
or U21844 (N_21844,N_21678,N_21700);
nand U21845 (N_21845,N_21558,N_21633);
or U21846 (N_21846,N_21617,N_21676);
nand U21847 (N_21847,N_21710,N_21502);
nor U21848 (N_21848,N_21513,N_21654);
nor U21849 (N_21849,N_21507,N_21539);
xor U21850 (N_21850,N_21568,N_21544);
nand U21851 (N_21851,N_21573,N_21683);
and U21852 (N_21852,N_21628,N_21588);
or U21853 (N_21853,N_21652,N_21723);
nand U21854 (N_21854,N_21619,N_21521);
xor U21855 (N_21855,N_21688,N_21620);
or U21856 (N_21856,N_21661,N_21741);
xnor U21857 (N_21857,N_21745,N_21557);
xnor U21858 (N_21858,N_21721,N_21643);
nor U21859 (N_21859,N_21563,N_21510);
nor U21860 (N_21860,N_21692,N_21560);
or U21861 (N_21861,N_21703,N_21559);
xor U21862 (N_21862,N_21719,N_21598);
xnor U21863 (N_21863,N_21744,N_21606);
or U21864 (N_21864,N_21663,N_21641);
xor U21865 (N_21865,N_21668,N_21662);
or U21866 (N_21866,N_21553,N_21590);
and U21867 (N_21867,N_21699,N_21500);
and U21868 (N_21868,N_21735,N_21522);
xor U21869 (N_21869,N_21693,N_21697);
nand U21870 (N_21870,N_21718,N_21538);
and U21871 (N_21871,N_21716,N_21506);
xnor U21872 (N_21872,N_21637,N_21677);
xor U21873 (N_21873,N_21749,N_21659);
nand U21874 (N_21874,N_21660,N_21580);
xnor U21875 (N_21875,N_21556,N_21730);
xnor U21876 (N_21876,N_21685,N_21635);
nand U21877 (N_21877,N_21684,N_21672);
xnor U21878 (N_21878,N_21560,N_21671);
xnor U21879 (N_21879,N_21570,N_21661);
nor U21880 (N_21880,N_21700,N_21606);
nand U21881 (N_21881,N_21709,N_21613);
nor U21882 (N_21882,N_21595,N_21528);
nor U21883 (N_21883,N_21625,N_21744);
and U21884 (N_21884,N_21723,N_21662);
nand U21885 (N_21885,N_21719,N_21642);
nor U21886 (N_21886,N_21550,N_21592);
nand U21887 (N_21887,N_21632,N_21577);
and U21888 (N_21888,N_21660,N_21717);
nand U21889 (N_21889,N_21568,N_21615);
nand U21890 (N_21890,N_21529,N_21511);
nand U21891 (N_21891,N_21577,N_21652);
xnor U21892 (N_21892,N_21700,N_21556);
xor U21893 (N_21893,N_21550,N_21567);
nor U21894 (N_21894,N_21697,N_21728);
or U21895 (N_21895,N_21630,N_21609);
xnor U21896 (N_21896,N_21630,N_21728);
and U21897 (N_21897,N_21508,N_21547);
and U21898 (N_21898,N_21703,N_21528);
and U21899 (N_21899,N_21604,N_21625);
or U21900 (N_21900,N_21518,N_21548);
nor U21901 (N_21901,N_21569,N_21672);
nor U21902 (N_21902,N_21732,N_21580);
and U21903 (N_21903,N_21740,N_21696);
nor U21904 (N_21904,N_21599,N_21583);
and U21905 (N_21905,N_21681,N_21636);
nor U21906 (N_21906,N_21687,N_21695);
nor U21907 (N_21907,N_21619,N_21724);
or U21908 (N_21908,N_21599,N_21624);
and U21909 (N_21909,N_21735,N_21550);
and U21910 (N_21910,N_21501,N_21731);
or U21911 (N_21911,N_21525,N_21657);
nand U21912 (N_21912,N_21583,N_21550);
and U21913 (N_21913,N_21546,N_21702);
nand U21914 (N_21914,N_21740,N_21631);
nor U21915 (N_21915,N_21524,N_21722);
nand U21916 (N_21916,N_21593,N_21687);
or U21917 (N_21917,N_21718,N_21590);
nand U21918 (N_21918,N_21638,N_21506);
nand U21919 (N_21919,N_21614,N_21653);
nor U21920 (N_21920,N_21610,N_21528);
and U21921 (N_21921,N_21594,N_21607);
nor U21922 (N_21922,N_21592,N_21672);
and U21923 (N_21923,N_21664,N_21508);
or U21924 (N_21924,N_21548,N_21744);
and U21925 (N_21925,N_21720,N_21678);
nand U21926 (N_21926,N_21640,N_21505);
nor U21927 (N_21927,N_21529,N_21681);
or U21928 (N_21928,N_21615,N_21585);
nor U21929 (N_21929,N_21622,N_21639);
nor U21930 (N_21930,N_21614,N_21607);
xnor U21931 (N_21931,N_21736,N_21690);
nand U21932 (N_21932,N_21546,N_21535);
xor U21933 (N_21933,N_21572,N_21563);
or U21934 (N_21934,N_21612,N_21577);
and U21935 (N_21935,N_21519,N_21713);
nor U21936 (N_21936,N_21707,N_21549);
nand U21937 (N_21937,N_21668,N_21661);
and U21938 (N_21938,N_21688,N_21578);
xor U21939 (N_21939,N_21562,N_21708);
xor U21940 (N_21940,N_21535,N_21536);
nor U21941 (N_21941,N_21598,N_21710);
xor U21942 (N_21942,N_21685,N_21640);
and U21943 (N_21943,N_21728,N_21693);
or U21944 (N_21944,N_21549,N_21604);
nand U21945 (N_21945,N_21508,N_21641);
or U21946 (N_21946,N_21699,N_21737);
nor U21947 (N_21947,N_21561,N_21502);
nand U21948 (N_21948,N_21569,N_21628);
nand U21949 (N_21949,N_21523,N_21683);
and U21950 (N_21950,N_21724,N_21622);
nand U21951 (N_21951,N_21642,N_21595);
and U21952 (N_21952,N_21714,N_21520);
or U21953 (N_21953,N_21599,N_21683);
nor U21954 (N_21954,N_21615,N_21511);
nor U21955 (N_21955,N_21634,N_21726);
nor U21956 (N_21956,N_21608,N_21641);
and U21957 (N_21957,N_21651,N_21723);
or U21958 (N_21958,N_21689,N_21527);
and U21959 (N_21959,N_21599,N_21743);
or U21960 (N_21960,N_21560,N_21660);
and U21961 (N_21961,N_21559,N_21502);
nor U21962 (N_21962,N_21634,N_21711);
xnor U21963 (N_21963,N_21688,N_21643);
and U21964 (N_21964,N_21500,N_21537);
nand U21965 (N_21965,N_21504,N_21572);
xor U21966 (N_21966,N_21604,N_21727);
or U21967 (N_21967,N_21539,N_21635);
xnor U21968 (N_21968,N_21509,N_21534);
xor U21969 (N_21969,N_21557,N_21615);
and U21970 (N_21970,N_21594,N_21640);
xor U21971 (N_21971,N_21506,N_21658);
nor U21972 (N_21972,N_21705,N_21597);
nor U21973 (N_21973,N_21534,N_21741);
nand U21974 (N_21974,N_21650,N_21532);
nor U21975 (N_21975,N_21613,N_21749);
xnor U21976 (N_21976,N_21642,N_21729);
nor U21977 (N_21977,N_21613,N_21645);
nand U21978 (N_21978,N_21725,N_21613);
or U21979 (N_21979,N_21540,N_21674);
xor U21980 (N_21980,N_21681,N_21536);
nor U21981 (N_21981,N_21501,N_21728);
or U21982 (N_21982,N_21514,N_21586);
or U21983 (N_21983,N_21663,N_21661);
or U21984 (N_21984,N_21718,N_21555);
and U21985 (N_21985,N_21527,N_21740);
xnor U21986 (N_21986,N_21530,N_21734);
xor U21987 (N_21987,N_21705,N_21515);
xor U21988 (N_21988,N_21707,N_21630);
nor U21989 (N_21989,N_21549,N_21724);
nand U21990 (N_21990,N_21508,N_21506);
nand U21991 (N_21991,N_21707,N_21579);
or U21992 (N_21992,N_21718,N_21716);
xnor U21993 (N_21993,N_21668,N_21575);
nand U21994 (N_21994,N_21679,N_21552);
nor U21995 (N_21995,N_21662,N_21738);
and U21996 (N_21996,N_21519,N_21600);
nor U21997 (N_21997,N_21712,N_21548);
nor U21998 (N_21998,N_21641,N_21549);
or U21999 (N_21999,N_21723,N_21562);
or U22000 (N_22000,N_21849,N_21843);
nor U22001 (N_22001,N_21980,N_21928);
and U22002 (N_22002,N_21850,N_21835);
and U22003 (N_22003,N_21870,N_21768);
nor U22004 (N_22004,N_21770,N_21769);
xor U22005 (N_22005,N_21898,N_21905);
and U22006 (N_22006,N_21948,N_21955);
xor U22007 (N_22007,N_21902,N_21956);
nor U22008 (N_22008,N_21848,N_21958);
xnor U22009 (N_22009,N_21767,N_21982);
nand U22010 (N_22010,N_21942,N_21775);
nor U22011 (N_22011,N_21764,N_21917);
nor U22012 (N_22012,N_21914,N_21951);
or U22013 (N_22013,N_21933,N_21924);
nor U22014 (N_22014,N_21784,N_21971);
and U22015 (N_22015,N_21871,N_21832);
xnor U22016 (N_22016,N_21973,N_21891);
and U22017 (N_22017,N_21961,N_21998);
nor U22018 (N_22018,N_21817,N_21861);
xnor U22019 (N_22019,N_21975,N_21864);
or U22020 (N_22020,N_21856,N_21904);
nor U22021 (N_22021,N_21972,N_21801);
xnor U22022 (N_22022,N_21766,N_21815);
nand U22023 (N_22023,N_21751,N_21908);
and U22024 (N_22024,N_21841,N_21992);
nor U22025 (N_22025,N_21798,N_21964);
nand U22026 (N_22026,N_21960,N_21869);
and U22027 (N_22027,N_21842,N_21903);
xnor U22028 (N_22028,N_21929,N_21776);
nand U22029 (N_22029,N_21878,N_21874);
nor U22030 (N_22030,N_21959,N_21943);
or U22031 (N_22031,N_21774,N_21920);
nor U22032 (N_22032,N_21834,N_21862);
nor U22033 (N_22033,N_21965,N_21937);
nand U22034 (N_22034,N_21762,N_21783);
and U22035 (N_22035,N_21896,N_21887);
or U22036 (N_22036,N_21811,N_21854);
nor U22037 (N_22037,N_21875,N_21820);
xnor U22038 (N_22038,N_21977,N_21799);
nand U22039 (N_22039,N_21840,N_21866);
or U22040 (N_22040,N_21909,N_21976);
and U22041 (N_22041,N_21863,N_21824);
nor U22042 (N_22042,N_21804,N_21922);
and U22043 (N_22043,N_21828,N_21771);
nand U22044 (N_22044,N_21830,N_21938);
and U22045 (N_22045,N_21996,N_21994);
xnor U22046 (N_22046,N_21808,N_21759);
nor U22047 (N_22047,N_21823,N_21906);
nand U22048 (N_22048,N_21995,N_21974);
xnor U22049 (N_22049,N_21950,N_21760);
xor U22050 (N_22050,N_21756,N_21868);
or U22051 (N_22051,N_21907,N_21797);
nor U22052 (N_22052,N_21763,N_21886);
xnor U22053 (N_22053,N_21931,N_21754);
xnor U22054 (N_22054,N_21919,N_21791);
nor U22055 (N_22055,N_21880,N_21802);
and U22056 (N_22056,N_21913,N_21939);
or U22057 (N_22057,N_21993,N_21836);
xor U22058 (N_22058,N_21847,N_21803);
nand U22059 (N_22059,N_21821,N_21912);
nor U22060 (N_22060,N_21758,N_21786);
xor U22061 (N_22061,N_21789,N_21860);
nand U22062 (N_22062,N_21921,N_21881);
xor U22063 (N_22063,N_21999,N_21852);
or U22064 (N_22064,N_21831,N_21845);
nor U22065 (N_22065,N_21925,N_21957);
xor U22066 (N_22066,N_21872,N_21916);
nand U22067 (N_22067,N_21989,N_21892);
or U22068 (N_22068,N_21941,N_21927);
nand U22069 (N_22069,N_21794,N_21779);
or U22070 (N_22070,N_21773,N_21788);
nor U22071 (N_22071,N_21936,N_21990);
xor U22072 (N_22072,N_21889,N_21792);
and U22073 (N_22073,N_21837,N_21893);
or U22074 (N_22074,N_21978,N_21926);
nand U22075 (N_22075,N_21827,N_21963);
nand U22076 (N_22076,N_21838,N_21986);
xnor U22077 (N_22077,N_21895,N_21790);
and U22078 (N_22078,N_21859,N_21879);
and U22079 (N_22079,N_21988,N_21777);
nand U22080 (N_22080,N_21882,N_21780);
xor U22081 (N_22081,N_21750,N_21983);
nor U22082 (N_22082,N_21953,N_21833);
nand U22083 (N_22083,N_21997,N_21873);
nor U22084 (N_22084,N_21765,N_21944);
and U22085 (N_22085,N_21839,N_21884);
or U22086 (N_22086,N_21962,N_21844);
nor U22087 (N_22087,N_21985,N_21781);
nor U22088 (N_22088,N_21979,N_21785);
nand U22089 (N_22089,N_21947,N_21778);
nor U22090 (N_22090,N_21813,N_21918);
nor U22091 (N_22091,N_21911,N_21816);
and U22092 (N_22092,N_21945,N_21814);
nand U22093 (N_22093,N_21888,N_21805);
or U22094 (N_22094,N_21899,N_21855);
nand U22095 (N_22095,N_21800,N_21987);
nand U22096 (N_22096,N_21755,N_21853);
or U22097 (N_22097,N_21901,N_21793);
xnor U22098 (N_22098,N_21900,N_21772);
nor U22099 (N_22099,N_21984,N_21930);
and U22100 (N_22100,N_21807,N_21946);
and U22101 (N_22101,N_21825,N_21952);
and U22102 (N_22102,N_21818,N_21822);
nand U22103 (N_22103,N_21969,N_21806);
nand U22104 (N_22104,N_21940,N_21981);
nor U22105 (N_22105,N_21753,N_21812);
nor U22106 (N_22106,N_21883,N_21846);
nand U22107 (N_22107,N_21782,N_21809);
nor U22108 (N_22108,N_21858,N_21970);
nor U22109 (N_22109,N_21910,N_21954);
or U22110 (N_22110,N_21894,N_21796);
or U22111 (N_22111,N_21867,N_21851);
xor U22112 (N_22112,N_21819,N_21915);
xnor U22113 (N_22113,N_21934,N_21857);
nor U22114 (N_22114,N_21932,N_21897);
and U22115 (N_22115,N_21877,N_21991);
and U22116 (N_22116,N_21968,N_21829);
or U22117 (N_22117,N_21787,N_21865);
xnor U22118 (N_22118,N_21949,N_21752);
nand U22119 (N_22119,N_21795,N_21935);
xnor U22120 (N_22120,N_21757,N_21966);
and U22121 (N_22121,N_21885,N_21826);
xnor U22122 (N_22122,N_21876,N_21810);
nand U22123 (N_22123,N_21761,N_21890);
or U22124 (N_22124,N_21923,N_21967);
or U22125 (N_22125,N_21869,N_21910);
nand U22126 (N_22126,N_21789,N_21934);
or U22127 (N_22127,N_21972,N_21850);
or U22128 (N_22128,N_21780,N_21856);
nor U22129 (N_22129,N_21862,N_21864);
or U22130 (N_22130,N_21965,N_21963);
or U22131 (N_22131,N_21876,N_21941);
xor U22132 (N_22132,N_21892,N_21921);
nor U22133 (N_22133,N_21915,N_21978);
nand U22134 (N_22134,N_21854,N_21765);
and U22135 (N_22135,N_21771,N_21820);
and U22136 (N_22136,N_21882,N_21894);
nor U22137 (N_22137,N_21807,N_21870);
nor U22138 (N_22138,N_21987,N_21966);
and U22139 (N_22139,N_21800,N_21836);
nor U22140 (N_22140,N_21811,N_21909);
nand U22141 (N_22141,N_21805,N_21784);
xnor U22142 (N_22142,N_21884,N_21865);
nor U22143 (N_22143,N_21832,N_21968);
nor U22144 (N_22144,N_21969,N_21867);
and U22145 (N_22145,N_21979,N_21924);
or U22146 (N_22146,N_21860,N_21977);
xor U22147 (N_22147,N_21858,N_21992);
or U22148 (N_22148,N_21797,N_21796);
or U22149 (N_22149,N_21938,N_21914);
and U22150 (N_22150,N_21862,N_21923);
xor U22151 (N_22151,N_21839,N_21831);
or U22152 (N_22152,N_21977,N_21888);
nand U22153 (N_22153,N_21945,N_21953);
or U22154 (N_22154,N_21842,N_21868);
nor U22155 (N_22155,N_21909,N_21793);
nor U22156 (N_22156,N_21763,N_21915);
xnor U22157 (N_22157,N_21959,N_21808);
xnor U22158 (N_22158,N_21801,N_21837);
xnor U22159 (N_22159,N_21891,N_21982);
and U22160 (N_22160,N_21868,N_21979);
or U22161 (N_22161,N_21842,N_21787);
or U22162 (N_22162,N_21910,N_21966);
nand U22163 (N_22163,N_21769,N_21894);
nand U22164 (N_22164,N_21942,N_21863);
nand U22165 (N_22165,N_21820,N_21836);
xor U22166 (N_22166,N_21971,N_21930);
xnor U22167 (N_22167,N_21925,N_21902);
nor U22168 (N_22168,N_21761,N_21897);
and U22169 (N_22169,N_21960,N_21882);
or U22170 (N_22170,N_21957,N_21857);
or U22171 (N_22171,N_21781,N_21874);
nand U22172 (N_22172,N_21857,N_21893);
or U22173 (N_22173,N_21780,N_21936);
xor U22174 (N_22174,N_21776,N_21821);
and U22175 (N_22175,N_21809,N_21975);
or U22176 (N_22176,N_21892,N_21931);
or U22177 (N_22177,N_21780,N_21992);
nor U22178 (N_22178,N_21855,N_21920);
nand U22179 (N_22179,N_21766,N_21780);
xor U22180 (N_22180,N_21983,N_21752);
xnor U22181 (N_22181,N_21831,N_21862);
or U22182 (N_22182,N_21940,N_21952);
xor U22183 (N_22183,N_21932,N_21818);
xor U22184 (N_22184,N_21780,N_21993);
xor U22185 (N_22185,N_21789,N_21863);
or U22186 (N_22186,N_21757,N_21994);
nand U22187 (N_22187,N_21947,N_21979);
nor U22188 (N_22188,N_21854,N_21780);
xnor U22189 (N_22189,N_21907,N_21795);
or U22190 (N_22190,N_21757,N_21989);
xnor U22191 (N_22191,N_21810,N_21768);
or U22192 (N_22192,N_21880,N_21788);
and U22193 (N_22193,N_21758,N_21883);
and U22194 (N_22194,N_21878,N_21959);
or U22195 (N_22195,N_21959,N_21978);
xnor U22196 (N_22196,N_21924,N_21819);
and U22197 (N_22197,N_21923,N_21954);
or U22198 (N_22198,N_21751,N_21868);
nor U22199 (N_22199,N_21781,N_21872);
xor U22200 (N_22200,N_21766,N_21799);
or U22201 (N_22201,N_21911,N_21937);
nand U22202 (N_22202,N_21893,N_21854);
or U22203 (N_22203,N_21957,N_21985);
nand U22204 (N_22204,N_21817,N_21820);
or U22205 (N_22205,N_21832,N_21945);
nor U22206 (N_22206,N_21760,N_21757);
xor U22207 (N_22207,N_21967,N_21796);
nand U22208 (N_22208,N_21799,N_21843);
xor U22209 (N_22209,N_21882,N_21766);
nand U22210 (N_22210,N_21922,N_21835);
nor U22211 (N_22211,N_21777,N_21975);
and U22212 (N_22212,N_21832,N_21884);
nand U22213 (N_22213,N_21966,N_21821);
nand U22214 (N_22214,N_21889,N_21865);
nand U22215 (N_22215,N_21768,N_21804);
xor U22216 (N_22216,N_21833,N_21849);
xnor U22217 (N_22217,N_21831,N_21843);
and U22218 (N_22218,N_21794,N_21826);
xor U22219 (N_22219,N_21785,N_21866);
or U22220 (N_22220,N_21772,N_21855);
nand U22221 (N_22221,N_21854,N_21806);
nor U22222 (N_22222,N_21997,N_21891);
xnor U22223 (N_22223,N_21822,N_21921);
nor U22224 (N_22224,N_21757,N_21776);
nand U22225 (N_22225,N_21769,N_21983);
and U22226 (N_22226,N_21887,N_21866);
or U22227 (N_22227,N_21826,N_21874);
xnor U22228 (N_22228,N_21775,N_21797);
and U22229 (N_22229,N_21774,N_21805);
xnor U22230 (N_22230,N_21995,N_21970);
nor U22231 (N_22231,N_21890,N_21854);
xor U22232 (N_22232,N_21950,N_21922);
or U22233 (N_22233,N_21878,N_21960);
and U22234 (N_22234,N_21915,N_21838);
nor U22235 (N_22235,N_21782,N_21784);
or U22236 (N_22236,N_21965,N_21856);
xor U22237 (N_22237,N_21924,N_21787);
nor U22238 (N_22238,N_21802,N_21983);
and U22239 (N_22239,N_21812,N_21981);
nand U22240 (N_22240,N_21892,N_21888);
nor U22241 (N_22241,N_21976,N_21754);
xor U22242 (N_22242,N_21860,N_21778);
and U22243 (N_22243,N_21863,N_21975);
and U22244 (N_22244,N_21891,N_21810);
xnor U22245 (N_22245,N_21979,N_21970);
nand U22246 (N_22246,N_21859,N_21887);
and U22247 (N_22247,N_21961,N_21902);
nand U22248 (N_22248,N_21802,N_21782);
xnor U22249 (N_22249,N_21969,N_21997);
nor U22250 (N_22250,N_22093,N_22208);
xor U22251 (N_22251,N_22149,N_22230);
or U22252 (N_22252,N_22231,N_22009);
or U22253 (N_22253,N_22058,N_22153);
nor U22254 (N_22254,N_22095,N_22119);
nand U22255 (N_22255,N_22057,N_22083);
nand U22256 (N_22256,N_22244,N_22146);
xnor U22257 (N_22257,N_22175,N_22090);
xor U22258 (N_22258,N_22236,N_22131);
and U22259 (N_22259,N_22063,N_22108);
xnor U22260 (N_22260,N_22213,N_22042);
nand U22261 (N_22261,N_22139,N_22245);
xnor U22262 (N_22262,N_22077,N_22008);
nor U22263 (N_22263,N_22140,N_22219);
nor U22264 (N_22264,N_22167,N_22045);
xor U22265 (N_22265,N_22118,N_22004);
nor U22266 (N_22266,N_22059,N_22136);
xor U22267 (N_22267,N_22056,N_22080);
xor U22268 (N_22268,N_22029,N_22151);
and U22269 (N_22269,N_22106,N_22122);
and U22270 (N_22270,N_22165,N_22053);
xnor U22271 (N_22271,N_22159,N_22068);
xor U22272 (N_22272,N_22210,N_22064);
nor U22273 (N_22273,N_22094,N_22086);
nand U22274 (N_22274,N_22242,N_22051);
nand U22275 (N_22275,N_22249,N_22246);
nand U22276 (N_22276,N_22007,N_22003);
nand U22277 (N_22277,N_22224,N_22241);
nand U22278 (N_22278,N_22105,N_22162);
or U22279 (N_22279,N_22134,N_22120);
nand U22280 (N_22280,N_22174,N_22043);
nand U22281 (N_22281,N_22019,N_22147);
or U22282 (N_22282,N_22070,N_22182);
and U22283 (N_22283,N_22141,N_22099);
and U22284 (N_22284,N_22016,N_22079);
xor U22285 (N_22285,N_22185,N_22110);
and U22286 (N_22286,N_22187,N_22235);
xor U22287 (N_22287,N_22065,N_22215);
or U22288 (N_22288,N_22037,N_22217);
nand U22289 (N_22289,N_22171,N_22025);
xor U22290 (N_22290,N_22178,N_22076);
nor U22291 (N_22291,N_22115,N_22001);
nor U22292 (N_22292,N_22000,N_22047);
xnor U22293 (N_22293,N_22107,N_22010);
or U22294 (N_22294,N_22156,N_22223);
and U22295 (N_22295,N_22145,N_22128);
nor U22296 (N_22296,N_22232,N_22170);
or U22297 (N_22297,N_22101,N_22052);
or U22298 (N_22298,N_22160,N_22143);
and U22299 (N_22299,N_22084,N_22015);
xnor U22300 (N_22300,N_22221,N_22155);
and U22301 (N_22301,N_22172,N_22133);
and U22302 (N_22302,N_22186,N_22197);
xor U22303 (N_22303,N_22032,N_22247);
nand U22304 (N_22304,N_22227,N_22188);
and U22305 (N_22305,N_22204,N_22117);
nand U22306 (N_22306,N_22096,N_22066);
or U22307 (N_22307,N_22098,N_22201);
nand U22308 (N_22308,N_22193,N_22179);
nor U22309 (N_22309,N_22206,N_22132);
and U22310 (N_22310,N_22028,N_22041);
and U22311 (N_22311,N_22126,N_22138);
nor U22312 (N_22312,N_22006,N_22233);
xnor U22313 (N_22313,N_22192,N_22209);
nand U22314 (N_22314,N_22112,N_22190);
nor U22315 (N_22315,N_22240,N_22154);
or U22316 (N_22316,N_22248,N_22100);
nor U22317 (N_22317,N_22049,N_22048);
and U22318 (N_22318,N_22237,N_22044);
xor U22319 (N_22319,N_22092,N_22013);
or U22320 (N_22320,N_22033,N_22129);
and U22321 (N_22321,N_22088,N_22239);
or U22322 (N_22322,N_22082,N_22198);
nand U22323 (N_22323,N_22169,N_22017);
and U22324 (N_22324,N_22113,N_22027);
and U22325 (N_22325,N_22243,N_22014);
or U22326 (N_22326,N_22046,N_22137);
and U22327 (N_22327,N_22002,N_22199);
and U22328 (N_22328,N_22050,N_22104);
nor U22329 (N_22329,N_22157,N_22228);
or U22330 (N_22330,N_22163,N_22135);
nand U22331 (N_22331,N_22189,N_22089);
xor U22332 (N_22332,N_22124,N_22055);
xor U22333 (N_22333,N_22150,N_22024);
nor U22334 (N_22334,N_22021,N_22023);
nand U22335 (N_22335,N_22097,N_22087);
nor U22336 (N_22336,N_22234,N_22012);
and U22337 (N_22337,N_22102,N_22207);
nand U22338 (N_22338,N_22121,N_22222);
nor U22339 (N_22339,N_22060,N_22074);
xnor U22340 (N_22340,N_22069,N_22130);
nand U22341 (N_22341,N_22072,N_22177);
nor U22342 (N_22342,N_22005,N_22091);
or U22343 (N_22343,N_22184,N_22195);
or U22344 (N_22344,N_22144,N_22200);
xnor U22345 (N_22345,N_22218,N_22173);
xor U22346 (N_22346,N_22109,N_22194);
or U22347 (N_22347,N_22035,N_22011);
or U22348 (N_22348,N_22111,N_22022);
nor U22349 (N_22349,N_22078,N_22226);
and U22350 (N_22350,N_22085,N_22229);
xor U22351 (N_22351,N_22203,N_22081);
nor U22352 (N_22352,N_22036,N_22020);
xnor U22353 (N_22353,N_22211,N_22181);
nor U22354 (N_22354,N_22191,N_22214);
nand U22355 (N_22355,N_22148,N_22038);
or U22356 (N_22356,N_22054,N_22062);
nor U22357 (N_22357,N_22040,N_22212);
nor U22358 (N_22358,N_22216,N_22125);
or U22359 (N_22359,N_22061,N_22176);
nor U22360 (N_22360,N_22158,N_22073);
nor U22361 (N_22361,N_22123,N_22026);
and U22362 (N_22362,N_22202,N_22018);
nand U22363 (N_22363,N_22168,N_22205);
and U22364 (N_22364,N_22103,N_22034);
and U22365 (N_22365,N_22127,N_22116);
nor U22366 (N_22366,N_22161,N_22142);
nor U22367 (N_22367,N_22238,N_22152);
or U22368 (N_22368,N_22030,N_22180);
nor U22369 (N_22369,N_22071,N_22067);
nor U22370 (N_22370,N_22031,N_22183);
and U22371 (N_22371,N_22075,N_22166);
xnor U22372 (N_22372,N_22039,N_22114);
nand U22373 (N_22373,N_22164,N_22220);
nand U22374 (N_22374,N_22225,N_22196);
and U22375 (N_22375,N_22171,N_22054);
nand U22376 (N_22376,N_22114,N_22220);
nand U22377 (N_22377,N_22098,N_22135);
or U22378 (N_22378,N_22183,N_22208);
xnor U22379 (N_22379,N_22095,N_22219);
nand U22380 (N_22380,N_22054,N_22231);
and U22381 (N_22381,N_22066,N_22230);
and U22382 (N_22382,N_22239,N_22182);
xnor U22383 (N_22383,N_22101,N_22049);
nor U22384 (N_22384,N_22022,N_22208);
or U22385 (N_22385,N_22044,N_22191);
or U22386 (N_22386,N_22185,N_22062);
and U22387 (N_22387,N_22176,N_22113);
nor U22388 (N_22388,N_22165,N_22054);
or U22389 (N_22389,N_22039,N_22011);
nand U22390 (N_22390,N_22179,N_22049);
nor U22391 (N_22391,N_22191,N_22150);
and U22392 (N_22392,N_22094,N_22003);
and U22393 (N_22393,N_22159,N_22222);
xor U22394 (N_22394,N_22021,N_22064);
nor U22395 (N_22395,N_22228,N_22007);
xor U22396 (N_22396,N_22196,N_22064);
and U22397 (N_22397,N_22079,N_22226);
nor U22398 (N_22398,N_22049,N_22056);
and U22399 (N_22399,N_22138,N_22186);
and U22400 (N_22400,N_22095,N_22024);
and U22401 (N_22401,N_22038,N_22017);
and U22402 (N_22402,N_22114,N_22068);
nor U22403 (N_22403,N_22029,N_22124);
and U22404 (N_22404,N_22248,N_22152);
and U22405 (N_22405,N_22220,N_22072);
or U22406 (N_22406,N_22118,N_22199);
nand U22407 (N_22407,N_22118,N_22053);
nor U22408 (N_22408,N_22238,N_22000);
and U22409 (N_22409,N_22141,N_22222);
xor U22410 (N_22410,N_22025,N_22013);
or U22411 (N_22411,N_22084,N_22012);
nand U22412 (N_22412,N_22216,N_22219);
nand U22413 (N_22413,N_22113,N_22223);
nand U22414 (N_22414,N_22002,N_22140);
xor U22415 (N_22415,N_22162,N_22076);
nor U22416 (N_22416,N_22098,N_22028);
or U22417 (N_22417,N_22238,N_22147);
xnor U22418 (N_22418,N_22186,N_22241);
nand U22419 (N_22419,N_22071,N_22008);
nand U22420 (N_22420,N_22036,N_22115);
nand U22421 (N_22421,N_22244,N_22059);
nor U22422 (N_22422,N_22161,N_22224);
nor U22423 (N_22423,N_22119,N_22089);
nor U22424 (N_22424,N_22148,N_22004);
nor U22425 (N_22425,N_22044,N_22062);
and U22426 (N_22426,N_22084,N_22104);
or U22427 (N_22427,N_22080,N_22040);
nor U22428 (N_22428,N_22123,N_22122);
xnor U22429 (N_22429,N_22188,N_22083);
nor U22430 (N_22430,N_22212,N_22123);
nor U22431 (N_22431,N_22239,N_22222);
and U22432 (N_22432,N_22140,N_22154);
and U22433 (N_22433,N_22002,N_22019);
and U22434 (N_22434,N_22200,N_22236);
nand U22435 (N_22435,N_22074,N_22186);
nand U22436 (N_22436,N_22122,N_22018);
nand U22437 (N_22437,N_22104,N_22032);
or U22438 (N_22438,N_22180,N_22064);
xnor U22439 (N_22439,N_22249,N_22204);
or U22440 (N_22440,N_22090,N_22118);
or U22441 (N_22441,N_22104,N_22109);
or U22442 (N_22442,N_22083,N_22143);
nor U22443 (N_22443,N_22055,N_22074);
nand U22444 (N_22444,N_22078,N_22082);
and U22445 (N_22445,N_22090,N_22088);
nand U22446 (N_22446,N_22214,N_22185);
xor U22447 (N_22447,N_22178,N_22097);
and U22448 (N_22448,N_22041,N_22119);
nand U22449 (N_22449,N_22077,N_22132);
and U22450 (N_22450,N_22160,N_22246);
nor U22451 (N_22451,N_22031,N_22215);
or U22452 (N_22452,N_22137,N_22014);
and U22453 (N_22453,N_22087,N_22012);
xor U22454 (N_22454,N_22240,N_22167);
or U22455 (N_22455,N_22088,N_22065);
and U22456 (N_22456,N_22165,N_22068);
nor U22457 (N_22457,N_22018,N_22060);
or U22458 (N_22458,N_22074,N_22128);
and U22459 (N_22459,N_22136,N_22151);
xnor U22460 (N_22460,N_22005,N_22081);
xor U22461 (N_22461,N_22014,N_22246);
nand U22462 (N_22462,N_22003,N_22169);
or U22463 (N_22463,N_22030,N_22161);
nand U22464 (N_22464,N_22015,N_22039);
nor U22465 (N_22465,N_22081,N_22029);
nor U22466 (N_22466,N_22164,N_22012);
nand U22467 (N_22467,N_22107,N_22126);
xor U22468 (N_22468,N_22134,N_22043);
or U22469 (N_22469,N_22066,N_22154);
or U22470 (N_22470,N_22206,N_22104);
nor U22471 (N_22471,N_22128,N_22087);
nand U22472 (N_22472,N_22101,N_22018);
and U22473 (N_22473,N_22239,N_22047);
xor U22474 (N_22474,N_22119,N_22130);
and U22475 (N_22475,N_22027,N_22174);
xor U22476 (N_22476,N_22171,N_22148);
nor U22477 (N_22477,N_22008,N_22015);
or U22478 (N_22478,N_22071,N_22159);
nor U22479 (N_22479,N_22024,N_22048);
nor U22480 (N_22480,N_22186,N_22058);
or U22481 (N_22481,N_22004,N_22194);
and U22482 (N_22482,N_22114,N_22010);
nand U22483 (N_22483,N_22212,N_22052);
or U22484 (N_22484,N_22022,N_22116);
or U22485 (N_22485,N_22025,N_22180);
nor U22486 (N_22486,N_22244,N_22071);
or U22487 (N_22487,N_22151,N_22105);
or U22488 (N_22488,N_22167,N_22080);
nand U22489 (N_22489,N_22030,N_22009);
and U22490 (N_22490,N_22190,N_22015);
nand U22491 (N_22491,N_22226,N_22006);
and U22492 (N_22492,N_22056,N_22109);
nor U22493 (N_22493,N_22248,N_22144);
nand U22494 (N_22494,N_22064,N_22162);
xor U22495 (N_22495,N_22152,N_22222);
and U22496 (N_22496,N_22008,N_22172);
and U22497 (N_22497,N_22117,N_22170);
nand U22498 (N_22498,N_22029,N_22209);
nand U22499 (N_22499,N_22198,N_22118);
nand U22500 (N_22500,N_22279,N_22435);
and U22501 (N_22501,N_22423,N_22466);
xnor U22502 (N_22502,N_22454,N_22339);
and U22503 (N_22503,N_22491,N_22283);
and U22504 (N_22504,N_22480,N_22386);
and U22505 (N_22505,N_22366,N_22291);
nor U22506 (N_22506,N_22318,N_22364);
and U22507 (N_22507,N_22262,N_22481);
or U22508 (N_22508,N_22275,N_22414);
and U22509 (N_22509,N_22444,N_22297);
or U22510 (N_22510,N_22400,N_22383);
nor U22511 (N_22511,N_22371,N_22267);
and U22512 (N_22512,N_22358,N_22314);
xnor U22513 (N_22513,N_22349,N_22378);
nand U22514 (N_22514,N_22406,N_22440);
nand U22515 (N_22515,N_22261,N_22348);
and U22516 (N_22516,N_22461,N_22344);
xnor U22517 (N_22517,N_22300,N_22257);
or U22518 (N_22518,N_22477,N_22379);
xor U22519 (N_22519,N_22418,N_22280);
nor U22520 (N_22520,N_22496,N_22368);
nor U22521 (N_22521,N_22375,N_22304);
or U22522 (N_22522,N_22473,N_22486);
nand U22523 (N_22523,N_22327,N_22252);
and U22524 (N_22524,N_22497,N_22484);
nor U22525 (N_22525,N_22258,N_22487);
nand U22526 (N_22526,N_22399,N_22431);
xor U22527 (N_22527,N_22436,N_22325);
xnor U22528 (N_22528,N_22299,N_22424);
or U22529 (N_22529,N_22485,N_22492);
or U22530 (N_22530,N_22351,N_22360);
or U22531 (N_22531,N_22405,N_22317);
nor U22532 (N_22532,N_22394,N_22359);
nand U22533 (N_22533,N_22441,N_22373);
and U22534 (N_22534,N_22316,N_22323);
xor U22535 (N_22535,N_22447,N_22362);
nand U22536 (N_22536,N_22456,N_22273);
xnor U22537 (N_22537,N_22263,N_22271);
nand U22538 (N_22538,N_22256,N_22421);
or U22539 (N_22539,N_22397,N_22255);
and U22540 (N_22540,N_22489,N_22471);
nand U22541 (N_22541,N_22369,N_22333);
xnor U22542 (N_22542,N_22446,N_22437);
nand U22543 (N_22543,N_22412,N_22286);
or U22544 (N_22544,N_22387,N_22250);
xnor U22545 (N_22545,N_22452,N_22465);
nand U22546 (N_22546,N_22409,N_22337);
and U22547 (N_22547,N_22415,N_22384);
and U22548 (N_22548,N_22393,N_22305);
or U22549 (N_22549,N_22347,N_22254);
nand U22550 (N_22550,N_22493,N_22476);
and U22551 (N_22551,N_22445,N_22478);
nor U22552 (N_22552,N_22322,N_22319);
nor U22553 (N_22553,N_22310,N_22342);
xor U22554 (N_22554,N_22468,N_22350);
nand U22555 (N_22555,N_22462,N_22425);
nand U22556 (N_22556,N_22479,N_22494);
xnor U22557 (N_22557,N_22268,N_22251);
xnor U22558 (N_22558,N_22433,N_22357);
nand U22559 (N_22559,N_22426,N_22451);
and U22560 (N_22560,N_22401,N_22303);
nand U22561 (N_22561,N_22392,N_22430);
nand U22562 (N_22562,N_22294,N_22259);
xnor U22563 (N_22563,N_22457,N_22274);
and U22564 (N_22564,N_22326,N_22289);
or U22565 (N_22565,N_22301,N_22346);
xor U22566 (N_22566,N_22296,N_22396);
or U22567 (N_22567,N_22408,N_22328);
or U22568 (N_22568,N_22352,N_22374);
and U22569 (N_22569,N_22427,N_22385);
and U22570 (N_22570,N_22302,N_22288);
xor U22571 (N_22571,N_22276,N_22464);
and U22572 (N_22572,N_22482,N_22432);
nand U22573 (N_22573,N_22388,N_22499);
nor U22574 (N_22574,N_22463,N_22356);
or U22575 (N_22575,N_22469,N_22449);
nor U22576 (N_22576,N_22495,N_22419);
and U22577 (N_22577,N_22284,N_22354);
or U22578 (N_22578,N_22306,N_22372);
nor U22579 (N_22579,N_22285,N_22411);
nor U22580 (N_22580,N_22260,N_22293);
xor U22581 (N_22581,N_22287,N_22353);
nand U22582 (N_22582,N_22309,N_22355);
nand U22583 (N_22583,N_22470,N_22343);
xnor U22584 (N_22584,N_22467,N_22340);
xnor U22585 (N_22585,N_22443,N_22330);
nor U22586 (N_22586,N_22341,N_22266);
nand U22587 (N_22587,N_22270,N_22404);
nor U22588 (N_22588,N_22455,N_22295);
and U22589 (N_22589,N_22265,N_22410);
xor U22590 (N_22590,N_22345,N_22367);
nor U22591 (N_22591,N_22311,N_22380);
and U22592 (N_22592,N_22417,N_22332);
nor U22593 (N_22593,N_22398,N_22269);
and U22594 (N_22594,N_22403,N_22395);
and U22595 (N_22595,N_22474,N_22498);
xor U22596 (N_22596,N_22490,N_22298);
and U22597 (N_22597,N_22434,N_22338);
nand U22598 (N_22598,N_22281,N_22329);
and U22599 (N_22599,N_22475,N_22450);
or U22600 (N_22600,N_22282,N_22413);
nor U22601 (N_22601,N_22389,N_22253);
nor U22602 (N_22602,N_22420,N_22365);
or U22603 (N_22603,N_22320,N_22290);
and U22604 (N_22604,N_22292,N_22382);
or U22605 (N_22605,N_22428,N_22390);
nand U22606 (N_22606,N_22381,N_22334);
nor U22607 (N_22607,N_22458,N_22278);
xor U22608 (N_22608,N_22448,N_22264);
nand U22609 (N_22609,N_22321,N_22453);
nand U22610 (N_22610,N_22488,N_22315);
xnor U22611 (N_22611,N_22336,N_22324);
nand U22612 (N_22612,N_22312,N_22308);
nor U22613 (N_22613,N_22370,N_22460);
nor U22614 (N_22614,N_22363,N_22459);
xnor U22615 (N_22615,N_22377,N_22313);
nand U22616 (N_22616,N_22472,N_22439);
and U22617 (N_22617,N_22429,N_22407);
and U22618 (N_22618,N_22331,N_22277);
and U22619 (N_22619,N_22416,N_22483);
nor U22620 (N_22620,N_22335,N_22376);
xor U22621 (N_22621,N_22442,N_22422);
nor U22622 (N_22622,N_22272,N_22391);
nand U22623 (N_22623,N_22307,N_22438);
nor U22624 (N_22624,N_22361,N_22402);
nand U22625 (N_22625,N_22338,N_22335);
nor U22626 (N_22626,N_22286,N_22462);
xor U22627 (N_22627,N_22277,N_22391);
and U22628 (N_22628,N_22463,N_22358);
nor U22629 (N_22629,N_22392,N_22473);
or U22630 (N_22630,N_22391,N_22336);
nor U22631 (N_22631,N_22314,N_22422);
xor U22632 (N_22632,N_22450,N_22380);
xor U22633 (N_22633,N_22473,N_22326);
or U22634 (N_22634,N_22386,N_22483);
nor U22635 (N_22635,N_22301,N_22435);
and U22636 (N_22636,N_22270,N_22331);
and U22637 (N_22637,N_22383,N_22360);
or U22638 (N_22638,N_22434,N_22370);
xor U22639 (N_22639,N_22472,N_22397);
xnor U22640 (N_22640,N_22252,N_22460);
nand U22641 (N_22641,N_22386,N_22347);
nand U22642 (N_22642,N_22427,N_22412);
or U22643 (N_22643,N_22334,N_22364);
xnor U22644 (N_22644,N_22461,N_22459);
or U22645 (N_22645,N_22499,N_22283);
or U22646 (N_22646,N_22473,N_22497);
nand U22647 (N_22647,N_22319,N_22472);
nand U22648 (N_22648,N_22257,N_22381);
xor U22649 (N_22649,N_22453,N_22390);
nand U22650 (N_22650,N_22492,N_22397);
or U22651 (N_22651,N_22307,N_22445);
xnor U22652 (N_22652,N_22256,N_22291);
or U22653 (N_22653,N_22326,N_22422);
xor U22654 (N_22654,N_22357,N_22293);
xnor U22655 (N_22655,N_22344,N_22372);
and U22656 (N_22656,N_22353,N_22484);
xnor U22657 (N_22657,N_22428,N_22263);
nor U22658 (N_22658,N_22271,N_22486);
or U22659 (N_22659,N_22350,N_22484);
and U22660 (N_22660,N_22381,N_22295);
nor U22661 (N_22661,N_22272,N_22458);
or U22662 (N_22662,N_22327,N_22456);
xnor U22663 (N_22663,N_22279,N_22496);
xor U22664 (N_22664,N_22436,N_22313);
and U22665 (N_22665,N_22460,N_22274);
nor U22666 (N_22666,N_22484,N_22406);
or U22667 (N_22667,N_22286,N_22330);
nand U22668 (N_22668,N_22369,N_22478);
nand U22669 (N_22669,N_22472,N_22308);
nand U22670 (N_22670,N_22298,N_22462);
nor U22671 (N_22671,N_22495,N_22452);
and U22672 (N_22672,N_22250,N_22283);
nand U22673 (N_22673,N_22348,N_22278);
nand U22674 (N_22674,N_22388,N_22468);
and U22675 (N_22675,N_22348,N_22254);
and U22676 (N_22676,N_22481,N_22415);
or U22677 (N_22677,N_22464,N_22284);
nor U22678 (N_22678,N_22289,N_22462);
nand U22679 (N_22679,N_22432,N_22429);
or U22680 (N_22680,N_22465,N_22495);
and U22681 (N_22681,N_22306,N_22250);
nor U22682 (N_22682,N_22408,N_22325);
xor U22683 (N_22683,N_22315,N_22446);
nor U22684 (N_22684,N_22280,N_22303);
nand U22685 (N_22685,N_22326,N_22370);
xor U22686 (N_22686,N_22426,N_22417);
xor U22687 (N_22687,N_22344,N_22280);
xnor U22688 (N_22688,N_22325,N_22267);
xnor U22689 (N_22689,N_22351,N_22487);
nor U22690 (N_22690,N_22261,N_22408);
xnor U22691 (N_22691,N_22405,N_22305);
nor U22692 (N_22692,N_22459,N_22361);
nand U22693 (N_22693,N_22384,N_22499);
nand U22694 (N_22694,N_22455,N_22266);
or U22695 (N_22695,N_22454,N_22260);
xnor U22696 (N_22696,N_22363,N_22267);
and U22697 (N_22697,N_22479,N_22456);
nor U22698 (N_22698,N_22266,N_22305);
nor U22699 (N_22699,N_22405,N_22319);
nand U22700 (N_22700,N_22329,N_22493);
or U22701 (N_22701,N_22265,N_22457);
nand U22702 (N_22702,N_22350,N_22401);
nor U22703 (N_22703,N_22313,N_22311);
or U22704 (N_22704,N_22352,N_22442);
xor U22705 (N_22705,N_22268,N_22253);
xor U22706 (N_22706,N_22314,N_22299);
and U22707 (N_22707,N_22431,N_22388);
xnor U22708 (N_22708,N_22405,N_22426);
or U22709 (N_22709,N_22463,N_22412);
or U22710 (N_22710,N_22478,N_22411);
or U22711 (N_22711,N_22313,N_22360);
nor U22712 (N_22712,N_22472,N_22341);
and U22713 (N_22713,N_22395,N_22447);
nor U22714 (N_22714,N_22417,N_22327);
xor U22715 (N_22715,N_22258,N_22417);
xor U22716 (N_22716,N_22381,N_22499);
and U22717 (N_22717,N_22449,N_22428);
or U22718 (N_22718,N_22412,N_22344);
nor U22719 (N_22719,N_22419,N_22287);
and U22720 (N_22720,N_22262,N_22400);
nor U22721 (N_22721,N_22274,N_22343);
xor U22722 (N_22722,N_22495,N_22318);
xor U22723 (N_22723,N_22289,N_22299);
xnor U22724 (N_22724,N_22274,N_22349);
xnor U22725 (N_22725,N_22411,N_22331);
xnor U22726 (N_22726,N_22278,N_22496);
nand U22727 (N_22727,N_22298,N_22444);
xnor U22728 (N_22728,N_22371,N_22370);
nor U22729 (N_22729,N_22426,N_22473);
or U22730 (N_22730,N_22341,N_22407);
or U22731 (N_22731,N_22446,N_22317);
nand U22732 (N_22732,N_22417,N_22303);
or U22733 (N_22733,N_22305,N_22486);
nand U22734 (N_22734,N_22310,N_22332);
nor U22735 (N_22735,N_22295,N_22414);
or U22736 (N_22736,N_22287,N_22468);
or U22737 (N_22737,N_22477,N_22499);
xnor U22738 (N_22738,N_22488,N_22497);
nor U22739 (N_22739,N_22280,N_22372);
nand U22740 (N_22740,N_22349,N_22425);
nand U22741 (N_22741,N_22371,N_22251);
xnor U22742 (N_22742,N_22282,N_22270);
nor U22743 (N_22743,N_22435,N_22313);
nor U22744 (N_22744,N_22355,N_22372);
xnor U22745 (N_22745,N_22449,N_22273);
nor U22746 (N_22746,N_22490,N_22346);
or U22747 (N_22747,N_22445,N_22258);
and U22748 (N_22748,N_22330,N_22255);
nor U22749 (N_22749,N_22288,N_22368);
nor U22750 (N_22750,N_22669,N_22592);
xnor U22751 (N_22751,N_22561,N_22746);
xnor U22752 (N_22752,N_22520,N_22586);
nand U22753 (N_22753,N_22580,N_22670);
xnor U22754 (N_22754,N_22594,N_22527);
nor U22755 (N_22755,N_22649,N_22579);
xnor U22756 (N_22756,N_22734,N_22727);
and U22757 (N_22757,N_22533,N_22713);
and U22758 (N_22758,N_22747,N_22552);
nor U22759 (N_22759,N_22578,N_22745);
nor U22760 (N_22760,N_22591,N_22684);
xor U22761 (N_22761,N_22554,N_22729);
nor U22762 (N_22762,N_22572,N_22528);
nand U22763 (N_22763,N_22665,N_22650);
or U22764 (N_22764,N_22557,N_22673);
nand U22765 (N_22765,N_22521,N_22716);
or U22766 (N_22766,N_22545,N_22524);
and U22767 (N_22767,N_22699,N_22706);
nand U22768 (N_22768,N_22530,N_22562);
or U22769 (N_22769,N_22659,N_22505);
nand U22770 (N_22770,N_22709,N_22531);
or U22771 (N_22771,N_22656,N_22648);
or U22772 (N_22772,N_22671,N_22574);
and U22773 (N_22773,N_22740,N_22596);
nor U22774 (N_22774,N_22525,N_22715);
nor U22775 (N_22775,N_22518,N_22685);
xnor U22776 (N_22776,N_22598,N_22725);
and U22777 (N_22777,N_22666,N_22507);
nor U22778 (N_22778,N_22697,N_22695);
nand U22779 (N_22779,N_22693,N_22582);
xnor U22780 (N_22780,N_22679,N_22575);
nand U22781 (N_22781,N_22587,N_22717);
nand U22782 (N_22782,N_22718,N_22732);
nor U22783 (N_22783,N_22658,N_22645);
or U22784 (N_22784,N_22742,N_22514);
xnor U22785 (N_22785,N_22712,N_22563);
nor U22786 (N_22786,N_22577,N_22733);
xnor U22787 (N_22787,N_22517,N_22631);
and U22788 (N_22788,N_22635,N_22647);
or U22789 (N_22789,N_22636,N_22642);
xnor U22790 (N_22790,N_22537,N_22630);
nor U22791 (N_22791,N_22682,N_22651);
nand U22792 (N_22792,N_22541,N_22519);
nand U22793 (N_22793,N_22700,N_22550);
and U22794 (N_22794,N_22613,N_22705);
nand U22795 (N_22795,N_22739,N_22628);
xnor U22796 (N_22796,N_22724,N_22597);
nor U22797 (N_22797,N_22609,N_22543);
and U22798 (N_22798,N_22619,N_22616);
nor U22799 (N_22799,N_22622,N_22620);
or U22800 (N_22800,N_22566,N_22694);
nor U22801 (N_22801,N_22637,N_22547);
xnor U22802 (N_22802,N_22504,N_22714);
or U22803 (N_22803,N_22526,N_22736);
nor U22804 (N_22804,N_22687,N_22680);
nor U22805 (N_22805,N_22568,N_22662);
or U22806 (N_22806,N_22653,N_22535);
xnor U22807 (N_22807,N_22604,N_22702);
and U22808 (N_22808,N_22617,N_22564);
and U22809 (N_22809,N_22721,N_22735);
xnor U22810 (N_22810,N_22556,N_22641);
or U22811 (N_22811,N_22611,N_22502);
nand U22812 (N_22812,N_22503,N_22544);
or U22813 (N_22813,N_22607,N_22626);
nor U22814 (N_22814,N_22612,N_22590);
and U22815 (N_22815,N_22744,N_22707);
and U22816 (N_22816,N_22560,N_22546);
nand U22817 (N_22817,N_22515,N_22614);
xnor U22818 (N_22818,N_22555,N_22640);
nor U22819 (N_22819,N_22608,N_22540);
xnor U22820 (N_22820,N_22688,N_22536);
or U22821 (N_22821,N_22660,N_22664);
nor U22822 (N_22822,N_22749,N_22573);
or U22823 (N_22823,N_22511,N_22708);
xor U22824 (N_22824,N_22567,N_22672);
or U22825 (N_22825,N_22539,N_22675);
nor U22826 (N_22826,N_22644,N_22501);
nor U22827 (N_22827,N_22523,N_22542);
and U22828 (N_22828,N_22661,N_22738);
and U22829 (N_22829,N_22674,N_22512);
and U22830 (N_22830,N_22610,N_22583);
nor U22831 (N_22831,N_22726,N_22516);
nor U22832 (N_22832,N_22696,N_22625);
or U22833 (N_22833,N_22730,N_22678);
or U22834 (N_22834,N_22606,N_22655);
nand U22835 (N_22835,N_22621,N_22618);
nand U22836 (N_22836,N_22677,N_22595);
and U22837 (N_22837,N_22634,N_22534);
nor U22838 (N_22838,N_22691,N_22711);
xnor U22839 (N_22839,N_22624,N_22500);
and U22840 (N_22840,N_22748,N_22548);
xor U22841 (N_22841,N_22603,N_22551);
xnor U22842 (N_22842,N_22599,N_22704);
or U22843 (N_22843,N_22570,N_22522);
or U22844 (N_22844,N_22558,N_22646);
and U22845 (N_22845,N_22667,N_22571);
or U22846 (N_22846,N_22588,N_22698);
nor U22847 (N_22847,N_22719,N_22602);
or U22848 (N_22848,N_22654,N_22565);
or U22849 (N_22849,N_22559,N_22720);
nor U22850 (N_22850,N_22532,N_22549);
nand U22851 (N_22851,N_22601,N_22633);
and U22852 (N_22852,N_22737,N_22627);
nand U22853 (N_22853,N_22538,N_22668);
and U22854 (N_22854,N_22690,N_22615);
nor U22855 (N_22855,N_22676,N_22741);
nor U22856 (N_22856,N_22681,N_22710);
and U22857 (N_22857,N_22569,N_22553);
nor U22858 (N_22858,N_22508,N_22585);
nand U22859 (N_22859,N_22657,N_22509);
or U22860 (N_22860,N_22643,N_22584);
or U22861 (N_22861,N_22652,N_22605);
or U22862 (N_22862,N_22728,N_22683);
and U22863 (N_22863,N_22722,N_22510);
or U22864 (N_22864,N_22686,N_22692);
or U22865 (N_22865,N_22513,N_22506);
nor U22866 (N_22866,N_22632,N_22529);
nor U22867 (N_22867,N_22638,N_22731);
or U22868 (N_22868,N_22689,N_22600);
or U22869 (N_22869,N_22703,N_22623);
xnor U22870 (N_22870,N_22629,N_22723);
nand U22871 (N_22871,N_22593,N_22663);
and U22872 (N_22872,N_22589,N_22639);
nor U22873 (N_22873,N_22701,N_22576);
nor U22874 (N_22874,N_22581,N_22743);
nand U22875 (N_22875,N_22704,N_22722);
xor U22876 (N_22876,N_22662,N_22538);
xor U22877 (N_22877,N_22582,N_22703);
and U22878 (N_22878,N_22674,N_22690);
and U22879 (N_22879,N_22722,N_22659);
nor U22880 (N_22880,N_22504,N_22695);
nand U22881 (N_22881,N_22607,N_22587);
or U22882 (N_22882,N_22681,N_22708);
xor U22883 (N_22883,N_22552,N_22647);
xor U22884 (N_22884,N_22639,N_22604);
nand U22885 (N_22885,N_22664,N_22691);
nor U22886 (N_22886,N_22529,N_22559);
or U22887 (N_22887,N_22599,N_22518);
or U22888 (N_22888,N_22702,N_22594);
xor U22889 (N_22889,N_22554,N_22633);
xor U22890 (N_22890,N_22561,N_22581);
and U22891 (N_22891,N_22520,N_22615);
nand U22892 (N_22892,N_22631,N_22619);
or U22893 (N_22893,N_22646,N_22637);
or U22894 (N_22894,N_22507,N_22619);
or U22895 (N_22895,N_22707,N_22553);
nand U22896 (N_22896,N_22544,N_22625);
or U22897 (N_22897,N_22607,N_22669);
and U22898 (N_22898,N_22532,N_22521);
and U22899 (N_22899,N_22616,N_22535);
nor U22900 (N_22900,N_22607,N_22642);
nand U22901 (N_22901,N_22743,N_22749);
nand U22902 (N_22902,N_22548,N_22728);
or U22903 (N_22903,N_22696,N_22589);
nor U22904 (N_22904,N_22594,N_22530);
xnor U22905 (N_22905,N_22558,N_22542);
nand U22906 (N_22906,N_22709,N_22552);
or U22907 (N_22907,N_22565,N_22636);
nand U22908 (N_22908,N_22652,N_22500);
or U22909 (N_22909,N_22676,N_22678);
nand U22910 (N_22910,N_22583,N_22649);
nand U22911 (N_22911,N_22707,N_22509);
and U22912 (N_22912,N_22610,N_22679);
or U22913 (N_22913,N_22652,N_22643);
nand U22914 (N_22914,N_22682,N_22737);
and U22915 (N_22915,N_22630,N_22542);
nor U22916 (N_22916,N_22669,N_22687);
nor U22917 (N_22917,N_22673,N_22572);
xor U22918 (N_22918,N_22737,N_22713);
nor U22919 (N_22919,N_22658,N_22692);
xor U22920 (N_22920,N_22614,N_22745);
or U22921 (N_22921,N_22664,N_22675);
or U22922 (N_22922,N_22716,N_22597);
and U22923 (N_22923,N_22693,N_22703);
or U22924 (N_22924,N_22613,N_22515);
or U22925 (N_22925,N_22703,N_22532);
or U22926 (N_22926,N_22532,N_22510);
or U22927 (N_22927,N_22574,N_22628);
and U22928 (N_22928,N_22700,N_22621);
nand U22929 (N_22929,N_22562,N_22549);
nor U22930 (N_22930,N_22509,N_22745);
xor U22931 (N_22931,N_22522,N_22651);
nand U22932 (N_22932,N_22739,N_22669);
and U22933 (N_22933,N_22718,N_22733);
nand U22934 (N_22934,N_22544,N_22611);
xor U22935 (N_22935,N_22533,N_22620);
nor U22936 (N_22936,N_22544,N_22609);
nor U22937 (N_22937,N_22661,N_22571);
nand U22938 (N_22938,N_22652,N_22602);
and U22939 (N_22939,N_22719,N_22664);
xor U22940 (N_22940,N_22700,N_22744);
or U22941 (N_22941,N_22621,N_22570);
nand U22942 (N_22942,N_22727,N_22579);
nor U22943 (N_22943,N_22623,N_22690);
and U22944 (N_22944,N_22534,N_22597);
nor U22945 (N_22945,N_22737,N_22628);
or U22946 (N_22946,N_22579,N_22684);
and U22947 (N_22947,N_22572,N_22670);
xor U22948 (N_22948,N_22609,N_22625);
and U22949 (N_22949,N_22663,N_22744);
or U22950 (N_22950,N_22549,N_22685);
and U22951 (N_22951,N_22510,N_22534);
xnor U22952 (N_22952,N_22525,N_22611);
nand U22953 (N_22953,N_22683,N_22525);
or U22954 (N_22954,N_22650,N_22619);
xor U22955 (N_22955,N_22716,N_22673);
xnor U22956 (N_22956,N_22609,N_22655);
xor U22957 (N_22957,N_22597,N_22570);
or U22958 (N_22958,N_22732,N_22588);
nor U22959 (N_22959,N_22552,N_22596);
nor U22960 (N_22960,N_22588,N_22645);
nand U22961 (N_22961,N_22614,N_22643);
nor U22962 (N_22962,N_22625,N_22536);
nor U22963 (N_22963,N_22602,N_22600);
nand U22964 (N_22964,N_22708,N_22723);
nor U22965 (N_22965,N_22637,N_22679);
and U22966 (N_22966,N_22693,N_22674);
nor U22967 (N_22967,N_22649,N_22744);
and U22968 (N_22968,N_22624,N_22557);
nand U22969 (N_22969,N_22561,N_22593);
nand U22970 (N_22970,N_22519,N_22593);
nand U22971 (N_22971,N_22615,N_22550);
and U22972 (N_22972,N_22643,N_22612);
xnor U22973 (N_22973,N_22617,N_22692);
and U22974 (N_22974,N_22705,N_22675);
or U22975 (N_22975,N_22690,N_22597);
and U22976 (N_22976,N_22733,N_22742);
xnor U22977 (N_22977,N_22748,N_22608);
or U22978 (N_22978,N_22660,N_22733);
and U22979 (N_22979,N_22629,N_22576);
nor U22980 (N_22980,N_22655,N_22564);
or U22981 (N_22981,N_22581,N_22630);
or U22982 (N_22982,N_22548,N_22665);
or U22983 (N_22983,N_22726,N_22528);
nand U22984 (N_22984,N_22619,N_22626);
and U22985 (N_22985,N_22575,N_22504);
xnor U22986 (N_22986,N_22643,N_22557);
nand U22987 (N_22987,N_22518,N_22656);
nand U22988 (N_22988,N_22708,N_22617);
xor U22989 (N_22989,N_22580,N_22708);
nor U22990 (N_22990,N_22662,N_22573);
nand U22991 (N_22991,N_22512,N_22644);
and U22992 (N_22992,N_22503,N_22512);
and U22993 (N_22993,N_22581,N_22583);
and U22994 (N_22994,N_22531,N_22726);
xnor U22995 (N_22995,N_22741,N_22598);
nand U22996 (N_22996,N_22705,N_22706);
xnor U22997 (N_22997,N_22623,N_22673);
xor U22998 (N_22998,N_22569,N_22540);
nand U22999 (N_22999,N_22706,N_22608);
nor U23000 (N_23000,N_22892,N_22822);
and U23001 (N_23001,N_22810,N_22828);
xnor U23002 (N_23002,N_22751,N_22921);
nor U23003 (N_23003,N_22850,N_22952);
nor U23004 (N_23004,N_22972,N_22969);
nor U23005 (N_23005,N_22791,N_22939);
or U23006 (N_23006,N_22855,N_22876);
and U23007 (N_23007,N_22973,N_22879);
nor U23008 (N_23008,N_22845,N_22956);
nor U23009 (N_23009,N_22912,N_22753);
xnor U23010 (N_23010,N_22967,N_22918);
xnor U23011 (N_23011,N_22861,N_22780);
xnor U23012 (N_23012,N_22786,N_22976);
nand U23013 (N_23013,N_22768,N_22797);
and U23014 (N_23014,N_22989,N_22925);
and U23015 (N_23015,N_22983,N_22994);
or U23016 (N_23016,N_22992,N_22763);
xor U23017 (N_23017,N_22764,N_22790);
and U23018 (N_23018,N_22907,N_22834);
nand U23019 (N_23019,N_22995,N_22801);
and U23020 (N_23020,N_22888,N_22777);
nor U23021 (N_23021,N_22882,N_22891);
xnor U23022 (N_23022,N_22755,N_22756);
and U23023 (N_23023,N_22830,N_22928);
xor U23024 (N_23024,N_22893,N_22905);
xor U23025 (N_23025,N_22958,N_22833);
or U23026 (N_23026,N_22919,N_22843);
nand U23027 (N_23027,N_22975,N_22785);
nand U23028 (N_23028,N_22949,N_22951);
and U23029 (N_23029,N_22823,N_22955);
nand U23030 (N_23030,N_22881,N_22897);
nand U23031 (N_23031,N_22904,N_22803);
xor U23032 (N_23032,N_22775,N_22903);
nor U23033 (N_23033,N_22809,N_22926);
or U23034 (N_23034,N_22761,N_22872);
nor U23035 (N_23035,N_22963,N_22874);
or U23036 (N_23036,N_22946,N_22851);
and U23037 (N_23037,N_22829,N_22859);
or U23038 (N_23038,N_22864,N_22767);
nor U23039 (N_23039,N_22922,N_22853);
nand U23040 (N_23040,N_22752,N_22932);
nor U23041 (N_23041,N_22831,N_22844);
xnor U23042 (N_23042,N_22782,N_22978);
xor U23043 (N_23043,N_22915,N_22865);
nand U23044 (N_23044,N_22981,N_22986);
nor U23045 (N_23045,N_22911,N_22894);
nor U23046 (N_23046,N_22940,N_22999);
and U23047 (N_23047,N_22982,N_22880);
or U23048 (N_23048,N_22910,N_22793);
and U23049 (N_23049,N_22868,N_22759);
nand U23050 (N_23050,N_22870,N_22877);
nor U23051 (N_23051,N_22953,N_22837);
or U23052 (N_23052,N_22862,N_22750);
and U23053 (N_23053,N_22947,N_22798);
nand U23054 (N_23054,N_22984,N_22966);
nor U23055 (N_23055,N_22991,N_22887);
nor U23056 (N_23056,N_22902,N_22799);
xor U23057 (N_23057,N_22979,N_22889);
xor U23058 (N_23058,N_22962,N_22895);
xor U23059 (N_23059,N_22890,N_22977);
nand U23060 (N_23060,N_22800,N_22929);
xnor U23061 (N_23061,N_22770,N_22885);
nor U23062 (N_23062,N_22954,N_22804);
or U23063 (N_23063,N_22988,N_22916);
nor U23064 (N_23064,N_22771,N_22818);
nand U23065 (N_23065,N_22993,N_22847);
and U23066 (N_23066,N_22838,N_22985);
nand U23067 (N_23067,N_22987,N_22772);
and U23068 (N_23068,N_22816,N_22937);
nand U23069 (N_23069,N_22835,N_22812);
nand U23070 (N_23070,N_22779,N_22968);
nor U23071 (N_23071,N_22927,N_22943);
and U23072 (N_23072,N_22974,N_22825);
or U23073 (N_23073,N_22832,N_22839);
xnor U23074 (N_23074,N_22841,N_22866);
or U23075 (N_23075,N_22842,N_22965);
nand U23076 (N_23076,N_22899,N_22858);
or U23077 (N_23077,N_22774,N_22900);
and U23078 (N_23078,N_22819,N_22941);
and U23079 (N_23079,N_22871,N_22964);
xor U23080 (N_23080,N_22781,N_22909);
and U23081 (N_23081,N_22827,N_22802);
nor U23082 (N_23082,N_22971,N_22863);
nor U23083 (N_23083,N_22826,N_22934);
or U23084 (N_23084,N_22784,N_22917);
xor U23085 (N_23085,N_22938,N_22787);
and U23086 (N_23086,N_22970,N_22997);
xnor U23087 (N_23087,N_22908,N_22950);
and U23088 (N_23088,N_22860,N_22886);
nand U23089 (N_23089,N_22896,N_22852);
xnor U23090 (N_23090,N_22788,N_22758);
nor U23091 (N_23091,N_22901,N_22854);
nand U23092 (N_23092,N_22945,N_22898);
or U23093 (N_23093,N_22933,N_22808);
nand U23094 (N_23094,N_22796,N_22765);
and U23095 (N_23095,N_22875,N_22878);
and U23096 (N_23096,N_22840,N_22960);
and U23097 (N_23097,N_22913,N_22998);
or U23098 (N_23098,N_22873,N_22980);
nand U23099 (N_23099,N_22884,N_22856);
and U23100 (N_23100,N_22957,N_22923);
nor U23101 (N_23101,N_22883,N_22857);
xnor U23102 (N_23102,N_22959,N_22813);
nand U23103 (N_23103,N_22776,N_22773);
nand U23104 (N_23104,N_22867,N_22848);
or U23105 (N_23105,N_22783,N_22906);
nor U23106 (N_23106,N_22944,N_22930);
and U23107 (N_23107,N_22757,N_22920);
or U23108 (N_23108,N_22805,N_22778);
or U23109 (N_23109,N_22942,N_22760);
or U23110 (N_23110,N_22914,N_22849);
and U23111 (N_23111,N_22807,N_22811);
or U23112 (N_23112,N_22806,N_22846);
nor U23113 (N_23113,N_22936,N_22794);
or U23114 (N_23114,N_22766,N_22931);
or U23115 (N_23115,N_22769,N_22792);
nand U23116 (N_23116,N_22836,N_22948);
nor U23117 (N_23117,N_22935,N_22824);
and U23118 (N_23118,N_22789,N_22924);
or U23119 (N_23119,N_22817,N_22869);
or U23120 (N_23120,N_22821,N_22795);
and U23121 (N_23121,N_22996,N_22762);
nor U23122 (N_23122,N_22820,N_22815);
or U23123 (N_23123,N_22814,N_22990);
nor U23124 (N_23124,N_22754,N_22961);
xor U23125 (N_23125,N_22789,N_22980);
and U23126 (N_23126,N_22885,N_22797);
nor U23127 (N_23127,N_22921,N_22917);
nand U23128 (N_23128,N_22906,N_22985);
nor U23129 (N_23129,N_22948,N_22817);
or U23130 (N_23130,N_22851,N_22818);
nand U23131 (N_23131,N_22888,N_22835);
nor U23132 (N_23132,N_22805,N_22903);
or U23133 (N_23133,N_22841,N_22918);
nor U23134 (N_23134,N_22805,N_22897);
or U23135 (N_23135,N_22791,N_22976);
and U23136 (N_23136,N_22949,N_22776);
xnor U23137 (N_23137,N_22789,N_22853);
and U23138 (N_23138,N_22896,N_22764);
and U23139 (N_23139,N_22963,N_22840);
xnor U23140 (N_23140,N_22812,N_22994);
and U23141 (N_23141,N_22959,N_22894);
and U23142 (N_23142,N_22975,N_22968);
nor U23143 (N_23143,N_22907,N_22790);
nand U23144 (N_23144,N_22783,N_22838);
or U23145 (N_23145,N_22791,N_22942);
nor U23146 (N_23146,N_22774,N_22934);
or U23147 (N_23147,N_22924,N_22872);
or U23148 (N_23148,N_22861,N_22890);
nor U23149 (N_23149,N_22849,N_22880);
nand U23150 (N_23150,N_22816,N_22813);
nor U23151 (N_23151,N_22759,N_22991);
nor U23152 (N_23152,N_22906,N_22866);
and U23153 (N_23153,N_22990,N_22829);
nand U23154 (N_23154,N_22863,N_22838);
or U23155 (N_23155,N_22975,N_22822);
or U23156 (N_23156,N_22853,N_22883);
nor U23157 (N_23157,N_22797,N_22782);
nor U23158 (N_23158,N_22833,N_22844);
or U23159 (N_23159,N_22790,N_22999);
and U23160 (N_23160,N_22982,N_22821);
xnor U23161 (N_23161,N_22861,N_22793);
nor U23162 (N_23162,N_22827,N_22983);
nor U23163 (N_23163,N_22982,N_22917);
and U23164 (N_23164,N_22847,N_22937);
and U23165 (N_23165,N_22887,N_22816);
nor U23166 (N_23166,N_22824,N_22971);
or U23167 (N_23167,N_22992,N_22912);
and U23168 (N_23168,N_22788,N_22800);
nand U23169 (N_23169,N_22997,N_22836);
xnor U23170 (N_23170,N_22934,N_22831);
xnor U23171 (N_23171,N_22858,N_22938);
xnor U23172 (N_23172,N_22770,N_22964);
or U23173 (N_23173,N_22905,N_22973);
xnor U23174 (N_23174,N_22772,N_22853);
nand U23175 (N_23175,N_22910,N_22769);
or U23176 (N_23176,N_22991,N_22982);
xnor U23177 (N_23177,N_22784,N_22794);
nand U23178 (N_23178,N_22759,N_22760);
xor U23179 (N_23179,N_22763,N_22944);
nand U23180 (N_23180,N_22978,N_22887);
xnor U23181 (N_23181,N_22945,N_22843);
nand U23182 (N_23182,N_22774,N_22781);
nand U23183 (N_23183,N_22885,N_22944);
and U23184 (N_23184,N_22887,N_22881);
or U23185 (N_23185,N_22857,N_22841);
nand U23186 (N_23186,N_22945,N_22963);
nor U23187 (N_23187,N_22866,N_22946);
xnor U23188 (N_23188,N_22750,N_22973);
nand U23189 (N_23189,N_22989,N_22981);
or U23190 (N_23190,N_22870,N_22964);
nor U23191 (N_23191,N_22902,N_22772);
nand U23192 (N_23192,N_22898,N_22856);
and U23193 (N_23193,N_22958,N_22915);
nor U23194 (N_23194,N_22964,N_22767);
or U23195 (N_23195,N_22949,N_22991);
nor U23196 (N_23196,N_22783,N_22896);
nor U23197 (N_23197,N_22892,N_22936);
nand U23198 (N_23198,N_22779,N_22786);
xor U23199 (N_23199,N_22964,N_22780);
xor U23200 (N_23200,N_22962,N_22792);
nor U23201 (N_23201,N_22772,N_22759);
nand U23202 (N_23202,N_22981,N_22806);
nor U23203 (N_23203,N_22835,N_22969);
and U23204 (N_23204,N_22928,N_22826);
nor U23205 (N_23205,N_22778,N_22974);
and U23206 (N_23206,N_22927,N_22850);
nor U23207 (N_23207,N_22886,N_22808);
xnor U23208 (N_23208,N_22787,N_22822);
and U23209 (N_23209,N_22830,N_22911);
or U23210 (N_23210,N_22876,N_22805);
xor U23211 (N_23211,N_22989,N_22947);
and U23212 (N_23212,N_22829,N_22790);
xor U23213 (N_23213,N_22757,N_22861);
xnor U23214 (N_23214,N_22757,N_22785);
nor U23215 (N_23215,N_22758,N_22833);
or U23216 (N_23216,N_22975,N_22862);
nor U23217 (N_23217,N_22884,N_22991);
nor U23218 (N_23218,N_22963,N_22962);
nand U23219 (N_23219,N_22767,N_22995);
nand U23220 (N_23220,N_22975,N_22864);
or U23221 (N_23221,N_22839,N_22852);
nand U23222 (N_23222,N_22879,N_22822);
xor U23223 (N_23223,N_22962,N_22884);
nand U23224 (N_23224,N_22817,N_22964);
and U23225 (N_23225,N_22851,N_22901);
xor U23226 (N_23226,N_22914,N_22968);
nor U23227 (N_23227,N_22855,N_22752);
and U23228 (N_23228,N_22954,N_22757);
and U23229 (N_23229,N_22889,N_22871);
or U23230 (N_23230,N_22775,N_22762);
nor U23231 (N_23231,N_22768,N_22793);
xor U23232 (N_23232,N_22968,N_22908);
and U23233 (N_23233,N_22985,N_22886);
xnor U23234 (N_23234,N_22800,N_22907);
nand U23235 (N_23235,N_22972,N_22769);
nand U23236 (N_23236,N_22984,N_22938);
nand U23237 (N_23237,N_22754,N_22839);
nor U23238 (N_23238,N_22925,N_22827);
nor U23239 (N_23239,N_22760,N_22880);
and U23240 (N_23240,N_22793,N_22938);
nand U23241 (N_23241,N_22885,N_22800);
and U23242 (N_23242,N_22840,N_22939);
nand U23243 (N_23243,N_22865,N_22890);
or U23244 (N_23244,N_22832,N_22831);
and U23245 (N_23245,N_22883,N_22772);
nand U23246 (N_23246,N_22828,N_22774);
or U23247 (N_23247,N_22766,N_22832);
nor U23248 (N_23248,N_22835,N_22972);
nor U23249 (N_23249,N_22775,N_22804);
xor U23250 (N_23250,N_23217,N_23189);
or U23251 (N_23251,N_23243,N_23050);
or U23252 (N_23252,N_23177,N_23114);
xor U23253 (N_23253,N_23150,N_23090);
nand U23254 (N_23254,N_23021,N_23009);
nor U23255 (N_23255,N_23010,N_23218);
and U23256 (N_23256,N_23229,N_23124);
xnor U23257 (N_23257,N_23220,N_23111);
nor U23258 (N_23258,N_23226,N_23160);
nor U23259 (N_23259,N_23195,N_23015);
or U23260 (N_23260,N_23076,N_23056);
or U23261 (N_23261,N_23247,N_23181);
nor U23262 (N_23262,N_23062,N_23190);
nand U23263 (N_23263,N_23157,N_23137);
or U23264 (N_23264,N_23162,N_23216);
nor U23265 (N_23265,N_23144,N_23075);
nand U23266 (N_23266,N_23054,N_23183);
xnor U23267 (N_23267,N_23240,N_23151);
xor U23268 (N_23268,N_23210,N_23084);
nor U23269 (N_23269,N_23244,N_23000);
nand U23270 (N_23270,N_23055,N_23155);
nand U23271 (N_23271,N_23225,N_23023);
nand U23272 (N_23272,N_23047,N_23078);
xor U23273 (N_23273,N_23202,N_23207);
or U23274 (N_23274,N_23239,N_23067);
xnor U23275 (N_23275,N_23208,N_23081);
and U23276 (N_23276,N_23206,N_23074);
or U23277 (N_23277,N_23094,N_23203);
and U23278 (N_23278,N_23173,N_23199);
nand U23279 (N_23279,N_23200,N_23082);
and U23280 (N_23280,N_23110,N_23066);
nor U23281 (N_23281,N_23099,N_23107);
and U23282 (N_23282,N_23087,N_23073);
xor U23283 (N_23283,N_23104,N_23233);
nand U23284 (N_23284,N_23086,N_23105);
nand U23285 (N_23285,N_23168,N_23201);
and U23286 (N_23286,N_23014,N_23020);
and U23287 (N_23287,N_23169,N_23095);
nor U23288 (N_23288,N_23184,N_23120);
and U23289 (N_23289,N_23235,N_23034);
xor U23290 (N_23290,N_23209,N_23089);
and U23291 (N_23291,N_23215,N_23079);
nor U23292 (N_23292,N_23163,N_23012);
nand U23293 (N_23293,N_23143,N_23222);
nor U23294 (N_23294,N_23064,N_23057);
and U23295 (N_23295,N_23098,N_23007);
nor U23296 (N_23296,N_23039,N_23140);
or U23297 (N_23297,N_23061,N_23172);
and U23298 (N_23298,N_23028,N_23156);
and U23299 (N_23299,N_23042,N_23219);
or U23300 (N_23300,N_23128,N_23170);
or U23301 (N_23301,N_23092,N_23179);
nand U23302 (N_23302,N_23204,N_23176);
nor U23303 (N_23303,N_23213,N_23122);
nor U23304 (N_23304,N_23123,N_23138);
nand U23305 (N_23305,N_23018,N_23148);
nand U23306 (N_23306,N_23024,N_23125);
nand U23307 (N_23307,N_23016,N_23129);
or U23308 (N_23308,N_23234,N_23197);
and U23309 (N_23309,N_23097,N_23117);
or U23310 (N_23310,N_23165,N_23040);
and U23311 (N_23311,N_23035,N_23146);
and U23312 (N_23312,N_23205,N_23223);
nor U23313 (N_23313,N_23025,N_23060);
nand U23314 (N_23314,N_23112,N_23096);
and U23315 (N_23315,N_23019,N_23182);
nor U23316 (N_23316,N_23232,N_23193);
nor U23317 (N_23317,N_23053,N_23051);
nand U23318 (N_23318,N_23154,N_23116);
or U23319 (N_23319,N_23109,N_23198);
nand U23320 (N_23320,N_23049,N_23006);
nand U23321 (N_23321,N_23072,N_23131);
and U23322 (N_23322,N_23118,N_23139);
nor U23323 (N_23323,N_23041,N_23212);
nand U23324 (N_23324,N_23101,N_23103);
nor U23325 (N_23325,N_23153,N_23065);
nor U23326 (N_23326,N_23026,N_23071);
xor U23327 (N_23327,N_23242,N_23052);
and U23328 (N_23328,N_23248,N_23038);
nand U23329 (N_23329,N_23017,N_23088);
xnor U23330 (N_23330,N_23147,N_23091);
nand U23331 (N_23331,N_23180,N_23048);
nor U23332 (N_23332,N_23191,N_23126);
xnor U23333 (N_23333,N_23186,N_23036);
nand U23334 (N_23334,N_23164,N_23136);
and U23335 (N_23335,N_23241,N_23158);
or U23336 (N_23336,N_23085,N_23211);
and U23337 (N_23337,N_23069,N_23002);
nor U23338 (N_23338,N_23231,N_23106);
nand U23339 (N_23339,N_23115,N_23196);
and U23340 (N_23340,N_23119,N_23044);
xnor U23341 (N_23341,N_23004,N_23030);
xor U23342 (N_23342,N_23022,N_23192);
and U23343 (N_23343,N_23077,N_23174);
nor U23344 (N_23344,N_23133,N_23063);
xor U23345 (N_23345,N_23142,N_23031);
and U23346 (N_23346,N_23058,N_23068);
nand U23347 (N_23347,N_23221,N_23132);
and U23348 (N_23348,N_23008,N_23245);
or U23349 (N_23349,N_23166,N_23230);
and U23350 (N_23350,N_23001,N_23224);
nand U23351 (N_23351,N_23045,N_23043);
nor U23352 (N_23352,N_23037,N_23130);
xnor U23353 (N_23353,N_23171,N_23059);
or U23354 (N_23354,N_23227,N_23100);
xor U23355 (N_23355,N_23033,N_23194);
nand U23356 (N_23356,N_23187,N_23159);
nor U23357 (N_23357,N_23228,N_23003);
nor U23358 (N_23358,N_23121,N_23178);
nor U23359 (N_23359,N_23236,N_23141);
xnor U23360 (N_23360,N_23134,N_23102);
and U23361 (N_23361,N_23027,N_23249);
nor U23362 (N_23362,N_23167,N_23032);
or U23363 (N_23363,N_23029,N_23185);
nand U23364 (N_23364,N_23135,N_23011);
or U23365 (N_23365,N_23005,N_23083);
or U23366 (N_23366,N_23113,N_23093);
xor U23367 (N_23367,N_23175,N_23127);
or U23368 (N_23368,N_23108,N_23149);
nor U23369 (N_23369,N_23161,N_23238);
nor U23370 (N_23370,N_23214,N_23080);
nor U23371 (N_23371,N_23070,N_23013);
or U23372 (N_23372,N_23188,N_23152);
xor U23373 (N_23373,N_23046,N_23145);
xnor U23374 (N_23374,N_23246,N_23237);
xnor U23375 (N_23375,N_23058,N_23147);
and U23376 (N_23376,N_23181,N_23095);
nand U23377 (N_23377,N_23048,N_23060);
or U23378 (N_23378,N_23057,N_23193);
and U23379 (N_23379,N_23122,N_23099);
or U23380 (N_23380,N_23158,N_23115);
xor U23381 (N_23381,N_23023,N_23012);
xor U23382 (N_23382,N_23161,N_23222);
nand U23383 (N_23383,N_23036,N_23205);
nor U23384 (N_23384,N_23218,N_23153);
or U23385 (N_23385,N_23057,N_23161);
nand U23386 (N_23386,N_23150,N_23117);
and U23387 (N_23387,N_23055,N_23104);
or U23388 (N_23388,N_23076,N_23214);
nand U23389 (N_23389,N_23120,N_23037);
or U23390 (N_23390,N_23078,N_23069);
or U23391 (N_23391,N_23214,N_23040);
and U23392 (N_23392,N_23056,N_23080);
and U23393 (N_23393,N_23039,N_23172);
xnor U23394 (N_23394,N_23074,N_23195);
nor U23395 (N_23395,N_23222,N_23041);
nor U23396 (N_23396,N_23005,N_23062);
and U23397 (N_23397,N_23171,N_23099);
and U23398 (N_23398,N_23013,N_23189);
nand U23399 (N_23399,N_23092,N_23135);
or U23400 (N_23400,N_23095,N_23005);
xor U23401 (N_23401,N_23092,N_23058);
nor U23402 (N_23402,N_23085,N_23129);
xor U23403 (N_23403,N_23022,N_23090);
or U23404 (N_23404,N_23028,N_23186);
xor U23405 (N_23405,N_23111,N_23153);
nand U23406 (N_23406,N_23038,N_23033);
nand U23407 (N_23407,N_23186,N_23111);
xnor U23408 (N_23408,N_23110,N_23045);
xnor U23409 (N_23409,N_23208,N_23045);
and U23410 (N_23410,N_23239,N_23125);
and U23411 (N_23411,N_23123,N_23093);
or U23412 (N_23412,N_23123,N_23059);
nor U23413 (N_23413,N_23199,N_23133);
nand U23414 (N_23414,N_23243,N_23178);
and U23415 (N_23415,N_23239,N_23196);
nand U23416 (N_23416,N_23168,N_23171);
or U23417 (N_23417,N_23180,N_23043);
nand U23418 (N_23418,N_23087,N_23119);
nand U23419 (N_23419,N_23232,N_23140);
and U23420 (N_23420,N_23034,N_23152);
and U23421 (N_23421,N_23020,N_23022);
xor U23422 (N_23422,N_23114,N_23168);
or U23423 (N_23423,N_23014,N_23160);
or U23424 (N_23424,N_23175,N_23106);
xnor U23425 (N_23425,N_23244,N_23231);
or U23426 (N_23426,N_23153,N_23119);
or U23427 (N_23427,N_23239,N_23039);
nand U23428 (N_23428,N_23220,N_23159);
or U23429 (N_23429,N_23096,N_23216);
nand U23430 (N_23430,N_23149,N_23236);
xor U23431 (N_23431,N_23123,N_23238);
and U23432 (N_23432,N_23102,N_23150);
and U23433 (N_23433,N_23221,N_23076);
nor U23434 (N_23434,N_23237,N_23005);
and U23435 (N_23435,N_23129,N_23248);
xnor U23436 (N_23436,N_23192,N_23136);
and U23437 (N_23437,N_23129,N_23203);
nor U23438 (N_23438,N_23184,N_23060);
and U23439 (N_23439,N_23105,N_23170);
or U23440 (N_23440,N_23131,N_23078);
xor U23441 (N_23441,N_23032,N_23220);
xnor U23442 (N_23442,N_23216,N_23175);
nand U23443 (N_23443,N_23146,N_23098);
nor U23444 (N_23444,N_23240,N_23058);
or U23445 (N_23445,N_23048,N_23059);
nor U23446 (N_23446,N_23160,N_23024);
xnor U23447 (N_23447,N_23072,N_23119);
xor U23448 (N_23448,N_23246,N_23025);
nand U23449 (N_23449,N_23050,N_23028);
or U23450 (N_23450,N_23156,N_23113);
or U23451 (N_23451,N_23127,N_23138);
nand U23452 (N_23452,N_23153,N_23123);
nor U23453 (N_23453,N_23131,N_23182);
or U23454 (N_23454,N_23073,N_23138);
and U23455 (N_23455,N_23171,N_23128);
xor U23456 (N_23456,N_23113,N_23110);
nor U23457 (N_23457,N_23119,N_23163);
nor U23458 (N_23458,N_23098,N_23202);
or U23459 (N_23459,N_23131,N_23137);
xor U23460 (N_23460,N_23153,N_23108);
or U23461 (N_23461,N_23103,N_23121);
and U23462 (N_23462,N_23191,N_23174);
xnor U23463 (N_23463,N_23064,N_23048);
nand U23464 (N_23464,N_23128,N_23216);
xnor U23465 (N_23465,N_23189,N_23233);
nor U23466 (N_23466,N_23114,N_23059);
nand U23467 (N_23467,N_23247,N_23191);
xor U23468 (N_23468,N_23030,N_23039);
or U23469 (N_23469,N_23054,N_23023);
and U23470 (N_23470,N_23058,N_23125);
xnor U23471 (N_23471,N_23105,N_23042);
nor U23472 (N_23472,N_23073,N_23083);
and U23473 (N_23473,N_23164,N_23170);
and U23474 (N_23474,N_23148,N_23198);
xor U23475 (N_23475,N_23158,N_23119);
nor U23476 (N_23476,N_23133,N_23028);
nor U23477 (N_23477,N_23074,N_23121);
and U23478 (N_23478,N_23062,N_23247);
nor U23479 (N_23479,N_23071,N_23165);
nand U23480 (N_23480,N_23051,N_23126);
nand U23481 (N_23481,N_23123,N_23074);
or U23482 (N_23482,N_23084,N_23079);
nor U23483 (N_23483,N_23086,N_23070);
and U23484 (N_23484,N_23095,N_23124);
nor U23485 (N_23485,N_23214,N_23098);
nand U23486 (N_23486,N_23036,N_23006);
xnor U23487 (N_23487,N_23222,N_23195);
nor U23488 (N_23488,N_23016,N_23122);
nor U23489 (N_23489,N_23188,N_23085);
and U23490 (N_23490,N_23102,N_23215);
nor U23491 (N_23491,N_23072,N_23020);
nor U23492 (N_23492,N_23085,N_23100);
and U23493 (N_23493,N_23138,N_23174);
xnor U23494 (N_23494,N_23053,N_23005);
and U23495 (N_23495,N_23229,N_23214);
nand U23496 (N_23496,N_23177,N_23243);
and U23497 (N_23497,N_23247,N_23046);
xnor U23498 (N_23498,N_23123,N_23184);
nand U23499 (N_23499,N_23163,N_23213);
or U23500 (N_23500,N_23385,N_23365);
nand U23501 (N_23501,N_23474,N_23269);
and U23502 (N_23502,N_23329,N_23302);
xnor U23503 (N_23503,N_23341,N_23340);
nand U23504 (N_23504,N_23483,N_23425);
nand U23505 (N_23505,N_23428,N_23421);
nor U23506 (N_23506,N_23306,N_23430);
xnor U23507 (N_23507,N_23445,N_23331);
or U23508 (N_23508,N_23380,N_23486);
and U23509 (N_23509,N_23360,N_23358);
or U23510 (N_23510,N_23296,N_23351);
xnor U23511 (N_23511,N_23357,N_23451);
nand U23512 (N_23512,N_23462,N_23459);
xor U23513 (N_23513,N_23333,N_23490);
or U23514 (N_23514,N_23390,N_23497);
or U23515 (N_23515,N_23349,N_23374);
nand U23516 (N_23516,N_23312,N_23378);
xor U23517 (N_23517,N_23263,N_23498);
nand U23518 (N_23518,N_23373,N_23308);
or U23519 (N_23519,N_23447,N_23408);
and U23520 (N_23520,N_23326,N_23250);
nand U23521 (N_23521,N_23295,N_23411);
xor U23522 (N_23522,N_23476,N_23396);
nor U23523 (N_23523,N_23362,N_23376);
or U23524 (N_23524,N_23482,N_23298);
xnor U23525 (N_23525,N_23437,N_23310);
and U23526 (N_23526,N_23400,N_23379);
nor U23527 (N_23527,N_23499,N_23332);
xnor U23528 (N_23528,N_23330,N_23352);
nand U23529 (N_23529,N_23392,N_23276);
or U23530 (N_23530,N_23288,N_23261);
xor U23531 (N_23531,N_23475,N_23456);
or U23532 (N_23532,N_23264,N_23265);
xor U23533 (N_23533,N_23485,N_23252);
nor U23534 (N_23534,N_23466,N_23383);
or U23535 (N_23535,N_23367,N_23393);
xnor U23536 (N_23536,N_23300,N_23453);
xor U23537 (N_23537,N_23464,N_23345);
or U23538 (N_23538,N_23371,N_23304);
nand U23539 (N_23539,N_23309,N_23446);
nor U23540 (N_23540,N_23450,N_23424);
nand U23541 (N_23541,N_23460,N_23394);
or U23542 (N_23542,N_23412,N_23384);
xor U23543 (N_23543,N_23353,N_23282);
and U23544 (N_23544,N_23364,N_23468);
xnor U23545 (N_23545,N_23318,N_23470);
nand U23546 (N_23546,N_23325,N_23492);
nor U23547 (N_23547,N_23431,N_23439);
or U23548 (N_23548,N_23496,N_23471);
xnor U23549 (N_23549,N_23368,N_23448);
xor U23550 (N_23550,N_23323,N_23370);
xor U23551 (N_23551,N_23372,N_23290);
nand U23552 (N_23552,N_23423,N_23401);
or U23553 (N_23553,N_23488,N_23443);
nand U23554 (N_23554,N_23441,N_23277);
or U23555 (N_23555,N_23472,N_23399);
nor U23556 (N_23556,N_23435,N_23343);
and U23557 (N_23557,N_23285,N_23275);
and U23558 (N_23558,N_23274,N_23256);
xor U23559 (N_23559,N_23494,N_23484);
xnor U23560 (N_23560,N_23272,N_23418);
nor U23561 (N_23561,N_23444,N_23283);
nand U23562 (N_23562,N_23317,N_23322);
and U23563 (N_23563,N_23432,N_23416);
or U23564 (N_23564,N_23347,N_23386);
nand U23565 (N_23565,N_23398,N_23388);
xnor U23566 (N_23566,N_23406,N_23355);
and U23567 (N_23567,N_23307,N_23342);
and U23568 (N_23568,N_23415,N_23420);
and U23569 (N_23569,N_23449,N_23452);
xor U23570 (N_23570,N_23267,N_23363);
nand U23571 (N_23571,N_23426,N_23395);
nor U23572 (N_23572,N_23389,N_23324);
nand U23573 (N_23573,N_23480,N_23427);
nand U23574 (N_23574,N_23478,N_23293);
nand U23575 (N_23575,N_23305,N_23258);
nor U23576 (N_23576,N_23254,N_23413);
xor U23577 (N_23577,N_23417,N_23438);
or U23578 (N_23578,N_23377,N_23260);
or U23579 (N_23579,N_23461,N_23436);
xor U23580 (N_23580,N_23495,N_23259);
xnor U23581 (N_23581,N_23409,N_23405);
and U23582 (N_23582,N_23348,N_23422);
xnor U23583 (N_23583,N_23489,N_23316);
nand U23584 (N_23584,N_23279,N_23284);
nand U23585 (N_23585,N_23253,N_23434);
nor U23586 (N_23586,N_23356,N_23465);
nor U23587 (N_23587,N_23366,N_23271);
nand U23588 (N_23588,N_23354,N_23287);
nor U23589 (N_23589,N_23402,N_23257);
nor U23590 (N_23590,N_23294,N_23419);
or U23591 (N_23591,N_23391,N_23381);
and U23592 (N_23592,N_23336,N_23369);
nand U23593 (N_23593,N_23328,N_23289);
nor U23594 (N_23594,N_23350,N_23255);
or U23595 (N_23595,N_23442,N_23278);
or U23596 (N_23596,N_23433,N_23491);
and U23597 (N_23597,N_23291,N_23280);
nor U23598 (N_23598,N_23397,N_23320);
nor U23599 (N_23599,N_23338,N_23321);
nor U23600 (N_23600,N_23493,N_23457);
or U23601 (N_23601,N_23327,N_23481);
nor U23602 (N_23602,N_23281,N_23458);
nor U23603 (N_23603,N_23311,N_23335);
or U23604 (N_23604,N_23266,N_23315);
or U23605 (N_23605,N_23334,N_23262);
and U23606 (N_23606,N_23314,N_23455);
or U23607 (N_23607,N_23410,N_23251);
or U23608 (N_23608,N_23403,N_23467);
xnor U23609 (N_23609,N_23404,N_23473);
or U23610 (N_23610,N_23286,N_23297);
nand U23611 (N_23611,N_23414,N_23292);
nand U23612 (N_23612,N_23382,N_23299);
nor U23613 (N_23613,N_23303,N_23387);
nor U23614 (N_23614,N_23454,N_23429);
nor U23615 (N_23615,N_23479,N_23313);
or U23616 (N_23616,N_23301,N_23270);
nand U23617 (N_23617,N_23319,N_23440);
nor U23618 (N_23618,N_23407,N_23344);
nand U23619 (N_23619,N_23339,N_23477);
nand U23620 (N_23620,N_23375,N_23337);
nor U23621 (N_23621,N_23361,N_23268);
nor U23622 (N_23622,N_23487,N_23359);
and U23623 (N_23623,N_23463,N_23469);
and U23624 (N_23624,N_23273,N_23346);
nor U23625 (N_23625,N_23431,N_23316);
or U23626 (N_23626,N_23332,N_23325);
and U23627 (N_23627,N_23288,N_23463);
and U23628 (N_23628,N_23349,N_23424);
or U23629 (N_23629,N_23464,N_23300);
or U23630 (N_23630,N_23303,N_23379);
nor U23631 (N_23631,N_23320,N_23394);
nor U23632 (N_23632,N_23433,N_23410);
xor U23633 (N_23633,N_23363,N_23389);
and U23634 (N_23634,N_23456,N_23252);
nor U23635 (N_23635,N_23280,N_23450);
or U23636 (N_23636,N_23306,N_23446);
and U23637 (N_23637,N_23486,N_23373);
nor U23638 (N_23638,N_23421,N_23431);
or U23639 (N_23639,N_23462,N_23413);
nor U23640 (N_23640,N_23261,N_23325);
and U23641 (N_23641,N_23345,N_23414);
xnor U23642 (N_23642,N_23370,N_23408);
or U23643 (N_23643,N_23451,N_23417);
or U23644 (N_23644,N_23414,N_23370);
or U23645 (N_23645,N_23280,N_23375);
xor U23646 (N_23646,N_23371,N_23268);
xnor U23647 (N_23647,N_23317,N_23408);
and U23648 (N_23648,N_23312,N_23429);
nand U23649 (N_23649,N_23421,N_23299);
nand U23650 (N_23650,N_23431,N_23360);
or U23651 (N_23651,N_23255,N_23408);
or U23652 (N_23652,N_23350,N_23311);
or U23653 (N_23653,N_23472,N_23293);
and U23654 (N_23654,N_23381,N_23450);
nor U23655 (N_23655,N_23420,N_23320);
and U23656 (N_23656,N_23463,N_23321);
or U23657 (N_23657,N_23398,N_23277);
and U23658 (N_23658,N_23266,N_23265);
or U23659 (N_23659,N_23405,N_23474);
nor U23660 (N_23660,N_23389,N_23342);
xor U23661 (N_23661,N_23280,N_23380);
nand U23662 (N_23662,N_23433,N_23253);
xnor U23663 (N_23663,N_23468,N_23320);
nor U23664 (N_23664,N_23366,N_23281);
or U23665 (N_23665,N_23367,N_23309);
nor U23666 (N_23666,N_23432,N_23282);
or U23667 (N_23667,N_23289,N_23280);
or U23668 (N_23668,N_23309,N_23311);
and U23669 (N_23669,N_23271,N_23326);
or U23670 (N_23670,N_23448,N_23359);
or U23671 (N_23671,N_23351,N_23390);
and U23672 (N_23672,N_23271,N_23253);
and U23673 (N_23673,N_23442,N_23295);
or U23674 (N_23674,N_23329,N_23366);
nand U23675 (N_23675,N_23294,N_23299);
nand U23676 (N_23676,N_23490,N_23269);
nor U23677 (N_23677,N_23299,N_23343);
or U23678 (N_23678,N_23498,N_23327);
and U23679 (N_23679,N_23497,N_23464);
nor U23680 (N_23680,N_23263,N_23320);
and U23681 (N_23681,N_23287,N_23487);
xor U23682 (N_23682,N_23396,N_23403);
and U23683 (N_23683,N_23253,N_23300);
and U23684 (N_23684,N_23426,N_23281);
or U23685 (N_23685,N_23393,N_23377);
or U23686 (N_23686,N_23471,N_23454);
and U23687 (N_23687,N_23279,N_23319);
nor U23688 (N_23688,N_23432,N_23307);
nor U23689 (N_23689,N_23300,N_23278);
nor U23690 (N_23690,N_23378,N_23478);
nor U23691 (N_23691,N_23407,N_23460);
nand U23692 (N_23692,N_23390,N_23360);
nor U23693 (N_23693,N_23374,N_23460);
nor U23694 (N_23694,N_23276,N_23394);
xnor U23695 (N_23695,N_23288,N_23480);
or U23696 (N_23696,N_23429,N_23406);
xor U23697 (N_23697,N_23491,N_23300);
xnor U23698 (N_23698,N_23365,N_23463);
and U23699 (N_23699,N_23251,N_23298);
nand U23700 (N_23700,N_23326,N_23300);
xor U23701 (N_23701,N_23445,N_23360);
nand U23702 (N_23702,N_23364,N_23269);
nand U23703 (N_23703,N_23435,N_23416);
and U23704 (N_23704,N_23491,N_23452);
or U23705 (N_23705,N_23388,N_23378);
nor U23706 (N_23706,N_23371,N_23466);
or U23707 (N_23707,N_23360,N_23259);
or U23708 (N_23708,N_23332,N_23340);
nand U23709 (N_23709,N_23446,N_23345);
or U23710 (N_23710,N_23468,N_23386);
xnor U23711 (N_23711,N_23474,N_23472);
and U23712 (N_23712,N_23294,N_23296);
and U23713 (N_23713,N_23377,N_23453);
nor U23714 (N_23714,N_23441,N_23464);
nand U23715 (N_23715,N_23445,N_23278);
nor U23716 (N_23716,N_23406,N_23343);
or U23717 (N_23717,N_23401,N_23314);
nand U23718 (N_23718,N_23346,N_23335);
and U23719 (N_23719,N_23400,N_23476);
xor U23720 (N_23720,N_23431,N_23462);
nand U23721 (N_23721,N_23335,N_23263);
and U23722 (N_23722,N_23381,N_23411);
nor U23723 (N_23723,N_23484,N_23454);
xnor U23724 (N_23724,N_23392,N_23299);
nand U23725 (N_23725,N_23376,N_23294);
and U23726 (N_23726,N_23347,N_23445);
nor U23727 (N_23727,N_23487,N_23357);
or U23728 (N_23728,N_23390,N_23486);
nor U23729 (N_23729,N_23376,N_23277);
and U23730 (N_23730,N_23471,N_23299);
and U23731 (N_23731,N_23383,N_23410);
nor U23732 (N_23732,N_23260,N_23379);
nor U23733 (N_23733,N_23482,N_23413);
nor U23734 (N_23734,N_23485,N_23349);
nand U23735 (N_23735,N_23443,N_23468);
or U23736 (N_23736,N_23329,N_23256);
nor U23737 (N_23737,N_23429,N_23493);
or U23738 (N_23738,N_23358,N_23488);
or U23739 (N_23739,N_23391,N_23283);
xnor U23740 (N_23740,N_23357,N_23334);
nor U23741 (N_23741,N_23419,N_23495);
nand U23742 (N_23742,N_23391,N_23312);
xnor U23743 (N_23743,N_23255,N_23456);
nand U23744 (N_23744,N_23274,N_23386);
nor U23745 (N_23745,N_23329,N_23269);
xor U23746 (N_23746,N_23315,N_23280);
xor U23747 (N_23747,N_23477,N_23381);
nor U23748 (N_23748,N_23336,N_23460);
xnor U23749 (N_23749,N_23435,N_23313);
or U23750 (N_23750,N_23585,N_23532);
xor U23751 (N_23751,N_23609,N_23633);
xnor U23752 (N_23752,N_23723,N_23626);
or U23753 (N_23753,N_23737,N_23652);
nand U23754 (N_23754,N_23548,N_23595);
nor U23755 (N_23755,N_23512,N_23549);
and U23756 (N_23756,N_23628,N_23598);
xor U23757 (N_23757,N_23565,N_23566);
or U23758 (N_23758,N_23550,N_23599);
and U23759 (N_23759,N_23584,N_23622);
or U23760 (N_23760,N_23644,N_23672);
and U23761 (N_23761,N_23574,N_23714);
nand U23762 (N_23762,N_23613,N_23625);
nand U23763 (N_23763,N_23665,N_23553);
xor U23764 (N_23764,N_23709,N_23591);
and U23765 (N_23765,N_23608,N_23510);
or U23766 (N_23766,N_23597,N_23736);
nand U23767 (N_23767,N_23729,N_23580);
nor U23768 (N_23768,N_23544,N_23513);
or U23769 (N_23769,N_23588,N_23743);
xnor U23770 (N_23770,N_23586,N_23635);
and U23771 (N_23771,N_23569,N_23690);
and U23772 (N_23772,N_23593,N_23698);
nand U23773 (N_23773,N_23692,N_23521);
or U23774 (N_23774,N_23528,N_23575);
and U23775 (N_23775,N_23707,N_23662);
nand U23776 (N_23776,N_23557,N_23686);
nand U23777 (N_23777,N_23687,N_23531);
xnor U23778 (N_23778,N_23541,N_23680);
or U23779 (N_23779,N_23722,N_23725);
or U23780 (N_23780,N_23660,N_23577);
xor U23781 (N_23781,N_23558,N_23651);
nand U23782 (N_23782,N_23711,N_23618);
xnor U23783 (N_23783,N_23708,N_23699);
nand U23784 (N_23784,N_23721,N_23715);
or U23785 (N_23785,N_23678,N_23562);
xor U23786 (N_23786,N_23675,N_23696);
nand U23787 (N_23787,N_23739,N_23555);
xnor U23788 (N_23788,N_23501,N_23610);
or U23789 (N_23789,N_23630,N_23554);
nand U23790 (N_23790,N_23646,N_23623);
nor U23791 (N_23791,N_23647,N_23694);
and U23792 (N_23792,N_23682,N_23502);
xor U23793 (N_23793,N_23620,N_23542);
or U23794 (N_23794,N_23604,N_23668);
or U23795 (N_23795,N_23650,N_23508);
or U23796 (N_23796,N_23522,N_23649);
or U23797 (N_23797,N_23543,N_23645);
nand U23798 (N_23798,N_23564,N_23602);
nor U23799 (N_23799,N_23615,N_23606);
nor U23800 (N_23800,N_23632,N_23648);
nand U23801 (N_23801,N_23621,N_23706);
nor U23802 (N_23802,N_23551,N_23570);
nor U23803 (N_23803,N_23735,N_23516);
and U23804 (N_23804,N_23518,N_23741);
xnor U23805 (N_23805,N_23547,N_23667);
or U23806 (N_23806,N_23624,N_23629);
nor U23807 (N_23807,N_23561,N_23563);
nand U23808 (N_23808,N_23744,N_23663);
nand U23809 (N_23809,N_23614,N_23713);
nor U23810 (N_23810,N_23681,N_23616);
and U23811 (N_23811,N_23504,N_23640);
nor U23812 (N_23812,N_23679,N_23530);
or U23813 (N_23813,N_23559,N_23573);
and U23814 (N_23814,N_23600,N_23677);
and U23815 (N_23815,N_23734,N_23517);
and U23816 (N_23816,N_23505,N_23590);
or U23817 (N_23817,N_23603,N_23703);
or U23818 (N_23818,N_23738,N_23740);
xor U23819 (N_23819,N_23742,N_23695);
and U23820 (N_23820,N_23693,N_23700);
and U23821 (N_23821,N_23654,N_23533);
and U23822 (N_23822,N_23611,N_23656);
xor U23823 (N_23823,N_23607,N_23534);
nand U23824 (N_23824,N_23581,N_23506);
nor U23825 (N_23825,N_23643,N_23655);
nor U23826 (N_23826,N_23592,N_23728);
nand U23827 (N_23827,N_23724,N_23638);
or U23828 (N_23828,N_23720,N_23529);
nor U23829 (N_23829,N_23568,N_23704);
and U23830 (N_23830,N_23636,N_23670);
nand U23831 (N_23831,N_23745,N_23579);
or U23832 (N_23832,N_23727,N_23748);
nor U23833 (N_23833,N_23674,N_23596);
or U23834 (N_23834,N_23671,N_23639);
nor U23835 (N_23835,N_23749,N_23688);
nor U23836 (N_23836,N_23526,N_23641);
and U23837 (N_23837,N_23691,N_23571);
xor U23838 (N_23838,N_23702,N_23537);
or U23839 (N_23839,N_23546,N_23732);
nand U23840 (N_23840,N_23627,N_23519);
nand U23841 (N_23841,N_23619,N_23589);
xnor U23842 (N_23842,N_23524,N_23684);
nand U23843 (N_23843,N_23523,N_23601);
xor U23844 (N_23844,N_23520,N_23500);
nor U23845 (N_23845,N_23637,N_23683);
nor U23846 (N_23846,N_23676,N_23669);
xor U23847 (N_23847,N_23661,N_23583);
or U23848 (N_23848,N_23572,N_23527);
nor U23849 (N_23849,N_23689,N_23747);
nor U23850 (N_23850,N_23718,N_23560);
xor U23851 (N_23851,N_23582,N_23605);
nor U23852 (N_23852,N_23716,N_23685);
nand U23853 (N_23853,N_23535,N_23664);
nor U23854 (N_23854,N_23507,N_23673);
nor U23855 (N_23855,N_23719,N_23659);
nor U23856 (N_23856,N_23701,N_23576);
or U23857 (N_23857,N_23514,N_23594);
nor U23858 (N_23858,N_23545,N_23705);
or U23859 (N_23859,N_23538,N_23634);
or U23860 (N_23860,N_23697,N_23511);
or U23861 (N_23861,N_23733,N_23525);
nand U23862 (N_23862,N_23631,N_23536);
xnor U23863 (N_23863,N_23617,N_23509);
nand U23864 (N_23864,N_23503,N_23552);
or U23865 (N_23865,N_23717,N_23657);
or U23866 (N_23866,N_23539,N_23556);
nand U23867 (N_23867,N_23726,N_23712);
nor U23868 (N_23868,N_23540,N_23658);
nor U23869 (N_23869,N_23666,N_23731);
nand U23870 (N_23870,N_23612,N_23730);
nand U23871 (N_23871,N_23515,N_23746);
nand U23872 (N_23872,N_23587,N_23710);
xnor U23873 (N_23873,N_23653,N_23642);
xor U23874 (N_23874,N_23578,N_23567);
nand U23875 (N_23875,N_23517,N_23741);
or U23876 (N_23876,N_23639,N_23705);
or U23877 (N_23877,N_23725,N_23693);
nor U23878 (N_23878,N_23675,N_23652);
or U23879 (N_23879,N_23710,N_23705);
or U23880 (N_23880,N_23558,N_23649);
xor U23881 (N_23881,N_23543,N_23646);
nand U23882 (N_23882,N_23598,N_23725);
nand U23883 (N_23883,N_23604,N_23629);
nand U23884 (N_23884,N_23749,N_23634);
xnor U23885 (N_23885,N_23615,N_23664);
or U23886 (N_23886,N_23716,N_23516);
xor U23887 (N_23887,N_23712,N_23650);
and U23888 (N_23888,N_23528,N_23709);
and U23889 (N_23889,N_23515,N_23523);
or U23890 (N_23890,N_23743,N_23606);
nand U23891 (N_23891,N_23647,N_23689);
nor U23892 (N_23892,N_23509,N_23605);
nor U23893 (N_23893,N_23506,N_23717);
nor U23894 (N_23894,N_23653,N_23587);
or U23895 (N_23895,N_23728,N_23533);
or U23896 (N_23896,N_23520,N_23590);
nand U23897 (N_23897,N_23742,N_23690);
nor U23898 (N_23898,N_23714,N_23579);
nand U23899 (N_23899,N_23739,N_23568);
nand U23900 (N_23900,N_23669,N_23690);
xnor U23901 (N_23901,N_23608,N_23691);
xnor U23902 (N_23902,N_23560,N_23743);
nand U23903 (N_23903,N_23645,N_23581);
or U23904 (N_23904,N_23732,N_23551);
nand U23905 (N_23905,N_23696,N_23503);
and U23906 (N_23906,N_23703,N_23556);
xnor U23907 (N_23907,N_23583,N_23655);
nand U23908 (N_23908,N_23699,N_23599);
xnor U23909 (N_23909,N_23521,N_23702);
and U23910 (N_23910,N_23627,N_23558);
and U23911 (N_23911,N_23649,N_23512);
nor U23912 (N_23912,N_23570,N_23522);
and U23913 (N_23913,N_23572,N_23649);
and U23914 (N_23914,N_23590,N_23689);
and U23915 (N_23915,N_23708,N_23698);
nand U23916 (N_23916,N_23708,N_23677);
xor U23917 (N_23917,N_23689,N_23547);
or U23918 (N_23918,N_23620,N_23587);
xnor U23919 (N_23919,N_23658,N_23537);
and U23920 (N_23920,N_23716,N_23618);
xor U23921 (N_23921,N_23655,N_23552);
or U23922 (N_23922,N_23606,N_23633);
nand U23923 (N_23923,N_23658,N_23657);
or U23924 (N_23924,N_23687,N_23649);
xnor U23925 (N_23925,N_23588,N_23534);
or U23926 (N_23926,N_23591,N_23668);
nor U23927 (N_23927,N_23571,N_23530);
and U23928 (N_23928,N_23564,N_23617);
xor U23929 (N_23929,N_23643,N_23520);
and U23930 (N_23930,N_23565,N_23655);
nand U23931 (N_23931,N_23608,N_23569);
nand U23932 (N_23932,N_23718,N_23613);
and U23933 (N_23933,N_23620,N_23681);
xor U23934 (N_23934,N_23508,N_23631);
nand U23935 (N_23935,N_23724,N_23513);
and U23936 (N_23936,N_23747,N_23615);
nand U23937 (N_23937,N_23649,N_23556);
xnor U23938 (N_23938,N_23500,N_23582);
nand U23939 (N_23939,N_23562,N_23512);
nor U23940 (N_23940,N_23569,N_23588);
and U23941 (N_23941,N_23617,N_23640);
xnor U23942 (N_23942,N_23603,N_23561);
or U23943 (N_23943,N_23540,N_23639);
and U23944 (N_23944,N_23594,N_23530);
nand U23945 (N_23945,N_23714,N_23515);
xnor U23946 (N_23946,N_23587,N_23616);
nor U23947 (N_23947,N_23719,N_23633);
xor U23948 (N_23948,N_23515,N_23504);
and U23949 (N_23949,N_23691,N_23749);
nand U23950 (N_23950,N_23504,N_23703);
xor U23951 (N_23951,N_23625,N_23707);
and U23952 (N_23952,N_23564,N_23655);
and U23953 (N_23953,N_23648,N_23560);
nor U23954 (N_23954,N_23703,N_23622);
xnor U23955 (N_23955,N_23587,N_23607);
and U23956 (N_23956,N_23736,N_23513);
nor U23957 (N_23957,N_23508,N_23656);
nand U23958 (N_23958,N_23569,N_23646);
xnor U23959 (N_23959,N_23623,N_23555);
nor U23960 (N_23960,N_23612,N_23698);
or U23961 (N_23961,N_23631,N_23550);
and U23962 (N_23962,N_23717,N_23515);
nor U23963 (N_23963,N_23632,N_23664);
and U23964 (N_23964,N_23674,N_23586);
xor U23965 (N_23965,N_23671,N_23627);
nor U23966 (N_23966,N_23685,N_23673);
nand U23967 (N_23967,N_23690,N_23734);
xor U23968 (N_23968,N_23703,N_23523);
nand U23969 (N_23969,N_23564,N_23517);
or U23970 (N_23970,N_23742,N_23623);
xor U23971 (N_23971,N_23582,N_23674);
nand U23972 (N_23972,N_23500,N_23646);
xnor U23973 (N_23973,N_23740,N_23571);
nor U23974 (N_23974,N_23720,N_23609);
xnor U23975 (N_23975,N_23645,N_23519);
and U23976 (N_23976,N_23740,N_23593);
and U23977 (N_23977,N_23536,N_23529);
nand U23978 (N_23978,N_23519,N_23690);
nand U23979 (N_23979,N_23579,N_23598);
and U23980 (N_23980,N_23738,N_23595);
nand U23981 (N_23981,N_23551,N_23703);
nand U23982 (N_23982,N_23526,N_23534);
and U23983 (N_23983,N_23656,N_23709);
xnor U23984 (N_23984,N_23564,N_23660);
nor U23985 (N_23985,N_23608,N_23686);
and U23986 (N_23986,N_23734,N_23623);
nor U23987 (N_23987,N_23516,N_23558);
nand U23988 (N_23988,N_23519,N_23674);
xor U23989 (N_23989,N_23543,N_23655);
and U23990 (N_23990,N_23532,N_23502);
and U23991 (N_23991,N_23523,N_23668);
and U23992 (N_23992,N_23705,N_23552);
nand U23993 (N_23993,N_23726,N_23562);
xnor U23994 (N_23994,N_23510,N_23743);
xnor U23995 (N_23995,N_23713,N_23730);
and U23996 (N_23996,N_23665,N_23747);
nand U23997 (N_23997,N_23607,N_23682);
xnor U23998 (N_23998,N_23714,N_23528);
xnor U23999 (N_23999,N_23547,N_23635);
nor U24000 (N_24000,N_23833,N_23815);
xor U24001 (N_24001,N_23884,N_23764);
or U24002 (N_24002,N_23806,N_23850);
xnor U24003 (N_24003,N_23978,N_23767);
nor U24004 (N_24004,N_23950,N_23779);
and U24005 (N_24005,N_23876,N_23887);
or U24006 (N_24006,N_23938,N_23894);
nor U24007 (N_24007,N_23924,N_23832);
and U24008 (N_24008,N_23939,N_23798);
nor U24009 (N_24009,N_23786,N_23760);
xor U24010 (N_24010,N_23891,N_23908);
nor U24011 (N_24011,N_23866,N_23947);
xor U24012 (N_24012,N_23948,N_23790);
nor U24013 (N_24013,N_23899,N_23890);
or U24014 (N_24014,N_23933,N_23913);
xnor U24015 (N_24015,N_23766,N_23919);
or U24016 (N_24016,N_23783,N_23882);
and U24017 (N_24017,N_23835,N_23991);
nor U24018 (N_24018,N_23784,N_23877);
or U24019 (N_24019,N_23812,N_23756);
nand U24020 (N_24020,N_23992,N_23911);
nand U24021 (N_24021,N_23980,N_23910);
nand U24022 (N_24022,N_23796,N_23925);
and U24023 (N_24023,N_23889,N_23984);
nor U24024 (N_24024,N_23903,N_23945);
xor U24025 (N_24025,N_23792,N_23974);
nor U24026 (N_24026,N_23958,N_23810);
and U24027 (N_24027,N_23907,N_23868);
and U24028 (N_24028,N_23937,N_23853);
and U24029 (N_24029,N_23966,N_23999);
nor U24030 (N_24030,N_23898,N_23780);
xor U24031 (N_24031,N_23915,N_23830);
nor U24032 (N_24032,N_23776,N_23820);
xnor U24033 (N_24033,N_23972,N_23967);
and U24034 (N_24034,N_23883,N_23785);
xor U24035 (N_24035,N_23775,N_23926);
or U24036 (N_24036,N_23782,N_23849);
nand U24037 (N_24037,N_23862,N_23989);
or U24038 (N_24038,N_23827,N_23920);
or U24039 (N_24039,N_23871,N_23879);
nand U24040 (N_24040,N_23901,N_23994);
nand U24041 (N_24041,N_23942,N_23755);
or U24042 (N_24042,N_23976,N_23927);
and U24043 (N_24043,N_23829,N_23804);
or U24044 (N_24044,N_23856,N_23874);
nand U24045 (N_24045,N_23841,N_23971);
or U24046 (N_24046,N_23988,N_23957);
and U24047 (N_24047,N_23824,N_23930);
nor U24048 (N_24048,N_23941,N_23761);
nor U24049 (N_24049,N_23765,N_23794);
nand U24050 (N_24050,N_23929,N_23808);
nand U24051 (N_24051,N_23961,N_23896);
and U24052 (N_24052,N_23912,N_23934);
nand U24053 (N_24053,N_23773,N_23970);
nand U24054 (N_24054,N_23855,N_23809);
nor U24055 (N_24055,N_23951,N_23789);
nand U24056 (N_24056,N_23818,N_23949);
or U24057 (N_24057,N_23787,N_23897);
and U24058 (N_24058,N_23923,N_23960);
xnor U24059 (N_24059,N_23778,N_23892);
nand U24060 (N_24060,N_23928,N_23763);
and U24061 (N_24061,N_23813,N_23895);
or U24062 (N_24062,N_23955,N_23921);
xor U24063 (N_24063,N_23822,N_23956);
nand U24064 (N_24064,N_23909,N_23881);
or U24065 (N_24065,N_23888,N_23837);
nor U24066 (N_24066,N_23793,N_23805);
xor U24067 (N_24067,N_23821,N_23772);
nor U24068 (N_24068,N_23838,N_23873);
and U24069 (N_24069,N_23834,N_23845);
nor U24070 (N_24070,N_23752,N_23878);
or U24071 (N_24071,N_23751,N_23981);
xnor U24072 (N_24072,N_23842,N_23854);
xnor U24073 (N_24073,N_23932,N_23823);
and U24074 (N_24074,N_23996,N_23817);
or U24075 (N_24075,N_23917,N_23825);
nand U24076 (N_24076,N_23916,N_23985);
nor U24077 (N_24077,N_23757,N_23803);
nor U24078 (N_24078,N_23982,N_23944);
nand U24079 (N_24079,N_23893,N_23847);
or U24080 (N_24080,N_23860,N_23900);
nand U24081 (N_24081,N_23997,N_23875);
nand U24082 (N_24082,N_23836,N_23931);
xor U24083 (N_24083,N_23762,N_23983);
nor U24084 (N_24084,N_23870,N_23774);
or U24085 (N_24085,N_23998,N_23859);
nand U24086 (N_24086,N_23819,N_23863);
nand U24087 (N_24087,N_23831,N_23811);
and U24088 (N_24088,N_23872,N_23979);
and U24089 (N_24089,N_23975,N_23946);
nor U24090 (N_24090,N_23777,N_23828);
or U24091 (N_24091,N_23839,N_23814);
or U24092 (N_24092,N_23840,N_23826);
nand U24093 (N_24093,N_23801,N_23987);
nand U24094 (N_24094,N_23906,N_23902);
nor U24095 (N_24095,N_23865,N_23962);
nand U24096 (N_24096,N_23965,N_23781);
or U24097 (N_24097,N_23952,N_23963);
nand U24098 (N_24098,N_23844,N_23990);
nor U24099 (N_24099,N_23986,N_23869);
nor U24100 (N_24100,N_23795,N_23807);
nor U24101 (N_24101,N_23769,N_23816);
nand U24102 (N_24102,N_23846,N_23753);
or U24103 (N_24103,N_23880,N_23768);
or U24104 (N_24104,N_23857,N_23918);
nand U24105 (N_24105,N_23867,N_23940);
or U24106 (N_24106,N_23964,N_23905);
xor U24107 (N_24107,N_23864,N_23968);
nand U24108 (N_24108,N_23969,N_23904);
or U24109 (N_24109,N_23758,N_23995);
or U24110 (N_24110,N_23943,N_23914);
and U24111 (N_24111,N_23959,N_23954);
xnor U24112 (N_24112,N_23799,N_23922);
or U24113 (N_24113,N_23843,N_23788);
and U24114 (N_24114,N_23885,N_23953);
and U24115 (N_24115,N_23770,N_23852);
nor U24116 (N_24116,N_23861,N_23848);
xor U24117 (N_24117,N_23977,N_23973);
nor U24118 (N_24118,N_23886,N_23800);
or U24119 (N_24119,N_23759,N_23802);
nand U24120 (N_24120,N_23797,N_23935);
nand U24121 (N_24121,N_23858,N_23936);
xnor U24122 (N_24122,N_23754,N_23771);
or U24123 (N_24123,N_23993,N_23791);
or U24124 (N_24124,N_23851,N_23750);
nand U24125 (N_24125,N_23896,N_23984);
nand U24126 (N_24126,N_23913,N_23765);
or U24127 (N_24127,N_23998,N_23933);
or U24128 (N_24128,N_23768,N_23826);
nand U24129 (N_24129,N_23998,N_23908);
xor U24130 (N_24130,N_23837,N_23842);
or U24131 (N_24131,N_23838,N_23864);
and U24132 (N_24132,N_23849,N_23851);
nor U24133 (N_24133,N_23851,N_23873);
xor U24134 (N_24134,N_23924,N_23939);
nor U24135 (N_24135,N_23804,N_23779);
nor U24136 (N_24136,N_23926,N_23822);
or U24137 (N_24137,N_23832,N_23857);
or U24138 (N_24138,N_23759,N_23818);
or U24139 (N_24139,N_23757,N_23829);
and U24140 (N_24140,N_23780,N_23851);
nor U24141 (N_24141,N_23793,N_23755);
nand U24142 (N_24142,N_23836,N_23922);
nand U24143 (N_24143,N_23939,N_23960);
nand U24144 (N_24144,N_23993,N_23819);
xor U24145 (N_24145,N_23794,N_23831);
and U24146 (N_24146,N_23779,N_23905);
or U24147 (N_24147,N_23938,N_23757);
and U24148 (N_24148,N_23762,N_23927);
xor U24149 (N_24149,N_23972,N_23759);
and U24150 (N_24150,N_23974,N_23772);
or U24151 (N_24151,N_23824,N_23981);
nor U24152 (N_24152,N_23867,N_23784);
or U24153 (N_24153,N_23899,N_23858);
nor U24154 (N_24154,N_23829,N_23855);
nor U24155 (N_24155,N_23811,N_23979);
xnor U24156 (N_24156,N_23792,N_23754);
or U24157 (N_24157,N_23781,N_23939);
and U24158 (N_24158,N_23766,N_23804);
xnor U24159 (N_24159,N_23828,N_23783);
and U24160 (N_24160,N_23814,N_23804);
xnor U24161 (N_24161,N_23946,N_23921);
and U24162 (N_24162,N_23816,N_23825);
nor U24163 (N_24163,N_23983,N_23823);
nor U24164 (N_24164,N_23972,N_23977);
xnor U24165 (N_24165,N_23841,N_23886);
xor U24166 (N_24166,N_23791,N_23883);
nand U24167 (N_24167,N_23832,N_23777);
and U24168 (N_24168,N_23991,N_23754);
and U24169 (N_24169,N_23794,N_23851);
nor U24170 (N_24170,N_23845,N_23994);
xnor U24171 (N_24171,N_23812,N_23893);
nor U24172 (N_24172,N_23757,N_23764);
xnor U24173 (N_24173,N_23788,N_23971);
xnor U24174 (N_24174,N_23890,N_23902);
xnor U24175 (N_24175,N_23906,N_23753);
xnor U24176 (N_24176,N_23882,N_23942);
xor U24177 (N_24177,N_23825,N_23924);
or U24178 (N_24178,N_23927,N_23899);
and U24179 (N_24179,N_23790,N_23870);
nand U24180 (N_24180,N_23918,N_23813);
and U24181 (N_24181,N_23820,N_23824);
or U24182 (N_24182,N_23951,N_23980);
or U24183 (N_24183,N_23807,N_23963);
nor U24184 (N_24184,N_23871,N_23973);
and U24185 (N_24185,N_23828,N_23935);
or U24186 (N_24186,N_23832,N_23905);
nor U24187 (N_24187,N_23987,N_23998);
or U24188 (N_24188,N_23832,N_23752);
nand U24189 (N_24189,N_23916,N_23864);
nor U24190 (N_24190,N_23767,N_23969);
or U24191 (N_24191,N_23856,N_23772);
nor U24192 (N_24192,N_23851,N_23988);
or U24193 (N_24193,N_23857,N_23896);
xnor U24194 (N_24194,N_23754,N_23831);
xnor U24195 (N_24195,N_23939,N_23870);
or U24196 (N_24196,N_23991,N_23827);
xnor U24197 (N_24197,N_23848,N_23967);
nand U24198 (N_24198,N_23967,N_23789);
or U24199 (N_24199,N_23932,N_23812);
nand U24200 (N_24200,N_23840,N_23919);
and U24201 (N_24201,N_23951,N_23891);
nor U24202 (N_24202,N_23817,N_23889);
nor U24203 (N_24203,N_23879,N_23884);
nor U24204 (N_24204,N_23799,N_23943);
xor U24205 (N_24205,N_23899,N_23885);
nand U24206 (N_24206,N_23832,N_23875);
xor U24207 (N_24207,N_23972,N_23940);
xnor U24208 (N_24208,N_23862,N_23891);
xnor U24209 (N_24209,N_23796,N_23969);
nand U24210 (N_24210,N_23986,N_23896);
and U24211 (N_24211,N_23941,N_23936);
xnor U24212 (N_24212,N_23799,N_23992);
nor U24213 (N_24213,N_23880,N_23849);
xnor U24214 (N_24214,N_23951,N_23858);
and U24215 (N_24215,N_23912,N_23939);
nand U24216 (N_24216,N_23914,N_23862);
xor U24217 (N_24217,N_23770,N_23906);
or U24218 (N_24218,N_23930,N_23871);
xnor U24219 (N_24219,N_23796,N_23887);
or U24220 (N_24220,N_23901,N_23885);
or U24221 (N_24221,N_23989,N_23798);
or U24222 (N_24222,N_23886,N_23758);
nor U24223 (N_24223,N_23960,N_23777);
and U24224 (N_24224,N_23970,N_23813);
nand U24225 (N_24225,N_23840,N_23920);
or U24226 (N_24226,N_23997,N_23947);
nand U24227 (N_24227,N_23945,N_23755);
nor U24228 (N_24228,N_23953,N_23990);
nand U24229 (N_24229,N_23873,N_23911);
or U24230 (N_24230,N_23808,N_23943);
and U24231 (N_24231,N_23840,N_23781);
nor U24232 (N_24232,N_23812,N_23834);
and U24233 (N_24233,N_23993,N_23793);
nor U24234 (N_24234,N_23842,N_23883);
nand U24235 (N_24235,N_23836,N_23981);
and U24236 (N_24236,N_23926,N_23796);
nor U24237 (N_24237,N_23893,N_23957);
nor U24238 (N_24238,N_23909,N_23840);
xnor U24239 (N_24239,N_23885,N_23775);
nor U24240 (N_24240,N_23926,N_23897);
nand U24241 (N_24241,N_23936,N_23995);
or U24242 (N_24242,N_23797,N_23819);
nand U24243 (N_24243,N_23845,N_23952);
xnor U24244 (N_24244,N_23780,N_23845);
nand U24245 (N_24245,N_23939,N_23755);
nor U24246 (N_24246,N_23762,N_23873);
and U24247 (N_24247,N_23867,N_23856);
nor U24248 (N_24248,N_23897,N_23904);
nand U24249 (N_24249,N_23884,N_23799);
xor U24250 (N_24250,N_24089,N_24087);
or U24251 (N_24251,N_24060,N_24152);
or U24252 (N_24252,N_24107,N_24239);
and U24253 (N_24253,N_24048,N_24074);
and U24254 (N_24254,N_24176,N_24177);
xnor U24255 (N_24255,N_24154,N_24221);
nand U24256 (N_24256,N_24077,N_24041);
nand U24257 (N_24257,N_24012,N_24081);
and U24258 (N_24258,N_24114,N_24182);
nand U24259 (N_24259,N_24170,N_24139);
nand U24260 (N_24260,N_24101,N_24019);
or U24261 (N_24261,N_24135,N_24179);
xor U24262 (N_24262,N_24066,N_24210);
nor U24263 (N_24263,N_24005,N_24134);
nand U24264 (N_24264,N_24249,N_24016);
nor U24265 (N_24265,N_24023,N_24213);
xor U24266 (N_24266,N_24008,N_24193);
and U24267 (N_24267,N_24243,N_24034);
xnor U24268 (N_24268,N_24248,N_24116);
xnor U24269 (N_24269,N_24209,N_24158);
nand U24270 (N_24270,N_24088,N_24211);
nor U24271 (N_24271,N_24229,N_24136);
or U24272 (N_24272,N_24159,N_24125);
xor U24273 (N_24273,N_24173,N_24190);
nand U24274 (N_24274,N_24029,N_24062);
and U24275 (N_24275,N_24076,N_24133);
nand U24276 (N_24276,N_24175,N_24061);
nand U24277 (N_24277,N_24043,N_24006);
nand U24278 (N_24278,N_24108,N_24242);
and U24279 (N_24279,N_24137,N_24247);
xor U24280 (N_24280,N_24132,N_24090);
xnor U24281 (N_24281,N_24241,N_24155);
or U24282 (N_24282,N_24082,N_24053);
xor U24283 (N_24283,N_24145,N_24014);
nand U24284 (N_24284,N_24004,N_24122);
nand U24285 (N_24285,N_24223,N_24202);
nand U24286 (N_24286,N_24162,N_24143);
xor U24287 (N_24287,N_24028,N_24102);
nand U24288 (N_24288,N_24010,N_24009);
nor U24289 (N_24289,N_24057,N_24113);
or U24290 (N_24290,N_24174,N_24044);
xor U24291 (N_24291,N_24217,N_24218);
or U24292 (N_24292,N_24171,N_24039);
xor U24293 (N_24293,N_24085,N_24083);
nand U24294 (N_24294,N_24104,N_24149);
nor U24295 (N_24295,N_24224,N_24234);
xnor U24296 (N_24296,N_24047,N_24126);
nor U24297 (N_24297,N_24235,N_24075);
xor U24298 (N_24298,N_24055,N_24232);
or U24299 (N_24299,N_24021,N_24205);
xnor U24300 (N_24300,N_24119,N_24115);
or U24301 (N_24301,N_24141,N_24204);
nand U24302 (N_24302,N_24203,N_24178);
and U24303 (N_24303,N_24227,N_24110);
and U24304 (N_24304,N_24096,N_24127);
xnor U24305 (N_24305,N_24112,N_24185);
nand U24306 (N_24306,N_24166,N_24165);
nand U24307 (N_24307,N_24036,N_24191);
nand U24308 (N_24308,N_24094,N_24022);
nand U24309 (N_24309,N_24184,N_24098);
nor U24310 (N_24310,N_24040,N_24188);
or U24311 (N_24311,N_24065,N_24002);
xor U24312 (N_24312,N_24198,N_24109);
nand U24313 (N_24313,N_24111,N_24099);
and U24314 (N_24314,N_24238,N_24097);
nand U24315 (N_24315,N_24045,N_24032);
xor U24316 (N_24316,N_24201,N_24144);
nand U24317 (N_24317,N_24206,N_24194);
nand U24318 (N_24318,N_24037,N_24128);
and U24319 (N_24319,N_24138,N_24220);
nand U24320 (N_24320,N_24146,N_24054);
or U24321 (N_24321,N_24068,N_24013);
xnor U24322 (N_24322,N_24049,N_24046);
or U24323 (N_24323,N_24142,N_24042);
nand U24324 (N_24324,N_24216,N_24086);
or U24325 (N_24325,N_24195,N_24180);
and U24326 (N_24326,N_24100,N_24000);
nor U24327 (N_24327,N_24093,N_24233);
nand U24328 (N_24328,N_24157,N_24091);
nor U24329 (N_24329,N_24129,N_24192);
and U24330 (N_24330,N_24199,N_24237);
and U24331 (N_24331,N_24078,N_24120);
or U24332 (N_24332,N_24130,N_24052);
nor U24333 (N_24333,N_24030,N_24225);
xnor U24334 (N_24334,N_24181,N_24072);
nand U24335 (N_24335,N_24236,N_24214);
xor U24336 (N_24336,N_24219,N_24151);
nor U24337 (N_24337,N_24208,N_24080);
xnor U24338 (N_24338,N_24033,N_24092);
and U24339 (N_24339,N_24200,N_24073);
and U24340 (N_24340,N_24105,N_24067);
and U24341 (N_24341,N_24160,N_24161);
and U24342 (N_24342,N_24035,N_24147);
nand U24343 (N_24343,N_24189,N_24207);
nand U24344 (N_24344,N_24063,N_24071);
nand U24345 (N_24345,N_24024,N_24124);
or U24346 (N_24346,N_24168,N_24018);
nand U24347 (N_24347,N_24003,N_24079);
and U24348 (N_24348,N_24020,N_24197);
and U24349 (N_24349,N_24027,N_24103);
and U24350 (N_24350,N_24051,N_24026);
nand U24351 (N_24351,N_24050,N_24007);
nor U24352 (N_24352,N_24069,N_24187);
xnor U24353 (N_24353,N_24017,N_24163);
and U24354 (N_24354,N_24172,N_24215);
xor U24355 (N_24355,N_24059,N_24231);
xor U24356 (N_24356,N_24245,N_24196);
nor U24357 (N_24357,N_24058,N_24153);
nand U24358 (N_24358,N_24240,N_24031);
nand U24359 (N_24359,N_24156,N_24212);
nor U24360 (N_24360,N_24228,N_24246);
nor U24361 (N_24361,N_24011,N_24222);
nor U24362 (N_24362,N_24084,N_24117);
nand U24363 (N_24363,N_24015,N_24150);
or U24364 (N_24364,N_24001,N_24164);
and U24365 (N_24365,N_24106,N_24056);
nand U24366 (N_24366,N_24169,N_24167);
nor U24367 (N_24367,N_24070,N_24025);
or U24368 (N_24368,N_24118,N_24226);
nor U24369 (N_24369,N_24038,N_24140);
xor U24370 (N_24370,N_24186,N_24244);
xor U24371 (N_24371,N_24131,N_24230);
and U24372 (N_24372,N_24123,N_24121);
and U24373 (N_24373,N_24064,N_24095);
nor U24374 (N_24374,N_24148,N_24183);
nor U24375 (N_24375,N_24110,N_24228);
nand U24376 (N_24376,N_24048,N_24237);
or U24377 (N_24377,N_24218,N_24097);
and U24378 (N_24378,N_24201,N_24118);
nand U24379 (N_24379,N_24005,N_24054);
nand U24380 (N_24380,N_24025,N_24227);
xnor U24381 (N_24381,N_24022,N_24101);
or U24382 (N_24382,N_24148,N_24007);
and U24383 (N_24383,N_24175,N_24039);
nand U24384 (N_24384,N_24036,N_24022);
and U24385 (N_24385,N_24009,N_24142);
nand U24386 (N_24386,N_24214,N_24137);
nor U24387 (N_24387,N_24172,N_24051);
and U24388 (N_24388,N_24012,N_24171);
nor U24389 (N_24389,N_24234,N_24117);
or U24390 (N_24390,N_24240,N_24075);
and U24391 (N_24391,N_24151,N_24239);
or U24392 (N_24392,N_24005,N_24239);
nor U24393 (N_24393,N_24081,N_24067);
nand U24394 (N_24394,N_24086,N_24124);
and U24395 (N_24395,N_24150,N_24070);
xor U24396 (N_24396,N_24016,N_24186);
and U24397 (N_24397,N_24219,N_24010);
and U24398 (N_24398,N_24178,N_24072);
nand U24399 (N_24399,N_24153,N_24009);
and U24400 (N_24400,N_24231,N_24195);
and U24401 (N_24401,N_24083,N_24247);
nor U24402 (N_24402,N_24113,N_24181);
xor U24403 (N_24403,N_24097,N_24223);
xnor U24404 (N_24404,N_24001,N_24195);
nor U24405 (N_24405,N_24036,N_24117);
nor U24406 (N_24406,N_24010,N_24066);
xor U24407 (N_24407,N_24122,N_24006);
and U24408 (N_24408,N_24180,N_24125);
xor U24409 (N_24409,N_24135,N_24111);
nand U24410 (N_24410,N_24104,N_24205);
nand U24411 (N_24411,N_24227,N_24028);
and U24412 (N_24412,N_24244,N_24191);
xnor U24413 (N_24413,N_24077,N_24119);
xnor U24414 (N_24414,N_24005,N_24188);
or U24415 (N_24415,N_24187,N_24144);
and U24416 (N_24416,N_24055,N_24249);
nand U24417 (N_24417,N_24127,N_24103);
xnor U24418 (N_24418,N_24141,N_24198);
xnor U24419 (N_24419,N_24248,N_24200);
nand U24420 (N_24420,N_24232,N_24207);
xnor U24421 (N_24421,N_24216,N_24044);
nor U24422 (N_24422,N_24228,N_24094);
nand U24423 (N_24423,N_24202,N_24142);
xor U24424 (N_24424,N_24174,N_24007);
or U24425 (N_24425,N_24240,N_24057);
nor U24426 (N_24426,N_24082,N_24131);
nand U24427 (N_24427,N_24176,N_24060);
xnor U24428 (N_24428,N_24025,N_24249);
or U24429 (N_24429,N_24021,N_24009);
and U24430 (N_24430,N_24068,N_24137);
or U24431 (N_24431,N_24174,N_24082);
and U24432 (N_24432,N_24249,N_24201);
and U24433 (N_24433,N_24044,N_24102);
and U24434 (N_24434,N_24163,N_24020);
or U24435 (N_24435,N_24097,N_24121);
nor U24436 (N_24436,N_24125,N_24181);
or U24437 (N_24437,N_24172,N_24060);
and U24438 (N_24438,N_24141,N_24245);
nor U24439 (N_24439,N_24057,N_24218);
nor U24440 (N_24440,N_24105,N_24050);
xor U24441 (N_24441,N_24008,N_24189);
and U24442 (N_24442,N_24223,N_24046);
xor U24443 (N_24443,N_24112,N_24219);
nand U24444 (N_24444,N_24031,N_24129);
or U24445 (N_24445,N_24175,N_24167);
and U24446 (N_24446,N_24233,N_24089);
nand U24447 (N_24447,N_24201,N_24131);
and U24448 (N_24448,N_24037,N_24023);
and U24449 (N_24449,N_24231,N_24171);
nand U24450 (N_24450,N_24049,N_24022);
nor U24451 (N_24451,N_24103,N_24160);
or U24452 (N_24452,N_24098,N_24018);
nand U24453 (N_24453,N_24234,N_24067);
nand U24454 (N_24454,N_24245,N_24027);
xnor U24455 (N_24455,N_24108,N_24015);
xor U24456 (N_24456,N_24115,N_24174);
or U24457 (N_24457,N_24139,N_24244);
nand U24458 (N_24458,N_24105,N_24182);
nand U24459 (N_24459,N_24167,N_24058);
and U24460 (N_24460,N_24241,N_24049);
and U24461 (N_24461,N_24201,N_24062);
nor U24462 (N_24462,N_24196,N_24046);
nand U24463 (N_24463,N_24204,N_24110);
nand U24464 (N_24464,N_24060,N_24147);
nand U24465 (N_24465,N_24148,N_24038);
xnor U24466 (N_24466,N_24135,N_24071);
nor U24467 (N_24467,N_24221,N_24204);
nand U24468 (N_24468,N_24079,N_24103);
or U24469 (N_24469,N_24167,N_24049);
nor U24470 (N_24470,N_24117,N_24155);
nand U24471 (N_24471,N_24112,N_24242);
nor U24472 (N_24472,N_24229,N_24108);
xnor U24473 (N_24473,N_24001,N_24068);
nand U24474 (N_24474,N_24178,N_24207);
and U24475 (N_24475,N_24126,N_24145);
nor U24476 (N_24476,N_24133,N_24134);
nand U24477 (N_24477,N_24105,N_24083);
nor U24478 (N_24478,N_24216,N_24184);
and U24479 (N_24479,N_24010,N_24006);
nor U24480 (N_24480,N_24049,N_24140);
and U24481 (N_24481,N_24189,N_24230);
nor U24482 (N_24482,N_24129,N_24138);
xnor U24483 (N_24483,N_24080,N_24013);
and U24484 (N_24484,N_24244,N_24243);
nor U24485 (N_24485,N_24136,N_24216);
nand U24486 (N_24486,N_24147,N_24144);
nor U24487 (N_24487,N_24075,N_24041);
nor U24488 (N_24488,N_24000,N_24178);
xor U24489 (N_24489,N_24094,N_24210);
or U24490 (N_24490,N_24140,N_24108);
nor U24491 (N_24491,N_24132,N_24135);
nand U24492 (N_24492,N_24225,N_24163);
nand U24493 (N_24493,N_24091,N_24176);
nand U24494 (N_24494,N_24051,N_24236);
nor U24495 (N_24495,N_24079,N_24217);
or U24496 (N_24496,N_24210,N_24143);
nand U24497 (N_24497,N_24022,N_24070);
nand U24498 (N_24498,N_24097,N_24098);
and U24499 (N_24499,N_24119,N_24054);
nor U24500 (N_24500,N_24385,N_24375);
or U24501 (N_24501,N_24289,N_24275);
nand U24502 (N_24502,N_24259,N_24312);
and U24503 (N_24503,N_24408,N_24478);
or U24504 (N_24504,N_24378,N_24483);
nor U24505 (N_24505,N_24474,N_24480);
and U24506 (N_24506,N_24469,N_24357);
xnor U24507 (N_24507,N_24351,N_24436);
nand U24508 (N_24508,N_24439,N_24290);
nor U24509 (N_24509,N_24489,N_24303);
or U24510 (N_24510,N_24374,N_24368);
or U24511 (N_24511,N_24499,N_24420);
nor U24512 (N_24512,N_24302,N_24257);
nor U24513 (N_24513,N_24421,N_24267);
xnor U24514 (N_24514,N_24459,N_24497);
or U24515 (N_24515,N_24423,N_24426);
nand U24516 (N_24516,N_24330,N_24438);
and U24517 (N_24517,N_24355,N_24435);
xnor U24518 (N_24518,N_24376,N_24437);
or U24519 (N_24519,N_24422,N_24444);
or U24520 (N_24520,N_24308,N_24453);
nor U24521 (N_24521,N_24442,N_24466);
nand U24522 (N_24522,N_24398,N_24293);
nor U24523 (N_24523,N_24406,N_24338);
nor U24524 (N_24524,N_24320,N_24460);
xnor U24525 (N_24525,N_24428,N_24292);
xnor U24526 (N_24526,N_24284,N_24416);
or U24527 (N_24527,N_24458,N_24317);
nor U24528 (N_24528,N_24325,N_24265);
or U24529 (N_24529,N_24481,N_24365);
nand U24530 (N_24530,N_24286,N_24433);
xor U24531 (N_24531,N_24496,N_24467);
or U24532 (N_24532,N_24276,N_24382);
or U24533 (N_24533,N_24470,N_24482);
nor U24534 (N_24534,N_24269,N_24372);
nor U24535 (N_24535,N_24395,N_24277);
xnor U24536 (N_24536,N_24305,N_24379);
xnor U24537 (N_24537,N_24354,N_24464);
nand U24538 (N_24538,N_24498,N_24394);
and U24539 (N_24539,N_24457,N_24323);
nand U24540 (N_24540,N_24488,N_24414);
xor U24541 (N_24541,N_24283,N_24333);
nand U24542 (N_24542,N_24287,N_24404);
and U24543 (N_24543,N_24484,N_24451);
nand U24544 (N_24544,N_24253,N_24328);
and U24545 (N_24545,N_24407,N_24358);
nand U24546 (N_24546,N_24295,N_24494);
nand U24547 (N_24547,N_24285,N_24367);
or U24548 (N_24548,N_24476,N_24341);
nor U24549 (N_24549,N_24359,N_24452);
nor U24550 (N_24550,N_24279,N_24311);
xor U24551 (N_24551,N_24288,N_24411);
xor U24552 (N_24552,N_24324,N_24319);
nand U24553 (N_24553,N_24380,N_24373);
or U24554 (N_24554,N_24432,N_24310);
xnor U24555 (N_24555,N_24396,N_24282);
nand U24556 (N_24556,N_24335,N_24252);
or U24557 (N_24557,N_24419,N_24493);
nand U24558 (N_24558,N_24261,N_24346);
and U24559 (N_24559,N_24350,N_24321);
nor U24560 (N_24560,N_24393,N_24402);
nor U24561 (N_24561,N_24315,N_24255);
xor U24562 (N_24562,N_24430,N_24445);
or U24563 (N_24563,N_24486,N_24446);
nand U24564 (N_24564,N_24399,N_24281);
xor U24565 (N_24565,N_24258,N_24417);
nand U24566 (N_24566,N_24434,N_24322);
xnor U24567 (N_24567,N_24316,N_24272);
or U24568 (N_24568,N_24254,N_24441);
and U24569 (N_24569,N_24266,N_24424);
and U24570 (N_24570,N_24371,N_24291);
nand U24571 (N_24571,N_24400,N_24256);
or U24572 (N_24572,N_24490,N_24440);
or U24573 (N_24573,N_24260,N_24413);
xor U24574 (N_24574,N_24301,N_24431);
nor U24575 (N_24575,N_24278,N_24262);
nor U24576 (N_24576,N_24427,N_24381);
and U24577 (N_24577,N_24314,N_24270);
nor U24578 (N_24578,N_24298,N_24369);
xnor U24579 (N_24579,N_24251,N_24472);
xnor U24580 (N_24580,N_24449,N_24479);
nand U24581 (N_24581,N_24273,N_24492);
nor U24582 (N_24582,N_24454,N_24384);
nand U24583 (N_24583,N_24342,N_24462);
nor U24584 (N_24584,N_24448,N_24300);
and U24585 (N_24585,N_24391,N_24347);
nand U24586 (N_24586,N_24401,N_24343);
or U24587 (N_24587,N_24429,N_24306);
and U24588 (N_24588,N_24487,N_24264);
and U24589 (N_24589,N_24304,N_24463);
and U24590 (N_24590,N_24471,N_24477);
or U24591 (N_24591,N_24461,N_24331);
and U24592 (N_24592,N_24409,N_24336);
xor U24593 (N_24593,N_24250,N_24309);
xnor U24594 (N_24594,N_24294,N_24405);
xor U24595 (N_24595,N_24268,N_24360);
nor U24596 (N_24596,N_24362,N_24352);
or U24597 (N_24597,N_24473,N_24299);
nor U24598 (N_24598,N_24339,N_24415);
or U24599 (N_24599,N_24491,N_24364);
and U24600 (N_24600,N_24389,N_24318);
nor U24601 (N_24601,N_24329,N_24274);
or U24602 (N_24602,N_24397,N_24386);
xor U24603 (N_24603,N_24332,N_24307);
or U24604 (N_24604,N_24370,N_24296);
nand U24605 (N_24605,N_24412,N_24377);
nand U24606 (N_24606,N_24447,N_24361);
xnor U24607 (N_24607,N_24313,N_24465);
and U24608 (N_24608,N_24334,N_24337);
nand U24609 (N_24609,N_24455,N_24387);
and U24610 (N_24610,N_24340,N_24356);
nor U24611 (N_24611,N_24349,N_24403);
nand U24612 (N_24612,N_24443,N_24297);
and U24613 (N_24613,N_24485,N_24450);
xnor U24614 (N_24614,N_24363,N_24366);
or U24615 (N_24615,N_24263,N_24353);
nor U24616 (N_24616,N_24425,N_24344);
nor U24617 (N_24617,N_24388,N_24418);
and U24618 (N_24618,N_24495,N_24383);
nand U24619 (N_24619,N_24348,N_24468);
and U24620 (N_24620,N_24280,N_24326);
nor U24621 (N_24621,N_24327,N_24271);
and U24622 (N_24622,N_24475,N_24392);
or U24623 (N_24623,N_24345,N_24456);
nand U24624 (N_24624,N_24410,N_24390);
xor U24625 (N_24625,N_24408,N_24440);
or U24626 (N_24626,N_24427,N_24320);
xnor U24627 (N_24627,N_24379,N_24410);
xor U24628 (N_24628,N_24465,N_24481);
and U24629 (N_24629,N_24367,N_24312);
and U24630 (N_24630,N_24406,N_24396);
and U24631 (N_24631,N_24402,N_24258);
xor U24632 (N_24632,N_24354,N_24413);
and U24633 (N_24633,N_24383,N_24376);
nand U24634 (N_24634,N_24330,N_24467);
and U24635 (N_24635,N_24252,N_24299);
xor U24636 (N_24636,N_24254,N_24379);
nor U24637 (N_24637,N_24423,N_24294);
xnor U24638 (N_24638,N_24279,N_24260);
nand U24639 (N_24639,N_24309,N_24359);
xnor U24640 (N_24640,N_24480,N_24449);
and U24641 (N_24641,N_24486,N_24267);
or U24642 (N_24642,N_24418,N_24386);
xnor U24643 (N_24643,N_24395,N_24473);
nor U24644 (N_24644,N_24374,N_24456);
nand U24645 (N_24645,N_24297,N_24419);
and U24646 (N_24646,N_24393,N_24380);
and U24647 (N_24647,N_24288,N_24318);
xnor U24648 (N_24648,N_24385,N_24331);
or U24649 (N_24649,N_24366,N_24402);
nor U24650 (N_24650,N_24384,N_24282);
or U24651 (N_24651,N_24378,N_24498);
nand U24652 (N_24652,N_24293,N_24259);
nor U24653 (N_24653,N_24406,N_24263);
nand U24654 (N_24654,N_24321,N_24329);
nor U24655 (N_24655,N_24415,N_24418);
and U24656 (N_24656,N_24347,N_24253);
or U24657 (N_24657,N_24277,N_24398);
nand U24658 (N_24658,N_24468,N_24291);
or U24659 (N_24659,N_24428,N_24387);
nor U24660 (N_24660,N_24399,N_24303);
or U24661 (N_24661,N_24379,N_24279);
nor U24662 (N_24662,N_24303,N_24461);
nand U24663 (N_24663,N_24258,N_24490);
xnor U24664 (N_24664,N_24267,N_24401);
xnor U24665 (N_24665,N_24358,N_24267);
nand U24666 (N_24666,N_24282,N_24441);
and U24667 (N_24667,N_24301,N_24377);
nand U24668 (N_24668,N_24437,N_24431);
and U24669 (N_24669,N_24289,N_24329);
xor U24670 (N_24670,N_24359,N_24495);
nand U24671 (N_24671,N_24381,N_24469);
nor U24672 (N_24672,N_24497,N_24384);
or U24673 (N_24673,N_24479,N_24332);
and U24674 (N_24674,N_24492,N_24499);
and U24675 (N_24675,N_24303,N_24368);
or U24676 (N_24676,N_24359,N_24270);
nand U24677 (N_24677,N_24418,N_24444);
and U24678 (N_24678,N_24252,N_24444);
or U24679 (N_24679,N_24307,N_24250);
and U24680 (N_24680,N_24394,N_24362);
or U24681 (N_24681,N_24438,N_24338);
xor U24682 (N_24682,N_24379,N_24354);
or U24683 (N_24683,N_24475,N_24333);
or U24684 (N_24684,N_24253,N_24276);
xnor U24685 (N_24685,N_24436,N_24407);
xnor U24686 (N_24686,N_24306,N_24273);
nor U24687 (N_24687,N_24363,N_24488);
and U24688 (N_24688,N_24328,N_24272);
xor U24689 (N_24689,N_24407,N_24396);
and U24690 (N_24690,N_24486,N_24285);
or U24691 (N_24691,N_24343,N_24484);
nand U24692 (N_24692,N_24465,N_24417);
nand U24693 (N_24693,N_24485,N_24495);
and U24694 (N_24694,N_24256,N_24430);
nand U24695 (N_24695,N_24397,N_24497);
or U24696 (N_24696,N_24315,N_24338);
xnor U24697 (N_24697,N_24350,N_24366);
xnor U24698 (N_24698,N_24408,N_24272);
xor U24699 (N_24699,N_24322,N_24285);
or U24700 (N_24700,N_24496,N_24353);
xnor U24701 (N_24701,N_24465,N_24397);
nor U24702 (N_24702,N_24399,N_24473);
or U24703 (N_24703,N_24367,N_24314);
xor U24704 (N_24704,N_24455,N_24263);
nor U24705 (N_24705,N_24340,N_24282);
or U24706 (N_24706,N_24331,N_24458);
and U24707 (N_24707,N_24399,N_24374);
or U24708 (N_24708,N_24427,N_24274);
nand U24709 (N_24709,N_24488,N_24471);
or U24710 (N_24710,N_24466,N_24417);
nand U24711 (N_24711,N_24354,N_24393);
or U24712 (N_24712,N_24495,N_24302);
and U24713 (N_24713,N_24441,N_24277);
and U24714 (N_24714,N_24491,N_24349);
nor U24715 (N_24715,N_24304,N_24318);
xor U24716 (N_24716,N_24413,N_24352);
or U24717 (N_24717,N_24402,N_24302);
and U24718 (N_24718,N_24448,N_24311);
and U24719 (N_24719,N_24293,N_24278);
xnor U24720 (N_24720,N_24345,N_24297);
xor U24721 (N_24721,N_24304,N_24392);
or U24722 (N_24722,N_24384,N_24319);
nor U24723 (N_24723,N_24488,N_24334);
and U24724 (N_24724,N_24424,N_24331);
nor U24725 (N_24725,N_24462,N_24473);
or U24726 (N_24726,N_24384,N_24299);
or U24727 (N_24727,N_24311,N_24294);
xor U24728 (N_24728,N_24442,N_24355);
and U24729 (N_24729,N_24273,N_24329);
nand U24730 (N_24730,N_24328,N_24284);
and U24731 (N_24731,N_24389,N_24287);
and U24732 (N_24732,N_24365,N_24455);
and U24733 (N_24733,N_24251,N_24354);
nor U24734 (N_24734,N_24316,N_24317);
nand U24735 (N_24735,N_24343,N_24409);
and U24736 (N_24736,N_24359,N_24290);
or U24737 (N_24737,N_24268,N_24333);
or U24738 (N_24738,N_24270,N_24468);
and U24739 (N_24739,N_24349,N_24424);
xor U24740 (N_24740,N_24256,N_24355);
or U24741 (N_24741,N_24252,N_24348);
nand U24742 (N_24742,N_24378,N_24313);
or U24743 (N_24743,N_24430,N_24401);
nand U24744 (N_24744,N_24409,N_24433);
or U24745 (N_24745,N_24462,N_24299);
or U24746 (N_24746,N_24419,N_24250);
or U24747 (N_24747,N_24290,N_24422);
xor U24748 (N_24748,N_24337,N_24256);
nand U24749 (N_24749,N_24351,N_24285);
xor U24750 (N_24750,N_24527,N_24725);
or U24751 (N_24751,N_24709,N_24526);
nor U24752 (N_24752,N_24696,N_24658);
and U24753 (N_24753,N_24684,N_24517);
or U24754 (N_24754,N_24729,N_24677);
xnor U24755 (N_24755,N_24613,N_24561);
or U24756 (N_24756,N_24650,N_24563);
nor U24757 (N_24757,N_24569,N_24548);
or U24758 (N_24758,N_24633,N_24547);
nor U24759 (N_24759,N_24701,N_24567);
xnor U24760 (N_24760,N_24745,N_24598);
or U24761 (N_24761,N_24646,N_24616);
or U24762 (N_24762,N_24659,N_24747);
or U24763 (N_24763,N_24609,N_24622);
or U24764 (N_24764,N_24726,N_24641);
nand U24765 (N_24765,N_24719,N_24566);
xnor U24766 (N_24766,N_24685,N_24558);
nor U24767 (N_24767,N_24578,N_24576);
or U24768 (N_24768,N_24509,N_24518);
xnor U24769 (N_24769,N_24668,N_24503);
and U24770 (N_24770,N_24597,N_24744);
nand U24771 (N_24771,N_24564,N_24520);
xor U24772 (N_24772,N_24557,N_24666);
nor U24773 (N_24773,N_24679,N_24608);
and U24774 (N_24774,N_24698,N_24501);
and U24775 (N_24775,N_24717,N_24675);
xnor U24776 (N_24776,N_24538,N_24645);
nor U24777 (N_24777,N_24652,N_24733);
and U24778 (N_24778,N_24721,N_24560);
xor U24779 (N_24779,N_24559,N_24507);
nand U24780 (N_24780,N_24512,N_24588);
and U24781 (N_24781,N_24690,N_24627);
nand U24782 (N_24782,N_24743,N_24740);
or U24783 (N_24783,N_24574,N_24615);
xnor U24784 (N_24784,N_24600,N_24577);
and U24785 (N_24785,N_24682,N_24692);
and U24786 (N_24786,N_24640,N_24586);
nor U24787 (N_24787,N_24704,N_24545);
nor U24788 (N_24788,N_24612,N_24625);
or U24789 (N_24789,N_24691,N_24516);
and U24790 (N_24790,N_24737,N_24632);
nor U24791 (N_24791,N_24595,N_24738);
xnor U24792 (N_24792,N_24594,N_24542);
and U24793 (N_24793,N_24746,N_24700);
and U24794 (N_24794,N_24619,N_24683);
or U24795 (N_24795,N_24637,N_24695);
and U24796 (N_24796,N_24504,N_24713);
nor U24797 (N_24797,N_24621,N_24506);
or U24798 (N_24798,N_24534,N_24669);
xnor U24799 (N_24799,N_24525,N_24749);
nor U24800 (N_24800,N_24727,N_24674);
nand U24801 (N_24801,N_24603,N_24537);
and U24802 (N_24802,N_24689,N_24541);
xor U24803 (N_24803,N_24553,N_24663);
nand U24804 (N_24804,N_24522,N_24720);
and U24805 (N_24805,N_24579,N_24723);
and U24806 (N_24806,N_24681,N_24552);
and U24807 (N_24807,N_24706,N_24549);
and U24808 (N_24808,N_24680,N_24667);
nand U24809 (N_24809,N_24571,N_24716);
nor U24810 (N_24810,N_24664,N_24617);
or U24811 (N_24811,N_24530,N_24589);
xnor U24812 (N_24812,N_24607,N_24556);
nand U24813 (N_24813,N_24546,N_24694);
or U24814 (N_24814,N_24635,N_24584);
nand U24815 (N_24815,N_24634,N_24722);
or U24816 (N_24816,N_24728,N_24630);
nor U24817 (N_24817,N_24732,N_24693);
nand U24818 (N_24818,N_24702,N_24550);
xor U24819 (N_24819,N_24573,N_24655);
and U24820 (N_24820,N_24735,N_24672);
nand U24821 (N_24821,N_24654,N_24532);
nand U24822 (N_24822,N_24724,N_24587);
xnor U24823 (N_24823,N_24585,N_24596);
nand U24824 (N_24824,N_24710,N_24629);
nor U24825 (N_24825,N_24510,N_24736);
and U24826 (N_24826,N_24741,N_24500);
or U24827 (N_24827,N_24642,N_24734);
xnor U24828 (N_24828,N_24620,N_24643);
or U24829 (N_24829,N_24593,N_24511);
and U24830 (N_24830,N_24697,N_24590);
and U24831 (N_24831,N_24656,N_24636);
nor U24832 (N_24832,N_24639,N_24686);
and U24833 (N_24833,N_24572,N_24565);
or U24834 (N_24834,N_24524,N_24688);
or U24835 (N_24835,N_24707,N_24555);
nand U24836 (N_24836,N_24624,N_24531);
or U24837 (N_24837,N_24602,N_24514);
nor U24838 (N_24838,N_24628,N_24610);
and U24839 (N_24839,N_24730,N_24583);
nor U24840 (N_24840,N_24678,N_24614);
or U24841 (N_24841,N_24551,N_24699);
or U24842 (N_24842,N_24535,N_24508);
or U24843 (N_24843,N_24581,N_24515);
nand U24844 (N_24844,N_24582,N_24539);
nand U24845 (N_24845,N_24731,N_24570);
nand U24846 (N_24846,N_24519,N_24739);
nand U24847 (N_24847,N_24653,N_24748);
and U24848 (N_24848,N_24708,N_24631);
xor U24849 (N_24849,N_24662,N_24742);
or U24850 (N_24850,N_24671,N_24676);
nor U24851 (N_24851,N_24592,N_24505);
or U24852 (N_24852,N_24544,N_24644);
and U24853 (N_24853,N_24651,N_24618);
xor U24854 (N_24854,N_24673,N_24703);
and U24855 (N_24855,N_24540,N_24523);
xnor U24856 (N_24856,N_24705,N_24647);
xor U24857 (N_24857,N_24536,N_24626);
xor U24858 (N_24858,N_24711,N_24606);
nand U24859 (N_24859,N_24568,N_24648);
nand U24860 (N_24860,N_24657,N_24623);
and U24861 (N_24861,N_24502,N_24661);
and U24862 (N_24862,N_24580,N_24543);
and U24863 (N_24863,N_24604,N_24575);
xnor U24864 (N_24864,N_24599,N_24712);
nand U24865 (N_24865,N_24529,N_24665);
nand U24866 (N_24866,N_24660,N_24718);
or U24867 (N_24867,N_24533,N_24601);
and U24868 (N_24868,N_24554,N_24521);
xnor U24869 (N_24869,N_24605,N_24638);
nor U24870 (N_24870,N_24611,N_24687);
nand U24871 (N_24871,N_24528,N_24513);
nand U24872 (N_24872,N_24649,N_24670);
or U24873 (N_24873,N_24715,N_24562);
xor U24874 (N_24874,N_24591,N_24714);
or U24875 (N_24875,N_24511,N_24687);
nand U24876 (N_24876,N_24748,N_24646);
and U24877 (N_24877,N_24526,N_24584);
xor U24878 (N_24878,N_24715,N_24612);
nand U24879 (N_24879,N_24594,N_24513);
or U24880 (N_24880,N_24582,N_24705);
nand U24881 (N_24881,N_24608,N_24651);
and U24882 (N_24882,N_24542,N_24621);
and U24883 (N_24883,N_24674,N_24506);
nor U24884 (N_24884,N_24660,N_24580);
nand U24885 (N_24885,N_24749,N_24650);
nand U24886 (N_24886,N_24632,N_24697);
nor U24887 (N_24887,N_24685,N_24681);
nor U24888 (N_24888,N_24660,N_24625);
or U24889 (N_24889,N_24656,N_24658);
and U24890 (N_24890,N_24720,N_24518);
xnor U24891 (N_24891,N_24703,N_24507);
or U24892 (N_24892,N_24603,N_24574);
and U24893 (N_24893,N_24619,N_24733);
xor U24894 (N_24894,N_24557,N_24646);
and U24895 (N_24895,N_24603,N_24628);
nor U24896 (N_24896,N_24648,N_24594);
or U24897 (N_24897,N_24685,N_24691);
xnor U24898 (N_24898,N_24620,N_24617);
and U24899 (N_24899,N_24695,N_24600);
nand U24900 (N_24900,N_24674,N_24713);
nand U24901 (N_24901,N_24685,N_24630);
nand U24902 (N_24902,N_24699,N_24740);
or U24903 (N_24903,N_24612,N_24733);
or U24904 (N_24904,N_24500,N_24625);
and U24905 (N_24905,N_24541,N_24631);
or U24906 (N_24906,N_24516,N_24618);
nor U24907 (N_24907,N_24737,N_24564);
nand U24908 (N_24908,N_24591,N_24742);
xnor U24909 (N_24909,N_24563,N_24636);
or U24910 (N_24910,N_24511,N_24581);
nor U24911 (N_24911,N_24609,N_24581);
and U24912 (N_24912,N_24583,N_24665);
and U24913 (N_24913,N_24544,N_24627);
nand U24914 (N_24914,N_24562,N_24630);
nand U24915 (N_24915,N_24587,N_24507);
or U24916 (N_24916,N_24509,N_24569);
or U24917 (N_24917,N_24599,N_24512);
xor U24918 (N_24918,N_24673,N_24534);
xnor U24919 (N_24919,N_24713,N_24698);
nor U24920 (N_24920,N_24537,N_24530);
nor U24921 (N_24921,N_24501,N_24515);
nand U24922 (N_24922,N_24681,N_24695);
and U24923 (N_24923,N_24657,N_24745);
nand U24924 (N_24924,N_24720,N_24613);
or U24925 (N_24925,N_24711,N_24527);
or U24926 (N_24926,N_24555,N_24636);
nor U24927 (N_24927,N_24723,N_24715);
nor U24928 (N_24928,N_24592,N_24735);
and U24929 (N_24929,N_24642,N_24695);
xnor U24930 (N_24930,N_24622,N_24645);
or U24931 (N_24931,N_24598,N_24521);
and U24932 (N_24932,N_24629,N_24746);
and U24933 (N_24933,N_24739,N_24647);
or U24934 (N_24934,N_24680,N_24594);
or U24935 (N_24935,N_24725,N_24632);
or U24936 (N_24936,N_24670,N_24613);
or U24937 (N_24937,N_24700,N_24628);
and U24938 (N_24938,N_24655,N_24678);
nand U24939 (N_24939,N_24593,N_24543);
or U24940 (N_24940,N_24538,N_24726);
and U24941 (N_24941,N_24726,N_24543);
nor U24942 (N_24942,N_24600,N_24699);
xor U24943 (N_24943,N_24504,N_24537);
and U24944 (N_24944,N_24733,N_24644);
nor U24945 (N_24945,N_24513,N_24553);
nor U24946 (N_24946,N_24698,N_24609);
nand U24947 (N_24947,N_24666,N_24559);
xnor U24948 (N_24948,N_24691,N_24715);
and U24949 (N_24949,N_24734,N_24505);
nor U24950 (N_24950,N_24684,N_24525);
nand U24951 (N_24951,N_24625,N_24606);
and U24952 (N_24952,N_24589,N_24615);
xnor U24953 (N_24953,N_24524,N_24584);
nor U24954 (N_24954,N_24740,N_24514);
xor U24955 (N_24955,N_24636,N_24739);
nor U24956 (N_24956,N_24740,N_24661);
nor U24957 (N_24957,N_24588,N_24508);
nor U24958 (N_24958,N_24567,N_24737);
or U24959 (N_24959,N_24657,N_24622);
nor U24960 (N_24960,N_24630,N_24545);
xnor U24961 (N_24961,N_24691,N_24663);
and U24962 (N_24962,N_24553,N_24659);
nand U24963 (N_24963,N_24600,N_24569);
or U24964 (N_24964,N_24671,N_24558);
or U24965 (N_24965,N_24589,N_24616);
or U24966 (N_24966,N_24500,N_24659);
nand U24967 (N_24967,N_24715,N_24502);
xor U24968 (N_24968,N_24512,N_24748);
nor U24969 (N_24969,N_24711,N_24516);
and U24970 (N_24970,N_24528,N_24623);
xnor U24971 (N_24971,N_24509,N_24624);
or U24972 (N_24972,N_24726,N_24739);
and U24973 (N_24973,N_24656,N_24574);
or U24974 (N_24974,N_24599,N_24559);
and U24975 (N_24975,N_24726,N_24613);
or U24976 (N_24976,N_24681,N_24650);
nor U24977 (N_24977,N_24560,N_24653);
or U24978 (N_24978,N_24626,N_24646);
and U24979 (N_24979,N_24703,N_24579);
and U24980 (N_24980,N_24739,N_24523);
and U24981 (N_24981,N_24529,N_24656);
or U24982 (N_24982,N_24621,N_24664);
or U24983 (N_24983,N_24640,N_24744);
nor U24984 (N_24984,N_24745,N_24539);
and U24985 (N_24985,N_24572,N_24543);
or U24986 (N_24986,N_24518,N_24715);
nand U24987 (N_24987,N_24662,N_24748);
nand U24988 (N_24988,N_24510,N_24691);
nor U24989 (N_24989,N_24501,N_24670);
or U24990 (N_24990,N_24568,N_24530);
nand U24991 (N_24991,N_24607,N_24705);
or U24992 (N_24992,N_24545,N_24715);
and U24993 (N_24993,N_24645,N_24560);
xor U24994 (N_24994,N_24519,N_24693);
nor U24995 (N_24995,N_24597,N_24701);
xor U24996 (N_24996,N_24582,N_24555);
xor U24997 (N_24997,N_24517,N_24605);
and U24998 (N_24998,N_24524,N_24622);
and U24999 (N_24999,N_24541,N_24511);
or UO_0 (O_0,N_24998,N_24869);
nand UO_1 (O_1,N_24877,N_24906);
and UO_2 (O_2,N_24895,N_24769);
xnor UO_3 (O_3,N_24999,N_24990);
nor UO_4 (O_4,N_24816,N_24861);
xnor UO_5 (O_5,N_24955,N_24919);
xnor UO_6 (O_6,N_24762,N_24922);
xnor UO_7 (O_7,N_24971,N_24873);
xor UO_8 (O_8,N_24767,N_24770);
xor UO_9 (O_9,N_24950,N_24864);
nor UO_10 (O_10,N_24857,N_24817);
nand UO_11 (O_11,N_24801,N_24792);
or UO_12 (O_12,N_24822,N_24995);
nand UO_13 (O_13,N_24893,N_24781);
nor UO_14 (O_14,N_24774,N_24884);
and UO_15 (O_15,N_24897,N_24917);
xor UO_16 (O_16,N_24820,N_24794);
nor UO_17 (O_17,N_24761,N_24963);
nand UO_18 (O_18,N_24848,N_24809);
nand UO_19 (O_19,N_24826,N_24982);
xnor UO_20 (O_20,N_24978,N_24789);
nor UO_21 (O_21,N_24989,N_24943);
or UO_22 (O_22,N_24850,N_24846);
nor UO_23 (O_23,N_24994,N_24968);
or UO_24 (O_24,N_24980,N_24765);
xnor UO_25 (O_25,N_24909,N_24925);
and UO_26 (O_26,N_24819,N_24904);
and UO_27 (O_27,N_24905,N_24900);
or UO_28 (O_28,N_24865,N_24983);
xnor UO_29 (O_29,N_24871,N_24992);
nand UO_30 (O_30,N_24868,N_24899);
xor UO_31 (O_31,N_24881,N_24754);
or UO_32 (O_32,N_24784,N_24876);
xor UO_33 (O_33,N_24966,N_24799);
and UO_34 (O_34,N_24973,N_24825);
and UO_35 (O_35,N_24827,N_24902);
and UO_36 (O_36,N_24987,N_24951);
or UO_37 (O_37,N_24967,N_24878);
or UO_38 (O_38,N_24785,N_24898);
xor UO_39 (O_39,N_24879,N_24824);
nor UO_40 (O_40,N_24815,N_24855);
and UO_41 (O_41,N_24757,N_24928);
nand UO_42 (O_42,N_24942,N_24993);
nand UO_43 (O_43,N_24914,N_24752);
or UO_44 (O_44,N_24964,N_24753);
nand UO_45 (O_45,N_24911,N_24800);
nand UO_46 (O_46,N_24796,N_24845);
nand UO_47 (O_47,N_24949,N_24853);
nor UO_48 (O_48,N_24933,N_24970);
nor UO_49 (O_49,N_24842,N_24930);
xnor UO_50 (O_50,N_24841,N_24953);
or UO_51 (O_51,N_24764,N_24772);
nand UO_52 (O_52,N_24874,N_24797);
or UO_53 (O_53,N_24975,N_24859);
or UO_54 (O_54,N_24870,N_24813);
xnor UO_55 (O_55,N_24939,N_24771);
nand UO_56 (O_56,N_24808,N_24838);
nand UO_57 (O_57,N_24924,N_24926);
or UO_58 (O_58,N_24768,N_24766);
or UO_59 (O_59,N_24843,N_24851);
nand UO_60 (O_60,N_24913,N_24798);
or UO_61 (O_61,N_24958,N_24823);
or UO_62 (O_62,N_24828,N_24903);
and UO_63 (O_63,N_24844,N_24831);
nor UO_64 (O_64,N_24810,N_24952);
or UO_65 (O_65,N_24920,N_24888);
nor UO_66 (O_66,N_24910,N_24821);
or UO_67 (O_67,N_24858,N_24915);
and UO_68 (O_68,N_24814,N_24974);
nand UO_69 (O_69,N_24986,N_24780);
nand UO_70 (O_70,N_24788,N_24880);
or UO_71 (O_71,N_24979,N_24847);
nand UO_72 (O_72,N_24889,N_24918);
or UO_73 (O_73,N_24887,N_24791);
xnor UO_74 (O_74,N_24901,N_24750);
nand UO_75 (O_75,N_24856,N_24991);
xor UO_76 (O_76,N_24976,N_24787);
nand UO_77 (O_77,N_24929,N_24938);
xnor UO_78 (O_78,N_24972,N_24882);
and UO_79 (O_79,N_24839,N_24946);
nor UO_80 (O_80,N_24927,N_24790);
xor UO_81 (O_81,N_24883,N_24778);
or UO_82 (O_82,N_24775,N_24829);
and UO_83 (O_83,N_24996,N_24985);
nand UO_84 (O_84,N_24830,N_24894);
and UO_85 (O_85,N_24834,N_24981);
and UO_86 (O_86,N_24934,N_24835);
or UO_87 (O_87,N_24776,N_24923);
and UO_88 (O_88,N_24954,N_24931);
or UO_89 (O_89,N_24977,N_24837);
and UO_90 (O_90,N_24751,N_24984);
nor UO_91 (O_91,N_24908,N_24782);
and UO_92 (O_92,N_24795,N_24806);
and UO_93 (O_93,N_24885,N_24965);
and UO_94 (O_94,N_24944,N_24760);
or UO_95 (O_95,N_24896,N_24892);
xor UO_96 (O_96,N_24803,N_24959);
nand UO_97 (O_97,N_24849,N_24860);
xor UO_98 (O_98,N_24805,N_24863);
or UO_99 (O_99,N_24759,N_24786);
nor UO_100 (O_100,N_24875,N_24763);
nand UO_101 (O_101,N_24969,N_24936);
nor UO_102 (O_102,N_24956,N_24862);
or UO_103 (O_103,N_24912,N_24777);
xor UO_104 (O_104,N_24921,N_24854);
and UO_105 (O_105,N_24886,N_24773);
nand UO_106 (O_106,N_24833,N_24840);
or UO_107 (O_107,N_24941,N_24812);
and UO_108 (O_108,N_24804,N_24935);
and UO_109 (O_109,N_24852,N_24807);
and UO_110 (O_110,N_24867,N_24793);
and UO_111 (O_111,N_24811,N_24907);
nand UO_112 (O_112,N_24758,N_24890);
and UO_113 (O_113,N_24945,N_24802);
nor UO_114 (O_114,N_24937,N_24891);
nand UO_115 (O_115,N_24988,N_24916);
and UO_116 (O_116,N_24932,N_24957);
nor UO_117 (O_117,N_24836,N_24866);
nand UO_118 (O_118,N_24997,N_24948);
nand UO_119 (O_119,N_24783,N_24756);
nand UO_120 (O_120,N_24947,N_24940);
and UO_121 (O_121,N_24832,N_24755);
or UO_122 (O_122,N_24872,N_24962);
nor UO_123 (O_123,N_24818,N_24960);
and UO_124 (O_124,N_24961,N_24779);
and UO_125 (O_125,N_24942,N_24845);
xnor UO_126 (O_126,N_24972,N_24799);
or UO_127 (O_127,N_24997,N_24927);
xor UO_128 (O_128,N_24806,N_24754);
nand UO_129 (O_129,N_24935,N_24778);
xor UO_130 (O_130,N_24905,N_24776);
and UO_131 (O_131,N_24992,N_24834);
nor UO_132 (O_132,N_24828,N_24957);
or UO_133 (O_133,N_24886,N_24954);
and UO_134 (O_134,N_24910,N_24768);
nand UO_135 (O_135,N_24950,N_24841);
or UO_136 (O_136,N_24878,N_24837);
and UO_137 (O_137,N_24825,N_24854);
nand UO_138 (O_138,N_24935,N_24785);
nor UO_139 (O_139,N_24970,N_24989);
and UO_140 (O_140,N_24908,N_24791);
and UO_141 (O_141,N_24962,N_24956);
nand UO_142 (O_142,N_24812,N_24953);
and UO_143 (O_143,N_24781,N_24877);
xnor UO_144 (O_144,N_24933,N_24964);
nand UO_145 (O_145,N_24844,N_24862);
xnor UO_146 (O_146,N_24810,N_24945);
nor UO_147 (O_147,N_24771,N_24930);
nand UO_148 (O_148,N_24975,N_24782);
nand UO_149 (O_149,N_24931,N_24819);
nor UO_150 (O_150,N_24854,N_24897);
or UO_151 (O_151,N_24872,N_24889);
nor UO_152 (O_152,N_24774,N_24757);
or UO_153 (O_153,N_24845,N_24868);
nand UO_154 (O_154,N_24822,N_24846);
and UO_155 (O_155,N_24777,N_24803);
nor UO_156 (O_156,N_24833,N_24780);
nor UO_157 (O_157,N_24833,N_24848);
or UO_158 (O_158,N_24802,N_24906);
xnor UO_159 (O_159,N_24805,N_24904);
xnor UO_160 (O_160,N_24901,N_24879);
or UO_161 (O_161,N_24835,N_24818);
nor UO_162 (O_162,N_24956,N_24965);
or UO_163 (O_163,N_24770,N_24762);
nor UO_164 (O_164,N_24860,N_24864);
nand UO_165 (O_165,N_24876,N_24911);
nand UO_166 (O_166,N_24882,N_24881);
nand UO_167 (O_167,N_24767,N_24894);
and UO_168 (O_168,N_24918,N_24851);
and UO_169 (O_169,N_24981,N_24919);
nor UO_170 (O_170,N_24966,N_24918);
or UO_171 (O_171,N_24890,N_24942);
nor UO_172 (O_172,N_24837,N_24793);
nand UO_173 (O_173,N_24852,N_24821);
xnor UO_174 (O_174,N_24936,N_24966);
nand UO_175 (O_175,N_24855,N_24925);
xor UO_176 (O_176,N_24817,N_24900);
or UO_177 (O_177,N_24898,N_24754);
nor UO_178 (O_178,N_24857,N_24774);
nand UO_179 (O_179,N_24822,N_24921);
nor UO_180 (O_180,N_24901,N_24787);
and UO_181 (O_181,N_24941,N_24767);
nor UO_182 (O_182,N_24762,N_24763);
nand UO_183 (O_183,N_24992,N_24911);
nor UO_184 (O_184,N_24866,N_24972);
or UO_185 (O_185,N_24771,N_24816);
xnor UO_186 (O_186,N_24971,N_24754);
nand UO_187 (O_187,N_24972,N_24833);
and UO_188 (O_188,N_24882,N_24959);
and UO_189 (O_189,N_24863,N_24871);
or UO_190 (O_190,N_24788,N_24864);
xnor UO_191 (O_191,N_24752,N_24919);
and UO_192 (O_192,N_24890,N_24787);
nor UO_193 (O_193,N_24961,N_24927);
and UO_194 (O_194,N_24816,N_24925);
nor UO_195 (O_195,N_24970,N_24834);
or UO_196 (O_196,N_24999,N_24979);
nor UO_197 (O_197,N_24913,N_24818);
xor UO_198 (O_198,N_24940,N_24852);
nor UO_199 (O_199,N_24766,N_24823);
nor UO_200 (O_200,N_24750,N_24785);
xor UO_201 (O_201,N_24945,N_24967);
and UO_202 (O_202,N_24957,N_24824);
and UO_203 (O_203,N_24933,N_24864);
nand UO_204 (O_204,N_24879,N_24827);
nor UO_205 (O_205,N_24764,N_24949);
nand UO_206 (O_206,N_24945,N_24979);
nor UO_207 (O_207,N_24784,N_24824);
or UO_208 (O_208,N_24967,N_24759);
and UO_209 (O_209,N_24852,N_24812);
nor UO_210 (O_210,N_24781,N_24752);
and UO_211 (O_211,N_24957,N_24901);
or UO_212 (O_212,N_24947,N_24857);
nand UO_213 (O_213,N_24906,N_24776);
or UO_214 (O_214,N_24959,N_24823);
nor UO_215 (O_215,N_24776,N_24926);
or UO_216 (O_216,N_24819,N_24869);
or UO_217 (O_217,N_24945,N_24868);
xnor UO_218 (O_218,N_24989,N_24934);
nor UO_219 (O_219,N_24904,N_24847);
nor UO_220 (O_220,N_24763,N_24840);
and UO_221 (O_221,N_24847,N_24924);
and UO_222 (O_222,N_24888,N_24884);
or UO_223 (O_223,N_24995,N_24872);
or UO_224 (O_224,N_24803,N_24904);
and UO_225 (O_225,N_24986,N_24854);
nand UO_226 (O_226,N_24834,N_24902);
nor UO_227 (O_227,N_24751,N_24850);
and UO_228 (O_228,N_24755,N_24917);
or UO_229 (O_229,N_24821,N_24911);
nor UO_230 (O_230,N_24902,N_24923);
and UO_231 (O_231,N_24873,N_24804);
nand UO_232 (O_232,N_24787,N_24792);
nor UO_233 (O_233,N_24876,N_24978);
nor UO_234 (O_234,N_24837,N_24895);
nor UO_235 (O_235,N_24983,N_24958);
and UO_236 (O_236,N_24935,N_24926);
nand UO_237 (O_237,N_24996,N_24861);
nor UO_238 (O_238,N_24773,N_24936);
nor UO_239 (O_239,N_24886,N_24820);
and UO_240 (O_240,N_24941,N_24903);
nor UO_241 (O_241,N_24959,N_24988);
xor UO_242 (O_242,N_24959,N_24798);
or UO_243 (O_243,N_24891,N_24847);
or UO_244 (O_244,N_24988,N_24946);
xor UO_245 (O_245,N_24833,N_24824);
and UO_246 (O_246,N_24904,N_24791);
nand UO_247 (O_247,N_24894,N_24959);
or UO_248 (O_248,N_24976,N_24857);
and UO_249 (O_249,N_24882,N_24975);
or UO_250 (O_250,N_24854,N_24954);
xor UO_251 (O_251,N_24792,N_24813);
or UO_252 (O_252,N_24832,N_24949);
nand UO_253 (O_253,N_24947,N_24932);
nand UO_254 (O_254,N_24875,N_24986);
xor UO_255 (O_255,N_24849,N_24880);
nand UO_256 (O_256,N_24919,N_24897);
nor UO_257 (O_257,N_24876,N_24958);
and UO_258 (O_258,N_24922,N_24780);
and UO_259 (O_259,N_24937,N_24919);
and UO_260 (O_260,N_24791,N_24882);
or UO_261 (O_261,N_24780,N_24913);
nand UO_262 (O_262,N_24880,N_24823);
xor UO_263 (O_263,N_24977,N_24989);
and UO_264 (O_264,N_24874,N_24775);
or UO_265 (O_265,N_24852,N_24937);
or UO_266 (O_266,N_24819,N_24814);
nor UO_267 (O_267,N_24908,N_24778);
or UO_268 (O_268,N_24990,N_24940);
and UO_269 (O_269,N_24848,N_24948);
and UO_270 (O_270,N_24955,N_24849);
nor UO_271 (O_271,N_24865,N_24930);
nand UO_272 (O_272,N_24843,N_24778);
xnor UO_273 (O_273,N_24785,N_24959);
xor UO_274 (O_274,N_24756,N_24917);
or UO_275 (O_275,N_24990,N_24776);
and UO_276 (O_276,N_24914,N_24755);
nand UO_277 (O_277,N_24889,N_24756);
nand UO_278 (O_278,N_24903,N_24907);
or UO_279 (O_279,N_24970,N_24779);
xnor UO_280 (O_280,N_24810,N_24989);
nand UO_281 (O_281,N_24946,N_24923);
or UO_282 (O_282,N_24983,N_24805);
nand UO_283 (O_283,N_24784,N_24940);
and UO_284 (O_284,N_24757,N_24771);
nor UO_285 (O_285,N_24915,N_24971);
or UO_286 (O_286,N_24916,N_24869);
xnor UO_287 (O_287,N_24846,N_24937);
nand UO_288 (O_288,N_24915,N_24796);
xnor UO_289 (O_289,N_24765,N_24951);
nand UO_290 (O_290,N_24979,N_24835);
or UO_291 (O_291,N_24941,N_24955);
or UO_292 (O_292,N_24973,N_24896);
nor UO_293 (O_293,N_24782,N_24915);
nand UO_294 (O_294,N_24894,N_24984);
xor UO_295 (O_295,N_24868,N_24870);
or UO_296 (O_296,N_24936,N_24876);
nand UO_297 (O_297,N_24763,N_24820);
or UO_298 (O_298,N_24824,N_24969);
nand UO_299 (O_299,N_24997,N_24849);
or UO_300 (O_300,N_24970,N_24788);
and UO_301 (O_301,N_24993,N_24924);
or UO_302 (O_302,N_24766,N_24953);
xnor UO_303 (O_303,N_24878,N_24888);
and UO_304 (O_304,N_24882,N_24860);
or UO_305 (O_305,N_24791,N_24781);
xnor UO_306 (O_306,N_24824,N_24929);
nand UO_307 (O_307,N_24763,N_24933);
and UO_308 (O_308,N_24886,N_24811);
xnor UO_309 (O_309,N_24965,N_24933);
or UO_310 (O_310,N_24816,N_24924);
and UO_311 (O_311,N_24761,N_24992);
nor UO_312 (O_312,N_24953,N_24756);
nand UO_313 (O_313,N_24793,N_24770);
and UO_314 (O_314,N_24920,N_24862);
xor UO_315 (O_315,N_24889,N_24927);
xnor UO_316 (O_316,N_24891,N_24956);
or UO_317 (O_317,N_24884,N_24934);
nand UO_318 (O_318,N_24998,N_24762);
nand UO_319 (O_319,N_24792,N_24969);
and UO_320 (O_320,N_24782,N_24886);
nor UO_321 (O_321,N_24768,N_24871);
or UO_322 (O_322,N_24987,N_24765);
nand UO_323 (O_323,N_24821,N_24974);
xnor UO_324 (O_324,N_24751,N_24857);
or UO_325 (O_325,N_24951,N_24946);
nor UO_326 (O_326,N_24995,N_24948);
nand UO_327 (O_327,N_24817,N_24798);
xor UO_328 (O_328,N_24916,N_24912);
and UO_329 (O_329,N_24840,N_24960);
and UO_330 (O_330,N_24802,N_24910);
and UO_331 (O_331,N_24941,N_24753);
nand UO_332 (O_332,N_24894,N_24881);
nand UO_333 (O_333,N_24982,N_24868);
nand UO_334 (O_334,N_24799,N_24949);
xor UO_335 (O_335,N_24844,N_24839);
xor UO_336 (O_336,N_24991,N_24981);
nand UO_337 (O_337,N_24900,N_24940);
xor UO_338 (O_338,N_24844,N_24921);
and UO_339 (O_339,N_24986,N_24848);
and UO_340 (O_340,N_24954,N_24938);
nand UO_341 (O_341,N_24852,N_24775);
or UO_342 (O_342,N_24833,N_24908);
nor UO_343 (O_343,N_24962,N_24849);
nor UO_344 (O_344,N_24793,N_24949);
xnor UO_345 (O_345,N_24882,N_24893);
nor UO_346 (O_346,N_24798,N_24849);
nand UO_347 (O_347,N_24782,N_24872);
or UO_348 (O_348,N_24844,N_24915);
nand UO_349 (O_349,N_24844,N_24841);
xnor UO_350 (O_350,N_24933,N_24927);
xnor UO_351 (O_351,N_24873,N_24996);
nand UO_352 (O_352,N_24752,N_24802);
and UO_353 (O_353,N_24987,N_24979);
xor UO_354 (O_354,N_24864,N_24960);
nand UO_355 (O_355,N_24767,N_24858);
nand UO_356 (O_356,N_24915,N_24875);
nor UO_357 (O_357,N_24913,N_24837);
or UO_358 (O_358,N_24906,N_24862);
or UO_359 (O_359,N_24912,N_24795);
or UO_360 (O_360,N_24992,N_24875);
and UO_361 (O_361,N_24950,N_24866);
or UO_362 (O_362,N_24975,N_24922);
xor UO_363 (O_363,N_24993,N_24910);
nor UO_364 (O_364,N_24825,N_24792);
and UO_365 (O_365,N_24906,N_24754);
nand UO_366 (O_366,N_24989,N_24882);
and UO_367 (O_367,N_24817,N_24870);
or UO_368 (O_368,N_24819,N_24805);
or UO_369 (O_369,N_24842,N_24941);
or UO_370 (O_370,N_24999,N_24792);
xnor UO_371 (O_371,N_24765,N_24846);
nand UO_372 (O_372,N_24797,N_24944);
and UO_373 (O_373,N_24766,N_24762);
or UO_374 (O_374,N_24912,N_24906);
xor UO_375 (O_375,N_24894,N_24941);
and UO_376 (O_376,N_24920,N_24842);
or UO_377 (O_377,N_24809,N_24851);
and UO_378 (O_378,N_24763,N_24967);
and UO_379 (O_379,N_24805,N_24807);
nand UO_380 (O_380,N_24989,N_24797);
xnor UO_381 (O_381,N_24796,N_24886);
or UO_382 (O_382,N_24764,N_24843);
nor UO_383 (O_383,N_24892,N_24917);
or UO_384 (O_384,N_24897,N_24959);
nand UO_385 (O_385,N_24760,N_24989);
or UO_386 (O_386,N_24790,N_24859);
and UO_387 (O_387,N_24779,N_24846);
or UO_388 (O_388,N_24997,N_24975);
or UO_389 (O_389,N_24876,N_24970);
or UO_390 (O_390,N_24756,N_24831);
or UO_391 (O_391,N_24974,N_24780);
or UO_392 (O_392,N_24777,N_24995);
or UO_393 (O_393,N_24966,N_24907);
nand UO_394 (O_394,N_24808,N_24870);
or UO_395 (O_395,N_24915,N_24770);
or UO_396 (O_396,N_24784,N_24973);
nand UO_397 (O_397,N_24906,N_24811);
xor UO_398 (O_398,N_24788,N_24977);
and UO_399 (O_399,N_24780,N_24846);
and UO_400 (O_400,N_24900,N_24913);
xor UO_401 (O_401,N_24987,N_24893);
nor UO_402 (O_402,N_24941,N_24788);
and UO_403 (O_403,N_24843,N_24797);
nand UO_404 (O_404,N_24824,N_24778);
nand UO_405 (O_405,N_24997,N_24942);
and UO_406 (O_406,N_24900,N_24939);
xor UO_407 (O_407,N_24761,N_24947);
or UO_408 (O_408,N_24931,N_24889);
or UO_409 (O_409,N_24899,N_24826);
or UO_410 (O_410,N_24903,N_24954);
xor UO_411 (O_411,N_24897,N_24802);
nor UO_412 (O_412,N_24777,N_24854);
nand UO_413 (O_413,N_24776,N_24828);
nand UO_414 (O_414,N_24852,N_24862);
xor UO_415 (O_415,N_24889,N_24871);
nor UO_416 (O_416,N_24764,N_24985);
nand UO_417 (O_417,N_24952,N_24758);
and UO_418 (O_418,N_24988,N_24765);
nand UO_419 (O_419,N_24854,N_24997);
xor UO_420 (O_420,N_24868,N_24909);
nor UO_421 (O_421,N_24792,N_24794);
and UO_422 (O_422,N_24915,N_24953);
nor UO_423 (O_423,N_24771,N_24768);
and UO_424 (O_424,N_24880,N_24786);
nor UO_425 (O_425,N_24937,N_24776);
xnor UO_426 (O_426,N_24941,N_24886);
nor UO_427 (O_427,N_24828,N_24774);
and UO_428 (O_428,N_24989,N_24902);
and UO_429 (O_429,N_24877,N_24783);
or UO_430 (O_430,N_24951,N_24950);
and UO_431 (O_431,N_24825,N_24990);
nand UO_432 (O_432,N_24993,N_24800);
and UO_433 (O_433,N_24892,N_24834);
and UO_434 (O_434,N_24755,N_24784);
xnor UO_435 (O_435,N_24974,N_24781);
xnor UO_436 (O_436,N_24816,N_24842);
nor UO_437 (O_437,N_24812,N_24979);
nor UO_438 (O_438,N_24750,N_24899);
nand UO_439 (O_439,N_24981,N_24929);
xnor UO_440 (O_440,N_24947,N_24853);
nor UO_441 (O_441,N_24828,N_24839);
and UO_442 (O_442,N_24971,N_24758);
or UO_443 (O_443,N_24998,N_24911);
nor UO_444 (O_444,N_24820,N_24912);
nor UO_445 (O_445,N_24855,N_24847);
or UO_446 (O_446,N_24964,N_24966);
or UO_447 (O_447,N_24825,N_24767);
or UO_448 (O_448,N_24956,N_24817);
nor UO_449 (O_449,N_24819,N_24852);
and UO_450 (O_450,N_24962,N_24972);
nand UO_451 (O_451,N_24857,N_24972);
or UO_452 (O_452,N_24758,N_24808);
and UO_453 (O_453,N_24836,N_24993);
and UO_454 (O_454,N_24887,N_24988);
nand UO_455 (O_455,N_24922,N_24990);
xor UO_456 (O_456,N_24841,N_24971);
and UO_457 (O_457,N_24971,N_24821);
xnor UO_458 (O_458,N_24829,N_24876);
xor UO_459 (O_459,N_24795,N_24999);
and UO_460 (O_460,N_24901,N_24862);
or UO_461 (O_461,N_24788,N_24762);
nor UO_462 (O_462,N_24963,N_24772);
nand UO_463 (O_463,N_24918,N_24873);
nand UO_464 (O_464,N_24850,N_24780);
xnor UO_465 (O_465,N_24859,N_24901);
xnor UO_466 (O_466,N_24822,N_24805);
and UO_467 (O_467,N_24810,N_24813);
nand UO_468 (O_468,N_24771,N_24846);
or UO_469 (O_469,N_24862,N_24980);
nor UO_470 (O_470,N_24897,N_24812);
and UO_471 (O_471,N_24897,N_24793);
or UO_472 (O_472,N_24892,N_24862);
nor UO_473 (O_473,N_24910,N_24871);
nand UO_474 (O_474,N_24967,N_24771);
nand UO_475 (O_475,N_24931,N_24759);
and UO_476 (O_476,N_24876,N_24839);
nand UO_477 (O_477,N_24975,N_24913);
xor UO_478 (O_478,N_24932,N_24887);
nand UO_479 (O_479,N_24976,N_24797);
xnor UO_480 (O_480,N_24925,N_24803);
or UO_481 (O_481,N_24784,N_24833);
nand UO_482 (O_482,N_24761,N_24920);
nor UO_483 (O_483,N_24984,N_24822);
xor UO_484 (O_484,N_24943,N_24913);
nand UO_485 (O_485,N_24912,N_24942);
and UO_486 (O_486,N_24927,N_24851);
nor UO_487 (O_487,N_24967,N_24975);
and UO_488 (O_488,N_24962,N_24756);
nor UO_489 (O_489,N_24935,N_24994);
or UO_490 (O_490,N_24918,N_24990);
xnor UO_491 (O_491,N_24902,N_24978);
nand UO_492 (O_492,N_24946,N_24848);
or UO_493 (O_493,N_24987,N_24766);
nor UO_494 (O_494,N_24777,N_24949);
or UO_495 (O_495,N_24960,N_24816);
or UO_496 (O_496,N_24954,N_24943);
nor UO_497 (O_497,N_24960,N_24823);
nor UO_498 (O_498,N_24753,N_24983);
xnor UO_499 (O_499,N_24882,N_24822);
or UO_500 (O_500,N_24849,N_24990);
nor UO_501 (O_501,N_24757,N_24980);
or UO_502 (O_502,N_24820,N_24931);
and UO_503 (O_503,N_24935,N_24909);
or UO_504 (O_504,N_24972,N_24899);
and UO_505 (O_505,N_24800,N_24752);
xor UO_506 (O_506,N_24921,N_24802);
nand UO_507 (O_507,N_24850,N_24753);
xor UO_508 (O_508,N_24982,N_24796);
and UO_509 (O_509,N_24937,N_24762);
nor UO_510 (O_510,N_24788,N_24846);
nand UO_511 (O_511,N_24987,N_24802);
nand UO_512 (O_512,N_24955,N_24895);
xnor UO_513 (O_513,N_24758,N_24893);
xnor UO_514 (O_514,N_24982,N_24781);
or UO_515 (O_515,N_24842,N_24773);
and UO_516 (O_516,N_24946,N_24766);
and UO_517 (O_517,N_24871,N_24993);
nand UO_518 (O_518,N_24892,N_24850);
and UO_519 (O_519,N_24897,N_24856);
or UO_520 (O_520,N_24955,N_24821);
nor UO_521 (O_521,N_24779,N_24880);
and UO_522 (O_522,N_24864,N_24907);
nor UO_523 (O_523,N_24901,N_24842);
xnor UO_524 (O_524,N_24954,N_24851);
nor UO_525 (O_525,N_24849,N_24775);
and UO_526 (O_526,N_24846,N_24998);
xor UO_527 (O_527,N_24994,N_24953);
xor UO_528 (O_528,N_24974,N_24763);
nand UO_529 (O_529,N_24845,N_24879);
xnor UO_530 (O_530,N_24788,N_24828);
xnor UO_531 (O_531,N_24966,N_24982);
and UO_532 (O_532,N_24969,N_24849);
or UO_533 (O_533,N_24962,N_24773);
or UO_534 (O_534,N_24885,N_24772);
or UO_535 (O_535,N_24952,N_24920);
xor UO_536 (O_536,N_24813,N_24791);
and UO_537 (O_537,N_24823,N_24797);
nand UO_538 (O_538,N_24965,N_24847);
and UO_539 (O_539,N_24885,N_24769);
nand UO_540 (O_540,N_24877,N_24986);
xnor UO_541 (O_541,N_24862,N_24908);
or UO_542 (O_542,N_24879,N_24828);
xor UO_543 (O_543,N_24761,N_24793);
and UO_544 (O_544,N_24955,N_24855);
and UO_545 (O_545,N_24908,N_24952);
and UO_546 (O_546,N_24757,N_24986);
or UO_547 (O_547,N_24845,N_24828);
nor UO_548 (O_548,N_24905,N_24992);
or UO_549 (O_549,N_24813,N_24789);
nor UO_550 (O_550,N_24853,N_24874);
xnor UO_551 (O_551,N_24919,N_24968);
xor UO_552 (O_552,N_24850,N_24999);
nand UO_553 (O_553,N_24770,N_24924);
or UO_554 (O_554,N_24812,N_24839);
nor UO_555 (O_555,N_24782,N_24924);
nand UO_556 (O_556,N_24796,N_24960);
nand UO_557 (O_557,N_24761,N_24989);
xnor UO_558 (O_558,N_24780,N_24950);
nand UO_559 (O_559,N_24959,N_24896);
or UO_560 (O_560,N_24967,N_24985);
nor UO_561 (O_561,N_24943,N_24805);
or UO_562 (O_562,N_24935,N_24972);
nor UO_563 (O_563,N_24914,N_24844);
and UO_564 (O_564,N_24754,N_24822);
nor UO_565 (O_565,N_24965,N_24904);
and UO_566 (O_566,N_24879,N_24937);
nand UO_567 (O_567,N_24803,N_24870);
and UO_568 (O_568,N_24761,N_24818);
and UO_569 (O_569,N_24954,N_24759);
xor UO_570 (O_570,N_24995,N_24879);
or UO_571 (O_571,N_24847,N_24966);
and UO_572 (O_572,N_24760,N_24974);
nor UO_573 (O_573,N_24998,N_24854);
and UO_574 (O_574,N_24951,N_24931);
or UO_575 (O_575,N_24839,N_24955);
and UO_576 (O_576,N_24892,N_24788);
nor UO_577 (O_577,N_24898,N_24958);
nand UO_578 (O_578,N_24948,N_24856);
or UO_579 (O_579,N_24926,N_24840);
xnor UO_580 (O_580,N_24937,N_24814);
nor UO_581 (O_581,N_24951,N_24869);
nor UO_582 (O_582,N_24866,N_24837);
or UO_583 (O_583,N_24991,N_24855);
xnor UO_584 (O_584,N_24990,N_24988);
xnor UO_585 (O_585,N_24790,N_24803);
and UO_586 (O_586,N_24844,N_24917);
or UO_587 (O_587,N_24902,N_24969);
nand UO_588 (O_588,N_24873,N_24857);
xnor UO_589 (O_589,N_24826,N_24777);
and UO_590 (O_590,N_24814,N_24811);
xor UO_591 (O_591,N_24910,N_24823);
nand UO_592 (O_592,N_24928,N_24989);
or UO_593 (O_593,N_24965,N_24999);
nor UO_594 (O_594,N_24759,N_24985);
nor UO_595 (O_595,N_24802,N_24770);
xor UO_596 (O_596,N_24799,N_24944);
nor UO_597 (O_597,N_24897,N_24756);
or UO_598 (O_598,N_24909,N_24929);
or UO_599 (O_599,N_24924,N_24841);
xnor UO_600 (O_600,N_24949,N_24878);
nand UO_601 (O_601,N_24825,N_24933);
nand UO_602 (O_602,N_24880,N_24887);
nand UO_603 (O_603,N_24858,N_24884);
or UO_604 (O_604,N_24944,N_24869);
xor UO_605 (O_605,N_24875,N_24826);
nand UO_606 (O_606,N_24882,N_24852);
or UO_607 (O_607,N_24958,N_24867);
nand UO_608 (O_608,N_24971,N_24894);
xor UO_609 (O_609,N_24912,N_24999);
xnor UO_610 (O_610,N_24792,N_24963);
and UO_611 (O_611,N_24853,N_24831);
nor UO_612 (O_612,N_24861,N_24976);
and UO_613 (O_613,N_24837,N_24830);
xor UO_614 (O_614,N_24832,N_24794);
or UO_615 (O_615,N_24992,N_24945);
and UO_616 (O_616,N_24949,N_24897);
and UO_617 (O_617,N_24874,N_24865);
and UO_618 (O_618,N_24958,N_24907);
nor UO_619 (O_619,N_24953,N_24847);
xor UO_620 (O_620,N_24899,N_24778);
nor UO_621 (O_621,N_24984,N_24953);
or UO_622 (O_622,N_24983,N_24893);
or UO_623 (O_623,N_24997,N_24993);
or UO_624 (O_624,N_24801,N_24930);
and UO_625 (O_625,N_24955,N_24983);
nor UO_626 (O_626,N_24810,N_24973);
xnor UO_627 (O_627,N_24775,N_24982);
nor UO_628 (O_628,N_24965,N_24944);
or UO_629 (O_629,N_24969,N_24861);
or UO_630 (O_630,N_24916,N_24850);
and UO_631 (O_631,N_24784,N_24858);
nor UO_632 (O_632,N_24969,N_24808);
and UO_633 (O_633,N_24990,N_24780);
or UO_634 (O_634,N_24971,N_24854);
or UO_635 (O_635,N_24822,N_24916);
nand UO_636 (O_636,N_24750,N_24801);
nor UO_637 (O_637,N_24779,N_24823);
nand UO_638 (O_638,N_24862,N_24836);
nand UO_639 (O_639,N_24842,N_24955);
xor UO_640 (O_640,N_24886,N_24837);
xor UO_641 (O_641,N_24802,N_24839);
or UO_642 (O_642,N_24756,N_24944);
nand UO_643 (O_643,N_24906,N_24951);
and UO_644 (O_644,N_24862,N_24835);
and UO_645 (O_645,N_24964,N_24999);
nand UO_646 (O_646,N_24847,N_24831);
or UO_647 (O_647,N_24804,N_24820);
and UO_648 (O_648,N_24927,N_24803);
xor UO_649 (O_649,N_24753,N_24853);
nor UO_650 (O_650,N_24775,N_24807);
or UO_651 (O_651,N_24789,N_24971);
xnor UO_652 (O_652,N_24861,N_24839);
nand UO_653 (O_653,N_24754,N_24921);
or UO_654 (O_654,N_24936,N_24814);
or UO_655 (O_655,N_24835,N_24911);
and UO_656 (O_656,N_24759,N_24890);
nor UO_657 (O_657,N_24825,N_24964);
nor UO_658 (O_658,N_24812,N_24855);
nand UO_659 (O_659,N_24792,N_24764);
nor UO_660 (O_660,N_24833,N_24993);
xor UO_661 (O_661,N_24917,N_24815);
nand UO_662 (O_662,N_24824,N_24894);
xor UO_663 (O_663,N_24993,N_24927);
or UO_664 (O_664,N_24799,N_24821);
nor UO_665 (O_665,N_24829,N_24855);
xnor UO_666 (O_666,N_24899,N_24923);
and UO_667 (O_667,N_24820,N_24962);
and UO_668 (O_668,N_24853,N_24982);
nand UO_669 (O_669,N_24771,N_24909);
and UO_670 (O_670,N_24926,N_24808);
xnor UO_671 (O_671,N_24948,N_24974);
xor UO_672 (O_672,N_24953,N_24990);
and UO_673 (O_673,N_24877,N_24788);
xnor UO_674 (O_674,N_24975,N_24981);
nand UO_675 (O_675,N_24886,N_24841);
nand UO_676 (O_676,N_24946,N_24966);
xor UO_677 (O_677,N_24956,N_24818);
xnor UO_678 (O_678,N_24975,N_24822);
nor UO_679 (O_679,N_24925,N_24950);
nand UO_680 (O_680,N_24814,N_24923);
xor UO_681 (O_681,N_24914,N_24986);
and UO_682 (O_682,N_24841,N_24984);
nand UO_683 (O_683,N_24768,N_24870);
nor UO_684 (O_684,N_24895,N_24876);
nor UO_685 (O_685,N_24788,N_24753);
or UO_686 (O_686,N_24818,N_24923);
xnor UO_687 (O_687,N_24821,N_24872);
xnor UO_688 (O_688,N_24940,N_24833);
nor UO_689 (O_689,N_24923,N_24983);
or UO_690 (O_690,N_24760,N_24926);
nand UO_691 (O_691,N_24841,N_24976);
nand UO_692 (O_692,N_24908,N_24977);
nand UO_693 (O_693,N_24990,N_24996);
and UO_694 (O_694,N_24885,N_24877);
or UO_695 (O_695,N_24845,N_24761);
or UO_696 (O_696,N_24893,N_24881);
or UO_697 (O_697,N_24938,N_24947);
nor UO_698 (O_698,N_24894,N_24819);
and UO_699 (O_699,N_24916,N_24889);
or UO_700 (O_700,N_24879,N_24997);
and UO_701 (O_701,N_24894,N_24899);
nor UO_702 (O_702,N_24768,N_24833);
nand UO_703 (O_703,N_24845,N_24985);
nand UO_704 (O_704,N_24762,N_24751);
nand UO_705 (O_705,N_24988,N_24927);
or UO_706 (O_706,N_24760,N_24887);
nor UO_707 (O_707,N_24899,N_24960);
nand UO_708 (O_708,N_24820,N_24873);
xor UO_709 (O_709,N_24930,N_24832);
and UO_710 (O_710,N_24832,N_24764);
xnor UO_711 (O_711,N_24958,N_24843);
and UO_712 (O_712,N_24866,N_24929);
xnor UO_713 (O_713,N_24933,N_24944);
xnor UO_714 (O_714,N_24846,N_24883);
nand UO_715 (O_715,N_24952,N_24796);
nand UO_716 (O_716,N_24931,N_24755);
nor UO_717 (O_717,N_24964,N_24814);
and UO_718 (O_718,N_24934,N_24976);
nor UO_719 (O_719,N_24848,N_24969);
nor UO_720 (O_720,N_24874,N_24903);
and UO_721 (O_721,N_24973,N_24897);
or UO_722 (O_722,N_24981,N_24800);
nand UO_723 (O_723,N_24762,N_24993);
nor UO_724 (O_724,N_24939,N_24767);
and UO_725 (O_725,N_24893,N_24773);
nor UO_726 (O_726,N_24852,N_24916);
and UO_727 (O_727,N_24782,N_24777);
nor UO_728 (O_728,N_24900,N_24789);
nand UO_729 (O_729,N_24754,N_24788);
xnor UO_730 (O_730,N_24914,N_24994);
or UO_731 (O_731,N_24891,N_24790);
or UO_732 (O_732,N_24889,N_24844);
and UO_733 (O_733,N_24822,N_24938);
nand UO_734 (O_734,N_24923,N_24907);
xor UO_735 (O_735,N_24851,N_24837);
nor UO_736 (O_736,N_24820,N_24812);
and UO_737 (O_737,N_24769,N_24751);
and UO_738 (O_738,N_24936,N_24867);
and UO_739 (O_739,N_24982,N_24899);
nand UO_740 (O_740,N_24944,N_24905);
nand UO_741 (O_741,N_24917,N_24954);
xor UO_742 (O_742,N_24917,N_24997);
xor UO_743 (O_743,N_24810,N_24853);
or UO_744 (O_744,N_24818,N_24943);
nand UO_745 (O_745,N_24995,N_24962);
and UO_746 (O_746,N_24994,N_24997);
nand UO_747 (O_747,N_24989,N_24992);
and UO_748 (O_748,N_24893,N_24925);
xor UO_749 (O_749,N_24967,N_24841);
and UO_750 (O_750,N_24826,N_24914);
nor UO_751 (O_751,N_24952,N_24779);
or UO_752 (O_752,N_24986,N_24755);
nand UO_753 (O_753,N_24776,N_24999);
and UO_754 (O_754,N_24841,N_24782);
nor UO_755 (O_755,N_24755,N_24951);
or UO_756 (O_756,N_24923,N_24816);
nand UO_757 (O_757,N_24831,N_24839);
nor UO_758 (O_758,N_24968,N_24952);
xor UO_759 (O_759,N_24762,N_24796);
xnor UO_760 (O_760,N_24757,N_24917);
and UO_761 (O_761,N_24905,N_24988);
nand UO_762 (O_762,N_24791,N_24999);
or UO_763 (O_763,N_24811,N_24767);
nand UO_764 (O_764,N_24765,N_24854);
and UO_765 (O_765,N_24753,N_24761);
xor UO_766 (O_766,N_24786,N_24979);
nor UO_767 (O_767,N_24770,N_24935);
nor UO_768 (O_768,N_24767,N_24840);
nand UO_769 (O_769,N_24898,N_24855);
nand UO_770 (O_770,N_24781,N_24999);
and UO_771 (O_771,N_24857,N_24932);
nand UO_772 (O_772,N_24918,N_24984);
nor UO_773 (O_773,N_24863,N_24937);
xnor UO_774 (O_774,N_24765,N_24750);
nand UO_775 (O_775,N_24971,N_24773);
xor UO_776 (O_776,N_24847,N_24814);
nand UO_777 (O_777,N_24770,N_24794);
nor UO_778 (O_778,N_24883,N_24895);
nor UO_779 (O_779,N_24865,N_24905);
or UO_780 (O_780,N_24751,N_24962);
xor UO_781 (O_781,N_24820,N_24971);
xor UO_782 (O_782,N_24809,N_24951);
nand UO_783 (O_783,N_24870,N_24782);
xnor UO_784 (O_784,N_24771,N_24999);
nor UO_785 (O_785,N_24939,N_24760);
or UO_786 (O_786,N_24903,N_24942);
and UO_787 (O_787,N_24933,N_24901);
xnor UO_788 (O_788,N_24963,N_24763);
nand UO_789 (O_789,N_24959,N_24850);
xor UO_790 (O_790,N_24870,N_24750);
nor UO_791 (O_791,N_24831,N_24771);
and UO_792 (O_792,N_24924,N_24927);
xor UO_793 (O_793,N_24791,N_24886);
and UO_794 (O_794,N_24959,N_24931);
nand UO_795 (O_795,N_24977,N_24966);
nor UO_796 (O_796,N_24978,N_24796);
or UO_797 (O_797,N_24888,N_24964);
nor UO_798 (O_798,N_24821,N_24908);
nor UO_799 (O_799,N_24817,N_24998);
nand UO_800 (O_800,N_24843,N_24918);
nand UO_801 (O_801,N_24807,N_24942);
nor UO_802 (O_802,N_24771,N_24804);
and UO_803 (O_803,N_24921,N_24907);
or UO_804 (O_804,N_24807,N_24950);
or UO_805 (O_805,N_24902,N_24926);
and UO_806 (O_806,N_24994,N_24897);
and UO_807 (O_807,N_24968,N_24878);
or UO_808 (O_808,N_24814,N_24985);
and UO_809 (O_809,N_24761,N_24974);
xnor UO_810 (O_810,N_24943,N_24982);
and UO_811 (O_811,N_24926,N_24930);
xor UO_812 (O_812,N_24909,N_24786);
or UO_813 (O_813,N_24986,N_24840);
and UO_814 (O_814,N_24823,N_24870);
nor UO_815 (O_815,N_24874,N_24790);
nand UO_816 (O_816,N_24862,N_24810);
and UO_817 (O_817,N_24859,N_24957);
xnor UO_818 (O_818,N_24941,N_24978);
or UO_819 (O_819,N_24806,N_24955);
xor UO_820 (O_820,N_24811,N_24809);
and UO_821 (O_821,N_24805,N_24833);
xor UO_822 (O_822,N_24894,N_24857);
and UO_823 (O_823,N_24831,N_24793);
or UO_824 (O_824,N_24767,N_24978);
or UO_825 (O_825,N_24822,N_24892);
or UO_826 (O_826,N_24961,N_24906);
nand UO_827 (O_827,N_24910,N_24927);
and UO_828 (O_828,N_24947,N_24804);
and UO_829 (O_829,N_24791,N_24848);
and UO_830 (O_830,N_24791,N_24866);
nand UO_831 (O_831,N_24755,N_24934);
nand UO_832 (O_832,N_24881,N_24788);
nor UO_833 (O_833,N_24987,N_24757);
nor UO_834 (O_834,N_24893,N_24762);
nor UO_835 (O_835,N_24821,N_24843);
nand UO_836 (O_836,N_24994,N_24956);
nor UO_837 (O_837,N_24902,N_24829);
xnor UO_838 (O_838,N_24848,N_24874);
xor UO_839 (O_839,N_24886,N_24784);
or UO_840 (O_840,N_24767,N_24867);
or UO_841 (O_841,N_24936,N_24794);
nor UO_842 (O_842,N_24959,N_24876);
nor UO_843 (O_843,N_24781,N_24873);
xor UO_844 (O_844,N_24890,N_24825);
nor UO_845 (O_845,N_24815,N_24766);
nor UO_846 (O_846,N_24910,N_24771);
or UO_847 (O_847,N_24863,N_24886);
and UO_848 (O_848,N_24966,N_24795);
or UO_849 (O_849,N_24798,N_24992);
xor UO_850 (O_850,N_24896,N_24913);
or UO_851 (O_851,N_24784,N_24794);
nand UO_852 (O_852,N_24849,N_24940);
and UO_853 (O_853,N_24900,N_24935);
nor UO_854 (O_854,N_24946,N_24987);
nor UO_855 (O_855,N_24776,N_24836);
nand UO_856 (O_856,N_24962,N_24923);
or UO_857 (O_857,N_24982,N_24926);
and UO_858 (O_858,N_24767,N_24926);
or UO_859 (O_859,N_24998,N_24913);
nand UO_860 (O_860,N_24860,N_24914);
nand UO_861 (O_861,N_24864,N_24803);
xor UO_862 (O_862,N_24760,N_24814);
nand UO_863 (O_863,N_24769,N_24817);
nand UO_864 (O_864,N_24894,N_24845);
and UO_865 (O_865,N_24864,N_24941);
xnor UO_866 (O_866,N_24900,N_24841);
and UO_867 (O_867,N_24913,N_24756);
nand UO_868 (O_868,N_24957,N_24753);
xnor UO_869 (O_869,N_24820,N_24995);
and UO_870 (O_870,N_24971,N_24964);
nor UO_871 (O_871,N_24861,N_24856);
nor UO_872 (O_872,N_24963,N_24794);
xnor UO_873 (O_873,N_24889,N_24934);
xnor UO_874 (O_874,N_24929,N_24888);
xor UO_875 (O_875,N_24944,N_24960);
nand UO_876 (O_876,N_24761,N_24787);
nand UO_877 (O_877,N_24937,N_24792);
and UO_878 (O_878,N_24753,N_24909);
xor UO_879 (O_879,N_24911,N_24810);
nand UO_880 (O_880,N_24788,N_24958);
nor UO_881 (O_881,N_24936,N_24882);
nor UO_882 (O_882,N_24952,N_24893);
nor UO_883 (O_883,N_24895,N_24872);
xnor UO_884 (O_884,N_24991,N_24841);
and UO_885 (O_885,N_24801,N_24762);
and UO_886 (O_886,N_24992,N_24839);
nand UO_887 (O_887,N_24794,N_24918);
xor UO_888 (O_888,N_24771,N_24894);
nand UO_889 (O_889,N_24984,N_24780);
nor UO_890 (O_890,N_24942,N_24918);
xor UO_891 (O_891,N_24861,N_24834);
or UO_892 (O_892,N_24972,N_24797);
nand UO_893 (O_893,N_24759,N_24971);
and UO_894 (O_894,N_24923,N_24823);
and UO_895 (O_895,N_24815,N_24994);
xnor UO_896 (O_896,N_24760,N_24761);
nand UO_897 (O_897,N_24905,N_24761);
nand UO_898 (O_898,N_24773,N_24862);
and UO_899 (O_899,N_24983,N_24898);
and UO_900 (O_900,N_24781,N_24952);
nor UO_901 (O_901,N_24928,N_24842);
nand UO_902 (O_902,N_24832,N_24825);
or UO_903 (O_903,N_24867,N_24881);
nor UO_904 (O_904,N_24969,N_24835);
nand UO_905 (O_905,N_24908,N_24996);
and UO_906 (O_906,N_24981,N_24997);
nand UO_907 (O_907,N_24767,N_24874);
or UO_908 (O_908,N_24956,N_24878);
xor UO_909 (O_909,N_24757,N_24792);
or UO_910 (O_910,N_24975,N_24784);
nor UO_911 (O_911,N_24825,N_24764);
xnor UO_912 (O_912,N_24883,N_24990);
or UO_913 (O_913,N_24970,N_24995);
nor UO_914 (O_914,N_24950,N_24996);
and UO_915 (O_915,N_24769,N_24822);
and UO_916 (O_916,N_24889,N_24857);
or UO_917 (O_917,N_24952,N_24775);
or UO_918 (O_918,N_24855,N_24838);
or UO_919 (O_919,N_24809,N_24916);
nor UO_920 (O_920,N_24835,N_24767);
nand UO_921 (O_921,N_24991,N_24902);
xor UO_922 (O_922,N_24929,N_24973);
or UO_923 (O_923,N_24858,N_24853);
nand UO_924 (O_924,N_24812,N_24827);
or UO_925 (O_925,N_24770,N_24862);
nor UO_926 (O_926,N_24923,N_24770);
nand UO_927 (O_927,N_24944,N_24938);
nor UO_928 (O_928,N_24750,N_24982);
nor UO_929 (O_929,N_24945,N_24923);
nand UO_930 (O_930,N_24832,N_24999);
nand UO_931 (O_931,N_24784,N_24952);
and UO_932 (O_932,N_24838,N_24969);
or UO_933 (O_933,N_24890,N_24874);
nand UO_934 (O_934,N_24787,N_24962);
xnor UO_935 (O_935,N_24786,N_24866);
and UO_936 (O_936,N_24992,N_24837);
and UO_937 (O_937,N_24803,N_24928);
nor UO_938 (O_938,N_24938,N_24914);
or UO_939 (O_939,N_24970,N_24865);
nor UO_940 (O_940,N_24803,N_24794);
xor UO_941 (O_941,N_24873,N_24875);
and UO_942 (O_942,N_24939,N_24982);
or UO_943 (O_943,N_24806,N_24973);
or UO_944 (O_944,N_24808,N_24846);
and UO_945 (O_945,N_24941,N_24942);
or UO_946 (O_946,N_24889,N_24863);
or UO_947 (O_947,N_24843,N_24969);
nand UO_948 (O_948,N_24889,N_24965);
xnor UO_949 (O_949,N_24980,N_24893);
nand UO_950 (O_950,N_24893,N_24785);
xnor UO_951 (O_951,N_24932,N_24774);
nand UO_952 (O_952,N_24970,N_24859);
xnor UO_953 (O_953,N_24959,N_24758);
nor UO_954 (O_954,N_24950,N_24885);
xor UO_955 (O_955,N_24751,N_24875);
xnor UO_956 (O_956,N_24878,N_24759);
or UO_957 (O_957,N_24889,N_24850);
and UO_958 (O_958,N_24955,N_24782);
and UO_959 (O_959,N_24963,N_24971);
nor UO_960 (O_960,N_24823,N_24811);
nand UO_961 (O_961,N_24871,N_24935);
nor UO_962 (O_962,N_24946,N_24961);
nand UO_963 (O_963,N_24936,N_24975);
nor UO_964 (O_964,N_24876,N_24885);
nand UO_965 (O_965,N_24847,N_24834);
or UO_966 (O_966,N_24994,N_24981);
or UO_967 (O_967,N_24979,N_24831);
or UO_968 (O_968,N_24868,N_24862);
nand UO_969 (O_969,N_24806,N_24830);
xnor UO_970 (O_970,N_24926,N_24786);
xor UO_971 (O_971,N_24921,N_24820);
or UO_972 (O_972,N_24783,N_24981);
xor UO_973 (O_973,N_24754,N_24901);
nand UO_974 (O_974,N_24947,N_24789);
xnor UO_975 (O_975,N_24825,N_24932);
xor UO_976 (O_976,N_24833,N_24891);
or UO_977 (O_977,N_24993,N_24940);
nand UO_978 (O_978,N_24883,N_24979);
and UO_979 (O_979,N_24868,N_24966);
xor UO_980 (O_980,N_24777,N_24865);
and UO_981 (O_981,N_24826,N_24989);
nand UO_982 (O_982,N_24757,N_24991);
nand UO_983 (O_983,N_24971,N_24868);
nor UO_984 (O_984,N_24822,N_24786);
or UO_985 (O_985,N_24857,N_24824);
nor UO_986 (O_986,N_24874,N_24880);
nor UO_987 (O_987,N_24857,N_24944);
nor UO_988 (O_988,N_24761,N_24770);
xor UO_989 (O_989,N_24993,N_24918);
nor UO_990 (O_990,N_24832,N_24874);
nand UO_991 (O_991,N_24816,N_24848);
nand UO_992 (O_992,N_24801,N_24894);
nor UO_993 (O_993,N_24762,N_24752);
nand UO_994 (O_994,N_24959,N_24996);
or UO_995 (O_995,N_24908,N_24934);
and UO_996 (O_996,N_24910,N_24827);
or UO_997 (O_997,N_24834,N_24859);
nand UO_998 (O_998,N_24940,N_24897);
xor UO_999 (O_999,N_24957,N_24960);
or UO_1000 (O_1000,N_24938,N_24851);
nand UO_1001 (O_1001,N_24971,N_24809);
nand UO_1002 (O_1002,N_24782,N_24878);
nor UO_1003 (O_1003,N_24830,N_24817);
nand UO_1004 (O_1004,N_24864,N_24938);
nand UO_1005 (O_1005,N_24946,N_24903);
or UO_1006 (O_1006,N_24841,N_24946);
or UO_1007 (O_1007,N_24829,N_24827);
nor UO_1008 (O_1008,N_24852,N_24886);
nand UO_1009 (O_1009,N_24912,N_24773);
xor UO_1010 (O_1010,N_24768,N_24907);
or UO_1011 (O_1011,N_24835,N_24850);
xnor UO_1012 (O_1012,N_24770,N_24985);
nor UO_1013 (O_1013,N_24833,N_24813);
nor UO_1014 (O_1014,N_24896,N_24856);
or UO_1015 (O_1015,N_24781,N_24935);
nand UO_1016 (O_1016,N_24783,N_24789);
or UO_1017 (O_1017,N_24861,N_24926);
or UO_1018 (O_1018,N_24940,N_24835);
nor UO_1019 (O_1019,N_24851,N_24947);
xor UO_1020 (O_1020,N_24782,N_24937);
or UO_1021 (O_1021,N_24854,N_24949);
nor UO_1022 (O_1022,N_24858,N_24765);
or UO_1023 (O_1023,N_24772,N_24986);
or UO_1024 (O_1024,N_24824,N_24807);
nand UO_1025 (O_1025,N_24940,N_24982);
xor UO_1026 (O_1026,N_24773,N_24775);
and UO_1027 (O_1027,N_24861,N_24925);
and UO_1028 (O_1028,N_24754,N_24946);
nor UO_1029 (O_1029,N_24870,N_24886);
nand UO_1030 (O_1030,N_24763,N_24809);
and UO_1031 (O_1031,N_24854,N_24936);
and UO_1032 (O_1032,N_24968,N_24785);
and UO_1033 (O_1033,N_24764,N_24909);
or UO_1034 (O_1034,N_24851,N_24901);
nor UO_1035 (O_1035,N_24799,N_24982);
nand UO_1036 (O_1036,N_24888,N_24872);
nor UO_1037 (O_1037,N_24889,N_24841);
xnor UO_1038 (O_1038,N_24752,N_24873);
and UO_1039 (O_1039,N_24756,N_24933);
xnor UO_1040 (O_1040,N_24911,N_24897);
or UO_1041 (O_1041,N_24920,N_24779);
or UO_1042 (O_1042,N_24896,N_24870);
and UO_1043 (O_1043,N_24890,N_24868);
nor UO_1044 (O_1044,N_24751,N_24766);
nor UO_1045 (O_1045,N_24896,N_24961);
or UO_1046 (O_1046,N_24797,N_24804);
nor UO_1047 (O_1047,N_24995,N_24846);
or UO_1048 (O_1048,N_24819,N_24785);
nand UO_1049 (O_1049,N_24864,N_24952);
and UO_1050 (O_1050,N_24813,N_24757);
nor UO_1051 (O_1051,N_24835,N_24755);
or UO_1052 (O_1052,N_24948,N_24872);
nor UO_1053 (O_1053,N_24815,N_24804);
nor UO_1054 (O_1054,N_24910,N_24946);
nand UO_1055 (O_1055,N_24978,N_24851);
or UO_1056 (O_1056,N_24848,N_24895);
nor UO_1057 (O_1057,N_24921,N_24841);
xnor UO_1058 (O_1058,N_24797,N_24964);
and UO_1059 (O_1059,N_24909,N_24906);
xnor UO_1060 (O_1060,N_24762,N_24761);
xnor UO_1061 (O_1061,N_24963,N_24954);
nor UO_1062 (O_1062,N_24876,N_24905);
nand UO_1063 (O_1063,N_24913,N_24931);
nand UO_1064 (O_1064,N_24763,N_24920);
nand UO_1065 (O_1065,N_24979,N_24953);
nand UO_1066 (O_1066,N_24813,N_24780);
nand UO_1067 (O_1067,N_24952,N_24772);
and UO_1068 (O_1068,N_24755,N_24945);
xnor UO_1069 (O_1069,N_24927,N_24953);
or UO_1070 (O_1070,N_24844,N_24985);
nor UO_1071 (O_1071,N_24918,N_24864);
xnor UO_1072 (O_1072,N_24903,N_24986);
xnor UO_1073 (O_1073,N_24824,N_24898);
nor UO_1074 (O_1074,N_24814,N_24765);
xnor UO_1075 (O_1075,N_24990,N_24764);
or UO_1076 (O_1076,N_24995,N_24892);
and UO_1077 (O_1077,N_24821,N_24820);
nor UO_1078 (O_1078,N_24904,N_24941);
and UO_1079 (O_1079,N_24862,N_24903);
and UO_1080 (O_1080,N_24997,N_24765);
and UO_1081 (O_1081,N_24989,N_24753);
nor UO_1082 (O_1082,N_24884,N_24775);
nor UO_1083 (O_1083,N_24898,N_24843);
or UO_1084 (O_1084,N_24800,N_24751);
nor UO_1085 (O_1085,N_24887,N_24778);
and UO_1086 (O_1086,N_24914,N_24801);
nor UO_1087 (O_1087,N_24838,N_24760);
nand UO_1088 (O_1088,N_24984,N_24813);
and UO_1089 (O_1089,N_24793,N_24765);
and UO_1090 (O_1090,N_24945,N_24866);
xnor UO_1091 (O_1091,N_24858,N_24989);
nor UO_1092 (O_1092,N_24811,N_24937);
nor UO_1093 (O_1093,N_24925,N_24936);
and UO_1094 (O_1094,N_24838,N_24872);
xnor UO_1095 (O_1095,N_24826,N_24833);
nor UO_1096 (O_1096,N_24969,N_24891);
nor UO_1097 (O_1097,N_24842,N_24782);
nand UO_1098 (O_1098,N_24871,N_24853);
nand UO_1099 (O_1099,N_24887,N_24909);
nor UO_1100 (O_1100,N_24834,N_24986);
and UO_1101 (O_1101,N_24767,N_24971);
or UO_1102 (O_1102,N_24960,N_24798);
and UO_1103 (O_1103,N_24903,N_24970);
xor UO_1104 (O_1104,N_24852,N_24771);
and UO_1105 (O_1105,N_24938,N_24926);
or UO_1106 (O_1106,N_24881,N_24986);
or UO_1107 (O_1107,N_24882,N_24907);
or UO_1108 (O_1108,N_24756,N_24762);
xnor UO_1109 (O_1109,N_24752,N_24857);
and UO_1110 (O_1110,N_24925,N_24790);
or UO_1111 (O_1111,N_24935,N_24793);
or UO_1112 (O_1112,N_24934,N_24839);
xor UO_1113 (O_1113,N_24935,N_24774);
nand UO_1114 (O_1114,N_24824,N_24869);
nor UO_1115 (O_1115,N_24810,N_24868);
nand UO_1116 (O_1116,N_24843,N_24914);
or UO_1117 (O_1117,N_24798,N_24928);
nand UO_1118 (O_1118,N_24767,N_24920);
xnor UO_1119 (O_1119,N_24844,N_24830);
nor UO_1120 (O_1120,N_24985,N_24942);
and UO_1121 (O_1121,N_24806,N_24961);
and UO_1122 (O_1122,N_24811,N_24768);
and UO_1123 (O_1123,N_24813,N_24995);
nor UO_1124 (O_1124,N_24798,N_24938);
nand UO_1125 (O_1125,N_24827,N_24825);
nor UO_1126 (O_1126,N_24979,N_24875);
or UO_1127 (O_1127,N_24773,N_24877);
xnor UO_1128 (O_1128,N_24885,N_24873);
nand UO_1129 (O_1129,N_24763,N_24943);
and UO_1130 (O_1130,N_24955,N_24887);
xnor UO_1131 (O_1131,N_24903,N_24911);
or UO_1132 (O_1132,N_24859,N_24921);
or UO_1133 (O_1133,N_24908,N_24923);
xor UO_1134 (O_1134,N_24911,N_24826);
nand UO_1135 (O_1135,N_24896,N_24865);
and UO_1136 (O_1136,N_24806,N_24982);
xnor UO_1137 (O_1137,N_24781,N_24838);
nand UO_1138 (O_1138,N_24753,N_24849);
nand UO_1139 (O_1139,N_24805,N_24830);
and UO_1140 (O_1140,N_24913,N_24979);
xor UO_1141 (O_1141,N_24968,N_24941);
and UO_1142 (O_1142,N_24854,N_24992);
or UO_1143 (O_1143,N_24880,N_24791);
nand UO_1144 (O_1144,N_24960,N_24765);
or UO_1145 (O_1145,N_24942,N_24755);
nor UO_1146 (O_1146,N_24952,N_24820);
and UO_1147 (O_1147,N_24762,N_24879);
xnor UO_1148 (O_1148,N_24784,N_24991);
or UO_1149 (O_1149,N_24807,N_24796);
or UO_1150 (O_1150,N_24978,N_24962);
nand UO_1151 (O_1151,N_24900,N_24950);
or UO_1152 (O_1152,N_24953,N_24968);
or UO_1153 (O_1153,N_24876,N_24931);
and UO_1154 (O_1154,N_24900,N_24867);
xnor UO_1155 (O_1155,N_24800,N_24872);
nor UO_1156 (O_1156,N_24924,N_24894);
xor UO_1157 (O_1157,N_24874,N_24944);
nor UO_1158 (O_1158,N_24951,N_24789);
or UO_1159 (O_1159,N_24980,N_24950);
nand UO_1160 (O_1160,N_24773,N_24997);
xnor UO_1161 (O_1161,N_24763,N_24797);
nor UO_1162 (O_1162,N_24779,N_24989);
xnor UO_1163 (O_1163,N_24922,N_24850);
and UO_1164 (O_1164,N_24834,N_24846);
and UO_1165 (O_1165,N_24835,N_24967);
nand UO_1166 (O_1166,N_24988,N_24960);
nor UO_1167 (O_1167,N_24824,N_24993);
nand UO_1168 (O_1168,N_24999,N_24800);
nor UO_1169 (O_1169,N_24784,N_24990);
xor UO_1170 (O_1170,N_24761,N_24979);
and UO_1171 (O_1171,N_24900,N_24930);
xor UO_1172 (O_1172,N_24753,N_24787);
xor UO_1173 (O_1173,N_24794,N_24796);
or UO_1174 (O_1174,N_24896,N_24842);
nor UO_1175 (O_1175,N_24777,N_24772);
nor UO_1176 (O_1176,N_24931,N_24845);
nand UO_1177 (O_1177,N_24977,N_24941);
or UO_1178 (O_1178,N_24832,N_24876);
nand UO_1179 (O_1179,N_24854,N_24787);
xor UO_1180 (O_1180,N_24751,N_24941);
xnor UO_1181 (O_1181,N_24780,N_24753);
nor UO_1182 (O_1182,N_24975,N_24934);
nor UO_1183 (O_1183,N_24862,N_24911);
and UO_1184 (O_1184,N_24965,N_24873);
nor UO_1185 (O_1185,N_24886,N_24912);
xor UO_1186 (O_1186,N_24780,N_24857);
xor UO_1187 (O_1187,N_24957,N_24914);
and UO_1188 (O_1188,N_24843,N_24857);
nand UO_1189 (O_1189,N_24915,N_24855);
or UO_1190 (O_1190,N_24866,N_24824);
or UO_1191 (O_1191,N_24906,N_24970);
nor UO_1192 (O_1192,N_24983,N_24751);
nand UO_1193 (O_1193,N_24852,N_24828);
xnor UO_1194 (O_1194,N_24792,N_24892);
and UO_1195 (O_1195,N_24767,N_24891);
xnor UO_1196 (O_1196,N_24984,N_24957);
xnor UO_1197 (O_1197,N_24756,N_24947);
nor UO_1198 (O_1198,N_24879,N_24811);
nor UO_1199 (O_1199,N_24780,N_24925);
nand UO_1200 (O_1200,N_24940,N_24823);
or UO_1201 (O_1201,N_24767,N_24962);
and UO_1202 (O_1202,N_24834,N_24905);
and UO_1203 (O_1203,N_24991,N_24955);
xor UO_1204 (O_1204,N_24800,N_24862);
xor UO_1205 (O_1205,N_24909,N_24893);
nor UO_1206 (O_1206,N_24878,N_24806);
xor UO_1207 (O_1207,N_24756,N_24869);
and UO_1208 (O_1208,N_24770,N_24910);
nor UO_1209 (O_1209,N_24788,N_24837);
nor UO_1210 (O_1210,N_24878,N_24810);
and UO_1211 (O_1211,N_24779,N_24979);
xnor UO_1212 (O_1212,N_24841,N_24859);
nor UO_1213 (O_1213,N_24845,N_24842);
nor UO_1214 (O_1214,N_24946,N_24849);
or UO_1215 (O_1215,N_24996,N_24806);
nor UO_1216 (O_1216,N_24765,N_24778);
xor UO_1217 (O_1217,N_24963,N_24879);
nand UO_1218 (O_1218,N_24851,N_24992);
or UO_1219 (O_1219,N_24784,N_24807);
xnor UO_1220 (O_1220,N_24994,N_24961);
and UO_1221 (O_1221,N_24915,N_24916);
or UO_1222 (O_1222,N_24755,N_24795);
nor UO_1223 (O_1223,N_24843,N_24893);
nand UO_1224 (O_1224,N_24752,N_24932);
nor UO_1225 (O_1225,N_24862,N_24957);
or UO_1226 (O_1226,N_24873,N_24967);
and UO_1227 (O_1227,N_24879,N_24872);
or UO_1228 (O_1228,N_24973,N_24750);
nor UO_1229 (O_1229,N_24771,N_24792);
or UO_1230 (O_1230,N_24854,N_24786);
xnor UO_1231 (O_1231,N_24760,N_24959);
and UO_1232 (O_1232,N_24789,N_24860);
and UO_1233 (O_1233,N_24782,N_24858);
and UO_1234 (O_1234,N_24878,N_24948);
nand UO_1235 (O_1235,N_24815,N_24788);
nand UO_1236 (O_1236,N_24839,N_24863);
xnor UO_1237 (O_1237,N_24978,N_24853);
or UO_1238 (O_1238,N_24866,N_24873);
nand UO_1239 (O_1239,N_24920,N_24924);
nand UO_1240 (O_1240,N_24981,N_24946);
nor UO_1241 (O_1241,N_24949,N_24959);
nor UO_1242 (O_1242,N_24789,N_24933);
and UO_1243 (O_1243,N_24858,N_24761);
and UO_1244 (O_1244,N_24902,N_24866);
nor UO_1245 (O_1245,N_24759,N_24921);
xnor UO_1246 (O_1246,N_24913,N_24831);
nor UO_1247 (O_1247,N_24855,N_24827);
nand UO_1248 (O_1248,N_24924,N_24791);
or UO_1249 (O_1249,N_24821,N_24897);
xnor UO_1250 (O_1250,N_24787,N_24848);
nand UO_1251 (O_1251,N_24935,N_24862);
nand UO_1252 (O_1252,N_24971,N_24892);
nor UO_1253 (O_1253,N_24766,N_24927);
xor UO_1254 (O_1254,N_24843,N_24982);
or UO_1255 (O_1255,N_24892,N_24967);
xnor UO_1256 (O_1256,N_24884,N_24892);
xnor UO_1257 (O_1257,N_24884,N_24849);
xnor UO_1258 (O_1258,N_24937,N_24874);
xor UO_1259 (O_1259,N_24857,N_24801);
or UO_1260 (O_1260,N_24937,N_24808);
or UO_1261 (O_1261,N_24782,N_24988);
nor UO_1262 (O_1262,N_24765,N_24836);
nor UO_1263 (O_1263,N_24877,N_24965);
and UO_1264 (O_1264,N_24973,N_24766);
xor UO_1265 (O_1265,N_24767,N_24854);
nor UO_1266 (O_1266,N_24931,N_24840);
and UO_1267 (O_1267,N_24841,N_24834);
or UO_1268 (O_1268,N_24800,N_24860);
or UO_1269 (O_1269,N_24936,N_24894);
nor UO_1270 (O_1270,N_24981,N_24802);
nand UO_1271 (O_1271,N_24972,N_24978);
nand UO_1272 (O_1272,N_24850,N_24856);
or UO_1273 (O_1273,N_24977,N_24930);
nand UO_1274 (O_1274,N_24795,N_24786);
nor UO_1275 (O_1275,N_24854,N_24991);
nand UO_1276 (O_1276,N_24939,N_24932);
or UO_1277 (O_1277,N_24927,N_24863);
xnor UO_1278 (O_1278,N_24992,N_24850);
and UO_1279 (O_1279,N_24898,N_24797);
or UO_1280 (O_1280,N_24853,N_24965);
and UO_1281 (O_1281,N_24987,N_24821);
or UO_1282 (O_1282,N_24895,N_24938);
nor UO_1283 (O_1283,N_24816,N_24822);
or UO_1284 (O_1284,N_24915,N_24882);
and UO_1285 (O_1285,N_24817,N_24824);
or UO_1286 (O_1286,N_24840,N_24906);
nor UO_1287 (O_1287,N_24764,N_24754);
and UO_1288 (O_1288,N_24881,N_24812);
or UO_1289 (O_1289,N_24799,N_24764);
xor UO_1290 (O_1290,N_24864,N_24795);
nor UO_1291 (O_1291,N_24776,N_24944);
xor UO_1292 (O_1292,N_24943,N_24762);
xor UO_1293 (O_1293,N_24755,N_24903);
nor UO_1294 (O_1294,N_24796,N_24781);
nand UO_1295 (O_1295,N_24940,N_24815);
nand UO_1296 (O_1296,N_24787,N_24999);
or UO_1297 (O_1297,N_24920,N_24811);
nor UO_1298 (O_1298,N_24792,N_24765);
or UO_1299 (O_1299,N_24864,N_24904);
and UO_1300 (O_1300,N_24831,N_24993);
and UO_1301 (O_1301,N_24857,N_24844);
and UO_1302 (O_1302,N_24945,N_24956);
nand UO_1303 (O_1303,N_24942,N_24955);
nand UO_1304 (O_1304,N_24883,N_24896);
nand UO_1305 (O_1305,N_24926,N_24855);
xor UO_1306 (O_1306,N_24959,N_24829);
xor UO_1307 (O_1307,N_24890,N_24928);
or UO_1308 (O_1308,N_24840,N_24954);
or UO_1309 (O_1309,N_24967,N_24893);
or UO_1310 (O_1310,N_24763,N_24882);
xor UO_1311 (O_1311,N_24841,N_24832);
or UO_1312 (O_1312,N_24975,N_24827);
and UO_1313 (O_1313,N_24899,N_24803);
or UO_1314 (O_1314,N_24854,N_24827);
xnor UO_1315 (O_1315,N_24960,N_24890);
xor UO_1316 (O_1316,N_24804,N_24967);
and UO_1317 (O_1317,N_24969,N_24789);
nand UO_1318 (O_1318,N_24839,N_24797);
and UO_1319 (O_1319,N_24956,N_24851);
nor UO_1320 (O_1320,N_24838,N_24903);
nor UO_1321 (O_1321,N_24806,N_24868);
or UO_1322 (O_1322,N_24930,N_24815);
and UO_1323 (O_1323,N_24923,N_24829);
nand UO_1324 (O_1324,N_24857,N_24821);
nor UO_1325 (O_1325,N_24795,N_24987);
xnor UO_1326 (O_1326,N_24958,N_24916);
and UO_1327 (O_1327,N_24864,N_24935);
and UO_1328 (O_1328,N_24845,N_24854);
xor UO_1329 (O_1329,N_24972,N_24821);
or UO_1330 (O_1330,N_24812,N_24920);
or UO_1331 (O_1331,N_24896,N_24934);
nand UO_1332 (O_1332,N_24947,N_24976);
xnor UO_1333 (O_1333,N_24855,N_24904);
nand UO_1334 (O_1334,N_24782,N_24772);
and UO_1335 (O_1335,N_24839,N_24961);
xnor UO_1336 (O_1336,N_24947,N_24869);
nand UO_1337 (O_1337,N_24896,N_24895);
nand UO_1338 (O_1338,N_24974,N_24955);
nor UO_1339 (O_1339,N_24997,N_24916);
nand UO_1340 (O_1340,N_24754,N_24866);
or UO_1341 (O_1341,N_24964,N_24750);
and UO_1342 (O_1342,N_24926,N_24944);
or UO_1343 (O_1343,N_24798,N_24844);
and UO_1344 (O_1344,N_24809,N_24822);
or UO_1345 (O_1345,N_24816,N_24767);
or UO_1346 (O_1346,N_24901,N_24966);
and UO_1347 (O_1347,N_24815,N_24877);
xor UO_1348 (O_1348,N_24892,N_24946);
nand UO_1349 (O_1349,N_24827,N_24837);
nand UO_1350 (O_1350,N_24828,N_24922);
or UO_1351 (O_1351,N_24837,N_24806);
or UO_1352 (O_1352,N_24955,N_24787);
xnor UO_1353 (O_1353,N_24908,N_24890);
nor UO_1354 (O_1354,N_24873,N_24922);
xnor UO_1355 (O_1355,N_24968,N_24787);
xnor UO_1356 (O_1356,N_24835,N_24837);
nor UO_1357 (O_1357,N_24967,N_24957);
or UO_1358 (O_1358,N_24862,N_24832);
nor UO_1359 (O_1359,N_24932,N_24962);
and UO_1360 (O_1360,N_24908,N_24917);
nor UO_1361 (O_1361,N_24831,N_24940);
or UO_1362 (O_1362,N_24962,N_24953);
and UO_1363 (O_1363,N_24891,N_24984);
or UO_1364 (O_1364,N_24947,N_24755);
xor UO_1365 (O_1365,N_24932,N_24998);
or UO_1366 (O_1366,N_24772,N_24854);
or UO_1367 (O_1367,N_24928,N_24889);
and UO_1368 (O_1368,N_24894,N_24804);
or UO_1369 (O_1369,N_24941,N_24827);
or UO_1370 (O_1370,N_24852,N_24770);
or UO_1371 (O_1371,N_24752,N_24854);
xor UO_1372 (O_1372,N_24881,N_24802);
nand UO_1373 (O_1373,N_24894,N_24883);
and UO_1374 (O_1374,N_24871,N_24954);
and UO_1375 (O_1375,N_24871,N_24763);
xnor UO_1376 (O_1376,N_24856,N_24835);
nand UO_1377 (O_1377,N_24900,N_24978);
nand UO_1378 (O_1378,N_24993,N_24956);
and UO_1379 (O_1379,N_24861,N_24972);
xor UO_1380 (O_1380,N_24987,N_24932);
nor UO_1381 (O_1381,N_24999,N_24940);
or UO_1382 (O_1382,N_24902,N_24974);
and UO_1383 (O_1383,N_24971,N_24838);
nand UO_1384 (O_1384,N_24904,N_24995);
and UO_1385 (O_1385,N_24792,N_24832);
and UO_1386 (O_1386,N_24879,N_24931);
nand UO_1387 (O_1387,N_24903,N_24931);
and UO_1388 (O_1388,N_24979,N_24944);
and UO_1389 (O_1389,N_24863,N_24821);
xnor UO_1390 (O_1390,N_24877,N_24874);
nor UO_1391 (O_1391,N_24963,N_24898);
and UO_1392 (O_1392,N_24756,N_24792);
xor UO_1393 (O_1393,N_24812,N_24907);
xor UO_1394 (O_1394,N_24903,N_24772);
nand UO_1395 (O_1395,N_24807,N_24753);
and UO_1396 (O_1396,N_24875,N_24783);
or UO_1397 (O_1397,N_24831,N_24800);
xor UO_1398 (O_1398,N_24835,N_24776);
xnor UO_1399 (O_1399,N_24859,N_24916);
and UO_1400 (O_1400,N_24752,N_24876);
xor UO_1401 (O_1401,N_24795,N_24908);
or UO_1402 (O_1402,N_24935,N_24938);
or UO_1403 (O_1403,N_24790,N_24812);
nor UO_1404 (O_1404,N_24832,N_24859);
or UO_1405 (O_1405,N_24768,N_24856);
nand UO_1406 (O_1406,N_24826,N_24865);
and UO_1407 (O_1407,N_24985,N_24983);
and UO_1408 (O_1408,N_24859,N_24986);
nor UO_1409 (O_1409,N_24867,N_24929);
xor UO_1410 (O_1410,N_24887,N_24777);
or UO_1411 (O_1411,N_24898,N_24895);
or UO_1412 (O_1412,N_24804,N_24882);
nand UO_1413 (O_1413,N_24973,N_24780);
nor UO_1414 (O_1414,N_24830,N_24793);
xnor UO_1415 (O_1415,N_24897,N_24930);
and UO_1416 (O_1416,N_24894,N_24761);
and UO_1417 (O_1417,N_24950,N_24905);
and UO_1418 (O_1418,N_24866,N_24978);
nor UO_1419 (O_1419,N_24785,N_24842);
nand UO_1420 (O_1420,N_24872,N_24975);
nor UO_1421 (O_1421,N_24988,N_24912);
xor UO_1422 (O_1422,N_24833,N_24753);
xor UO_1423 (O_1423,N_24751,N_24932);
and UO_1424 (O_1424,N_24950,N_24974);
nor UO_1425 (O_1425,N_24802,N_24842);
nand UO_1426 (O_1426,N_24765,N_24986);
nand UO_1427 (O_1427,N_24977,N_24906);
or UO_1428 (O_1428,N_24887,N_24827);
or UO_1429 (O_1429,N_24877,N_24891);
xor UO_1430 (O_1430,N_24866,N_24893);
or UO_1431 (O_1431,N_24879,N_24894);
nand UO_1432 (O_1432,N_24874,N_24816);
nor UO_1433 (O_1433,N_24881,N_24984);
nor UO_1434 (O_1434,N_24876,N_24847);
or UO_1435 (O_1435,N_24967,N_24944);
nor UO_1436 (O_1436,N_24880,N_24994);
or UO_1437 (O_1437,N_24963,N_24755);
nor UO_1438 (O_1438,N_24783,N_24819);
nand UO_1439 (O_1439,N_24995,N_24862);
or UO_1440 (O_1440,N_24901,N_24776);
or UO_1441 (O_1441,N_24813,N_24843);
nor UO_1442 (O_1442,N_24966,N_24797);
nor UO_1443 (O_1443,N_24764,N_24866);
nor UO_1444 (O_1444,N_24973,N_24815);
nand UO_1445 (O_1445,N_24948,N_24765);
nand UO_1446 (O_1446,N_24773,N_24858);
nor UO_1447 (O_1447,N_24849,N_24982);
and UO_1448 (O_1448,N_24942,N_24946);
nor UO_1449 (O_1449,N_24903,N_24861);
xnor UO_1450 (O_1450,N_24888,N_24859);
nor UO_1451 (O_1451,N_24833,N_24876);
nand UO_1452 (O_1452,N_24845,N_24999);
or UO_1453 (O_1453,N_24787,N_24965);
or UO_1454 (O_1454,N_24952,N_24999);
nand UO_1455 (O_1455,N_24803,N_24930);
nor UO_1456 (O_1456,N_24949,N_24901);
and UO_1457 (O_1457,N_24917,N_24982);
and UO_1458 (O_1458,N_24757,N_24924);
and UO_1459 (O_1459,N_24894,N_24940);
and UO_1460 (O_1460,N_24913,N_24866);
nor UO_1461 (O_1461,N_24840,N_24900);
xor UO_1462 (O_1462,N_24910,N_24988);
and UO_1463 (O_1463,N_24974,N_24890);
xnor UO_1464 (O_1464,N_24852,N_24835);
xnor UO_1465 (O_1465,N_24820,N_24905);
nand UO_1466 (O_1466,N_24787,N_24959);
xnor UO_1467 (O_1467,N_24754,N_24792);
xnor UO_1468 (O_1468,N_24840,N_24878);
and UO_1469 (O_1469,N_24980,N_24936);
nor UO_1470 (O_1470,N_24960,N_24978);
xnor UO_1471 (O_1471,N_24910,N_24955);
or UO_1472 (O_1472,N_24864,N_24842);
or UO_1473 (O_1473,N_24959,N_24939);
or UO_1474 (O_1474,N_24780,N_24926);
or UO_1475 (O_1475,N_24937,N_24941);
and UO_1476 (O_1476,N_24865,N_24789);
nor UO_1477 (O_1477,N_24824,N_24859);
xnor UO_1478 (O_1478,N_24909,N_24961);
xor UO_1479 (O_1479,N_24764,N_24942);
and UO_1480 (O_1480,N_24868,N_24783);
xor UO_1481 (O_1481,N_24810,N_24931);
or UO_1482 (O_1482,N_24964,N_24796);
or UO_1483 (O_1483,N_24883,N_24922);
nor UO_1484 (O_1484,N_24953,N_24922);
nand UO_1485 (O_1485,N_24870,N_24917);
and UO_1486 (O_1486,N_24851,N_24997);
xor UO_1487 (O_1487,N_24902,N_24760);
xor UO_1488 (O_1488,N_24834,N_24940);
nand UO_1489 (O_1489,N_24810,N_24763);
nor UO_1490 (O_1490,N_24839,N_24826);
nand UO_1491 (O_1491,N_24945,N_24880);
nor UO_1492 (O_1492,N_24796,N_24895);
and UO_1493 (O_1493,N_24750,N_24862);
nor UO_1494 (O_1494,N_24984,N_24792);
xor UO_1495 (O_1495,N_24799,N_24856);
or UO_1496 (O_1496,N_24872,N_24846);
and UO_1497 (O_1497,N_24823,N_24991);
nor UO_1498 (O_1498,N_24942,N_24816);
and UO_1499 (O_1499,N_24943,N_24803);
xnor UO_1500 (O_1500,N_24849,N_24777);
xnor UO_1501 (O_1501,N_24953,N_24933);
xnor UO_1502 (O_1502,N_24948,N_24934);
xor UO_1503 (O_1503,N_24914,N_24753);
or UO_1504 (O_1504,N_24817,N_24889);
nor UO_1505 (O_1505,N_24907,N_24818);
xnor UO_1506 (O_1506,N_24975,N_24828);
and UO_1507 (O_1507,N_24837,N_24978);
and UO_1508 (O_1508,N_24837,N_24762);
nand UO_1509 (O_1509,N_24807,N_24869);
or UO_1510 (O_1510,N_24806,N_24871);
nand UO_1511 (O_1511,N_24839,N_24841);
nor UO_1512 (O_1512,N_24964,N_24987);
nand UO_1513 (O_1513,N_24879,N_24771);
and UO_1514 (O_1514,N_24910,N_24919);
nand UO_1515 (O_1515,N_24795,N_24962);
xor UO_1516 (O_1516,N_24762,N_24858);
nor UO_1517 (O_1517,N_24752,N_24995);
nor UO_1518 (O_1518,N_24851,N_24835);
xor UO_1519 (O_1519,N_24946,N_24856);
nand UO_1520 (O_1520,N_24825,N_24931);
or UO_1521 (O_1521,N_24912,N_24914);
xnor UO_1522 (O_1522,N_24870,N_24797);
nand UO_1523 (O_1523,N_24895,N_24937);
xor UO_1524 (O_1524,N_24878,N_24901);
xor UO_1525 (O_1525,N_24795,N_24751);
xor UO_1526 (O_1526,N_24971,N_24804);
or UO_1527 (O_1527,N_24767,N_24832);
and UO_1528 (O_1528,N_24798,N_24954);
nand UO_1529 (O_1529,N_24915,N_24992);
and UO_1530 (O_1530,N_24833,N_24937);
or UO_1531 (O_1531,N_24875,N_24893);
nand UO_1532 (O_1532,N_24915,N_24752);
nand UO_1533 (O_1533,N_24935,N_24880);
nor UO_1534 (O_1534,N_24816,N_24776);
or UO_1535 (O_1535,N_24775,N_24967);
and UO_1536 (O_1536,N_24937,N_24951);
xnor UO_1537 (O_1537,N_24809,N_24910);
nand UO_1538 (O_1538,N_24872,N_24934);
nand UO_1539 (O_1539,N_24989,N_24874);
or UO_1540 (O_1540,N_24826,N_24785);
and UO_1541 (O_1541,N_24965,N_24981);
and UO_1542 (O_1542,N_24844,N_24875);
xor UO_1543 (O_1543,N_24902,N_24985);
nor UO_1544 (O_1544,N_24956,N_24964);
nand UO_1545 (O_1545,N_24954,N_24909);
nand UO_1546 (O_1546,N_24902,N_24860);
nand UO_1547 (O_1547,N_24920,N_24821);
xor UO_1548 (O_1548,N_24794,N_24839);
and UO_1549 (O_1549,N_24884,N_24981);
or UO_1550 (O_1550,N_24853,N_24957);
or UO_1551 (O_1551,N_24992,N_24897);
nand UO_1552 (O_1552,N_24807,N_24966);
and UO_1553 (O_1553,N_24963,N_24825);
or UO_1554 (O_1554,N_24864,N_24993);
xor UO_1555 (O_1555,N_24802,N_24903);
xor UO_1556 (O_1556,N_24908,N_24997);
nor UO_1557 (O_1557,N_24946,N_24998);
nand UO_1558 (O_1558,N_24989,N_24838);
and UO_1559 (O_1559,N_24849,N_24913);
and UO_1560 (O_1560,N_24987,N_24982);
nor UO_1561 (O_1561,N_24784,N_24770);
nor UO_1562 (O_1562,N_24903,N_24928);
xnor UO_1563 (O_1563,N_24978,N_24783);
or UO_1564 (O_1564,N_24931,N_24862);
nor UO_1565 (O_1565,N_24854,N_24849);
xnor UO_1566 (O_1566,N_24803,N_24901);
or UO_1567 (O_1567,N_24910,N_24944);
or UO_1568 (O_1568,N_24950,N_24965);
nand UO_1569 (O_1569,N_24934,N_24756);
nand UO_1570 (O_1570,N_24874,N_24841);
or UO_1571 (O_1571,N_24883,N_24768);
and UO_1572 (O_1572,N_24762,N_24776);
and UO_1573 (O_1573,N_24811,N_24868);
nor UO_1574 (O_1574,N_24944,N_24919);
nor UO_1575 (O_1575,N_24884,N_24827);
nand UO_1576 (O_1576,N_24796,N_24920);
and UO_1577 (O_1577,N_24898,N_24985);
or UO_1578 (O_1578,N_24910,N_24868);
nand UO_1579 (O_1579,N_24787,N_24778);
nor UO_1580 (O_1580,N_24920,N_24829);
nor UO_1581 (O_1581,N_24846,N_24858);
nand UO_1582 (O_1582,N_24991,N_24974);
xnor UO_1583 (O_1583,N_24793,N_24941);
and UO_1584 (O_1584,N_24932,N_24758);
xor UO_1585 (O_1585,N_24941,N_24764);
xnor UO_1586 (O_1586,N_24879,N_24925);
or UO_1587 (O_1587,N_24965,N_24756);
xnor UO_1588 (O_1588,N_24811,N_24939);
nand UO_1589 (O_1589,N_24837,N_24841);
xor UO_1590 (O_1590,N_24998,N_24879);
nand UO_1591 (O_1591,N_24892,N_24820);
nor UO_1592 (O_1592,N_24858,N_24866);
xor UO_1593 (O_1593,N_24831,N_24830);
nand UO_1594 (O_1594,N_24872,N_24902);
nand UO_1595 (O_1595,N_24915,N_24938);
and UO_1596 (O_1596,N_24918,N_24981);
xor UO_1597 (O_1597,N_24826,N_24792);
nand UO_1598 (O_1598,N_24777,N_24939);
or UO_1599 (O_1599,N_24904,N_24903);
nand UO_1600 (O_1600,N_24872,N_24896);
or UO_1601 (O_1601,N_24823,N_24920);
nor UO_1602 (O_1602,N_24853,N_24898);
or UO_1603 (O_1603,N_24781,N_24950);
or UO_1604 (O_1604,N_24961,N_24897);
nand UO_1605 (O_1605,N_24791,N_24948);
nor UO_1606 (O_1606,N_24926,N_24810);
xor UO_1607 (O_1607,N_24886,N_24927);
nand UO_1608 (O_1608,N_24899,N_24998);
and UO_1609 (O_1609,N_24989,N_24771);
xor UO_1610 (O_1610,N_24860,N_24825);
nand UO_1611 (O_1611,N_24755,N_24898);
or UO_1612 (O_1612,N_24918,N_24992);
nor UO_1613 (O_1613,N_24807,N_24792);
nor UO_1614 (O_1614,N_24965,N_24765);
nand UO_1615 (O_1615,N_24766,N_24993);
and UO_1616 (O_1616,N_24756,N_24887);
and UO_1617 (O_1617,N_24787,N_24793);
xor UO_1618 (O_1618,N_24771,N_24899);
and UO_1619 (O_1619,N_24977,N_24891);
nand UO_1620 (O_1620,N_24899,N_24933);
xnor UO_1621 (O_1621,N_24864,N_24845);
nor UO_1622 (O_1622,N_24931,N_24968);
nand UO_1623 (O_1623,N_24754,N_24807);
and UO_1624 (O_1624,N_24919,N_24939);
xor UO_1625 (O_1625,N_24759,N_24771);
xnor UO_1626 (O_1626,N_24771,N_24821);
and UO_1627 (O_1627,N_24959,N_24786);
xor UO_1628 (O_1628,N_24900,N_24885);
or UO_1629 (O_1629,N_24780,N_24792);
nor UO_1630 (O_1630,N_24770,N_24825);
and UO_1631 (O_1631,N_24810,N_24941);
xor UO_1632 (O_1632,N_24795,N_24775);
nor UO_1633 (O_1633,N_24775,N_24784);
or UO_1634 (O_1634,N_24937,N_24768);
nor UO_1635 (O_1635,N_24835,N_24780);
nand UO_1636 (O_1636,N_24948,N_24775);
xor UO_1637 (O_1637,N_24960,N_24767);
xnor UO_1638 (O_1638,N_24801,N_24798);
and UO_1639 (O_1639,N_24790,N_24786);
nor UO_1640 (O_1640,N_24969,N_24885);
xor UO_1641 (O_1641,N_24831,N_24818);
or UO_1642 (O_1642,N_24921,N_24956);
nor UO_1643 (O_1643,N_24756,N_24856);
or UO_1644 (O_1644,N_24788,N_24855);
or UO_1645 (O_1645,N_24981,N_24832);
nor UO_1646 (O_1646,N_24988,N_24992);
xnor UO_1647 (O_1647,N_24961,N_24932);
nor UO_1648 (O_1648,N_24823,N_24824);
nand UO_1649 (O_1649,N_24965,N_24804);
xnor UO_1650 (O_1650,N_24780,N_24995);
nor UO_1651 (O_1651,N_24864,N_24810);
xnor UO_1652 (O_1652,N_24954,N_24841);
nand UO_1653 (O_1653,N_24818,N_24766);
nor UO_1654 (O_1654,N_24947,N_24859);
and UO_1655 (O_1655,N_24882,N_24819);
and UO_1656 (O_1656,N_24944,N_24806);
nand UO_1657 (O_1657,N_24912,N_24975);
or UO_1658 (O_1658,N_24945,N_24946);
nand UO_1659 (O_1659,N_24833,N_24838);
nor UO_1660 (O_1660,N_24791,N_24994);
xor UO_1661 (O_1661,N_24949,N_24863);
xnor UO_1662 (O_1662,N_24875,N_24753);
nor UO_1663 (O_1663,N_24979,N_24869);
nor UO_1664 (O_1664,N_24813,N_24808);
nand UO_1665 (O_1665,N_24826,N_24830);
and UO_1666 (O_1666,N_24905,N_24908);
nor UO_1667 (O_1667,N_24816,N_24847);
xor UO_1668 (O_1668,N_24797,N_24983);
and UO_1669 (O_1669,N_24950,N_24886);
nor UO_1670 (O_1670,N_24769,N_24911);
and UO_1671 (O_1671,N_24905,N_24839);
nor UO_1672 (O_1672,N_24890,N_24769);
and UO_1673 (O_1673,N_24995,N_24960);
xnor UO_1674 (O_1674,N_24900,N_24875);
xor UO_1675 (O_1675,N_24993,N_24775);
xnor UO_1676 (O_1676,N_24917,N_24788);
nand UO_1677 (O_1677,N_24802,N_24954);
nand UO_1678 (O_1678,N_24940,N_24950);
nor UO_1679 (O_1679,N_24840,N_24806);
nand UO_1680 (O_1680,N_24974,N_24751);
or UO_1681 (O_1681,N_24789,N_24771);
nor UO_1682 (O_1682,N_24840,N_24957);
nor UO_1683 (O_1683,N_24854,N_24776);
nand UO_1684 (O_1684,N_24765,N_24806);
and UO_1685 (O_1685,N_24944,N_24843);
or UO_1686 (O_1686,N_24912,N_24924);
nor UO_1687 (O_1687,N_24872,N_24772);
and UO_1688 (O_1688,N_24769,N_24859);
xnor UO_1689 (O_1689,N_24935,N_24752);
xor UO_1690 (O_1690,N_24978,N_24785);
nor UO_1691 (O_1691,N_24773,N_24866);
nand UO_1692 (O_1692,N_24915,N_24761);
nor UO_1693 (O_1693,N_24872,N_24978);
nor UO_1694 (O_1694,N_24914,N_24830);
or UO_1695 (O_1695,N_24915,N_24997);
nand UO_1696 (O_1696,N_24977,N_24762);
or UO_1697 (O_1697,N_24994,N_24941);
xor UO_1698 (O_1698,N_24902,N_24999);
xor UO_1699 (O_1699,N_24810,N_24846);
nand UO_1700 (O_1700,N_24883,N_24970);
nand UO_1701 (O_1701,N_24787,N_24911);
and UO_1702 (O_1702,N_24753,N_24922);
xnor UO_1703 (O_1703,N_24991,N_24772);
or UO_1704 (O_1704,N_24940,N_24901);
nor UO_1705 (O_1705,N_24924,N_24859);
nand UO_1706 (O_1706,N_24852,N_24789);
nand UO_1707 (O_1707,N_24852,N_24893);
nor UO_1708 (O_1708,N_24786,N_24899);
and UO_1709 (O_1709,N_24786,N_24843);
and UO_1710 (O_1710,N_24825,N_24756);
nor UO_1711 (O_1711,N_24799,N_24908);
and UO_1712 (O_1712,N_24892,N_24798);
or UO_1713 (O_1713,N_24967,N_24787);
and UO_1714 (O_1714,N_24888,N_24857);
and UO_1715 (O_1715,N_24778,N_24943);
or UO_1716 (O_1716,N_24968,N_24758);
nand UO_1717 (O_1717,N_24998,N_24939);
nand UO_1718 (O_1718,N_24988,N_24847);
and UO_1719 (O_1719,N_24858,N_24964);
or UO_1720 (O_1720,N_24948,N_24864);
nor UO_1721 (O_1721,N_24887,N_24951);
and UO_1722 (O_1722,N_24812,N_24801);
nand UO_1723 (O_1723,N_24799,N_24947);
nand UO_1724 (O_1724,N_24993,N_24991);
and UO_1725 (O_1725,N_24870,N_24936);
and UO_1726 (O_1726,N_24868,N_24987);
nor UO_1727 (O_1727,N_24825,N_24855);
nor UO_1728 (O_1728,N_24940,N_24977);
nand UO_1729 (O_1729,N_24933,N_24875);
nor UO_1730 (O_1730,N_24884,N_24906);
nor UO_1731 (O_1731,N_24906,N_24992);
or UO_1732 (O_1732,N_24918,N_24835);
nor UO_1733 (O_1733,N_24971,N_24823);
xor UO_1734 (O_1734,N_24955,N_24860);
or UO_1735 (O_1735,N_24980,N_24902);
xor UO_1736 (O_1736,N_24846,N_24868);
or UO_1737 (O_1737,N_24939,N_24833);
nand UO_1738 (O_1738,N_24779,N_24876);
or UO_1739 (O_1739,N_24872,N_24919);
and UO_1740 (O_1740,N_24892,N_24948);
and UO_1741 (O_1741,N_24842,N_24776);
and UO_1742 (O_1742,N_24965,N_24753);
nand UO_1743 (O_1743,N_24865,N_24828);
nor UO_1744 (O_1744,N_24843,N_24776);
nand UO_1745 (O_1745,N_24790,N_24817);
nor UO_1746 (O_1746,N_24829,N_24905);
or UO_1747 (O_1747,N_24969,N_24780);
xor UO_1748 (O_1748,N_24976,N_24836);
and UO_1749 (O_1749,N_24803,N_24775);
and UO_1750 (O_1750,N_24936,N_24772);
or UO_1751 (O_1751,N_24799,N_24841);
or UO_1752 (O_1752,N_24913,N_24779);
nand UO_1753 (O_1753,N_24784,N_24898);
and UO_1754 (O_1754,N_24803,N_24860);
xnor UO_1755 (O_1755,N_24840,N_24949);
or UO_1756 (O_1756,N_24784,N_24948);
xor UO_1757 (O_1757,N_24794,N_24826);
and UO_1758 (O_1758,N_24912,N_24995);
nand UO_1759 (O_1759,N_24799,N_24941);
and UO_1760 (O_1760,N_24907,N_24837);
xor UO_1761 (O_1761,N_24804,N_24773);
or UO_1762 (O_1762,N_24964,N_24760);
nor UO_1763 (O_1763,N_24872,N_24917);
xor UO_1764 (O_1764,N_24985,N_24853);
and UO_1765 (O_1765,N_24829,N_24976);
xor UO_1766 (O_1766,N_24795,N_24849);
xnor UO_1767 (O_1767,N_24962,N_24992);
nand UO_1768 (O_1768,N_24923,N_24889);
nor UO_1769 (O_1769,N_24787,N_24760);
or UO_1770 (O_1770,N_24935,N_24827);
nor UO_1771 (O_1771,N_24982,N_24894);
or UO_1772 (O_1772,N_24976,N_24782);
nor UO_1773 (O_1773,N_24969,N_24766);
and UO_1774 (O_1774,N_24757,N_24968);
xnor UO_1775 (O_1775,N_24989,N_24834);
xor UO_1776 (O_1776,N_24903,N_24805);
and UO_1777 (O_1777,N_24778,N_24789);
nand UO_1778 (O_1778,N_24986,N_24931);
and UO_1779 (O_1779,N_24853,N_24904);
or UO_1780 (O_1780,N_24751,N_24996);
or UO_1781 (O_1781,N_24754,N_24935);
and UO_1782 (O_1782,N_24932,N_24805);
xor UO_1783 (O_1783,N_24824,N_24940);
nor UO_1784 (O_1784,N_24978,N_24995);
nand UO_1785 (O_1785,N_24827,N_24959);
and UO_1786 (O_1786,N_24935,N_24823);
xnor UO_1787 (O_1787,N_24819,N_24775);
and UO_1788 (O_1788,N_24860,N_24899);
nand UO_1789 (O_1789,N_24843,N_24879);
or UO_1790 (O_1790,N_24951,N_24808);
or UO_1791 (O_1791,N_24875,N_24956);
or UO_1792 (O_1792,N_24768,N_24939);
xor UO_1793 (O_1793,N_24750,N_24972);
nand UO_1794 (O_1794,N_24885,N_24793);
xnor UO_1795 (O_1795,N_24869,N_24898);
or UO_1796 (O_1796,N_24933,N_24932);
and UO_1797 (O_1797,N_24815,N_24843);
and UO_1798 (O_1798,N_24982,N_24755);
and UO_1799 (O_1799,N_24953,N_24834);
and UO_1800 (O_1800,N_24976,N_24901);
and UO_1801 (O_1801,N_24785,N_24816);
and UO_1802 (O_1802,N_24906,N_24851);
nand UO_1803 (O_1803,N_24889,N_24792);
xor UO_1804 (O_1804,N_24834,N_24808);
xnor UO_1805 (O_1805,N_24959,N_24790);
or UO_1806 (O_1806,N_24912,N_24908);
or UO_1807 (O_1807,N_24930,N_24989);
nor UO_1808 (O_1808,N_24848,N_24893);
xor UO_1809 (O_1809,N_24799,N_24806);
or UO_1810 (O_1810,N_24869,N_24954);
and UO_1811 (O_1811,N_24847,N_24796);
and UO_1812 (O_1812,N_24951,N_24933);
nor UO_1813 (O_1813,N_24925,N_24839);
or UO_1814 (O_1814,N_24952,N_24847);
and UO_1815 (O_1815,N_24762,N_24851);
nor UO_1816 (O_1816,N_24991,N_24846);
and UO_1817 (O_1817,N_24895,N_24830);
nor UO_1818 (O_1818,N_24829,N_24981);
or UO_1819 (O_1819,N_24835,N_24762);
or UO_1820 (O_1820,N_24828,N_24945);
nor UO_1821 (O_1821,N_24876,N_24848);
xnor UO_1822 (O_1822,N_24846,N_24758);
or UO_1823 (O_1823,N_24908,N_24779);
nand UO_1824 (O_1824,N_24977,N_24910);
xnor UO_1825 (O_1825,N_24833,N_24806);
and UO_1826 (O_1826,N_24971,N_24975);
and UO_1827 (O_1827,N_24921,N_24852);
nand UO_1828 (O_1828,N_24792,N_24815);
xnor UO_1829 (O_1829,N_24798,N_24975);
and UO_1830 (O_1830,N_24962,N_24971);
or UO_1831 (O_1831,N_24857,N_24957);
or UO_1832 (O_1832,N_24904,N_24949);
nand UO_1833 (O_1833,N_24986,N_24874);
xor UO_1834 (O_1834,N_24755,N_24981);
and UO_1835 (O_1835,N_24754,N_24923);
and UO_1836 (O_1836,N_24930,N_24952);
xnor UO_1837 (O_1837,N_24955,N_24935);
nor UO_1838 (O_1838,N_24895,N_24763);
xnor UO_1839 (O_1839,N_24809,N_24898);
and UO_1840 (O_1840,N_24755,N_24955);
and UO_1841 (O_1841,N_24755,N_24911);
or UO_1842 (O_1842,N_24769,N_24836);
nand UO_1843 (O_1843,N_24989,N_24794);
and UO_1844 (O_1844,N_24755,N_24980);
xor UO_1845 (O_1845,N_24981,N_24949);
nand UO_1846 (O_1846,N_24863,N_24779);
and UO_1847 (O_1847,N_24834,N_24991);
nor UO_1848 (O_1848,N_24964,N_24872);
nor UO_1849 (O_1849,N_24885,N_24916);
xor UO_1850 (O_1850,N_24896,N_24878);
and UO_1851 (O_1851,N_24996,N_24876);
or UO_1852 (O_1852,N_24870,N_24924);
nor UO_1853 (O_1853,N_24764,N_24826);
xnor UO_1854 (O_1854,N_24985,N_24756);
xnor UO_1855 (O_1855,N_24977,N_24990);
nand UO_1856 (O_1856,N_24830,N_24945);
nand UO_1857 (O_1857,N_24752,N_24785);
and UO_1858 (O_1858,N_24963,N_24989);
nand UO_1859 (O_1859,N_24853,N_24996);
xor UO_1860 (O_1860,N_24773,N_24883);
nor UO_1861 (O_1861,N_24826,N_24809);
and UO_1862 (O_1862,N_24954,N_24982);
xnor UO_1863 (O_1863,N_24940,N_24822);
nand UO_1864 (O_1864,N_24855,N_24846);
nand UO_1865 (O_1865,N_24915,N_24988);
and UO_1866 (O_1866,N_24913,N_24823);
nand UO_1867 (O_1867,N_24755,N_24973);
nand UO_1868 (O_1868,N_24902,N_24837);
nand UO_1869 (O_1869,N_24933,N_24818);
nor UO_1870 (O_1870,N_24750,N_24955);
and UO_1871 (O_1871,N_24753,N_24762);
nand UO_1872 (O_1872,N_24805,N_24995);
nand UO_1873 (O_1873,N_24819,N_24779);
nand UO_1874 (O_1874,N_24878,N_24937);
and UO_1875 (O_1875,N_24760,N_24848);
or UO_1876 (O_1876,N_24830,N_24974);
nand UO_1877 (O_1877,N_24985,N_24850);
or UO_1878 (O_1878,N_24936,N_24837);
nor UO_1879 (O_1879,N_24821,N_24817);
xnor UO_1880 (O_1880,N_24892,N_24860);
xnor UO_1881 (O_1881,N_24779,N_24955);
and UO_1882 (O_1882,N_24955,N_24871);
or UO_1883 (O_1883,N_24975,N_24916);
and UO_1884 (O_1884,N_24751,N_24980);
and UO_1885 (O_1885,N_24843,N_24873);
xnor UO_1886 (O_1886,N_24845,N_24915);
or UO_1887 (O_1887,N_24770,N_24757);
nand UO_1888 (O_1888,N_24875,N_24841);
and UO_1889 (O_1889,N_24890,N_24969);
and UO_1890 (O_1890,N_24929,N_24895);
nand UO_1891 (O_1891,N_24826,N_24772);
nor UO_1892 (O_1892,N_24967,N_24852);
nand UO_1893 (O_1893,N_24947,N_24844);
nor UO_1894 (O_1894,N_24756,N_24806);
xnor UO_1895 (O_1895,N_24781,N_24887);
and UO_1896 (O_1896,N_24903,N_24801);
xnor UO_1897 (O_1897,N_24806,N_24875);
nand UO_1898 (O_1898,N_24960,N_24930);
or UO_1899 (O_1899,N_24754,N_24994);
or UO_1900 (O_1900,N_24863,N_24780);
xor UO_1901 (O_1901,N_24944,N_24861);
xor UO_1902 (O_1902,N_24760,N_24762);
xnor UO_1903 (O_1903,N_24877,N_24966);
and UO_1904 (O_1904,N_24771,N_24977);
nand UO_1905 (O_1905,N_24814,N_24940);
and UO_1906 (O_1906,N_24947,N_24893);
nand UO_1907 (O_1907,N_24812,N_24770);
or UO_1908 (O_1908,N_24896,N_24780);
nand UO_1909 (O_1909,N_24942,N_24752);
and UO_1910 (O_1910,N_24976,N_24772);
or UO_1911 (O_1911,N_24856,N_24842);
nand UO_1912 (O_1912,N_24860,N_24814);
nor UO_1913 (O_1913,N_24852,N_24825);
nand UO_1914 (O_1914,N_24797,N_24877);
nor UO_1915 (O_1915,N_24777,N_24967);
xor UO_1916 (O_1916,N_24943,N_24890);
and UO_1917 (O_1917,N_24798,N_24845);
nor UO_1918 (O_1918,N_24839,N_24888);
nor UO_1919 (O_1919,N_24910,N_24766);
and UO_1920 (O_1920,N_24888,N_24984);
xnor UO_1921 (O_1921,N_24992,N_24972);
and UO_1922 (O_1922,N_24800,N_24845);
or UO_1923 (O_1923,N_24939,N_24954);
or UO_1924 (O_1924,N_24928,N_24885);
or UO_1925 (O_1925,N_24941,N_24754);
nand UO_1926 (O_1926,N_24920,N_24846);
nor UO_1927 (O_1927,N_24981,N_24888);
xor UO_1928 (O_1928,N_24759,N_24875);
nor UO_1929 (O_1929,N_24832,N_24800);
xnor UO_1930 (O_1930,N_24922,N_24933);
and UO_1931 (O_1931,N_24761,N_24802);
and UO_1932 (O_1932,N_24889,N_24777);
xnor UO_1933 (O_1933,N_24812,N_24906);
nand UO_1934 (O_1934,N_24801,N_24867);
nor UO_1935 (O_1935,N_24923,N_24917);
or UO_1936 (O_1936,N_24853,N_24942);
xor UO_1937 (O_1937,N_24901,N_24791);
or UO_1938 (O_1938,N_24850,N_24757);
nand UO_1939 (O_1939,N_24988,N_24769);
or UO_1940 (O_1940,N_24915,N_24890);
and UO_1941 (O_1941,N_24767,N_24910);
nand UO_1942 (O_1942,N_24767,N_24967);
xor UO_1943 (O_1943,N_24825,N_24895);
and UO_1944 (O_1944,N_24978,N_24997);
nor UO_1945 (O_1945,N_24856,N_24969);
nand UO_1946 (O_1946,N_24805,N_24781);
and UO_1947 (O_1947,N_24912,N_24761);
nand UO_1948 (O_1948,N_24856,N_24932);
and UO_1949 (O_1949,N_24938,N_24754);
nor UO_1950 (O_1950,N_24942,N_24907);
or UO_1951 (O_1951,N_24891,N_24943);
xor UO_1952 (O_1952,N_24798,N_24829);
or UO_1953 (O_1953,N_24920,N_24817);
nor UO_1954 (O_1954,N_24848,N_24818);
or UO_1955 (O_1955,N_24940,N_24918);
or UO_1956 (O_1956,N_24819,N_24802);
xnor UO_1957 (O_1957,N_24884,N_24940);
xnor UO_1958 (O_1958,N_24991,N_24882);
and UO_1959 (O_1959,N_24883,N_24853);
nor UO_1960 (O_1960,N_24824,N_24899);
or UO_1961 (O_1961,N_24799,N_24934);
and UO_1962 (O_1962,N_24939,N_24935);
xnor UO_1963 (O_1963,N_24872,N_24761);
or UO_1964 (O_1964,N_24859,N_24836);
and UO_1965 (O_1965,N_24760,N_24978);
nor UO_1966 (O_1966,N_24923,N_24757);
nor UO_1967 (O_1967,N_24857,N_24909);
nand UO_1968 (O_1968,N_24942,N_24848);
nand UO_1969 (O_1969,N_24863,N_24875);
and UO_1970 (O_1970,N_24947,N_24842);
or UO_1971 (O_1971,N_24819,N_24847);
xnor UO_1972 (O_1972,N_24979,N_24942);
or UO_1973 (O_1973,N_24972,N_24762);
nand UO_1974 (O_1974,N_24950,N_24876);
nor UO_1975 (O_1975,N_24913,N_24954);
or UO_1976 (O_1976,N_24971,N_24813);
xnor UO_1977 (O_1977,N_24908,N_24773);
xnor UO_1978 (O_1978,N_24980,N_24877);
nor UO_1979 (O_1979,N_24857,N_24797);
and UO_1980 (O_1980,N_24794,N_24779);
nand UO_1981 (O_1981,N_24884,N_24855);
or UO_1982 (O_1982,N_24828,N_24909);
nand UO_1983 (O_1983,N_24964,N_24877);
nand UO_1984 (O_1984,N_24901,N_24956);
nor UO_1985 (O_1985,N_24754,N_24815);
nand UO_1986 (O_1986,N_24953,N_24934);
or UO_1987 (O_1987,N_24915,N_24880);
nand UO_1988 (O_1988,N_24904,N_24876);
or UO_1989 (O_1989,N_24952,N_24951);
nand UO_1990 (O_1990,N_24877,N_24887);
xnor UO_1991 (O_1991,N_24908,N_24852);
or UO_1992 (O_1992,N_24853,N_24928);
or UO_1993 (O_1993,N_24804,N_24822);
and UO_1994 (O_1994,N_24799,N_24811);
and UO_1995 (O_1995,N_24850,N_24772);
nor UO_1996 (O_1996,N_24832,N_24906);
and UO_1997 (O_1997,N_24803,N_24964);
and UO_1998 (O_1998,N_24935,N_24912);
nand UO_1999 (O_1999,N_24784,N_24766);
xor UO_2000 (O_2000,N_24936,N_24795);
or UO_2001 (O_2001,N_24983,N_24789);
nor UO_2002 (O_2002,N_24853,N_24961);
nand UO_2003 (O_2003,N_24823,N_24993);
nand UO_2004 (O_2004,N_24836,N_24877);
nor UO_2005 (O_2005,N_24783,N_24820);
nor UO_2006 (O_2006,N_24923,N_24879);
or UO_2007 (O_2007,N_24871,N_24890);
and UO_2008 (O_2008,N_24997,N_24856);
nand UO_2009 (O_2009,N_24778,N_24751);
xor UO_2010 (O_2010,N_24811,N_24869);
nor UO_2011 (O_2011,N_24876,N_24759);
xor UO_2012 (O_2012,N_24966,N_24929);
and UO_2013 (O_2013,N_24926,N_24888);
xnor UO_2014 (O_2014,N_24798,N_24851);
nor UO_2015 (O_2015,N_24761,N_24774);
nand UO_2016 (O_2016,N_24982,N_24864);
xnor UO_2017 (O_2017,N_24856,N_24880);
or UO_2018 (O_2018,N_24753,N_24978);
and UO_2019 (O_2019,N_24820,N_24904);
xnor UO_2020 (O_2020,N_24967,N_24909);
and UO_2021 (O_2021,N_24855,N_24843);
xor UO_2022 (O_2022,N_24752,N_24870);
nand UO_2023 (O_2023,N_24886,N_24961);
nand UO_2024 (O_2024,N_24949,N_24963);
nor UO_2025 (O_2025,N_24889,N_24778);
nor UO_2026 (O_2026,N_24802,N_24838);
nand UO_2027 (O_2027,N_24866,N_24832);
and UO_2028 (O_2028,N_24895,N_24880);
nor UO_2029 (O_2029,N_24753,N_24894);
and UO_2030 (O_2030,N_24790,N_24798);
nor UO_2031 (O_2031,N_24961,N_24872);
and UO_2032 (O_2032,N_24975,N_24943);
or UO_2033 (O_2033,N_24891,N_24789);
nor UO_2034 (O_2034,N_24807,N_24871);
nand UO_2035 (O_2035,N_24832,N_24953);
nor UO_2036 (O_2036,N_24856,N_24765);
or UO_2037 (O_2037,N_24828,N_24861);
or UO_2038 (O_2038,N_24960,N_24758);
or UO_2039 (O_2039,N_24808,N_24980);
or UO_2040 (O_2040,N_24753,N_24867);
nor UO_2041 (O_2041,N_24832,N_24937);
xnor UO_2042 (O_2042,N_24761,N_24909);
xor UO_2043 (O_2043,N_24869,N_24787);
or UO_2044 (O_2044,N_24756,N_24890);
xnor UO_2045 (O_2045,N_24964,N_24843);
or UO_2046 (O_2046,N_24971,N_24911);
nor UO_2047 (O_2047,N_24831,N_24935);
nand UO_2048 (O_2048,N_24818,N_24794);
nand UO_2049 (O_2049,N_24775,N_24900);
or UO_2050 (O_2050,N_24924,N_24972);
or UO_2051 (O_2051,N_24883,N_24931);
or UO_2052 (O_2052,N_24850,N_24871);
and UO_2053 (O_2053,N_24823,N_24822);
nor UO_2054 (O_2054,N_24821,N_24754);
xor UO_2055 (O_2055,N_24927,N_24921);
nor UO_2056 (O_2056,N_24851,N_24875);
nor UO_2057 (O_2057,N_24969,N_24819);
and UO_2058 (O_2058,N_24989,N_24995);
nand UO_2059 (O_2059,N_24952,N_24972);
and UO_2060 (O_2060,N_24978,N_24877);
and UO_2061 (O_2061,N_24767,N_24841);
or UO_2062 (O_2062,N_24903,N_24783);
xor UO_2063 (O_2063,N_24861,N_24842);
and UO_2064 (O_2064,N_24870,N_24795);
and UO_2065 (O_2065,N_24758,N_24841);
and UO_2066 (O_2066,N_24805,N_24813);
nand UO_2067 (O_2067,N_24944,N_24931);
nor UO_2068 (O_2068,N_24782,N_24810);
and UO_2069 (O_2069,N_24904,N_24830);
nand UO_2070 (O_2070,N_24809,N_24751);
nand UO_2071 (O_2071,N_24904,N_24810);
and UO_2072 (O_2072,N_24751,N_24987);
nand UO_2073 (O_2073,N_24939,N_24875);
xor UO_2074 (O_2074,N_24852,N_24996);
or UO_2075 (O_2075,N_24881,N_24981);
and UO_2076 (O_2076,N_24757,N_24935);
nor UO_2077 (O_2077,N_24842,N_24952);
or UO_2078 (O_2078,N_24794,N_24947);
nor UO_2079 (O_2079,N_24945,N_24989);
nand UO_2080 (O_2080,N_24951,N_24900);
or UO_2081 (O_2081,N_24767,N_24922);
and UO_2082 (O_2082,N_24856,N_24804);
or UO_2083 (O_2083,N_24860,N_24909);
nor UO_2084 (O_2084,N_24754,N_24795);
xnor UO_2085 (O_2085,N_24828,N_24758);
xor UO_2086 (O_2086,N_24881,N_24988);
nand UO_2087 (O_2087,N_24867,N_24787);
and UO_2088 (O_2088,N_24795,N_24968);
nor UO_2089 (O_2089,N_24890,N_24897);
and UO_2090 (O_2090,N_24762,N_24755);
xor UO_2091 (O_2091,N_24983,N_24964);
nor UO_2092 (O_2092,N_24807,N_24994);
or UO_2093 (O_2093,N_24831,N_24995);
nand UO_2094 (O_2094,N_24853,N_24873);
nand UO_2095 (O_2095,N_24913,N_24909);
and UO_2096 (O_2096,N_24886,N_24808);
xnor UO_2097 (O_2097,N_24903,N_24973);
nand UO_2098 (O_2098,N_24901,N_24963);
nand UO_2099 (O_2099,N_24891,N_24998);
or UO_2100 (O_2100,N_24914,N_24953);
nor UO_2101 (O_2101,N_24910,N_24974);
xor UO_2102 (O_2102,N_24852,N_24857);
nor UO_2103 (O_2103,N_24988,N_24930);
or UO_2104 (O_2104,N_24791,N_24895);
and UO_2105 (O_2105,N_24975,N_24937);
and UO_2106 (O_2106,N_24768,N_24822);
or UO_2107 (O_2107,N_24814,N_24973);
and UO_2108 (O_2108,N_24798,N_24874);
or UO_2109 (O_2109,N_24975,N_24791);
or UO_2110 (O_2110,N_24824,N_24986);
and UO_2111 (O_2111,N_24832,N_24979);
xnor UO_2112 (O_2112,N_24968,N_24763);
or UO_2113 (O_2113,N_24751,N_24882);
nor UO_2114 (O_2114,N_24760,N_24855);
nor UO_2115 (O_2115,N_24902,N_24839);
xnor UO_2116 (O_2116,N_24954,N_24822);
xnor UO_2117 (O_2117,N_24878,N_24942);
nor UO_2118 (O_2118,N_24793,N_24991);
nand UO_2119 (O_2119,N_24983,N_24971);
nor UO_2120 (O_2120,N_24909,N_24880);
nor UO_2121 (O_2121,N_24823,N_24953);
xnor UO_2122 (O_2122,N_24957,N_24860);
nand UO_2123 (O_2123,N_24998,N_24770);
and UO_2124 (O_2124,N_24844,N_24871);
nor UO_2125 (O_2125,N_24825,N_24799);
nand UO_2126 (O_2126,N_24862,N_24863);
xnor UO_2127 (O_2127,N_24983,N_24907);
nor UO_2128 (O_2128,N_24755,N_24900);
and UO_2129 (O_2129,N_24816,N_24999);
nand UO_2130 (O_2130,N_24795,N_24851);
nor UO_2131 (O_2131,N_24965,N_24862);
nand UO_2132 (O_2132,N_24848,N_24879);
or UO_2133 (O_2133,N_24831,N_24896);
nor UO_2134 (O_2134,N_24960,N_24891);
nor UO_2135 (O_2135,N_24839,N_24865);
nand UO_2136 (O_2136,N_24786,N_24859);
and UO_2137 (O_2137,N_24985,N_24914);
or UO_2138 (O_2138,N_24795,N_24899);
nor UO_2139 (O_2139,N_24818,N_24938);
or UO_2140 (O_2140,N_24840,N_24800);
or UO_2141 (O_2141,N_24821,N_24846);
nand UO_2142 (O_2142,N_24977,N_24843);
or UO_2143 (O_2143,N_24886,N_24840);
or UO_2144 (O_2144,N_24894,N_24877);
and UO_2145 (O_2145,N_24815,N_24820);
nand UO_2146 (O_2146,N_24752,N_24985);
or UO_2147 (O_2147,N_24785,N_24804);
nand UO_2148 (O_2148,N_24808,N_24850);
nor UO_2149 (O_2149,N_24820,N_24998);
nand UO_2150 (O_2150,N_24993,N_24882);
xor UO_2151 (O_2151,N_24870,N_24848);
xor UO_2152 (O_2152,N_24847,N_24824);
or UO_2153 (O_2153,N_24755,N_24843);
xor UO_2154 (O_2154,N_24961,N_24898);
or UO_2155 (O_2155,N_24846,N_24971);
nand UO_2156 (O_2156,N_24868,N_24963);
and UO_2157 (O_2157,N_24752,N_24831);
and UO_2158 (O_2158,N_24762,N_24991);
nand UO_2159 (O_2159,N_24988,N_24767);
or UO_2160 (O_2160,N_24789,N_24981);
nand UO_2161 (O_2161,N_24955,N_24802);
xnor UO_2162 (O_2162,N_24806,N_24847);
xnor UO_2163 (O_2163,N_24845,N_24989);
xnor UO_2164 (O_2164,N_24982,N_24999);
nor UO_2165 (O_2165,N_24821,N_24980);
nand UO_2166 (O_2166,N_24761,N_24778);
nand UO_2167 (O_2167,N_24878,N_24794);
nand UO_2168 (O_2168,N_24773,N_24859);
nor UO_2169 (O_2169,N_24796,N_24763);
nand UO_2170 (O_2170,N_24943,N_24998);
nor UO_2171 (O_2171,N_24818,N_24931);
and UO_2172 (O_2172,N_24972,N_24776);
and UO_2173 (O_2173,N_24861,N_24798);
nor UO_2174 (O_2174,N_24777,N_24911);
nor UO_2175 (O_2175,N_24993,N_24990);
nand UO_2176 (O_2176,N_24784,N_24932);
nand UO_2177 (O_2177,N_24851,N_24805);
and UO_2178 (O_2178,N_24952,N_24766);
nand UO_2179 (O_2179,N_24840,N_24762);
nand UO_2180 (O_2180,N_24980,N_24960);
nand UO_2181 (O_2181,N_24848,N_24762);
or UO_2182 (O_2182,N_24752,N_24862);
nand UO_2183 (O_2183,N_24893,N_24959);
or UO_2184 (O_2184,N_24890,N_24879);
or UO_2185 (O_2185,N_24895,N_24900);
xnor UO_2186 (O_2186,N_24873,N_24814);
nor UO_2187 (O_2187,N_24777,N_24874);
nor UO_2188 (O_2188,N_24750,N_24881);
or UO_2189 (O_2189,N_24835,N_24989);
and UO_2190 (O_2190,N_24812,N_24891);
or UO_2191 (O_2191,N_24977,N_24808);
nor UO_2192 (O_2192,N_24962,N_24780);
nand UO_2193 (O_2193,N_24787,N_24759);
xor UO_2194 (O_2194,N_24926,N_24884);
nand UO_2195 (O_2195,N_24950,N_24759);
xor UO_2196 (O_2196,N_24967,N_24790);
or UO_2197 (O_2197,N_24780,N_24858);
nor UO_2198 (O_2198,N_24803,N_24796);
or UO_2199 (O_2199,N_24952,N_24795);
nand UO_2200 (O_2200,N_24788,N_24750);
nor UO_2201 (O_2201,N_24854,N_24818);
and UO_2202 (O_2202,N_24784,N_24985);
xnor UO_2203 (O_2203,N_24855,N_24830);
xnor UO_2204 (O_2204,N_24845,N_24871);
xor UO_2205 (O_2205,N_24798,N_24907);
nand UO_2206 (O_2206,N_24925,N_24885);
nor UO_2207 (O_2207,N_24859,N_24977);
nor UO_2208 (O_2208,N_24822,N_24982);
and UO_2209 (O_2209,N_24819,N_24764);
xor UO_2210 (O_2210,N_24900,N_24949);
nand UO_2211 (O_2211,N_24910,N_24776);
xor UO_2212 (O_2212,N_24924,N_24761);
nand UO_2213 (O_2213,N_24996,N_24863);
xnor UO_2214 (O_2214,N_24766,N_24947);
nor UO_2215 (O_2215,N_24792,N_24970);
and UO_2216 (O_2216,N_24998,N_24931);
nor UO_2217 (O_2217,N_24891,N_24823);
and UO_2218 (O_2218,N_24890,N_24822);
nand UO_2219 (O_2219,N_24754,N_24926);
xor UO_2220 (O_2220,N_24992,N_24960);
nand UO_2221 (O_2221,N_24911,N_24868);
or UO_2222 (O_2222,N_24958,N_24772);
and UO_2223 (O_2223,N_24962,N_24897);
and UO_2224 (O_2224,N_24937,N_24752);
xnor UO_2225 (O_2225,N_24936,N_24851);
or UO_2226 (O_2226,N_24999,N_24860);
nand UO_2227 (O_2227,N_24994,N_24959);
nand UO_2228 (O_2228,N_24877,N_24803);
nand UO_2229 (O_2229,N_24751,N_24837);
nand UO_2230 (O_2230,N_24881,N_24910);
or UO_2231 (O_2231,N_24956,N_24978);
nand UO_2232 (O_2232,N_24792,N_24822);
or UO_2233 (O_2233,N_24884,N_24985);
xnor UO_2234 (O_2234,N_24890,N_24797);
nand UO_2235 (O_2235,N_24934,N_24841);
or UO_2236 (O_2236,N_24939,N_24778);
nand UO_2237 (O_2237,N_24917,N_24777);
nand UO_2238 (O_2238,N_24865,N_24913);
xor UO_2239 (O_2239,N_24978,N_24891);
xnor UO_2240 (O_2240,N_24902,N_24753);
nand UO_2241 (O_2241,N_24935,N_24923);
xor UO_2242 (O_2242,N_24767,N_24794);
xnor UO_2243 (O_2243,N_24918,N_24823);
nand UO_2244 (O_2244,N_24999,N_24948);
and UO_2245 (O_2245,N_24984,N_24983);
nor UO_2246 (O_2246,N_24996,N_24957);
nand UO_2247 (O_2247,N_24981,N_24932);
or UO_2248 (O_2248,N_24774,N_24816);
xnor UO_2249 (O_2249,N_24780,N_24987);
nor UO_2250 (O_2250,N_24848,N_24764);
xor UO_2251 (O_2251,N_24966,N_24775);
or UO_2252 (O_2252,N_24920,N_24754);
xnor UO_2253 (O_2253,N_24843,N_24952);
or UO_2254 (O_2254,N_24897,N_24943);
nor UO_2255 (O_2255,N_24888,N_24937);
and UO_2256 (O_2256,N_24781,N_24864);
nor UO_2257 (O_2257,N_24997,N_24957);
xor UO_2258 (O_2258,N_24770,N_24881);
and UO_2259 (O_2259,N_24821,N_24879);
xnor UO_2260 (O_2260,N_24775,N_24814);
nor UO_2261 (O_2261,N_24804,N_24794);
nand UO_2262 (O_2262,N_24928,N_24908);
or UO_2263 (O_2263,N_24901,N_24979);
and UO_2264 (O_2264,N_24960,N_24768);
nand UO_2265 (O_2265,N_24983,N_24913);
and UO_2266 (O_2266,N_24785,N_24882);
xnor UO_2267 (O_2267,N_24826,N_24959);
xnor UO_2268 (O_2268,N_24796,N_24832);
and UO_2269 (O_2269,N_24884,N_24825);
nor UO_2270 (O_2270,N_24803,N_24830);
xor UO_2271 (O_2271,N_24815,N_24863);
nand UO_2272 (O_2272,N_24926,N_24995);
and UO_2273 (O_2273,N_24987,N_24944);
xor UO_2274 (O_2274,N_24912,N_24765);
nor UO_2275 (O_2275,N_24809,N_24912);
and UO_2276 (O_2276,N_24945,N_24926);
or UO_2277 (O_2277,N_24891,N_24900);
nor UO_2278 (O_2278,N_24763,N_24868);
xnor UO_2279 (O_2279,N_24920,N_24803);
nand UO_2280 (O_2280,N_24860,N_24928);
xnor UO_2281 (O_2281,N_24961,N_24760);
or UO_2282 (O_2282,N_24938,N_24795);
or UO_2283 (O_2283,N_24868,N_24840);
nor UO_2284 (O_2284,N_24867,N_24975);
nand UO_2285 (O_2285,N_24851,N_24881);
xor UO_2286 (O_2286,N_24866,N_24818);
xnor UO_2287 (O_2287,N_24820,N_24762);
nand UO_2288 (O_2288,N_24951,N_24871);
nor UO_2289 (O_2289,N_24992,N_24766);
xnor UO_2290 (O_2290,N_24946,N_24762);
xnor UO_2291 (O_2291,N_24923,N_24957);
nor UO_2292 (O_2292,N_24860,N_24843);
nand UO_2293 (O_2293,N_24827,N_24869);
xnor UO_2294 (O_2294,N_24984,N_24999);
and UO_2295 (O_2295,N_24817,N_24809);
and UO_2296 (O_2296,N_24911,N_24805);
or UO_2297 (O_2297,N_24828,N_24812);
and UO_2298 (O_2298,N_24802,N_24999);
or UO_2299 (O_2299,N_24921,N_24948);
nor UO_2300 (O_2300,N_24932,N_24913);
nand UO_2301 (O_2301,N_24795,N_24839);
nand UO_2302 (O_2302,N_24974,N_24918);
nand UO_2303 (O_2303,N_24946,N_24824);
and UO_2304 (O_2304,N_24756,N_24891);
nand UO_2305 (O_2305,N_24975,N_24878);
and UO_2306 (O_2306,N_24908,N_24893);
xnor UO_2307 (O_2307,N_24985,N_24936);
xor UO_2308 (O_2308,N_24941,N_24975);
and UO_2309 (O_2309,N_24866,N_24975);
and UO_2310 (O_2310,N_24760,N_24877);
or UO_2311 (O_2311,N_24755,N_24826);
and UO_2312 (O_2312,N_24849,N_24964);
and UO_2313 (O_2313,N_24926,N_24823);
nand UO_2314 (O_2314,N_24843,N_24853);
xnor UO_2315 (O_2315,N_24837,N_24897);
nor UO_2316 (O_2316,N_24894,N_24955);
nand UO_2317 (O_2317,N_24907,N_24955);
nand UO_2318 (O_2318,N_24876,N_24834);
nand UO_2319 (O_2319,N_24966,N_24761);
or UO_2320 (O_2320,N_24764,N_24817);
nor UO_2321 (O_2321,N_24952,N_24874);
or UO_2322 (O_2322,N_24920,N_24851);
nor UO_2323 (O_2323,N_24899,N_24801);
nor UO_2324 (O_2324,N_24799,N_24918);
and UO_2325 (O_2325,N_24957,N_24893);
nand UO_2326 (O_2326,N_24978,N_24865);
nor UO_2327 (O_2327,N_24780,N_24791);
nor UO_2328 (O_2328,N_24766,N_24903);
and UO_2329 (O_2329,N_24888,N_24844);
nand UO_2330 (O_2330,N_24879,N_24854);
and UO_2331 (O_2331,N_24798,N_24828);
xnor UO_2332 (O_2332,N_24791,N_24897);
nand UO_2333 (O_2333,N_24941,N_24982);
or UO_2334 (O_2334,N_24904,N_24897);
xor UO_2335 (O_2335,N_24954,N_24807);
xor UO_2336 (O_2336,N_24809,N_24887);
xor UO_2337 (O_2337,N_24815,N_24862);
or UO_2338 (O_2338,N_24994,N_24930);
nand UO_2339 (O_2339,N_24792,N_24991);
nand UO_2340 (O_2340,N_24764,N_24956);
nor UO_2341 (O_2341,N_24844,N_24873);
or UO_2342 (O_2342,N_24784,N_24979);
xnor UO_2343 (O_2343,N_24987,N_24886);
xor UO_2344 (O_2344,N_24838,N_24908);
nand UO_2345 (O_2345,N_24791,N_24971);
nand UO_2346 (O_2346,N_24866,N_24769);
nor UO_2347 (O_2347,N_24986,N_24992);
xnor UO_2348 (O_2348,N_24842,N_24962);
or UO_2349 (O_2349,N_24781,N_24957);
and UO_2350 (O_2350,N_24819,N_24752);
or UO_2351 (O_2351,N_24990,N_24944);
nor UO_2352 (O_2352,N_24976,N_24854);
or UO_2353 (O_2353,N_24764,N_24978);
or UO_2354 (O_2354,N_24969,N_24752);
nor UO_2355 (O_2355,N_24991,N_24943);
xnor UO_2356 (O_2356,N_24886,N_24767);
or UO_2357 (O_2357,N_24960,N_24973);
and UO_2358 (O_2358,N_24864,N_24999);
and UO_2359 (O_2359,N_24751,N_24887);
nor UO_2360 (O_2360,N_24820,N_24772);
nand UO_2361 (O_2361,N_24922,N_24901);
xnor UO_2362 (O_2362,N_24789,N_24994);
nor UO_2363 (O_2363,N_24912,N_24770);
xor UO_2364 (O_2364,N_24778,N_24860);
nor UO_2365 (O_2365,N_24845,N_24858);
xor UO_2366 (O_2366,N_24753,N_24829);
xor UO_2367 (O_2367,N_24990,N_24817);
and UO_2368 (O_2368,N_24955,N_24857);
nand UO_2369 (O_2369,N_24967,N_24896);
nor UO_2370 (O_2370,N_24939,N_24793);
or UO_2371 (O_2371,N_24903,N_24864);
xor UO_2372 (O_2372,N_24751,N_24985);
nor UO_2373 (O_2373,N_24887,N_24831);
xnor UO_2374 (O_2374,N_24803,N_24941);
nand UO_2375 (O_2375,N_24851,N_24816);
and UO_2376 (O_2376,N_24836,N_24946);
and UO_2377 (O_2377,N_24923,N_24789);
xor UO_2378 (O_2378,N_24928,N_24976);
xnor UO_2379 (O_2379,N_24835,N_24905);
or UO_2380 (O_2380,N_24930,N_24978);
nand UO_2381 (O_2381,N_24970,N_24769);
and UO_2382 (O_2382,N_24897,N_24840);
and UO_2383 (O_2383,N_24811,N_24998);
or UO_2384 (O_2384,N_24993,N_24853);
and UO_2385 (O_2385,N_24825,N_24883);
xnor UO_2386 (O_2386,N_24988,N_24879);
nand UO_2387 (O_2387,N_24873,N_24798);
or UO_2388 (O_2388,N_24786,N_24753);
and UO_2389 (O_2389,N_24937,N_24885);
and UO_2390 (O_2390,N_24979,N_24790);
and UO_2391 (O_2391,N_24975,N_24862);
or UO_2392 (O_2392,N_24912,N_24830);
xnor UO_2393 (O_2393,N_24852,N_24871);
xor UO_2394 (O_2394,N_24875,N_24953);
xnor UO_2395 (O_2395,N_24906,N_24822);
xor UO_2396 (O_2396,N_24845,N_24818);
or UO_2397 (O_2397,N_24771,N_24917);
and UO_2398 (O_2398,N_24804,N_24911);
nor UO_2399 (O_2399,N_24807,N_24949);
nand UO_2400 (O_2400,N_24776,N_24827);
nand UO_2401 (O_2401,N_24811,N_24983);
and UO_2402 (O_2402,N_24919,N_24959);
nor UO_2403 (O_2403,N_24973,N_24829);
nand UO_2404 (O_2404,N_24766,N_24904);
nand UO_2405 (O_2405,N_24931,N_24853);
nand UO_2406 (O_2406,N_24928,N_24980);
xor UO_2407 (O_2407,N_24878,N_24908);
or UO_2408 (O_2408,N_24857,N_24807);
xor UO_2409 (O_2409,N_24852,N_24806);
or UO_2410 (O_2410,N_24763,N_24805);
and UO_2411 (O_2411,N_24769,N_24764);
and UO_2412 (O_2412,N_24753,N_24751);
xnor UO_2413 (O_2413,N_24853,N_24844);
and UO_2414 (O_2414,N_24878,N_24911);
xnor UO_2415 (O_2415,N_24798,N_24797);
nor UO_2416 (O_2416,N_24851,N_24802);
nand UO_2417 (O_2417,N_24888,N_24895);
nor UO_2418 (O_2418,N_24935,N_24934);
xnor UO_2419 (O_2419,N_24846,N_24861);
and UO_2420 (O_2420,N_24849,N_24867);
and UO_2421 (O_2421,N_24919,N_24834);
nand UO_2422 (O_2422,N_24762,N_24769);
and UO_2423 (O_2423,N_24911,N_24834);
xor UO_2424 (O_2424,N_24837,N_24758);
nand UO_2425 (O_2425,N_24970,N_24964);
and UO_2426 (O_2426,N_24982,N_24968);
or UO_2427 (O_2427,N_24818,N_24894);
and UO_2428 (O_2428,N_24803,N_24926);
or UO_2429 (O_2429,N_24878,N_24978);
or UO_2430 (O_2430,N_24857,N_24910);
and UO_2431 (O_2431,N_24864,N_24984);
or UO_2432 (O_2432,N_24882,N_24973);
nor UO_2433 (O_2433,N_24962,N_24807);
and UO_2434 (O_2434,N_24941,N_24832);
nor UO_2435 (O_2435,N_24895,N_24935);
xnor UO_2436 (O_2436,N_24946,N_24986);
and UO_2437 (O_2437,N_24960,N_24786);
and UO_2438 (O_2438,N_24976,N_24924);
nor UO_2439 (O_2439,N_24796,N_24981);
nand UO_2440 (O_2440,N_24788,N_24765);
and UO_2441 (O_2441,N_24928,N_24847);
and UO_2442 (O_2442,N_24869,N_24837);
and UO_2443 (O_2443,N_24930,N_24850);
nor UO_2444 (O_2444,N_24931,N_24870);
nor UO_2445 (O_2445,N_24757,N_24865);
nor UO_2446 (O_2446,N_24815,N_24904);
xor UO_2447 (O_2447,N_24945,N_24877);
xor UO_2448 (O_2448,N_24861,N_24992);
xor UO_2449 (O_2449,N_24957,N_24845);
or UO_2450 (O_2450,N_24981,N_24833);
nand UO_2451 (O_2451,N_24809,N_24945);
nand UO_2452 (O_2452,N_24992,N_24982);
nand UO_2453 (O_2453,N_24821,N_24789);
nand UO_2454 (O_2454,N_24948,N_24883);
nor UO_2455 (O_2455,N_24859,N_24844);
nor UO_2456 (O_2456,N_24837,N_24816);
or UO_2457 (O_2457,N_24901,N_24821);
or UO_2458 (O_2458,N_24911,N_24752);
and UO_2459 (O_2459,N_24784,N_24935);
or UO_2460 (O_2460,N_24995,N_24761);
nor UO_2461 (O_2461,N_24853,N_24834);
nand UO_2462 (O_2462,N_24977,N_24846);
xnor UO_2463 (O_2463,N_24816,N_24880);
xnor UO_2464 (O_2464,N_24910,N_24900);
nor UO_2465 (O_2465,N_24795,N_24813);
nor UO_2466 (O_2466,N_24840,N_24971);
and UO_2467 (O_2467,N_24776,N_24956);
xor UO_2468 (O_2468,N_24769,N_24759);
or UO_2469 (O_2469,N_24954,N_24937);
nor UO_2470 (O_2470,N_24820,N_24878);
and UO_2471 (O_2471,N_24817,N_24936);
or UO_2472 (O_2472,N_24881,N_24924);
xnor UO_2473 (O_2473,N_24841,N_24838);
nand UO_2474 (O_2474,N_24896,N_24873);
nand UO_2475 (O_2475,N_24839,N_24952);
and UO_2476 (O_2476,N_24861,N_24774);
nor UO_2477 (O_2477,N_24805,N_24981);
and UO_2478 (O_2478,N_24808,N_24777);
nand UO_2479 (O_2479,N_24799,N_24933);
or UO_2480 (O_2480,N_24857,N_24896);
xnor UO_2481 (O_2481,N_24988,N_24943);
xnor UO_2482 (O_2482,N_24842,N_24767);
nor UO_2483 (O_2483,N_24986,N_24951);
nor UO_2484 (O_2484,N_24753,N_24938);
nor UO_2485 (O_2485,N_24932,N_24931);
and UO_2486 (O_2486,N_24837,N_24750);
and UO_2487 (O_2487,N_24780,N_24870);
xor UO_2488 (O_2488,N_24936,N_24962);
nand UO_2489 (O_2489,N_24895,N_24856);
and UO_2490 (O_2490,N_24954,N_24992);
nor UO_2491 (O_2491,N_24759,N_24811);
or UO_2492 (O_2492,N_24976,N_24793);
nand UO_2493 (O_2493,N_24842,N_24751);
xnor UO_2494 (O_2494,N_24901,N_24756);
or UO_2495 (O_2495,N_24905,N_24986);
and UO_2496 (O_2496,N_24795,N_24957);
xnor UO_2497 (O_2497,N_24833,N_24998);
nand UO_2498 (O_2498,N_24920,N_24996);
xor UO_2499 (O_2499,N_24807,N_24839);
or UO_2500 (O_2500,N_24853,N_24960);
nor UO_2501 (O_2501,N_24810,N_24893);
or UO_2502 (O_2502,N_24773,N_24938);
nor UO_2503 (O_2503,N_24825,N_24779);
nand UO_2504 (O_2504,N_24767,N_24755);
and UO_2505 (O_2505,N_24947,N_24772);
nor UO_2506 (O_2506,N_24977,N_24925);
or UO_2507 (O_2507,N_24784,N_24892);
nor UO_2508 (O_2508,N_24869,N_24812);
or UO_2509 (O_2509,N_24872,N_24875);
or UO_2510 (O_2510,N_24793,N_24790);
and UO_2511 (O_2511,N_24905,N_24883);
and UO_2512 (O_2512,N_24924,N_24899);
and UO_2513 (O_2513,N_24956,N_24896);
nand UO_2514 (O_2514,N_24859,N_24807);
nand UO_2515 (O_2515,N_24764,N_24875);
xor UO_2516 (O_2516,N_24794,N_24845);
nand UO_2517 (O_2517,N_24920,N_24831);
nand UO_2518 (O_2518,N_24808,N_24782);
xor UO_2519 (O_2519,N_24914,N_24858);
and UO_2520 (O_2520,N_24881,N_24891);
nand UO_2521 (O_2521,N_24760,N_24952);
xor UO_2522 (O_2522,N_24879,N_24907);
nand UO_2523 (O_2523,N_24858,N_24930);
nand UO_2524 (O_2524,N_24890,N_24821);
nand UO_2525 (O_2525,N_24856,N_24803);
nand UO_2526 (O_2526,N_24767,N_24897);
nor UO_2527 (O_2527,N_24845,N_24929);
nand UO_2528 (O_2528,N_24798,N_24768);
and UO_2529 (O_2529,N_24816,N_24801);
or UO_2530 (O_2530,N_24924,N_24767);
and UO_2531 (O_2531,N_24968,N_24823);
or UO_2532 (O_2532,N_24927,N_24880);
xnor UO_2533 (O_2533,N_24813,N_24936);
nand UO_2534 (O_2534,N_24952,N_24832);
xor UO_2535 (O_2535,N_24925,N_24869);
or UO_2536 (O_2536,N_24916,N_24762);
xor UO_2537 (O_2537,N_24818,N_24985);
xor UO_2538 (O_2538,N_24965,N_24811);
nor UO_2539 (O_2539,N_24948,N_24942);
nand UO_2540 (O_2540,N_24814,N_24916);
xnor UO_2541 (O_2541,N_24966,N_24980);
nor UO_2542 (O_2542,N_24840,N_24933);
and UO_2543 (O_2543,N_24998,N_24761);
xor UO_2544 (O_2544,N_24840,N_24988);
or UO_2545 (O_2545,N_24816,N_24784);
or UO_2546 (O_2546,N_24927,N_24978);
and UO_2547 (O_2547,N_24835,N_24794);
xnor UO_2548 (O_2548,N_24809,N_24960);
nand UO_2549 (O_2549,N_24985,N_24918);
nand UO_2550 (O_2550,N_24880,N_24804);
xnor UO_2551 (O_2551,N_24914,N_24987);
or UO_2552 (O_2552,N_24927,N_24984);
nor UO_2553 (O_2553,N_24836,N_24806);
or UO_2554 (O_2554,N_24794,N_24806);
nor UO_2555 (O_2555,N_24866,N_24963);
nand UO_2556 (O_2556,N_24970,N_24770);
xnor UO_2557 (O_2557,N_24959,N_24825);
xnor UO_2558 (O_2558,N_24870,N_24889);
and UO_2559 (O_2559,N_24858,N_24950);
xor UO_2560 (O_2560,N_24836,N_24921);
xnor UO_2561 (O_2561,N_24836,N_24914);
xor UO_2562 (O_2562,N_24779,N_24969);
nand UO_2563 (O_2563,N_24889,N_24767);
or UO_2564 (O_2564,N_24833,N_24782);
nand UO_2565 (O_2565,N_24907,N_24991);
and UO_2566 (O_2566,N_24819,N_24940);
nand UO_2567 (O_2567,N_24753,N_24996);
nand UO_2568 (O_2568,N_24895,N_24863);
and UO_2569 (O_2569,N_24827,N_24907);
nand UO_2570 (O_2570,N_24885,N_24808);
nor UO_2571 (O_2571,N_24856,N_24805);
nand UO_2572 (O_2572,N_24910,N_24989);
nor UO_2573 (O_2573,N_24803,N_24868);
xnor UO_2574 (O_2574,N_24920,N_24768);
or UO_2575 (O_2575,N_24811,N_24752);
or UO_2576 (O_2576,N_24905,N_24936);
and UO_2577 (O_2577,N_24807,N_24894);
or UO_2578 (O_2578,N_24885,N_24832);
and UO_2579 (O_2579,N_24852,N_24773);
nor UO_2580 (O_2580,N_24902,N_24853);
nor UO_2581 (O_2581,N_24881,N_24898);
or UO_2582 (O_2582,N_24854,N_24857);
nor UO_2583 (O_2583,N_24940,N_24956);
and UO_2584 (O_2584,N_24936,N_24789);
xnor UO_2585 (O_2585,N_24841,N_24755);
and UO_2586 (O_2586,N_24874,N_24896);
nand UO_2587 (O_2587,N_24884,N_24861);
xor UO_2588 (O_2588,N_24997,N_24767);
nand UO_2589 (O_2589,N_24823,N_24937);
or UO_2590 (O_2590,N_24765,N_24795);
nand UO_2591 (O_2591,N_24867,N_24770);
xor UO_2592 (O_2592,N_24835,N_24829);
nor UO_2593 (O_2593,N_24787,N_24857);
and UO_2594 (O_2594,N_24820,N_24895);
or UO_2595 (O_2595,N_24891,N_24829);
or UO_2596 (O_2596,N_24798,N_24923);
xnor UO_2597 (O_2597,N_24759,N_24834);
nand UO_2598 (O_2598,N_24754,N_24830);
or UO_2599 (O_2599,N_24771,N_24963);
nand UO_2600 (O_2600,N_24926,N_24940);
or UO_2601 (O_2601,N_24889,N_24828);
nand UO_2602 (O_2602,N_24998,N_24829);
xor UO_2603 (O_2603,N_24965,N_24764);
nor UO_2604 (O_2604,N_24975,N_24946);
or UO_2605 (O_2605,N_24840,N_24976);
or UO_2606 (O_2606,N_24823,N_24976);
nor UO_2607 (O_2607,N_24984,N_24843);
nand UO_2608 (O_2608,N_24830,N_24832);
nor UO_2609 (O_2609,N_24764,N_24865);
nor UO_2610 (O_2610,N_24762,N_24888);
nor UO_2611 (O_2611,N_24813,N_24937);
xor UO_2612 (O_2612,N_24984,N_24830);
nand UO_2613 (O_2613,N_24886,N_24896);
xnor UO_2614 (O_2614,N_24752,N_24962);
xor UO_2615 (O_2615,N_24965,N_24779);
or UO_2616 (O_2616,N_24964,N_24845);
or UO_2617 (O_2617,N_24843,N_24777);
nor UO_2618 (O_2618,N_24854,N_24796);
or UO_2619 (O_2619,N_24938,N_24973);
or UO_2620 (O_2620,N_24803,N_24865);
or UO_2621 (O_2621,N_24987,N_24984);
nand UO_2622 (O_2622,N_24908,N_24982);
xor UO_2623 (O_2623,N_24757,N_24858);
nor UO_2624 (O_2624,N_24892,N_24842);
xor UO_2625 (O_2625,N_24936,N_24928);
or UO_2626 (O_2626,N_24817,N_24806);
nor UO_2627 (O_2627,N_24942,N_24971);
nand UO_2628 (O_2628,N_24835,N_24910);
and UO_2629 (O_2629,N_24827,N_24996);
nand UO_2630 (O_2630,N_24860,N_24806);
nor UO_2631 (O_2631,N_24823,N_24804);
nand UO_2632 (O_2632,N_24868,N_24949);
xnor UO_2633 (O_2633,N_24773,N_24947);
nand UO_2634 (O_2634,N_24940,N_24786);
nand UO_2635 (O_2635,N_24896,N_24927);
nor UO_2636 (O_2636,N_24750,N_24919);
xnor UO_2637 (O_2637,N_24926,N_24961);
nand UO_2638 (O_2638,N_24981,N_24880);
nor UO_2639 (O_2639,N_24879,N_24847);
nor UO_2640 (O_2640,N_24834,N_24894);
nand UO_2641 (O_2641,N_24850,N_24758);
nor UO_2642 (O_2642,N_24953,N_24999);
nand UO_2643 (O_2643,N_24910,N_24897);
and UO_2644 (O_2644,N_24812,N_24942);
nor UO_2645 (O_2645,N_24775,N_24995);
nor UO_2646 (O_2646,N_24934,N_24893);
and UO_2647 (O_2647,N_24875,N_24998);
nand UO_2648 (O_2648,N_24773,N_24788);
and UO_2649 (O_2649,N_24762,N_24815);
or UO_2650 (O_2650,N_24780,N_24971);
nor UO_2651 (O_2651,N_24902,N_24873);
nand UO_2652 (O_2652,N_24998,N_24848);
nand UO_2653 (O_2653,N_24761,N_24888);
or UO_2654 (O_2654,N_24975,N_24877);
and UO_2655 (O_2655,N_24767,N_24908);
or UO_2656 (O_2656,N_24790,N_24807);
xnor UO_2657 (O_2657,N_24966,N_24988);
or UO_2658 (O_2658,N_24933,N_24851);
xnor UO_2659 (O_2659,N_24750,N_24950);
or UO_2660 (O_2660,N_24765,N_24942);
and UO_2661 (O_2661,N_24762,N_24982);
xnor UO_2662 (O_2662,N_24919,N_24969);
and UO_2663 (O_2663,N_24755,N_24760);
xnor UO_2664 (O_2664,N_24962,N_24906);
and UO_2665 (O_2665,N_24907,N_24949);
or UO_2666 (O_2666,N_24866,N_24798);
xor UO_2667 (O_2667,N_24999,N_24893);
xor UO_2668 (O_2668,N_24934,N_24945);
xnor UO_2669 (O_2669,N_24995,N_24795);
nor UO_2670 (O_2670,N_24961,N_24928);
and UO_2671 (O_2671,N_24915,N_24859);
nor UO_2672 (O_2672,N_24846,N_24918);
nor UO_2673 (O_2673,N_24841,N_24751);
or UO_2674 (O_2674,N_24901,N_24953);
and UO_2675 (O_2675,N_24868,N_24777);
or UO_2676 (O_2676,N_24756,N_24850);
and UO_2677 (O_2677,N_24866,N_24839);
nor UO_2678 (O_2678,N_24790,N_24843);
or UO_2679 (O_2679,N_24850,N_24989);
nor UO_2680 (O_2680,N_24946,N_24944);
nor UO_2681 (O_2681,N_24809,N_24868);
and UO_2682 (O_2682,N_24985,N_24959);
and UO_2683 (O_2683,N_24836,N_24809);
and UO_2684 (O_2684,N_24884,N_24936);
nor UO_2685 (O_2685,N_24767,N_24758);
or UO_2686 (O_2686,N_24884,N_24920);
or UO_2687 (O_2687,N_24793,N_24819);
and UO_2688 (O_2688,N_24949,N_24806);
and UO_2689 (O_2689,N_24975,N_24800);
nand UO_2690 (O_2690,N_24939,N_24870);
nor UO_2691 (O_2691,N_24969,N_24908);
and UO_2692 (O_2692,N_24952,N_24878);
and UO_2693 (O_2693,N_24993,N_24937);
or UO_2694 (O_2694,N_24816,N_24986);
or UO_2695 (O_2695,N_24869,N_24879);
xor UO_2696 (O_2696,N_24763,N_24855);
or UO_2697 (O_2697,N_24952,N_24971);
and UO_2698 (O_2698,N_24969,N_24901);
and UO_2699 (O_2699,N_24884,N_24893);
nor UO_2700 (O_2700,N_24904,N_24790);
xor UO_2701 (O_2701,N_24845,N_24882);
xnor UO_2702 (O_2702,N_24866,N_24842);
nand UO_2703 (O_2703,N_24861,N_24965);
or UO_2704 (O_2704,N_24786,N_24945);
nand UO_2705 (O_2705,N_24792,N_24956);
nor UO_2706 (O_2706,N_24949,N_24780);
or UO_2707 (O_2707,N_24757,N_24981);
and UO_2708 (O_2708,N_24752,N_24908);
and UO_2709 (O_2709,N_24854,N_24783);
or UO_2710 (O_2710,N_24846,N_24794);
xnor UO_2711 (O_2711,N_24905,N_24904);
xor UO_2712 (O_2712,N_24922,N_24915);
nor UO_2713 (O_2713,N_24999,N_24994);
and UO_2714 (O_2714,N_24791,N_24984);
xnor UO_2715 (O_2715,N_24776,N_24769);
nand UO_2716 (O_2716,N_24839,N_24962);
xnor UO_2717 (O_2717,N_24868,N_24897);
xnor UO_2718 (O_2718,N_24821,N_24978);
and UO_2719 (O_2719,N_24838,N_24850);
nor UO_2720 (O_2720,N_24785,N_24912);
nor UO_2721 (O_2721,N_24868,N_24969);
and UO_2722 (O_2722,N_24884,N_24913);
xor UO_2723 (O_2723,N_24887,N_24801);
or UO_2724 (O_2724,N_24933,N_24835);
nor UO_2725 (O_2725,N_24847,N_24789);
or UO_2726 (O_2726,N_24943,N_24838);
nor UO_2727 (O_2727,N_24832,N_24750);
nor UO_2728 (O_2728,N_24896,N_24756);
nand UO_2729 (O_2729,N_24841,N_24779);
and UO_2730 (O_2730,N_24826,N_24938);
nand UO_2731 (O_2731,N_24954,N_24922);
and UO_2732 (O_2732,N_24790,N_24983);
or UO_2733 (O_2733,N_24795,N_24858);
xnor UO_2734 (O_2734,N_24915,N_24940);
or UO_2735 (O_2735,N_24897,N_24831);
nand UO_2736 (O_2736,N_24977,N_24839);
xnor UO_2737 (O_2737,N_24752,N_24922);
nor UO_2738 (O_2738,N_24927,N_24817);
and UO_2739 (O_2739,N_24966,N_24938);
and UO_2740 (O_2740,N_24983,N_24930);
nor UO_2741 (O_2741,N_24764,N_24750);
xnor UO_2742 (O_2742,N_24954,N_24804);
nand UO_2743 (O_2743,N_24890,N_24995);
xnor UO_2744 (O_2744,N_24971,N_24771);
or UO_2745 (O_2745,N_24885,N_24971);
and UO_2746 (O_2746,N_24921,N_24880);
and UO_2747 (O_2747,N_24906,N_24919);
and UO_2748 (O_2748,N_24960,N_24778);
or UO_2749 (O_2749,N_24904,N_24891);
or UO_2750 (O_2750,N_24930,N_24821);
and UO_2751 (O_2751,N_24936,N_24804);
nand UO_2752 (O_2752,N_24861,N_24935);
nor UO_2753 (O_2753,N_24754,N_24991);
xnor UO_2754 (O_2754,N_24974,N_24828);
nand UO_2755 (O_2755,N_24819,N_24840);
and UO_2756 (O_2756,N_24821,N_24947);
or UO_2757 (O_2757,N_24858,N_24776);
or UO_2758 (O_2758,N_24956,N_24894);
nand UO_2759 (O_2759,N_24976,N_24808);
and UO_2760 (O_2760,N_24797,N_24762);
and UO_2761 (O_2761,N_24987,N_24969);
and UO_2762 (O_2762,N_24896,N_24916);
or UO_2763 (O_2763,N_24875,N_24968);
nor UO_2764 (O_2764,N_24931,N_24894);
and UO_2765 (O_2765,N_24945,N_24841);
or UO_2766 (O_2766,N_24861,N_24850);
or UO_2767 (O_2767,N_24831,N_24948);
or UO_2768 (O_2768,N_24792,N_24805);
xor UO_2769 (O_2769,N_24784,N_24843);
nand UO_2770 (O_2770,N_24865,N_24965);
or UO_2771 (O_2771,N_24935,N_24903);
xnor UO_2772 (O_2772,N_24846,N_24963);
and UO_2773 (O_2773,N_24963,N_24931);
xnor UO_2774 (O_2774,N_24867,N_24903);
and UO_2775 (O_2775,N_24775,N_24964);
or UO_2776 (O_2776,N_24852,N_24766);
nand UO_2777 (O_2777,N_24968,N_24768);
xnor UO_2778 (O_2778,N_24823,N_24896);
nand UO_2779 (O_2779,N_24834,N_24862);
or UO_2780 (O_2780,N_24902,N_24973);
or UO_2781 (O_2781,N_24962,N_24868);
nor UO_2782 (O_2782,N_24792,N_24852);
or UO_2783 (O_2783,N_24920,N_24975);
nand UO_2784 (O_2784,N_24820,N_24855);
nor UO_2785 (O_2785,N_24834,N_24931);
nand UO_2786 (O_2786,N_24875,N_24865);
xor UO_2787 (O_2787,N_24997,N_24936);
or UO_2788 (O_2788,N_24889,N_24915);
or UO_2789 (O_2789,N_24759,N_24817);
and UO_2790 (O_2790,N_24950,N_24937);
nor UO_2791 (O_2791,N_24818,N_24802);
nor UO_2792 (O_2792,N_24801,N_24938);
xnor UO_2793 (O_2793,N_24950,N_24993);
nor UO_2794 (O_2794,N_24973,N_24955);
nor UO_2795 (O_2795,N_24902,N_24851);
xnor UO_2796 (O_2796,N_24985,N_24830);
nand UO_2797 (O_2797,N_24928,N_24809);
nor UO_2798 (O_2798,N_24861,N_24795);
nand UO_2799 (O_2799,N_24950,N_24819);
nand UO_2800 (O_2800,N_24820,N_24911);
nand UO_2801 (O_2801,N_24955,N_24869);
nor UO_2802 (O_2802,N_24844,N_24807);
xnor UO_2803 (O_2803,N_24963,N_24983);
nor UO_2804 (O_2804,N_24978,N_24825);
nand UO_2805 (O_2805,N_24835,N_24775);
and UO_2806 (O_2806,N_24844,N_24783);
xnor UO_2807 (O_2807,N_24952,N_24865);
nor UO_2808 (O_2808,N_24921,N_24853);
xnor UO_2809 (O_2809,N_24757,N_24808);
nor UO_2810 (O_2810,N_24966,N_24992);
and UO_2811 (O_2811,N_24797,N_24832);
or UO_2812 (O_2812,N_24915,N_24928);
nor UO_2813 (O_2813,N_24921,N_24760);
nand UO_2814 (O_2814,N_24818,N_24979);
or UO_2815 (O_2815,N_24981,N_24842);
nand UO_2816 (O_2816,N_24957,N_24835);
xnor UO_2817 (O_2817,N_24757,N_24895);
and UO_2818 (O_2818,N_24772,N_24942);
and UO_2819 (O_2819,N_24818,N_24942);
and UO_2820 (O_2820,N_24991,N_24818);
xnor UO_2821 (O_2821,N_24784,N_24982);
nand UO_2822 (O_2822,N_24957,N_24994);
or UO_2823 (O_2823,N_24761,N_24828);
xnor UO_2824 (O_2824,N_24827,N_24777);
or UO_2825 (O_2825,N_24804,N_24950);
and UO_2826 (O_2826,N_24751,N_24836);
nor UO_2827 (O_2827,N_24807,N_24951);
nand UO_2828 (O_2828,N_24825,N_24967);
and UO_2829 (O_2829,N_24802,N_24939);
xor UO_2830 (O_2830,N_24869,N_24864);
nor UO_2831 (O_2831,N_24779,N_24885);
xnor UO_2832 (O_2832,N_24866,N_24977);
nand UO_2833 (O_2833,N_24789,N_24801);
xnor UO_2834 (O_2834,N_24907,N_24928);
nand UO_2835 (O_2835,N_24847,N_24938);
nor UO_2836 (O_2836,N_24827,N_24978);
xnor UO_2837 (O_2837,N_24952,N_24914);
xor UO_2838 (O_2838,N_24916,N_24967);
or UO_2839 (O_2839,N_24777,N_24992);
and UO_2840 (O_2840,N_24807,N_24780);
and UO_2841 (O_2841,N_24963,N_24902);
nor UO_2842 (O_2842,N_24805,N_24817);
or UO_2843 (O_2843,N_24868,N_24967);
xor UO_2844 (O_2844,N_24830,N_24979);
or UO_2845 (O_2845,N_24961,N_24904);
nor UO_2846 (O_2846,N_24973,N_24835);
or UO_2847 (O_2847,N_24962,N_24772);
and UO_2848 (O_2848,N_24866,N_24948);
nor UO_2849 (O_2849,N_24911,N_24891);
or UO_2850 (O_2850,N_24773,N_24921);
nor UO_2851 (O_2851,N_24832,N_24871);
xnor UO_2852 (O_2852,N_24990,N_24983);
nand UO_2853 (O_2853,N_24775,N_24848);
and UO_2854 (O_2854,N_24858,N_24955);
xor UO_2855 (O_2855,N_24766,N_24873);
nand UO_2856 (O_2856,N_24758,N_24995);
nor UO_2857 (O_2857,N_24816,N_24997);
nor UO_2858 (O_2858,N_24766,N_24942);
xor UO_2859 (O_2859,N_24863,N_24842);
nand UO_2860 (O_2860,N_24849,N_24987);
or UO_2861 (O_2861,N_24878,N_24839);
and UO_2862 (O_2862,N_24830,N_24821);
xor UO_2863 (O_2863,N_24971,N_24851);
nor UO_2864 (O_2864,N_24950,N_24796);
or UO_2865 (O_2865,N_24869,N_24856);
or UO_2866 (O_2866,N_24857,N_24759);
nand UO_2867 (O_2867,N_24899,N_24812);
or UO_2868 (O_2868,N_24987,N_24905);
nor UO_2869 (O_2869,N_24800,N_24878);
nand UO_2870 (O_2870,N_24901,N_24896);
and UO_2871 (O_2871,N_24756,N_24798);
nand UO_2872 (O_2872,N_24781,N_24797);
or UO_2873 (O_2873,N_24781,N_24947);
and UO_2874 (O_2874,N_24844,N_24881);
or UO_2875 (O_2875,N_24777,N_24966);
and UO_2876 (O_2876,N_24884,N_24946);
and UO_2877 (O_2877,N_24938,N_24870);
nand UO_2878 (O_2878,N_24943,N_24879);
nand UO_2879 (O_2879,N_24820,N_24896);
or UO_2880 (O_2880,N_24781,N_24750);
nand UO_2881 (O_2881,N_24793,N_24805);
or UO_2882 (O_2882,N_24993,N_24909);
nand UO_2883 (O_2883,N_24802,N_24840);
nand UO_2884 (O_2884,N_24960,N_24753);
nor UO_2885 (O_2885,N_24920,N_24962);
and UO_2886 (O_2886,N_24759,N_24842);
nor UO_2887 (O_2887,N_24776,N_24889);
xnor UO_2888 (O_2888,N_24826,N_24946);
nor UO_2889 (O_2889,N_24953,N_24865);
nor UO_2890 (O_2890,N_24863,N_24834);
or UO_2891 (O_2891,N_24785,N_24994);
nor UO_2892 (O_2892,N_24934,N_24914);
xor UO_2893 (O_2893,N_24839,N_24849);
and UO_2894 (O_2894,N_24956,N_24805);
xor UO_2895 (O_2895,N_24983,N_24794);
or UO_2896 (O_2896,N_24922,N_24905);
nor UO_2897 (O_2897,N_24928,N_24801);
nor UO_2898 (O_2898,N_24794,N_24790);
nor UO_2899 (O_2899,N_24832,N_24961);
nor UO_2900 (O_2900,N_24813,N_24806);
nand UO_2901 (O_2901,N_24815,N_24770);
nand UO_2902 (O_2902,N_24827,N_24818);
nor UO_2903 (O_2903,N_24824,N_24840);
nor UO_2904 (O_2904,N_24833,N_24943);
and UO_2905 (O_2905,N_24750,N_24930);
or UO_2906 (O_2906,N_24862,N_24907);
and UO_2907 (O_2907,N_24853,N_24932);
and UO_2908 (O_2908,N_24868,N_24832);
nor UO_2909 (O_2909,N_24850,N_24837);
and UO_2910 (O_2910,N_24793,N_24969);
nand UO_2911 (O_2911,N_24769,N_24889);
xnor UO_2912 (O_2912,N_24805,N_24804);
or UO_2913 (O_2913,N_24842,N_24772);
or UO_2914 (O_2914,N_24900,N_24917);
and UO_2915 (O_2915,N_24886,N_24849);
nand UO_2916 (O_2916,N_24845,N_24760);
nor UO_2917 (O_2917,N_24888,N_24787);
nand UO_2918 (O_2918,N_24751,N_24943);
nand UO_2919 (O_2919,N_24812,N_24928);
xnor UO_2920 (O_2920,N_24762,N_24988);
and UO_2921 (O_2921,N_24939,N_24889);
xor UO_2922 (O_2922,N_24938,N_24893);
or UO_2923 (O_2923,N_24873,N_24931);
or UO_2924 (O_2924,N_24845,N_24960);
or UO_2925 (O_2925,N_24876,N_24835);
nor UO_2926 (O_2926,N_24954,N_24845);
or UO_2927 (O_2927,N_24763,N_24766);
nand UO_2928 (O_2928,N_24823,N_24756);
nor UO_2929 (O_2929,N_24858,N_24907);
xor UO_2930 (O_2930,N_24897,N_24893);
or UO_2931 (O_2931,N_24936,N_24953);
and UO_2932 (O_2932,N_24788,N_24763);
nand UO_2933 (O_2933,N_24931,N_24765);
nor UO_2934 (O_2934,N_24868,N_24796);
nor UO_2935 (O_2935,N_24904,N_24983);
and UO_2936 (O_2936,N_24805,N_24757);
nand UO_2937 (O_2937,N_24941,N_24780);
xnor UO_2938 (O_2938,N_24872,N_24950);
nand UO_2939 (O_2939,N_24834,N_24762);
xnor UO_2940 (O_2940,N_24867,N_24907);
xnor UO_2941 (O_2941,N_24945,N_24906);
xor UO_2942 (O_2942,N_24949,N_24809);
nor UO_2943 (O_2943,N_24941,N_24825);
nor UO_2944 (O_2944,N_24876,N_24993);
or UO_2945 (O_2945,N_24999,N_24785);
nor UO_2946 (O_2946,N_24947,N_24929);
or UO_2947 (O_2947,N_24906,N_24978);
nor UO_2948 (O_2948,N_24858,N_24929);
or UO_2949 (O_2949,N_24876,N_24915);
or UO_2950 (O_2950,N_24970,N_24899);
xnor UO_2951 (O_2951,N_24786,N_24817);
and UO_2952 (O_2952,N_24825,N_24811);
and UO_2953 (O_2953,N_24974,N_24876);
nand UO_2954 (O_2954,N_24793,N_24788);
or UO_2955 (O_2955,N_24950,N_24894);
xnor UO_2956 (O_2956,N_24982,N_24944);
or UO_2957 (O_2957,N_24830,N_24802);
xor UO_2958 (O_2958,N_24925,N_24881);
nand UO_2959 (O_2959,N_24760,N_24936);
nor UO_2960 (O_2960,N_24804,N_24910);
nand UO_2961 (O_2961,N_24789,N_24912);
nand UO_2962 (O_2962,N_24824,N_24758);
xnor UO_2963 (O_2963,N_24995,N_24936);
nand UO_2964 (O_2964,N_24915,N_24989);
xnor UO_2965 (O_2965,N_24915,N_24887);
xor UO_2966 (O_2966,N_24896,N_24906);
nand UO_2967 (O_2967,N_24959,N_24907);
nor UO_2968 (O_2968,N_24940,N_24812);
or UO_2969 (O_2969,N_24959,N_24813);
xnor UO_2970 (O_2970,N_24974,N_24962);
and UO_2971 (O_2971,N_24816,N_24977);
or UO_2972 (O_2972,N_24855,N_24975);
nor UO_2973 (O_2973,N_24827,N_24844);
nand UO_2974 (O_2974,N_24835,N_24753);
nand UO_2975 (O_2975,N_24982,N_24924);
nand UO_2976 (O_2976,N_24977,N_24984);
xor UO_2977 (O_2977,N_24835,N_24879);
nor UO_2978 (O_2978,N_24983,N_24812);
nand UO_2979 (O_2979,N_24882,N_24871);
nand UO_2980 (O_2980,N_24928,N_24969);
and UO_2981 (O_2981,N_24907,N_24944);
nor UO_2982 (O_2982,N_24778,N_24915);
nand UO_2983 (O_2983,N_24776,N_24825);
or UO_2984 (O_2984,N_24942,N_24950);
and UO_2985 (O_2985,N_24798,N_24893);
xnor UO_2986 (O_2986,N_24801,N_24771);
xor UO_2987 (O_2987,N_24969,N_24976);
or UO_2988 (O_2988,N_24972,N_24850);
xnor UO_2989 (O_2989,N_24985,N_24773);
xor UO_2990 (O_2990,N_24938,N_24896);
and UO_2991 (O_2991,N_24860,N_24927);
or UO_2992 (O_2992,N_24992,N_24893);
nor UO_2993 (O_2993,N_24800,N_24998);
nor UO_2994 (O_2994,N_24913,N_24813);
and UO_2995 (O_2995,N_24807,N_24895);
nand UO_2996 (O_2996,N_24885,N_24816);
or UO_2997 (O_2997,N_24823,N_24980);
nor UO_2998 (O_2998,N_24822,N_24760);
or UO_2999 (O_2999,N_24892,N_24751);
endmodule