module basic_2000_20000_2500_10_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1093,In_1479);
nor U1 (N_1,In_1471,In_1758);
and U2 (N_2,In_804,In_335);
or U3 (N_3,In_692,In_1456);
nor U4 (N_4,In_664,In_729);
nand U5 (N_5,In_432,In_530);
or U6 (N_6,In_747,In_1344);
and U7 (N_7,In_1185,In_854);
and U8 (N_8,In_1882,In_737);
nand U9 (N_9,In_370,In_1929);
nand U10 (N_10,In_332,In_543);
nor U11 (N_11,In_1951,In_1794);
nand U12 (N_12,In_1740,In_888);
xnor U13 (N_13,In_589,In_436);
nor U14 (N_14,In_1457,In_1394);
nor U15 (N_15,In_1886,In_36);
or U16 (N_16,In_859,In_643);
nand U17 (N_17,In_1778,In_1950);
nand U18 (N_18,In_1139,In_1339);
nand U19 (N_19,In_608,In_241);
or U20 (N_20,In_306,In_27);
and U21 (N_21,In_455,In_886);
and U22 (N_22,In_1106,In_666);
xnor U23 (N_23,In_1572,In_333);
nand U24 (N_24,In_0,In_1698);
nand U25 (N_25,In_911,In_1591);
nand U26 (N_26,In_1253,In_1055);
and U27 (N_27,In_350,In_1648);
and U28 (N_28,In_388,In_1472);
nand U29 (N_29,In_1840,In_1984);
or U30 (N_30,In_959,In_1352);
nand U31 (N_31,In_1395,In_919);
nor U32 (N_32,In_529,In_1001);
xnor U33 (N_33,In_1205,In_305);
nand U34 (N_34,In_1030,In_1700);
and U35 (N_35,In_553,In_550);
and U36 (N_36,In_1904,In_1604);
xor U37 (N_37,In_1310,In_1076);
or U38 (N_38,In_825,In_1451);
and U39 (N_39,In_979,In_1616);
and U40 (N_40,In_1593,In_1252);
and U41 (N_41,In_938,In_978);
xor U42 (N_42,In_746,In_456);
nand U43 (N_43,In_1668,In_1598);
and U44 (N_44,In_1993,In_1420);
nand U45 (N_45,In_883,In_1008);
or U46 (N_46,In_1731,In_740);
nand U47 (N_47,In_1889,In_670);
or U48 (N_48,In_488,In_1866);
or U49 (N_49,In_185,In_1645);
nor U50 (N_50,In_1602,In_205);
xor U51 (N_51,In_472,In_743);
nand U52 (N_52,In_569,In_1192);
and U53 (N_53,In_1627,In_154);
and U54 (N_54,In_482,In_372);
xor U55 (N_55,In_1815,In_1034);
nand U56 (N_56,In_1974,In_1662);
nand U57 (N_57,In_1626,In_1266);
nor U58 (N_58,In_789,In_1169);
xnor U59 (N_59,In_114,In_1379);
and U60 (N_60,In_1982,In_940);
nor U61 (N_61,In_1547,In_1579);
nor U62 (N_62,In_1475,In_1697);
and U63 (N_63,In_1632,In_423);
and U64 (N_64,In_1194,In_1552);
nand U65 (N_65,In_1635,In_240);
nor U66 (N_66,In_1608,In_136);
and U67 (N_67,In_1224,In_540);
and U68 (N_68,In_1495,In_147);
nand U69 (N_69,In_1018,In_1070);
and U70 (N_70,In_1907,In_982);
or U71 (N_71,In_1002,In_866);
nor U72 (N_72,In_41,In_948);
or U73 (N_73,In_704,In_770);
and U74 (N_74,In_1198,In_1195);
nand U75 (N_75,In_312,In_1980);
and U76 (N_76,In_1784,In_95);
and U77 (N_77,In_1149,In_1745);
xor U78 (N_78,In_1998,In_447);
xnor U79 (N_79,In_1704,In_784);
nand U80 (N_80,In_239,In_1623);
nand U81 (N_81,In_25,In_12);
nor U82 (N_82,In_945,In_586);
xnor U83 (N_83,In_1927,In_646);
nand U84 (N_84,In_1611,In_1753);
nand U85 (N_85,In_385,In_431);
or U86 (N_86,In_212,In_1836);
nor U87 (N_87,In_709,In_578);
xor U88 (N_88,In_815,In_92);
nor U89 (N_89,In_444,In_62);
and U90 (N_90,In_1330,In_887);
nand U91 (N_91,In_435,In_1393);
nand U92 (N_92,In_951,In_590);
nor U93 (N_93,In_1959,In_1193);
nor U94 (N_94,In_930,In_1737);
and U95 (N_95,In_1268,In_823);
nor U96 (N_96,In_840,In_427);
xnor U97 (N_97,In_195,In_1426);
or U98 (N_98,In_1706,In_52);
or U99 (N_99,In_277,In_884);
or U100 (N_100,In_612,In_853);
or U101 (N_101,In_1213,In_725);
and U102 (N_102,In_1234,In_1090);
and U103 (N_103,In_268,In_227);
nand U104 (N_104,In_1216,In_899);
nor U105 (N_105,In_440,In_1518);
and U106 (N_106,In_1655,In_1082);
nor U107 (N_107,In_1481,In_649);
and U108 (N_108,In_1617,In_1414);
nand U109 (N_109,In_1750,In_1869);
nor U110 (N_110,In_1187,In_1003);
nor U111 (N_111,In_1883,In_1212);
and U112 (N_112,In_976,In_1497);
or U113 (N_113,In_123,In_1023);
nand U114 (N_114,In_572,In_871);
xor U115 (N_115,In_1690,In_1500);
or U116 (N_116,In_1621,In_399);
and U117 (N_117,In_603,In_1587);
xnor U118 (N_118,In_767,In_1735);
or U119 (N_119,In_741,In_426);
nand U120 (N_120,In_762,In_1845);
nand U121 (N_121,In_1658,In_921);
or U122 (N_122,In_1992,In_623);
xnor U123 (N_123,In_1669,In_1038);
xnor U124 (N_124,In_1743,In_1321);
and U125 (N_125,In_942,In_952);
and U126 (N_126,In_594,In_248);
nand U127 (N_127,In_11,In_857);
nor U128 (N_128,In_523,In_127);
nor U129 (N_129,In_1986,In_1484);
and U130 (N_130,In_1118,In_1359);
nand U131 (N_131,In_1351,In_960);
nand U132 (N_132,In_1926,In_1620);
or U133 (N_133,In_1120,In_330);
and U134 (N_134,In_1772,In_772);
xnor U135 (N_135,In_496,In_1249);
nand U136 (N_136,In_1649,In_1112);
nand U137 (N_137,In_1361,In_1200);
nor U138 (N_138,In_1806,In_1548);
or U139 (N_139,In_182,In_1583);
or U140 (N_140,In_1524,In_500);
nor U141 (N_141,In_499,In_562);
or U142 (N_142,In_410,In_1981);
nor U143 (N_143,In_882,In_953);
and U144 (N_144,In_1975,In_1808);
and U145 (N_145,In_975,In_476);
and U146 (N_146,In_1525,In_599);
or U147 (N_147,In_1117,In_1783);
nand U148 (N_148,In_336,In_779);
nand U149 (N_149,In_793,In_7);
nand U150 (N_150,In_1087,In_1970);
nor U151 (N_151,In_1837,In_1787);
nor U152 (N_152,In_9,In_687);
nand U153 (N_153,In_571,In_294);
or U154 (N_154,In_81,In_902);
nand U155 (N_155,In_1831,In_856);
and U156 (N_156,In_1862,In_1116);
or U157 (N_157,In_1629,In_491);
nand U158 (N_158,In_1368,In_1418);
xnor U159 (N_159,In_547,In_785);
or U160 (N_160,In_1546,In_61);
or U161 (N_161,In_1235,In_1086);
nor U162 (N_162,In_1651,In_1404);
and U163 (N_163,In_1461,In_1590);
and U164 (N_164,In_1757,In_880);
or U165 (N_165,In_1121,In_987);
or U166 (N_166,In_460,In_164);
nor U167 (N_167,In_1115,In_252);
and U168 (N_168,In_1191,In_1292);
or U169 (N_169,In_1222,In_568);
nor U170 (N_170,In_808,In_1782);
nor U171 (N_171,In_601,In_1133);
or U172 (N_172,In_1734,In_1720);
nand U173 (N_173,In_1014,In_255);
and U174 (N_174,In_1307,In_78);
nor U175 (N_175,In_282,In_364);
nand U176 (N_176,In_1453,In_1328);
or U177 (N_177,In_378,In_359);
nand U178 (N_178,In_107,In_573);
nor U179 (N_179,In_1920,In_1910);
and U180 (N_180,In_188,In_796);
xnor U181 (N_181,In_1853,In_821);
nor U182 (N_182,In_1505,In_108);
nor U183 (N_183,In_698,In_759);
or U184 (N_184,In_997,In_171);
nand U185 (N_185,In_820,In_1380);
xor U186 (N_186,In_1176,In_1802);
nand U187 (N_187,In_1966,In_727);
nor U188 (N_188,In_609,In_1541);
nor U189 (N_189,In_72,In_801);
or U190 (N_190,In_483,In_387);
nor U191 (N_191,In_29,In_1374);
or U192 (N_192,In_329,In_877);
nand U193 (N_193,In_1108,In_1719);
and U194 (N_194,In_818,In_84);
or U195 (N_195,In_858,In_146);
or U196 (N_196,In_77,In_1103);
nor U197 (N_197,In_102,In_1536);
nand U198 (N_198,In_1256,In_313);
nand U199 (N_199,In_106,In_1389);
or U200 (N_200,In_792,In_1857);
or U201 (N_201,In_520,In_990);
nor U202 (N_202,In_393,In_703);
nor U203 (N_203,In_1458,In_1146);
nor U204 (N_204,In_1065,In_627);
nor U205 (N_205,In_645,In_527);
or U206 (N_206,In_1932,In_1281);
and U207 (N_207,In_231,In_130);
nor U208 (N_208,In_844,In_705);
nor U209 (N_209,In_1941,In_973);
nand U210 (N_210,In_453,In_1375);
nand U211 (N_211,In_618,In_276);
or U212 (N_212,In_96,In_140);
xor U213 (N_213,In_1665,In_1282);
or U214 (N_214,In_860,In_1206);
nand U215 (N_215,In_629,In_1179);
nand U216 (N_216,In_1147,In_85);
nor U217 (N_217,In_383,In_1596);
nand U218 (N_218,In_1523,In_957);
and U219 (N_219,In_1040,In_802);
nor U220 (N_220,In_1860,In_1102);
or U221 (N_221,In_449,In_1708);
nor U222 (N_222,In_441,In_261);
or U223 (N_223,In_962,In_538);
or U224 (N_224,In_546,In_280);
and U225 (N_225,In_145,In_218);
nor U226 (N_226,In_728,In_1994);
nand U227 (N_227,In_234,In_1296);
nor U228 (N_228,In_655,In_824);
nand U229 (N_229,In_517,In_1677);
nor U230 (N_230,In_971,In_714);
nand U231 (N_231,In_69,In_1295);
nor U232 (N_232,In_1259,In_1263);
or U233 (N_233,In_1051,In_865);
nor U234 (N_234,In_1849,In_1835);
or U235 (N_235,In_1080,In_1721);
nand U236 (N_236,In_794,In_906);
nand U237 (N_237,In_237,In_1832);
nand U238 (N_238,In_903,In_774);
and U239 (N_239,In_912,In_1452);
nand U240 (N_240,In_531,In_376);
nor U241 (N_241,In_1371,In_1908);
and U242 (N_242,In_738,In_606);
and U243 (N_243,In_199,In_250);
and U244 (N_244,In_44,In_889);
nor U245 (N_245,In_838,In_1397);
and U246 (N_246,In_26,In_1672);
nor U247 (N_247,In_1696,In_1048);
nand U248 (N_248,In_309,In_157);
or U249 (N_249,In_1972,In_1531);
nor U250 (N_250,In_1534,In_137);
nor U251 (N_251,In_1843,In_300);
nand U252 (N_252,In_1124,In_1610);
or U253 (N_253,In_1699,In_1961);
nor U254 (N_254,In_461,In_1675);
nor U255 (N_255,In_833,In_1110);
or U256 (N_256,In_1245,In_56);
xor U257 (N_257,In_904,In_1279);
nor U258 (N_258,In_1299,In_551);
and U259 (N_259,In_1633,In_259);
or U260 (N_260,In_303,In_139);
or U261 (N_261,In_454,In_1983);
or U262 (N_262,In_1613,In_1791);
nor U263 (N_263,In_907,In_730);
nand U264 (N_264,In_718,In_1558);
and U265 (N_265,In_1449,In_356);
or U266 (N_266,In_1607,In_1269);
xor U267 (N_267,In_65,In_1006);
nand U268 (N_268,In_1807,In_1277);
nand U269 (N_269,In_1965,In_1923);
nand U270 (N_270,In_1214,In_289);
nand U271 (N_271,In_870,In_1370);
nor U272 (N_272,In_1248,In_225);
nor U273 (N_273,In_260,In_661);
xor U274 (N_274,In_1431,In_1417);
and U275 (N_275,In_293,In_323);
and U276 (N_276,In_122,In_1542);
and U277 (N_277,In_54,In_99);
or U278 (N_278,In_894,In_1510);
nand U279 (N_279,In_1968,In_473);
nand U280 (N_280,In_1202,In_638);
and U281 (N_281,In_120,In_2);
nor U282 (N_282,In_315,In_1016);
or U283 (N_283,In_94,In_658);
or U284 (N_284,In_1298,In_34);
or U285 (N_285,In_626,In_1842);
and U286 (N_286,In_209,In_466);
and U287 (N_287,In_1997,In_893);
nand U288 (N_288,In_1841,In_428);
nor U289 (N_289,In_1094,In_885);
nor U290 (N_290,In_1010,In_545);
and U291 (N_291,In_1334,In_691);
nor U292 (N_292,In_1798,In_1673);
and U293 (N_293,In_272,In_873);
or U294 (N_294,In_344,In_1874);
and U295 (N_295,In_1877,In_660);
or U296 (N_296,In_284,In_1976);
nand U297 (N_297,In_295,In_701);
nand U298 (N_298,In_1319,In_55);
or U299 (N_299,In_999,In_1520);
nand U300 (N_300,In_1682,In_1428);
and U301 (N_301,In_1589,In_1811);
xnor U302 (N_302,In_148,In_1508);
nand U303 (N_303,In_1501,In_339);
and U304 (N_304,In_192,In_1340);
xnor U305 (N_305,In_519,In_1575);
or U306 (N_306,In_1775,In_696);
and U307 (N_307,In_1795,In_434);
xor U308 (N_308,In_1346,In_712);
and U309 (N_309,In_595,In_1032);
nor U310 (N_310,In_686,In_262);
nor U311 (N_311,In_1262,In_1438);
nor U312 (N_312,In_1095,In_565);
nand U313 (N_313,In_1163,In_849);
nor U314 (N_314,In_1494,In_1289);
and U315 (N_315,In_963,In_1412);
nand U316 (N_316,In_757,In_1027);
or U317 (N_317,In_1460,In_809);
xor U318 (N_318,In_1223,In_1180);
nor U319 (N_319,In_672,In_1887);
nand U320 (N_320,In_841,In_1915);
nor U321 (N_321,In_1151,In_47);
and U322 (N_322,In_32,In_1683);
nor U323 (N_323,In_1123,In_1056);
xor U324 (N_324,In_1448,In_694);
nor U325 (N_325,In_1868,In_1160);
or U326 (N_326,In_1780,In_1674);
nand U327 (N_327,In_1320,In_509);
and U328 (N_328,In_533,In_699);
nor U329 (N_329,In_1209,In_1844);
nor U330 (N_330,In_1396,In_1897);
nor U331 (N_331,In_1278,In_909);
or U332 (N_332,In_377,In_862);
or U333 (N_333,In_819,In_1741);
nand U334 (N_334,In_949,In_1324);
nor U335 (N_335,In_813,In_1063);
nor U336 (N_336,In_1891,In_582);
or U337 (N_337,In_731,In_1852);
and U338 (N_338,In_70,In_579);
and U339 (N_339,In_1640,In_1364);
nand U340 (N_340,In_352,In_715);
nand U341 (N_341,In_177,In_1401);
nand U342 (N_342,In_574,In_1432);
and U343 (N_343,In_1423,In_258);
and U344 (N_344,In_1440,In_1430);
or U345 (N_345,In_1145,In_211);
and U346 (N_346,In_1990,In_17);
nor U347 (N_347,In_150,In_1688);
and U348 (N_348,In_524,In_1689);
nand U349 (N_349,In_141,In_1411);
xnor U350 (N_350,In_1876,In_20);
nor U351 (N_351,In_156,In_1301);
xor U352 (N_352,In_1846,In_634);
nor U353 (N_353,In_810,In_1391);
and U354 (N_354,In_630,In_722);
nand U355 (N_355,In_1636,In_1964);
nor U356 (N_356,In_1353,In_155);
and U357 (N_357,In_1378,In_98);
nand U358 (N_358,In_285,In_1348);
and U359 (N_359,In_181,In_935);
and U360 (N_360,In_944,In_318);
nand U361 (N_361,In_394,In_1469);
or U362 (N_362,In_1527,In_1126);
nor U363 (N_363,In_104,In_1267);
and U364 (N_364,In_1365,In_1820);
or U365 (N_365,In_468,In_1517);
and U366 (N_366,In_1751,In_166);
or U367 (N_367,In_1712,In_901);
and U368 (N_368,In_790,In_816);
nor U369 (N_369,In_1302,In_682);
and U370 (N_370,In_671,In_763);
and U371 (N_371,In_659,In_1482);
nand U372 (N_372,In_652,In_924);
or U373 (N_373,In_1854,In_1530);
xor U374 (N_374,In_1563,In_1347);
or U375 (N_375,In_1503,In_898);
or U376 (N_376,In_1555,In_561);
xor U377 (N_377,In_213,In_1250);
or U378 (N_378,In_970,In_1088);
or U379 (N_379,In_908,In_220);
xor U380 (N_380,In_1489,In_995);
nor U381 (N_381,In_1382,In_1363);
and U382 (N_382,In_1229,In_63);
nor U383 (N_383,In_442,In_1512);
or U384 (N_384,In_619,In_1275);
or U385 (N_385,In_642,In_265);
or U386 (N_386,In_679,In_560);
nand U387 (N_387,In_1424,In_950);
and U388 (N_388,In_1387,In_1233);
or U389 (N_389,In_402,In_274);
nand U390 (N_390,In_557,In_97);
nand U391 (N_391,In_1614,In_507);
xor U392 (N_392,In_839,In_1599);
or U393 (N_393,In_494,In_1276);
or U394 (N_394,In_1099,In_187);
and U395 (N_395,In_23,In_644);
nor U396 (N_396,In_929,In_878);
xnor U397 (N_397,In_799,In_1019);
or U398 (N_398,In_1476,In_628);
nor U399 (N_399,In_768,In_100);
and U400 (N_400,In_1366,In_577);
nor U401 (N_401,In_283,In_125);
or U402 (N_402,In_1297,In_1089);
and U403 (N_403,In_1153,In_1748);
and U404 (N_404,In_173,In_319);
nand U405 (N_405,In_787,In_1814);
nand U406 (N_406,In_1800,In_1464);
and U407 (N_407,In_783,In_286);
nor U408 (N_408,In_1178,In_1024);
xor U409 (N_409,In_467,In_144);
and U410 (N_410,In_1367,In_302);
nand U411 (N_411,In_1190,In_693);
and U412 (N_412,In_1119,In_1963);
nand U413 (N_413,In_1101,In_1083);
nand U414 (N_414,In_1122,In_710);
nor U415 (N_415,In_28,In_826);
or U416 (N_416,In_1634,In_1935);
and U417 (N_417,In_832,In_1075);
and U418 (N_418,In_269,In_1601);
nand U419 (N_419,In_1046,In_484);
nand U420 (N_420,In_87,In_310);
or U421 (N_421,In_1399,In_1141);
and U422 (N_422,In_1226,In_1052);
nand U423 (N_423,In_1666,In_707);
or U424 (N_424,In_1933,In_1676);
xnor U425 (N_425,In_937,In_1989);
nor U426 (N_426,In_1726,In_1144);
or U427 (N_427,In_503,In_625);
nand U428 (N_428,In_414,In_1477);
and U429 (N_429,In_1025,In_477);
nand U430 (N_430,In_4,In_674);
and U431 (N_431,In_1261,In_1906);
and U432 (N_432,In_1136,In_943);
or U433 (N_433,In_614,In_475);
nor U434 (N_434,In_851,In_1447);
and U435 (N_435,In_1433,In_521);
or U436 (N_436,In_1071,In_15);
nand U437 (N_437,In_724,In_1474);
and U438 (N_438,In_1540,In_1532);
and U439 (N_439,In_189,In_129);
nand U440 (N_440,In_162,In_993);
xor U441 (N_441,In_396,In_992);
or U442 (N_442,In_1755,In_1012);
or U443 (N_443,In_1204,In_867);
nand U444 (N_444,In_1559,In_1100);
nor U445 (N_445,In_1188,In_233);
and U446 (N_446,In_13,In_1855);
and U447 (N_447,In_1381,In_57);
and U448 (N_448,In_1005,In_1954);
or U449 (N_449,In_489,In_965);
nand U450 (N_450,In_1343,In_109);
or U451 (N_451,In_900,In_1437);
or U452 (N_452,In_1739,In_1333);
and U453 (N_453,In_716,In_662);
nand U454 (N_454,In_1054,In_1659);
and U455 (N_455,In_1560,In_1392);
and U456 (N_456,In_1577,In_1174);
nor U457 (N_457,In_235,In_534);
and U458 (N_458,In_24,In_1148);
nor U459 (N_459,In_1529,In_417);
and U460 (N_460,In_695,In_621);
nor U461 (N_461,In_1528,In_1667);
and U462 (N_462,In_1053,In_1728);
and U463 (N_463,In_721,In_1917);
or U464 (N_464,In_1158,In_1356);
nor U465 (N_465,In_548,In_864);
or U466 (N_466,In_1656,In_287);
nand U467 (N_467,In_1884,In_1044);
nor U468 (N_468,In_505,In_822);
and U469 (N_469,In_1097,In_689);
or U470 (N_470,In_1492,In_1550);
xor U471 (N_471,In_1826,In_46);
nand U472 (N_472,In_381,In_1839);
nand U473 (N_473,In_1013,In_184);
nand U474 (N_474,In_602,In_91);
nor U475 (N_475,In_1488,In_827);
nor U476 (N_476,In_204,In_281);
and U477 (N_477,In_1419,In_528);
xor U478 (N_478,In_1823,In_1624);
or U479 (N_479,In_271,In_765);
nor U480 (N_480,In_321,In_1561);
nor U481 (N_481,In_665,In_1759);
or U482 (N_482,In_1225,In_1043);
nor U483 (N_483,In_640,In_1684);
nor U484 (N_484,In_169,In_115);
or U485 (N_485,In_1221,In_1723);
or U486 (N_486,In_279,In_1092);
and U487 (N_487,In_1628,In_1916);
and U488 (N_488,In_1638,In_490);
or U489 (N_489,In_1196,In_67);
nand U490 (N_490,In_739,In_913);
and U491 (N_491,In_1322,In_1405);
or U492 (N_492,In_1554,In_1864);
nor U493 (N_493,In_868,In_1805);
nand U494 (N_494,In_744,In_1317);
xor U495 (N_495,In_984,In_736);
nor U496 (N_496,In_134,In_1900);
nand U497 (N_497,In_201,In_1872);
nand U498 (N_498,In_1402,In_411);
nand U499 (N_499,In_1435,In_1422);
and U500 (N_500,In_1127,In_40);
nand U501 (N_501,In_1217,In_717);
nand U502 (N_502,In_508,In_392);
nor U503 (N_503,In_1037,In_1445);
and U504 (N_504,In_539,In_863);
nand U505 (N_505,In_723,In_761);
nand U506 (N_506,In_1967,In_345);
nor U507 (N_507,In_1625,In_1265);
and U508 (N_508,In_1165,In_1057);
nor U509 (N_509,In_776,In_1663);
or U510 (N_510,In_366,In_1777);
or U511 (N_511,In_1637,In_760);
nor U512 (N_512,In_135,In_536);
nand U513 (N_513,In_64,In_928);
or U514 (N_514,In_941,In_834);
or U515 (N_515,In_914,In_1851);
nand U516 (N_516,In_931,In_1239);
and U517 (N_517,In_617,In_439);
nor U518 (N_518,In_1588,In_170);
or U519 (N_519,In_327,In_256);
or U520 (N_520,In_121,In_373);
or U521 (N_521,In_1863,In_947);
nor U522 (N_522,In_358,In_143);
nor U523 (N_523,In_1557,In_245);
xnor U524 (N_524,In_126,In_734);
nor U525 (N_525,In_648,In_1171);
nor U526 (N_526,In_1442,In_570);
nand U527 (N_527,In_934,In_238);
and U528 (N_528,In_409,In_1770);
nor U529 (N_529,In_1930,In_554);
nor U530 (N_530,In_925,In_298);
or U531 (N_531,In_1164,In_273);
and U532 (N_532,In_35,In_1166);
nor U533 (N_533,In_1254,In_1824);
or U534 (N_534,In_492,In_1571);
nor U535 (N_535,In_684,In_264);
nor U536 (N_536,In_478,In_420);
or U537 (N_537,In_1280,In_1064);
nand U538 (N_538,In_457,In_1388);
and U539 (N_539,In_1098,In_1376);
and U540 (N_540,In_1944,In_1600);
nor U541 (N_541,In_88,In_1246);
and U542 (N_542,In_79,In_175);
or U543 (N_543,In_1940,In_1644);
or U544 (N_544,In_1881,In_487);
nor U545 (N_545,In_632,In_3);
nand U546 (N_546,In_133,In_588);
or U547 (N_547,In_549,In_1237);
nand U548 (N_548,In_1979,In_958);
nor U549 (N_549,In_1504,In_1231);
and U550 (N_550,In_879,In_1184);
nor U551 (N_551,In_1513,In_1274);
nand U552 (N_552,In_5,In_1208);
nand U553 (N_553,In_1303,In_1385);
or U554 (N_554,In_1756,In_1969);
nor U555 (N_555,In_1227,In_656);
nand U556 (N_556,In_1797,In_516);
or U557 (N_557,In_994,In_1228);
or U558 (N_558,In_430,In_1308);
and U559 (N_559,In_1140,In_386);
and U560 (N_560,In_1809,In_1861);
or U561 (N_561,In_1948,In_480);
and U562 (N_562,In_346,In_1175);
or U563 (N_563,In_90,In_1776);
or U564 (N_564,In_1349,In_397);
nand U565 (N_565,In_1186,In_76);
nand U566 (N_566,In_153,In_1793);
and U567 (N_567,In_1362,In_663);
xor U568 (N_568,In_1605,In_1714);
nor U569 (N_569,In_1850,In_416);
and U570 (N_570,In_117,In_1924);
nor U571 (N_571,In_732,In_343);
or U572 (N_572,In_1074,In_1009);
nor U573 (N_573,In_31,In_1870);
and U574 (N_574,In_1358,In_916);
and U575 (N_575,In_1183,In_1403);
nor U576 (N_576,In_814,In_675);
and U577 (N_577,In_795,In_1270);
nor U578 (N_578,In_308,In_450);
nand U579 (N_579,In_847,In_750);
xor U580 (N_580,In_362,In_1020);
nand U581 (N_581,In_964,In_1657);
or U582 (N_582,In_1441,In_607);
xnor U583 (N_583,In_1670,In_1957);
or U584 (N_584,In_1818,In_1060);
nor U585 (N_585,In_685,In_391);
nand U586 (N_586,In_812,In_168);
xor U587 (N_587,In_1498,In_425);
and U588 (N_588,In_526,In_1332);
or U589 (N_589,In_1733,In_611);
nor U590 (N_590,In_1425,In_1565);
nand U591 (N_591,In_1710,In_668);
and U592 (N_592,In_1316,In_1511);
nand U593 (N_593,In_1985,In_1996);
or U594 (N_594,In_459,In_592);
or U595 (N_595,In_518,In_502);
or U596 (N_596,In_1913,In_1473);
nand U597 (N_597,In_955,In_1902);
nor U598 (N_598,In_563,In_1096);
and U599 (N_599,In_555,In_1746);
and U600 (N_600,In_1409,In_216);
or U601 (N_601,In_116,In_68);
and U602 (N_602,In_1152,In_405);
nand U603 (N_603,In_180,In_1161);
nor U604 (N_604,In_933,In_830);
and U605 (N_605,In_998,In_542);
and U606 (N_606,In_221,In_249);
nor U607 (N_607,In_1515,In_1764);
nor U608 (N_608,In_836,In_1300);
and U609 (N_609,In_733,In_1952);
xor U610 (N_610,In_1491,In_1360);
and U611 (N_611,In_1875,In_1580);
and U612 (N_612,In_633,In_1566);
and U613 (N_613,In_486,In_497);
nor U614 (N_614,In_1283,In_1687);
or U615 (N_615,In_236,In_1537);
nand U616 (N_616,In_232,In_374);
nand U617 (N_617,In_1643,In_1413);
and U618 (N_618,In_1905,In_1847);
nand U619 (N_619,In_535,In_254);
nor U620 (N_620,In_1896,In_1914);
or U621 (N_621,In_178,In_82);
or U622 (N_622,In_415,In_1181);
xor U623 (N_623,In_631,In_564);
nor U624 (N_624,In_1129,In_1724);
nand U625 (N_625,In_101,In_1134);
and U626 (N_626,In_1812,In_320);
nand U627 (N_627,In_1960,In_855);
xor U628 (N_628,In_16,In_1871);
nor U629 (N_629,In_1264,In_412);
nand U630 (N_630,In_1919,In_1691);
or U631 (N_631,In_989,In_708);
and U632 (N_632,In_1199,In_465);
nor U633 (N_633,In_753,In_1526);
nand U634 (N_634,In_1582,In_75);
nor U635 (N_635,In_406,In_290);
and U636 (N_636,In_700,In_980);
or U637 (N_637,In_1466,In_1592);
or U638 (N_638,In_1285,In_1955);
and U639 (N_639,In_1945,In_591);
nand U640 (N_640,In_504,In_1912);
nor U641 (N_641,In_1230,In_1732);
and U642 (N_642,In_1722,In_1893);
xnor U643 (N_643,In_1066,In_1062);
nor U644 (N_644,In_1830,In_1949);
and U645 (N_645,In_1692,In_197);
or U646 (N_646,In_1068,In_1671);
or U647 (N_647,In_342,In_1921);
or U648 (N_648,In_1177,In_86);
xor U649 (N_649,In_230,In_1829);
nor U650 (N_650,In_522,In_1031);
xor U651 (N_651,In_961,In_207);
nand U652 (N_652,In_1067,In_74);
nand U653 (N_653,In_1765,In_1584);
nand U654 (N_654,In_1315,In_1744);
nand U655 (N_655,In_226,In_537);
nand U656 (N_656,In_920,In_755);
nor U657 (N_657,In_365,In_10);
or U658 (N_658,In_1061,In_861);
and U659 (N_659,In_1958,In_1693);
xor U660 (N_660,In_1789,In_749);
or U661 (N_661,In_706,In_1618);
nor U662 (N_662,In_1664,In_1077);
or U663 (N_663,In_890,In_1335);
nor U664 (N_664,In_1,In_1899);
and U665 (N_665,In_647,In_1130);
and U666 (N_666,In_1774,In_1091);
or U667 (N_667,In_217,In_895);
nand U668 (N_668,In_1567,In_1128);
or U669 (N_669,In_1415,In_1991);
nor U670 (N_670,In_1509,In_1939);
nor U671 (N_671,In_1258,In_683);
and U672 (N_672,In_58,In_1465);
or U673 (N_673,In_161,In_1398);
xor U674 (N_674,In_1942,In_326);
xor U675 (N_675,In_118,In_1416);
nand U676 (N_676,In_193,In_1232);
or U677 (N_677,In_316,In_382);
nor U678 (N_678,In_202,In_1408);
nor U679 (N_679,In_932,In_1729);
nor U680 (N_680,In_1170,In_1312);
nand U681 (N_681,In_196,In_1042);
or U682 (N_682,In_30,In_510);
nor U683 (N_683,In_1154,In_915);
nor U684 (N_684,In_458,In_1521);
or U685 (N_685,In_1015,In_1779);
nand U686 (N_686,In_1922,In_702);
and U687 (N_687,In_1903,In_636);
xnor U688 (N_688,In_93,In_1597);
nor U689 (N_689,In_1790,In_463);
nand U690 (N_690,In_1619,In_1257);
nand U691 (N_691,In_1490,In_1715);
and U692 (N_692,In_1111,In_331);
or U693 (N_693,In_243,In_341);
and U694 (N_694,In_48,In_1803);
xnor U695 (N_695,In_1995,In_1182);
nor U696 (N_696,In_918,In_224);
nor U697 (N_697,In_576,In_969);
nor U698 (N_698,In_1342,In_1142);
nor U699 (N_699,In_375,In_748);
or U700 (N_700,In_142,In_1543);
xor U701 (N_701,In_1962,In_1859);
nand U702 (N_702,In_720,In_1218);
or U703 (N_703,In_1045,In_1036);
nand U704 (N_704,In_443,In_1240);
xor U705 (N_705,In_1338,In_1026);
nor U706 (N_706,In_1702,In_1928);
nor U707 (N_707,In_452,In_613);
or U708 (N_708,In_1455,In_1742);
or U709 (N_709,In_59,In_1646);
or U710 (N_710,In_1821,In_317);
and U711 (N_711,In_798,In_1241);
or U712 (N_712,In_1576,In_673);
or U713 (N_713,In_1211,In_1858);
nor U714 (N_714,In_690,In_1642);
nor U715 (N_715,In_278,In_1131);
nor U716 (N_716,In_1892,In_288);
and U717 (N_717,In_1443,In_1946);
xnor U718 (N_718,In_1827,In_1207);
nand U719 (N_719,In_1502,In_575);
nand U720 (N_720,In_1242,In_1306);
nand U721 (N_721,In_1647,In_513);
or U722 (N_722,In_1943,In_881);
nor U723 (N_723,In_1586,In_1470);
nand U724 (N_724,In_917,In_996);
xor U725 (N_725,In_1819,In_437);
nand U726 (N_726,In_775,In_1848);
and U727 (N_727,In_429,In_669);
nand U728 (N_728,In_805,In_581);
or U729 (N_729,In_1107,In_596);
nor U730 (N_730,In_384,In_113);
nor U731 (N_731,In_1386,In_357);
and U732 (N_732,In_1918,In_1763);
and U733 (N_733,In_719,In_905);
nor U734 (N_734,In_263,In_469);
or U735 (N_735,In_1890,In_1000);
and U736 (N_736,In_892,In_1653);
nor U737 (N_737,In_138,In_1384);
nor U738 (N_738,In_1041,In_1717);
nor U739 (N_739,In_641,In_1694);
nand U740 (N_740,In_846,In_266);
nor U741 (N_741,In_307,In_1695);
and U742 (N_742,In_1595,In_1911);
or U743 (N_743,In_1769,In_1654);
nor U744 (N_744,In_1125,In_756);
nor U745 (N_745,In_848,In_742);
and U746 (N_746,In_936,In_111);
and U747 (N_747,In_1804,In_1377);
and U748 (N_748,In_270,In_493);
or U749 (N_749,In_831,In_1084);
nand U750 (N_750,In_1318,In_433);
or U751 (N_751,In_80,In_1788);
or U752 (N_752,In_872,In_1834);
xor U753 (N_753,In_347,In_1459);
or U754 (N_754,In_1516,In_132);
nand U755 (N_755,In_1894,In_251);
and U756 (N_756,In_1813,In_128);
nand U757 (N_757,In_1817,In_51);
or U758 (N_758,In_446,In_1007);
and U759 (N_759,In_349,In_778);
nor U760 (N_760,In_1022,In_1796);
and U761 (N_761,In_676,In_837);
nand U762 (N_762,In_1585,In_781);
nor U763 (N_763,In_680,In_754);
or U764 (N_764,In_1017,In_1109);
xnor U765 (N_765,In_325,In_1641);
nor U766 (N_766,In_605,In_33);
and U767 (N_767,In_1711,In_1493);
xnor U768 (N_768,In_1773,In_1701);
nand U769 (N_769,In_348,In_1159);
xor U770 (N_770,In_1243,In_1716);
nor U771 (N_771,In_165,In_1244);
nand U772 (N_772,In_780,In_407);
nand U773 (N_773,In_292,In_751);
nand U774 (N_774,In_1327,In_1999);
nand U775 (N_775,In_1369,In_1685);
nor U776 (N_776,In_1215,In_1357);
nor U777 (N_777,In_1661,In_1873);
nor U778 (N_778,In_1081,In_1931);
and U779 (N_779,In_361,In_1569);
and U780 (N_780,In_807,In_119);
and U781 (N_781,In_1703,In_610);
nand U782 (N_782,In_1485,In_8);
or U783 (N_783,In_1167,In_584);
or U784 (N_784,In_1522,In_1936);
and U785 (N_785,In_1004,In_194);
xor U786 (N_786,In_923,In_1507);
or U787 (N_787,In_1311,In_1947);
nand U788 (N_788,In_1898,In_215);
or U789 (N_789,In_1885,In_1828);
nand U790 (N_790,In_559,In_1201);
xnor U791 (N_791,In_445,In_1568);
nor U792 (N_792,In_1436,In_1519);
and U793 (N_793,In_131,In_471);
nor U794 (N_794,In_37,In_1029);
xor U795 (N_795,In_1514,In_1938);
and U796 (N_796,In_615,In_758);
or U797 (N_797,In_875,In_967);
or U798 (N_798,In_1162,In_1681);
nand U799 (N_799,In_985,In_511);
nor U800 (N_800,In_991,In_1157);
and U801 (N_801,In_580,In_296);
nand U802 (N_802,In_620,In_1762);
nor U803 (N_803,In_1168,In_797);
nand U804 (N_804,In_1467,In_1273);
or U805 (N_805,In_1761,In_83);
or U806 (N_806,In_208,In_1909);
xnor U807 (N_807,In_1331,In_1747);
and U808 (N_808,In_922,In_939);
or U809 (N_809,In_635,In_1901);
nand U810 (N_810,In_481,In_291);
nor U811 (N_811,In_1480,In_874);
or U812 (N_812,In_1973,In_1792);
or U813 (N_813,In_360,In_328);
xnor U814 (N_814,In_1113,In_541);
nand U815 (N_815,In_438,In_788);
or U816 (N_816,In_1203,In_1236);
or U817 (N_817,In_1350,In_1035);
nor U818 (N_818,In_791,In_1615);
nand U819 (N_819,In_1287,In_1679);
nand U820 (N_820,In_593,In_421);
or U821 (N_821,In_424,In_1730);
xor U822 (N_822,In_1345,In_1172);
nand U823 (N_823,In_337,In_512);
nor U824 (N_824,In_558,In_498);
nand U825 (N_825,In_1650,In_966);
nor U826 (N_826,In_124,In_1533);
or U827 (N_827,In_1538,In_567);
nand U828 (N_828,In_1603,In_1462);
xnor U829 (N_829,In_650,In_1059);
nand U830 (N_830,In_474,In_203);
nor U831 (N_831,In_6,In_198);
nor U832 (N_832,In_222,In_624);
and U833 (N_833,In_1400,In_1446);
or U834 (N_834,In_681,In_1573);
nor U835 (N_835,In_850,In_1173);
nor U836 (N_836,In_956,In_1838);
nor U837 (N_837,In_1718,In_828);
nor U838 (N_838,In_103,In_651);
nor U839 (N_839,In_1544,In_1801);
or U840 (N_840,In_334,In_408);
nand U841 (N_841,In_404,In_267);
nor U842 (N_842,In_1372,In_566);
nand U843 (N_843,In_556,In_1556);
nor U844 (N_844,In_1132,In_1768);
and U845 (N_845,In_1606,In_598);
and U846 (N_846,In_803,In_544);
and U847 (N_847,In_1197,In_1879);
and U848 (N_848,In_299,In_1639);
and U849 (N_849,In_604,In_1049);
nand U850 (N_850,In_773,In_1150);
xnor U851 (N_851,In_1407,In_1652);
nor U852 (N_852,In_1078,In_1570);
nand U853 (N_853,In_1079,In_151);
xnor U854 (N_854,In_1271,In_1325);
nand U855 (N_855,In_1630,In_174);
or U856 (N_856,In_45,In_1156);
nor U857 (N_857,In_413,In_418);
and U858 (N_858,In_448,In_1294);
xnor U859 (N_859,In_244,In_229);
or U860 (N_860,In_1535,In_1260);
nor U861 (N_861,In_786,In_1373);
nand U862 (N_862,In_1578,In_422);
and U863 (N_863,In_1705,In_1925);
and U864 (N_864,In_974,In_191);
and U865 (N_865,In_876,In_1786);
nor U866 (N_866,In_1073,In_1736);
nor U867 (N_867,In_1799,In_369);
or U868 (N_868,In_246,In_1410);
or U869 (N_869,In_1336,In_1255);
or U870 (N_870,In_713,In_401);
or U871 (N_871,In_843,In_379);
nor U872 (N_872,In_228,In_1304);
and U873 (N_873,In_112,In_1506);
and U874 (N_874,In_752,In_66);
nand U875 (N_875,In_811,In_1766);
nand U876 (N_876,In_1314,In_371);
nor U877 (N_877,In_1104,In_1988);
xnor U878 (N_878,In_653,In_1895);
nor U879 (N_879,In_1155,In_159);
xor U880 (N_880,In_1594,In_1880);
nor U881 (N_881,In_1977,In_1888);
or U882 (N_882,In_1463,In_829);
or U883 (N_883,In_89,In_735);
nand U884 (N_884,In_1220,In_1551);
xnor U885 (N_885,In_43,In_1867);
or U886 (N_886,In_1956,In_322);
and U887 (N_887,In_1678,In_354);
or U888 (N_888,In_73,In_800);
xnor U889 (N_889,In_304,In_1251);
xnor U890 (N_890,In_1953,In_1286);
nand U891 (N_891,In_400,In_766);
or U892 (N_892,In_14,In_977);
nand U893 (N_893,In_19,In_1069);
and U894 (N_894,In_485,In_340);
and U895 (N_895,In_60,In_1421);
or U896 (N_896,In_1137,In_183);
xor U897 (N_897,In_1707,In_637);
or U898 (N_898,In_891,In_110);
or U899 (N_899,In_1468,In_1272);
nand U900 (N_900,In_1326,In_50);
xor U901 (N_901,In_1033,In_697);
xnor U902 (N_902,In_552,In_1021);
nand U903 (N_903,In_1293,In_1427);
nand U904 (N_904,In_1865,In_464);
or U905 (N_905,In_1028,In_1383);
or U906 (N_906,In_247,In_1406);
and U907 (N_907,In_1749,In_1138);
and U908 (N_908,In_1496,In_910);
nand U909 (N_909,In_1738,In_1329);
or U910 (N_910,In_223,In_1754);
xnor U911 (N_911,In_71,In_1355);
xor U912 (N_912,In_22,In_389);
and U913 (N_913,In_1309,In_1454);
xor U914 (N_914,In_654,In_219);
or U915 (N_915,In_1219,In_395);
nand U916 (N_916,In_506,In_1058);
nor U917 (N_917,In_1039,In_968);
or U918 (N_918,In_927,In_764);
xor U919 (N_919,In_257,In_21);
and U920 (N_920,In_896,In_1499);
nand U921 (N_921,In_1631,In_18);
and U922 (N_922,In_1781,In_190);
nand U923 (N_923,In_470,In_1553);
xor U924 (N_924,In_380,In_179);
and U925 (N_925,In_817,In_1483);
nand U926 (N_926,In_1011,In_1760);
nand U927 (N_927,In_585,In_1767);
nor U928 (N_928,In_1609,In_160);
nand U929 (N_929,In_1135,In_1210);
nor U930 (N_930,In_1622,In_1612);
and U931 (N_931,In_53,In_954);
and U932 (N_932,In_1539,In_1833);
xor U933 (N_933,In_988,In_176);
or U934 (N_934,In_42,In_324);
nor U935 (N_935,In_1752,In_616);
nor U936 (N_936,In_842,In_451);
nand U937 (N_937,In_351,In_1050);
nor U938 (N_938,In_771,In_587);
nor U939 (N_939,In_1987,In_338);
and U940 (N_940,In_186,In_1247);
nand U941 (N_941,In_1305,In_301);
nand U942 (N_942,In_242,In_1478);
and U943 (N_943,In_1450,In_639);
or U944 (N_944,In_1686,In_745);
xor U945 (N_945,In_525,In_200);
or U946 (N_946,In_253,In_1978);
or U947 (N_947,In_214,In_210);
and U948 (N_948,In_622,In_677);
nand U949 (N_949,In_1713,In_1878);
nand U950 (N_950,In_769,In_1284);
or U951 (N_951,In_172,In_419);
or U952 (N_952,In_158,In_297);
nor U953 (N_953,In_1816,In_845);
nor U954 (N_954,In_1444,In_983);
nand U955 (N_955,In_1549,In_600);
or U956 (N_956,In_206,In_398);
nor U957 (N_957,In_390,In_462);
and U958 (N_958,In_1323,In_1771);
nor U959 (N_959,In_1934,In_1238);
nor U960 (N_960,In_972,In_355);
nand U961 (N_961,In_1487,In_1937);
nand U962 (N_962,In_105,In_1143);
and U963 (N_963,In_532,In_1725);
nand U964 (N_964,In_1545,In_1439);
nand U965 (N_965,In_368,In_946);
and U966 (N_966,In_1114,In_1856);
and U967 (N_967,In_501,In_1810);
nand U968 (N_968,In_926,In_1313);
nand U969 (N_969,In_986,In_1291);
nor U970 (N_970,In_49,In_1047);
and U971 (N_971,In_678,In_149);
nand U972 (N_972,In_1574,In_495);
and U973 (N_973,In_403,In_1288);
and U974 (N_974,In_367,In_1105);
and U975 (N_975,In_583,In_657);
nand U976 (N_976,In_667,In_869);
nand U977 (N_977,In_835,In_726);
and U978 (N_978,In_1341,In_1680);
and U979 (N_979,In_1825,In_1429);
nor U980 (N_980,In_515,In_167);
or U981 (N_981,In_163,In_688);
and U982 (N_982,In_1660,In_981);
nor U983 (N_983,In_353,In_1562);
nand U984 (N_984,In_1486,In_711);
and U985 (N_985,In_39,In_479);
nor U986 (N_986,In_363,In_1354);
nor U987 (N_987,In_152,In_597);
nor U988 (N_988,In_1434,In_1337);
nand U989 (N_989,In_275,In_1072);
and U990 (N_990,In_1727,In_1709);
and U991 (N_991,In_1290,In_514);
and U992 (N_992,In_1822,In_852);
and U993 (N_993,In_782,In_1581);
and U994 (N_994,In_777,In_1785);
and U995 (N_995,In_1564,In_806);
nand U996 (N_996,In_314,In_38);
or U997 (N_997,In_1390,In_1189);
nor U998 (N_998,In_1971,In_897);
nor U999 (N_999,In_311,In_1085);
and U1000 (N_1000,In_1840,In_64);
nand U1001 (N_1001,In_1193,In_379);
nor U1002 (N_1002,In_205,In_181);
xor U1003 (N_1003,In_1176,In_1780);
or U1004 (N_1004,In_1748,In_742);
nor U1005 (N_1005,In_1021,In_1404);
and U1006 (N_1006,In_653,In_1576);
xnor U1007 (N_1007,In_1738,In_249);
nand U1008 (N_1008,In_1033,In_1226);
nand U1009 (N_1009,In_574,In_360);
and U1010 (N_1010,In_862,In_1920);
nand U1011 (N_1011,In_1321,In_1438);
or U1012 (N_1012,In_1582,In_516);
xor U1013 (N_1013,In_959,In_359);
xor U1014 (N_1014,In_981,In_1262);
nor U1015 (N_1015,In_915,In_162);
and U1016 (N_1016,In_498,In_871);
nor U1017 (N_1017,In_199,In_626);
nand U1018 (N_1018,In_1073,In_152);
or U1019 (N_1019,In_246,In_1275);
nor U1020 (N_1020,In_1170,In_488);
and U1021 (N_1021,In_1214,In_1924);
xnor U1022 (N_1022,In_1014,In_1303);
or U1023 (N_1023,In_1211,In_603);
or U1024 (N_1024,In_500,In_952);
or U1025 (N_1025,In_1718,In_837);
xnor U1026 (N_1026,In_616,In_222);
nor U1027 (N_1027,In_1687,In_423);
nand U1028 (N_1028,In_1807,In_1292);
or U1029 (N_1029,In_775,In_876);
and U1030 (N_1030,In_1695,In_1514);
or U1031 (N_1031,In_1973,In_1507);
nor U1032 (N_1032,In_1791,In_1206);
nand U1033 (N_1033,In_1952,In_241);
nor U1034 (N_1034,In_194,In_1601);
nand U1035 (N_1035,In_1770,In_1450);
nor U1036 (N_1036,In_1463,In_45);
xnor U1037 (N_1037,In_519,In_851);
and U1038 (N_1038,In_846,In_637);
or U1039 (N_1039,In_190,In_294);
nand U1040 (N_1040,In_82,In_884);
nand U1041 (N_1041,In_1738,In_1141);
nor U1042 (N_1042,In_689,In_590);
nor U1043 (N_1043,In_332,In_693);
and U1044 (N_1044,In_662,In_907);
and U1045 (N_1045,In_42,In_1717);
or U1046 (N_1046,In_1411,In_1268);
or U1047 (N_1047,In_90,In_990);
or U1048 (N_1048,In_214,In_235);
or U1049 (N_1049,In_697,In_19);
and U1050 (N_1050,In_1498,In_133);
or U1051 (N_1051,In_1653,In_1931);
nor U1052 (N_1052,In_1797,In_369);
and U1053 (N_1053,In_904,In_977);
or U1054 (N_1054,In_1480,In_974);
nor U1055 (N_1055,In_619,In_300);
or U1056 (N_1056,In_1809,In_412);
xnor U1057 (N_1057,In_850,In_1379);
nor U1058 (N_1058,In_1402,In_1336);
nor U1059 (N_1059,In_1652,In_212);
and U1060 (N_1060,In_843,In_743);
and U1061 (N_1061,In_1139,In_1189);
and U1062 (N_1062,In_1951,In_1749);
or U1063 (N_1063,In_1581,In_243);
nand U1064 (N_1064,In_1503,In_1381);
or U1065 (N_1065,In_1126,In_259);
or U1066 (N_1066,In_1890,In_587);
nor U1067 (N_1067,In_249,In_619);
or U1068 (N_1068,In_1395,In_1998);
xnor U1069 (N_1069,In_1864,In_1904);
or U1070 (N_1070,In_1216,In_1645);
xnor U1071 (N_1071,In_1706,In_1266);
nor U1072 (N_1072,In_256,In_66);
nor U1073 (N_1073,In_491,In_1686);
or U1074 (N_1074,In_322,In_146);
nor U1075 (N_1075,In_1975,In_1155);
nand U1076 (N_1076,In_241,In_717);
nand U1077 (N_1077,In_797,In_1950);
nor U1078 (N_1078,In_439,In_849);
xor U1079 (N_1079,In_1990,In_846);
nor U1080 (N_1080,In_367,In_1918);
nor U1081 (N_1081,In_1056,In_463);
nor U1082 (N_1082,In_1211,In_751);
nand U1083 (N_1083,In_1922,In_176);
and U1084 (N_1084,In_1266,In_592);
or U1085 (N_1085,In_895,In_1113);
xor U1086 (N_1086,In_1564,In_148);
nor U1087 (N_1087,In_539,In_1109);
and U1088 (N_1088,In_1251,In_1215);
and U1089 (N_1089,In_782,In_950);
nand U1090 (N_1090,In_1938,In_1220);
or U1091 (N_1091,In_791,In_712);
nand U1092 (N_1092,In_693,In_1408);
and U1093 (N_1093,In_695,In_1701);
and U1094 (N_1094,In_643,In_714);
nand U1095 (N_1095,In_894,In_629);
nand U1096 (N_1096,In_361,In_883);
and U1097 (N_1097,In_1184,In_123);
nor U1098 (N_1098,In_1896,In_234);
nor U1099 (N_1099,In_666,In_1989);
nand U1100 (N_1100,In_46,In_203);
nand U1101 (N_1101,In_529,In_406);
nand U1102 (N_1102,In_1004,In_1193);
and U1103 (N_1103,In_873,In_191);
xor U1104 (N_1104,In_1281,In_1218);
nor U1105 (N_1105,In_519,In_947);
and U1106 (N_1106,In_611,In_255);
xor U1107 (N_1107,In_1599,In_1031);
nand U1108 (N_1108,In_1453,In_475);
or U1109 (N_1109,In_917,In_313);
or U1110 (N_1110,In_1670,In_89);
nor U1111 (N_1111,In_1535,In_334);
xor U1112 (N_1112,In_1994,In_346);
xor U1113 (N_1113,In_170,In_1486);
nand U1114 (N_1114,In_1559,In_1532);
nor U1115 (N_1115,In_672,In_653);
nand U1116 (N_1116,In_1568,In_1017);
and U1117 (N_1117,In_308,In_1224);
nor U1118 (N_1118,In_756,In_1750);
xor U1119 (N_1119,In_1554,In_209);
or U1120 (N_1120,In_692,In_1019);
nor U1121 (N_1121,In_1103,In_1368);
nor U1122 (N_1122,In_379,In_286);
nor U1123 (N_1123,In_541,In_1971);
nand U1124 (N_1124,In_799,In_316);
or U1125 (N_1125,In_1370,In_59);
nand U1126 (N_1126,In_599,In_375);
and U1127 (N_1127,In_582,In_242);
nand U1128 (N_1128,In_528,In_1568);
and U1129 (N_1129,In_115,In_634);
and U1130 (N_1130,In_1829,In_1070);
nand U1131 (N_1131,In_1827,In_1197);
nand U1132 (N_1132,In_1946,In_1387);
xor U1133 (N_1133,In_770,In_1303);
or U1134 (N_1134,In_1044,In_784);
nor U1135 (N_1135,In_919,In_130);
and U1136 (N_1136,In_662,In_890);
or U1137 (N_1137,In_1125,In_841);
nor U1138 (N_1138,In_541,In_1461);
and U1139 (N_1139,In_188,In_1364);
nor U1140 (N_1140,In_244,In_18);
xnor U1141 (N_1141,In_875,In_137);
or U1142 (N_1142,In_489,In_1513);
or U1143 (N_1143,In_1679,In_711);
and U1144 (N_1144,In_1420,In_1833);
nand U1145 (N_1145,In_315,In_1468);
xor U1146 (N_1146,In_112,In_1372);
nor U1147 (N_1147,In_1017,In_586);
nand U1148 (N_1148,In_927,In_755);
or U1149 (N_1149,In_390,In_513);
or U1150 (N_1150,In_1067,In_1078);
or U1151 (N_1151,In_994,In_1054);
or U1152 (N_1152,In_1763,In_1578);
nand U1153 (N_1153,In_1653,In_964);
and U1154 (N_1154,In_1264,In_1868);
or U1155 (N_1155,In_1973,In_1609);
nand U1156 (N_1156,In_875,In_1645);
xor U1157 (N_1157,In_1943,In_393);
nand U1158 (N_1158,In_1578,In_1869);
nor U1159 (N_1159,In_1176,In_1864);
xor U1160 (N_1160,In_1703,In_162);
nor U1161 (N_1161,In_1928,In_457);
and U1162 (N_1162,In_1435,In_247);
or U1163 (N_1163,In_1359,In_1273);
nor U1164 (N_1164,In_1405,In_1036);
nand U1165 (N_1165,In_1364,In_761);
nor U1166 (N_1166,In_1821,In_672);
or U1167 (N_1167,In_41,In_1191);
nand U1168 (N_1168,In_264,In_1931);
and U1169 (N_1169,In_919,In_937);
nor U1170 (N_1170,In_1062,In_109);
and U1171 (N_1171,In_5,In_201);
or U1172 (N_1172,In_727,In_1071);
or U1173 (N_1173,In_332,In_269);
or U1174 (N_1174,In_1327,In_258);
and U1175 (N_1175,In_1739,In_456);
nand U1176 (N_1176,In_1448,In_351);
and U1177 (N_1177,In_1261,In_1884);
and U1178 (N_1178,In_692,In_1724);
or U1179 (N_1179,In_173,In_1166);
and U1180 (N_1180,In_94,In_545);
and U1181 (N_1181,In_728,In_466);
nand U1182 (N_1182,In_1899,In_603);
nor U1183 (N_1183,In_535,In_514);
nand U1184 (N_1184,In_1358,In_421);
nand U1185 (N_1185,In_1286,In_212);
nand U1186 (N_1186,In_411,In_1893);
nor U1187 (N_1187,In_671,In_1602);
nor U1188 (N_1188,In_1990,In_595);
or U1189 (N_1189,In_263,In_244);
nor U1190 (N_1190,In_551,In_427);
nor U1191 (N_1191,In_846,In_1128);
or U1192 (N_1192,In_1507,In_224);
and U1193 (N_1193,In_1696,In_1396);
xnor U1194 (N_1194,In_630,In_57);
and U1195 (N_1195,In_883,In_895);
or U1196 (N_1196,In_1368,In_1998);
and U1197 (N_1197,In_837,In_1919);
or U1198 (N_1198,In_1337,In_1125);
and U1199 (N_1199,In_975,In_168);
nor U1200 (N_1200,In_1620,In_9);
nor U1201 (N_1201,In_1875,In_855);
or U1202 (N_1202,In_227,In_408);
nand U1203 (N_1203,In_1826,In_159);
or U1204 (N_1204,In_1248,In_1664);
nand U1205 (N_1205,In_18,In_705);
or U1206 (N_1206,In_780,In_574);
or U1207 (N_1207,In_172,In_1117);
nor U1208 (N_1208,In_195,In_1087);
nor U1209 (N_1209,In_698,In_679);
nand U1210 (N_1210,In_1885,In_289);
or U1211 (N_1211,In_708,In_1604);
nor U1212 (N_1212,In_298,In_1151);
xnor U1213 (N_1213,In_815,In_1493);
or U1214 (N_1214,In_878,In_356);
nor U1215 (N_1215,In_1782,In_173);
nand U1216 (N_1216,In_1266,In_198);
xor U1217 (N_1217,In_100,In_375);
nand U1218 (N_1218,In_1461,In_927);
or U1219 (N_1219,In_1070,In_365);
and U1220 (N_1220,In_689,In_1665);
nor U1221 (N_1221,In_1725,In_1064);
or U1222 (N_1222,In_294,In_1336);
nand U1223 (N_1223,In_1579,In_1451);
nand U1224 (N_1224,In_1630,In_400);
nand U1225 (N_1225,In_208,In_687);
nor U1226 (N_1226,In_516,In_1482);
nand U1227 (N_1227,In_186,In_1339);
nor U1228 (N_1228,In_18,In_644);
and U1229 (N_1229,In_1694,In_149);
or U1230 (N_1230,In_680,In_347);
xor U1231 (N_1231,In_23,In_737);
nand U1232 (N_1232,In_1565,In_499);
nor U1233 (N_1233,In_1824,In_1784);
and U1234 (N_1234,In_1212,In_1214);
or U1235 (N_1235,In_54,In_671);
nor U1236 (N_1236,In_141,In_1324);
nand U1237 (N_1237,In_738,In_926);
nand U1238 (N_1238,In_854,In_901);
xnor U1239 (N_1239,In_1039,In_803);
and U1240 (N_1240,In_114,In_1421);
nand U1241 (N_1241,In_1807,In_1699);
and U1242 (N_1242,In_44,In_1276);
nand U1243 (N_1243,In_1511,In_550);
or U1244 (N_1244,In_609,In_1920);
or U1245 (N_1245,In_521,In_1528);
nor U1246 (N_1246,In_177,In_1045);
or U1247 (N_1247,In_115,In_4);
nor U1248 (N_1248,In_1675,In_764);
or U1249 (N_1249,In_1930,In_985);
xnor U1250 (N_1250,In_414,In_1736);
or U1251 (N_1251,In_370,In_231);
xnor U1252 (N_1252,In_1080,In_117);
and U1253 (N_1253,In_1250,In_1962);
xor U1254 (N_1254,In_506,In_1716);
nand U1255 (N_1255,In_20,In_1590);
or U1256 (N_1256,In_939,In_405);
nand U1257 (N_1257,In_1594,In_403);
xor U1258 (N_1258,In_907,In_547);
or U1259 (N_1259,In_833,In_914);
or U1260 (N_1260,In_1494,In_991);
nor U1261 (N_1261,In_711,In_670);
and U1262 (N_1262,In_1482,In_1388);
nand U1263 (N_1263,In_802,In_1432);
nor U1264 (N_1264,In_1343,In_1700);
nand U1265 (N_1265,In_1525,In_1103);
nand U1266 (N_1266,In_1742,In_1673);
nor U1267 (N_1267,In_819,In_1733);
nor U1268 (N_1268,In_1829,In_1482);
or U1269 (N_1269,In_935,In_1974);
nor U1270 (N_1270,In_717,In_1267);
and U1271 (N_1271,In_602,In_287);
nor U1272 (N_1272,In_113,In_1121);
or U1273 (N_1273,In_1673,In_1196);
nand U1274 (N_1274,In_891,In_533);
nand U1275 (N_1275,In_1701,In_617);
or U1276 (N_1276,In_731,In_390);
nand U1277 (N_1277,In_699,In_921);
xnor U1278 (N_1278,In_981,In_1357);
nand U1279 (N_1279,In_1137,In_766);
and U1280 (N_1280,In_174,In_1392);
or U1281 (N_1281,In_644,In_1238);
and U1282 (N_1282,In_530,In_894);
nor U1283 (N_1283,In_1288,In_1052);
and U1284 (N_1284,In_897,In_998);
or U1285 (N_1285,In_219,In_185);
nand U1286 (N_1286,In_838,In_1860);
nand U1287 (N_1287,In_1021,In_329);
nand U1288 (N_1288,In_1704,In_1212);
nor U1289 (N_1289,In_1036,In_1418);
nor U1290 (N_1290,In_1199,In_1078);
nand U1291 (N_1291,In_1870,In_799);
nand U1292 (N_1292,In_590,In_1860);
nor U1293 (N_1293,In_1666,In_191);
or U1294 (N_1294,In_284,In_165);
and U1295 (N_1295,In_1454,In_1230);
xor U1296 (N_1296,In_656,In_857);
and U1297 (N_1297,In_980,In_974);
nand U1298 (N_1298,In_115,In_1712);
nand U1299 (N_1299,In_617,In_1788);
and U1300 (N_1300,In_1990,In_1917);
and U1301 (N_1301,In_336,In_1683);
nand U1302 (N_1302,In_1767,In_1963);
nand U1303 (N_1303,In_723,In_1366);
and U1304 (N_1304,In_995,In_1481);
or U1305 (N_1305,In_796,In_1351);
and U1306 (N_1306,In_1123,In_1317);
and U1307 (N_1307,In_1541,In_221);
nand U1308 (N_1308,In_671,In_1994);
nand U1309 (N_1309,In_507,In_1092);
and U1310 (N_1310,In_16,In_1213);
nand U1311 (N_1311,In_569,In_1201);
xnor U1312 (N_1312,In_1110,In_489);
and U1313 (N_1313,In_1198,In_1387);
or U1314 (N_1314,In_425,In_200);
and U1315 (N_1315,In_1266,In_1196);
xnor U1316 (N_1316,In_1306,In_318);
nand U1317 (N_1317,In_929,In_458);
nand U1318 (N_1318,In_405,In_1604);
or U1319 (N_1319,In_1719,In_711);
or U1320 (N_1320,In_1992,In_503);
and U1321 (N_1321,In_849,In_1849);
or U1322 (N_1322,In_1255,In_148);
nor U1323 (N_1323,In_1227,In_563);
or U1324 (N_1324,In_660,In_278);
nand U1325 (N_1325,In_1657,In_875);
nand U1326 (N_1326,In_1463,In_1079);
or U1327 (N_1327,In_143,In_1181);
and U1328 (N_1328,In_311,In_805);
nor U1329 (N_1329,In_1364,In_1540);
nor U1330 (N_1330,In_1588,In_1751);
xor U1331 (N_1331,In_1485,In_728);
nor U1332 (N_1332,In_124,In_1306);
nand U1333 (N_1333,In_1888,In_1550);
nor U1334 (N_1334,In_776,In_1320);
or U1335 (N_1335,In_1262,In_435);
and U1336 (N_1336,In_455,In_406);
nand U1337 (N_1337,In_1235,In_1056);
or U1338 (N_1338,In_389,In_325);
nand U1339 (N_1339,In_147,In_174);
nor U1340 (N_1340,In_193,In_518);
nand U1341 (N_1341,In_1503,In_77);
or U1342 (N_1342,In_344,In_713);
nand U1343 (N_1343,In_663,In_518);
nor U1344 (N_1344,In_1384,In_57);
and U1345 (N_1345,In_361,In_1726);
nand U1346 (N_1346,In_1138,In_714);
xnor U1347 (N_1347,In_827,In_1642);
nand U1348 (N_1348,In_622,In_159);
or U1349 (N_1349,In_399,In_1783);
nor U1350 (N_1350,In_1226,In_1593);
or U1351 (N_1351,In_898,In_1715);
nor U1352 (N_1352,In_1762,In_738);
nor U1353 (N_1353,In_1006,In_1467);
and U1354 (N_1354,In_710,In_1186);
nand U1355 (N_1355,In_1393,In_1272);
and U1356 (N_1356,In_697,In_91);
nor U1357 (N_1357,In_1554,In_585);
nand U1358 (N_1358,In_180,In_168);
nor U1359 (N_1359,In_1219,In_1723);
or U1360 (N_1360,In_1241,In_825);
nor U1361 (N_1361,In_1166,In_521);
and U1362 (N_1362,In_138,In_1472);
nand U1363 (N_1363,In_1145,In_654);
or U1364 (N_1364,In_606,In_376);
nor U1365 (N_1365,In_1753,In_1961);
xor U1366 (N_1366,In_1046,In_714);
xor U1367 (N_1367,In_450,In_778);
and U1368 (N_1368,In_1801,In_1082);
nand U1369 (N_1369,In_83,In_351);
nand U1370 (N_1370,In_1797,In_1162);
or U1371 (N_1371,In_824,In_609);
nor U1372 (N_1372,In_1358,In_1371);
or U1373 (N_1373,In_1601,In_1802);
or U1374 (N_1374,In_1583,In_1348);
nor U1375 (N_1375,In_1430,In_1561);
xnor U1376 (N_1376,In_1408,In_432);
nand U1377 (N_1377,In_860,In_1651);
or U1378 (N_1378,In_1428,In_1056);
nand U1379 (N_1379,In_1603,In_634);
nand U1380 (N_1380,In_693,In_1055);
nor U1381 (N_1381,In_307,In_1502);
and U1382 (N_1382,In_8,In_417);
or U1383 (N_1383,In_1546,In_1251);
xor U1384 (N_1384,In_492,In_52);
and U1385 (N_1385,In_654,In_402);
nor U1386 (N_1386,In_1416,In_1739);
nand U1387 (N_1387,In_217,In_649);
nor U1388 (N_1388,In_978,In_628);
and U1389 (N_1389,In_842,In_1824);
nand U1390 (N_1390,In_1550,In_197);
nor U1391 (N_1391,In_947,In_1442);
nand U1392 (N_1392,In_745,In_1718);
nor U1393 (N_1393,In_1347,In_358);
nand U1394 (N_1394,In_533,In_1883);
or U1395 (N_1395,In_507,In_154);
nand U1396 (N_1396,In_341,In_533);
nand U1397 (N_1397,In_1241,In_593);
or U1398 (N_1398,In_1064,In_119);
or U1399 (N_1399,In_545,In_1761);
or U1400 (N_1400,In_628,In_1089);
nor U1401 (N_1401,In_377,In_1330);
nor U1402 (N_1402,In_1418,In_1038);
nor U1403 (N_1403,In_502,In_389);
and U1404 (N_1404,In_1596,In_754);
xnor U1405 (N_1405,In_664,In_1962);
and U1406 (N_1406,In_483,In_1606);
nand U1407 (N_1407,In_189,In_764);
xnor U1408 (N_1408,In_1297,In_754);
and U1409 (N_1409,In_903,In_1102);
and U1410 (N_1410,In_341,In_1294);
nand U1411 (N_1411,In_957,In_1682);
or U1412 (N_1412,In_63,In_356);
nor U1413 (N_1413,In_299,In_960);
nand U1414 (N_1414,In_1137,In_1473);
or U1415 (N_1415,In_1846,In_115);
nor U1416 (N_1416,In_1805,In_770);
nor U1417 (N_1417,In_1796,In_195);
and U1418 (N_1418,In_658,In_1740);
nand U1419 (N_1419,In_1392,In_1448);
or U1420 (N_1420,In_1589,In_771);
or U1421 (N_1421,In_276,In_42);
nor U1422 (N_1422,In_1814,In_1380);
and U1423 (N_1423,In_1296,In_1104);
and U1424 (N_1424,In_1355,In_658);
nor U1425 (N_1425,In_362,In_404);
nor U1426 (N_1426,In_1264,In_597);
or U1427 (N_1427,In_1437,In_281);
xnor U1428 (N_1428,In_1658,In_1043);
or U1429 (N_1429,In_332,In_49);
nand U1430 (N_1430,In_622,In_688);
nand U1431 (N_1431,In_1242,In_332);
nand U1432 (N_1432,In_1769,In_1373);
xnor U1433 (N_1433,In_1215,In_674);
or U1434 (N_1434,In_1961,In_1737);
nor U1435 (N_1435,In_1305,In_350);
and U1436 (N_1436,In_154,In_1746);
and U1437 (N_1437,In_12,In_569);
or U1438 (N_1438,In_107,In_884);
or U1439 (N_1439,In_1755,In_1903);
or U1440 (N_1440,In_1664,In_758);
nand U1441 (N_1441,In_1175,In_1201);
nand U1442 (N_1442,In_1017,In_1043);
or U1443 (N_1443,In_1205,In_243);
or U1444 (N_1444,In_1389,In_1218);
nor U1445 (N_1445,In_920,In_1914);
nand U1446 (N_1446,In_1893,In_1934);
nand U1447 (N_1447,In_384,In_1038);
xnor U1448 (N_1448,In_1056,In_1418);
xor U1449 (N_1449,In_1297,In_1145);
nor U1450 (N_1450,In_1865,In_1936);
nor U1451 (N_1451,In_1668,In_1662);
and U1452 (N_1452,In_747,In_1486);
nor U1453 (N_1453,In_1576,In_460);
or U1454 (N_1454,In_1315,In_1510);
nand U1455 (N_1455,In_834,In_270);
nor U1456 (N_1456,In_1644,In_1643);
nor U1457 (N_1457,In_210,In_165);
nand U1458 (N_1458,In_14,In_1643);
and U1459 (N_1459,In_1472,In_1654);
or U1460 (N_1460,In_1929,In_225);
or U1461 (N_1461,In_602,In_355);
and U1462 (N_1462,In_374,In_1027);
xor U1463 (N_1463,In_1516,In_1920);
or U1464 (N_1464,In_66,In_16);
and U1465 (N_1465,In_783,In_182);
nand U1466 (N_1466,In_1777,In_1927);
or U1467 (N_1467,In_1267,In_562);
nand U1468 (N_1468,In_1377,In_556);
nor U1469 (N_1469,In_326,In_1023);
or U1470 (N_1470,In_933,In_517);
and U1471 (N_1471,In_526,In_1710);
nor U1472 (N_1472,In_1314,In_335);
xor U1473 (N_1473,In_599,In_1159);
nand U1474 (N_1474,In_1891,In_1739);
nor U1475 (N_1475,In_646,In_1837);
nand U1476 (N_1476,In_1291,In_1850);
and U1477 (N_1477,In_1579,In_171);
or U1478 (N_1478,In_573,In_615);
or U1479 (N_1479,In_1737,In_625);
or U1480 (N_1480,In_1944,In_374);
or U1481 (N_1481,In_1212,In_269);
nor U1482 (N_1482,In_948,In_1878);
nand U1483 (N_1483,In_1513,In_1313);
and U1484 (N_1484,In_1967,In_1988);
nor U1485 (N_1485,In_546,In_729);
nor U1486 (N_1486,In_561,In_362);
nor U1487 (N_1487,In_553,In_1323);
xnor U1488 (N_1488,In_37,In_911);
and U1489 (N_1489,In_778,In_786);
nand U1490 (N_1490,In_95,In_503);
or U1491 (N_1491,In_178,In_1962);
and U1492 (N_1492,In_218,In_1967);
or U1493 (N_1493,In_632,In_1272);
nand U1494 (N_1494,In_1159,In_1223);
nand U1495 (N_1495,In_1016,In_1116);
and U1496 (N_1496,In_446,In_1512);
or U1497 (N_1497,In_1668,In_1026);
and U1498 (N_1498,In_653,In_212);
and U1499 (N_1499,In_1510,In_1472);
nor U1500 (N_1500,In_316,In_1171);
nand U1501 (N_1501,In_185,In_1530);
nand U1502 (N_1502,In_451,In_1955);
and U1503 (N_1503,In_918,In_213);
nand U1504 (N_1504,In_767,In_85);
and U1505 (N_1505,In_1987,In_1622);
or U1506 (N_1506,In_1962,In_1111);
nor U1507 (N_1507,In_135,In_1159);
nand U1508 (N_1508,In_670,In_809);
or U1509 (N_1509,In_1012,In_1196);
nand U1510 (N_1510,In_534,In_1469);
and U1511 (N_1511,In_121,In_183);
and U1512 (N_1512,In_859,In_757);
nor U1513 (N_1513,In_897,In_702);
xnor U1514 (N_1514,In_1512,In_927);
and U1515 (N_1515,In_1361,In_751);
xor U1516 (N_1516,In_520,In_1274);
nor U1517 (N_1517,In_636,In_751);
nor U1518 (N_1518,In_296,In_1925);
nand U1519 (N_1519,In_337,In_55);
nand U1520 (N_1520,In_1881,In_1852);
nand U1521 (N_1521,In_869,In_1872);
nor U1522 (N_1522,In_1120,In_284);
nor U1523 (N_1523,In_152,In_1008);
nor U1524 (N_1524,In_1616,In_1040);
xor U1525 (N_1525,In_1766,In_368);
nor U1526 (N_1526,In_57,In_1726);
nor U1527 (N_1527,In_698,In_128);
xor U1528 (N_1528,In_1631,In_211);
and U1529 (N_1529,In_531,In_1326);
nand U1530 (N_1530,In_1760,In_157);
xor U1531 (N_1531,In_1258,In_633);
nor U1532 (N_1532,In_217,In_1043);
or U1533 (N_1533,In_699,In_1726);
or U1534 (N_1534,In_1912,In_795);
and U1535 (N_1535,In_1429,In_1942);
xor U1536 (N_1536,In_172,In_179);
nor U1537 (N_1537,In_1423,In_1064);
nand U1538 (N_1538,In_1571,In_137);
nand U1539 (N_1539,In_1179,In_153);
or U1540 (N_1540,In_83,In_1388);
nor U1541 (N_1541,In_1704,In_802);
nand U1542 (N_1542,In_869,In_42);
xor U1543 (N_1543,In_987,In_1212);
and U1544 (N_1544,In_1770,In_519);
xor U1545 (N_1545,In_1524,In_1152);
nor U1546 (N_1546,In_1260,In_1915);
or U1547 (N_1547,In_135,In_1153);
nor U1548 (N_1548,In_1060,In_339);
nor U1549 (N_1549,In_1002,In_1285);
and U1550 (N_1550,In_1083,In_922);
or U1551 (N_1551,In_1117,In_1163);
nand U1552 (N_1552,In_1193,In_1168);
xor U1553 (N_1553,In_1723,In_60);
or U1554 (N_1554,In_305,In_1266);
nor U1555 (N_1555,In_1046,In_886);
and U1556 (N_1556,In_1400,In_432);
nand U1557 (N_1557,In_86,In_932);
and U1558 (N_1558,In_1611,In_1767);
nand U1559 (N_1559,In_1010,In_1846);
and U1560 (N_1560,In_897,In_1206);
nand U1561 (N_1561,In_828,In_1874);
nand U1562 (N_1562,In_1959,In_1497);
or U1563 (N_1563,In_1828,In_576);
nand U1564 (N_1564,In_486,In_1326);
nor U1565 (N_1565,In_1632,In_1532);
or U1566 (N_1566,In_349,In_745);
nor U1567 (N_1567,In_1318,In_821);
nand U1568 (N_1568,In_1522,In_995);
and U1569 (N_1569,In_51,In_1319);
nor U1570 (N_1570,In_613,In_987);
nand U1571 (N_1571,In_1771,In_110);
nor U1572 (N_1572,In_553,In_401);
nand U1573 (N_1573,In_1464,In_836);
nor U1574 (N_1574,In_1810,In_938);
nor U1575 (N_1575,In_1713,In_706);
or U1576 (N_1576,In_153,In_888);
or U1577 (N_1577,In_1292,In_5);
and U1578 (N_1578,In_332,In_630);
nand U1579 (N_1579,In_583,In_586);
or U1580 (N_1580,In_1025,In_211);
nand U1581 (N_1581,In_1337,In_1515);
and U1582 (N_1582,In_788,In_517);
xor U1583 (N_1583,In_674,In_1252);
nor U1584 (N_1584,In_1686,In_489);
or U1585 (N_1585,In_513,In_218);
or U1586 (N_1586,In_1972,In_705);
nor U1587 (N_1587,In_1538,In_382);
and U1588 (N_1588,In_1502,In_1755);
and U1589 (N_1589,In_1817,In_1033);
nor U1590 (N_1590,In_1022,In_627);
or U1591 (N_1591,In_1586,In_1049);
nor U1592 (N_1592,In_539,In_876);
nor U1593 (N_1593,In_25,In_990);
or U1594 (N_1594,In_1678,In_1644);
nor U1595 (N_1595,In_992,In_1767);
nand U1596 (N_1596,In_1075,In_450);
or U1597 (N_1597,In_958,In_613);
and U1598 (N_1598,In_17,In_1844);
and U1599 (N_1599,In_1972,In_1104);
and U1600 (N_1600,In_832,In_42);
xor U1601 (N_1601,In_1687,In_1822);
or U1602 (N_1602,In_1907,In_825);
and U1603 (N_1603,In_1977,In_1835);
nand U1604 (N_1604,In_998,In_8);
and U1605 (N_1605,In_422,In_35);
and U1606 (N_1606,In_508,In_236);
and U1607 (N_1607,In_902,In_1820);
and U1608 (N_1608,In_1597,In_101);
xnor U1609 (N_1609,In_536,In_1192);
and U1610 (N_1610,In_1309,In_1320);
or U1611 (N_1611,In_1019,In_1417);
xnor U1612 (N_1612,In_1312,In_365);
and U1613 (N_1613,In_930,In_842);
nor U1614 (N_1614,In_841,In_492);
nand U1615 (N_1615,In_437,In_1228);
or U1616 (N_1616,In_719,In_385);
nand U1617 (N_1617,In_1410,In_253);
xnor U1618 (N_1618,In_1987,In_90);
nor U1619 (N_1619,In_696,In_824);
nand U1620 (N_1620,In_543,In_707);
nand U1621 (N_1621,In_128,In_1538);
or U1622 (N_1622,In_1312,In_1566);
and U1623 (N_1623,In_481,In_1187);
and U1624 (N_1624,In_338,In_1836);
or U1625 (N_1625,In_991,In_1537);
nor U1626 (N_1626,In_1247,In_458);
nand U1627 (N_1627,In_489,In_397);
nand U1628 (N_1628,In_135,In_250);
and U1629 (N_1629,In_1565,In_1501);
and U1630 (N_1630,In_1406,In_1917);
nor U1631 (N_1631,In_845,In_119);
nor U1632 (N_1632,In_223,In_1147);
or U1633 (N_1633,In_1070,In_776);
nor U1634 (N_1634,In_1192,In_517);
nor U1635 (N_1635,In_626,In_489);
and U1636 (N_1636,In_226,In_1476);
and U1637 (N_1637,In_1992,In_1572);
or U1638 (N_1638,In_1367,In_1920);
or U1639 (N_1639,In_382,In_1904);
and U1640 (N_1640,In_1686,In_512);
and U1641 (N_1641,In_1357,In_975);
or U1642 (N_1642,In_1974,In_1841);
or U1643 (N_1643,In_558,In_696);
or U1644 (N_1644,In_1405,In_1637);
nor U1645 (N_1645,In_1304,In_1939);
nor U1646 (N_1646,In_429,In_763);
or U1647 (N_1647,In_342,In_876);
and U1648 (N_1648,In_82,In_1869);
nor U1649 (N_1649,In_699,In_882);
nand U1650 (N_1650,In_1248,In_1725);
xnor U1651 (N_1651,In_620,In_1824);
nand U1652 (N_1652,In_937,In_1637);
and U1653 (N_1653,In_1202,In_1918);
nor U1654 (N_1654,In_239,In_348);
nand U1655 (N_1655,In_445,In_1546);
or U1656 (N_1656,In_1462,In_468);
nand U1657 (N_1657,In_27,In_1621);
nor U1658 (N_1658,In_1301,In_543);
or U1659 (N_1659,In_239,In_642);
nand U1660 (N_1660,In_1331,In_1777);
nand U1661 (N_1661,In_768,In_995);
nand U1662 (N_1662,In_1970,In_354);
and U1663 (N_1663,In_1510,In_1168);
xor U1664 (N_1664,In_1331,In_1291);
nor U1665 (N_1665,In_183,In_88);
nand U1666 (N_1666,In_1664,In_1083);
nor U1667 (N_1667,In_349,In_1192);
or U1668 (N_1668,In_400,In_722);
and U1669 (N_1669,In_1615,In_1073);
nand U1670 (N_1670,In_803,In_581);
or U1671 (N_1671,In_1720,In_1198);
or U1672 (N_1672,In_1795,In_1744);
nand U1673 (N_1673,In_1008,In_1273);
or U1674 (N_1674,In_52,In_1979);
and U1675 (N_1675,In_257,In_932);
or U1676 (N_1676,In_1055,In_595);
or U1677 (N_1677,In_1458,In_607);
nor U1678 (N_1678,In_1625,In_1360);
nor U1679 (N_1679,In_1414,In_995);
and U1680 (N_1680,In_576,In_451);
and U1681 (N_1681,In_1188,In_1754);
nor U1682 (N_1682,In_1476,In_892);
nor U1683 (N_1683,In_727,In_1006);
or U1684 (N_1684,In_1034,In_1918);
or U1685 (N_1685,In_491,In_844);
nor U1686 (N_1686,In_1203,In_846);
xnor U1687 (N_1687,In_9,In_1633);
and U1688 (N_1688,In_712,In_1828);
or U1689 (N_1689,In_1471,In_108);
and U1690 (N_1690,In_1968,In_1162);
and U1691 (N_1691,In_1960,In_1585);
and U1692 (N_1692,In_337,In_1468);
nor U1693 (N_1693,In_1610,In_1299);
nor U1694 (N_1694,In_908,In_126);
nand U1695 (N_1695,In_1681,In_334);
xor U1696 (N_1696,In_630,In_499);
and U1697 (N_1697,In_1056,In_575);
and U1698 (N_1698,In_1486,In_1288);
nor U1699 (N_1699,In_100,In_1689);
or U1700 (N_1700,In_1972,In_1987);
and U1701 (N_1701,In_1160,In_1741);
nor U1702 (N_1702,In_1937,In_1821);
or U1703 (N_1703,In_1274,In_657);
and U1704 (N_1704,In_353,In_565);
and U1705 (N_1705,In_1646,In_1564);
nor U1706 (N_1706,In_1322,In_1130);
or U1707 (N_1707,In_842,In_1919);
and U1708 (N_1708,In_971,In_672);
and U1709 (N_1709,In_1409,In_812);
nand U1710 (N_1710,In_869,In_1009);
or U1711 (N_1711,In_1936,In_1834);
and U1712 (N_1712,In_1470,In_5);
nor U1713 (N_1713,In_841,In_450);
or U1714 (N_1714,In_61,In_1073);
nor U1715 (N_1715,In_1113,In_1716);
and U1716 (N_1716,In_443,In_1806);
nand U1717 (N_1717,In_516,In_58);
nand U1718 (N_1718,In_1352,In_1379);
nand U1719 (N_1719,In_692,In_1984);
nand U1720 (N_1720,In_1176,In_168);
and U1721 (N_1721,In_1342,In_1155);
xor U1722 (N_1722,In_790,In_1922);
or U1723 (N_1723,In_879,In_1553);
or U1724 (N_1724,In_1735,In_748);
xor U1725 (N_1725,In_1361,In_1108);
nor U1726 (N_1726,In_1924,In_1467);
or U1727 (N_1727,In_1019,In_688);
nand U1728 (N_1728,In_1574,In_773);
or U1729 (N_1729,In_1337,In_31);
nand U1730 (N_1730,In_310,In_8);
nor U1731 (N_1731,In_1261,In_1215);
nor U1732 (N_1732,In_1731,In_1453);
nand U1733 (N_1733,In_975,In_1633);
nor U1734 (N_1734,In_1500,In_1422);
nand U1735 (N_1735,In_156,In_1615);
and U1736 (N_1736,In_1650,In_775);
nor U1737 (N_1737,In_1456,In_1031);
xnor U1738 (N_1738,In_760,In_1791);
or U1739 (N_1739,In_505,In_1302);
and U1740 (N_1740,In_1284,In_364);
nor U1741 (N_1741,In_1211,In_1191);
and U1742 (N_1742,In_757,In_838);
and U1743 (N_1743,In_392,In_1097);
or U1744 (N_1744,In_1361,In_302);
nor U1745 (N_1745,In_1212,In_587);
and U1746 (N_1746,In_1153,In_110);
nor U1747 (N_1747,In_1180,In_1684);
or U1748 (N_1748,In_69,In_1575);
nand U1749 (N_1749,In_921,In_91);
and U1750 (N_1750,In_824,In_1510);
or U1751 (N_1751,In_1571,In_1721);
nand U1752 (N_1752,In_1216,In_1840);
and U1753 (N_1753,In_1095,In_703);
and U1754 (N_1754,In_1458,In_652);
and U1755 (N_1755,In_444,In_1916);
nand U1756 (N_1756,In_155,In_75);
nor U1757 (N_1757,In_1608,In_848);
nand U1758 (N_1758,In_292,In_740);
nand U1759 (N_1759,In_323,In_65);
and U1760 (N_1760,In_1520,In_384);
nand U1761 (N_1761,In_1118,In_1292);
nand U1762 (N_1762,In_310,In_658);
and U1763 (N_1763,In_355,In_1781);
nand U1764 (N_1764,In_1232,In_326);
or U1765 (N_1765,In_371,In_198);
and U1766 (N_1766,In_612,In_173);
xor U1767 (N_1767,In_1030,In_1047);
xor U1768 (N_1768,In_899,In_987);
and U1769 (N_1769,In_1073,In_1116);
nand U1770 (N_1770,In_1143,In_1251);
nand U1771 (N_1771,In_1264,In_254);
and U1772 (N_1772,In_61,In_444);
and U1773 (N_1773,In_1180,In_1425);
nor U1774 (N_1774,In_342,In_1295);
or U1775 (N_1775,In_1704,In_228);
or U1776 (N_1776,In_653,In_537);
nand U1777 (N_1777,In_868,In_65);
or U1778 (N_1778,In_483,In_1540);
nor U1779 (N_1779,In_864,In_1703);
nand U1780 (N_1780,In_1916,In_828);
xnor U1781 (N_1781,In_1825,In_403);
nand U1782 (N_1782,In_790,In_1032);
nor U1783 (N_1783,In_981,In_1580);
nor U1784 (N_1784,In_1453,In_1875);
nand U1785 (N_1785,In_1811,In_419);
and U1786 (N_1786,In_1838,In_344);
nand U1787 (N_1787,In_1024,In_1477);
and U1788 (N_1788,In_1711,In_1008);
nand U1789 (N_1789,In_1832,In_589);
or U1790 (N_1790,In_873,In_436);
or U1791 (N_1791,In_57,In_593);
nor U1792 (N_1792,In_812,In_56);
or U1793 (N_1793,In_1818,In_1522);
nor U1794 (N_1794,In_1402,In_741);
or U1795 (N_1795,In_1351,In_819);
xor U1796 (N_1796,In_297,In_1284);
and U1797 (N_1797,In_1028,In_705);
and U1798 (N_1798,In_1846,In_269);
xor U1799 (N_1799,In_159,In_1810);
or U1800 (N_1800,In_1556,In_1021);
nor U1801 (N_1801,In_819,In_779);
or U1802 (N_1802,In_1553,In_518);
and U1803 (N_1803,In_1030,In_1289);
nand U1804 (N_1804,In_1645,In_795);
and U1805 (N_1805,In_1820,In_1270);
nand U1806 (N_1806,In_514,In_1083);
or U1807 (N_1807,In_406,In_94);
or U1808 (N_1808,In_1194,In_1544);
and U1809 (N_1809,In_305,In_672);
or U1810 (N_1810,In_782,In_1306);
nand U1811 (N_1811,In_1983,In_614);
and U1812 (N_1812,In_442,In_1185);
nor U1813 (N_1813,In_1789,In_543);
xor U1814 (N_1814,In_1365,In_369);
xnor U1815 (N_1815,In_1440,In_488);
nand U1816 (N_1816,In_938,In_1449);
and U1817 (N_1817,In_164,In_993);
nand U1818 (N_1818,In_1853,In_1736);
nor U1819 (N_1819,In_477,In_700);
nor U1820 (N_1820,In_1957,In_1520);
nand U1821 (N_1821,In_1271,In_1582);
nand U1822 (N_1822,In_1073,In_1265);
nor U1823 (N_1823,In_1657,In_1909);
nor U1824 (N_1824,In_1777,In_778);
or U1825 (N_1825,In_1103,In_1596);
or U1826 (N_1826,In_56,In_938);
nand U1827 (N_1827,In_1198,In_1473);
and U1828 (N_1828,In_73,In_228);
or U1829 (N_1829,In_1492,In_1481);
or U1830 (N_1830,In_483,In_1293);
nor U1831 (N_1831,In_1682,In_1852);
nor U1832 (N_1832,In_52,In_336);
nor U1833 (N_1833,In_797,In_1353);
nor U1834 (N_1834,In_331,In_209);
nor U1835 (N_1835,In_1120,In_476);
nor U1836 (N_1836,In_1723,In_1786);
nand U1837 (N_1837,In_14,In_619);
nand U1838 (N_1838,In_197,In_1999);
and U1839 (N_1839,In_819,In_1291);
nand U1840 (N_1840,In_1414,In_1421);
xnor U1841 (N_1841,In_690,In_1517);
nand U1842 (N_1842,In_624,In_1761);
and U1843 (N_1843,In_633,In_1961);
or U1844 (N_1844,In_1852,In_1929);
nand U1845 (N_1845,In_1945,In_1450);
and U1846 (N_1846,In_1308,In_499);
nand U1847 (N_1847,In_1549,In_607);
nand U1848 (N_1848,In_1062,In_768);
nand U1849 (N_1849,In_1957,In_1112);
nand U1850 (N_1850,In_682,In_1890);
and U1851 (N_1851,In_434,In_1146);
nand U1852 (N_1852,In_1367,In_1430);
nor U1853 (N_1853,In_1444,In_1506);
and U1854 (N_1854,In_1379,In_984);
xnor U1855 (N_1855,In_1255,In_636);
xnor U1856 (N_1856,In_0,In_66);
nand U1857 (N_1857,In_1126,In_374);
nand U1858 (N_1858,In_743,In_252);
nand U1859 (N_1859,In_708,In_615);
or U1860 (N_1860,In_1216,In_1716);
nand U1861 (N_1861,In_1756,In_1595);
xnor U1862 (N_1862,In_1814,In_1866);
nor U1863 (N_1863,In_1844,In_1720);
or U1864 (N_1864,In_390,In_306);
nand U1865 (N_1865,In_69,In_1197);
and U1866 (N_1866,In_1640,In_601);
nor U1867 (N_1867,In_324,In_892);
nand U1868 (N_1868,In_149,In_897);
nor U1869 (N_1869,In_1306,In_1706);
or U1870 (N_1870,In_1735,In_259);
or U1871 (N_1871,In_840,In_826);
nand U1872 (N_1872,In_1125,In_1080);
and U1873 (N_1873,In_618,In_1858);
nor U1874 (N_1874,In_141,In_1869);
xnor U1875 (N_1875,In_442,In_1749);
xor U1876 (N_1876,In_1345,In_573);
and U1877 (N_1877,In_240,In_1196);
or U1878 (N_1878,In_1694,In_1687);
or U1879 (N_1879,In_969,In_1023);
nand U1880 (N_1880,In_613,In_1274);
nand U1881 (N_1881,In_18,In_723);
and U1882 (N_1882,In_1600,In_1830);
nor U1883 (N_1883,In_1619,In_81);
or U1884 (N_1884,In_1812,In_1286);
nand U1885 (N_1885,In_1778,In_1617);
nor U1886 (N_1886,In_362,In_1537);
nand U1887 (N_1887,In_1481,In_673);
nor U1888 (N_1888,In_1133,In_1588);
xnor U1889 (N_1889,In_1457,In_496);
nand U1890 (N_1890,In_496,In_419);
nor U1891 (N_1891,In_970,In_1307);
nand U1892 (N_1892,In_1040,In_633);
xnor U1893 (N_1893,In_1245,In_657);
nand U1894 (N_1894,In_1975,In_10);
or U1895 (N_1895,In_1195,In_1580);
nor U1896 (N_1896,In_919,In_1044);
nand U1897 (N_1897,In_1973,In_1970);
and U1898 (N_1898,In_63,In_261);
and U1899 (N_1899,In_111,In_566);
nor U1900 (N_1900,In_1855,In_1205);
nand U1901 (N_1901,In_891,In_1628);
nor U1902 (N_1902,In_103,In_878);
xor U1903 (N_1903,In_1634,In_71);
or U1904 (N_1904,In_1162,In_1000);
xnor U1905 (N_1905,In_1472,In_1560);
nor U1906 (N_1906,In_521,In_1726);
or U1907 (N_1907,In_1684,In_1886);
or U1908 (N_1908,In_586,In_1859);
nor U1909 (N_1909,In_993,In_1260);
and U1910 (N_1910,In_317,In_1834);
nor U1911 (N_1911,In_586,In_1660);
nand U1912 (N_1912,In_714,In_1218);
or U1913 (N_1913,In_544,In_603);
nor U1914 (N_1914,In_992,In_180);
xnor U1915 (N_1915,In_1225,In_384);
nand U1916 (N_1916,In_711,In_1816);
or U1917 (N_1917,In_453,In_855);
or U1918 (N_1918,In_151,In_1282);
and U1919 (N_1919,In_1716,In_1729);
and U1920 (N_1920,In_1008,In_132);
and U1921 (N_1921,In_502,In_1140);
and U1922 (N_1922,In_619,In_759);
nor U1923 (N_1923,In_1631,In_1733);
nand U1924 (N_1924,In_1126,In_350);
nand U1925 (N_1925,In_1906,In_1315);
nand U1926 (N_1926,In_114,In_1106);
nor U1927 (N_1927,In_1226,In_220);
nor U1928 (N_1928,In_801,In_1572);
and U1929 (N_1929,In_280,In_301);
nor U1930 (N_1930,In_1198,In_747);
and U1931 (N_1931,In_1109,In_1652);
xor U1932 (N_1932,In_1271,In_961);
nor U1933 (N_1933,In_1853,In_1047);
nor U1934 (N_1934,In_348,In_1522);
and U1935 (N_1935,In_325,In_1535);
nor U1936 (N_1936,In_444,In_1782);
nor U1937 (N_1937,In_1101,In_1879);
nor U1938 (N_1938,In_326,In_1708);
and U1939 (N_1939,In_515,In_968);
nand U1940 (N_1940,In_1004,In_291);
nor U1941 (N_1941,In_1915,In_1513);
xnor U1942 (N_1942,In_1815,In_895);
or U1943 (N_1943,In_490,In_1985);
nor U1944 (N_1944,In_1551,In_479);
nor U1945 (N_1945,In_23,In_1987);
nor U1946 (N_1946,In_1362,In_1223);
or U1947 (N_1947,In_1406,In_377);
and U1948 (N_1948,In_1611,In_828);
xor U1949 (N_1949,In_373,In_1183);
nand U1950 (N_1950,In_426,In_644);
or U1951 (N_1951,In_529,In_198);
nand U1952 (N_1952,In_276,In_1789);
and U1953 (N_1953,In_1733,In_1555);
and U1954 (N_1954,In_1887,In_1740);
or U1955 (N_1955,In_1664,In_559);
nand U1956 (N_1956,In_1570,In_1617);
nor U1957 (N_1957,In_540,In_788);
nand U1958 (N_1958,In_1923,In_1924);
nand U1959 (N_1959,In_986,In_1100);
and U1960 (N_1960,In_1849,In_707);
nor U1961 (N_1961,In_29,In_1926);
or U1962 (N_1962,In_252,In_897);
or U1963 (N_1963,In_1105,In_282);
and U1964 (N_1964,In_1048,In_1551);
or U1965 (N_1965,In_227,In_1133);
nor U1966 (N_1966,In_908,In_1553);
nor U1967 (N_1967,In_52,In_137);
xnor U1968 (N_1968,In_445,In_1940);
and U1969 (N_1969,In_1985,In_1146);
or U1970 (N_1970,In_1497,In_631);
nand U1971 (N_1971,In_978,In_409);
xor U1972 (N_1972,In_1052,In_1453);
nor U1973 (N_1973,In_360,In_911);
or U1974 (N_1974,In_690,In_241);
nand U1975 (N_1975,In_232,In_263);
xnor U1976 (N_1976,In_1093,In_570);
nand U1977 (N_1977,In_1710,In_855);
nand U1978 (N_1978,In_1031,In_862);
or U1979 (N_1979,In_1175,In_1089);
xor U1980 (N_1980,In_1313,In_687);
and U1981 (N_1981,In_1494,In_871);
and U1982 (N_1982,In_314,In_1010);
xor U1983 (N_1983,In_856,In_340);
nor U1984 (N_1984,In_1250,In_905);
and U1985 (N_1985,In_1131,In_1629);
and U1986 (N_1986,In_979,In_740);
or U1987 (N_1987,In_360,In_219);
xnor U1988 (N_1988,In_132,In_1270);
xor U1989 (N_1989,In_1461,In_1133);
nor U1990 (N_1990,In_135,In_162);
nand U1991 (N_1991,In_1233,In_1950);
or U1992 (N_1992,In_1957,In_747);
and U1993 (N_1993,In_1118,In_899);
and U1994 (N_1994,In_662,In_1994);
nand U1995 (N_1995,In_1530,In_1488);
and U1996 (N_1996,In_1234,In_1564);
and U1997 (N_1997,In_448,In_812);
nand U1998 (N_1998,In_493,In_339);
xnor U1999 (N_1999,In_585,In_1924);
and U2000 (N_2000,N_1023,N_900);
or U2001 (N_2001,N_1809,N_865);
nand U2002 (N_2002,N_1434,N_35);
nand U2003 (N_2003,N_1416,N_97);
nand U2004 (N_2004,N_369,N_1149);
and U2005 (N_2005,N_1052,N_1264);
and U2006 (N_2006,N_281,N_661);
nand U2007 (N_2007,N_786,N_464);
nand U2008 (N_2008,N_156,N_1516);
or U2009 (N_2009,N_303,N_546);
nand U2010 (N_2010,N_1639,N_1127);
or U2011 (N_2011,N_1688,N_1100);
nor U2012 (N_2012,N_1588,N_750);
and U2013 (N_2013,N_1738,N_270);
nand U2014 (N_2014,N_1184,N_532);
or U2015 (N_2015,N_267,N_1774);
nor U2016 (N_2016,N_1800,N_1016);
xnor U2017 (N_2017,N_1144,N_1124);
and U2018 (N_2018,N_1551,N_645);
and U2019 (N_2019,N_187,N_98);
and U2020 (N_2020,N_757,N_1054);
and U2021 (N_2021,N_1439,N_1563);
and U2022 (N_2022,N_1213,N_1285);
and U2023 (N_2023,N_1346,N_400);
and U2024 (N_2024,N_344,N_130);
nor U2025 (N_2025,N_899,N_590);
xor U2026 (N_2026,N_869,N_765);
nor U2027 (N_2027,N_1869,N_1519);
nand U2028 (N_2028,N_1719,N_808);
and U2029 (N_2029,N_1091,N_1922);
and U2030 (N_2030,N_1497,N_1482);
and U2031 (N_2031,N_66,N_1546);
nor U2032 (N_2032,N_990,N_725);
nand U2033 (N_2033,N_30,N_1320);
or U2034 (N_2034,N_818,N_712);
nor U2035 (N_2035,N_1938,N_381);
and U2036 (N_2036,N_289,N_1543);
or U2037 (N_2037,N_1520,N_1002);
nand U2038 (N_2038,N_135,N_1778);
or U2039 (N_2039,N_128,N_1772);
or U2040 (N_2040,N_150,N_1697);
nand U2041 (N_2041,N_326,N_1804);
xor U2042 (N_2042,N_413,N_345);
nor U2043 (N_2043,N_184,N_1846);
nor U2044 (N_2044,N_1401,N_160);
nor U2045 (N_2045,N_901,N_257);
and U2046 (N_2046,N_279,N_134);
or U2047 (N_2047,N_678,N_81);
nor U2048 (N_2048,N_908,N_1703);
and U2049 (N_2049,N_877,N_685);
nor U2050 (N_2050,N_236,N_1567);
or U2051 (N_2051,N_827,N_767);
nand U2052 (N_2052,N_789,N_352);
nand U2053 (N_2053,N_1132,N_1750);
or U2054 (N_2054,N_1968,N_719);
xnor U2055 (N_2055,N_537,N_198);
and U2056 (N_2056,N_1629,N_1930);
and U2057 (N_2057,N_1428,N_738);
nor U2058 (N_2058,N_742,N_577);
nor U2059 (N_2059,N_953,N_1090);
or U2060 (N_2060,N_860,N_633);
nand U2061 (N_2061,N_103,N_237);
or U2062 (N_2062,N_36,N_1097);
or U2063 (N_2063,N_245,N_1308);
nor U2064 (N_2064,N_701,N_843);
nand U2065 (N_2065,N_1397,N_788);
nor U2066 (N_2066,N_74,N_620);
nor U2067 (N_2067,N_598,N_6);
or U2068 (N_2068,N_567,N_784);
or U2069 (N_2069,N_1518,N_318);
and U2070 (N_2070,N_583,N_215);
xnor U2071 (N_2071,N_1284,N_1559);
nand U2072 (N_2072,N_1610,N_675);
or U2073 (N_2073,N_434,N_1895);
and U2074 (N_2074,N_365,N_1408);
or U2075 (N_2075,N_111,N_1775);
or U2076 (N_2076,N_1523,N_906);
xor U2077 (N_2077,N_1553,N_1229);
xor U2078 (N_2078,N_1542,N_86);
and U2079 (N_2079,N_1392,N_1530);
xnor U2080 (N_2080,N_528,N_129);
nor U2081 (N_2081,N_116,N_1910);
nand U2082 (N_2082,N_1390,N_399);
or U2083 (N_2083,N_649,N_1965);
or U2084 (N_2084,N_1709,N_353);
or U2085 (N_2085,N_1012,N_161);
nor U2086 (N_2086,N_787,N_1374);
and U2087 (N_2087,N_1803,N_1407);
nor U2088 (N_2088,N_1472,N_96);
nor U2089 (N_2089,N_1698,N_561);
nand U2090 (N_2090,N_166,N_447);
nand U2091 (N_2091,N_1872,N_1584);
xor U2092 (N_2092,N_1524,N_1795);
nand U2093 (N_2093,N_1594,N_846);
xnor U2094 (N_2094,N_1433,N_1333);
or U2095 (N_2095,N_1598,N_163);
nor U2096 (N_2096,N_201,N_987);
xor U2097 (N_2097,N_1662,N_1010);
nor U2098 (N_2098,N_1780,N_1391);
nor U2099 (N_2099,N_254,N_662);
and U2100 (N_2100,N_1783,N_1625);
nand U2101 (N_2101,N_1048,N_1825);
nor U2102 (N_2102,N_1493,N_1249);
xnor U2103 (N_2103,N_991,N_211);
nand U2104 (N_2104,N_898,N_230);
xor U2105 (N_2105,N_722,N_558);
nor U2106 (N_2106,N_466,N_624);
nor U2107 (N_2107,N_1668,N_1621);
and U2108 (N_2108,N_132,N_515);
xor U2109 (N_2109,N_829,N_456);
nand U2110 (N_2110,N_1821,N_1175);
and U2111 (N_2111,N_210,N_1962);
nor U2112 (N_2112,N_1202,N_33);
and U2113 (N_2113,N_1381,N_1105);
or U2114 (N_2114,N_1086,N_1852);
nor U2115 (N_2115,N_259,N_1989);
nand U2116 (N_2116,N_133,N_605);
nor U2117 (N_2117,N_179,N_938);
nand U2118 (N_2118,N_1166,N_1145);
and U2119 (N_2119,N_1254,N_1395);
nor U2120 (N_2120,N_1337,N_266);
or U2121 (N_2121,N_555,N_1443);
nand U2122 (N_2122,N_856,N_142);
xor U2123 (N_2123,N_1875,N_285);
xor U2124 (N_2124,N_917,N_582);
nor U2125 (N_2125,N_239,N_1713);
xor U2126 (N_2126,N_394,N_739);
and U2127 (N_2127,N_518,N_28);
nor U2128 (N_2128,N_1951,N_1237);
or U2129 (N_2129,N_554,N_1599);
and U2130 (N_2130,N_1736,N_1440);
or U2131 (N_2131,N_798,N_999);
nor U2132 (N_2132,N_51,N_146);
nand U2133 (N_2133,N_1212,N_770);
or U2134 (N_2134,N_1690,N_1691);
and U2135 (N_2135,N_1609,N_440);
and U2136 (N_2136,N_1334,N_57);
nor U2137 (N_2137,N_1777,N_492);
and U2138 (N_2138,N_1011,N_1661);
or U2139 (N_2139,N_942,N_88);
and U2140 (N_2140,N_1506,N_71);
or U2141 (N_2141,N_1812,N_1914);
nor U2142 (N_2142,N_1197,N_1365);
and U2143 (N_2143,N_273,N_1295);
nand U2144 (N_2144,N_931,N_397);
and U2145 (N_2145,N_506,N_1238);
or U2146 (N_2146,N_795,N_1566);
or U2147 (N_2147,N_659,N_1163);
nand U2148 (N_2148,N_1928,N_1529);
and U2149 (N_2149,N_1708,N_1502);
nor U2150 (N_2150,N_148,N_252);
or U2151 (N_2151,N_1014,N_589);
and U2152 (N_2152,N_1402,N_1160);
nand U2153 (N_2153,N_1767,N_1223);
or U2154 (N_2154,N_1796,N_1741);
and U2155 (N_2155,N_1555,N_436);
or U2156 (N_2156,N_1918,N_1554);
or U2157 (N_2157,N_1611,N_1865);
nand U2158 (N_2158,N_206,N_1317);
nand U2159 (N_2159,N_337,N_534);
and U2160 (N_2160,N_115,N_1169);
nor U2161 (N_2161,N_277,N_423);
nand U2162 (N_2162,N_668,N_370);
nand U2163 (N_2163,N_1283,N_797);
xor U2164 (N_2164,N_1387,N_1373);
or U2165 (N_2165,N_92,N_1185);
and U2166 (N_2166,N_1060,N_102);
nor U2167 (N_2167,N_993,N_527);
nor U2168 (N_2168,N_34,N_861);
or U2169 (N_2169,N_1527,N_62);
or U2170 (N_2170,N_175,N_1031);
and U2171 (N_2171,N_327,N_806);
and U2172 (N_2172,N_233,N_510);
nand U2173 (N_2173,N_626,N_976);
nor U2174 (N_2174,N_1255,N_1253);
or U2175 (N_2175,N_1168,N_835);
and U2176 (N_2176,N_1075,N_979);
nor U2177 (N_2177,N_138,N_501);
xor U2178 (N_2178,N_1890,N_793);
nor U2179 (N_2179,N_1481,N_1470);
and U2180 (N_2180,N_1029,N_1987);
nand U2181 (N_2181,N_1752,N_1514);
or U2182 (N_2182,N_1819,N_731);
and U2183 (N_2183,N_38,N_1004);
nand U2184 (N_2184,N_1332,N_1612);
and U2185 (N_2185,N_1233,N_1537);
and U2186 (N_2186,N_780,N_648);
xor U2187 (N_2187,N_242,N_1787);
nand U2188 (N_2188,N_1125,N_1595);
or U2189 (N_2189,N_1517,N_875);
nand U2190 (N_2190,N_1855,N_190);
xnor U2191 (N_2191,N_570,N_1905);
or U2192 (N_2192,N_1486,N_830);
and U2193 (N_2193,N_680,N_1837);
and U2194 (N_2194,N_55,N_517);
nor U2195 (N_2195,N_1119,N_1972);
nand U2196 (N_2196,N_568,N_499);
nand U2197 (N_2197,N_614,N_1991);
nand U2198 (N_2198,N_1062,N_1321);
xor U2199 (N_2199,N_1158,N_1758);
or U2200 (N_2200,N_1248,N_1154);
and U2201 (N_2201,N_1976,N_841);
or U2202 (N_2202,N_1560,N_287);
nor U2203 (N_2203,N_1384,N_1526);
nand U2204 (N_2204,N_87,N_304);
and U2205 (N_2205,N_1769,N_984);
or U2206 (N_2206,N_692,N_1005);
nand U2207 (N_2207,N_696,N_982);
and U2208 (N_2208,N_1178,N_1096);
nand U2209 (N_2209,N_1376,N_973);
or U2210 (N_2210,N_151,N_530);
nand U2211 (N_2211,N_1570,N_1994);
and U2212 (N_2212,N_264,N_941);
and U2213 (N_2213,N_791,N_320);
nor U2214 (N_2214,N_361,N_1114);
and U2215 (N_2215,N_1579,N_2);
or U2216 (N_2216,N_1483,N_154);
nor U2217 (N_2217,N_1521,N_507);
or U2218 (N_2218,N_1207,N_358);
nor U2219 (N_2219,N_1288,N_1901);
nand U2220 (N_2220,N_606,N_1307);
and U2221 (N_2221,N_1650,N_241);
and U2222 (N_2222,N_1165,N_26);
nand U2223 (N_2223,N_7,N_1418);
nor U2224 (N_2224,N_1235,N_1722);
nor U2225 (N_2225,N_1663,N_595);
or U2226 (N_2226,N_222,N_1360);
nand U2227 (N_2227,N_978,N_1270);
or U2228 (N_2228,N_193,N_774);
or U2229 (N_2229,N_1082,N_885);
nand U2230 (N_2230,N_1632,N_936);
or U2231 (N_2231,N_1366,N_228);
nor U2232 (N_2232,N_69,N_123);
nor U2233 (N_2233,N_964,N_1919);
nand U2234 (N_2234,N_1068,N_1730);
and U2235 (N_2235,N_862,N_800);
nor U2236 (N_2236,N_359,N_1456);
nand U2237 (N_2237,N_278,N_1265);
nand U2238 (N_2238,N_110,N_1351);
and U2239 (N_2239,N_801,N_1071);
xor U2240 (N_2240,N_455,N_101);
nor U2241 (N_2241,N_1676,N_1773);
nand U2242 (N_2242,N_1940,N_505);
nor U2243 (N_2243,N_173,N_700);
and U2244 (N_2244,N_905,N_1490);
nand U2245 (N_2245,N_1534,N_1686);
nand U2246 (N_2246,N_73,N_349);
and U2247 (N_2247,N_1049,N_1934);
nor U2248 (N_2248,N_391,N_27);
nor U2249 (N_2249,N_1271,N_824);
and U2250 (N_2250,N_693,N_1535);
and U2251 (N_2251,N_366,N_751);
or U2252 (N_2252,N_1904,N_691);
or U2253 (N_2253,N_1451,N_486);
or U2254 (N_2254,N_164,N_954);
nor U2255 (N_2255,N_1246,N_1492);
or U2256 (N_2256,N_377,N_1389);
xor U2257 (N_2257,N_1619,N_269);
and U2258 (N_2258,N_83,N_522);
or U2259 (N_2259,N_1247,N_1834);
or U2260 (N_2260,N_430,N_1179);
or U2261 (N_2261,N_802,N_374);
nor U2262 (N_2262,N_169,N_821);
xor U2263 (N_2263,N_1377,N_1172);
nand U2264 (N_2264,N_826,N_1720);
nand U2265 (N_2265,N_78,N_911);
and U2266 (N_2266,N_481,N_1866);
xor U2267 (N_2267,N_435,N_588);
nand U2268 (N_2268,N_1108,N_1427);
xor U2269 (N_2269,N_415,N_104);
nand U2270 (N_2270,N_1471,N_468);
nor U2271 (N_2271,N_1889,N_574);
nor U2272 (N_2272,N_1358,N_1932);
nand U2273 (N_2273,N_416,N_1412);
nand U2274 (N_2274,N_232,N_526);
and U2275 (N_2275,N_1980,N_213);
and U2276 (N_2276,N_769,N_1467);
or U2277 (N_2277,N_1893,N_820);
nand U2278 (N_2278,N_748,N_1653);
and U2279 (N_2279,N_596,N_642);
nor U2280 (N_2280,N_1117,N_1139);
xor U2281 (N_2281,N_43,N_579);
and U2282 (N_2282,N_1743,N_876);
or U2283 (N_2283,N_533,N_811);
nor U2284 (N_2284,N_168,N_32);
nor U2285 (N_2285,N_1615,N_282);
nor U2286 (N_2286,N_1626,N_1022);
or U2287 (N_2287,N_321,N_1279);
or U2288 (N_2288,N_1756,N_839);
nor U2289 (N_2289,N_1177,N_195);
nand U2290 (N_2290,N_749,N_1324);
and U2291 (N_2291,N_998,N_641);
and U2292 (N_2292,N_708,N_197);
or U2293 (N_2293,N_1099,N_362);
nand U2294 (N_2294,N_593,N_1239);
xnor U2295 (N_2295,N_1019,N_286);
nor U2296 (N_2296,N_1256,N_1654);
nand U2297 (N_2297,N_909,N_790);
nand U2298 (N_2298,N_1251,N_1590);
nor U2299 (N_2299,N_39,N_1208);
and U2300 (N_2300,N_1357,N_1845);
and U2301 (N_2301,N_1072,N_1779);
nand U2302 (N_2302,N_258,N_170);
or U2303 (N_2303,N_1380,N_1695);
or U2304 (N_2304,N_341,N_90);
nand U2305 (N_2305,N_472,N_873);
or U2306 (N_2306,N_1876,N_1643);
or U2307 (N_2307,N_776,N_1963);
nor U2308 (N_2308,N_1969,N_1533);
nand U2309 (N_2309,N_1445,N_716);
and U2310 (N_2310,N_1372,N_666);
or U2311 (N_2311,N_1996,N_1182);
nor U2312 (N_2312,N_837,N_1435);
or U2313 (N_2313,N_144,N_200);
and U2314 (N_2314,N_1282,N_1310);
and U2315 (N_2315,N_1788,N_1926);
or U2316 (N_2316,N_189,N_1180);
xnor U2317 (N_2317,N_22,N_1808);
nand U2318 (N_2318,N_833,N_45);
nand U2319 (N_2319,N_1051,N_1102);
and U2320 (N_2320,N_405,N_350);
nor U2321 (N_2321,N_562,N_1327);
or U2322 (N_2322,N_732,N_323);
or U2323 (N_2323,N_652,N_336);
nor U2324 (N_2324,N_325,N_294);
nand U2325 (N_2325,N_1089,N_771);
nand U2326 (N_2326,N_1419,N_172);
nand U2327 (N_2327,N_409,N_403);
nand U2328 (N_2328,N_699,N_1340);
nor U2329 (N_2329,N_575,N_1155);
nor U2330 (N_2330,N_916,N_1015);
or U2331 (N_2331,N_1272,N_225);
xor U2332 (N_2332,N_1647,N_1129);
or U2333 (N_2333,N_1781,N_1651);
nand U2334 (N_2334,N_1126,N_223);
nand U2335 (N_2335,N_1268,N_1147);
or U2336 (N_2336,N_915,N_311);
nor U2337 (N_2337,N_1457,N_1494);
and U2338 (N_2338,N_773,N_1913);
and U2339 (N_2339,N_1188,N_1701);
and U2340 (N_2340,N_346,N_1681);
or U2341 (N_2341,N_1092,N_77);
and U2342 (N_2342,N_1735,N_1261);
nand U2343 (N_2343,N_1525,N_244);
and U2344 (N_2344,N_1061,N_997);
nand U2345 (N_2345,N_1881,N_1740);
or U2346 (N_2346,N_470,N_108);
and U2347 (N_2347,N_737,N_1322);
nor U2348 (N_2348,N_857,N_1449);
and U2349 (N_2349,N_1911,N_376);
and U2350 (N_2350,N_1400,N_141);
nand U2351 (N_2351,N_24,N_1198);
or U2352 (N_2352,N_1136,N_11);
or U2353 (N_2353,N_935,N_1243);
or U2354 (N_2354,N_18,N_729);
or U2355 (N_2355,N_753,N_946);
or U2356 (N_2356,N_1488,N_432);
nand U2357 (N_2357,N_717,N_1694);
xnor U2358 (N_2358,N_112,N_1053);
xnor U2359 (N_2359,N_1763,N_319);
xnor U2360 (N_2360,N_247,N_1966);
or U2361 (N_2361,N_1263,N_1915);
or U2362 (N_2362,N_1081,N_989);
xnor U2363 (N_2363,N_721,N_1747);
nand U2364 (N_2364,N_1103,N_1847);
nor U2365 (N_2365,N_1411,N_450);
and U2366 (N_2366,N_385,N_1896);
or U2367 (N_2367,N_1868,N_995);
or U2368 (N_2368,N_969,N_1296);
nand U2369 (N_2369,N_186,N_1157);
or U2370 (N_2370,N_1798,N_1880);
nor U2371 (N_2371,N_819,N_832);
nand U2372 (N_2372,N_1133,N_778);
xnor U2373 (N_2373,N_1485,N_126);
nand U2374 (N_2374,N_99,N_1792);
nand U2375 (N_2375,N_1162,N_0);
or U2376 (N_2376,N_1274,N_958);
or U2377 (N_2377,N_392,N_1156);
nand U2378 (N_2378,N_1689,N_157);
nor U2379 (N_2379,N_1806,N_1835);
nand U2380 (N_2380,N_713,N_1454);
or U2381 (N_2381,N_752,N_1326);
or U2382 (N_2382,N_1547,N_1899);
nand U2383 (N_2383,N_672,N_566);
nor U2384 (N_2384,N_634,N_585);
or U2385 (N_2385,N_1027,N_1167);
nand U2386 (N_2386,N_1776,N_1093);
nand U2387 (N_2387,N_1173,N_1718);
xnor U2388 (N_2388,N_76,N_478);
or U2389 (N_2389,N_1228,N_1441);
or U2390 (N_2390,N_1964,N_919);
nand U2391 (N_2391,N_1013,N_602);
nor U2392 (N_2392,N_17,N_1649);
xnor U2393 (N_2393,N_924,N_1205);
xor U2394 (N_2394,N_474,N_1058);
and U2395 (N_2395,N_107,N_1503);
xor U2396 (N_2396,N_364,N_697);
xor U2397 (N_2397,N_262,N_1903);
nand U2398 (N_2398,N_1830,N_469);
xor U2399 (N_2399,N_887,N_1276);
xor U2400 (N_2400,N_1059,N_647);
and U2401 (N_2401,N_4,N_1020);
and U2402 (N_2402,N_961,N_1887);
xnor U2403 (N_2403,N_1844,N_1764);
or U2404 (N_2404,N_1946,N_1413);
or U2405 (N_2405,N_1396,N_1544);
nor U2406 (N_2406,N_601,N_667);
nor U2407 (N_2407,N_1040,N_1083);
nand U2408 (N_2408,N_411,N_1363);
or U2409 (N_2409,N_484,N_1323);
nor U2410 (N_2410,N_1608,N_1035);
or U2411 (N_2411,N_1312,N_192);
nand U2412 (N_2412,N_204,N_1328);
and U2413 (N_2413,N_50,N_893);
nand U2414 (N_2414,N_971,N_1917);
nand U2415 (N_2415,N_914,N_730);
nor U2416 (N_2416,N_373,N_1286);
or U2417 (N_2417,N_834,N_1631);
or U2418 (N_2418,N_454,N_1665);
nand U2419 (N_2419,N_1696,N_1080);
and U2420 (N_2420,N_1039,N_1531);
xor U2421 (N_2421,N_448,N_1827);
nor U2422 (N_2422,N_497,N_1267);
xnor U2423 (N_2423,N_1771,N_445);
or U2424 (N_2424,N_1123,N_1448);
and U2425 (N_2425,N_1085,N_1836);
nand U2426 (N_2426,N_1583,N_1414);
nor U2427 (N_2427,N_580,N_1260);
and U2428 (N_2428,N_420,N_21);
nand U2429 (N_2429,N_695,N_139);
nor U2430 (N_2430,N_334,N_525);
and U2431 (N_2431,N_308,N_382);
or U2432 (N_2432,N_607,N_1672);
xor U2433 (N_2433,N_967,N_889);
nand U2434 (N_2434,N_1843,N_1464);
and U2435 (N_2435,N_523,N_882);
and U2436 (N_2436,N_1603,N_429);
or U2437 (N_2437,N_932,N_433);
and U2438 (N_2438,N_1909,N_202);
and U2439 (N_2439,N_714,N_1799);
and U2440 (N_2440,N_1591,N_145);
nor U2441 (N_2441,N_60,N_458);
nor U2442 (N_2442,N_581,N_1225);
xnor U2443 (N_2443,N_490,N_1680);
and U2444 (N_2444,N_733,N_1556);
nand U2445 (N_2445,N_944,N_89);
or U2446 (N_2446,N_947,N_1159);
nor U2447 (N_2447,N_631,N_855);
nand U2448 (N_2448,N_1148,N_1298);
nor U2449 (N_2449,N_943,N_387);
and U2450 (N_2450,N_950,N_105);
and U2451 (N_2451,N_970,N_1863);
nand U2452 (N_2452,N_754,N_1578);
xor U2453 (N_2453,N_1110,N_1122);
nand U2454 (N_2454,N_1728,N_255);
or U2455 (N_2455,N_1245,N_1368);
nor U2456 (N_2456,N_660,N_1107);
nand U2457 (N_2457,N_1459,N_246);
and U2458 (N_2458,N_386,N_1305);
nand U2459 (N_2459,N_1006,N_1532);
xnor U2460 (N_2460,N_1755,N_3);
nand U2461 (N_2461,N_292,N_1386);
nand U2462 (N_2462,N_628,N_892);
nand U2463 (N_2463,N_1854,N_512);
nand U2464 (N_2464,N_1942,N_1884);
or U2465 (N_2465,N_70,N_854);
or U2466 (N_2466,N_1988,N_923);
nor U2467 (N_2467,N_53,N_137);
and U2468 (N_2468,N_952,N_59);
nand U2469 (N_2469,N_298,N_351);
and U2470 (N_2470,N_147,N_272);
nor U2471 (N_2471,N_155,N_84);
and U2472 (N_2472,N_1498,N_1751);
and U2473 (N_2473,N_1982,N_331);
nand U2474 (N_2474,N_1871,N_1912);
or U2475 (N_2475,N_1765,N_1768);
and U2476 (N_2476,N_182,N_1431);
nor U2477 (N_2477,N_1897,N_1929);
and U2478 (N_2478,N_1187,N_487);
nand U2479 (N_2479,N_1316,N_1714);
and U2480 (N_2480,N_1294,N_457);
nor U2481 (N_2481,N_868,N_1141);
and U2482 (N_2482,N_449,N_1641);
and U2483 (N_2483,N_1923,N_1955);
nor U2484 (N_2484,N_564,N_1944);
nand U2485 (N_2485,N_1415,N_1558);
nor U2486 (N_2486,N_300,N_880);
and U2487 (N_2487,N_1329,N_1000);
and U2488 (N_2488,N_1601,N_438);
nor U2489 (N_2489,N_888,N_578);
nand U2490 (N_2490,N_746,N_1309);
and U2491 (N_2491,N_207,N_1648);
xor U2492 (N_2492,N_1269,N_1444);
nor U2493 (N_2493,N_723,N_473);
or U2494 (N_2494,N_1215,N_1879);
and U2495 (N_2495,N_951,N_879);
nor U2496 (N_2496,N_992,N_1146);
nor U2497 (N_2497,N_619,N_1447);
and U2498 (N_2498,N_1084,N_597);
or U2499 (N_2499,N_167,N_1504);
or U2500 (N_2500,N_1784,N_912);
or U2501 (N_2501,N_1352,N_1183);
nor U2502 (N_2502,N_1813,N_493);
nand U2503 (N_2503,N_792,N_406);
xor U2504 (N_2504,N_329,N_1815);
or U2505 (N_2505,N_1860,N_1353);
and U2506 (N_2506,N_963,N_1927);
or U2507 (N_2507,N_710,N_965);
nand U2508 (N_2508,N_238,N_1682);
and U2509 (N_2509,N_1618,N_1637);
or U2510 (N_2510,N_328,N_1937);
and U2511 (N_2511,N_1950,N_1839);
or U2512 (N_2512,N_1424,N_1109);
nand U2513 (N_2513,N_1707,N_371);
and U2514 (N_2514,N_758,N_674);
and U2515 (N_2515,N_867,N_521);
or U2516 (N_2516,N_480,N_871);
nand U2517 (N_2517,N_58,N_996);
nor U2518 (N_2518,N_1958,N_844);
nor U2519 (N_2519,N_1112,N_1685);
or U2520 (N_2520,N_380,N_479);
or U2521 (N_2521,N_1473,N_1677);
and U2522 (N_2522,N_1453,N_1607);
nand U2523 (N_2523,N_1138,N_772);
nor U2524 (N_2524,N_1231,N_1505);
or U2525 (N_2525,N_460,N_980);
nand U2526 (N_2526,N_1992,N_840);
xnor U2527 (N_2527,N_23,N_1240);
or U2528 (N_2528,N_1509,N_886);
nor U2529 (N_2529,N_1345,N_1571);
nand U2530 (N_2530,N_442,N_1151);
or U2531 (N_2531,N_1883,N_524);
or U2532 (N_2532,N_630,N_859);
nor U2533 (N_2533,N_265,N_599);
and U2534 (N_2534,N_894,N_342);
nor U2535 (N_2535,N_1581,N_632);
nor U2536 (N_2536,N_918,N_1920);
or U2537 (N_2537,N_1699,N_1826);
nor U2538 (N_2538,N_1857,N_939);
nor U2539 (N_2539,N_520,N_1200);
or U2540 (N_2540,N_1737,N_1540);
nor U2541 (N_2541,N_745,N_1287);
and U2542 (N_2542,N_1194,N_1477);
or U2543 (N_2543,N_1131,N_673);
and U2544 (N_2544,N_1580,N_476);
nor U2545 (N_2545,N_1902,N_1297);
or U2546 (N_2546,N_592,N_1028);
or U2547 (N_2547,N_1393,N_694);
nor U2548 (N_2548,N_288,N_1042);
nand U2549 (N_2549,N_1828,N_610);
nand U2550 (N_2550,N_1266,N_1350);
or U2551 (N_2551,N_500,N_679);
nand U2552 (N_2552,N_261,N_726);
nand U2553 (N_2553,N_890,N_419);
nor U2554 (N_2554,N_925,N_1704);
and U2555 (N_2555,N_848,N_1971);
or U2556 (N_2556,N_12,N_307);
nand U2557 (N_2557,N_1589,N_418);
nor U2558 (N_2558,N_937,N_689);
or U2559 (N_2559,N_1931,N_1805);
nand U2560 (N_2560,N_19,N_1410);
nand U2561 (N_2561,N_1638,N_1802);
nor U2562 (N_2562,N_1954,N_706);
or U2563 (N_2563,N_594,N_437);
nand U2564 (N_2564,N_1257,N_755);
nand U2565 (N_2565,N_571,N_1731);
nor U2566 (N_2566,N_1303,N_176);
nor U2567 (N_2567,N_1717,N_682);
and U2568 (N_2568,N_1655,N_569);
nor U2569 (N_2569,N_849,N_1164);
nand U2570 (N_2570,N_1450,N_547);
and U2571 (N_2571,N_687,N_807);
or U2572 (N_2572,N_275,N_1193);
and U2573 (N_2573,N_1293,N_1760);
xnor U2574 (N_2574,N_744,N_1087);
nor U2575 (N_2575,N_274,N_10);
and U2576 (N_2576,N_1500,N_1189);
or U2577 (N_2577,N_1790,N_203);
and U2578 (N_2578,N_249,N_1104);
xnor U2579 (N_2579,N_1113,N_15);
nor U2580 (N_2580,N_1073,N_813);
xor U2581 (N_2581,N_426,N_1403);
or U2582 (N_2582,N_251,N_759);
and U2583 (N_2583,N_462,N_1820);
and U2584 (N_2584,N_657,N_1398);
or U2585 (N_2585,N_529,N_1512);
and U2586 (N_2586,N_1220,N_1593);
or U2587 (N_2587,N_872,N_1423);
and U2588 (N_2588,N_777,N_794);
nand U2589 (N_2589,N_482,N_1782);
xnor U2590 (N_2590,N_1945,N_1949);
xnor U2591 (N_2591,N_1037,N_650);
nor U2592 (N_2592,N_1227,N_178);
nand U2593 (N_2593,N_1056,N_221);
xnor U2594 (N_2594,N_1562,N_1636);
or U2595 (N_2595,N_1628,N_1121);
or U2596 (N_2596,N_1216,N_1959);
nand U2597 (N_2597,N_1007,N_496);
and U2598 (N_2598,N_283,N_56);
nor U2599 (N_2599,N_1900,N_1838);
or U2600 (N_2600,N_1577,N_519);
xor U2601 (N_2601,N_904,N_783);
nand U2602 (N_2602,N_1361,N_1936);
and U2603 (N_2603,N_535,N_629);
or U2604 (N_2604,N_1409,N_1644);
nor U2605 (N_2605,N_930,N_1549);
or U2606 (N_2606,N_1452,N_1226);
nor U2607 (N_2607,N_1916,N_1851);
nand U2608 (N_2608,N_1032,N_735);
xnor U2609 (N_2609,N_149,N_1711);
and U2610 (N_2610,N_1613,N_1375);
nand U2611 (N_2611,N_119,N_962);
nand U2612 (N_2612,N_705,N_1742);
nand U2613 (N_2613,N_1793,N_1422);
nor U2614 (N_2614,N_355,N_831);
and U2615 (N_2615,N_842,N_29);
and U2616 (N_2616,N_1399,N_728);
nor U2617 (N_2617,N_1687,N_981);
nand U2618 (N_2618,N_960,N_100);
or U2619 (N_2619,N_1956,N_1822);
and U2620 (N_2620,N_1548,N_1630);
or U2621 (N_2621,N_1705,N_616);
nor U2622 (N_2622,N_118,N_1234);
xnor U2623 (N_2623,N_637,N_1436);
and U2624 (N_2624,N_983,N_1379);
nand U2625 (N_2625,N_1466,N_404);
xnor U2626 (N_2626,N_63,N_698);
xnor U2627 (N_2627,N_498,N_782);
or U2628 (N_2628,N_1744,N_1442);
nand U2629 (N_2629,N_1,N_1842);
nand U2630 (N_2630,N_550,N_240);
and U2631 (N_2631,N_216,N_422);
or U2632 (N_2632,N_1475,N_1678);
xnor U2633 (N_2633,N_219,N_870);
and U2634 (N_2634,N_1315,N_1635);
nor U2635 (N_2635,N_1501,N_1191);
nor U2636 (N_2636,N_718,N_1468);
nand U2637 (N_2637,N_1095,N_1766);
xnor U2638 (N_2638,N_20,N_1242);
and U2639 (N_2639,N_1078,N_741);
nor U2640 (N_2640,N_177,N_1118);
and U2641 (N_2641,N_1356,N_1645);
and U2642 (N_2642,N_1437,N_878);
nor U2643 (N_2643,N_1885,N_425);
or U2644 (N_2644,N_676,N_707);
nand U2645 (N_2645,N_5,N_1633);
nand U2646 (N_2646,N_301,N_850);
or U2647 (N_2647,N_1617,N_143);
nor U2648 (N_2648,N_314,N_451);
nor U2649 (N_2649,N_1658,N_340);
and U2650 (N_2650,N_1176,N_256);
nor U2651 (N_2651,N_49,N_617);
nor U2652 (N_2652,N_1978,N_1230);
or U2653 (N_2653,N_227,N_485);
nand U2654 (N_2654,N_664,N_412);
nand U2655 (N_2655,N_158,N_929);
nor U2656 (N_2656,N_1620,N_1438);
and U2657 (N_2657,N_263,N_231);
xnor U2658 (N_2658,N_883,N_243);
nand U2659 (N_2659,N_853,N_1511);
and U2660 (N_2660,N_1348,N_293);
nand U2661 (N_2661,N_125,N_1487);
nand U2662 (N_2662,N_302,N_235);
or U2663 (N_2663,N_1673,N_1275);
and U2664 (N_2664,N_354,N_643);
and U2665 (N_2665,N_1420,N_75);
and U2666 (N_2666,N_828,N_1861);
nor U2667 (N_2667,N_1794,N_106);
nand U2668 (N_2668,N_1935,N_1161);
or U2669 (N_2669,N_511,N_688);
or U2670 (N_2670,N_1134,N_1977);
nand U2671 (N_2671,N_410,N_902);
nor U2672 (N_2672,N_720,N_671);
xor U2673 (N_2673,N_79,N_1550);
nor U2674 (N_2674,N_891,N_1961);
nor U2675 (N_2675,N_443,N_669);
nor U2676 (N_2676,N_625,N_805);
or U2677 (N_2677,N_838,N_1939);
nand U2678 (N_2678,N_1762,N_1406);
nand U2679 (N_2679,N_417,N_740);
nand U2680 (N_2680,N_1034,N_1066);
and U2681 (N_2681,N_609,N_375);
nand U2682 (N_2682,N_1829,N_1646);
nor U2683 (N_2683,N_646,N_1967);
nand U2684 (N_2684,N_1044,N_544);
and U2685 (N_2685,N_280,N_903);
or U2686 (N_2686,N_1576,N_1602);
or U2687 (N_2687,N_1634,N_804);
xor U2688 (N_2688,N_542,N_1908);
xor U2689 (N_2689,N_1853,N_85);
xnor U2690 (N_2690,N_1761,N_1724);
nor U2691 (N_2691,N_312,N_1569);
nand U2692 (N_2692,N_428,N_1181);
nand U2693 (N_2693,N_638,N_8);
xnor U2694 (N_2694,N_852,N_1970);
and U2695 (N_2695,N_1364,N_623);
nand U2696 (N_2696,N_1417,N_948);
xor U2697 (N_2697,N_13,N_874);
or U2698 (N_2698,N_940,N_1224);
nor U2699 (N_2699,N_1429,N_1292);
or U2700 (N_2700,N_1943,N_1921);
and U2701 (N_2701,N_441,N_61);
nand U2702 (N_2702,N_1300,N_747);
or U2703 (N_2703,N_68,N_549);
nor U2704 (N_2704,N_1446,N_654);
and U2705 (N_2705,N_1088,N_363);
or U2706 (N_2706,N_1383,N_703);
nand U2707 (N_2707,N_396,N_316);
or U2708 (N_2708,N_545,N_1786);
xor U2709 (N_2709,N_46,N_1674);
nand U2710 (N_2710,N_1941,N_64);
and U2711 (N_2711,N_922,N_1150);
nand U2712 (N_2712,N_44,N_313);
or U2713 (N_2713,N_1354,N_1754);
nand U2714 (N_2714,N_1201,N_208);
nor U2715 (N_2715,N_1281,N_1280);
or U2716 (N_2716,N_47,N_516);
and U2717 (N_2717,N_557,N_209);
or U2718 (N_2718,N_1186,N_1495);
or U2719 (N_2719,N_1573,N_226);
and U2720 (N_2720,N_690,N_1306);
and U2721 (N_2721,N_1670,N_803);
nor U2722 (N_2722,N_1998,N_1886);
or U2723 (N_2723,N_1130,N_1465);
or U2724 (N_2724,N_553,N_1196);
nor U2725 (N_2725,N_453,N_768);
nand U2726 (N_2726,N_1301,N_655);
nand U2727 (N_2727,N_229,N_1195);
nor U2728 (N_2728,N_764,N_467);
and U2729 (N_2729,N_1513,N_603);
or U2730 (N_2730,N_1614,N_1604);
nand U2731 (N_2731,N_1236,N_309);
xnor U2732 (N_2732,N_171,N_1906);
nand U2733 (N_2733,N_743,N_810);
and U2734 (N_2734,N_1343,N_1811);
nand U2735 (N_2735,N_1596,N_1539);
and U2736 (N_2736,N_896,N_556);
nor U2737 (N_2737,N_907,N_1404);
nor U2738 (N_2738,N_48,N_715);
xnor U2739 (N_2739,N_618,N_347);
nor U2740 (N_2740,N_762,N_1026);
nand U2741 (N_2741,N_1867,N_584);
and U2742 (N_2742,N_1862,N_986);
and U2743 (N_2743,N_1669,N_1370);
nor U2744 (N_2744,N_1757,N_686);
nor U2745 (N_2745,N_1209,N_196);
xor U2746 (N_2746,N_217,N_1816);
or U2747 (N_2747,N_1041,N_1848);
xor U2748 (N_2748,N_1657,N_1499);
and U2749 (N_2749,N_1021,N_1727);
nand U2750 (N_2750,N_926,N_1627);
nor U2751 (N_2751,N_1748,N_656);
or U2752 (N_2752,N_1721,N_1432);
or U2753 (N_2753,N_1349,N_1063);
xnor U2754 (N_2754,N_1565,N_799);
and U2755 (N_2755,N_1111,N_1367);
or U2756 (N_2756,N_174,N_1426);
or U2757 (N_2757,N_1508,N_763);
or U2758 (N_2758,N_1211,N_1710);
nand U2759 (N_2759,N_1960,N_1001);
or U2760 (N_2760,N_1585,N_1342);
nor U2761 (N_2761,N_921,N_1652);
or U2762 (N_2762,N_1749,N_1046);
nand U2763 (N_2763,N_548,N_1671);
nand U2764 (N_2764,N_1008,N_218);
and U2765 (N_2765,N_9,N_1347);
xor U2766 (N_2766,N_724,N_1759);
and U2767 (N_2767,N_1142,N_966);
nor U2768 (N_2768,N_1979,N_1458);
and U2769 (N_2769,N_1640,N_1476);
or U2770 (N_2770,N_766,N_1564);
or U2771 (N_2771,N_1101,N_185);
nor U2772 (N_2772,N_615,N_1907);
nand U2773 (N_2773,N_305,N_1070);
nand U2774 (N_2774,N_1232,N_957);
nor U2775 (N_2775,N_1814,N_604);
nor U2776 (N_2776,N_1203,N_477);
nand U2777 (N_2777,N_120,N_536);
nand U2778 (N_2778,N_165,N_93);
xor U2779 (N_2779,N_494,N_560);
nor U2780 (N_2780,N_1336,N_822);
nand U2781 (N_2781,N_920,N_681);
xor U2782 (N_2782,N_956,N_1038);
and U2783 (N_2783,N_1474,N_1810);
nor U2784 (N_2784,N_1557,N_1953);
nor U2785 (N_2785,N_37,N_1259);
nand U2786 (N_2786,N_390,N_847);
or U2787 (N_2787,N_1017,N_884);
nand U2788 (N_2788,N_587,N_1217);
and U2789 (N_2789,N_291,N_268);
or U2790 (N_2790,N_504,N_540);
xnor U2791 (N_2791,N_401,N_1898);
or U2792 (N_2792,N_1461,N_974);
and U2793 (N_2793,N_612,N_205);
and U2794 (N_2794,N_1304,N_194);
nor U2795 (N_2795,N_509,N_1210);
nor U2796 (N_2796,N_586,N_1789);
and U2797 (N_2797,N_199,N_543);
nand U2798 (N_2798,N_945,N_1933);
nor U2799 (N_2799,N_1702,N_446);
nor U2800 (N_2800,N_1120,N_483);
or U2801 (N_2801,N_1575,N_372);
or U2802 (N_2802,N_576,N_1925);
nand U2803 (N_2803,N_1043,N_1878);
and U2804 (N_2804,N_756,N_1250);
nand U2805 (N_2805,N_290,N_1055);
and U2806 (N_2806,N_836,N_1425);
nor U2807 (N_2807,N_1993,N_317);
or U2808 (N_2808,N_1106,N_812);
nor U2809 (N_2809,N_1079,N_40);
nand U2810 (N_2810,N_658,N_1858);
and U2811 (N_2811,N_297,N_1214);
xor U2812 (N_2812,N_1170,N_933);
and U2813 (N_2813,N_736,N_1341);
xor U2814 (N_2814,N_378,N_683);
nor U2815 (N_2815,N_1859,N_785);
and U2816 (N_2816,N_1479,N_224);
nand U2817 (N_2817,N_91,N_761);
nor U2818 (N_2818,N_414,N_1050);
and U2819 (N_2819,N_1302,N_1262);
and U2820 (N_2820,N_183,N_1683);
nor U2821 (N_2821,N_1997,N_1064);
nor U2822 (N_2822,N_1204,N_271);
nor U2823 (N_2823,N_421,N_1864);
or U2824 (N_2824,N_1716,N_1362);
and U2825 (N_2825,N_1791,N_41);
nand U2826 (N_2826,N_1378,N_402);
or U2827 (N_2827,N_1974,N_1817);
nand U2828 (N_2828,N_1463,N_389);
and U2829 (N_2829,N_1192,N_1258);
or U2830 (N_2830,N_14,N_1199);
nand U2831 (N_2831,N_471,N_1153);
xnor U2832 (N_2832,N_1947,N_1489);
or U2833 (N_2833,N_1624,N_191);
nand U2834 (N_2834,N_444,N_324);
and U2835 (N_2835,N_1592,N_122);
or U2836 (N_2836,N_1715,N_968);
and U2837 (N_2837,N_640,N_339);
nand U2838 (N_2838,N_121,N_781);
and U2839 (N_2839,N_1057,N_42);
and U2840 (N_2840,N_1319,N_653);
nand U2841 (N_2841,N_1801,N_1984);
nor U2842 (N_2842,N_1622,N_1385);
nor U2843 (N_2843,N_611,N_565);
or U2844 (N_2844,N_82,N_927);
nand U2845 (N_2845,N_709,N_644);
nand U2846 (N_2846,N_1770,N_131);
nand U2847 (N_2847,N_383,N_398);
nor U2848 (N_2848,N_809,N_127);
xor U2849 (N_2849,N_825,N_1605);
xor U2850 (N_2850,N_1318,N_1094);
nand U2851 (N_2851,N_1277,N_600);
and U2852 (N_2852,N_1355,N_1874);
nand U2853 (N_2853,N_306,N_1732);
and U2854 (N_2854,N_1561,N_94);
and U2855 (N_2855,N_220,N_1313);
nand U2856 (N_2856,N_1797,N_1491);
nor U2857 (N_2857,N_985,N_367);
nor U2858 (N_2858,N_972,N_1995);
nor U2859 (N_2859,N_1069,N_1515);
nor U2860 (N_2860,N_234,N_1850);
or U2861 (N_2861,N_895,N_627);
xor U2862 (N_2862,N_1536,N_1222);
or U2863 (N_2863,N_1818,N_408);
or U2864 (N_2864,N_823,N_52);
nor U2865 (N_2865,N_684,N_1831);
or U2866 (N_2866,N_541,N_338);
and U2867 (N_2867,N_379,N_994);
xnor U2868 (N_2868,N_452,N_1656);
nor U2869 (N_2869,N_1823,N_95);
nand U2870 (N_2870,N_1660,N_1076);
and U2871 (N_2871,N_1462,N_1870);
or U2872 (N_2872,N_357,N_734);
nand U2873 (N_2873,N_461,N_1840);
or U2874 (N_2874,N_1009,N_1679);
and U2875 (N_2875,N_1725,N_25);
nor U2876 (N_2876,N_760,N_16);
and U2877 (N_2877,N_1371,N_1325);
nand U2878 (N_2878,N_1700,N_1218);
nand U2879 (N_2879,N_1975,N_608);
and U2880 (N_2880,N_1745,N_1030);
xor U2881 (N_2881,N_180,N_1985);
nand U2882 (N_2882,N_1586,N_1036);
nor U2883 (N_2883,N_299,N_1856);
nor U2884 (N_2884,N_1174,N_1616);
and U2885 (N_2885,N_1405,N_1659);
and U2886 (N_2886,N_775,N_613);
xor U2887 (N_2887,N_1291,N_665);
or U2888 (N_2888,N_1330,N_1597);
nor U2889 (N_2889,N_1469,N_181);
or U2890 (N_2890,N_573,N_368);
or U2891 (N_2891,N_296,N_113);
and U2892 (N_2892,N_1973,N_1299);
nor U2893 (N_2893,N_559,N_1666);
and U2894 (N_2894,N_214,N_863);
or U2895 (N_2895,N_1480,N_343);
nand U2896 (N_2896,N_1706,N_1545);
or U2897 (N_2897,N_384,N_1455);
nand U2898 (N_2898,N_1241,N_1785);
or U2899 (N_2899,N_1552,N_531);
nor U2900 (N_2900,N_463,N_54);
and U2901 (N_2901,N_817,N_1832);
or U2902 (N_2902,N_1278,N_248);
nor U2903 (N_2903,N_388,N_1252);
nor U2904 (N_2904,N_1244,N_1344);
nand U2905 (N_2905,N_1045,N_1574);
nand U2906 (N_2906,N_1171,N_845);
nor U2907 (N_2907,N_489,N_1746);
nor U2908 (N_2908,N_1338,N_1143);
and U2909 (N_2909,N_315,N_702);
and U2910 (N_2910,N_677,N_1952);
nand U2911 (N_2911,N_330,N_1582);
xnor U2912 (N_2912,N_514,N_284);
or U2913 (N_2913,N_212,N_815);
nand U2914 (N_2914,N_897,N_495);
nor U2915 (N_2915,N_295,N_1873);
nor U2916 (N_2916,N_1999,N_1712);
or U2917 (N_2917,N_1568,N_1137);
nor U2918 (N_2918,N_502,N_188);
nand U2919 (N_2919,N_1290,N_1877);
xnor U2920 (N_2920,N_1128,N_572);
nor U2921 (N_2921,N_1623,N_1115);
xor U2922 (N_2922,N_465,N_1894);
nand U2923 (N_2923,N_949,N_356);
nand U2924 (N_2924,N_1734,N_1587);
nand U2925 (N_2925,N_1067,N_727);
or U2926 (N_2926,N_621,N_136);
or U2927 (N_2927,N_1359,N_563);
nor U2928 (N_2928,N_1116,N_407);
and U2929 (N_2929,N_1882,N_508);
xnor U2930 (N_2930,N_1206,N_1693);
or U2931 (N_2931,N_1065,N_332);
nor U2932 (N_2932,N_814,N_1600);
and U2933 (N_2933,N_651,N_1541);
nand U2934 (N_2934,N_1221,N_1723);
or U2935 (N_2935,N_977,N_988);
or U2936 (N_2936,N_1098,N_427);
nand U2937 (N_2937,N_1394,N_1311);
or U2938 (N_2938,N_1841,N_335);
nand U2939 (N_2939,N_1948,N_928);
xnor U2940 (N_2940,N_503,N_475);
nor U2941 (N_2941,N_140,N_779);
and U2942 (N_2942,N_1003,N_250);
xor U2943 (N_2943,N_67,N_1421);
nand U2944 (N_2944,N_360,N_1667);
or U2945 (N_2945,N_1190,N_109);
and U2946 (N_2946,N_796,N_1990);
nor U2947 (N_2947,N_72,N_1510);
or U2948 (N_2948,N_459,N_310);
and U2949 (N_2949,N_1957,N_1606);
or U2950 (N_2950,N_1047,N_153);
xor U2951 (N_2951,N_1507,N_1382);
and U2952 (N_2952,N_959,N_1692);
xnor U2953 (N_2953,N_864,N_663);
nand U2954 (N_2954,N_1140,N_551);
nand U2955 (N_2955,N_1729,N_260);
and U2956 (N_2956,N_31,N_1849);
nor U2957 (N_2957,N_858,N_65);
and U2958 (N_2958,N_1314,N_1496);
nand U2959 (N_2959,N_934,N_539);
nor U2960 (N_2960,N_117,N_913);
or U2961 (N_2961,N_159,N_1572);
and U2962 (N_2962,N_1983,N_1981);
and U2963 (N_2963,N_670,N_622);
or U2964 (N_2964,N_1888,N_591);
nor U2965 (N_2965,N_1664,N_1528);
nand U2966 (N_2966,N_114,N_1339);
xnor U2967 (N_2967,N_1460,N_1025);
nor U2968 (N_2968,N_955,N_124);
or U2969 (N_2969,N_1484,N_322);
and U2970 (N_2970,N_1833,N_1986);
nor U2971 (N_2971,N_1219,N_333);
nor U2972 (N_2972,N_253,N_1726);
xor U2973 (N_2973,N_552,N_152);
nand U2974 (N_2974,N_393,N_635);
and U2975 (N_2975,N_1753,N_1135);
and U2976 (N_2976,N_491,N_1289);
or U2977 (N_2977,N_1684,N_1675);
or U2978 (N_2978,N_816,N_1739);
nand U2979 (N_2979,N_276,N_711);
and U2980 (N_2980,N_1924,N_975);
xnor U2981 (N_2981,N_1522,N_488);
and U2982 (N_2982,N_881,N_1430);
nand U2983 (N_2983,N_910,N_1369);
nor U2984 (N_2984,N_348,N_1733);
and U2985 (N_2985,N_1077,N_639);
and U2986 (N_2986,N_1074,N_1642);
nor U2987 (N_2987,N_1891,N_1273);
and U2988 (N_2988,N_538,N_1152);
xnor U2989 (N_2989,N_704,N_1331);
nand U2990 (N_2990,N_1824,N_851);
nand U2991 (N_2991,N_80,N_1018);
or U2992 (N_2992,N_1033,N_395);
and U2993 (N_2993,N_1388,N_513);
and U2994 (N_2994,N_439,N_1335);
or U2995 (N_2995,N_636,N_1807);
nand U2996 (N_2996,N_1892,N_424);
nor U2997 (N_2997,N_162,N_1024);
xnor U2998 (N_2998,N_431,N_1478);
or U2999 (N_2999,N_1538,N_866);
nor U3000 (N_3000,N_247,N_959);
and U3001 (N_3001,N_312,N_1818);
and U3002 (N_3002,N_1735,N_1206);
xnor U3003 (N_3003,N_1429,N_429);
or U3004 (N_3004,N_269,N_1176);
and U3005 (N_3005,N_231,N_1557);
or U3006 (N_3006,N_577,N_865);
nand U3007 (N_3007,N_701,N_345);
or U3008 (N_3008,N_1822,N_250);
xnor U3009 (N_3009,N_869,N_48);
and U3010 (N_3010,N_1843,N_169);
or U3011 (N_3011,N_1711,N_974);
and U3012 (N_3012,N_1722,N_971);
nand U3013 (N_3013,N_316,N_1844);
nor U3014 (N_3014,N_1051,N_122);
or U3015 (N_3015,N_343,N_120);
nor U3016 (N_3016,N_1392,N_1377);
nand U3017 (N_3017,N_1862,N_535);
nor U3018 (N_3018,N_1427,N_545);
nand U3019 (N_3019,N_1146,N_91);
or U3020 (N_3020,N_1378,N_581);
nor U3021 (N_3021,N_690,N_1668);
or U3022 (N_3022,N_388,N_9);
nor U3023 (N_3023,N_1870,N_1523);
nor U3024 (N_3024,N_934,N_1142);
and U3025 (N_3025,N_233,N_288);
and U3026 (N_3026,N_1049,N_1898);
or U3027 (N_3027,N_1983,N_1140);
or U3028 (N_3028,N_1301,N_1513);
or U3029 (N_3029,N_1394,N_712);
nor U3030 (N_3030,N_1685,N_712);
and U3031 (N_3031,N_1698,N_514);
nand U3032 (N_3032,N_677,N_1212);
nand U3033 (N_3033,N_1296,N_765);
and U3034 (N_3034,N_1672,N_60);
or U3035 (N_3035,N_1571,N_298);
or U3036 (N_3036,N_1974,N_1553);
nor U3037 (N_3037,N_179,N_551);
nand U3038 (N_3038,N_939,N_240);
and U3039 (N_3039,N_248,N_1488);
nand U3040 (N_3040,N_1822,N_1162);
nor U3041 (N_3041,N_560,N_699);
or U3042 (N_3042,N_658,N_1280);
or U3043 (N_3043,N_223,N_1365);
xor U3044 (N_3044,N_1722,N_1221);
and U3045 (N_3045,N_600,N_111);
nor U3046 (N_3046,N_1513,N_1322);
or U3047 (N_3047,N_1508,N_882);
and U3048 (N_3048,N_1279,N_1270);
and U3049 (N_3049,N_501,N_1212);
nand U3050 (N_3050,N_1373,N_286);
or U3051 (N_3051,N_1520,N_1018);
nand U3052 (N_3052,N_171,N_1777);
nand U3053 (N_3053,N_18,N_195);
nor U3054 (N_3054,N_214,N_1369);
nor U3055 (N_3055,N_1951,N_900);
nor U3056 (N_3056,N_1984,N_112);
and U3057 (N_3057,N_1204,N_875);
and U3058 (N_3058,N_1813,N_1746);
nor U3059 (N_3059,N_158,N_1846);
or U3060 (N_3060,N_1764,N_438);
and U3061 (N_3061,N_1085,N_161);
xor U3062 (N_3062,N_1231,N_426);
and U3063 (N_3063,N_1257,N_4);
nor U3064 (N_3064,N_1967,N_660);
or U3065 (N_3065,N_385,N_1174);
and U3066 (N_3066,N_191,N_992);
or U3067 (N_3067,N_1194,N_831);
nand U3068 (N_3068,N_840,N_278);
or U3069 (N_3069,N_1039,N_302);
xor U3070 (N_3070,N_1857,N_1116);
and U3071 (N_3071,N_550,N_1862);
xor U3072 (N_3072,N_1340,N_12);
nor U3073 (N_3073,N_1782,N_681);
and U3074 (N_3074,N_498,N_538);
and U3075 (N_3075,N_580,N_1490);
nor U3076 (N_3076,N_1107,N_1686);
or U3077 (N_3077,N_1000,N_541);
nand U3078 (N_3078,N_999,N_931);
or U3079 (N_3079,N_1525,N_1415);
xnor U3080 (N_3080,N_662,N_499);
and U3081 (N_3081,N_928,N_1901);
nand U3082 (N_3082,N_937,N_978);
or U3083 (N_3083,N_1566,N_1509);
nor U3084 (N_3084,N_293,N_107);
and U3085 (N_3085,N_1250,N_81);
nor U3086 (N_3086,N_1430,N_122);
and U3087 (N_3087,N_1570,N_1575);
xnor U3088 (N_3088,N_996,N_1015);
nor U3089 (N_3089,N_1535,N_1370);
nor U3090 (N_3090,N_1475,N_145);
nor U3091 (N_3091,N_1888,N_216);
nand U3092 (N_3092,N_1858,N_1580);
or U3093 (N_3093,N_1501,N_672);
nor U3094 (N_3094,N_1646,N_38);
nand U3095 (N_3095,N_1763,N_490);
nand U3096 (N_3096,N_1196,N_513);
nand U3097 (N_3097,N_774,N_1768);
nor U3098 (N_3098,N_126,N_501);
and U3099 (N_3099,N_119,N_1969);
xor U3100 (N_3100,N_1371,N_417);
and U3101 (N_3101,N_1873,N_535);
nand U3102 (N_3102,N_594,N_810);
nor U3103 (N_3103,N_1207,N_1323);
and U3104 (N_3104,N_1324,N_693);
or U3105 (N_3105,N_102,N_456);
nor U3106 (N_3106,N_699,N_12);
and U3107 (N_3107,N_583,N_1976);
nand U3108 (N_3108,N_676,N_786);
nor U3109 (N_3109,N_130,N_1045);
nand U3110 (N_3110,N_1969,N_155);
or U3111 (N_3111,N_601,N_1146);
or U3112 (N_3112,N_104,N_627);
nor U3113 (N_3113,N_112,N_1676);
or U3114 (N_3114,N_807,N_1866);
and U3115 (N_3115,N_808,N_1336);
nand U3116 (N_3116,N_852,N_1702);
and U3117 (N_3117,N_1535,N_68);
nand U3118 (N_3118,N_1956,N_1946);
or U3119 (N_3119,N_663,N_1570);
nor U3120 (N_3120,N_1818,N_884);
xor U3121 (N_3121,N_430,N_239);
and U3122 (N_3122,N_128,N_1026);
and U3123 (N_3123,N_1189,N_33);
or U3124 (N_3124,N_738,N_996);
or U3125 (N_3125,N_969,N_59);
or U3126 (N_3126,N_69,N_162);
and U3127 (N_3127,N_934,N_1812);
or U3128 (N_3128,N_284,N_1322);
or U3129 (N_3129,N_270,N_1023);
and U3130 (N_3130,N_8,N_31);
or U3131 (N_3131,N_374,N_1830);
and U3132 (N_3132,N_413,N_884);
nor U3133 (N_3133,N_1556,N_448);
nand U3134 (N_3134,N_876,N_1923);
or U3135 (N_3135,N_1416,N_1195);
nor U3136 (N_3136,N_17,N_1825);
nor U3137 (N_3137,N_249,N_427);
nand U3138 (N_3138,N_1900,N_861);
or U3139 (N_3139,N_645,N_1627);
or U3140 (N_3140,N_1514,N_798);
or U3141 (N_3141,N_1522,N_823);
and U3142 (N_3142,N_1344,N_446);
or U3143 (N_3143,N_504,N_933);
or U3144 (N_3144,N_26,N_1394);
nand U3145 (N_3145,N_275,N_626);
xor U3146 (N_3146,N_754,N_682);
and U3147 (N_3147,N_3,N_1997);
and U3148 (N_3148,N_1417,N_1766);
nand U3149 (N_3149,N_80,N_1685);
xor U3150 (N_3150,N_921,N_1618);
and U3151 (N_3151,N_1841,N_1657);
and U3152 (N_3152,N_942,N_1395);
and U3153 (N_3153,N_1346,N_1599);
or U3154 (N_3154,N_1345,N_1984);
nor U3155 (N_3155,N_1343,N_1130);
nand U3156 (N_3156,N_1263,N_1078);
xnor U3157 (N_3157,N_793,N_49);
and U3158 (N_3158,N_172,N_1466);
or U3159 (N_3159,N_1159,N_1505);
nor U3160 (N_3160,N_1277,N_1111);
xnor U3161 (N_3161,N_1219,N_14);
or U3162 (N_3162,N_1842,N_1971);
nand U3163 (N_3163,N_1313,N_1651);
nand U3164 (N_3164,N_64,N_1118);
nand U3165 (N_3165,N_1185,N_192);
nor U3166 (N_3166,N_1375,N_13);
nor U3167 (N_3167,N_114,N_27);
nor U3168 (N_3168,N_816,N_110);
nor U3169 (N_3169,N_604,N_125);
or U3170 (N_3170,N_731,N_27);
xor U3171 (N_3171,N_1986,N_198);
nor U3172 (N_3172,N_540,N_125);
or U3173 (N_3173,N_1877,N_1965);
nor U3174 (N_3174,N_960,N_1393);
nor U3175 (N_3175,N_1551,N_1929);
and U3176 (N_3176,N_1590,N_1115);
nand U3177 (N_3177,N_1970,N_502);
nand U3178 (N_3178,N_731,N_380);
and U3179 (N_3179,N_1799,N_1493);
nor U3180 (N_3180,N_808,N_1650);
xor U3181 (N_3181,N_1057,N_210);
or U3182 (N_3182,N_120,N_1190);
or U3183 (N_3183,N_1947,N_1173);
nand U3184 (N_3184,N_32,N_673);
and U3185 (N_3185,N_272,N_430);
nor U3186 (N_3186,N_525,N_1213);
or U3187 (N_3187,N_1502,N_1106);
nor U3188 (N_3188,N_1428,N_1589);
nand U3189 (N_3189,N_708,N_1162);
and U3190 (N_3190,N_220,N_1949);
nor U3191 (N_3191,N_1520,N_170);
and U3192 (N_3192,N_1806,N_1729);
nor U3193 (N_3193,N_1234,N_1958);
and U3194 (N_3194,N_519,N_418);
and U3195 (N_3195,N_749,N_1944);
and U3196 (N_3196,N_112,N_1220);
or U3197 (N_3197,N_497,N_1053);
or U3198 (N_3198,N_1878,N_1299);
and U3199 (N_3199,N_1654,N_150);
or U3200 (N_3200,N_1020,N_1727);
or U3201 (N_3201,N_242,N_540);
nand U3202 (N_3202,N_1214,N_1992);
nor U3203 (N_3203,N_1218,N_1864);
xor U3204 (N_3204,N_197,N_1555);
and U3205 (N_3205,N_749,N_1492);
xnor U3206 (N_3206,N_1779,N_1148);
or U3207 (N_3207,N_687,N_486);
and U3208 (N_3208,N_1457,N_781);
and U3209 (N_3209,N_1636,N_55);
or U3210 (N_3210,N_845,N_1206);
and U3211 (N_3211,N_242,N_375);
nor U3212 (N_3212,N_1704,N_1897);
nand U3213 (N_3213,N_1061,N_1824);
and U3214 (N_3214,N_1907,N_1480);
nand U3215 (N_3215,N_708,N_961);
nand U3216 (N_3216,N_363,N_1952);
xor U3217 (N_3217,N_940,N_1056);
nor U3218 (N_3218,N_1249,N_1350);
nand U3219 (N_3219,N_506,N_265);
nand U3220 (N_3220,N_1134,N_1905);
nand U3221 (N_3221,N_1485,N_693);
or U3222 (N_3222,N_1729,N_1758);
and U3223 (N_3223,N_700,N_550);
nand U3224 (N_3224,N_1860,N_497);
or U3225 (N_3225,N_1327,N_129);
nand U3226 (N_3226,N_160,N_1640);
xnor U3227 (N_3227,N_1235,N_109);
nand U3228 (N_3228,N_1154,N_1782);
or U3229 (N_3229,N_440,N_1340);
xor U3230 (N_3230,N_1503,N_1214);
or U3231 (N_3231,N_1588,N_1550);
nor U3232 (N_3232,N_859,N_801);
or U3233 (N_3233,N_124,N_874);
and U3234 (N_3234,N_705,N_1148);
or U3235 (N_3235,N_116,N_1540);
nand U3236 (N_3236,N_1832,N_1312);
or U3237 (N_3237,N_793,N_776);
nand U3238 (N_3238,N_256,N_1256);
nor U3239 (N_3239,N_1784,N_438);
and U3240 (N_3240,N_129,N_1048);
xnor U3241 (N_3241,N_1746,N_210);
nand U3242 (N_3242,N_849,N_1366);
xor U3243 (N_3243,N_1275,N_965);
and U3244 (N_3244,N_1114,N_532);
nand U3245 (N_3245,N_1100,N_405);
and U3246 (N_3246,N_324,N_1694);
and U3247 (N_3247,N_1062,N_92);
or U3248 (N_3248,N_1176,N_56);
or U3249 (N_3249,N_19,N_1157);
and U3250 (N_3250,N_329,N_1792);
or U3251 (N_3251,N_1980,N_1582);
or U3252 (N_3252,N_191,N_861);
nand U3253 (N_3253,N_1691,N_376);
and U3254 (N_3254,N_806,N_127);
nor U3255 (N_3255,N_828,N_41);
and U3256 (N_3256,N_494,N_1275);
xor U3257 (N_3257,N_529,N_51);
nor U3258 (N_3258,N_291,N_245);
nand U3259 (N_3259,N_44,N_1869);
nand U3260 (N_3260,N_403,N_1910);
or U3261 (N_3261,N_600,N_1956);
nand U3262 (N_3262,N_192,N_112);
xnor U3263 (N_3263,N_1233,N_1199);
or U3264 (N_3264,N_673,N_15);
nor U3265 (N_3265,N_655,N_1536);
or U3266 (N_3266,N_1673,N_1753);
nand U3267 (N_3267,N_1639,N_906);
and U3268 (N_3268,N_1659,N_1430);
nor U3269 (N_3269,N_895,N_154);
nand U3270 (N_3270,N_1882,N_912);
and U3271 (N_3271,N_54,N_600);
nand U3272 (N_3272,N_1285,N_1338);
xnor U3273 (N_3273,N_745,N_951);
or U3274 (N_3274,N_1234,N_585);
nor U3275 (N_3275,N_538,N_570);
and U3276 (N_3276,N_900,N_424);
and U3277 (N_3277,N_203,N_227);
nor U3278 (N_3278,N_1267,N_1052);
and U3279 (N_3279,N_1708,N_232);
nand U3280 (N_3280,N_744,N_556);
and U3281 (N_3281,N_1506,N_1718);
and U3282 (N_3282,N_138,N_795);
nand U3283 (N_3283,N_475,N_205);
nand U3284 (N_3284,N_1404,N_1333);
nor U3285 (N_3285,N_793,N_78);
or U3286 (N_3286,N_119,N_190);
nor U3287 (N_3287,N_802,N_1824);
nand U3288 (N_3288,N_1933,N_333);
and U3289 (N_3289,N_1798,N_1692);
nand U3290 (N_3290,N_1549,N_815);
and U3291 (N_3291,N_1975,N_1039);
and U3292 (N_3292,N_1775,N_1902);
or U3293 (N_3293,N_1663,N_1706);
nand U3294 (N_3294,N_854,N_507);
nor U3295 (N_3295,N_1791,N_232);
and U3296 (N_3296,N_1004,N_1526);
nand U3297 (N_3297,N_1765,N_1025);
nor U3298 (N_3298,N_1964,N_1366);
nor U3299 (N_3299,N_1812,N_749);
nand U3300 (N_3300,N_217,N_916);
nand U3301 (N_3301,N_1445,N_1024);
xor U3302 (N_3302,N_654,N_439);
xor U3303 (N_3303,N_656,N_1098);
nor U3304 (N_3304,N_105,N_1198);
xnor U3305 (N_3305,N_1001,N_1595);
or U3306 (N_3306,N_543,N_82);
or U3307 (N_3307,N_1158,N_125);
nor U3308 (N_3308,N_451,N_751);
nor U3309 (N_3309,N_1901,N_66);
nand U3310 (N_3310,N_124,N_440);
xor U3311 (N_3311,N_428,N_1559);
nor U3312 (N_3312,N_1454,N_687);
nand U3313 (N_3313,N_136,N_518);
and U3314 (N_3314,N_1980,N_372);
nand U3315 (N_3315,N_1476,N_1030);
and U3316 (N_3316,N_616,N_105);
nor U3317 (N_3317,N_1969,N_1304);
or U3318 (N_3318,N_331,N_1032);
or U3319 (N_3319,N_1450,N_518);
nand U3320 (N_3320,N_814,N_501);
and U3321 (N_3321,N_676,N_353);
or U3322 (N_3322,N_170,N_849);
or U3323 (N_3323,N_116,N_1372);
nand U3324 (N_3324,N_433,N_1910);
xnor U3325 (N_3325,N_898,N_19);
or U3326 (N_3326,N_318,N_1951);
and U3327 (N_3327,N_521,N_637);
nand U3328 (N_3328,N_235,N_1638);
xor U3329 (N_3329,N_1532,N_1358);
nand U3330 (N_3330,N_80,N_1613);
nand U3331 (N_3331,N_108,N_254);
nor U3332 (N_3332,N_1676,N_1347);
or U3333 (N_3333,N_1451,N_1907);
nor U3334 (N_3334,N_1031,N_1613);
nand U3335 (N_3335,N_731,N_900);
nand U3336 (N_3336,N_1102,N_578);
nor U3337 (N_3337,N_518,N_1017);
nand U3338 (N_3338,N_207,N_324);
and U3339 (N_3339,N_1763,N_1285);
nand U3340 (N_3340,N_1963,N_855);
nor U3341 (N_3341,N_1296,N_562);
nor U3342 (N_3342,N_557,N_581);
xnor U3343 (N_3343,N_493,N_1271);
nand U3344 (N_3344,N_1512,N_1325);
nand U3345 (N_3345,N_486,N_1355);
xor U3346 (N_3346,N_1169,N_1667);
nor U3347 (N_3347,N_1775,N_549);
nand U3348 (N_3348,N_1386,N_1776);
nor U3349 (N_3349,N_786,N_991);
nor U3350 (N_3350,N_94,N_1063);
nand U3351 (N_3351,N_404,N_1584);
nand U3352 (N_3352,N_1123,N_1980);
nand U3353 (N_3353,N_1589,N_1011);
or U3354 (N_3354,N_1728,N_535);
or U3355 (N_3355,N_1529,N_410);
xor U3356 (N_3356,N_1412,N_322);
nor U3357 (N_3357,N_294,N_1271);
or U3358 (N_3358,N_547,N_1256);
nor U3359 (N_3359,N_630,N_1451);
nand U3360 (N_3360,N_832,N_622);
xnor U3361 (N_3361,N_325,N_680);
nand U3362 (N_3362,N_534,N_252);
nand U3363 (N_3363,N_1767,N_876);
and U3364 (N_3364,N_825,N_23);
nand U3365 (N_3365,N_1812,N_505);
and U3366 (N_3366,N_455,N_375);
nor U3367 (N_3367,N_1481,N_1519);
nor U3368 (N_3368,N_1803,N_387);
nand U3369 (N_3369,N_123,N_356);
nand U3370 (N_3370,N_739,N_1561);
nand U3371 (N_3371,N_641,N_1444);
nand U3372 (N_3372,N_303,N_1609);
or U3373 (N_3373,N_1064,N_321);
and U3374 (N_3374,N_1699,N_641);
xnor U3375 (N_3375,N_1732,N_798);
nor U3376 (N_3376,N_1744,N_59);
xor U3377 (N_3377,N_1055,N_1242);
xnor U3378 (N_3378,N_308,N_267);
xnor U3379 (N_3379,N_972,N_214);
and U3380 (N_3380,N_1749,N_1829);
or U3381 (N_3381,N_371,N_473);
and U3382 (N_3382,N_124,N_264);
nor U3383 (N_3383,N_926,N_1593);
or U3384 (N_3384,N_1328,N_871);
nand U3385 (N_3385,N_1156,N_1304);
nor U3386 (N_3386,N_1435,N_1690);
or U3387 (N_3387,N_1743,N_1868);
or U3388 (N_3388,N_722,N_412);
or U3389 (N_3389,N_1341,N_973);
nand U3390 (N_3390,N_93,N_831);
and U3391 (N_3391,N_517,N_915);
xnor U3392 (N_3392,N_1107,N_1996);
xor U3393 (N_3393,N_1528,N_12);
nor U3394 (N_3394,N_1611,N_1162);
or U3395 (N_3395,N_1150,N_1934);
or U3396 (N_3396,N_1680,N_1076);
and U3397 (N_3397,N_977,N_1141);
and U3398 (N_3398,N_673,N_1838);
or U3399 (N_3399,N_669,N_1903);
nor U3400 (N_3400,N_784,N_1070);
nor U3401 (N_3401,N_1943,N_210);
nor U3402 (N_3402,N_1332,N_1252);
nand U3403 (N_3403,N_1038,N_533);
or U3404 (N_3404,N_97,N_1376);
nand U3405 (N_3405,N_850,N_1933);
nor U3406 (N_3406,N_592,N_700);
or U3407 (N_3407,N_175,N_1380);
or U3408 (N_3408,N_101,N_612);
xor U3409 (N_3409,N_1270,N_628);
nand U3410 (N_3410,N_171,N_327);
and U3411 (N_3411,N_1337,N_1410);
or U3412 (N_3412,N_444,N_100);
and U3413 (N_3413,N_874,N_147);
and U3414 (N_3414,N_1613,N_1435);
nand U3415 (N_3415,N_1192,N_1161);
or U3416 (N_3416,N_1220,N_328);
or U3417 (N_3417,N_1858,N_603);
nand U3418 (N_3418,N_1522,N_1424);
or U3419 (N_3419,N_538,N_173);
nand U3420 (N_3420,N_193,N_351);
nand U3421 (N_3421,N_101,N_1045);
or U3422 (N_3422,N_170,N_135);
or U3423 (N_3423,N_255,N_295);
xor U3424 (N_3424,N_473,N_182);
xor U3425 (N_3425,N_141,N_1514);
nand U3426 (N_3426,N_1310,N_894);
and U3427 (N_3427,N_768,N_1125);
or U3428 (N_3428,N_1839,N_272);
and U3429 (N_3429,N_1615,N_25);
or U3430 (N_3430,N_617,N_1482);
nand U3431 (N_3431,N_694,N_1591);
or U3432 (N_3432,N_1453,N_863);
and U3433 (N_3433,N_1531,N_267);
and U3434 (N_3434,N_456,N_959);
xnor U3435 (N_3435,N_1025,N_1614);
and U3436 (N_3436,N_421,N_587);
and U3437 (N_3437,N_113,N_1410);
or U3438 (N_3438,N_549,N_285);
nand U3439 (N_3439,N_877,N_551);
and U3440 (N_3440,N_1133,N_1017);
xnor U3441 (N_3441,N_1431,N_1331);
or U3442 (N_3442,N_1451,N_129);
xnor U3443 (N_3443,N_1722,N_385);
nand U3444 (N_3444,N_1882,N_221);
nor U3445 (N_3445,N_1246,N_36);
nor U3446 (N_3446,N_1050,N_323);
xnor U3447 (N_3447,N_1138,N_1180);
nand U3448 (N_3448,N_1337,N_1838);
nor U3449 (N_3449,N_949,N_533);
nor U3450 (N_3450,N_1394,N_1365);
nand U3451 (N_3451,N_1598,N_1021);
and U3452 (N_3452,N_1752,N_685);
xnor U3453 (N_3453,N_1144,N_553);
and U3454 (N_3454,N_1647,N_703);
nand U3455 (N_3455,N_499,N_95);
xor U3456 (N_3456,N_1074,N_1252);
xnor U3457 (N_3457,N_823,N_1858);
nand U3458 (N_3458,N_1677,N_1055);
or U3459 (N_3459,N_130,N_865);
and U3460 (N_3460,N_128,N_1233);
and U3461 (N_3461,N_1032,N_155);
and U3462 (N_3462,N_792,N_1564);
nor U3463 (N_3463,N_623,N_255);
or U3464 (N_3464,N_714,N_1927);
and U3465 (N_3465,N_56,N_1253);
or U3466 (N_3466,N_1626,N_1230);
and U3467 (N_3467,N_936,N_159);
nand U3468 (N_3468,N_474,N_145);
xnor U3469 (N_3469,N_1171,N_1525);
xor U3470 (N_3470,N_307,N_1874);
or U3471 (N_3471,N_107,N_1692);
nand U3472 (N_3472,N_1817,N_698);
and U3473 (N_3473,N_191,N_1527);
or U3474 (N_3474,N_1304,N_221);
and U3475 (N_3475,N_855,N_1813);
nand U3476 (N_3476,N_1841,N_362);
nor U3477 (N_3477,N_613,N_1009);
and U3478 (N_3478,N_269,N_766);
xnor U3479 (N_3479,N_118,N_1155);
or U3480 (N_3480,N_24,N_90);
or U3481 (N_3481,N_1695,N_1805);
xnor U3482 (N_3482,N_1233,N_115);
nor U3483 (N_3483,N_823,N_1133);
or U3484 (N_3484,N_594,N_1313);
nor U3485 (N_3485,N_466,N_516);
nand U3486 (N_3486,N_775,N_1499);
and U3487 (N_3487,N_913,N_1251);
and U3488 (N_3488,N_1174,N_1654);
and U3489 (N_3489,N_1382,N_1380);
or U3490 (N_3490,N_284,N_383);
nor U3491 (N_3491,N_1088,N_1282);
and U3492 (N_3492,N_1533,N_1914);
or U3493 (N_3493,N_1299,N_856);
nor U3494 (N_3494,N_483,N_936);
and U3495 (N_3495,N_578,N_591);
xnor U3496 (N_3496,N_965,N_976);
nor U3497 (N_3497,N_1702,N_249);
and U3498 (N_3498,N_1097,N_216);
and U3499 (N_3499,N_1541,N_1722);
or U3500 (N_3500,N_247,N_1578);
or U3501 (N_3501,N_1636,N_1432);
and U3502 (N_3502,N_1533,N_1697);
or U3503 (N_3503,N_23,N_182);
or U3504 (N_3504,N_90,N_1610);
nand U3505 (N_3505,N_755,N_481);
and U3506 (N_3506,N_1708,N_1806);
nor U3507 (N_3507,N_352,N_1030);
and U3508 (N_3508,N_630,N_1116);
or U3509 (N_3509,N_1408,N_1781);
or U3510 (N_3510,N_1393,N_1032);
and U3511 (N_3511,N_889,N_953);
nor U3512 (N_3512,N_1530,N_19);
nor U3513 (N_3513,N_293,N_1556);
nand U3514 (N_3514,N_1301,N_83);
nor U3515 (N_3515,N_572,N_587);
and U3516 (N_3516,N_1639,N_994);
nand U3517 (N_3517,N_445,N_459);
nor U3518 (N_3518,N_839,N_1811);
nor U3519 (N_3519,N_21,N_930);
and U3520 (N_3520,N_1799,N_1232);
or U3521 (N_3521,N_739,N_421);
and U3522 (N_3522,N_1709,N_674);
nand U3523 (N_3523,N_962,N_114);
nor U3524 (N_3524,N_486,N_1583);
nor U3525 (N_3525,N_1957,N_961);
or U3526 (N_3526,N_147,N_150);
xnor U3527 (N_3527,N_1562,N_1595);
or U3528 (N_3528,N_1489,N_1641);
and U3529 (N_3529,N_1654,N_661);
nand U3530 (N_3530,N_1491,N_1805);
nand U3531 (N_3531,N_263,N_800);
and U3532 (N_3532,N_1674,N_1683);
nor U3533 (N_3533,N_663,N_209);
and U3534 (N_3534,N_55,N_665);
nor U3535 (N_3535,N_598,N_758);
or U3536 (N_3536,N_605,N_1694);
or U3537 (N_3537,N_217,N_289);
or U3538 (N_3538,N_182,N_1864);
xor U3539 (N_3539,N_1497,N_400);
or U3540 (N_3540,N_1556,N_1700);
and U3541 (N_3541,N_542,N_1098);
and U3542 (N_3542,N_1341,N_903);
nand U3543 (N_3543,N_1662,N_1092);
and U3544 (N_3544,N_1799,N_1189);
or U3545 (N_3545,N_66,N_498);
nand U3546 (N_3546,N_727,N_746);
xnor U3547 (N_3547,N_1255,N_1586);
nand U3548 (N_3548,N_456,N_1097);
or U3549 (N_3549,N_739,N_1347);
xnor U3550 (N_3550,N_84,N_1722);
nor U3551 (N_3551,N_206,N_384);
nor U3552 (N_3552,N_1146,N_756);
or U3553 (N_3553,N_1932,N_1480);
nor U3554 (N_3554,N_1715,N_1579);
and U3555 (N_3555,N_734,N_467);
nor U3556 (N_3556,N_254,N_444);
nor U3557 (N_3557,N_1811,N_45);
nor U3558 (N_3558,N_715,N_391);
nand U3559 (N_3559,N_1766,N_47);
or U3560 (N_3560,N_487,N_167);
nand U3561 (N_3561,N_851,N_1101);
nand U3562 (N_3562,N_297,N_649);
nand U3563 (N_3563,N_1351,N_1760);
nor U3564 (N_3564,N_266,N_666);
and U3565 (N_3565,N_1524,N_752);
nor U3566 (N_3566,N_644,N_350);
and U3567 (N_3567,N_1403,N_242);
nor U3568 (N_3568,N_697,N_1055);
and U3569 (N_3569,N_673,N_1213);
and U3570 (N_3570,N_1420,N_1553);
or U3571 (N_3571,N_227,N_235);
and U3572 (N_3572,N_1050,N_1469);
or U3573 (N_3573,N_1419,N_488);
xnor U3574 (N_3574,N_626,N_1010);
and U3575 (N_3575,N_306,N_1121);
nand U3576 (N_3576,N_1692,N_1181);
and U3577 (N_3577,N_379,N_1394);
xor U3578 (N_3578,N_1254,N_1000);
or U3579 (N_3579,N_780,N_1167);
xor U3580 (N_3580,N_1316,N_1855);
nand U3581 (N_3581,N_1885,N_423);
nor U3582 (N_3582,N_1001,N_692);
and U3583 (N_3583,N_1159,N_194);
or U3584 (N_3584,N_313,N_1067);
or U3585 (N_3585,N_195,N_1963);
nor U3586 (N_3586,N_1930,N_593);
nor U3587 (N_3587,N_1096,N_152);
and U3588 (N_3588,N_28,N_1874);
and U3589 (N_3589,N_968,N_1820);
nor U3590 (N_3590,N_447,N_632);
and U3591 (N_3591,N_1497,N_264);
nor U3592 (N_3592,N_1705,N_1071);
and U3593 (N_3593,N_1422,N_37);
or U3594 (N_3594,N_833,N_663);
nor U3595 (N_3595,N_175,N_1900);
nand U3596 (N_3596,N_223,N_160);
nand U3597 (N_3597,N_58,N_1424);
xnor U3598 (N_3598,N_765,N_1922);
nor U3599 (N_3599,N_293,N_1871);
and U3600 (N_3600,N_1185,N_752);
or U3601 (N_3601,N_63,N_138);
and U3602 (N_3602,N_420,N_1275);
xnor U3603 (N_3603,N_603,N_1146);
or U3604 (N_3604,N_710,N_681);
nor U3605 (N_3605,N_1751,N_1507);
nand U3606 (N_3606,N_1369,N_860);
or U3607 (N_3607,N_1780,N_806);
nor U3608 (N_3608,N_1594,N_588);
nand U3609 (N_3609,N_1111,N_715);
or U3610 (N_3610,N_199,N_6);
and U3611 (N_3611,N_203,N_1832);
nand U3612 (N_3612,N_822,N_1387);
nor U3613 (N_3613,N_1633,N_1134);
and U3614 (N_3614,N_65,N_1108);
nand U3615 (N_3615,N_1391,N_522);
or U3616 (N_3616,N_1952,N_130);
nand U3617 (N_3617,N_796,N_966);
or U3618 (N_3618,N_1512,N_1415);
and U3619 (N_3619,N_577,N_1960);
and U3620 (N_3620,N_1602,N_937);
xnor U3621 (N_3621,N_1198,N_131);
or U3622 (N_3622,N_1058,N_776);
nor U3623 (N_3623,N_1216,N_540);
nor U3624 (N_3624,N_180,N_1118);
nand U3625 (N_3625,N_522,N_828);
nand U3626 (N_3626,N_1505,N_336);
nor U3627 (N_3627,N_1424,N_963);
or U3628 (N_3628,N_739,N_495);
or U3629 (N_3629,N_713,N_1006);
xor U3630 (N_3630,N_1853,N_973);
and U3631 (N_3631,N_683,N_1438);
nand U3632 (N_3632,N_1389,N_352);
nor U3633 (N_3633,N_1424,N_1410);
or U3634 (N_3634,N_598,N_1981);
and U3635 (N_3635,N_690,N_1678);
or U3636 (N_3636,N_1151,N_704);
nand U3637 (N_3637,N_180,N_27);
or U3638 (N_3638,N_1455,N_496);
nand U3639 (N_3639,N_956,N_732);
xnor U3640 (N_3640,N_419,N_1023);
and U3641 (N_3641,N_1409,N_1949);
nand U3642 (N_3642,N_848,N_210);
or U3643 (N_3643,N_297,N_516);
and U3644 (N_3644,N_762,N_228);
nand U3645 (N_3645,N_1945,N_145);
nand U3646 (N_3646,N_151,N_1874);
nor U3647 (N_3647,N_968,N_1521);
and U3648 (N_3648,N_746,N_1530);
nand U3649 (N_3649,N_1959,N_861);
and U3650 (N_3650,N_760,N_1951);
and U3651 (N_3651,N_1441,N_36);
and U3652 (N_3652,N_1974,N_336);
nand U3653 (N_3653,N_352,N_1408);
xor U3654 (N_3654,N_1286,N_1429);
and U3655 (N_3655,N_601,N_1095);
and U3656 (N_3656,N_1684,N_1336);
or U3657 (N_3657,N_141,N_1612);
nand U3658 (N_3658,N_1031,N_1086);
and U3659 (N_3659,N_608,N_759);
nor U3660 (N_3660,N_539,N_1027);
nor U3661 (N_3661,N_1899,N_140);
nand U3662 (N_3662,N_773,N_1024);
and U3663 (N_3663,N_1084,N_1047);
xnor U3664 (N_3664,N_919,N_827);
and U3665 (N_3665,N_209,N_1157);
or U3666 (N_3666,N_1121,N_1470);
and U3667 (N_3667,N_1556,N_71);
and U3668 (N_3668,N_628,N_80);
nand U3669 (N_3669,N_613,N_270);
or U3670 (N_3670,N_383,N_970);
or U3671 (N_3671,N_432,N_1024);
nand U3672 (N_3672,N_1908,N_649);
xor U3673 (N_3673,N_142,N_82);
nand U3674 (N_3674,N_851,N_706);
or U3675 (N_3675,N_86,N_1966);
xor U3676 (N_3676,N_1649,N_920);
and U3677 (N_3677,N_931,N_640);
and U3678 (N_3678,N_557,N_1532);
and U3679 (N_3679,N_1649,N_1947);
xor U3680 (N_3680,N_1235,N_622);
nand U3681 (N_3681,N_608,N_1206);
nor U3682 (N_3682,N_368,N_1607);
or U3683 (N_3683,N_498,N_315);
xor U3684 (N_3684,N_1875,N_892);
or U3685 (N_3685,N_1593,N_1802);
nor U3686 (N_3686,N_1498,N_1998);
or U3687 (N_3687,N_1706,N_474);
or U3688 (N_3688,N_16,N_958);
or U3689 (N_3689,N_172,N_943);
nand U3690 (N_3690,N_1927,N_269);
nor U3691 (N_3691,N_1670,N_1960);
or U3692 (N_3692,N_791,N_1382);
and U3693 (N_3693,N_114,N_306);
or U3694 (N_3694,N_1806,N_1917);
or U3695 (N_3695,N_1221,N_1459);
and U3696 (N_3696,N_905,N_767);
nand U3697 (N_3697,N_349,N_551);
nor U3698 (N_3698,N_1767,N_1472);
nor U3699 (N_3699,N_1298,N_1891);
nor U3700 (N_3700,N_297,N_1649);
and U3701 (N_3701,N_1658,N_1939);
nand U3702 (N_3702,N_496,N_1);
and U3703 (N_3703,N_471,N_1098);
xnor U3704 (N_3704,N_800,N_620);
and U3705 (N_3705,N_790,N_557);
or U3706 (N_3706,N_185,N_1481);
nand U3707 (N_3707,N_971,N_421);
nor U3708 (N_3708,N_312,N_1347);
nand U3709 (N_3709,N_732,N_1924);
and U3710 (N_3710,N_118,N_1736);
and U3711 (N_3711,N_860,N_1101);
or U3712 (N_3712,N_1491,N_1998);
nand U3713 (N_3713,N_306,N_1004);
or U3714 (N_3714,N_1503,N_1705);
or U3715 (N_3715,N_1517,N_768);
and U3716 (N_3716,N_1923,N_1944);
and U3717 (N_3717,N_1242,N_1701);
nand U3718 (N_3718,N_1430,N_1611);
nand U3719 (N_3719,N_274,N_764);
nor U3720 (N_3720,N_1637,N_1577);
nor U3721 (N_3721,N_765,N_1135);
or U3722 (N_3722,N_1712,N_1640);
or U3723 (N_3723,N_1691,N_1560);
nor U3724 (N_3724,N_615,N_92);
nand U3725 (N_3725,N_893,N_11);
or U3726 (N_3726,N_1073,N_1052);
nor U3727 (N_3727,N_250,N_1802);
or U3728 (N_3728,N_1817,N_1856);
or U3729 (N_3729,N_1653,N_152);
and U3730 (N_3730,N_1160,N_1812);
and U3731 (N_3731,N_1502,N_746);
nand U3732 (N_3732,N_725,N_1039);
and U3733 (N_3733,N_1371,N_882);
nor U3734 (N_3734,N_741,N_1153);
nand U3735 (N_3735,N_264,N_231);
nor U3736 (N_3736,N_1126,N_1676);
or U3737 (N_3737,N_1032,N_1834);
nor U3738 (N_3738,N_1472,N_1845);
or U3739 (N_3739,N_1340,N_1953);
and U3740 (N_3740,N_1773,N_302);
xor U3741 (N_3741,N_400,N_265);
or U3742 (N_3742,N_1014,N_1015);
nand U3743 (N_3743,N_897,N_348);
and U3744 (N_3744,N_840,N_1562);
or U3745 (N_3745,N_1000,N_579);
and U3746 (N_3746,N_895,N_328);
nand U3747 (N_3747,N_1286,N_1257);
or U3748 (N_3748,N_445,N_1578);
or U3749 (N_3749,N_290,N_577);
nand U3750 (N_3750,N_543,N_554);
and U3751 (N_3751,N_957,N_1400);
nor U3752 (N_3752,N_148,N_1061);
xnor U3753 (N_3753,N_127,N_1183);
and U3754 (N_3754,N_1448,N_253);
or U3755 (N_3755,N_1,N_630);
nor U3756 (N_3756,N_817,N_1721);
nand U3757 (N_3757,N_1728,N_1451);
or U3758 (N_3758,N_1571,N_1084);
nor U3759 (N_3759,N_1013,N_1964);
or U3760 (N_3760,N_1906,N_1313);
and U3761 (N_3761,N_1280,N_886);
and U3762 (N_3762,N_441,N_1329);
nand U3763 (N_3763,N_867,N_267);
or U3764 (N_3764,N_1565,N_1721);
or U3765 (N_3765,N_1148,N_1794);
xor U3766 (N_3766,N_335,N_1368);
or U3767 (N_3767,N_349,N_1168);
or U3768 (N_3768,N_41,N_189);
nor U3769 (N_3769,N_1538,N_1068);
nand U3770 (N_3770,N_71,N_974);
nor U3771 (N_3771,N_1183,N_652);
nand U3772 (N_3772,N_174,N_1947);
and U3773 (N_3773,N_473,N_1177);
and U3774 (N_3774,N_754,N_636);
nor U3775 (N_3775,N_1695,N_560);
nor U3776 (N_3776,N_1522,N_1483);
nor U3777 (N_3777,N_441,N_1586);
nand U3778 (N_3778,N_1541,N_1565);
nor U3779 (N_3779,N_943,N_1144);
or U3780 (N_3780,N_1145,N_1283);
or U3781 (N_3781,N_1719,N_590);
nor U3782 (N_3782,N_1465,N_883);
nor U3783 (N_3783,N_1030,N_807);
or U3784 (N_3784,N_730,N_438);
or U3785 (N_3785,N_750,N_866);
or U3786 (N_3786,N_1585,N_499);
nand U3787 (N_3787,N_1031,N_1622);
nand U3788 (N_3788,N_1757,N_2);
xnor U3789 (N_3789,N_756,N_1223);
nand U3790 (N_3790,N_1550,N_1640);
xor U3791 (N_3791,N_409,N_662);
and U3792 (N_3792,N_974,N_941);
and U3793 (N_3793,N_1929,N_291);
or U3794 (N_3794,N_222,N_352);
nor U3795 (N_3795,N_531,N_57);
nand U3796 (N_3796,N_1688,N_427);
nand U3797 (N_3797,N_611,N_680);
and U3798 (N_3798,N_713,N_1838);
nor U3799 (N_3799,N_1150,N_1059);
nor U3800 (N_3800,N_1783,N_1165);
nor U3801 (N_3801,N_639,N_300);
nor U3802 (N_3802,N_5,N_1223);
xnor U3803 (N_3803,N_403,N_726);
nand U3804 (N_3804,N_750,N_120);
and U3805 (N_3805,N_135,N_1316);
and U3806 (N_3806,N_546,N_1032);
or U3807 (N_3807,N_1364,N_1774);
or U3808 (N_3808,N_258,N_766);
nor U3809 (N_3809,N_484,N_1003);
nor U3810 (N_3810,N_100,N_678);
or U3811 (N_3811,N_1215,N_932);
nor U3812 (N_3812,N_1200,N_1294);
nand U3813 (N_3813,N_827,N_718);
and U3814 (N_3814,N_1534,N_91);
or U3815 (N_3815,N_855,N_592);
nand U3816 (N_3816,N_1903,N_487);
nor U3817 (N_3817,N_479,N_673);
nand U3818 (N_3818,N_1705,N_971);
nor U3819 (N_3819,N_640,N_243);
or U3820 (N_3820,N_1745,N_1224);
nand U3821 (N_3821,N_419,N_1848);
or U3822 (N_3822,N_28,N_1709);
or U3823 (N_3823,N_566,N_386);
nand U3824 (N_3824,N_705,N_1945);
and U3825 (N_3825,N_909,N_1771);
and U3826 (N_3826,N_42,N_1253);
nor U3827 (N_3827,N_1209,N_1352);
and U3828 (N_3828,N_1471,N_1303);
or U3829 (N_3829,N_1901,N_40);
or U3830 (N_3830,N_559,N_287);
xnor U3831 (N_3831,N_1790,N_885);
nand U3832 (N_3832,N_285,N_1107);
nor U3833 (N_3833,N_5,N_662);
or U3834 (N_3834,N_40,N_15);
nand U3835 (N_3835,N_1369,N_543);
and U3836 (N_3836,N_1946,N_59);
nor U3837 (N_3837,N_1005,N_508);
nand U3838 (N_3838,N_418,N_924);
nand U3839 (N_3839,N_1077,N_181);
nand U3840 (N_3840,N_1704,N_1875);
or U3841 (N_3841,N_877,N_169);
nor U3842 (N_3842,N_290,N_1987);
xor U3843 (N_3843,N_1871,N_1651);
or U3844 (N_3844,N_1582,N_1212);
and U3845 (N_3845,N_553,N_193);
nand U3846 (N_3846,N_1217,N_920);
and U3847 (N_3847,N_644,N_1830);
or U3848 (N_3848,N_825,N_1254);
xnor U3849 (N_3849,N_1043,N_477);
or U3850 (N_3850,N_1159,N_1209);
or U3851 (N_3851,N_270,N_457);
nand U3852 (N_3852,N_327,N_44);
nor U3853 (N_3853,N_1974,N_708);
nand U3854 (N_3854,N_1813,N_334);
or U3855 (N_3855,N_1497,N_1588);
or U3856 (N_3856,N_789,N_1568);
or U3857 (N_3857,N_875,N_393);
or U3858 (N_3858,N_720,N_1153);
nor U3859 (N_3859,N_401,N_1531);
xor U3860 (N_3860,N_1492,N_300);
xor U3861 (N_3861,N_998,N_394);
nand U3862 (N_3862,N_1205,N_697);
and U3863 (N_3863,N_1754,N_198);
nor U3864 (N_3864,N_1267,N_191);
nand U3865 (N_3865,N_1939,N_1979);
and U3866 (N_3866,N_428,N_1351);
xnor U3867 (N_3867,N_1369,N_1565);
or U3868 (N_3868,N_565,N_1563);
and U3869 (N_3869,N_1647,N_1515);
nand U3870 (N_3870,N_1656,N_760);
or U3871 (N_3871,N_1602,N_1004);
and U3872 (N_3872,N_1193,N_1227);
nand U3873 (N_3873,N_1732,N_1002);
and U3874 (N_3874,N_992,N_664);
nand U3875 (N_3875,N_1967,N_1558);
and U3876 (N_3876,N_236,N_1020);
and U3877 (N_3877,N_903,N_1879);
and U3878 (N_3878,N_1985,N_1844);
or U3879 (N_3879,N_1284,N_395);
nand U3880 (N_3880,N_1610,N_765);
nor U3881 (N_3881,N_818,N_110);
nor U3882 (N_3882,N_1703,N_969);
or U3883 (N_3883,N_1365,N_1263);
nor U3884 (N_3884,N_993,N_363);
or U3885 (N_3885,N_923,N_1796);
nor U3886 (N_3886,N_1466,N_1664);
nor U3887 (N_3887,N_970,N_787);
nor U3888 (N_3888,N_376,N_635);
and U3889 (N_3889,N_637,N_1984);
and U3890 (N_3890,N_784,N_95);
nand U3891 (N_3891,N_1513,N_1266);
xor U3892 (N_3892,N_1650,N_1472);
nor U3893 (N_3893,N_521,N_1934);
nand U3894 (N_3894,N_362,N_535);
nand U3895 (N_3895,N_766,N_449);
nand U3896 (N_3896,N_887,N_234);
and U3897 (N_3897,N_1547,N_671);
and U3898 (N_3898,N_1132,N_594);
nor U3899 (N_3899,N_556,N_496);
xor U3900 (N_3900,N_1390,N_658);
nand U3901 (N_3901,N_930,N_1666);
and U3902 (N_3902,N_606,N_895);
nand U3903 (N_3903,N_1923,N_948);
nor U3904 (N_3904,N_278,N_1297);
and U3905 (N_3905,N_812,N_82);
nor U3906 (N_3906,N_1608,N_494);
xnor U3907 (N_3907,N_701,N_1253);
nand U3908 (N_3908,N_617,N_1401);
nor U3909 (N_3909,N_1279,N_1513);
nor U3910 (N_3910,N_1282,N_448);
and U3911 (N_3911,N_1129,N_660);
and U3912 (N_3912,N_1243,N_656);
nand U3913 (N_3913,N_1805,N_622);
xor U3914 (N_3914,N_107,N_1714);
or U3915 (N_3915,N_1036,N_1929);
xor U3916 (N_3916,N_1527,N_1063);
or U3917 (N_3917,N_530,N_766);
nand U3918 (N_3918,N_1750,N_1265);
nand U3919 (N_3919,N_1186,N_412);
and U3920 (N_3920,N_223,N_410);
nor U3921 (N_3921,N_1864,N_567);
xnor U3922 (N_3922,N_1532,N_216);
or U3923 (N_3923,N_269,N_255);
nor U3924 (N_3924,N_1394,N_451);
or U3925 (N_3925,N_1886,N_455);
xnor U3926 (N_3926,N_1251,N_976);
xor U3927 (N_3927,N_252,N_289);
nand U3928 (N_3928,N_30,N_1206);
and U3929 (N_3929,N_945,N_505);
nand U3930 (N_3930,N_1214,N_837);
xor U3931 (N_3931,N_846,N_1170);
nand U3932 (N_3932,N_496,N_701);
nand U3933 (N_3933,N_316,N_1874);
xor U3934 (N_3934,N_1278,N_1131);
xnor U3935 (N_3935,N_590,N_1798);
or U3936 (N_3936,N_1263,N_1259);
or U3937 (N_3937,N_1997,N_731);
and U3938 (N_3938,N_1392,N_1449);
and U3939 (N_3939,N_1247,N_645);
xnor U3940 (N_3940,N_1083,N_1121);
xor U3941 (N_3941,N_1069,N_1274);
xor U3942 (N_3942,N_324,N_469);
and U3943 (N_3943,N_915,N_0);
or U3944 (N_3944,N_323,N_177);
or U3945 (N_3945,N_27,N_936);
and U3946 (N_3946,N_1453,N_1912);
or U3947 (N_3947,N_1529,N_1860);
nand U3948 (N_3948,N_284,N_863);
nand U3949 (N_3949,N_1356,N_1050);
nand U3950 (N_3950,N_814,N_791);
nand U3951 (N_3951,N_1080,N_1875);
or U3952 (N_3952,N_1662,N_377);
nor U3953 (N_3953,N_1362,N_40);
and U3954 (N_3954,N_1852,N_1254);
nand U3955 (N_3955,N_23,N_574);
xnor U3956 (N_3956,N_6,N_91);
xor U3957 (N_3957,N_643,N_755);
and U3958 (N_3958,N_704,N_1209);
or U3959 (N_3959,N_665,N_255);
and U3960 (N_3960,N_504,N_251);
nor U3961 (N_3961,N_377,N_1858);
or U3962 (N_3962,N_486,N_30);
or U3963 (N_3963,N_578,N_1856);
and U3964 (N_3964,N_208,N_519);
nand U3965 (N_3965,N_1507,N_798);
xnor U3966 (N_3966,N_823,N_708);
nor U3967 (N_3967,N_438,N_306);
nand U3968 (N_3968,N_66,N_212);
and U3969 (N_3969,N_126,N_1581);
and U3970 (N_3970,N_1931,N_906);
and U3971 (N_3971,N_1489,N_62);
or U3972 (N_3972,N_783,N_1863);
nand U3973 (N_3973,N_152,N_679);
nor U3974 (N_3974,N_1815,N_171);
or U3975 (N_3975,N_1556,N_183);
nand U3976 (N_3976,N_1025,N_1357);
or U3977 (N_3977,N_1517,N_1356);
nand U3978 (N_3978,N_1108,N_1151);
nand U3979 (N_3979,N_1452,N_526);
or U3980 (N_3980,N_1486,N_576);
and U3981 (N_3981,N_1759,N_732);
nor U3982 (N_3982,N_1510,N_642);
or U3983 (N_3983,N_770,N_1429);
and U3984 (N_3984,N_825,N_91);
and U3985 (N_3985,N_67,N_95);
xor U3986 (N_3986,N_1665,N_1374);
nand U3987 (N_3987,N_1236,N_677);
nand U3988 (N_3988,N_1019,N_236);
and U3989 (N_3989,N_852,N_1233);
or U3990 (N_3990,N_91,N_558);
nor U3991 (N_3991,N_1339,N_1081);
nand U3992 (N_3992,N_977,N_1495);
nor U3993 (N_3993,N_756,N_1215);
xnor U3994 (N_3994,N_1680,N_1562);
nor U3995 (N_3995,N_1400,N_1188);
nand U3996 (N_3996,N_1204,N_1763);
nor U3997 (N_3997,N_755,N_1139);
or U3998 (N_3998,N_1624,N_546);
or U3999 (N_3999,N_912,N_1911);
or U4000 (N_4000,N_2578,N_2825);
nand U4001 (N_4001,N_2741,N_3855);
or U4002 (N_4002,N_2414,N_2826);
and U4003 (N_4003,N_2447,N_2655);
or U4004 (N_4004,N_3922,N_3055);
nand U4005 (N_4005,N_2165,N_3865);
nand U4006 (N_4006,N_2601,N_3021);
or U4007 (N_4007,N_2040,N_2900);
xor U4008 (N_4008,N_3116,N_3435);
nand U4009 (N_4009,N_3837,N_3051);
xor U4010 (N_4010,N_2435,N_2445);
nand U4011 (N_4011,N_3065,N_2292);
or U4012 (N_4012,N_3285,N_3164);
nor U4013 (N_4013,N_2373,N_2336);
or U4014 (N_4014,N_2609,N_3247);
nor U4015 (N_4015,N_3686,N_3890);
and U4016 (N_4016,N_3458,N_3776);
nor U4017 (N_4017,N_3591,N_3223);
or U4018 (N_4018,N_3919,N_3942);
and U4019 (N_4019,N_3347,N_2961);
nor U4020 (N_4020,N_2914,N_3460);
nor U4021 (N_4021,N_3887,N_3044);
nor U4022 (N_4022,N_2619,N_2369);
and U4023 (N_4023,N_3530,N_3235);
nor U4024 (N_4024,N_3396,N_3770);
or U4025 (N_4025,N_2988,N_3599);
or U4026 (N_4026,N_3367,N_2598);
and U4027 (N_4027,N_3420,N_2288);
nand U4028 (N_4028,N_3277,N_2028);
nor U4029 (N_4029,N_3513,N_3613);
nor U4030 (N_4030,N_3796,N_2811);
or U4031 (N_4031,N_3238,N_2696);
and U4032 (N_4032,N_3624,N_2842);
or U4033 (N_4033,N_2047,N_3709);
nor U4034 (N_4034,N_2658,N_3846);
nor U4035 (N_4035,N_2958,N_3201);
or U4036 (N_4036,N_2936,N_3958);
xnor U4037 (N_4037,N_2925,N_3813);
and U4038 (N_4038,N_2260,N_3150);
nor U4039 (N_4039,N_2903,N_2691);
and U4040 (N_4040,N_3313,N_3804);
nand U4041 (N_4041,N_2909,N_2636);
nor U4042 (N_4042,N_3035,N_2289);
and U4043 (N_4043,N_3782,N_2401);
nand U4044 (N_4044,N_2162,N_3068);
or U4045 (N_4045,N_3619,N_2891);
and U4046 (N_4046,N_2890,N_3830);
nand U4047 (N_4047,N_3622,N_2230);
nand U4048 (N_4048,N_3618,N_3973);
nor U4049 (N_4049,N_3444,N_2623);
or U4050 (N_4050,N_3412,N_2948);
and U4051 (N_4051,N_3766,N_2795);
and U4052 (N_4052,N_3082,N_3853);
xnor U4053 (N_4053,N_2234,N_2018);
nor U4054 (N_4054,N_2740,N_3754);
xor U4055 (N_4055,N_3646,N_3414);
xor U4056 (N_4056,N_3243,N_3240);
nand U4057 (N_4057,N_2546,N_3097);
nand U4058 (N_4058,N_2526,N_2202);
xnor U4059 (N_4059,N_2736,N_2629);
xor U4060 (N_4060,N_3215,N_3042);
and U4061 (N_4061,N_3126,N_2938);
nand U4062 (N_4062,N_3557,N_3436);
nor U4063 (N_4063,N_3349,N_2261);
nor U4064 (N_4064,N_2307,N_2461);
and U4065 (N_4065,N_3468,N_3857);
nor U4066 (N_4066,N_3230,N_3724);
nor U4067 (N_4067,N_3951,N_2644);
nand U4068 (N_4068,N_2072,N_2487);
or U4069 (N_4069,N_3262,N_2415);
or U4070 (N_4070,N_3812,N_2413);
and U4071 (N_4071,N_3673,N_3476);
or U4072 (N_4072,N_2228,N_2284);
or U4073 (N_4073,N_2592,N_3045);
or U4074 (N_4074,N_2215,N_3652);
and U4075 (N_4075,N_2033,N_3621);
nor U4076 (N_4076,N_2384,N_3779);
and U4077 (N_4077,N_2160,N_3514);
or U4078 (N_4078,N_2127,N_3493);
xnor U4079 (N_4079,N_2013,N_2743);
and U4080 (N_4080,N_2268,N_2400);
and U4081 (N_4081,N_3840,N_2888);
nor U4082 (N_4082,N_3981,N_3090);
nor U4083 (N_4083,N_2638,N_3699);
and U4084 (N_4084,N_2597,N_3250);
nor U4085 (N_4085,N_2978,N_3029);
nor U4086 (N_4086,N_3986,N_2507);
and U4087 (N_4087,N_3936,N_3140);
nand U4088 (N_4088,N_2784,N_2171);
nor U4089 (N_4089,N_2320,N_3426);
nor U4090 (N_4090,N_3397,N_2761);
or U4091 (N_4091,N_3688,N_3715);
xnor U4092 (N_4092,N_2466,N_2739);
and U4093 (N_4093,N_3935,N_3982);
nor U4094 (N_4094,N_3987,N_2087);
nand U4095 (N_4095,N_3685,N_2392);
and U4096 (N_4096,N_3604,N_3502);
or U4097 (N_4097,N_3665,N_3927);
nor U4098 (N_4098,N_2079,N_3010);
or U4099 (N_4099,N_3077,N_2590);
or U4100 (N_4100,N_3096,N_2068);
nor U4101 (N_4101,N_3969,N_2679);
nand U4102 (N_4102,N_3542,N_3428);
nor U4103 (N_4103,N_3245,N_3020);
nor U4104 (N_4104,N_3115,N_3399);
nand U4105 (N_4105,N_3635,N_2050);
nor U4106 (N_4106,N_2015,N_3907);
or U4107 (N_4107,N_3898,N_2627);
or U4108 (N_4108,N_3566,N_3667);
nor U4109 (N_4109,N_3564,N_3968);
and U4110 (N_4110,N_2799,N_2570);
nor U4111 (N_4111,N_2243,N_2659);
xnor U4112 (N_4112,N_3264,N_3036);
or U4113 (N_4113,N_2272,N_2731);
nand U4114 (N_4114,N_3048,N_3595);
nand U4115 (N_4115,N_2448,N_2910);
and U4116 (N_4116,N_2820,N_3291);
and U4117 (N_4117,N_3382,N_3616);
nor U4118 (N_4118,N_2553,N_3679);
and U4119 (N_4119,N_3216,N_3344);
and U4120 (N_4120,N_2967,N_2617);
nor U4121 (N_4121,N_2934,N_3944);
nand U4122 (N_4122,N_2966,N_3343);
and U4123 (N_4123,N_2287,N_2429);
nand U4124 (N_4124,N_2531,N_3778);
nand U4125 (N_4125,N_3177,N_3429);
nor U4126 (N_4126,N_3901,N_2084);
nand U4127 (N_4127,N_2703,N_3902);
nand U4128 (N_4128,N_3132,N_3369);
xnor U4129 (N_4129,N_3455,N_2879);
or U4130 (N_4130,N_2264,N_3141);
nor U4131 (N_4131,N_2338,N_3500);
xnor U4132 (N_4132,N_2575,N_3854);
nor U4133 (N_4133,N_3790,N_3729);
and U4134 (N_4134,N_2712,N_2439);
and U4135 (N_4135,N_2863,N_3976);
xor U4136 (N_4136,N_2587,N_3886);
and U4137 (N_4137,N_3047,N_2633);
or U4138 (N_4138,N_3832,N_2115);
nand U4139 (N_4139,N_3009,N_2962);
nor U4140 (N_4140,N_3208,N_2303);
and U4141 (N_4141,N_2545,N_3324);
nor U4142 (N_4142,N_3188,N_2042);
and U4143 (N_4143,N_2662,N_2204);
nand U4144 (N_4144,N_3627,N_2785);
nor U4145 (N_4145,N_3228,N_3341);
or U4146 (N_4146,N_2455,N_3548);
nor U4147 (N_4147,N_2019,N_3966);
or U4148 (N_4148,N_3878,N_2045);
and U4149 (N_4149,N_3822,N_3231);
or U4150 (N_4150,N_2122,N_3008);
or U4151 (N_4151,N_2669,N_2552);
or U4152 (N_4152,N_3841,N_3317);
nor U4153 (N_4153,N_3254,N_2744);
or U4154 (N_4154,N_3301,N_2494);
xor U4155 (N_4155,N_2219,N_2245);
nor U4156 (N_4156,N_2498,N_2959);
and U4157 (N_4157,N_3915,N_2342);
nand U4158 (N_4158,N_2821,N_2156);
and U4159 (N_4159,N_3427,N_3520);
or U4160 (N_4160,N_2408,N_2027);
nand U4161 (N_4161,N_3824,N_2346);
or U4162 (N_4162,N_2975,N_3979);
or U4163 (N_4163,N_3167,N_2536);
nor U4164 (N_4164,N_2725,N_2880);
or U4165 (N_4165,N_2972,N_3834);
and U4166 (N_4166,N_3598,N_2329);
xor U4167 (N_4167,N_3783,N_3847);
or U4168 (N_4168,N_2104,N_3883);
xor U4169 (N_4169,N_2341,N_3615);
nand U4170 (N_4170,N_3517,N_3753);
xnor U4171 (N_4171,N_3198,N_3539);
xnor U4172 (N_4172,N_3536,N_2901);
nor U4173 (N_4173,N_3109,N_3743);
xnor U4174 (N_4174,N_2049,N_3028);
nand U4175 (N_4175,N_3448,N_2174);
nor U4176 (N_4176,N_3328,N_2090);
nand U4177 (N_4177,N_2647,N_2167);
xnor U4178 (N_4178,N_2358,N_3971);
and U4179 (N_4179,N_3316,N_2912);
nand U4180 (N_4180,N_2273,N_3512);
nor U4181 (N_4181,N_3144,N_3255);
and U4182 (N_4182,N_2310,N_2995);
and U4183 (N_4183,N_2332,N_3123);
nand U4184 (N_4184,N_2351,N_2857);
nor U4185 (N_4185,N_2130,N_2702);
and U4186 (N_4186,N_3510,N_2618);
nand U4187 (N_4187,N_3292,N_2709);
nand U4188 (N_4188,N_2353,N_3532);
and U4189 (N_4189,N_3092,N_2349);
nand U4190 (N_4190,N_3166,N_2881);
nor U4191 (N_4191,N_3803,N_2294);
or U4192 (N_4192,N_3389,N_2304);
or U4193 (N_4193,N_2678,N_2684);
or U4194 (N_4194,N_2100,N_2947);
nor U4195 (N_4195,N_2152,N_2670);
xor U4196 (N_4196,N_3746,N_3997);
and U4197 (N_4197,N_2957,N_3212);
or U4198 (N_4198,N_2168,N_2993);
nor U4199 (N_4199,N_3845,N_3637);
and U4200 (N_4200,N_3148,N_2613);
nor U4201 (N_4201,N_2089,N_2527);
nor U4202 (N_4202,N_2252,N_2453);
or U4203 (N_4203,N_2490,N_3495);
nand U4204 (N_4204,N_3903,N_2665);
nand U4205 (N_4205,N_3693,N_2161);
and U4206 (N_4206,N_2181,N_2577);
nor U4207 (N_4207,N_2897,N_2950);
and U4208 (N_4208,N_2768,N_3664);
nor U4209 (N_4209,N_3678,N_3360);
nor U4210 (N_4210,N_2144,N_2055);
nand U4211 (N_4211,N_3340,N_3385);
and U4212 (N_4212,N_3617,N_2225);
and U4213 (N_4213,N_2295,N_2123);
xnor U4214 (N_4214,N_2532,N_2321);
nand U4215 (N_4215,N_2265,N_2838);
nand U4216 (N_4216,N_2782,N_3070);
nor U4217 (N_4217,N_3653,N_2191);
and U4218 (N_4218,N_3300,N_2639);
nor U4219 (N_4219,N_3704,N_3759);
and U4220 (N_4220,N_3511,N_3183);
nand U4221 (N_4221,N_3073,N_3118);
or U4222 (N_4222,N_2694,N_3642);
nor U4223 (N_4223,N_2675,N_2073);
or U4224 (N_4224,N_3383,N_2126);
nor U4225 (N_4225,N_2356,N_3603);
nand U4226 (N_4226,N_3309,N_2529);
and U4227 (N_4227,N_2212,N_3763);
or U4228 (N_4228,N_3745,N_3459);
and U4229 (N_4229,N_2423,N_2023);
xnor U4230 (N_4230,N_2990,N_3153);
nor U4231 (N_4231,N_2020,N_2125);
nor U4232 (N_4232,N_2078,N_3839);
nand U4233 (N_4233,N_2076,N_2685);
and U4234 (N_4234,N_3287,N_2451);
and U4235 (N_4235,N_3716,N_2555);
or U4236 (N_4236,N_2110,N_3134);
and U4237 (N_4237,N_2119,N_3333);
and U4238 (N_4238,N_3998,N_3643);
nand U4239 (N_4239,N_3992,N_3308);
and U4240 (N_4240,N_3259,N_2322);
nor U4241 (N_4241,N_3422,N_2190);
and U4242 (N_4242,N_2333,N_2386);
nor U4243 (N_4243,N_3527,N_3221);
nand U4244 (N_4244,N_2483,N_2108);
nand U4245 (N_4245,N_3952,N_2954);
and U4246 (N_4246,N_3103,N_2008);
nor U4247 (N_4247,N_2989,N_3283);
nor U4248 (N_4248,N_3000,N_3737);
or U4249 (N_4249,N_3424,N_2229);
or U4250 (N_4250,N_3991,N_3807);
xnor U4251 (N_4251,N_3970,N_2921);
and U4252 (N_4252,N_2754,N_2029);
xor U4253 (N_4253,N_2381,N_2688);
and U4254 (N_4254,N_2985,N_3735);
nand U4255 (N_4255,N_2753,N_2773);
or U4256 (N_4256,N_2098,N_2390);
and U4257 (N_4257,N_3191,N_3127);
nor U4258 (N_4258,N_2614,N_3974);
or U4259 (N_4259,N_3411,N_3761);
nor U4260 (N_4260,N_2025,N_3496);
nor U4261 (N_4261,N_2470,N_2977);
or U4262 (N_4262,N_2622,N_2365);
or U4263 (N_4263,N_3381,N_2118);
nor U4264 (N_4264,N_2205,N_3798);
or U4265 (N_4265,N_3559,N_3634);
nor U4266 (N_4266,N_3636,N_3911);
and U4267 (N_4267,N_3727,N_2651);
or U4268 (N_4268,N_3178,N_2733);
nor U4269 (N_4269,N_3039,N_2635);
or U4270 (N_4270,N_2893,N_3101);
xor U4271 (N_4271,N_2139,N_2851);
nor U4272 (N_4272,N_3180,N_2195);
or U4273 (N_4273,N_3355,N_2766);
and U4274 (N_4274,N_2363,N_2861);
or U4275 (N_4275,N_2145,N_3639);
or U4276 (N_4276,N_3815,N_2819);
xnor U4277 (N_4277,N_3346,N_3592);
and U4278 (N_4278,N_3863,N_3996);
xor U4279 (N_4279,N_3366,N_2790);
nand U4280 (N_4280,N_3083,N_2812);
and U4281 (N_4281,N_3787,N_2537);
nand U4282 (N_4282,N_3279,N_2048);
nor U4283 (N_4283,N_2833,N_2681);
nand U4284 (N_4284,N_2634,N_2091);
nor U4285 (N_4285,N_2796,N_3268);
nor U4286 (N_4286,N_2308,N_3326);
and U4287 (N_4287,N_2482,N_3239);
nor U4288 (N_4288,N_3645,N_3494);
nor U4289 (N_4289,N_3711,N_2297);
nand U4290 (N_4290,N_2339,N_3195);
or U4291 (N_4291,N_2412,N_3905);
and U4292 (N_4292,N_3474,N_3151);
and U4293 (N_4293,N_3288,N_2603);
nor U4294 (N_4294,N_2596,N_3297);
xnor U4295 (N_4295,N_3370,N_3146);
nand U4296 (N_4296,N_3380,N_3362);
and U4297 (N_4297,N_2132,N_2282);
or U4298 (N_4298,N_2649,N_3608);
xnor U4299 (N_4299,N_2194,N_2965);
nor U4300 (N_4300,N_2615,N_2937);
or U4301 (N_4301,N_3274,N_3576);
nand U4302 (N_4302,N_2374,N_3567);
and U4303 (N_4303,N_3315,N_3858);
or U4304 (N_4304,N_2846,N_2830);
and U4305 (N_4305,N_3242,N_3960);
nor U4306 (N_4306,N_3491,N_2530);
xnor U4307 (N_4307,N_2767,N_2660);
or U4308 (N_4308,N_3554,N_3695);
or U4309 (N_4309,N_3137,N_3058);
nand U4310 (N_4310,N_2422,N_2301);
or U4311 (N_4311,N_2565,N_2113);
nor U4312 (N_4312,N_3540,N_2533);
and U4313 (N_4313,N_2514,N_3323);
nor U4314 (N_4314,N_3069,N_3352);
and U4315 (N_4315,N_2722,N_3924);
or U4316 (N_4316,N_2915,N_2579);
nand U4317 (N_4317,N_3589,N_2683);
and U4318 (N_4318,N_3012,N_2387);
xnor U4319 (N_4319,N_2668,N_3278);
nand U4320 (N_4320,N_3676,N_3625);
xnor U4321 (N_4321,N_3738,N_2066);
nand U4322 (N_4322,N_3657,N_2855);
and U4323 (N_4323,N_3108,N_3296);
and U4324 (N_4324,N_3168,N_3914);
or U4325 (N_4325,N_3220,N_3670);
and U4326 (N_4326,N_3516,N_3789);
or U4327 (N_4327,N_2293,N_3106);
or U4328 (N_4328,N_2153,N_3139);
nand U4329 (N_4329,N_2562,N_2518);
or U4330 (N_4330,N_2437,N_2411);
xor U4331 (N_4331,N_2862,N_2460);
and U4332 (N_4332,N_2463,N_2805);
nand U4333 (N_4333,N_3049,N_2330);
and U4334 (N_4334,N_2941,N_3294);
and U4335 (N_4335,N_2515,N_2699);
nand U4336 (N_4336,N_2366,N_2757);
nand U4337 (N_4337,N_2886,N_2142);
xnor U4338 (N_4338,N_3063,N_3701);
nor U4339 (N_4339,N_3571,N_3361);
nor U4340 (N_4340,N_2426,N_2124);
or U4341 (N_4341,N_3913,N_3056);
nor U4342 (N_4342,N_3303,N_3094);
nand U4343 (N_4343,N_2640,N_2462);
or U4344 (N_4344,N_2086,N_3187);
or U4345 (N_4345,N_2478,N_2468);
nor U4346 (N_4346,N_3176,N_2102);
or U4347 (N_4347,N_3888,N_3172);
or U4348 (N_4348,N_3024,N_3365);
or U4349 (N_4349,N_3433,N_3462);
nor U4350 (N_4350,N_3655,N_2041);
or U4351 (N_4351,N_3658,N_2186);
or U4352 (N_4352,N_3454,N_3764);
or U4353 (N_4353,N_3192,N_2255);
nand U4354 (N_4354,N_2452,N_3479);
nor U4355 (N_4355,N_3722,N_3876);
nor U4356 (N_4356,N_2652,N_2641);
or U4357 (N_4357,N_2802,N_2714);
nor U4358 (N_4358,N_3980,N_2700);
or U4359 (N_4359,N_2238,N_2380);
nor U4360 (N_4360,N_2208,N_2899);
and U4361 (N_4361,N_3675,N_3747);
or U4362 (N_4362,N_2602,N_3408);
xnor U4363 (N_4363,N_3121,N_3504);
nand U4364 (N_4364,N_3768,N_3773);
nor U4365 (N_4365,N_3572,N_2378);
nor U4366 (N_4366,N_2198,N_3733);
nand U4367 (N_4367,N_3648,N_3896);
or U4368 (N_4368,N_3125,N_2864);
and U4369 (N_4369,N_2200,N_3415);
and U4370 (N_4370,N_2556,N_3486);
and U4371 (N_4371,N_2667,N_2038);
nand U4372 (N_4372,N_3842,N_2892);
xnor U4373 (N_4373,N_3714,N_3224);
nand U4374 (N_4374,N_3080,N_2749);
or U4375 (N_4375,N_2189,N_3473);
or U4376 (N_4376,N_2420,N_2718);
nor U4377 (N_4377,N_2464,N_3384);
and U4378 (N_4378,N_3629,N_3260);
nand U4379 (N_4379,N_2882,N_3152);
or U4380 (N_4380,N_3295,N_3989);
nor U4381 (N_4381,N_2564,N_3821);
nor U4382 (N_4382,N_3407,N_2248);
xnor U4383 (N_4383,N_3614,N_3644);
xor U4384 (N_4384,N_2371,N_2403);
and U4385 (N_4385,N_2956,N_3314);
nand U4386 (N_4386,N_3793,N_3207);
nand U4387 (N_4387,N_3921,N_2410);
or U4388 (N_4388,N_2509,N_2516);
nor U4389 (N_4389,N_3769,N_2164);
and U4390 (N_4390,N_2585,N_3043);
or U4391 (N_4391,N_3529,N_3034);
xnor U4392 (N_4392,N_3641,N_2017);
xnor U4393 (N_4393,N_2246,N_2711);
nand U4394 (N_4394,N_3609,N_3920);
nor U4395 (N_4395,N_3957,N_2524);
nor U4396 (N_4396,N_2479,N_3013);
and U4397 (N_4397,N_3556,N_3871);
and U4398 (N_4398,N_3794,N_2362);
and U4399 (N_4399,N_2535,N_3961);
nand U4400 (N_4400,N_2822,N_3792);
or U4401 (N_4401,N_3222,N_3165);
or U4402 (N_4402,N_3498,N_2600);
or U4403 (N_4403,N_3662,N_3910);
and U4404 (N_4404,N_3431,N_2783);
nor U4405 (N_4405,N_3033,N_3075);
nor U4406 (N_4406,N_3777,N_2044);
nand U4407 (N_4407,N_3702,N_3395);
nand U4408 (N_4408,N_3953,N_3712);
nand U4409 (N_4409,N_3038,N_3682);
or U4410 (N_4410,N_2939,N_3805);
or U4411 (N_4411,N_2706,N_3471);
xor U4412 (N_4412,N_3066,N_2856);
or U4413 (N_4413,N_3467,N_2986);
and U4414 (N_4414,N_2715,N_3378);
and U4415 (N_4415,N_3289,N_3321);
and U4416 (N_4416,N_2443,N_2742);
nand U4417 (N_4417,N_2331,N_2140);
nand U4418 (N_4418,N_3105,N_2405);
nand U4419 (N_4419,N_2263,N_3851);
nor U4420 (N_4420,N_2022,N_2723);
and U4421 (N_4421,N_2541,N_3100);
or U4422 (N_4422,N_2421,N_2136);
and U4423 (N_4423,N_2801,N_3451);
nand U4424 (N_4424,N_2419,N_3692);
and U4425 (N_4425,N_2214,N_3868);
or U4426 (N_4426,N_2067,N_2327);
nand U4427 (N_4427,N_3909,N_2866);
xnor U4428 (N_4428,N_3154,N_2393);
nand U4429 (N_4429,N_2778,N_3443);
and U4430 (N_4430,N_2896,N_3593);
nor U4431 (N_4431,N_2275,N_3590);
and U4432 (N_4432,N_3788,N_2488);
or U4433 (N_4433,N_3757,N_3136);
and U4434 (N_4434,N_2317,N_2444);
and U4435 (N_4435,N_2328,N_3507);
nor U4436 (N_4436,N_2251,N_2155);
nor U4437 (N_4437,N_2610,N_3440);
and U4438 (N_4438,N_2438,N_3350);
and U4439 (N_4439,N_2236,N_2569);
nor U4440 (N_4440,N_2542,N_3052);
and U4441 (N_4441,N_2898,N_2368);
nand U4442 (N_4442,N_2183,N_2159);
nor U4443 (N_4443,N_2557,N_2605);
and U4444 (N_4444,N_3774,N_3633);
and U4445 (N_4445,N_2996,N_3112);
and U4446 (N_4446,N_2059,N_3710);
nor U4447 (N_4447,N_2149,N_3452);
nand U4448 (N_4448,N_2844,N_2813);
nand U4449 (N_4449,N_2496,N_3475);
nand U4450 (N_4450,N_2991,N_3488);
and U4451 (N_4451,N_3182,N_2469);
and U4452 (N_4452,N_2756,N_3196);
nor U4453 (N_4453,N_3142,N_3663);
and U4454 (N_4454,N_3135,N_2759);
and U4455 (N_4455,N_2673,N_2584);
or U4456 (N_4456,N_2729,N_3133);
nand U4457 (N_4457,N_2456,N_3232);
and U4458 (N_4458,N_2755,N_3418);
and U4459 (N_4459,N_2276,N_3930);
nand U4460 (N_4460,N_3205,N_2824);
nand U4461 (N_4461,N_3949,N_3213);
or U4462 (N_4462,N_2769,N_2326);
nor U4463 (N_4463,N_2839,N_3681);
nor U4464 (N_4464,N_3817,N_3059);
xnor U4465 (N_4465,N_3405,N_2082);
or U4466 (N_4466,N_3931,N_3870);
and U4467 (N_4467,N_3897,N_2831);
nor U4468 (N_4468,N_2572,N_2919);
or U4469 (N_4469,N_2418,N_3445);
nand U4470 (N_4470,N_3640,N_2648);
nor U4471 (N_4471,N_3481,N_3299);
and U4472 (N_4472,N_2279,N_2539);
and U4473 (N_4473,N_3526,N_3423);
nor U4474 (N_4474,N_2434,N_2497);
nand U4475 (N_4475,N_2944,N_3419);
or U4476 (N_4476,N_3550,N_2549);
nor U4477 (N_4477,N_3401,N_3585);
nor U4478 (N_4478,N_3131,N_3271);
and U4479 (N_4479,N_3304,N_3257);
nor U4480 (N_4480,N_3272,N_2751);
xnor U4481 (N_4481,N_2166,N_3553);
and U4482 (N_4482,N_3705,N_2472);
nor U4483 (N_4483,N_2278,N_3356);
nor U4484 (N_4484,N_3490,N_2760);
or U4485 (N_4485,N_2877,N_2146);
nand U4486 (N_4486,N_3583,N_3461);
or U4487 (N_4487,N_2203,N_2120);
nor U4488 (N_4488,N_2354,N_2998);
and U4489 (N_4489,N_2026,N_2789);
or U4490 (N_4490,N_2474,N_2873);
and U4491 (N_4491,N_3844,N_3535);
nand U4492 (N_4492,N_3917,N_2876);
and U4493 (N_4493,N_2547,N_3660);
nor U4494 (N_4494,N_3760,N_3908);
xor U4495 (N_4495,N_2114,N_2807);
or U4496 (N_4496,N_3162,N_3521);
and U4497 (N_4497,N_2253,N_3827);
and U4498 (N_4498,N_3402,N_3524);
or U4499 (N_4499,N_3823,N_2306);
and U4500 (N_4500,N_2457,N_3575);
and U4501 (N_4501,N_3866,N_2604);
or U4502 (N_4502,N_3661,N_2323);
or U4503 (N_4503,N_2734,N_2150);
or U4504 (N_4504,N_3270,N_3470);
nor U4505 (N_4505,N_2036,N_2708);
and U4506 (N_4506,N_3062,N_3189);
nor U4507 (N_4507,N_2506,N_3081);
nand U4508 (N_4508,N_3508,N_3197);
or U4509 (N_4509,N_2064,N_3027);
nand U4510 (N_4510,N_2735,N_2775);
nor U4511 (N_4511,N_3484,N_3725);
nor U4512 (N_4512,N_3005,N_2946);
xnor U4513 (N_4513,N_3739,N_3706);
nand U4514 (N_4514,N_2997,N_2994);
and U4515 (N_4515,N_3157,N_3780);
xnor U4516 (N_4516,N_3843,N_2436);
or U4517 (N_4517,N_2016,N_2720);
nor U4518 (N_4518,N_3900,N_3750);
xnor U4519 (N_4519,N_2291,N_2383);
nand U4520 (N_4520,N_3983,N_2475);
or U4521 (N_4521,N_3744,N_2674);
nor U4522 (N_4522,N_3707,N_2467);
and U4523 (N_4523,N_2913,N_3456);
or U4524 (N_4524,N_2963,N_2316);
nand U4525 (N_4525,N_2105,N_2319);
nor U4526 (N_4526,N_3275,N_3649);
or U4527 (N_4527,N_3579,N_3872);
nor U4528 (N_4528,N_3117,N_3666);
and U4529 (N_4529,N_3130,N_3859);
nor U4530 (N_4530,N_3269,N_2220);
or U4531 (N_4531,N_2521,N_2427);
and U4532 (N_4532,N_3104,N_2980);
nor U4533 (N_4533,N_3533,N_2302);
and U4534 (N_4534,N_3214,N_3102);
nor U4535 (N_4535,N_2732,N_3398);
and U4536 (N_4536,N_2424,N_3569);
nand U4537 (N_4537,N_2088,N_3873);
xnor U4538 (N_4538,N_3826,N_3522);
nor U4539 (N_4539,N_2367,N_2682);
nor U4540 (N_4540,N_3956,N_2184);
and U4541 (N_4541,N_3160,N_3449);
nor U4542 (N_4542,N_2781,N_2607);
nand U4543 (N_4543,N_3684,N_2179);
nor U4544 (N_4544,N_2357,N_2477);
or U4545 (N_4545,N_3421,N_2738);
and U4546 (N_4546,N_2503,N_3124);
or U4547 (N_4547,N_2296,N_3555);
nand U4548 (N_4548,N_2827,N_3311);
nor U4549 (N_4549,N_2491,N_2106);
and U4550 (N_4550,N_2473,N_2705);
or U4551 (N_4551,N_2631,N_2777);
xor U4552 (N_4552,N_3934,N_3204);
nand U4553 (N_4553,N_2970,N_2449);
and U4554 (N_4554,N_3432,N_2054);
xnor U4555 (N_4555,N_2836,N_2823);
and U4556 (N_4556,N_3339,N_2835);
and U4557 (N_4557,N_2788,N_3014);
xnor U4558 (N_4558,N_2442,N_3811);
nor U4559 (N_4559,N_2257,N_2907);
or U4560 (N_4560,N_2653,N_3586);
nand U4561 (N_4561,N_3948,N_3375);
or U4562 (N_4562,N_3962,N_2630);
and U4563 (N_4563,N_2247,N_2335);
and U4564 (N_4564,N_2730,N_3810);
and U4565 (N_4565,N_3785,N_3120);
nor U4566 (N_4566,N_2176,N_2250);
and U4567 (N_4567,N_3057,N_2624);
or U4568 (N_4568,N_2591,N_3248);
xor U4569 (N_4569,N_2428,N_2538);
or U4570 (N_4570,N_2030,N_3085);
xor U4571 (N_4571,N_2007,N_3501);
or U4572 (N_4572,N_2070,N_2840);
and U4573 (N_4573,N_2837,N_2918);
and U4574 (N_4574,N_3972,N_2904);
nor U4575 (N_4575,N_3087,N_2484);
or U4576 (N_4576,N_3377,N_2485);
nor U4577 (N_4577,N_2154,N_3489);
xor U4578 (N_4578,N_2271,N_3442);
nor U4579 (N_4579,N_2350,N_3721);
nand U4580 (N_4580,N_3577,N_2083);
and U4581 (N_4581,N_2312,N_2034);
or U4582 (N_4582,N_2493,N_3325);
nor U4583 (N_4583,N_3371,N_3054);
and U4584 (N_4584,N_2492,N_2221);
and U4585 (N_4585,N_3916,N_2489);
nand U4586 (N_4586,N_3026,N_2232);
nand U4587 (N_4587,N_2834,N_3233);
or U4588 (N_4588,N_2286,N_2148);
nor U4589 (N_4589,N_2446,N_2583);
xor U4590 (N_4590,N_2096,N_3409);
nor U4591 (N_4591,N_2399,N_3284);
nor U4592 (N_4592,N_3767,N_3318);
and U4593 (N_4593,N_3391,N_2726);
nand U4594 (N_4594,N_2574,N_3388);
nor U4595 (N_4595,N_2804,N_2262);
nor U4596 (N_4596,N_3515,N_3551);
xnor U4597 (N_4597,N_2693,N_3546);
or U4598 (N_4598,N_2012,N_3893);
and U4599 (N_4599,N_2037,N_3802);
nor U4600 (N_4600,N_2828,N_2060);
nand U4601 (N_4601,N_3879,N_2525);
or U4602 (N_4602,N_3046,N_3061);
nor U4603 (N_4603,N_2780,N_2141);
or U4604 (N_4604,N_3833,N_3404);
nand U4605 (N_4605,N_2075,N_2077);
and U4606 (N_4606,N_2809,N_3623);
nor U4607 (N_4607,N_3185,N_2750);
nand U4608 (N_4608,N_3964,N_3659);
nor U4609 (N_4609,N_3651,N_2843);
nand U4610 (N_4610,N_2097,N_3610);
xor U4611 (N_4611,N_3190,N_2209);
nor U4612 (N_4612,N_2391,N_2344);
nand U4613 (N_4613,N_3582,N_3528);
nor U4614 (N_4614,N_3691,N_2724);
nand U4615 (N_4615,N_2707,N_2112);
or U4616 (N_4616,N_3263,N_2964);
or U4617 (N_4617,N_3717,N_2905);
xor U4618 (N_4618,N_2594,N_2052);
nand U4619 (N_4619,N_3331,N_3718);
xor U4620 (N_4620,N_3654,N_2847);
and U4621 (N_4621,N_2360,N_2256);
nor U4622 (N_4622,N_3446,N_3538);
or U4623 (N_4623,N_3963,N_2981);
or U4624 (N_4624,N_3017,N_3206);
and U4625 (N_4625,N_2134,N_3023);
and U4626 (N_4626,N_2277,N_2661);
or U4627 (N_4627,N_2143,N_3732);
nor U4628 (N_4628,N_2803,N_2011);
nor U4629 (N_4629,N_3015,N_3899);
nand U4630 (N_4630,N_2573,N_3266);
nor U4631 (N_4631,N_3273,N_3406);
nor U4632 (N_4632,N_3434,N_3694);
and U4633 (N_4633,N_2758,N_3003);
or U4634 (N_4634,N_2151,N_2274);
and U4635 (N_4635,N_3831,N_3373);
or U4636 (N_4636,N_2713,N_3327);
nand U4637 (N_4637,N_2001,N_2666);
nand U4638 (N_4638,N_3932,N_3227);
and U4639 (N_4639,N_3672,N_2170);
or U4640 (N_4640,N_3574,N_2692);
or U4641 (N_4641,N_2698,N_2394);
xor U4642 (N_4642,N_3001,N_2109);
xnor U4643 (N_4643,N_2337,N_3880);
nor U4644 (N_4644,N_2786,N_3862);
nand U4645 (N_4645,N_3007,N_3089);
or U4646 (N_4646,N_2971,N_3611);
nor U4647 (N_4647,N_2787,N_2290);
nand U4648 (N_4648,N_2315,N_2701);
nand U4649 (N_4649,N_2450,N_2244);
nor U4650 (N_4650,N_3018,N_3977);
nand U4651 (N_4651,N_3147,N_2853);
nand U4652 (N_4652,N_3933,N_2239);
nor U4653 (N_4653,N_2314,N_3093);
or U4654 (N_4654,N_2625,N_3161);
or U4655 (N_4655,N_3358,N_2960);
or U4656 (N_4656,N_2309,N_3984);
and U4657 (N_4657,N_2677,N_3256);
or U4658 (N_4658,N_3806,N_3492);
nand U4659 (N_4659,N_2576,N_2973);
nor U4660 (N_4660,N_3856,N_2311);
nor U4661 (N_4661,N_3713,N_3762);
nor U4662 (N_4662,N_3549,N_2883);
and U4663 (N_4663,N_2922,N_2559);
nor U4664 (N_4664,N_2841,N_3485);
nand U4665 (N_4665,N_2197,N_2476);
xnor U4666 (N_4666,N_2748,N_2798);
or U4667 (N_4667,N_3156,N_2207);
nand U4668 (N_4668,N_3669,N_2911);
and U4669 (N_4669,N_2425,N_3889);
and U4670 (N_4670,N_2095,N_3861);
and U4671 (N_4671,N_2854,N_3606);
and U4672 (N_4672,N_2009,N_3671);
nand U4673 (N_4673,N_3011,N_3808);
xor U4674 (N_4674,N_2177,N_2481);
xnor U4675 (N_4675,N_2002,N_2376);
or U4676 (N_4676,N_2000,N_3002);
xor U4677 (N_4677,N_3891,N_2721);
nor U4678 (N_4678,N_2717,N_2505);
nor U4679 (N_4679,N_2924,N_3158);
nand U4680 (N_4680,N_2432,N_3967);
nor U4681 (N_4681,N_3882,N_2581);
nor U4682 (N_4682,N_3940,N_2599);
xor U4683 (N_4683,N_3482,N_2258);
nand U4684 (N_4684,N_2887,N_3163);
or U4685 (N_4685,N_2407,N_3955);
nand U4686 (N_4686,N_3376,N_2933);
nor U4687 (N_4687,N_2388,N_3253);
xnor U4688 (N_4688,N_3509,N_2626);
nand U4689 (N_4689,N_2999,N_2031);
xnor U4690 (N_4690,N_3417,N_3689);
and U4691 (N_4691,N_3472,N_2231);
nor U4692 (N_4692,N_3267,N_3519);
xnor U4693 (N_4693,N_2211,N_2968);
nand U4694 (N_4694,N_2502,N_3600);
nor U4695 (N_4695,N_3219,N_2058);
nand U4696 (N_4696,N_3752,N_2566);
nand U4697 (N_4697,N_3946,N_3019);
nand U4698 (N_4698,N_2551,N_2370);
or U4699 (N_4699,N_3252,N_2249);
xnor U4700 (N_4700,N_3169,N_2417);
nand U4701 (N_4701,N_3925,N_3647);
nor U4702 (N_4702,N_3884,N_2003);
or U4703 (N_4703,N_2865,N_3394);
and U4704 (N_4704,N_2406,N_2719);
nand U4705 (N_4705,N_3179,N_2074);
nand U4706 (N_4706,N_2065,N_3107);
nor U4707 (N_4707,N_3173,N_3487);
or U4708 (N_4708,N_2348,N_3403);
xor U4709 (N_4709,N_2544,N_2135);
and U4710 (N_4710,N_3372,N_3416);
and U4711 (N_4711,N_3363,N_2188);
nor U4712 (N_4712,N_2953,N_3775);
nor U4713 (N_4713,N_2645,N_3067);
nand U4714 (N_4714,N_3877,N_3016);
xor U4715 (N_4715,N_3708,N_2955);
nor U4716 (N_4716,N_3990,N_2728);
xor U4717 (N_4717,N_2737,N_2196);
nor U4718 (N_4718,N_3943,N_3829);
xnor U4719 (N_4719,N_3441,N_2389);
nor U4720 (N_4720,N_3393,N_2808);
nand U4721 (N_4721,N_3797,N_3994);
nor U4722 (N_4722,N_3719,N_3561);
nor U4723 (N_4723,N_3174,N_2024);
or U4724 (N_4724,N_3364,N_3544);
and U4725 (N_4725,N_2182,N_2588);
or U4726 (N_4726,N_3801,N_3307);
nor U4727 (N_4727,N_3580,N_2859);
nor U4728 (N_4728,N_2765,N_3537);
or U4729 (N_4729,N_3541,N_2554);
nand U4730 (N_4730,N_3965,N_2175);
nand U4731 (N_4731,N_3740,N_3074);
and U4732 (N_4732,N_2218,N_2053);
and U4733 (N_4733,N_2254,N_2829);
nand U4734 (N_4734,N_2223,N_2942);
and U4735 (N_4735,N_2894,N_3939);
and U4736 (N_4736,N_3742,N_3098);
nand U4737 (N_4737,N_2871,N_3078);
and U4738 (N_4738,N_2501,N_2643);
or U4739 (N_4739,N_2858,N_2364);
and U4740 (N_4740,N_3155,N_2716);
nor U4741 (N_4741,N_2379,N_3499);
xor U4742 (N_4742,N_2672,N_3720);
and U4743 (N_4743,N_3929,N_2324);
and U4744 (N_4744,N_2895,N_3881);
nor U4745 (N_4745,N_2057,N_2241);
and U4746 (N_4746,N_3906,N_3241);
or U4747 (N_4747,N_2885,N_3119);
nor U4748 (N_4748,N_2628,N_2916);
xnor U4749 (N_4749,N_3869,N_3226);
xnor U4750 (N_4750,N_3560,N_2173);
or U4751 (N_4751,N_2300,N_2224);
and U4752 (N_4752,N_2697,N_2632);
xnor U4753 (N_4753,N_2906,N_2763);
or U4754 (N_4754,N_2878,N_2686);
or U4755 (N_4755,N_3336,N_3217);
and U4756 (N_4756,N_3941,N_3723);
and U4757 (N_4757,N_3578,N_3186);
nor U4758 (N_4758,N_3690,N_3730);
nor U4759 (N_4759,N_2650,N_2345);
or U4760 (N_4760,N_3290,N_2772);
nand U4761 (N_4761,N_3596,N_3631);
or U4762 (N_4762,N_2138,N_3286);
or U4763 (N_4763,N_3756,N_3060);
nor U4764 (N_4764,N_2131,N_2347);
nand U4765 (N_4765,N_3748,N_3453);
nor U4766 (N_4766,N_2416,N_2611);
xor U4767 (N_4767,N_2259,N_2797);
and U4768 (N_4768,N_3978,N_3450);
nor U4769 (N_4769,N_3607,N_3570);
or U4770 (N_4770,N_2465,N_3022);
or U4771 (N_4771,N_3478,N_3795);
nand U4772 (N_4772,N_2480,N_3181);
nand U4773 (N_4773,N_2318,N_3193);
nand U4774 (N_4774,N_3892,N_2512);
or U4775 (N_4775,N_3597,N_2334);
nand U4776 (N_4776,N_3687,N_3895);
and U4777 (N_4777,N_3079,N_2727);
nand U4778 (N_4778,N_2664,N_2932);
or U4779 (N_4779,N_3348,N_3923);
or U4780 (N_4780,N_3447,N_3601);
and U4781 (N_4781,N_2129,N_2889);
nor U4782 (N_4782,N_3584,N_3265);
or U4783 (N_4783,N_2237,N_3400);
or U4784 (N_4784,N_3626,N_3650);
nor U4785 (N_4785,N_3938,N_3159);
nand U4786 (N_4786,N_2663,N_2213);
nor U4787 (N_4787,N_3552,N_2983);
and U4788 (N_4788,N_2222,N_3076);
nor U4789 (N_4789,N_3928,N_2032);
or U4790 (N_4790,N_2471,N_2520);
and U4791 (N_4791,N_3261,N_3305);
xnor U4792 (N_4792,N_3312,N_2441);
nor U4793 (N_4793,N_2800,N_3697);
nand U4794 (N_4794,N_2952,N_3006);
or U4795 (N_4795,N_2226,N_3683);
nand U4796 (N_4796,N_2361,N_3280);
xor U4797 (N_4797,N_2283,N_2774);
and U4798 (N_4798,N_3337,N_2210);
or U4799 (N_4799,N_2582,N_2540);
or U4800 (N_4800,N_3031,N_2128);
xor U4801 (N_4801,N_2908,N_3091);
or U4802 (N_4802,N_3342,N_3465);
nand U4803 (N_4803,N_3828,N_3413);
or U4804 (N_4804,N_2305,N_2092);
and U4805 (N_4805,N_3122,N_2517);
or U4806 (N_4806,N_2242,N_2111);
nand U4807 (N_4807,N_3731,N_3322);
nor U4808 (N_4808,N_2608,N_2343);
or U4809 (N_4809,N_3149,N_3668);
and U4810 (N_4810,N_3477,N_2433);
nand U4811 (N_4811,N_2010,N_2593);
nand U4812 (N_4812,N_2794,N_3072);
and U4813 (N_4813,N_2216,N_2656);
or U4814 (N_4814,N_2637,N_2548);
and U4815 (N_4815,N_2560,N_3032);
and U4816 (N_4816,N_2704,N_2849);
nor U4817 (N_4817,N_2902,N_2269);
nor U4818 (N_4818,N_2872,N_2192);
and U4819 (N_4819,N_3864,N_2440);
nand U4820 (N_4820,N_2867,N_3558);
and U4821 (N_4821,N_3088,N_3357);
nor U4822 (N_4822,N_3656,N_2005);
nor U4823 (N_4823,N_2325,N_2917);
nand U4824 (N_4824,N_3587,N_2680);
and U4825 (N_4825,N_2137,N_3410);
or U4826 (N_4826,N_2206,N_3251);
xnor U4827 (N_4827,N_2035,N_2006);
xnor U4828 (N_4828,N_3988,N_2121);
nand U4829 (N_4829,N_2567,N_2157);
or U4830 (N_4830,N_3995,N_2459);
or U4831 (N_4831,N_2923,N_2431);
nand U4832 (N_4832,N_2375,N_3945);
nor U4833 (N_4833,N_2930,N_3071);
and U4834 (N_4834,N_3437,N_2752);
nor U4835 (N_4835,N_3612,N_3306);
nor U4836 (N_4836,N_2987,N_3547);
nand U4837 (N_4837,N_3497,N_3771);
nor U4838 (N_4838,N_3959,N_2085);
and U4839 (N_4839,N_2511,N_3145);
nand U4840 (N_4840,N_3620,N_2528);
nor U4841 (N_4841,N_3040,N_3781);
nor U4842 (N_4842,N_2779,N_2690);
nand U4843 (N_4843,N_2580,N_3867);
xor U4844 (N_4844,N_2508,N_2061);
or U4845 (N_4845,N_3430,N_3765);
nor U4846 (N_4846,N_2976,N_2832);
nand U4847 (N_4847,N_2227,N_3562);
or U4848 (N_4848,N_2818,N_2039);
xor U4849 (N_4849,N_2402,N_2101);
nand U4850 (N_4850,N_2043,N_2687);
or U4851 (N_4851,N_3736,N_3480);
or U4852 (N_4852,N_3875,N_2949);
and U4853 (N_4853,N_3602,N_2056);
and U4854 (N_4854,N_2927,N_2815);
nand U4855 (N_4855,N_2193,N_3726);
nor U4856 (N_4856,N_3386,N_3860);
nor U4857 (N_4857,N_2654,N_2409);
nor U4858 (N_4858,N_2945,N_2094);
nand U4859 (N_4859,N_3819,N_2791);
xor U4860 (N_4860,N_2169,N_3302);
and U4861 (N_4861,N_3874,N_2621);
and U4862 (N_4862,N_2984,N_2240);
or U4863 (N_4863,N_3469,N_2395);
or U4864 (N_4864,N_2814,N_3351);
and U4865 (N_4865,N_3696,N_2063);
and U4866 (N_4866,N_2747,N_3379);
and U4867 (N_4867,N_2523,N_2116);
or U4868 (N_4868,N_2616,N_2051);
nor U4869 (N_4869,N_2852,N_3438);
nor U4870 (N_4870,N_3320,N_3199);
or U4871 (N_4871,N_3758,N_2817);
and U4872 (N_4872,N_3466,N_2870);
and U4873 (N_4873,N_2201,N_3310);
nor U4874 (N_4874,N_3581,N_2771);
or U4875 (N_4875,N_3209,N_3086);
nand U4876 (N_4876,N_3143,N_2178);
nand U4877 (N_4877,N_3523,N_3565);
xnor U4878 (N_4878,N_3849,N_3791);
and U4879 (N_4879,N_3293,N_2558);
and U4880 (N_4880,N_3772,N_2398);
or U4881 (N_4881,N_3374,N_3353);
or U4882 (N_4882,N_2671,N_2359);
and U4883 (N_4883,N_2776,N_3298);
and U4884 (N_4884,N_3110,N_3425);
nand U4885 (N_4885,N_2561,N_3809);
and U4886 (N_4886,N_2816,N_2874);
nand U4887 (N_4887,N_3800,N_3518);
nand U4888 (N_4888,N_2884,N_2299);
or U4889 (N_4889,N_3335,N_3894);
and U4890 (N_4890,N_2298,N_3836);
xnor U4891 (N_4891,N_3632,N_2806);
and U4892 (N_4892,N_2163,N_2519);
or U4893 (N_4893,N_3218,N_2267);
nor U4894 (N_4894,N_3354,N_2793);
and U4895 (N_4895,N_3171,N_2396);
and U4896 (N_4896,N_3680,N_2107);
or U4897 (N_4897,N_2499,N_3184);
and U4898 (N_4898,N_2069,N_3319);
xnor U4899 (N_4899,N_2589,N_2534);
nand U4900 (N_4900,N_2158,N_2689);
xnor U4901 (N_4901,N_2568,N_2982);
nand U4902 (N_4902,N_3138,N_2185);
and U4903 (N_4903,N_2746,N_3918);
xnor U4904 (N_4904,N_2646,N_3950);
or U4905 (N_4905,N_3543,N_3755);
and U4906 (N_4906,N_2612,N_2404);
and U4907 (N_4907,N_3203,N_2770);
nor U4908 (N_4908,N_2875,N_3113);
nor U4909 (N_4909,N_3545,N_3330);
nor U4910 (N_4910,N_3200,N_2382);
and U4911 (N_4911,N_3084,N_3345);
and U4912 (N_4912,N_2046,N_3503);
or U4913 (N_4913,N_3594,N_3848);
and U4914 (N_4914,N_2845,N_3175);
nor U4915 (N_4915,N_2071,N_3099);
or U4916 (N_4916,N_2147,N_2021);
and U4917 (N_4917,N_3904,N_3464);
nor U4918 (N_4918,N_3338,N_3728);
nand U4919 (N_4919,N_3210,N_2926);
and U4920 (N_4920,N_2285,N_2920);
and U4921 (N_4921,N_3359,N_2850);
nand U4922 (N_4922,N_2792,N_3505);
nor U4923 (N_4923,N_2377,N_2940);
nor U4924 (N_4924,N_2280,N_3975);
nor U4925 (N_4925,N_3030,N_2928);
nor U4926 (N_4926,N_2620,N_3751);
or U4927 (N_4927,N_2869,N_3947);
nor U4928 (N_4928,N_3041,N_3734);
and U4929 (N_4929,N_2430,N_3534);
and U4930 (N_4930,N_2642,N_2550);
or U4931 (N_4931,N_3786,N_3999);
and U4932 (N_4932,N_3211,N_2199);
nor U4933 (N_4933,N_3703,N_3698);
xor U4934 (N_4934,N_3820,N_3237);
nor U4935 (N_4935,N_3926,N_3677);
nor U4936 (N_4936,N_3246,N_2979);
and U4937 (N_4937,N_2266,N_2014);
nand U4938 (N_4938,N_3390,N_2172);
or U4939 (N_4939,N_2951,N_3129);
nor U4940 (N_4940,N_3605,N_3850);
xor U4941 (N_4941,N_2340,N_2563);
nor U4942 (N_4942,N_2495,N_3229);
nor U4943 (N_4943,N_2710,N_2510);
or U4944 (N_4944,N_2522,N_3170);
nand U4945 (N_4945,N_2810,N_2868);
xor U4946 (N_4946,N_2372,N_3568);
and U4947 (N_4947,N_3749,N_3838);
or U4948 (N_4948,N_2187,N_2486);
nor U4949 (N_4949,N_3281,N_3937);
and U4950 (N_4950,N_3111,N_3799);
nand U4951 (N_4951,N_2586,N_3825);
nor U4952 (N_4952,N_3202,N_3037);
nand U4953 (N_4953,N_3885,N_2764);
and U4954 (N_4954,N_2595,N_3329);
and U4955 (N_4955,N_2745,N_3095);
nand U4956 (N_4956,N_3282,N_2571);
nor U4957 (N_4957,N_2081,N_3816);
nor U4958 (N_4958,N_3638,N_2762);
or U4959 (N_4959,N_2504,N_3784);
nand U4960 (N_4960,N_3050,N_2974);
and U4961 (N_4961,N_3531,N_2848);
nor U4962 (N_4962,N_2235,N_2352);
or U4963 (N_4963,N_2004,N_3258);
nand U4964 (N_4964,N_3064,N_3588);
xor U4965 (N_4965,N_3194,N_2500);
xnor U4966 (N_4966,N_3128,N_2676);
nor U4967 (N_4967,N_3985,N_3741);
nand U4968 (N_4968,N_3954,N_3483);
nand U4969 (N_4969,N_3439,N_2513);
nor U4970 (N_4970,N_2099,N_3225);
nand U4971 (N_4971,N_2860,N_3334);
nor U4972 (N_4972,N_3463,N_3912);
nor U4973 (N_4973,N_2217,N_3674);
nor U4974 (N_4974,N_3563,N_3506);
xor U4975 (N_4975,N_2969,N_3457);
and U4976 (N_4976,N_2313,N_2657);
xor U4977 (N_4977,N_2133,N_3234);
or U4978 (N_4978,N_3814,N_2180);
or U4979 (N_4979,N_3630,N_2093);
nor U4980 (N_4980,N_2695,N_3387);
nor U4981 (N_4981,N_3244,N_2281);
or U4982 (N_4982,N_3573,N_2931);
or U4983 (N_4983,N_2929,N_3249);
and U4984 (N_4984,N_2458,N_3276);
or U4985 (N_4985,N_3332,N_3114);
nor U4986 (N_4986,N_3993,N_2606);
nand U4987 (N_4987,N_2543,N_3236);
and U4988 (N_4988,N_2062,N_2397);
and U4989 (N_4989,N_3835,N_3025);
or U4990 (N_4990,N_2233,N_2454);
xor U4991 (N_4991,N_3368,N_2103);
and U4992 (N_4992,N_3525,N_3392);
nor U4993 (N_4993,N_3053,N_2935);
nor U4994 (N_4994,N_2270,N_2080);
nor U4995 (N_4995,N_3852,N_3700);
xor U4996 (N_4996,N_2992,N_2355);
or U4997 (N_4997,N_3628,N_2943);
nand U4998 (N_4998,N_3004,N_2117);
and U4999 (N_4999,N_2385,N_3818);
nand U5000 (N_5000,N_2580,N_3067);
and U5001 (N_5001,N_2389,N_2677);
and U5002 (N_5002,N_2786,N_3635);
and U5003 (N_5003,N_2639,N_3931);
xnor U5004 (N_5004,N_3331,N_3629);
xnor U5005 (N_5005,N_2389,N_2510);
nand U5006 (N_5006,N_3737,N_3209);
nor U5007 (N_5007,N_3190,N_2314);
or U5008 (N_5008,N_2070,N_2116);
nand U5009 (N_5009,N_2927,N_2242);
nand U5010 (N_5010,N_3223,N_3536);
or U5011 (N_5011,N_3318,N_3402);
nand U5012 (N_5012,N_3169,N_2409);
nand U5013 (N_5013,N_2984,N_2542);
nor U5014 (N_5014,N_2857,N_3105);
xor U5015 (N_5015,N_3528,N_2125);
nor U5016 (N_5016,N_2240,N_3576);
and U5017 (N_5017,N_2527,N_2253);
nor U5018 (N_5018,N_2379,N_2946);
or U5019 (N_5019,N_3532,N_2891);
nor U5020 (N_5020,N_3559,N_3691);
or U5021 (N_5021,N_2243,N_2613);
nor U5022 (N_5022,N_2059,N_2287);
nand U5023 (N_5023,N_3155,N_3618);
and U5024 (N_5024,N_2146,N_3733);
xnor U5025 (N_5025,N_3883,N_2243);
nor U5026 (N_5026,N_3246,N_3452);
xor U5027 (N_5027,N_3459,N_2269);
nor U5028 (N_5028,N_3622,N_2276);
nor U5029 (N_5029,N_3615,N_3288);
or U5030 (N_5030,N_3208,N_3205);
and U5031 (N_5031,N_2880,N_2669);
nand U5032 (N_5032,N_3309,N_3882);
and U5033 (N_5033,N_3847,N_3286);
nor U5034 (N_5034,N_3120,N_2471);
nand U5035 (N_5035,N_2876,N_2213);
xor U5036 (N_5036,N_2395,N_3062);
nor U5037 (N_5037,N_2114,N_2204);
xor U5038 (N_5038,N_3018,N_3702);
and U5039 (N_5039,N_3167,N_2057);
xnor U5040 (N_5040,N_3678,N_3790);
nand U5041 (N_5041,N_2586,N_2915);
or U5042 (N_5042,N_2293,N_2497);
or U5043 (N_5043,N_2823,N_3663);
nor U5044 (N_5044,N_2717,N_3835);
nor U5045 (N_5045,N_3545,N_3805);
or U5046 (N_5046,N_2026,N_3215);
and U5047 (N_5047,N_3872,N_2438);
nor U5048 (N_5048,N_2587,N_2452);
nand U5049 (N_5049,N_2595,N_2834);
xnor U5050 (N_5050,N_3205,N_2951);
or U5051 (N_5051,N_3292,N_3710);
nor U5052 (N_5052,N_3262,N_3353);
and U5053 (N_5053,N_2525,N_2197);
or U5054 (N_5054,N_3440,N_2493);
nand U5055 (N_5055,N_2748,N_3964);
or U5056 (N_5056,N_2273,N_2426);
xor U5057 (N_5057,N_2422,N_3925);
and U5058 (N_5058,N_3838,N_2693);
xor U5059 (N_5059,N_2375,N_2590);
nor U5060 (N_5060,N_3066,N_2973);
nor U5061 (N_5061,N_3167,N_3968);
xor U5062 (N_5062,N_2539,N_3537);
and U5063 (N_5063,N_2500,N_3792);
and U5064 (N_5064,N_2221,N_2731);
nor U5065 (N_5065,N_2671,N_3037);
nand U5066 (N_5066,N_2770,N_3082);
or U5067 (N_5067,N_2591,N_2946);
nor U5068 (N_5068,N_2606,N_3911);
or U5069 (N_5069,N_3663,N_2540);
xnor U5070 (N_5070,N_2430,N_3582);
nand U5071 (N_5071,N_2648,N_2231);
xnor U5072 (N_5072,N_2407,N_2403);
nor U5073 (N_5073,N_3990,N_3767);
and U5074 (N_5074,N_2908,N_2471);
nand U5075 (N_5075,N_3254,N_2262);
and U5076 (N_5076,N_3467,N_2859);
nor U5077 (N_5077,N_3677,N_2099);
or U5078 (N_5078,N_2807,N_3831);
or U5079 (N_5079,N_3332,N_2324);
or U5080 (N_5080,N_3348,N_3667);
nand U5081 (N_5081,N_3292,N_2001);
nand U5082 (N_5082,N_3568,N_2003);
and U5083 (N_5083,N_3506,N_2030);
nand U5084 (N_5084,N_2315,N_2206);
nand U5085 (N_5085,N_3539,N_2606);
and U5086 (N_5086,N_2860,N_2566);
nor U5087 (N_5087,N_2403,N_2712);
and U5088 (N_5088,N_2796,N_3324);
or U5089 (N_5089,N_3138,N_2174);
or U5090 (N_5090,N_3486,N_3493);
nand U5091 (N_5091,N_3876,N_3840);
xor U5092 (N_5092,N_2019,N_3192);
or U5093 (N_5093,N_3732,N_3815);
or U5094 (N_5094,N_2859,N_2247);
or U5095 (N_5095,N_2891,N_3021);
nor U5096 (N_5096,N_2575,N_3919);
xor U5097 (N_5097,N_2773,N_3779);
nand U5098 (N_5098,N_2327,N_2721);
or U5099 (N_5099,N_2846,N_3378);
nand U5100 (N_5100,N_2640,N_2314);
nor U5101 (N_5101,N_2807,N_3001);
nor U5102 (N_5102,N_3557,N_3349);
nand U5103 (N_5103,N_3227,N_3438);
xor U5104 (N_5104,N_3241,N_2485);
xor U5105 (N_5105,N_3971,N_3340);
or U5106 (N_5106,N_2099,N_2958);
or U5107 (N_5107,N_2736,N_3401);
or U5108 (N_5108,N_3529,N_3019);
nand U5109 (N_5109,N_3753,N_3109);
nand U5110 (N_5110,N_2940,N_2034);
or U5111 (N_5111,N_3052,N_2240);
or U5112 (N_5112,N_2868,N_2256);
or U5113 (N_5113,N_2675,N_2304);
and U5114 (N_5114,N_3471,N_3762);
nor U5115 (N_5115,N_2830,N_3227);
xnor U5116 (N_5116,N_3072,N_2178);
nand U5117 (N_5117,N_2843,N_3925);
nor U5118 (N_5118,N_3084,N_3752);
nand U5119 (N_5119,N_2496,N_3976);
and U5120 (N_5120,N_2852,N_2450);
and U5121 (N_5121,N_2171,N_3356);
nor U5122 (N_5122,N_3860,N_3259);
xor U5123 (N_5123,N_2032,N_2649);
and U5124 (N_5124,N_2653,N_2934);
nand U5125 (N_5125,N_3511,N_3856);
xnor U5126 (N_5126,N_3482,N_2571);
or U5127 (N_5127,N_3694,N_2789);
nand U5128 (N_5128,N_3953,N_2254);
nand U5129 (N_5129,N_3719,N_3590);
xnor U5130 (N_5130,N_2259,N_3079);
nor U5131 (N_5131,N_2475,N_3758);
or U5132 (N_5132,N_3698,N_3637);
xor U5133 (N_5133,N_3418,N_3528);
xnor U5134 (N_5134,N_2473,N_2853);
or U5135 (N_5135,N_2923,N_2094);
nor U5136 (N_5136,N_3939,N_3300);
nor U5137 (N_5137,N_3984,N_3919);
or U5138 (N_5138,N_3560,N_3127);
nand U5139 (N_5139,N_3230,N_3499);
nand U5140 (N_5140,N_3115,N_3407);
or U5141 (N_5141,N_3748,N_2925);
or U5142 (N_5142,N_2650,N_2535);
and U5143 (N_5143,N_2459,N_3906);
nor U5144 (N_5144,N_3905,N_3321);
or U5145 (N_5145,N_2005,N_3785);
nor U5146 (N_5146,N_2749,N_2082);
or U5147 (N_5147,N_2924,N_3594);
nand U5148 (N_5148,N_2590,N_2854);
nand U5149 (N_5149,N_3082,N_2454);
and U5150 (N_5150,N_3677,N_3907);
and U5151 (N_5151,N_2204,N_2454);
nand U5152 (N_5152,N_3444,N_3327);
and U5153 (N_5153,N_2404,N_2691);
nand U5154 (N_5154,N_2745,N_3167);
nor U5155 (N_5155,N_3974,N_2311);
or U5156 (N_5156,N_3344,N_2253);
nand U5157 (N_5157,N_2444,N_3257);
xnor U5158 (N_5158,N_3080,N_3347);
nand U5159 (N_5159,N_3490,N_2745);
nand U5160 (N_5160,N_3215,N_2163);
nand U5161 (N_5161,N_2858,N_2720);
nand U5162 (N_5162,N_3327,N_2084);
nand U5163 (N_5163,N_2490,N_3475);
nand U5164 (N_5164,N_3772,N_2569);
nand U5165 (N_5165,N_3213,N_3960);
xor U5166 (N_5166,N_3401,N_3720);
and U5167 (N_5167,N_2517,N_2105);
or U5168 (N_5168,N_2920,N_2181);
or U5169 (N_5169,N_2047,N_3647);
and U5170 (N_5170,N_3286,N_3899);
nor U5171 (N_5171,N_2621,N_2169);
nand U5172 (N_5172,N_3980,N_2662);
nand U5173 (N_5173,N_3935,N_3041);
or U5174 (N_5174,N_2792,N_2250);
nand U5175 (N_5175,N_3939,N_3959);
nand U5176 (N_5176,N_3916,N_3596);
and U5177 (N_5177,N_2825,N_3100);
and U5178 (N_5178,N_2296,N_2649);
or U5179 (N_5179,N_3795,N_2909);
nand U5180 (N_5180,N_3537,N_3003);
xor U5181 (N_5181,N_2286,N_3115);
nand U5182 (N_5182,N_3924,N_2123);
nand U5183 (N_5183,N_2718,N_2601);
xnor U5184 (N_5184,N_3756,N_3435);
nand U5185 (N_5185,N_3710,N_3169);
nand U5186 (N_5186,N_3959,N_3010);
and U5187 (N_5187,N_2426,N_2927);
and U5188 (N_5188,N_3688,N_3422);
or U5189 (N_5189,N_3275,N_3330);
or U5190 (N_5190,N_3349,N_3376);
or U5191 (N_5191,N_2845,N_3487);
nor U5192 (N_5192,N_2793,N_3207);
nand U5193 (N_5193,N_2398,N_2979);
xnor U5194 (N_5194,N_3312,N_3987);
xnor U5195 (N_5195,N_2418,N_3847);
or U5196 (N_5196,N_2950,N_2435);
and U5197 (N_5197,N_2231,N_2472);
and U5198 (N_5198,N_2903,N_2703);
nor U5199 (N_5199,N_2568,N_2784);
or U5200 (N_5200,N_3751,N_3701);
or U5201 (N_5201,N_3529,N_3237);
xor U5202 (N_5202,N_2910,N_2029);
nand U5203 (N_5203,N_3637,N_3366);
or U5204 (N_5204,N_2681,N_3087);
xnor U5205 (N_5205,N_3391,N_3843);
nand U5206 (N_5206,N_2885,N_3137);
and U5207 (N_5207,N_2691,N_3261);
and U5208 (N_5208,N_3108,N_2760);
nor U5209 (N_5209,N_2604,N_3383);
nor U5210 (N_5210,N_3326,N_3019);
and U5211 (N_5211,N_3396,N_2998);
nor U5212 (N_5212,N_3730,N_2839);
nand U5213 (N_5213,N_2363,N_3095);
or U5214 (N_5214,N_2004,N_2883);
nor U5215 (N_5215,N_3849,N_3987);
or U5216 (N_5216,N_3095,N_2888);
xor U5217 (N_5217,N_3313,N_2013);
nor U5218 (N_5218,N_3130,N_2164);
nand U5219 (N_5219,N_3182,N_2498);
nor U5220 (N_5220,N_2466,N_2366);
nor U5221 (N_5221,N_3515,N_2643);
nor U5222 (N_5222,N_2547,N_3665);
xor U5223 (N_5223,N_3540,N_2697);
xor U5224 (N_5224,N_2040,N_2091);
and U5225 (N_5225,N_3247,N_2713);
and U5226 (N_5226,N_2100,N_3835);
or U5227 (N_5227,N_2033,N_2268);
and U5228 (N_5228,N_3182,N_2701);
nor U5229 (N_5229,N_2997,N_2003);
and U5230 (N_5230,N_3945,N_3775);
nor U5231 (N_5231,N_3918,N_2497);
nor U5232 (N_5232,N_3650,N_3188);
or U5233 (N_5233,N_2596,N_3448);
or U5234 (N_5234,N_3515,N_2051);
and U5235 (N_5235,N_2388,N_3103);
nand U5236 (N_5236,N_3201,N_3033);
nand U5237 (N_5237,N_2846,N_3757);
xnor U5238 (N_5238,N_2785,N_2966);
and U5239 (N_5239,N_3689,N_2554);
nor U5240 (N_5240,N_3000,N_2284);
nand U5241 (N_5241,N_2212,N_2598);
or U5242 (N_5242,N_3722,N_3631);
or U5243 (N_5243,N_2469,N_3436);
and U5244 (N_5244,N_3443,N_3111);
or U5245 (N_5245,N_3111,N_2428);
nand U5246 (N_5246,N_3795,N_3398);
and U5247 (N_5247,N_2196,N_2906);
or U5248 (N_5248,N_2161,N_3752);
and U5249 (N_5249,N_3772,N_3865);
nand U5250 (N_5250,N_3665,N_2816);
nand U5251 (N_5251,N_2178,N_3890);
and U5252 (N_5252,N_2127,N_3899);
nand U5253 (N_5253,N_3796,N_2679);
nor U5254 (N_5254,N_3215,N_2022);
or U5255 (N_5255,N_3326,N_2115);
xor U5256 (N_5256,N_3482,N_3005);
and U5257 (N_5257,N_3263,N_2149);
or U5258 (N_5258,N_3472,N_2297);
and U5259 (N_5259,N_3043,N_2410);
nand U5260 (N_5260,N_3421,N_3891);
nor U5261 (N_5261,N_2346,N_3008);
nor U5262 (N_5262,N_3632,N_3819);
xor U5263 (N_5263,N_2989,N_3116);
or U5264 (N_5264,N_2192,N_2720);
or U5265 (N_5265,N_2474,N_2618);
nand U5266 (N_5266,N_3720,N_2844);
or U5267 (N_5267,N_2547,N_2078);
and U5268 (N_5268,N_2692,N_2329);
and U5269 (N_5269,N_2107,N_2100);
nand U5270 (N_5270,N_2093,N_3899);
nor U5271 (N_5271,N_3141,N_3485);
nor U5272 (N_5272,N_2321,N_3666);
and U5273 (N_5273,N_2625,N_3353);
and U5274 (N_5274,N_2748,N_3723);
nand U5275 (N_5275,N_3962,N_3993);
xor U5276 (N_5276,N_3180,N_2522);
nor U5277 (N_5277,N_2143,N_2515);
and U5278 (N_5278,N_2163,N_2511);
and U5279 (N_5279,N_3369,N_2624);
nand U5280 (N_5280,N_3080,N_3234);
nand U5281 (N_5281,N_2176,N_3630);
nor U5282 (N_5282,N_2243,N_3438);
or U5283 (N_5283,N_2853,N_3503);
nor U5284 (N_5284,N_2903,N_3400);
or U5285 (N_5285,N_2472,N_2078);
or U5286 (N_5286,N_3586,N_2637);
xnor U5287 (N_5287,N_3378,N_2801);
xnor U5288 (N_5288,N_2258,N_3643);
or U5289 (N_5289,N_3011,N_3291);
nand U5290 (N_5290,N_2653,N_2725);
nand U5291 (N_5291,N_3691,N_2574);
nor U5292 (N_5292,N_3335,N_3149);
or U5293 (N_5293,N_2858,N_3860);
nor U5294 (N_5294,N_2327,N_3399);
xnor U5295 (N_5295,N_2618,N_2038);
or U5296 (N_5296,N_3949,N_3125);
or U5297 (N_5297,N_3954,N_2494);
xor U5298 (N_5298,N_2906,N_2938);
and U5299 (N_5299,N_3548,N_2094);
nand U5300 (N_5300,N_2666,N_3300);
xor U5301 (N_5301,N_3195,N_2527);
or U5302 (N_5302,N_2928,N_3174);
nor U5303 (N_5303,N_3546,N_3263);
and U5304 (N_5304,N_3885,N_2619);
nor U5305 (N_5305,N_3619,N_2549);
nand U5306 (N_5306,N_3332,N_2509);
nor U5307 (N_5307,N_2112,N_3569);
and U5308 (N_5308,N_3044,N_2668);
nand U5309 (N_5309,N_3612,N_2841);
or U5310 (N_5310,N_2215,N_3248);
and U5311 (N_5311,N_3383,N_3471);
nand U5312 (N_5312,N_3273,N_2352);
nor U5313 (N_5313,N_3441,N_3216);
nor U5314 (N_5314,N_2689,N_3606);
and U5315 (N_5315,N_2860,N_3256);
and U5316 (N_5316,N_3052,N_2915);
nand U5317 (N_5317,N_2661,N_2981);
or U5318 (N_5318,N_2267,N_2802);
and U5319 (N_5319,N_2922,N_2255);
nor U5320 (N_5320,N_2485,N_2731);
xor U5321 (N_5321,N_3525,N_2052);
nor U5322 (N_5322,N_2115,N_3280);
and U5323 (N_5323,N_3480,N_3248);
nand U5324 (N_5324,N_2426,N_3530);
nor U5325 (N_5325,N_3327,N_3945);
and U5326 (N_5326,N_2606,N_2211);
or U5327 (N_5327,N_3882,N_3807);
nand U5328 (N_5328,N_2247,N_3722);
or U5329 (N_5329,N_2027,N_3500);
or U5330 (N_5330,N_3305,N_2586);
or U5331 (N_5331,N_3287,N_2368);
nor U5332 (N_5332,N_3178,N_2831);
nor U5333 (N_5333,N_3417,N_2422);
or U5334 (N_5334,N_2171,N_3987);
nor U5335 (N_5335,N_2388,N_3099);
nand U5336 (N_5336,N_3080,N_2412);
and U5337 (N_5337,N_2924,N_3123);
and U5338 (N_5338,N_3543,N_3222);
or U5339 (N_5339,N_2209,N_3709);
nor U5340 (N_5340,N_2592,N_2314);
nor U5341 (N_5341,N_3619,N_3779);
and U5342 (N_5342,N_2536,N_2646);
and U5343 (N_5343,N_2526,N_2826);
nor U5344 (N_5344,N_3174,N_2001);
nand U5345 (N_5345,N_2882,N_2140);
nand U5346 (N_5346,N_3523,N_2937);
or U5347 (N_5347,N_3833,N_2941);
nor U5348 (N_5348,N_2549,N_2628);
nor U5349 (N_5349,N_2139,N_2294);
and U5350 (N_5350,N_2889,N_2350);
nand U5351 (N_5351,N_2571,N_2444);
xor U5352 (N_5352,N_2007,N_3927);
nand U5353 (N_5353,N_3633,N_3930);
nand U5354 (N_5354,N_3461,N_3570);
nand U5355 (N_5355,N_2913,N_2507);
and U5356 (N_5356,N_2938,N_2110);
nand U5357 (N_5357,N_3861,N_3858);
nand U5358 (N_5358,N_2987,N_3834);
or U5359 (N_5359,N_2429,N_3385);
or U5360 (N_5360,N_2857,N_2076);
and U5361 (N_5361,N_2459,N_3533);
nand U5362 (N_5362,N_3540,N_2599);
nand U5363 (N_5363,N_3236,N_3842);
and U5364 (N_5364,N_3547,N_3335);
nand U5365 (N_5365,N_2356,N_2128);
nor U5366 (N_5366,N_2234,N_3155);
or U5367 (N_5367,N_3465,N_3304);
or U5368 (N_5368,N_3989,N_2036);
or U5369 (N_5369,N_3576,N_2537);
nand U5370 (N_5370,N_3986,N_2575);
or U5371 (N_5371,N_3413,N_2654);
xnor U5372 (N_5372,N_2598,N_3158);
and U5373 (N_5373,N_3616,N_2444);
and U5374 (N_5374,N_3671,N_2892);
or U5375 (N_5375,N_3128,N_3351);
nand U5376 (N_5376,N_2421,N_3094);
nor U5377 (N_5377,N_3302,N_2983);
or U5378 (N_5378,N_2992,N_2261);
xor U5379 (N_5379,N_3066,N_3505);
or U5380 (N_5380,N_3031,N_2322);
xnor U5381 (N_5381,N_3909,N_3512);
or U5382 (N_5382,N_2854,N_2075);
nand U5383 (N_5383,N_2105,N_3728);
nand U5384 (N_5384,N_3104,N_2307);
nand U5385 (N_5385,N_2247,N_3515);
or U5386 (N_5386,N_2566,N_2886);
or U5387 (N_5387,N_2888,N_3306);
xnor U5388 (N_5388,N_3122,N_3726);
or U5389 (N_5389,N_2569,N_3433);
nor U5390 (N_5390,N_3565,N_3869);
or U5391 (N_5391,N_2276,N_3363);
nor U5392 (N_5392,N_2072,N_3109);
and U5393 (N_5393,N_2344,N_2196);
or U5394 (N_5394,N_3567,N_3027);
and U5395 (N_5395,N_2419,N_3296);
nor U5396 (N_5396,N_3112,N_3475);
nand U5397 (N_5397,N_3641,N_3589);
xnor U5398 (N_5398,N_3560,N_3243);
or U5399 (N_5399,N_3001,N_2721);
nand U5400 (N_5400,N_3786,N_3624);
and U5401 (N_5401,N_2841,N_2236);
xnor U5402 (N_5402,N_3933,N_2397);
or U5403 (N_5403,N_2645,N_2843);
and U5404 (N_5404,N_2631,N_3760);
nand U5405 (N_5405,N_2007,N_2182);
nand U5406 (N_5406,N_2194,N_2616);
nor U5407 (N_5407,N_3861,N_2203);
or U5408 (N_5408,N_3191,N_2863);
or U5409 (N_5409,N_2324,N_3858);
nor U5410 (N_5410,N_2944,N_3415);
xor U5411 (N_5411,N_2282,N_2618);
and U5412 (N_5412,N_2713,N_3169);
nor U5413 (N_5413,N_2118,N_2131);
nor U5414 (N_5414,N_3604,N_2388);
nor U5415 (N_5415,N_2902,N_3747);
xor U5416 (N_5416,N_2803,N_2189);
or U5417 (N_5417,N_2984,N_2020);
and U5418 (N_5418,N_2680,N_3593);
or U5419 (N_5419,N_3378,N_3544);
or U5420 (N_5420,N_3856,N_2675);
and U5421 (N_5421,N_2567,N_3427);
and U5422 (N_5422,N_2841,N_2949);
nand U5423 (N_5423,N_2220,N_2518);
and U5424 (N_5424,N_2995,N_3554);
nand U5425 (N_5425,N_3556,N_2642);
or U5426 (N_5426,N_2015,N_3518);
nor U5427 (N_5427,N_2562,N_3562);
xor U5428 (N_5428,N_2357,N_2467);
nor U5429 (N_5429,N_3235,N_3861);
nand U5430 (N_5430,N_2134,N_2351);
nand U5431 (N_5431,N_2731,N_3694);
or U5432 (N_5432,N_3020,N_2072);
nand U5433 (N_5433,N_2888,N_2085);
and U5434 (N_5434,N_3933,N_2793);
nor U5435 (N_5435,N_2833,N_2437);
nor U5436 (N_5436,N_3900,N_2944);
and U5437 (N_5437,N_3324,N_3824);
xnor U5438 (N_5438,N_3458,N_2910);
or U5439 (N_5439,N_2818,N_2493);
nand U5440 (N_5440,N_3160,N_3283);
or U5441 (N_5441,N_3112,N_3148);
or U5442 (N_5442,N_3454,N_2534);
and U5443 (N_5443,N_3676,N_2214);
nand U5444 (N_5444,N_3696,N_2910);
nand U5445 (N_5445,N_2541,N_3939);
nor U5446 (N_5446,N_3706,N_2751);
nor U5447 (N_5447,N_3349,N_3798);
and U5448 (N_5448,N_2429,N_3686);
and U5449 (N_5449,N_3948,N_3428);
or U5450 (N_5450,N_3454,N_2563);
nand U5451 (N_5451,N_3532,N_2916);
nor U5452 (N_5452,N_2086,N_3925);
or U5453 (N_5453,N_2113,N_3380);
or U5454 (N_5454,N_2284,N_2571);
nor U5455 (N_5455,N_2738,N_2185);
xnor U5456 (N_5456,N_2124,N_3699);
xor U5457 (N_5457,N_3421,N_3954);
or U5458 (N_5458,N_3310,N_3430);
nand U5459 (N_5459,N_2493,N_3139);
and U5460 (N_5460,N_2311,N_3998);
or U5461 (N_5461,N_2386,N_3937);
nor U5462 (N_5462,N_3764,N_2153);
and U5463 (N_5463,N_2936,N_2179);
nand U5464 (N_5464,N_3484,N_3950);
and U5465 (N_5465,N_3717,N_2301);
nand U5466 (N_5466,N_3569,N_2534);
and U5467 (N_5467,N_3668,N_2649);
nand U5468 (N_5468,N_3919,N_2822);
xnor U5469 (N_5469,N_3026,N_3238);
or U5470 (N_5470,N_2050,N_3326);
xnor U5471 (N_5471,N_3792,N_3134);
nand U5472 (N_5472,N_3444,N_3465);
nor U5473 (N_5473,N_3712,N_2862);
nand U5474 (N_5474,N_2567,N_2106);
nand U5475 (N_5475,N_3869,N_2494);
or U5476 (N_5476,N_3726,N_3871);
and U5477 (N_5477,N_3265,N_2802);
or U5478 (N_5478,N_2078,N_2925);
and U5479 (N_5479,N_3812,N_3413);
nor U5480 (N_5480,N_3773,N_3377);
nand U5481 (N_5481,N_2699,N_3660);
nand U5482 (N_5482,N_2013,N_2548);
nor U5483 (N_5483,N_3512,N_2528);
nand U5484 (N_5484,N_2207,N_3471);
nor U5485 (N_5485,N_3825,N_3761);
or U5486 (N_5486,N_3066,N_3069);
nor U5487 (N_5487,N_2561,N_3867);
or U5488 (N_5488,N_2653,N_3571);
nor U5489 (N_5489,N_3800,N_2636);
nand U5490 (N_5490,N_2712,N_2028);
and U5491 (N_5491,N_3658,N_3862);
nand U5492 (N_5492,N_2311,N_3352);
nand U5493 (N_5493,N_3460,N_2106);
or U5494 (N_5494,N_2669,N_2881);
or U5495 (N_5495,N_3907,N_2208);
and U5496 (N_5496,N_3159,N_2222);
or U5497 (N_5497,N_3107,N_3234);
nand U5498 (N_5498,N_3891,N_3871);
or U5499 (N_5499,N_3833,N_2820);
nor U5500 (N_5500,N_3523,N_3798);
nand U5501 (N_5501,N_2439,N_3322);
and U5502 (N_5502,N_3248,N_3622);
or U5503 (N_5503,N_2023,N_2620);
or U5504 (N_5504,N_3561,N_2895);
nor U5505 (N_5505,N_3465,N_2922);
and U5506 (N_5506,N_3737,N_3118);
nor U5507 (N_5507,N_3025,N_3107);
nand U5508 (N_5508,N_2578,N_3207);
xnor U5509 (N_5509,N_2933,N_2113);
nor U5510 (N_5510,N_3801,N_2420);
or U5511 (N_5511,N_2409,N_2048);
or U5512 (N_5512,N_2738,N_2389);
nor U5513 (N_5513,N_3237,N_3103);
or U5514 (N_5514,N_2862,N_2645);
or U5515 (N_5515,N_2659,N_2161);
or U5516 (N_5516,N_3476,N_3380);
nor U5517 (N_5517,N_2185,N_2971);
nand U5518 (N_5518,N_3556,N_3012);
nor U5519 (N_5519,N_2295,N_2999);
and U5520 (N_5520,N_3882,N_2953);
and U5521 (N_5521,N_3504,N_3909);
and U5522 (N_5522,N_3321,N_3126);
or U5523 (N_5523,N_3877,N_3855);
or U5524 (N_5524,N_2343,N_3584);
nor U5525 (N_5525,N_3066,N_3497);
and U5526 (N_5526,N_3575,N_2872);
nand U5527 (N_5527,N_2077,N_2688);
or U5528 (N_5528,N_2063,N_2148);
nor U5529 (N_5529,N_2261,N_3455);
or U5530 (N_5530,N_2594,N_3711);
nor U5531 (N_5531,N_3378,N_3078);
nor U5532 (N_5532,N_2107,N_2364);
or U5533 (N_5533,N_3847,N_2732);
xor U5534 (N_5534,N_2711,N_3966);
nand U5535 (N_5535,N_3386,N_3819);
and U5536 (N_5536,N_3223,N_2962);
xnor U5537 (N_5537,N_3763,N_3167);
nand U5538 (N_5538,N_2585,N_2786);
nand U5539 (N_5539,N_2661,N_3346);
nor U5540 (N_5540,N_2726,N_2228);
nand U5541 (N_5541,N_2915,N_2647);
or U5542 (N_5542,N_2471,N_2732);
xor U5543 (N_5543,N_3864,N_2596);
xor U5544 (N_5544,N_3382,N_2822);
nand U5545 (N_5545,N_3748,N_3897);
and U5546 (N_5546,N_2779,N_2737);
and U5547 (N_5547,N_3670,N_3027);
or U5548 (N_5548,N_3199,N_3131);
xor U5549 (N_5549,N_3271,N_2513);
or U5550 (N_5550,N_3231,N_2132);
or U5551 (N_5551,N_3552,N_2481);
nand U5552 (N_5552,N_2719,N_3752);
xnor U5553 (N_5553,N_2537,N_3529);
xnor U5554 (N_5554,N_2337,N_2877);
nand U5555 (N_5555,N_2900,N_2956);
nand U5556 (N_5556,N_3422,N_2975);
xor U5557 (N_5557,N_2442,N_2424);
and U5558 (N_5558,N_3280,N_3760);
or U5559 (N_5559,N_3494,N_3590);
nor U5560 (N_5560,N_3666,N_3192);
nor U5561 (N_5561,N_3018,N_2671);
xor U5562 (N_5562,N_2185,N_2803);
nor U5563 (N_5563,N_3426,N_2876);
and U5564 (N_5564,N_2170,N_2652);
nor U5565 (N_5565,N_2192,N_3873);
nand U5566 (N_5566,N_2127,N_3234);
and U5567 (N_5567,N_2915,N_3176);
xor U5568 (N_5568,N_3550,N_2895);
nor U5569 (N_5569,N_2657,N_2561);
nor U5570 (N_5570,N_2345,N_2872);
and U5571 (N_5571,N_3071,N_3518);
or U5572 (N_5572,N_3983,N_3221);
nand U5573 (N_5573,N_2497,N_3598);
nor U5574 (N_5574,N_2027,N_3140);
nand U5575 (N_5575,N_3071,N_3009);
nand U5576 (N_5576,N_2534,N_2827);
xor U5577 (N_5577,N_2617,N_2705);
nor U5578 (N_5578,N_3335,N_3072);
nor U5579 (N_5579,N_3180,N_3693);
or U5580 (N_5580,N_3152,N_3142);
nor U5581 (N_5581,N_2694,N_2506);
or U5582 (N_5582,N_3380,N_2132);
xnor U5583 (N_5583,N_2333,N_3237);
or U5584 (N_5584,N_2244,N_2584);
nand U5585 (N_5585,N_3429,N_2607);
nand U5586 (N_5586,N_3828,N_3015);
nor U5587 (N_5587,N_2031,N_3470);
nand U5588 (N_5588,N_3650,N_3703);
nor U5589 (N_5589,N_2337,N_2874);
or U5590 (N_5590,N_2722,N_3552);
nand U5591 (N_5591,N_3243,N_3848);
and U5592 (N_5592,N_2282,N_2390);
nand U5593 (N_5593,N_3439,N_2336);
or U5594 (N_5594,N_2607,N_2701);
xor U5595 (N_5595,N_3122,N_2738);
or U5596 (N_5596,N_2126,N_3397);
or U5597 (N_5597,N_3919,N_2030);
and U5598 (N_5598,N_2020,N_3625);
nand U5599 (N_5599,N_3182,N_3110);
and U5600 (N_5600,N_3048,N_2435);
nor U5601 (N_5601,N_2948,N_3337);
nand U5602 (N_5602,N_3303,N_2399);
xnor U5603 (N_5603,N_2503,N_3327);
and U5604 (N_5604,N_2491,N_2878);
and U5605 (N_5605,N_2967,N_2951);
nor U5606 (N_5606,N_3638,N_2099);
nor U5607 (N_5607,N_2545,N_3580);
nand U5608 (N_5608,N_3783,N_2328);
nor U5609 (N_5609,N_2785,N_3908);
nor U5610 (N_5610,N_2647,N_3158);
nor U5611 (N_5611,N_2995,N_3239);
or U5612 (N_5612,N_3650,N_2322);
xnor U5613 (N_5613,N_3389,N_3330);
or U5614 (N_5614,N_3531,N_3196);
or U5615 (N_5615,N_2621,N_2074);
and U5616 (N_5616,N_3267,N_3200);
and U5617 (N_5617,N_3158,N_3830);
nor U5618 (N_5618,N_3066,N_3855);
or U5619 (N_5619,N_3585,N_3908);
or U5620 (N_5620,N_3411,N_2619);
nor U5621 (N_5621,N_3221,N_2291);
or U5622 (N_5622,N_2697,N_3802);
or U5623 (N_5623,N_2280,N_3826);
and U5624 (N_5624,N_2840,N_3954);
nor U5625 (N_5625,N_3666,N_2917);
nand U5626 (N_5626,N_2494,N_3916);
nand U5627 (N_5627,N_3304,N_2733);
and U5628 (N_5628,N_2029,N_2645);
nor U5629 (N_5629,N_3571,N_3061);
nor U5630 (N_5630,N_2455,N_3777);
xnor U5631 (N_5631,N_2219,N_2523);
or U5632 (N_5632,N_2750,N_3579);
and U5633 (N_5633,N_3627,N_3163);
nand U5634 (N_5634,N_2798,N_2298);
nand U5635 (N_5635,N_3570,N_3614);
or U5636 (N_5636,N_3819,N_2752);
nor U5637 (N_5637,N_2825,N_3296);
nor U5638 (N_5638,N_3110,N_2613);
and U5639 (N_5639,N_2530,N_2588);
nor U5640 (N_5640,N_2706,N_3535);
nor U5641 (N_5641,N_3176,N_2261);
nand U5642 (N_5642,N_2559,N_3938);
and U5643 (N_5643,N_3671,N_2185);
and U5644 (N_5644,N_2550,N_3532);
and U5645 (N_5645,N_2093,N_3765);
nand U5646 (N_5646,N_3528,N_3382);
and U5647 (N_5647,N_3001,N_3538);
and U5648 (N_5648,N_3706,N_2689);
xnor U5649 (N_5649,N_2204,N_2072);
nor U5650 (N_5650,N_3216,N_3225);
nor U5651 (N_5651,N_2921,N_3439);
or U5652 (N_5652,N_2530,N_3075);
or U5653 (N_5653,N_3562,N_2886);
xor U5654 (N_5654,N_2734,N_3684);
nand U5655 (N_5655,N_2289,N_3409);
and U5656 (N_5656,N_2279,N_2130);
nor U5657 (N_5657,N_3065,N_2153);
or U5658 (N_5658,N_3148,N_3053);
nand U5659 (N_5659,N_3219,N_3249);
or U5660 (N_5660,N_3370,N_2296);
xnor U5661 (N_5661,N_3509,N_3699);
or U5662 (N_5662,N_2383,N_2697);
and U5663 (N_5663,N_2105,N_3131);
or U5664 (N_5664,N_2000,N_3019);
xnor U5665 (N_5665,N_3376,N_3950);
xor U5666 (N_5666,N_3654,N_3294);
nor U5667 (N_5667,N_2015,N_2569);
or U5668 (N_5668,N_3940,N_3953);
or U5669 (N_5669,N_3850,N_3935);
and U5670 (N_5670,N_3895,N_2323);
or U5671 (N_5671,N_2861,N_2426);
nor U5672 (N_5672,N_2352,N_3575);
and U5673 (N_5673,N_2498,N_2351);
nor U5674 (N_5674,N_3693,N_3635);
and U5675 (N_5675,N_3806,N_3172);
xnor U5676 (N_5676,N_2699,N_2405);
or U5677 (N_5677,N_2776,N_3558);
nand U5678 (N_5678,N_2629,N_2678);
nand U5679 (N_5679,N_2513,N_3208);
or U5680 (N_5680,N_2989,N_3018);
xor U5681 (N_5681,N_3524,N_3534);
and U5682 (N_5682,N_3439,N_3866);
nor U5683 (N_5683,N_2867,N_2791);
nor U5684 (N_5684,N_3065,N_3354);
nor U5685 (N_5685,N_3870,N_2340);
nand U5686 (N_5686,N_3712,N_3276);
and U5687 (N_5687,N_2893,N_2286);
and U5688 (N_5688,N_3315,N_2972);
or U5689 (N_5689,N_3019,N_2259);
xor U5690 (N_5690,N_2262,N_2346);
nand U5691 (N_5691,N_3747,N_3151);
nor U5692 (N_5692,N_2367,N_2807);
and U5693 (N_5693,N_2702,N_2192);
xnor U5694 (N_5694,N_2123,N_2795);
and U5695 (N_5695,N_3295,N_3019);
and U5696 (N_5696,N_3560,N_3895);
nand U5697 (N_5697,N_3688,N_3602);
nor U5698 (N_5698,N_3843,N_2428);
nand U5699 (N_5699,N_3010,N_3394);
and U5700 (N_5700,N_2128,N_3528);
nand U5701 (N_5701,N_2708,N_2497);
and U5702 (N_5702,N_3259,N_3639);
xor U5703 (N_5703,N_3888,N_2784);
and U5704 (N_5704,N_3431,N_3136);
nand U5705 (N_5705,N_3995,N_3543);
nand U5706 (N_5706,N_3039,N_2805);
nor U5707 (N_5707,N_3584,N_3236);
nor U5708 (N_5708,N_3454,N_2205);
and U5709 (N_5709,N_2616,N_2941);
nand U5710 (N_5710,N_2753,N_2545);
xor U5711 (N_5711,N_2652,N_2606);
nor U5712 (N_5712,N_2682,N_3568);
nor U5713 (N_5713,N_2281,N_2162);
or U5714 (N_5714,N_2589,N_3033);
nor U5715 (N_5715,N_3652,N_3876);
nand U5716 (N_5716,N_3122,N_3722);
nor U5717 (N_5717,N_3794,N_3761);
xnor U5718 (N_5718,N_2806,N_2227);
nor U5719 (N_5719,N_2007,N_2143);
or U5720 (N_5720,N_2900,N_3744);
nand U5721 (N_5721,N_3045,N_2277);
xor U5722 (N_5722,N_3213,N_2397);
and U5723 (N_5723,N_2182,N_2269);
and U5724 (N_5724,N_2551,N_3749);
and U5725 (N_5725,N_3532,N_3688);
and U5726 (N_5726,N_3147,N_3360);
and U5727 (N_5727,N_2976,N_2983);
nor U5728 (N_5728,N_3518,N_2351);
and U5729 (N_5729,N_3356,N_2157);
xnor U5730 (N_5730,N_3822,N_3721);
nand U5731 (N_5731,N_3930,N_2378);
nor U5732 (N_5732,N_3688,N_2929);
nor U5733 (N_5733,N_2616,N_3536);
xnor U5734 (N_5734,N_2466,N_2735);
or U5735 (N_5735,N_2723,N_2502);
nor U5736 (N_5736,N_3863,N_2716);
nor U5737 (N_5737,N_2837,N_2178);
nor U5738 (N_5738,N_2918,N_3255);
nor U5739 (N_5739,N_3902,N_2487);
nor U5740 (N_5740,N_3307,N_3923);
or U5741 (N_5741,N_3808,N_3668);
and U5742 (N_5742,N_3212,N_2455);
or U5743 (N_5743,N_3820,N_3912);
nand U5744 (N_5744,N_2225,N_3942);
nand U5745 (N_5745,N_3325,N_2688);
xnor U5746 (N_5746,N_2750,N_2506);
nor U5747 (N_5747,N_2636,N_3216);
and U5748 (N_5748,N_2279,N_3730);
nand U5749 (N_5749,N_2979,N_3271);
nor U5750 (N_5750,N_2924,N_2541);
and U5751 (N_5751,N_2952,N_2836);
or U5752 (N_5752,N_3635,N_3160);
or U5753 (N_5753,N_2389,N_2655);
and U5754 (N_5754,N_2198,N_3602);
nor U5755 (N_5755,N_2196,N_3936);
or U5756 (N_5756,N_2885,N_2918);
or U5757 (N_5757,N_3118,N_3912);
and U5758 (N_5758,N_2024,N_2552);
nor U5759 (N_5759,N_2406,N_2677);
nand U5760 (N_5760,N_3689,N_2801);
nand U5761 (N_5761,N_2520,N_2413);
and U5762 (N_5762,N_3882,N_3461);
and U5763 (N_5763,N_2421,N_3961);
and U5764 (N_5764,N_3089,N_3132);
nor U5765 (N_5765,N_3822,N_3602);
xnor U5766 (N_5766,N_2673,N_3436);
nor U5767 (N_5767,N_3871,N_2255);
and U5768 (N_5768,N_3237,N_2550);
and U5769 (N_5769,N_2130,N_3801);
nand U5770 (N_5770,N_2856,N_3095);
and U5771 (N_5771,N_2447,N_2805);
nand U5772 (N_5772,N_2952,N_2700);
nand U5773 (N_5773,N_2939,N_2897);
or U5774 (N_5774,N_3856,N_2826);
nand U5775 (N_5775,N_2934,N_2341);
and U5776 (N_5776,N_2077,N_2461);
or U5777 (N_5777,N_3001,N_2269);
or U5778 (N_5778,N_3483,N_3856);
and U5779 (N_5779,N_3309,N_2094);
and U5780 (N_5780,N_3548,N_2538);
or U5781 (N_5781,N_3104,N_3666);
xnor U5782 (N_5782,N_3072,N_2079);
and U5783 (N_5783,N_2174,N_2960);
or U5784 (N_5784,N_2946,N_3664);
nor U5785 (N_5785,N_3111,N_3115);
or U5786 (N_5786,N_3105,N_2076);
and U5787 (N_5787,N_3001,N_2838);
nor U5788 (N_5788,N_3218,N_3424);
and U5789 (N_5789,N_3699,N_3498);
or U5790 (N_5790,N_3832,N_2586);
or U5791 (N_5791,N_2749,N_2659);
or U5792 (N_5792,N_3209,N_2082);
xor U5793 (N_5793,N_2016,N_3465);
nand U5794 (N_5794,N_2447,N_2489);
and U5795 (N_5795,N_3929,N_3369);
nor U5796 (N_5796,N_2732,N_3784);
nand U5797 (N_5797,N_2410,N_2399);
or U5798 (N_5798,N_3269,N_3631);
xor U5799 (N_5799,N_3903,N_2003);
nand U5800 (N_5800,N_2483,N_2622);
or U5801 (N_5801,N_3403,N_2123);
nand U5802 (N_5802,N_2702,N_2133);
and U5803 (N_5803,N_2552,N_3412);
and U5804 (N_5804,N_3661,N_3900);
nand U5805 (N_5805,N_3632,N_2101);
or U5806 (N_5806,N_2588,N_3075);
or U5807 (N_5807,N_2735,N_2322);
or U5808 (N_5808,N_3850,N_2609);
or U5809 (N_5809,N_2019,N_3436);
xor U5810 (N_5810,N_2089,N_3107);
and U5811 (N_5811,N_3642,N_3482);
xor U5812 (N_5812,N_2477,N_3561);
or U5813 (N_5813,N_2778,N_2354);
xnor U5814 (N_5814,N_3937,N_2729);
nor U5815 (N_5815,N_3601,N_3282);
or U5816 (N_5816,N_2239,N_3820);
and U5817 (N_5817,N_3887,N_2046);
nand U5818 (N_5818,N_2376,N_3275);
and U5819 (N_5819,N_2979,N_2558);
nand U5820 (N_5820,N_3482,N_3569);
or U5821 (N_5821,N_2411,N_3560);
and U5822 (N_5822,N_3657,N_2289);
xnor U5823 (N_5823,N_3567,N_3242);
nand U5824 (N_5824,N_2391,N_3679);
nand U5825 (N_5825,N_2073,N_3474);
or U5826 (N_5826,N_2334,N_2897);
and U5827 (N_5827,N_2788,N_3002);
and U5828 (N_5828,N_3388,N_2464);
or U5829 (N_5829,N_2059,N_2008);
and U5830 (N_5830,N_3490,N_3530);
xnor U5831 (N_5831,N_2797,N_2021);
and U5832 (N_5832,N_2766,N_2253);
nor U5833 (N_5833,N_2535,N_2521);
and U5834 (N_5834,N_3835,N_2644);
nand U5835 (N_5835,N_2341,N_3852);
or U5836 (N_5836,N_3892,N_3180);
nor U5837 (N_5837,N_2296,N_3638);
nor U5838 (N_5838,N_2524,N_3440);
nor U5839 (N_5839,N_3677,N_2939);
nand U5840 (N_5840,N_3764,N_2293);
or U5841 (N_5841,N_2093,N_3875);
nand U5842 (N_5842,N_2578,N_3874);
and U5843 (N_5843,N_3967,N_3933);
xor U5844 (N_5844,N_3782,N_2181);
nand U5845 (N_5845,N_3317,N_3282);
or U5846 (N_5846,N_2889,N_2877);
nand U5847 (N_5847,N_2219,N_3501);
nand U5848 (N_5848,N_3201,N_2296);
or U5849 (N_5849,N_2430,N_2078);
or U5850 (N_5850,N_3036,N_2344);
nand U5851 (N_5851,N_3415,N_2202);
nor U5852 (N_5852,N_3591,N_2703);
and U5853 (N_5853,N_3774,N_3560);
xnor U5854 (N_5854,N_3708,N_2600);
xnor U5855 (N_5855,N_2314,N_2119);
xnor U5856 (N_5856,N_2273,N_3360);
nor U5857 (N_5857,N_3354,N_2059);
or U5858 (N_5858,N_3014,N_3133);
nand U5859 (N_5859,N_3514,N_3298);
or U5860 (N_5860,N_3215,N_2885);
and U5861 (N_5861,N_2634,N_2368);
nand U5862 (N_5862,N_3373,N_3262);
nor U5863 (N_5863,N_3314,N_2834);
and U5864 (N_5864,N_2894,N_3890);
or U5865 (N_5865,N_2360,N_2188);
xor U5866 (N_5866,N_3511,N_2620);
or U5867 (N_5867,N_2883,N_3863);
nor U5868 (N_5868,N_2699,N_3371);
nor U5869 (N_5869,N_2948,N_2987);
and U5870 (N_5870,N_2869,N_3768);
or U5871 (N_5871,N_3454,N_2564);
xor U5872 (N_5872,N_2350,N_2466);
or U5873 (N_5873,N_3603,N_2619);
nand U5874 (N_5874,N_2215,N_3501);
nor U5875 (N_5875,N_3059,N_3231);
nor U5876 (N_5876,N_2090,N_2046);
and U5877 (N_5877,N_3324,N_2354);
and U5878 (N_5878,N_3405,N_2305);
nand U5879 (N_5879,N_2678,N_2378);
and U5880 (N_5880,N_3213,N_3531);
xor U5881 (N_5881,N_2690,N_2270);
xor U5882 (N_5882,N_3769,N_2215);
nor U5883 (N_5883,N_3959,N_3800);
nand U5884 (N_5884,N_2599,N_2837);
and U5885 (N_5885,N_3994,N_3962);
nand U5886 (N_5886,N_2604,N_2147);
or U5887 (N_5887,N_2868,N_3981);
and U5888 (N_5888,N_2132,N_3028);
and U5889 (N_5889,N_2523,N_3454);
nor U5890 (N_5890,N_2251,N_3613);
and U5891 (N_5891,N_3826,N_3997);
nor U5892 (N_5892,N_3377,N_2869);
nand U5893 (N_5893,N_3119,N_3927);
nor U5894 (N_5894,N_2351,N_2370);
and U5895 (N_5895,N_2482,N_2836);
nand U5896 (N_5896,N_3810,N_2905);
nand U5897 (N_5897,N_2963,N_3502);
and U5898 (N_5898,N_3698,N_2327);
xor U5899 (N_5899,N_3828,N_2028);
nand U5900 (N_5900,N_3737,N_2601);
and U5901 (N_5901,N_2440,N_3456);
and U5902 (N_5902,N_2879,N_2544);
xor U5903 (N_5903,N_3428,N_2372);
and U5904 (N_5904,N_3811,N_2155);
and U5905 (N_5905,N_3983,N_2685);
nand U5906 (N_5906,N_2041,N_2125);
nor U5907 (N_5907,N_3710,N_3213);
nand U5908 (N_5908,N_3026,N_2808);
or U5909 (N_5909,N_2629,N_3915);
nand U5910 (N_5910,N_3749,N_2974);
nor U5911 (N_5911,N_3637,N_3428);
and U5912 (N_5912,N_3015,N_2140);
and U5913 (N_5913,N_2416,N_3138);
nand U5914 (N_5914,N_3031,N_3721);
or U5915 (N_5915,N_2592,N_3148);
or U5916 (N_5916,N_2985,N_2401);
or U5917 (N_5917,N_3804,N_3827);
nor U5918 (N_5918,N_2976,N_2595);
nor U5919 (N_5919,N_3998,N_2335);
or U5920 (N_5920,N_2279,N_2687);
nand U5921 (N_5921,N_3989,N_2426);
nor U5922 (N_5922,N_3394,N_3106);
or U5923 (N_5923,N_2578,N_2755);
or U5924 (N_5924,N_3902,N_3057);
and U5925 (N_5925,N_3155,N_2694);
xor U5926 (N_5926,N_3244,N_2849);
nor U5927 (N_5927,N_2960,N_3502);
nor U5928 (N_5928,N_3179,N_2503);
nand U5929 (N_5929,N_2821,N_3534);
or U5930 (N_5930,N_3702,N_2095);
nand U5931 (N_5931,N_3254,N_3348);
nand U5932 (N_5932,N_2112,N_3263);
xor U5933 (N_5933,N_3659,N_2033);
or U5934 (N_5934,N_2019,N_3115);
nor U5935 (N_5935,N_2976,N_3153);
and U5936 (N_5936,N_3056,N_2256);
xnor U5937 (N_5937,N_3037,N_3753);
nor U5938 (N_5938,N_3919,N_3756);
or U5939 (N_5939,N_3728,N_2700);
or U5940 (N_5940,N_3253,N_3195);
nand U5941 (N_5941,N_2463,N_2758);
xnor U5942 (N_5942,N_3987,N_2688);
nor U5943 (N_5943,N_2711,N_2251);
nand U5944 (N_5944,N_3445,N_3235);
nor U5945 (N_5945,N_2393,N_2274);
and U5946 (N_5946,N_2684,N_3196);
nand U5947 (N_5947,N_2663,N_2397);
or U5948 (N_5948,N_2644,N_3786);
nor U5949 (N_5949,N_2046,N_3040);
nor U5950 (N_5950,N_2646,N_3971);
nand U5951 (N_5951,N_2307,N_3368);
or U5952 (N_5952,N_2626,N_3736);
nor U5953 (N_5953,N_2836,N_2408);
xnor U5954 (N_5954,N_2773,N_3407);
nand U5955 (N_5955,N_3071,N_3174);
nor U5956 (N_5956,N_3415,N_2902);
or U5957 (N_5957,N_2408,N_3077);
or U5958 (N_5958,N_3235,N_3822);
nand U5959 (N_5959,N_2020,N_2668);
or U5960 (N_5960,N_2432,N_3518);
nand U5961 (N_5961,N_3668,N_2519);
xor U5962 (N_5962,N_2598,N_2630);
nand U5963 (N_5963,N_3344,N_2418);
nor U5964 (N_5964,N_3757,N_2777);
nand U5965 (N_5965,N_3486,N_3846);
xnor U5966 (N_5966,N_3480,N_2996);
nor U5967 (N_5967,N_2401,N_2784);
nand U5968 (N_5968,N_2257,N_3532);
and U5969 (N_5969,N_2848,N_3105);
nor U5970 (N_5970,N_3589,N_3401);
nand U5971 (N_5971,N_2753,N_3191);
or U5972 (N_5972,N_3727,N_2957);
or U5973 (N_5973,N_2297,N_2353);
nand U5974 (N_5974,N_3235,N_3042);
and U5975 (N_5975,N_3814,N_3399);
and U5976 (N_5976,N_2806,N_3942);
and U5977 (N_5977,N_2258,N_3221);
and U5978 (N_5978,N_2380,N_2852);
or U5979 (N_5979,N_2951,N_3571);
nand U5980 (N_5980,N_2957,N_2586);
nor U5981 (N_5981,N_3980,N_2362);
and U5982 (N_5982,N_3960,N_3076);
nand U5983 (N_5983,N_3862,N_2014);
and U5984 (N_5984,N_2516,N_3045);
and U5985 (N_5985,N_2054,N_3306);
nor U5986 (N_5986,N_3748,N_3785);
nor U5987 (N_5987,N_2219,N_2298);
nand U5988 (N_5988,N_3283,N_3542);
nand U5989 (N_5989,N_3837,N_2555);
nand U5990 (N_5990,N_2933,N_2907);
or U5991 (N_5991,N_2248,N_3269);
nor U5992 (N_5992,N_2696,N_2049);
xor U5993 (N_5993,N_3999,N_3683);
or U5994 (N_5994,N_3923,N_3002);
or U5995 (N_5995,N_3199,N_2660);
xnor U5996 (N_5996,N_3677,N_3480);
nand U5997 (N_5997,N_3316,N_3187);
or U5998 (N_5998,N_3825,N_3945);
and U5999 (N_5999,N_2650,N_2658);
and U6000 (N_6000,N_5379,N_5228);
nand U6001 (N_6001,N_5568,N_4970);
or U6002 (N_6002,N_4434,N_4689);
or U6003 (N_6003,N_5393,N_5767);
xnor U6004 (N_6004,N_4167,N_5240);
and U6005 (N_6005,N_4107,N_5171);
and U6006 (N_6006,N_4867,N_5942);
nand U6007 (N_6007,N_5303,N_4288);
and U6008 (N_6008,N_4808,N_5002);
and U6009 (N_6009,N_5217,N_5743);
nand U6010 (N_6010,N_4038,N_4232);
or U6011 (N_6011,N_5365,N_4761);
nand U6012 (N_6012,N_4591,N_5902);
and U6013 (N_6013,N_4893,N_4600);
nand U6014 (N_6014,N_4493,N_5052);
nor U6015 (N_6015,N_4848,N_4063);
nand U6016 (N_6016,N_5371,N_5138);
nor U6017 (N_6017,N_5233,N_4791);
and U6018 (N_6018,N_4877,N_5456);
and U6019 (N_6019,N_4148,N_4869);
and U6020 (N_6020,N_4551,N_4767);
nor U6021 (N_6021,N_5208,N_4269);
and U6022 (N_6022,N_5594,N_5358);
xnor U6023 (N_6023,N_4704,N_4996);
and U6024 (N_6024,N_5064,N_4678);
nor U6025 (N_6025,N_5739,N_5609);
or U6026 (N_6026,N_5253,N_4500);
nor U6027 (N_6027,N_4323,N_4881);
xor U6028 (N_6028,N_4222,N_4174);
xor U6029 (N_6029,N_5604,N_4283);
and U6030 (N_6030,N_5291,N_5910);
xor U6031 (N_6031,N_4208,N_5372);
nor U6032 (N_6032,N_5547,N_4006);
nand U6033 (N_6033,N_5298,N_4213);
and U6034 (N_6034,N_4637,N_4401);
or U6035 (N_6035,N_5949,N_4136);
nand U6036 (N_6036,N_5308,N_4954);
and U6037 (N_6037,N_4999,N_5343);
or U6038 (N_6038,N_5294,N_4099);
and U6039 (N_6039,N_5563,N_4062);
and U6040 (N_6040,N_5309,N_5092);
or U6041 (N_6041,N_4947,N_4571);
and U6042 (N_6042,N_5293,N_4168);
or U6043 (N_6043,N_5601,N_5356);
nand U6044 (N_6044,N_5473,N_4523);
xor U6045 (N_6045,N_5118,N_5627);
nor U6046 (N_6046,N_4366,N_4139);
and U6047 (N_6047,N_5225,N_5960);
nor U6048 (N_6048,N_5034,N_5694);
xnor U6049 (N_6049,N_5445,N_4393);
or U6050 (N_6050,N_4976,N_5194);
or U6051 (N_6051,N_5238,N_4708);
nand U6052 (N_6052,N_4741,N_4642);
xnor U6053 (N_6053,N_4550,N_4246);
nand U6054 (N_6054,N_4948,N_5053);
or U6055 (N_6055,N_4749,N_5311);
and U6056 (N_6056,N_4302,N_4952);
nand U6057 (N_6057,N_4077,N_5271);
or U6058 (N_6058,N_4928,N_4435);
xnor U6059 (N_6059,N_4601,N_5099);
and U6060 (N_6060,N_5079,N_5723);
nor U6061 (N_6061,N_5415,N_4456);
nor U6062 (N_6062,N_4982,N_5447);
nand U6063 (N_6063,N_5981,N_5510);
or U6064 (N_6064,N_5252,N_5660);
nor U6065 (N_6065,N_4409,N_4703);
or U6066 (N_6066,N_5448,N_5494);
nand U6067 (N_6067,N_4821,N_5847);
nor U6068 (N_6068,N_4919,N_5903);
nand U6069 (N_6069,N_5410,N_4781);
nand U6070 (N_6070,N_4610,N_5734);
or U6071 (N_6071,N_5121,N_4912);
nor U6072 (N_6072,N_5145,N_5350);
nor U6073 (N_6073,N_4487,N_5057);
and U6074 (N_6074,N_5459,N_4300);
nand U6075 (N_6075,N_4529,N_4587);
nand U6076 (N_6076,N_4513,N_5236);
or U6077 (N_6077,N_5526,N_4911);
or U6078 (N_6078,N_5501,N_5579);
xnor U6079 (N_6079,N_4763,N_5581);
and U6080 (N_6080,N_4901,N_5745);
and U6081 (N_6081,N_5668,N_5403);
nand U6082 (N_6082,N_4340,N_4764);
nand U6083 (N_6083,N_5747,N_4215);
xnor U6084 (N_6084,N_4843,N_5110);
nand U6085 (N_6085,N_5128,N_4756);
nand U6086 (N_6086,N_5848,N_5182);
nand U6087 (N_6087,N_4926,N_5474);
or U6088 (N_6088,N_5540,N_5724);
nor U6089 (N_6089,N_5658,N_4747);
xor U6090 (N_6090,N_4310,N_4719);
and U6091 (N_6091,N_4070,N_4701);
nand U6092 (N_6092,N_4913,N_4295);
nor U6093 (N_6093,N_5994,N_5490);
and U6094 (N_6094,N_4207,N_5257);
nand U6095 (N_6095,N_5987,N_5058);
nor U6096 (N_6096,N_4512,N_4992);
nand U6097 (N_6097,N_5261,N_4440);
or U6098 (N_6098,N_4790,N_5421);
xnor U6099 (N_6099,N_4639,N_5738);
nor U6100 (N_6100,N_4072,N_5499);
nor U6101 (N_6101,N_4073,N_4087);
or U6102 (N_6102,N_5504,N_4515);
and U6103 (N_6103,N_5400,N_5742);
and U6104 (N_6104,N_5210,N_4676);
or U6105 (N_6105,N_4120,N_4477);
or U6106 (N_6106,N_4622,N_4809);
nand U6107 (N_6107,N_5800,N_4303);
nor U6108 (N_6108,N_5882,N_5589);
nand U6109 (N_6109,N_5636,N_5032);
or U6110 (N_6110,N_5664,N_4503);
or U6111 (N_6111,N_5429,N_4617);
or U6112 (N_6112,N_5561,N_4542);
nand U6113 (N_6113,N_4615,N_5634);
nor U6114 (N_6114,N_5159,N_5527);
and U6115 (N_6115,N_4036,N_4424);
or U6116 (N_6116,N_5856,N_5564);
nand U6117 (N_6117,N_5854,N_5245);
nor U6118 (N_6118,N_5509,N_5783);
nand U6119 (N_6119,N_5885,N_5908);
nor U6120 (N_6120,N_4675,N_5255);
nor U6121 (N_6121,N_4548,N_4307);
and U6122 (N_6122,N_5152,N_4154);
nor U6123 (N_6123,N_5431,N_5251);
nor U6124 (N_6124,N_4290,N_4309);
nand U6125 (N_6125,N_5460,N_4430);
xnor U6126 (N_6126,N_5809,N_5321);
nand U6127 (N_6127,N_5711,N_4231);
nor U6128 (N_6128,N_5083,N_4325);
and U6129 (N_6129,N_4431,N_5899);
nand U6130 (N_6130,N_5316,N_5206);
nand U6131 (N_6131,N_5835,N_4308);
and U6132 (N_6132,N_4329,N_4349);
nor U6133 (N_6133,N_4203,N_4140);
xor U6134 (N_6134,N_4380,N_4720);
or U6135 (N_6135,N_4443,N_5129);
nor U6136 (N_6136,N_4552,N_4485);
nor U6137 (N_6137,N_5368,N_4138);
and U6138 (N_6138,N_5575,N_5176);
xnor U6139 (N_6139,N_4680,N_5939);
and U6140 (N_6140,N_5818,N_4454);
or U6141 (N_6141,N_5794,N_5907);
nand U6142 (N_6142,N_4988,N_4414);
xor U6143 (N_6143,N_5242,N_5435);
nor U6144 (N_6144,N_5823,N_5953);
nand U6145 (N_6145,N_5498,N_4359);
nand U6146 (N_6146,N_5131,N_5243);
nand U6147 (N_6147,N_5405,N_5966);
nor U6148 (N_6148,N_4461,N_4384);
and U6149 (N_6149,N_4182,N_5630);
and U6150 (N_6150,N_4093,N_4693);
and U6151 (N_6151,N_5962,N_5774);
nand U6152 (N_6152,N_5707,N_5808);
or U6153 (N_6153,N_5141,N_4449);
nand U6154 (N_6154,N_4827,N_4026);
nor U6155 (N_6155,N_5884,N_5496);
and U6156 (N_6156,N_4738,N_5156);
or U6157 (N_6157,N_4248,N_4267);
nor U6158 (N_6158,N_5227,N_4888);
or U6159 (N_6159,N_4626,N_5605);
nand U6160 (N_6160,N_4549,N_4711);
nand U6161 (N_6161,N_4007,N_5492);
nor U6162 (N_6162,N_5751,N_5729);
nand U6163 (N_6163,N_4373,N_5394);
xor U6164 (N_6164,N_5478,N_4623);
or U6165 (N_6165,N_4799,N_4990);
and U6166 (N_6166,N_4682,N_4371);
or U6167 (N_6167,N_5820,N_5952);
and U6168 (N_6168,N_4220,N_5346);
or U6169 (N_6169,N_5114,N_4031);
nor U6170 (N_6170,N_5262,N_4458);
nor U6171 (N_6171,N_5248,N_5682);
and U6172 (N_6172,N_5482,N_4321);
and U6173 (N_6173,N_4653,N_4949);
or U6174 (N_6174,N_5582,N_4211);
or U6175 (N_6175,N_5222,N_4488);
and U6176 (N_6176,N_4080,N_4352);
or U6177 (N_6177,N_4511,N_4603);
nor U6178 (N_6178,N_4852,N_4051);
xor U6179 (N_6179,N_5810,N_5554);
or U6180 (N_6180,N_5877,N_5263);
or U6181 (N_6181,N_4909,N_5637);
nor U6182 (N_6182,N_4934,N_4406);
and U6183 (N_6183,N_4097,N_5043);
nand U6184 (N_6184,N_5387,N_4668);
or U6185 (N_6185,N_5990,N_4645);
and U6186 (N_6186,N_5548,N_4650);
or U6187 (N_6187,N_5635,N_5135);
and U6188 (N_6188,N_5607,N_4876);
and U6189 (N_6189,N_4593,N_4452);
nor U6190 (N_6190,N_5891,N_5631);
and U6191 (N_6191,N_4611,N_5777);
or U6192 (N_6192,N_5659,N_5184);
nor U6193 (N_6193,N_4636,N_5934);
or U6194 (N_6194,N_4102,N_4633);
nand U6195 (N_6195,N_5537,N_5706);
and U6196 (N_6196,N_4491,N_4890);
or U6197 (N_6197,N_5111,N_5420);
and U6198 (N_6198,N_5798,N_5412);
and U6199 (N_6199,N_4906,N_4543);
nand U6200 (N_6200,N_5716,N_4684);
or U6201 (N_6201,N_5827,N_5109);
and U6202 (N_6202,N_4266,N_5229);
nor U6203 (N_6203,N_5805,N_5331);
or U6204 (N_6204,N_5599,N_4201);
xnor U6205 (N_6205,N_5784,N_5381);
or U6206 (N_6206,N_5787,N_5771);
nand U6207 (N_6207,N_4586,N_4698);
nand U6208 (N_6208,N_5922,N_4972);
and U6209 (N_6209,N_4795,N_4021);
nand U6210 (N_6210,N_5532,N_4433);
or U6211 (N_6211,N_4939,N_5106);
nand U6212 (N_6212,N_5825,N_4450);
nor U6213 (N_6213,N_5427,N_4173);
nand U6214 (N_6214,N_5649,N_4473);
or U6215 (N_6215,N_4058,N_4181);
and U6216 (N_6216,N_4836,N_4171);
or U6217 (N_6217,N_4332,N_4334);
and U6218 (N_6218,N_4740,N_5108);
and U6219 (N_6219,N_4779,N_4002);
and U6220 (N_6220,N_5201,N_5380);
nand U6221 (N_6221,N_5216,N_5434);
xnor U6222 (N_6222,N_5452,N_5895);
or U6223 (N_6223,N_4429,N_5082);
or U6224 (N_6224,N_5299,N_5187);
nor U6225 (N_6225,N_4152,N_5726);
xnor U6226 (N_6226,N_5041,N_4894);
nand U6227 (N_6227,N_5779,N_5849);
or U6228 (N_6228,N_5086,N_5397);
nand U6229 (N_6229,N_4100,N_5692);
or U6230 (N_6230,N_5918,N_5090);
nor U6231 (N_6231,N_4853,N_4261);
xor U6232 (N_6232,N_4640,N_5084);
nor U6233 (N_6233,N_5688,N_5551);
nor U6234 (N_6234,N_4572,N_4664);
nor U6235 (N_6235,N_5542,N_4963);
nor U6236 (N_6236,N_4158,N_4457);
nand U6237 (N_6237,N_5154,N_5234);
or U6238 (N_6238,N_5195,N_4936);
nor U6239 (N_6239,N_5807,N_4566);
nand U6240 (N_6240,N_5102,N_4262);
and U6241 (N_6241,N_5383,N_5833);
nand U6242 (N_6242,N_5753,N_5495);
or U6243 (N_6243,N_4306,N_4367);
nand U6244 (N_6244,N_5686,N_5022);
nor U6245 (N_6245,N_5440,N_4736);
nor U6246 (N_6246,N_5911,N_4824);
nand U6247 (N_6247,N_4277,N_4768);
nor U6248 (N_6248,N_5552,N_4797);
and U6249 (N_6249,N_5388,N_4276);
nor U6250 (N_6250,N_4737,N_4382);
or U6251 (N_6251,N_4157,N_5972);
nor U6252 (N_6252,N_4218,N_5016);
and U6253 (N_6253,N_4592,N_5602);
or U6254 (N_6254,N_4620,N_5756);
nand U6255 (N_6255,N_4599,N_4233);
nand U6256 (N_6256,N_5192,N_4563);
or U6257 (N_6257,N_4339,N_5158);
and U6258 (N_6258,N_4621,N_5212);
or U6259 (N_6259,N_4304,N_4442);
or U6260 (N_6260,N_4212,N_5180);
nor U6261 (N_6261,N_5676,N_4699);
nand U6262 (N_6262,N_5663,N_4933);
and U6263 (N_6263,N_4643,N_5219);
and U6264 (N_6264,N_5438,N_4391);
xor U6265 (N_6265,N_4921,N_4750);
xnor U6266 (N_6266,N_4722,N_5571);
or U6267 (N_6267,N_5488,N_5161);
and U6268 (N_6268,N_4607,N_5608);
nand U6269 (N_6269,N_4804,N_4345);
and U6270 (N_6270,N_4465,N_4818);
nand U6271 (N_6271,N_5035,N_5363);
nand U6272 (N_6272,N_4146,N_5348);
nand U6273 (N_6273,N_4811,N_4268);
nor U6274 (N_6274,N_4354,N_5355);
nand U6275 (N_6275,N_5009,N_5585);
or U6276 (N_6276,N_4180,N_5932);
nor U6277 (N_6277,N_4343,N_5703);
nand U6278 (N_6278,N_5773,N_4882);
nand U6279 (N_6279,N_5274,N_5731);
or U6280 (N_6280,N_4765,N_5978);
or U6281 (N_6281,N_4053,N_4368);
nand U6282 (N_6282,N_5324,N_4113);
xnor U6283 (N_6283,N_5570,N_5620);
or U6284 (N_6284,N_4064,N_5112);
or U6285 (N_6285,N_5375,N_5497);
or U6286 (N_6286,N_4855,N_4247);
and U6287 (N_6287,N_4376,N_5370);
nand U6288 (N_6288,N_5334,N_4445);
or U6289 (N_6289,N_4534,N_5572);
nand U6290 (N_6290,N_4028,N_4658);
and U6291 (N_6291,N_4482,N_5048);
nand U6292 (N_6292,N_5886,N_4553);
and U6293 (N_6293,N_5012,N_4423);
and U6294 (N_6294,N_5179,N_5287);
and U6295 (N_6295,N_4987,N_5300);
nand U6296 (N_6296,N_5183,N_4792);
and U6297 (N_6297,N_5615,N_4149);
nand U6298 (N_6298,N_5481,N_4287);
or U6299 (N_6299,N_4418,N_5669);
and U6300 (N_6300,N_5033,N_5469);
and U6301 (N_6301,N_4713,N_4715);
nand U6302 (N_6302,N_4669,N_4257);
or U6303 (N_6303,N_4386,N_5288);
or U6304 (N_6304,N_4472,N_5733);
nand U6305 (N_6305,N_4994,N_4880);
and U6306 (N_6306,N_4396,N_5975);
and U6307 (N_6307,N_4902,N_5980);
nand U6308 (N_6308,N_5887,N_4924);
xnor U6309 (N_6309,N_5611,N_4614);
nand U6310 (N_6310,N_4725,N_5999);
nand U6311 (N_6311,N_5565,N_5712);
xnor U6312 (N_6312,N_5720,N_5218);
or U6313 (N_6313,N_4151,N_5905);
and U6314 (N_6314,N_4015,N_5323);
or U6315 (N_6315,N_5275,N_5020);
and U6316 (N_6316,N_4962,N_5389);
nand U6317 (N_6317,N_5404,N_4665);
or U6318 (N_6318,N_5466,N_5970);
or U6319 (N_6319,N_4789,N_5428);
nor U6320 (N_6320,N_5741,N_4597);
nand U6321 (N_6321,N_5765,N_5095);
or U6322 (N_6322,N_5116,N_5764);
nand U6323 (N_6323,N_5367,N_5878);
nand U6324 (N_6324,N_5947,N_4466);
or U6325 (N_6325,N_5089,N_5120);
and U6326 (N_6326,N_4870,N_4872);
nand U6327 (N_6327,N_4499,N_5824);
and U6328 (N_6328,N_5622,N_4832);
nor U6329 (N_6329,N_4042,N_5595);
or U6330 (N_6330,N_5133,N_4925);
nor U6331 (N_6331,N_4350,N_4816);
nand U6332 (N_6332,N_5977,N_4706);
or U6333 (N_6333,N_5204,N_5858);
and U6334 (N_6334,N_4864,N_4039);
nor U6335 (N_6335,N_4469,N_5164);
or U6336 (N_6336,N_4094,N_4317);
or U6337 (N_6337,N_5104,N_5178);
or U6338 (N_6338,N_4337,N_4574);
nor U6339 (N_6339,N_4712,N_4776);
nor U6340 (N_6340,N_4125,N_4326);
and U6341 (N_6341,N_4116,N_5347);
and U6342 (N_6342,N_5819,N_4444);
or U6343 (N_6343,N_4083,N_5541);
nor U6344 (N_6344,N_5443,N_5312);
or U6345 (N_6345,N_4724,N_4132);
and U6346 (N_6346,N_4969,N_4065);
nand U6347 (N_6347,N_5401,N_5004);
or U6348 (N_6348,N_4530,N_4427);
and U6349 (N_6349,N_5470,N_4479);
nand U6350 (N_6350,N_4953,N_4109);
and U6351 (N_6351,N_5385,N_5047);
or U6352 (N_6352,N_5072,N_4686);
nand U6353 (N_6353,N_4106,N_4279);
nand U6354 (N_6354,N_5265,N_4375);
and U6355 (N_6355,N_4993,N_5979);
xnor U6356 (N_6356,N_5521,N_5283);
or U6357 (N_6357,N_4787,N_4786);
and U6358 (N_6358,N_5444,N_5744);
xnor U6359 (N_6359,N_5377,N_5361);
nand U6360 (N_6360,N_5603,N_5992);
xnor U6361 (N_6361,N_5569,N_5317);
or U6362 (N_6362,N_5476,N_5430);
or U6363 (N_6363,N_4090,N_5273);
xor U6364 (N_6364,N_4191,N_5066);
nor U6365 (N_6365,N_4470,N_5101);
and U6366 (N_6366,N_4944,N_4219);
and U6367 (N_6367,N_4716,N_4519);
nor U6368 (N_6368,N_5305,N_4481);
or U6369 (N_6369,N_5446,N_5454);
nand U6370 (N_6370,N_4942,N_5754);
or U6371 (N_6371,N_5489,N_4286);
or U6372 (N_6372,N_5797,N_5039);
nor U6373 (N_6373,N_5718,N_4648);
nand U6374 (N_6374,N_5221,N_5890);
nand U6375 (N_6375,N_4897,N_4961);
or U6376 (N_6376,N_5650,N_5418);
and U6377 (N_6377,N_5149,N_4502);
and U6378 (N_6378,N_4568,N_4946);
nand U6379 (N_6379,N_4577,N_4766);
nand U6380 (N_6380,N_4661,N_5702);
and U6381 (N_6381,N_5984,N_5717);
nand U6382 (N_6382,N_4825,N_5531);
nand U6383 (N_6383,N_5357,N_4504);
nor U6384 (N_6384,N_5632,N_5614);
nand U6385 (N_6385,N_4390,N_5677);
and U6386 (N_6386,N_4164,N_4865);
or U6387 (N_6387,N_4034,N_5130);
nand U6388 (N_6388,N_4627,N_5689);
or U6389 (N_6389,N_4751,N_5071);
or U6390 (N_6390,N_4258,N_5719);
nand U6391 (N_6391,N_5125,N_5924);
nand U6392 (N_6392,N_4474,N_4535);
or U6393 (N_6393,N_5730,N_4820);
or U6394 (N_6394,N_4092,N_4527);
nor U6395 (N_6395,N_5276,N_4830);
or U6396 (N_6396,N_4363,N_5748);
nand U6397 (N_6397,N_5736,N_4278);
nor U6398 (N_6398,N_4397,N_4197);
or U6399 (N_6399,N_5883,N_5487);
nand U6400 (N_6400,N_4108,N_4696);
or U6401 (N_6401,N_5591,N_4873);
and U6402 (N_6402,N_5577,N_5416);
nor U6403 (N_6403,N_5369,N_4404);
xor U6404 (N_6404,N_4398,N_4748);
nor U6405 (N_6405,N_5811,N_5266);
nand U6406 (N_6406,N_4141,N_4644);
nor U6407 (N_6407,N_4695,N_5480);
nand U6408 (N_6408,N_5529,N_4618);
nor U6409 (N_6409,N_5453,N_4837);
nor U6410 (N_6410,N_5518,N_5074);
and U6411 (N_6411,N_5969,N_4575);
nor U6412 (N_6412,N_4531,N_5354);
or U6413 (N_6413,N_5871,N_5044);
nor U6414 (N_6414,N_5536,N_5037);
and U6415 (N_6415,N_5770,N_4823);
nand U6416 (N_6416,N_4263,N_5055);
or U6417 (N_6417,N_5560,N_5107);
nand U6418 (N_6418,N_5423,N_5913);
nand U6419 (N_6419,N_4416,N_5640);
nor U6420 (N_6420,N_5338,N_4192);
nor U6421 (N_6421,N_4629,N_5307);
or U6422 (N_6422,N_4649,N_5535);
nor U6423 (N_6423,N_4459,N_5181);
or U6424 (N_6424,N_4646,N_5398);
and U6425 (N_6425,N_5003,N_5793);
and U6426 (N_6426,N_4803,N_4342);
nor U6427 (N_6427,N_5366,N_5322);
nand U6428 (N_6428,N_4112,N_5342);
and U6429 (N_6429,N_4845,N_4221);
nor U6430 (N_6430,N_5714,N_4495);
nand U6431 (N_6431,N_5061,N_5998);
nor U6432 (N_6432,N_4565,N_4679);
and U6433 (N_6433,N_4322,N_5610);
nor U6434 (N_6434,N_5633,N_5926);
or U6435 (N_6435,N_5834,N_5506);
xor U6436 (N_6436,N_5562,N_5938);
and U6437 (N_6437,N_5001,N_4255);
and U6438 (N_6438,N_5433,N_5127);
or U6439 (N_6439,N_4613,N_4560);
or U6440 (N_6440,N_5249,N_5458);
or U6441 (N_6441,N_5314,N_4358);
and U6442 (N_6442,N_5524,N_5687);
and U6443 (N_6443,N_4674,N_5968);
nand U6444 (N_6444,N_4585,N_5040);
and U6445 (N_6445,N_5619,N_4193);
or U6446 (N_6446,N_5483,N_4462);
and U6447 (N_6447,N_4123,N_5740);
nor U6448 (N_6448,N_5018,N_5573);
nand U6449 (N_6449,N_4273,N_5318);
nor U6450 (N_6450,N_5442,N_5936);
and U6451 (N_6451,N_5486,N_4372);
and U6452 (N_6452,N_4666,N_4777);
or U6453 (N_6453,N_4009,N_5378);
nand U6454 (N_6454,N_5162,N_4555);
nor U6455 (N_6455,N_4252,N_5502);
nor U6456 (N_6456,N_4150,N_5362);
nand U6457 (N_6457,N_4583,N_4717);
nand U6458 (N_6458,N_4041,N_5277);
and U6459 (N_6459,N_4866,N_4598);
or U6460 (N_6460,N_4985,N_4353);
or U6461 (N_6461,N_5831,N_4453);
nor U6462 (N_6462,N_4032,N_4705);
and U6463 (N_6463,N_5169,N_5073);
nor U6464 (N_6464,N_4179,N_5786);
or U6465 (N_6465,N_5737,N_4616);
and U6466 (N_6466,N_5235,N_4341);
nor U6467 (N_6467,N_4922,N_5203);
and U6468 (N_6468,N_4723,N_5320);
nand U6469 (N_6469,N_5749,N_5746);
and U6470 (N_6470,N_5762,N_4085);
nand U6471 (N_6471,N_4846,N_4033);
nand U6472 (N_6472,N_4995,N_4480);
or U6473 (N_6473,N_4984,N_5959);
and U6474 (N_6474,N_5451,N_5685);
nor U6475 (N_6475,N_5134,N_4849);
and U6476 (N_6476,N_5710,N_5479);
nand U6477 (N_6477,N_5008,N_4670);
and U6478 (N_6478,N_4189,N_4681);
or U6479 (N_6479,N_4851,N_4172);
nand U6480 (N_6480,N_5051,N_5559);
nor U6481 (N_6481,N_4710,N_5123);
nor U6482 (N_6482,N_5198,N_4205);
and U6483 (N_6483,N_5188,N_5643);
and U6484 (N_6484,N_4652,N_5259);
nand U6485 (N_6485,N_4812,N_4950);
and U6486 (N_6486,N_5103,N_5813);
and U6487 (N_6487,N_4918,N_4753);
and U6488 (N_6488,N_5491,N_5921);
or U6489 (N_6489,N_4111,N_5900);
nor U6490 (N_6490,N_4859,N_5792);
nor U6491 (N_6491,N_4000,N_4169);
nor U6492 (N_6492,N_4293,N_4402);
nor U6493 (N_6493,N_4735,N_4121);
nor U6494 (N_6494,N_4559,N_4506);
nor U6495 (N_6495,N_4634,N_4486);
nand U6496 (N_6496,N_4718,N_5097);
and U6497 (N_6497,N_5457,N_4244);
or U6498 (N_6498,N_4541,N_5645);
xnor U6499 (N_6499,N_5174,N_4428);
or U6500 (N_6500,N_5270,N_5826);
nand U6501 (N_6501,N_5391,N_5115);
or U6502 (N_6502,N_4929,N_5246);
nand U6503 (N_6503,N_4580,N_4436);
and U6504 (N_6504,N_4755,N_4128);
and U6505 (N_6505,N_5247,N_4426);
or U6506 (N_6506,N_4335,N_5530);
nand U6507 (N_6507,N_4476,N_5580);
xnor U6508 (N_6508,N_4573,N_5533);
and U6509 (N_6509,N_5988,N_4226);
nand U6510 (N_6510,N_4986,N_4594);
nand U6511 (N_6511,N_5596,N_4019);
nor U6512 (N_6512,N_5642,N_4324);
or U6513 (N_6513,N_4537,N_5864);
and U6514 (N_6514,N_4292,N_5485);
nand U6515 (N_6515,N_4916,N_5030);
nand U6516 (N_6516,N_4096,N_4004);
xor U6517 (N_6517,N_4732,N_4509);
nand U6518 (N_6518,N_5339,N_5750);
xor U6519 (N_6519,N_5782,N_5328);
and U6520 (N_6520,N_5177,N_5463);
nor U6521 (N_6521,N_4012,N_5075);
nor U6522 (N_6522,N_5861,N_4822);
nand U6523 (N_6523,N_5815,N_4259);
and U6524 (N_6524,N_5160,N_4828);
and U6525 (N_6525,N_4981,N_4539);
nor U6526 (N_6526,N_5091,N_5028);
nor U6527 (N_6527,N_5780,N_5665);
and U6528 (N_6528,N_4314,N_4561);
or U6529 (N_6529,N_5772,N_4819);
and U6530 (N_6530,N_4413,N_5105);
or U6531 (N_6531,N_4588,N_4410);
nand U6532 (N_6532,N_5725,N_4989);
nand U6533 (N_6533,N_4010,N_4241);
and U6534 (N_6534,N_4762,N_4657);
or U6535 (N_6535,N_5841,N_5172);
nor U6536 (N_6536,N_5407,N_5704);
xnor U6537 (N_6537,N_5758,N_5829);
or U6538 (N_6538,N_4250,N_4439);
or U6539 (N_6539,N_5344,N_5426);
nand U6540 (N_6540,N_4091,N_4299);
xor U6541 (N_6541,N_4931,N_5417);
nand U6542 (N_6542,N_5471,N_5029);
and U6543 (N_6543,N_4011,N_5189);
or U6544 (N_6544,N_5657,N_4842);
or U6545 (N_6545,N_5396,N_4806);
xor U6546 (N_6546,N_4518,N_5327);
nand U6547 (N_6547,N_4214,N_5140);
nor U6548 (N_6548,N_5837,N_4850);
nand U6549 (N_6549,N_4044,N_5644);
nand U6550 (N_6550,N_5545,N_4361);
or U6551 (N_6551,N_5011,N_4965);
nand U6552 (N_6552,N_4417,N_5906);
nand U6553 (N_6553,N_4857,N_5661);
nor U6554 (N_6554,N_5822,N_4907);
nor U6555 (N_6555,N_4496,N_4291);
nor U6556 (N_6556,N_4145,N_5759);
nor U6557 (N_6557,N_4043,N_4796);
and U6558 (N_6558,N_5695,N_5186);
and U6559 (N_6559,N_4392,N_5310);
and U6560 (N_6560,N_5000,N_4672);
nand U6561 (N_6561,N_4405,N_5424);
and U6562 (N_6562,N_4887,N_5892);
or U6563 (N_6563,N_5965,N_4813);
or U6564 (N_6564,N_5876,N_4862);
or U6565 (N_6565,N_5647,N_5543);
and U6566 (N_6566,N_5788,N_4878);
or U6567 (N_6567,N_4311,N_4810);
nor U6568 (N_6568,N_5576,N_4333);
nand U6569 (N_6569,N_4023,N_4389);
nand U6570 (N_6570,N_5666,N_5390);
and U6571 (N_6571,N_5296,N_4022);
nand U6572 (N_6572,N_5844,N_4115);
or U6573 (N_6573,N_5930,N_5943);
nor U6574 (N_6574,N_4892,N_4508);
and U6575 (N_6575,N_5117,N_5983);
xor U6576 (N_6576,N_5628,N_5302);
nor U6577 (N_6577,N_5042,N_4730);
or U6578 (N_6578,N_4379,N_5757);
or U6579 (N_6579,N_4794,N_4275);
or U6580 (N_6580,N_4369,N_4841);
and U6581 (N_6581,N_4697,N_5727);
and U6582 (N_6582,N_5013,N_4886);
or U6583 (N_6583,N_5673,N_5897);
nor U6584 (N_6584,N_4858,N_5098);
or U6585 (N_6585,N_4579,N_4831);
nor U6586 (N_6586,N_5113,N_4937);
or U6587 (N_6587,N_5191,N_5587);
nor U6588 (N_6588,N_4960,N_4505);
and U6589 (N_6589,N_5909,N_4294);
and U6590 (N_6590,N_4190,N_5295);
nand U6591 (N_6591,N_4175,N_5063);
and U6592 (N_6592,N_5364,N_5641);
nor U6593 (N_6593,N_4687,N_5708);
xnor U6594 (N_6594,N_4742,N_4833);
xor U6595 (N_6595,N_5578,N_5197);
and U6596 (N_6596,N_4223,N_4484);
and U6597 (N_6597,N_5699,N_4131);
nor U6598 (N_6598,N_5292,N_4957);
xor U6599 (N_6599,N_5985,N_5196);
nor U6600 (N_6600,N_4975,N_4251);
or U6601 (N_6601,N_5528,N_4069);
or U6602 (N_6602,N_4874,N_5795);
and U6603 (N_6603,N_5523,N_4076);
and U6604 (N_6604,N_5167,N_5336);
nand U6605 (N_6605,N_4973,N_4683);
nor U6606 (N_6606,N_5971,N_4497);
or U6607 (N_6607,N_5359,N_4526);
or U6608 (N_6608,N_4045,N_5679);
or U6609 (N_6609,N_5790,N_5144);
nand U6610 (N_6610,N_4501,N_4967);
and U6611 (N_6611,N_4758,N_4871);
or U6612 (N_6612,N_4312,N_4773);
nor U6613 (N_6613,N_4914,N_4050);
nor U6614 (N_6614,N_4854,N_4142);
or U6615 (N_6615,N_5828,N_5205);
and U6616 (N_6616,N_4264,N_5215);
or U6617 (N_6617,N_4119,N_4714);
nor U6618 (N_6618,N_5024,N_4159);
nor U6619 (N_6619,N_4979,N_5865);
nor U6620 (N_6620,N_5137,N_4861);
and U6621 (N_6621,N_4356,N_4020);
or U6622 (N_6622,N_4320,N_5917);
nor U6623 (N_6623,N_4447,N_4377);
or U6624 (N_6624,N_4057,N_4166);
xor U6625 (N_6625,N_4336,N_5625);
or U6626 (N_6626,N_5606,N_5955);
nand U6627 (N_6627,N_5873,N_4930);
or U6628 (N_6628,N_4927,N_4798);
and U6629 (N_6629,N_5213,N_4478);
nand U6630 (N_6630,N_5766,N_4037);
and U6631 (N_6631,N_5209,N_5132);
nor U6632 (N_6632,N_5651,N_5555);
or U6633 (N_6633,N_5735,N_5330);
or U6634 (N_6634,N_4071,N_5214);
nand U6635 (N_6635,N_5525,N_4253);
nor U6636 (N_6636,N_5850,N_5721);
nor U6637 (N_6637,N_5286,N_5335);
or U6638 (N_6638,N_4691,N_5341);
nor U6639 (N_6639,N_5549,N_4008);
or U6640 (N_6640,N_4517,N_5804);
or U6641 (N_6641,N_4143,N_4357);
nor U6642 (N_6642,N_5306,N_5190);
nor U6643 (N_6643,N_5211,N_5337);
and U6644 (N_6644,N_5049,N_5626);
and U6645 (N_6645,N_5076,N_4210);
nor U6646 (N_6646,N_5700,N_4688);
nand U6647 (N_6647,N_5006,N_4641);
nand U6648 (N_6648,N_5769,N_4826);
xnor U6649 (N_6649,N_5867,N_4360);
nor U6650 (N_6650,N_5840,N_5586);
xnor U6651 (N_6651,N_4860,N_4098);
or U6652 (N_6652,N_4200,N_4745);
or U6653 (N_6653,N_5094,N_5923);
nor U6654 (N_6654,N_5507,N_5613);
and U6655 (N_6655,N_5232,N_5974);
nor U6656 (N_6656,N_4018,N_4785);
or U6657 (N_6657,N_5653,N_5280);
nand U6658 (N_6658,N_4362,N_4743);
and U6659 (N_6659,N_5954,N_5230);
nand U6660 (N_6660,N_4204,N_4455);
or U6661 (N_6661,N_4217,N_5928);
and U6662 (N_6662,N_5546,N_5776);
nor U6663 (N_6663,N_4815,N_4524);
and U6664 (N_6664,N_4202,N_4977);
xor U6665 (N_6665,N_4104,N_4782);
and U6666 (N_6666,N_5279,N_5493);
nand U6667 (N_6667,N_4770,N_5851);
nor U6668 (N_6668,N_5508,N_5516);
nand U6669 (N_6669,N_4655,N_4702);
or U6670 (N_6670,N_5567,N_4619);
nand U6671 (N_6671,N_4562,N_5683);
nand U6672 (N_6672,N_4667,N_5200);
nand U6673 (N_6673,N_4692,N_5078);
or U6674 (N_6674,N_4467,N_4059);
xor U6675 (N_6675,N_4569,N_5450);
and U6676 (N_6676,N_4991,N_5461);
or U6677 (N_6677,N_4165,N_4029);
or U6678 (N_6678,N_5207,N_4974);
xor U6679 (N_6679,N_5406,N_4441);
xor U6680 (N_6680,N_4160,N_5693);
nand U6681 (N_6681,N_5588,N_4654);
and U6682 (N_6682,N_5254,N_5691);
and U6683 (N_6683,N_4422,N_5511);
or U6684 (N_6684,N_4908,N_5465);
or U6685 (N_6685,N_4879,N_5146);
nand U6686 (N_6686,N_5021,N_5901);
or U6687 (N_6687,N_4134,N_5888);
nand U6688 (N_6688,N_4707,N_5441);
nand U6689 (N_6689,N_4898,N_4003);
nand U6690 (N_6690,N_5284,N_5360);
and U6691 (N_6691,N_5832,N_4254);
and U6692 (N_6692,N_4608,N_5124);
nor U6693 (N_6693,N_5503,N_4726);
nor U6694 (N_6694,N_5945,N_5654);
or U6695 (N_6695,N_4318,N_5163);
and U6696 (N_6696,N_4086,N_5173);
or U6697 (N_6697,N_4101,N_5898);
nand U6698 (N_6698,N_5638,N_4133);
nor U6699 (N_6699,N_4105,N_4448);
nor U6700 (N_6700,N_5863,N_5333);
nand U6701 (N_6701,N_5297,N_4216);
nand U6702 (N_6702,N_4046,N_5713);
and U6703 (N_6703,N_5325,N_5268);
xor U6704 (N_6704,N_4068,N_4532);
nor U6705 (N_6705,N_5224,N_5056);
nor U6706 (N_6706,N_5920,N_4671);
and U6707 (N_6707,N_5881,N_4938);
nor U6708 (N_6708,N_5153,N_4895);
xnor U6709 (N_6709,N_4582,N_5799);
xor U6710 (N_6710,N_4547,N_5629);
and U6711 (N_6711,N_5472,N_4074);
nor U6712 (N_6712,N_5646,N_5019);
nor U6713 (N_6713,N_4540,N_5087);
or U6714 (N_6714,N_5862,N_4904);
or U6715 (N_6715,N_4209,N_4331);
nand U6716 (N_6716,N_5096,N_5648);
nand U6717 (N_6717,N_4186,N_4868);
and U6718 (N_6718,N_4196,N_4771);
and U6719 (N_6719,N_5267,N_4581);
and U6720 (N_6720,N_4365,N_5425);
nand U6721 (N_6721,N_5413,N_4606);
and U6722 (N_6722,N_5916,N_5329);
and U6723 (N_6723,N_5624,N_5872);
nand U6724 (N_6724,N_4829,N_4721);
or U6725 (N_6725,N_5550,N_4319);
and U6726 (N_6726,N_4178,N_4460);
or U6727 (N_6727,N_5467,N_4628);
nor U6728 (N_6728,N_5522,N_5373);
nor U6729 (N_6729,N_5986,N_4066);
nand U6730 (N_6730,N_4498,N_4659);
xor U6731 (N_6731,N_5148,N_4137);
xnor U6732 (N_6732,N_4399,N_5889);
nand U6733 (N_6733,N_4772,N_4387);
nor U6734 (N_6734,N_5411,N_4746);
nand U6735 (N_6735,N_5301,N_5995);
nor U6736 (N_6736,N_4917,N_5059);
nor U6737 (N_6737,N_5026,N_4395);
xor U6738 (N_6738,N_5583,N_4421);
and U6739 (N_6739,N_5991,N_5077);
or U6740 (N_6740,N_4514,N_4144);
nor U6741 (N_6741,N_4590,N_4631);
or U6742 (N_6742,N_4079,N_4147);
nor U6743 (N_6743,N_5946,N_4346);
nor U6744 (N_6744,N_5781,N_4225);
xnor U6745 (N_6745,N_5556,N_4049);
xor U6746 (N_6746,N_4759,N_4570);
and U6747 (N_6747,N_4437,N_4915);
nor U6748 (N_6748,N_5593,N_4662);
and U6749 (N_6749,N_4489,N_5399);
and U6750 (N_6750,N_4955,N_5763);
nand U6751 (N_6751,N_4844,N_4187);
and U6752 (N_6752,N_4733,N_5500);
or U6753 (N_6753,N_4891,N_5964);
and U6754 (N_6754,N_5853,N_4817);
nor U6755 (N_6755,N_5846,N_4016);
nor U6756 (N_6756,N_5119,N_5239);
nor U6757 (N_6757,N_4945,N_5590);
and U6758 (N_6758,N_4760,N_5600);
nand U6759 (N_6759,N_4793,N_5752);
or U6760 (N_6760,N_5806,N_5933);
or U6761 (N_6761,N_5031,N_4313);
nor U6762 (N_6762,N_4971,N_5623);
nand U6763 (N_6763,N_5812,N_5761);
or U6764 (N_6764,N_4538,N_4728);
nor U6765 (N_6765,N_5655,N_4612);
and U6766 (N_6766,N_5639,N_5870);
and U6767 (N_6767,N_4001,N_4556);
and U6768 (N_6768,N_4536,N_4305);
nor U6769 (N_6769,N_4638,N_5462);
or U6770 (N_6770,N_4463,N_4966);
or U6771 (N_6771,N_5919,N_5937);
nand U6772 (N_6772,N_4040,N_4875);
and U6773 (N_6773,N_4554,N_5732);
nand U6774 (N_6774,N_4920,N_4968);
and U6775 (N_6775,N_5353,N_5170);
nor U6776 (N_6776,N_5705,N_5760);
and U6777 (N_6777,N_4420,N_4814);
xor U6778 (N_6778,N_4412,N_4245);
nand U6779 (N_6779,N_5778,N_4774);
xor U6780 (N_6780,N_4896,N_4475);
nand U6781 (N_6781,N_4394,N_4905);
xnor U6782 (N_6782,N_4110,N_5538);
or U6783 (N_6783,N_4807,N_4381);
and U6784 (N_6784,N_4660,N_5621);
and U6785 (N_6785,N_4883,N_5285);
nor U6786 (N_6786,N_5802,N_5796);
and U6787 (N_6787,N_4625,N_4135);
xor U6788 (N_6788,N_5226,N_4176);
nand U6789 (N_6789,N_4052,N_4425);
and U6790 (N_6790,N_4240,N_5816);
nand U6791 (N_6791,N_4978,N_5068);
or U6792 (N_6792,N_5455,N_5351);
or U6793 (N_6793,N_4419,N_5845);
nand U6794 (N_6794,N_5231,N_5514);
nor U6795 (N_6795,N_4432,N_5392);
nand U6796 (N_6796,N_4297,N_5439);
and U6797 (N_6797,N_4510,N_4673);
or U6798 (N_6798,N_5142,N_4089);
nor U6799 (N_6799,N_5904,N_5290);
nor U6800 (N_6800,N_4647,N_5935);
nand U6801 (N_6801,N_4055,N_5278);
xor U6802 (N_6802,N_4769,N_5386);
or U6803 (N_6803,N_4082,N_4017);
and U6804 (N_6804,N_5422,N_4651);
and U6805 (N_6805,N_4483,N_4129);
nand U6806 (N_6806,N_5062,N_5505);
or U6807 (N_6807,N_5675,N_4964);
and U6808 (N_6808,N_4383,N_5715);
nor U6809 (N_6809,N_4236,N_4727);
nor U6810 (N_6810,N_5027,N_4492);
nor U6811 (N_6811,N_4075,N_5690);
nor U6812 (N_6812,N_4494,N_5519);
xnor U6813 (N_6813,N_4237,N_5951);
or U6814 (N_6814,N_4885,N_4910);
and U6815 (N_6815,N_5617,N_4471);
nor U6816 (N_6816,N_4084,N_5264);
nor U6817 (N_6817,N_5612,N_4940);
nor U6818 (N_6818,N_5941,N_4281);
or U6819 (N_6819,N_4838,N_5674);
and U6820 (N_6820,N_4576,N_5915);
or U6821 (N_6821,N_4163,N_4265);
or U6822 (N_6822,N_4403,N_5652);
and U6823 (N_6823,N_5319,N_5768);
and U6824 (N_6824,N_4124,N_5408);
xor U6825 (N_6825,N_5958,N_4184);
nand U6826 (N_6826,N_4752,N_5672);
nor U6827 (N_6827,N_4126,N_4558);
or U6828 (N_6828,N_5830,N_4282);
or U6829 (N_6829,N_5382,N_5963);
nand U6830 (N_6830,N_4378,N_4161);
or U6831 (N_6831,N_4155,N_5054);
nor U6832 (N_6832,N_5662,N_4663);
and U6833 (N_6833,N_5728,N_5374);
nor U6834 (N_6834,N_4694,N_5875);
nand U6835 (N_6835,N_5880,N_4239);
or U6836 (N_6836,N_4856,N_5857);
nand U6837 (N_6837,N_4932,N_5993);
and U6838 (N_6838,N_5484,N_5050);
xor U6839 (N_6839,N_5855,N_5223);
and U6840 (N_6840,N_5244,N_5409);
or U6841 (N_6841,N_5667,N_5574);
and U6842 (N_6842,N_4630,N_5976);
nand U6843 (N_6843,N_5513,N_5126);
or U6844 (N_6844,N_4374,N_5598);
or U6845 (N_6845,N_4557,N_5282);
or U6846 (N_6846,N_4959,N_5202);
nor U6847 (N_6847,N_4355,N_4081);
nor U6848 (N_6848,N_4700,N_4238);
nand U6849 (N_6849,N_5775,N_4602);
and U6850 (N_6850,N_5896,N_4400);
or U6851 (N_6851,N_5914,N_5956);
xor U6852 (N_6852,N_4054,N_4364);
nor U6853 (N_6853,N_5684,N_5067);
nand U6854 (N_6854,N_5477,N_4095);
nand U6855 (N_6855,N_4521,N_5241);
or U6856 (N_6856,N_5155,N_5045);
and U6857 (N_6857,N_5345,N_5996);
and U6858 (N_6858,N_5512,N_4162);
and U6859 (N_6859,N_4235,N_4889);
xor U6860 (N_6860,N_4185,N_5340);
or U6861 (N_6861,N_5534,N_4025);
nand U6862 (N_6862,N_4013,N_5616);
nand U6863 (N_6863,N_5384,N_4899);
nor U6864 (N_6864,N_4229,N_5803);
xnor U6865 (N_6865,N_5157,N_5566);
nand U6866 (N_6866,N_5289,N_5852);
or U6867 (N_6867,N_5940,N_4958);
nand U6868 (N_6868,N_4754,N_5866);
nand U6869 (N_6869,N_5879,N_5017);
nand U6870 (N_6870,N_4941,N_4884);
nor U6871 (N_6871,N_5927,N_5100);
nor U6872 (N_6872,N_4677,N_4271);
and U6873 (N_6873,N_4578,N_5395);
nand U6874 (N_6874,N_4243,N_5014);
and U6875 (N_6875,N_4328,N_4805);
nor U6876 (N_6876,N_4595,N_4014);
nand U6877 (N_6877,N_5814,N_5839);
xor U6878 (N_6878,N_4839,N_4330);
or U6879 (N_6879,N_4438,N_4533);
or U6880 (N_6880,N_4118,N_5950);
nor U6881 (N_6881,N_4520,N_5670);
and U6882 (N_6882,N_5237,N_4800);
and U6883 (N_6883,N_5326,N_5272);
or U6884 (N_6884,N_4775,N_4935);
nand U6885 (N_6885,N_5256,N_4951);
xnor U6886 (N_6886,N_4739,N_5982);
nor U6887 (N_6887,N_5136,N_5449);
or U6888 (N_6888,N_4451,N_5838);
xnor U6889 (N_6889,N_5698,N_4114);
nand U6890 (N_6890,N_4005,N_4998);
nor U6891 (N_6891,N_5869,N_5038);
and U6892 (N_6892,N_4546,N_4943);
and U6893 (N_6893,N_5260,N_4234);
or U6894 (N_6894,N_4117,N_5025);
nor U6895 (N_6895,N_5817,N_4411);
nand U6896 (N_6896,N_5122,N_4734);
and U6897 (N_6897,N_4801,N_4784);
or U6898 (N_6898,N_4122,N_4256);
and U6899 (N_6899,N_4272,N_5944);
and U6900 (N_6900,N_4316,N_5414);
nand U6901 (N_6901,N_5553,N_4249);
nor U6902 (N_6902,N_4298,N_4731);
nor U6903 (N_6903,N_4596,N_4047);
nand U6904 (N_6904,N_4060,N_4757);
and U6905 (N_6905,N_4840,N_5515);
and U6906 (N_6906,N_5558,N_4242);
or U6907 (N_6907,N_4315,N_5349);
and U6908 (N_6908,N_4834,N_4567);
nand U6909 (N_6909,N_5671,N_4528);
nand U6910 (N_6910,N_5315,N_5520);
nor U6911 (N_6911,N_4900,N_4327);
nand U6912 (N_6912,N_5168,N_5680);
nand U6913 (N_6913,N_4522,N_5060);
nor U6914 (N_6914,N_5093,N_5618);
or U6915 (N_6915,N_5801,N_4464);
or U6916 (N_6916,N_5836,N_4156);
nor U6917 (N_6917,N_5678,N_4690);
or U6918 (N_6918,N_5046,N_5656);
nor U6919 (N_6919,N_4301,N_4338);
nand U6920 (N_6920,N_5175,N_4835);
or U6921 (N_6921,N_5436,N_5894);
and U6922 (N_6922,N_4078,N_5036);
and U6923 (N_6923,N_5432,N_5007);
and U6924 (N_6924,N_5005,N_4183);
or U6925 (N_6925,N_4778,N_4656);
nand U6926 (N_6926,N_5250,N_4088);
or U6927 (N_6927,N_5258,N_4632);
nor U6928 (N_6928,N_4605,N_5821);
nand U6929 (N_6929,N_4127,N_5475);
or U6930 (N_6930,N_4685,N_5859);
and U6931 (N_6931,N_5165,N_4609);
and U6932 (N_6932,N_4544,N_4035);
and U6933 (N_6933,N_4507,N_4385);
or U6934 (N_6934,N_5544,N_5468);
nand U6935 (N_6935,N_5313,N_5143);
or U6936 (N_6936,N_5464,N_4198);
and U6937 (N_6937,N_4285,N_4370);
and U6938 (N_6938,N_4344,N_4997);
xnor U6939 (N_6939,N_5332,N_5893);
nand U6940 (N_6940,N_5304,N_5791);
nor U6941 (N_6941,N_5069,N_4516);
nor U6942 (N_6942,N_5957,N_5070);
or U6943 (N_6943,N_4188,N_4103);
or U6944 (N_6944,N_4260,N_5419);
and U6945 (N_6945,N_4130,N_5402);
and U6946 (N_6946,N_4709,N_5085);
nand U6947 (N_6947,N_4199,N_4289);
nand U6948 (N_6948,N_4415,N_5755);
or U6949 (N_6949,N_4783,N_5789);
and U6950 (N_6950,N_5842,N_4230);
nand U6951 (N_6951,N_5929,N_5925);
nor U6952 (N_6952,N_4351,N_4194);
nor U6953 (N_6953,N_5592,N_4923);
or U6954 (N_6954,N_4048,N_5584);
nand U6955 (N_6955,N_5080,N_5709);
and U6956 (N_6956,N_5722,N_4956);
xnor U6957 (N_6957,N_4206,N_4274);
or U6958 (N_6958,N_4227,N_5912);
nand U6959 (N_6959,N_5860,N_5681);
nor U6960 (N_6960,N_5065,N_4635);
nand U6961 (N_6961,N_5185,N_5697);
and U6962 (N_6962,N_4564,N_5023);
nor U6963 (N_6963,N_5269,N_5701);
and U6964 (N_6964,N_5220,N_4863);
nor U6965 (N_6965,N_4195,N_4788);
xnor U6966 (N_6966,N_4027,N_5843);
and U6967 (N_6967,N_4348,N_4407);
nor U6968 (N_6968,N_4847,N_4980);
and U6969 (N_6969,N_5010,N_5437);
xor U6970 (N_6970,N_5517,N_4624);
nand U6971 (N_6971,N_5193,N_4228);
xnor U6972 (N_6972,N_4903,N_4525);
and U6973 (N_6973,N_4584,N_5015);
and U6974 (N_6974,N_4177,N_5967);
nand U6975 (N_6975,N_5597,N_4030);
and U6976 (N_6976,N_4983,N_4468);
or U6977 (N_6977,N_4729,N_4280);
xor U6978 (N_6978,N_4604,N_5376);
xor U6979 (N_6979,N_5081,N_5539);
nor U6980 (N_6980,N_4744,N_4224);
nor U6981 (N_6981,N_5874,N_5147);
and U6982 (N_6982,N_5139,N_5199);
nor U6983 (N_6983,N_5931,N_4284);
or U6984 (N_6984,N_5352,N_4589);
nand U6985 (N_6985,N_5150,N_5989);
or U6986 (N_6986,N_4446,N_4490);
nor U6987 (N_6987,N_4067,N_5696);
nand U6988 (N_6988,N_5088,N_4296);
nor U6989 (N_6989,N_5281,N_4170);
nor U6990 (N_6990,N_4270,N_4408);
nand U6991 (N_6991,N_5973,N_5997);
and U6992 (N_6992,N_4780,N_4545);
and U6993 (N_6993,N_4024,N_5151);
and U6994 (N_6994,N_4153,N_4388);
nor U6995 (N_6995,N_5557,N_5948);
and U6996 (N_6996,N_5166,N_4347);
xnor U6997 (N_6997,N_5961,N_5868);
nor U6998 (N_6998,N_5785,N_4056);
or U6999 (N_6999,N_4802,N_4061);
nand U7000 (N_7000,N_4209,N_4868);
xor U7001 (N_7001,N_5852,N_5660);
xnor U7002 (N_7002,N_5220,N_5075);
nand U7003 (N_7003,N_4537,N_4261);
and U7004 (N_7004,N_5337,N_5233);
or U7005 (N_7005,N_4493,N_5382);
or U7006 (N_7006,N_5679,N_4516);
xor U7007 (N_7007,N_4810,N_5300);
and U7008 (N_7008,N_5198,N_5622);
nor U7009 (N_7009,N_4935,N_4139);
xnor U7010 (N_7010,N_4231,N_5440);
and U7011 (N_7011,N_4489,N_5339);
and U7012 (N_7012,N_4003,N_4466);
or U7013 (N_7013,N_5205,N_4760);
nand U7014 (N_7014,N_4632,N_5667);
nor U7015 (N_7015,N_5509,N_5042);
and U7016 (N_7016,N_4667,N_4349);
nor U7017 (N_7017,N_4277,N_5815);
nand U7018 (N_7018,N_4279,N_5932);
or U7019 (N_7019,N_5733,N_4367);
and U7020 (N_7020,N_5457,N_4714);
nand U7021 (N_7021,N_4632,N_4854);
nor U7022 (N_7022,N_4976,N_5276);
or U7023 (N_7023,N_5452,N_5422);
nand U7024 (N_7024,N_4505,N_4791);
and U7025 (N_7025,N_4805,N_5674);
nor U7026 (N_7026,N_4272,N_4434);
nand U7027 (N_7027,N_5889,N_4618);
and U7028 (N_7028,N_4702,N_4129);
or U7029 (N_7029,N_5282,N_4371);
xor U7030 (N_7030,N_4147,N_5866);
nand U7031 (N_7031,N_4307,N_4926);
and U7032 (N_7032,N_5974,N_4240);
and U7033 (N_7033,N_4407,N_5716);
nor U7034 (N_7034,N_4222,N_4676);
nand U7035 (N_7035,N_4721,N_4966);
and U7036 (N_7036,N_4342,N_5699);
nor U7037 (N_7037,N_5437,N_5003);
xor U7038 (N_7038,N_4551,N_4002);
and U7039 (N_7039,N_4635,N_5794);
nor U7040 (N_7040,N_4397,N_5111);
nor U7041 (N_7041,N_4959,N_4969);
nand U7042 (N_7042,N_4253,N_5609);
nand U7043 (N_7043,N_5935,N_5949);
nor U7044 (N_7044,N_5154,N_5075);
xnor U7045 (N_7045,N_4663,N_5311);
nand U7046 (N_7046,N_5792,N_5691);
nand U7047 (N_7047,N_5228,N_5767);
or U7048 (N_7048,N_4276,N_4283);
or U7049 (N_7049,N_4423,N_5921);
and U7050 (N_7050,N_4749,N_5498);
nor U7051 (N_7051,N_5003,N_5264);
or U7052 (N_7052,N_4197,N_4432);
nor U7053 (N_7053,N_5520,N_5818);
nand U7054 (N_7054,N_5314,N_5626);
or U7055 (N_7055,N_4270,N_4741);
and U7056 (N_7056,N_4896,N_4232);
nor U7057 (N_7057,N_5941,N_4830);
xor U7058 (N_7058,N_4382,N_4107);
nor U7059 (N_7059,N_4317,N_5851);
nand U7060 (N_7060,N_4767,N_5286);
or U7061 (N_7061,N_4955,N_5812);
and U7062 (N_7062,N_5613,N_5081);
and U7063 (N_7063,N_5914,N_4626);
or U7064 (N_7064,N_4746,N_4835);
or U7065 (N_7065,N_4958,N_4178);
xnor U7066 (N_7066,N_4112,N_5013);
and U7067 (N_7067,N_4773,N_5601);
and U7068 (N_7068,N_4345,N_5828);
nor U7069 (N_7069,N_5315,N_5473);
and U7070 (N_7070,N_5129,N_5372);
nand U7071 (N_7071,N_5876,N_4520);
and U7072 (N_7072,N_4569,N_4801);
nor U7073 (N_7073,N_5587,N_4374);
xor U7074 (N_7074,N_4389,N_4133);
or U7075 (N_7075,N_4275,N_4143);
nand U7076 (N_7076,N_5314,N_4958);
nor U7077 (N_7077,N_5047,N_4032);
or U7078 (N_7078,N_4254,N_5952);
nand U7079 (N_7079,N_4132,N_4409);
or U7080 (N_7080,N_5636,N_4104);
nand U7081 (N_7081,N_4363,N_5125);
nor U7082 (N_7082,N_4377,N_5576);
xor U7083 (N_7083,N_4098,N_4740);
nor U7084 (N_7084,N_5224,N_5138);
nand U7085 (N_7085,N_5025,N_5647);
xnor U7086 (N_7086,N_5385,N_4284);
and U7087 (N_7087,N_5272,N_5709);
nand U7088 (N_7088,N_5485,N_4867);
and U7089 (N_7089,N_4530,N_5774);
nand U7090 (N_7090,N_5926,N_4152);
nor U7091 (N_7091,N_4123,N_4202);
and U7092 (N_7092,N_4718,N_4005);
nor U7093 (N_7093,N_5589,N_4769);
nand U7094 (N_7094,N_4796,N_4874);
or U7095 (N_7095,N_5758,N_5198);
nand U7096 (N_7096,N_4761,N_4466);
xnor U7097 (N_7097,N_4423,N_4648);
nor U7098 (N_7098,N_4328,N_5388);
nor U7099 (N_7099,N_4326,N_4386);
nand U7100 (N_7100,N_4998,N_4540);
nor U7101 (N_7101,N_5683,N_5050);
and U7102 (N_7102,N_5519,N_5437);
nand U7103 (N_7103,N_5230,N_5248);
or U7104 (N_7104,N_4238,N_4114);
nand U7105 (N_7105,N_4240,N_5753);
and U7106 (N_7106,N_4079,N_5877);
nor U7107 (N_7107,N_5494,N_5112);
nor U7108 (N_7108,N_4943,N_4079);
nand U7109 (N_7109,N_4923,N_5256);
nand U7110 (N_7110,N_5420,N_4148);
or U7111 (N_7111,N_4840,N_5758);
nor U7112 (N_7112,N_4433,N_4397);
nor U7113 (N_7113,N_5658,N_5792);
and U7114 (N_7114,N_4590,N_5389);
or U7115 (N_7115,N_5354,N_5762);
and U7116 (N_7116,N_4148,N_5519);
or U7117 (N_7117,N_5165,N_4676);
nor U7118 (N_7118,N_4695,N_5251);
or U7119 (N_7119,N_4249,N_4378);
and U7120 (N_7120,N_5058,N_4790);
or U7121 (N_7121,N_4677,N_4418);
nor U7122 (N_7122,N_4151,N_4995);
nand U7123 (N_7123,N_4354,N_4099);
or U7124 (N_7124,N_4852,N_4656);
nand U7125 (N_7125,N_5566,N_5894);
nand U7126 (N_7126,N_4064,N_5544);
nor U7127 (N_7127,N_5182,N_5411);
nor U7128 (N_7128,N_4493,N_4017);
or U7129 (N_7129,N_5573,N_4697);
and U7130 (N_7130,N_4103,N_4075);
or U7131 (N_7131,N_5082,N_5767);
or U7132 (N_7132,N_4944,N_5098);
nor U7133 (N_7133,N_5991,N_5402);
or U7134 (N_7134,N_5498,N_5126);
xnor U7135 (N_7135,N_5924,N_5762);
nand U7136 (N_7136,N_5048,N_5301);
or U7137 (N_7137,N_4453,N_4707);
nand U7138 (N_7138,N_4364,N_4636);
nand U7139 (N_7139,N_4960,N_5390);
and U7140 (N_7140,N_5498,N_5307);
xnor U7141 (N_7141,N_5643,N_5926);
and U7142 (N_7142,N_5562,N_5698);
and U7143 (N_7143,N_4688,N_4624);
nor U7144 (N_7144,N_5404,N_5736);
nand U7145 (N_7145,N_5033,N_5555);
and U7146 (N_7146,N_4704,N_4636);
nor U7147 (N_7147,N_4605,N_4053);
and U7148 (N_7148,N_5293,N_4886);
xnor U7149 (N_7149,N_4483,N_4645);
nor U7150 (N_7150,N_4628,N_4623);
nand U7151 (N_7151,N_4752,N_4621);
and U7152 (N_7152,N_4043,N_4025);
nand U7153 (N_7153,N_5890,N_4776);
nor U7154 (N_7154,N_5333,N_4468);
or U7155 (N_7155,N_5834,N_4569);
nand U7156 (N_7156,N_5742,N_4297);
xnor U7157 (N_7157,N_5395,N_5055);
or U7158 (N_7158,N_4353,N_5339);
xnor U7159 (N_7159,N_5237,N_4536);
nor U7160 (N_7160,N_4273,N_4376);
nand U7161 (N_7161,N_5500,N_4066);
and U7162 (N_7162,N_5311,N_4176);
nor U7163 (N_7163,N_4645,N_4157);
xnor U7164 (N_7164,N_4307,N_4837);
nor U7165 (N_7165,N_4971,N_5289);
nand U7166 (N_7166,N_5845,N_4452);
nand U7167 (N_7167,N_5828,N_4074);
nor U7168 (N_7168,N_5857,N_5652);
nor U7169 (N_7169,N_4811,N_4761);
and U7170 (N_7170,N_5359,N_4600);
and U7171 (N_7171,N_4093,N_4004);
or U7172 (N_7172,N_4907,N_5982);
nor U7173 (N_7173,N_4196,N_4397);
nand U7174 (N_7174,N_4405,N_5661);
and U7175 (N_7175,N_4088,N_5738);
or U7176 (N_7176,N_5177,N_5644);
and U7177 (N_7177,N_5022,N_5007);
nand U7178 (N_7178,N_4431,N_4650);
xor U7179 (N_7179,N_5147,N_4322);
and U7180 (N_7180,N_4051,N_4842);
xor U7181 (N_7181,N_5410,N_5082);
or U7182 (N_7182,N_5362,N_4691);
nor U7183 (N_7183,N_4069,N_4858);
or U7184 (N_7184,N_5096,N_4522);
or U7185 (N_7185,N_4902,N_5835);
or U7186 (N_7186,N_5968,N_4460);
nor U7187 (N_7187,N_4255,N_4613);
nor U7188 (N_7188,N_5287,N_4926);
and U7189 (N_7189,N_4176,N_5277);
xnor U7190 (N_7190,N_4642,N_5247);
or U7191 (N_7191,N_5678,N_5863);
nor U7192 (N_7192,N_5778,N_5515);
or U7193 (N_7193,N_4213,N_4286);
and U7194 (N_7194,N_4502,N_4756);
xnor U7195 (N_7195,N_4382,N_4541);
xor U7196 (N_7196,N_5998,N_5572);
nand U7197 (N_7197,N_4256,N_4942);
nor U7198 (N_7198,N_4701,N_5930);
nand U7199 (N_7199,N_4796,N_5331);
and U7200 (N_7200,N_4610,N_4062);
nand U7201 (N_7201,N_5245,N_5442);
or U7202 (N_7202,N_4113,N_5567);
or U7203 (N_7203,N_4476,N_5715);
nand U7204 (N_7204,N_4755,N_4763);
or U7205 (N_7205,N_5546,N_5881);
nand U7206 (N_7206,N_4843,N_5023);
and U7207 (N_7207,N_5442,N_5737);
nand U7208 (N_7208,N_4137,N_5427);
and U7209 (N_7209,N_5071,N_5927);
nor U7210 (N_7210,N_5503,N_4992);
or U7211 (N_7211,N_4302,N_4503);
nand U7212 (N_7212,N_4853,N_4809);
and U7213 (N_7213,N_4558,N_5664);
nand U7214 (N_7214,N_4369,N_4809);
and U7215 (N_7215,N_5008,N_5270);
nand U7216 (N_7216,N_5362,N_4529);
or U7217 (N_7217,N_4465,N_4788);
and U7218 (N_7218,N_5833,N_5205);
nand U7219 (N_7219,N_5694,N_4850);
and U7220 (N_7220,N_5166,N_4616);
nor U7221 (N_7221,N_4941,N_5537);
nand U7222 (N_7222,N_4327,N_4220);
and U7223 (N_7223,N_5451,N_5697);
and U7224 (N_7224,N_5869,N_4969);
or U7225 (N_7225,N_4789,N_5115);
or U7226 (N_7226,N_4365,N_4141);
nor U7227 (N_7227,N_5065,N_5928);
and U7228 (N_7228,N_5136,N_5166);
xnor U7229 (N_7229,N_5835,N_5364);
nand U7230 (N_7230,N_5576,N_5629);
nor U7231 (N_7231,N_4946,N_5907);
xnor U7232 (N_7232,N_5837,N_4778);
or U7233 (N_7233,N_5060,N_4682);
or U7234 (N_7234,N_5824,N_4646);
and U7235 (N_7235,N_5459,N_5888);
nand U7236 (N_7236,N_4305,N_4155);
nor U7237 (N_7237,N_4349,N_5900);
or U7238 (N_7238,N_4415,N_4458);
xnor U7239 (N_7239,N_5197,N_5670);
and U7240 (N_7240,N_4442,N_5952);
xor U7241 (N_7241,N_5252,N_4544);
nand U7242 (N_7242,N_4052,N_5057);
or U7243 (N_7243,N_4092,N_5346);
nor U7244 (N_7244,N_4428,N_4943);
nor U7245 (N_7245,N_5786,N_5830);
nor U7246 (N_7246,N_5963,N_5977);
and U7247 (N_7247,N_5352,N_4500);
nor U7248 (N_7248,N_5291,N_4304);
nor U7249 (N_7249,N_4143,N_5147);
and U7250 (N_7250,N_4939,N_4259);
and U7251 (N_7251,N_5509,N_4664);
or U7252 (N_7252,N_5377,N_5035);
nand U7253 (N_7253,N_5919,N_5377);
or U7254 (N_7254,N_4910,N_5809);
nor U7255 (N_7255,N_5802,N_5067);
nand U7256 (N_7256,N_5365,N_4183);
or U7257 (N_7257,N_5105,N_5050);
and U7258 (N_7258,N_4668,N_5197);
or U7259 (N_7259,N_4085,N_4618);
and U7260 (N_7260,N_4364,N_4824);
or U7261 (N_7261,N_5576,N_4960);
or U7262 (N_7262,N_5510,N_5232);
nand U7263 (N_7263,N_5396,N_4315);
nand U7264 (N_7264,N_5009,N_5711);
and U7265 (N_7265,N_4307,N_5787);
nand U7266 (N_7266,N_5680,N_4691);
nor U7267 (N_7267,N_4308,N_5944);
xnor U7268 (N_7268,N_5334,N_4336);
xnor U7269 (N_7269,N_4989,N_4979);
or U7270 (N_7270,N_4595,N_5238);
nand U7271 (N_7271,N_5246,N_5911);
and U7272 (N_7272,N_4316,N_4666);
nor U7273 (N_7273,N_4365,N_4049);
nor U7274 (N_7274,N_4103,N_4171);
and U7275 (N_7275,N_5360,N_5630);
and U7276 (N_7276,N_5888,N_5255);
and U7277 (N_7277,N_5362,N_4047);
or U7278 (N_7278,N_4896,N_4329);
and U7279 (N_7279,N_5944,N_5091);
nor U7280 (N_7280,N_5154,N_5903);
xnor U7281 (N_7281,N_4248,N_5331);
xnor U7282 (N_7282,N_4458,N_5395);
nand U7283 (N_7283,N_5613,N_4564);
xnor U7284 (N_7284,N_5655,N_4198);
or U7285 (N_7285,N_5892,N_5174);
or U7286 (N_7286,N_5812,N_4548);
nand U7287 (N_7287,N_5756,N_5973);
or U7288 (N_7288,N_4154,N_4727);
nand U7289 (N_7289,N_4349,N_5036);
nand U7290 (N_7290,N_4745,N_4273);
and U7291 (N_7291,N_4703,N_4250);
nor U7292 (N_7292,N_4784,N_4284);
and U7293 (N_7293,N_5836,N_4761);
and U7294 (N_7294,N_4471,N_4763);
and U7295 (N_7295,N_4292,N_4879);
nor U7296 (N_7296,N_5920,N_5968);
or U7297 (N_7297,N_4268,N_5228);
and U7298 (N_7298,N_4593,N_5046);
or U7299 (N_7299,N_4590,N_5823);
or U7300 (N_7300,N_4043,N_5291);
nand U7301 (N_7301,N_4693,N_5229);
nor U7302 (N_7302,N_5108,N_5142);
nor U7303 (N_7303,N_4999,N_4593);
nor U7304 (N_7304,N_4292,N_4101);
or U7305 (N_7305,N_5795,N_5953);
nor U7306 (N_7306,N_4305,N_5421);
nor U7307 (N_7307,N_5567,N_5435);
and U7308 (N_7308,N_5615,N_5210);
or U7309 (N_7309,N_4505,N_5894);
nand U7310 (N_7310,N_5901,N_4840);
or U7311 (N_7311,N_5206,N_5551);
or U7312 (N_7312,N_5932,N_5437);
nor U7313 (N_7313,N_5550,N_5429);
nand U7314 (N_7314,N_5148,N_5223);
nor U7315 (N_7315,N_4121,N_4065);
or U7316 (N_7316,N_5839,N_5401);
nand U7317 (N_7317,N_4475,N_5971);
and U7318 (N_7318,N_5282,N_5805);
or U7319 (N_7319,N_5457,N_4609);
nand U7320 (N_7320,N_5451,N_5012);
xor U7321 (N_7321,N_5223,N_4275);
xor U7322 (N_7322,N_4770,N_4278);
xor U7323 (N_7323,N_4852,N_4469);
and U7324 (N_7324,N_4259,N_4172);
nand U7325 (N_7325,N_5365,N_5541);
nand U7326 (N_7326,N_5284,N_4548);
nor U7327 (N_7327,N_4273,N_5035);
and U7328 (N_7328,N_4498,N_4078);
nand U7329 (N_7329,N_5659,N_4052);
xor U7330 (N_7330,N_5970,N_4925);
nor U7331 (N_7331,N_5349,N_5031);
or U7332 (N_7332,N_4745,N_4525);
xor U7333 (N_7333,N_5857,N_5203);
or U7334 (N_7334,N_4907,N_5364);
nand U7335 (N_7335,N_4451,N_5862);
or U7336 (N_7336,N_4359,N_4227);
or U7337 (N_7337,N_5496,N_5419);
or U7338 (N_7338,N_5557,N_4326);
and U7339 (N_7339,N_5183,N_4127);
nor U7340 (N_7340,N_5881,N_5242);
and U7341 (N_7341,N_4364,N_4757);
or U7342 (N_7342,N_4341,N_5513);
or U7343 (N_7343,N_5021,N_4771);
or U7344 (N_7344,N_4996,N_5100);
nor U7345 (N_7345,N_5952,N_4489);
and U7346 (N_7346,N_5781,N_5130);
nor U7347 (N_7347,N_4801,N_5196);
nand U7348 (N_7348,N_4866,N_4349);
xor U7349 (N_7349,N_5913,N_4844);
xor U7350 (N_7350,N_5588,N_4384);
and U7351 (N_7351,N_4344,N_5499);
and U7352 (N_7352,N_4912,N_4245);
and U7353 (N_7353,N_4115,N_5640);
nand U7354 (N_7354,N_5344,N_5084);
xor U7355 (N_7355,N_4733,N_4214);
and U7356 (N_7356,N_4928,N_5250);
nor U7357 (N_7357,N_5363,N_4977);
or U7358 (N_7358,N_5689,N_4866);
nand U7359 (N_7359,N_4283,N_4404);
nor U7360 (N_7360,N_5066,N_5184);
nand U7361 (N_7361,N_4608,N_5104);
nand U7362 (N_7362,N_5815,N_5588);
and U7363 (N_7363,N_5901,N_5000);
nand U7364 (N_7364,N_4085,N_4760);
or U7365 (N_7365,N_5324,N_5087);
nand U7366 (N_7366,N_4649,N_4826);
xor U7367 (N_7367,N_4106,N_4118);
or U7368 (N_7368,N_5920,N_5284);
xor U7369 (N_7369,N_4195,N_5899);
or U7370 (N_7370,N_4307,N_4903);
nor U7371 (N_7371,N_5920,N_4586);
nor U7372 (N_7372,N_4228,N_5370);
or U7373 (N_7373,N_5875,N_5587);
nand U7374 (N_7374,N_4671,N_5410);
nand U7375 (N_7375,N_4754,N_5496);
nor U7376 (N_7376,N_5902,N_4011);
nand U7377 (N_7377,N_5737,N_4002);
nand U7378 (N_7378,N_5631,N_5001);
nor U7379 (N_7379,N_5006,N_5547);
nand U7380 (N_7380,N_4991,N_5089);
nand U7381 (N_7381,N_5353,N_5358);
and U7382 (N_7382,N_5048,N_4264);
nor U7383 (N_7383,N_4816,N_4811);
nand U7384 (N_7384,N_4969,N_5953);
nand U7385 (N_7385,N_5361,N_4472);
nand U7386 (N_7386,N_4968,N_5332);
nor U7387 (N_7387,N_4158,N_4277);
nor U7388 (N_7388,N_4086,N_4088);
nand U7389 (N_7389,N_4638,N_5764);
or U7390 (N_7390,N_4092,N_5103);
nor U7391 (N_7391,N_5757,N_4608);
nand U7392 (N_7392,N_4896,N_5571);
and U7393 (N_7393,N_5885,N_4368);
nand U7394 (N_7394,N_4572,N_4741);
or U7395 (N_7395,N_5117,N_5725);
nand U7396 (N_7396,N_4566,N_5052);
xor U7397 (N_7397,N_4620,N_4969);
nand U7398 (N_7398,N_4831,N_5791);
and U7399 (N_7399,N_4019,N_4924);
nor U7400 (N_7400,N_4099,N_4695);
nor U7401 (N_7401,N_4493,N_4175);
or U7402 (N_7402,N_5352,N_4592);
nor U7403 (N_7403,N_4154,N_5211);
nor U7404 (N_7404,N_4116,N_4489);
and U7405 (N_7405,N_4075,N_5471);
nor U7406 (N_7406,N_5424,N_5457);
and U7407 (N_7407,N_5857,N_4970);
or U7408 (N_7408,N_5963,N_5338);
and U7409 (N_7409,N_4831,N_4617);
xnor U7410 (N_7410,N_5067,N_4848);
nand U7411 (N_7411,N_5792,N_4690);
or U7412 (N_7412,N_4865,N_4885);
or U7413 (N_7413,N_4184,N_4077);
and U7414 (N_7414,N_4236,N_4800);
nand U7415 (N_7415,N_5691,N_4475);
or U7416 (N_7416,N_4607,N_5003);
nand U7417 (N_7417,N_4510,N_4726);
or U7418 (N_7418,N_5184,N_4684);
xnor U7419 (N_7419,N_4376,N_5353);
and U7420 (N_7420,N_5631,N_5444);
and U7421 (N_7421,N_5944,N_4106);
and U7422 (N_7422,N_5815,N_4661);
or U7423 (N_7423,N_5127,N_5391);
nand U7424 (N_7424,N_5609,N_4193);
nor U7425 (N_7425,N_5880,N_4515);
nor U7426 (N_7426,N_5649,N_4315);
and U7427 (N_7427,N_5006,N_5420);
nand U7428 (N_7428,N_4412,N_5383);
or U7429 (N_7429,N_4651,N_4014);
and U7430 (N_7430,N_4845,N_4496);
and U7431 (N_7431,N_4512,N_4483);
nor U7432 (N_7432,N_4731,N_4039);
or U7433 (N_7433,N_4115,N_4616);
nor U7434 (N_7434,N_5226,N_4267);
nor U7435 (N_7435,N_4304,N_4102);
nand U7436 (N_7436,N_5715,N_4272);
and U7437 (N_7437,N_4116,N_5473);
xnor U7438 (N_7438,N_5575,N_4901);
or U7439 (N_7439,N_5063,N_4231);
nor U7440 (N_7440,N_4968,N_5234);
or U7441 (N_7441,N_4132,N_5341);
nand U7442 (N_7442,N_4690,N_4886);
nor U7443 (N_7443,N_4041,N_5517);
nor U7444 (N_7444,N_4605,N_5645);
and U7445 (N_7445,N_5392,N_5578);
nand U7446 (N_7446,N_5671,N_4306);
nor U7447 (N_7447,N_5284,N_4975);
nand U7448 (N_7448,N_4387,N_5642);
nor U7449 (N_7449,N_4073,N_5708);
or U7450 (N_7450,N_5186,N_4029);
and U7451 (N_7451,N_5484,N_4425);
and U7452 (N_7452,N_4756,N_4250);
or U7453 (N_7453,N_5372,N_5808);
or U7454 (N_7454,N_5319,N_4898);
and U7455 (N_7455,N_5235,N_5716);
nand U7456 (N_7456,N_4615,N_5785);
and U7457 (N_7457,N_5195,N_4210);
and U7458 (N_7458,N_4648,N_4800);
xor U7459 (N_7459,N_4700,N_4375);
xor U7460 (N_7460,N_5205,N_5467);
nand U7461 (N_7461,N_4489,N_5453);
and U7462 (N_7462,N_5423,N_5507);
nand U7463 (N_7463,N_5753,N_5555);
and U7464 (N_7464,N_4175,N_5423);
nand U7465 (N_7465,N_4140,N_4281);
nor U7466 (N_7466,N_4556,N_5318);
and U7467 (N_7467,N_5238,N_5543);
or U7468 (N_7468,N_5719,N_5218);
nor U7469 (N_7469,N_4303,N_4551);
and U7470 (N_7470,N_5482,N_4152);
nand U7471 (N_7471,N_4575,N_4628);
and U7472 (N_7472,N_4750,N_5908);
nand U7473 (N_7473,N_4891,N_5521);
nor U7474 (N_7474,N_5476,N_4153);
and U7475 (N_7475,N_5495,N_4898);
and U7476 (N_7476,N_5861,N_4566);
or U7477 (N_7477,N_5042,N_4708);
or U7478 (N_7478,N_4660,N_5234);
and U7479 (N_7479,N_5586,N_4768);
nor U7480 (N_7480,N_5271,N_5327);
and U7481 (N_7481,N_4153,N_4969);
nor U7482 (N_7482,N_4325,N_4343);
nand U7483 (N_7483,N_5114,N_5218);
xnor U7484 (N_7484,N_4041,N_5266);
or U7485 (N_7485,N_4157,N_5130);
or U7486 (N_7486,N_5625,N_5307);
nor U7487 (N_7487,N_5605,N_4661);
or U7488 (N_7488,N_5331,N_4708);
nand U7489 (N_7489,N_4480,N_5226);
and U7490 (N_7490,N_5900,N_5694);
nor U7491 (N_7491,N_4728,N_4600);
nand U7492 (N_7492,N_4787,N_4863);
or U7493 (N_7493,N_5493,N_5457);
nor U7494 (N_7494,N_4890,N_4116);
xnor U7495 (N_7495,N_5849,N_4161);
nor U7496 (N_7496,N_5062,N_4693);
nor U7497 (N_7497,N_4343,N_4486);
nand U7498 (N_7498,N_4945,N_4509);
and U7499 (N_7499,N_4558,N_5714);
nand U7500 (N_7500,N_4781,N_4951);
nand U7501 (N_7501,N_5096,N_4076);
nand U7502 (N_7502,N_5038,N_5039);
and U7503 (N_7503,N_5256,N_5212);
and U7504 (N_7504,N_5339,N_4784);
nand U7505 (N_7505,N_5977,N_4347);
nor U7506 (N_7506,N_4536,N_5425);
or U7507 (N_7507,N_4653,N_5346);
and U7508 (N_7508,N_5813,N_4510);
xor U7509 (N_7509,N_4627,N_5404);
or U7510 (N_7510,N_4060,N_4658);
and U7511 (N_7511,N_5033,N_5636);
and U7512 (N_7512,N_5853,N_4934);
nand U7513 (N_7513,N_4506,N_5562);
or U7514 (N_7514,N_5340,N_5091);
or U7515 (N_7515,N_4533,N_5648);
or U7516 (N_7516,N_5438,N_4677);
or U7517 (N_7517,N_4636,N_4791);
or U7518 (N_7518,N_5504,N_5389);
and U7519 (N_7519,N_5342,N_4947);
xor U7520 (N_7520,N_5466,N_4574);
or U7521 (N_7521,N_4435,N_4766);
xnor U7522 (N_7522,N_4064,N_4361);
nand U7523 (N_7523,N_4702,N_4126);
xor U7524 (N_7524,N_5715,N_5963);
or U7525 (N_7525,N_5387,N_5710);
nor U7526 (N_7526,N_4581,N_4894);
or U7527 (N_7527,N_5846,N_4311);
nand U7528 (N_7528,N_5249,N_4058);
and U7529 (N_7529,N_5701,N_5774);
and U7530 (N_7530,N_4406,N_4488);
or U7531 (N_7531,N_4290,N_4682);
nand U7532 (N_7532,N_4628,N_4081);
and U7533 (N_7533,N_4413,N_4572);
xor U7534 (N_7534,N_4093,N_5458);
nor U7535 (N_7535,N_5677,N_5250);
or U7536 (N_7536,N_4130,N_5720);
and U7537 (N_7537,N_5565,N_4217);
nand U7538 (N_7538,N_4103,N_5592);
or U7539 (N_7539,N_4048,N_4547);
nand U7540 (N_7540,N_4482,N_5227);
or U7541 (N_7541,N_4630,N_5748);
or U7542 (N_7542,N_4605,N_5902);
nand U7543 (N_7543,N_5222,N_5070);
and U7544 (N_7544,N_4078,N_4440);
nor U7545 (N_7545,N_4007,N_5081);
nor U7546 (N_7546,N_5572,N_4403);
nor U7547 (N_7547,N_4301,N_5807);
nor U7548 (N_7548,N_5220,N_5699);
or U7549 (N_7549,N_4048,N_4272);
or U7550 (N_7550,N_5175,N_5289);
xor U7551 (N_7551,N_5103,N_4842);
nor U7552 (N_7552,N_4588,N_5884);
and U7553 (N_7553,N_5432,N_5882);
nor U7554 (N_7554,N_4581,N_5675);
nor U7555 (N_7555,N_5516,N_4487);
or U7556 (N_7556,N_4449,N_5116);
nor U7557 (N_7557,N_4710,N_4737);
and U7558 (N_7558,N_5416,N_5931);
nor U7559 (N_7559,N_5384,N_4135);
or U7560 (N_7560,N_4976,N_5545);
nand U7561 (N_7561,N_4126,N_4723);
or U7562 (N_7562,N_5814,N_4690);
nor U7563 (N_7563,N_5676,N_5596);
nor U7564 (N_7564,N_4591,N_5470);
nand U7565 (N_7565,N_4278,N_5268);
nand U7566 (N_7566,N_5996,N_5542);
or U7567 (N_7567,N_4762,N_4803);
nor U7568 (N_7568,N_4339,N_5176);
nor U7569 (N_7569,N_4351,N_4537);
nor U7570 (N_7570,N_4793,N_5769);
nand U7571 (N_7571,N_4628,N_4929);
nor U7572 (N_7572,N_5255,N_4912);
and U7573 (N_7573,N_5968,N_5840);
and U7574 (N_7574,N_4307,N_5330);
xor U7575 (N_7575,N_4271,N_4600);
or U7576 (N_7576,N_5795,N_5437);
nor U7577 (N_7577,N_4381,N_5964);
nor U7578 (N_7578,N_5709,N_5657);
nand U7579 (N_7579,N_5666,N_4236);
xnor U7580 (N_7580,N_5099,N_5317);
nand U7581 (N_7581,N_4252,N_5782);
or U7582 (N_7582,N_4657,N_4446);
nor U7583 (N_7583,N_4915,N_4470);
or U7584 (N_7584,N_4374,N_4062);
nor U7585 (N_7585,N_4004,N_5402);
nand U7586 (N_7586,N_5742,N_4496);
and U7587 (N_7587,N_4876,N_4393);
or U7588 (N_7588,N_5945,N_4634);
nor U7589 (N_7589,N_4131,N_5732);
xor U7590 (N_7590,N_4630,N_5320);
or U7591 (N_7591,N_5711,N_5942);
or U7592 (N_7592,N_4062,N_5916);
nor U7593 (N_7593,N_4087,N_5281);
and U7594 (N_7594,N_4377,N_5137);
nand U7595 (N_7595,N_5221,N_5785);
xor U7596 (N_7596,N_4390,N_5598);
nor U7597 (N_7597,N_4041,N_4221);
nand U7598 (N_7598,N_5021,N_4743);
nand U7599 (N_7599,N_5386,N_4195);
and U7600 (N_7600,N_5318,N_4748);
nand U7601 (N_7601,N_4528,N_4044);
or U7602 (N_7602,N_5267,N_5023);
xor U7603 (N_7603,N_4963,N_4294);
nand U7604 (N_7604,N_5353,N_5735);
nand U7605 (N_7605,N_4588,N_4272);
and U7606 (N_7606,N_4997,N_5366);
nor U7607 (N_7607,N_4964,N_4311);
nand U7608 (N_7608,N_5594,N_4448);
xnor U7609 (N_7609,N_5202,N_5985);
nand U7610 (N_7610,N_4903,N_5620);
or U7611 (N_7611,N_5252,N_5905);
nand U7612 (N_7612,N_5721,N_5453);
nand U7613 (N_7613,N_5256,N_5967);
or U7614 (N_7614,N_4014,N_4864);
xnor U7615 (N_7615,N_4138,N_5150);
xor U7616 (N_7616,N_4354,N_4072);
nor U7617 (N_7617,N_4318,N_5684);
nor U7618 (N_7618,N_5478,N_5358);
nor U7619 (N_7619,N_4874,N_5730);
nor U7620 (N_7620,N_5328,N_4546);
or U7621 (N_7621,N_5846,N_5943);
and U7622 (N_7622,N_4093,N_5920);
nor U7623 (N_7623,N_4265,N_5339);
and U7624 (N_7624,N_5095,N_5709);
nor U7625 (N_7625,N_5107,N_4797);
or U7626 (N_7626,N_4951,N_4676);
nand U7627 (N_7627,N_5148,N_4849);
and U7628 (N_7628,N_5670,N_5013);
nor U7629 (N_7629,N_4104,N_5773);
and U7630 (N_7630,N_4172,N_4492);
or U7631 (N_7631,N_5102,N_4939);
xor U7632 (N_7632,N_4173,N_5190);
or U7633 (N_7633,N_4495,N_4577);
nor U7634 (N_7634,N_4187,N_4351);
xor U7635 (N_7635,N_4743,N_5085);
and U7636 (N_7636,N_4055,N_5561);
nand U7637 (N_7637,N_5718,N_5418);
or U7638 (N_7638,N_5968,N_5130);
nor U7639 (N_7639,N_5320,N_4456);
and U7640 (N_7640,N_5526,N_4863);
and U7641 (N_7641,N_4480,N_4331);
and U7642 (N_7642,N_5502,N_4968);
nor U7643 (N_7643,N_4340,N_5001);
nand U7644 (N_7644,N_5831,N_5113);
nand U7645 (N_7645,N_5007,N_5358);
nor U7646 (N_7646,N_4722,N_5004);
and U7647 (N_7647,N_5099,N_4749);
nor U7648 (N_7648,N_5814,N_4377);
or U7649 (N_7649,N_4666,N_4370);
nor U7650 (N_7650,N_4938,N_5706);
nor U7651 (N_7651,N_4784,N_4531);
nand U7652 (N_7652,N_5311,N_5190);
or U7653 (N_7653,N_5090,N_4797);
nor U7654 (N_7654,N_5924,N_4604);
and U7655 (N_7655,N_4601,N_4586);
and U7656 (N_7656,N_4191,N_4461);
and U7657 (N_7657,N_4088,N_4050);
nor U7658 (N_7658,N_5918,N_4116);
xor U7659 (N_7659,N_5699,N_4905);
or U7660 (N_7660,N_5447,N_4099);
and U7661 (N_7661,N_5358,N_4857);
nor U7662 (N_7662,N_5049,N_4034);
nor U7663 (N_7663,N_5425,N_5023);
nor U7664 (N_7664,N_5882,N_4666);
nand U7665 (N_7665,N_5869,N_5583);
xor U7666 (N_7666,N_4261,N_5351);
xor U7667 (N_7667,N_4750,N_5634);
or U7668 (N_7668,N_5042,N_4607);
and U7669 (N_7669,N_5962,N_5309);
nor U7670 (N_7670,N_5272,N_4501);
xnor U7671 (N_7671,N_5101,N_4854);
and U7672 (N_7672,N_4295,N_5046);
or U7673 (N_7673,N_5235,N_4525);
or U7674 (N_7674,N_5161,N_5192);
nor U7675 (N_7675,N_5877,N_4587);
and U7676 (N_7676,N_4386,N_5560);
nand U7677 (N_7677,N_5532,N_5405);
nor U7678 (N_7678,N_5892,N_4309);
and U7679 (N_7679,N_5349,N_4658);
nand U7680 (N_7680,N_4461,N_5465);
nand U7681 (N_7681,N_4935,N_5622);
xor U7682 (N_7682,N_5375,N_5495);
and U7683 (N_7683,N_5028,N_4803);
nor U7684 (N_7684,N_4984,N_4658);
and U7685 (N_7685,N_5615,N_4852);
or U7686 (N_7686,N_4121,N_4284);
nand U7687 (N_7687,N_4909,N_5338);
nor U7688 (N_7688,N_4912,N_4886);
and U7689 (N_7689,N_4174,N_4061);
or U7690 (N_7690,N_5365,N_5378);
or U7691 (N_7691,N_4334,N_4408);
nor U7692 (N_7692,N_5631,N_4278);
and U7693 (N_7693,N_4425,N_4302);
or U7694 (N_7694,N_5765,N_5755);
and U7695 (N_7695,N_4946,N_4897);
nor U7696 (N_7696,N_4593,N_4806);
xnor U7697 (N_7697,N_4422,N_5129);
nor U7698 (N_7698,N_5070,N_5285);
or U7699 (N_7699,N_5103,N_4718);
or U7700 (N_7700,N_5864,N_5177);
nand U7701 (N_7701,N_4128,N_5348);
and U7702 (N_7702,N_4146,N_4960);
or U7703 (N_7703,N_4593,N_4446);
nand U7704 (N_7704,N_5283,N_4312);
nand U7705 (N_7705,N_4362,N_5354);
and U7706 (N_7706,N_4994,N_5073);
xor U7707 (N_7707,N_5168,N_4713);
nand U7708 (N_7708,N_5217,N_5888);
nor U7709 (N_7709,N_4755,N_4546);
or U7710 (N_7710,N_4510,N_4176);
or U7711 (N_7711,N_5528,N_4704);
nand U7712 (N_7712,N_4845,N_4497);
nand U7713 (N_7713,N_4047,N_5935);
nor U7714 (N_7714,N_5150,N_4910);
and U7715 (N_7715,N_5346,N_5415);
or U7716 (N_7716,N_4558,N_5717);
xnor U7717 (N_7717,N_5730,N_4450);
nand U7718 (N_7718,N_5017,N_5389);
nand U7719 (N_7719,N_4152,N_4762);
nor U7720 (N_7720,N_4390,N_4872);
and U7721 (N_7721,N_5185,N_4794);
xnor U7722 (N_7722,N_4125,N_4348);
nor U7723 (N_7723,N_4016,N_4933);
nor U7724 (N_7724,N_4833,N_5156);
nor U7725 (N_7725,N_4247,N_5635);
or U7726 (N_7726,N_4167,N_4216);
nand U7727 (N_7727,N_4522,N_5734);
nand U7728 (N_7728,N_4114,N_4668);
and U7729 (N_7729,N_4251,N_5055);
nand U7730 (N_7730,N_5319,N_4166);
nand U7731 (N_7731,N_4142,N_4304);
and U7732 (N_7732,N_4277,N_5142);
and U7733 (N_7733,N_5273,N_4738);
or U7734 (N_7734,N_5776,N_5779);
or U7735 (N_7735,N_4793,N_5755);
and U7736 (N_7736,N_4374,N_5017);
nor U7737 (N_7737,N_5553,N_4613);
nand U7738 (N_7738,N_4444,N_5953);
nand U7739 (N_7739,N_5483,N_5626);
nor U7740 (N_7740,N_5579,N_5756);
nor U7741 (N_7741,N_5883,N_5804);
and U7742 (N_7742,N_5905,N_5871);
and U7743 (N_7743,N_5715,N_4651);
nor U7744 (N_7744,N_4251,N_5051);
or U7745 (N_7745,N_5233,N_5758);
or U7746 (N_7746,N_4333,N_5802);
nor U7747 (N_7747,N_5470,N_4449);
nand U7748 (N_7748,N_4378,N_4721);
nor U7749 (N_7749,N_5075,N_4660);
nand U7750 (N_7750,N_4358,N_4217);
xor U7751 (N_7751,N_4522,N_4660);
and U7752 (N_7752,N_4628,N_4688);
nor U7753 (N_7753,N_4286,N_4644);
nor U7754 (N_7754,N_5065,N_5711);
and U7755 (N_7755,N_5570,N_4983);
and U7756 (N_7756,N_4124,N_4608);
nor U7757 (N_7757,N_4345,N_4346);
or U7758 (N_7758,N_5201,N_4741);
xnor U7759 (N_7759,N_5309,N_5267);
xor U7760 (N_7760,N_4671,N_4021);
xor U7761 (N_7761,N_4844,N_5851);
nand U7762 (N_7762,N_5699,N_5355);
xor U7763 (N_7763,N_4283,N_5712);
xor U7764 (N_7764,N_5477,N_5489);
and U7765 (N_7765,N_5791,N_4207);
or U7766 (N_7766,N_5224,N_5356);
or U7767 (N_7767,N_5878,N_5187);
or U7768 (N_7768,N_4165,N_5219);
nor U7769 (N_7769,N_4226,N_4903);
nand U7770 (N_7770,N_4097,N_4243);
and U7771 (N_7771,N_5413,N_4192);
and U7772 (N_7772,N_4064,N_5562);
nand U7773 (N_7773,N_4710,N_5216);
or U7774 (N_7774,N_5588,N_5483);
xor U7775 (N_7775,N_4778,N_5693);
and U7776 (N_7776,N_4665,N_5684);
and U7777 (N_7777,N_4542,N_5264);
or U7778 (N_7778,N_4915,N_4840);
nor U7779 (N_7779,N_5399,N_5931);
and U7780 (N_7780,N_4167,N_5193);
nor U7781 (N_7781,N_4907,N_4082);
or U7782 (N_7782,N_5084,N_5175);
and U7783 (N_7783,N_5468,N_4248);
and U7784 (N_7784,N_4028,N_5046);
nand U7785 (N_7785,N_5161,N_4128);
or U7786 (N_7786,N_4273,N_4174);
nor U7787 (N_7787,N_5461,N_5715);
nand U7788 (N_7788,N_4087,N_5580);
or U7789 (N_7789,N_4113,N_4031);
or U7790 (N_7790,N_4760,N_4208);
nor U7791 (N_7791,N_5245,N_4676);
nor U7792 (N_7792,N_4409,N_4863);
or U7793 (N_7793,N_4744,N_4923);
or U7794 (N_7794,N_5798,N_4980);
nand U7795 (N_7795,N_4678,N_5738);
and U7796 (N_7796,N_5563,N_4026);
nand U7797 (N_7797,N_4065,N_4228);
or U7798 (N_7798,N_4664,N_5049);
xnor U7799 (N_7799,N_5091,N_4641);
nor U7800 (N_7800,N_5465,N_4981);
or U7801 (N_7801,N_5444,N_5934);
nand U7802 (N_7802,N_4192,N_5909);
and U7803 (N_7803,N_5680,N_4724);
nand U7804 (N_7804,N_4993,N_4809);
and U7805 (N_7805,N_4970,N_5979);
or U7806 (N_7806,N_5734,N_4186);
nand U7807 (N_7807,N_5398,N_5579);
nand U7808 (N_7808,N_5602,N_5575);
and U7809 (N_7809,N_4383,N_5545);
and U7810 (N_7810,N_5461,N_4195);
nor U7811 (N_7811,N_5886,N_5429);
nand U7812 (N_7812,N_4557,N_5244);
and U7813 (N_7813,N_4458,N_4764);
nand U7814 (N_7814,N_5984,N_5796);
nor U7815 (N_7815,N_4585,N_4654);
nor U7816 (N_7816,N_5911,N_4996);
or U7817 (N_7817,N_5735,N_5606);
and U7818 (N_7818,N_5317,N_5661);
nand U7819 (N_7819,N_4544,N_5860);
nor U7820 (N_7820,N_5422,N_5219);
and U7821 (N_7821,N_4358,N_5813);
nand U7822 (N_7822,N_5890,N_5398);
nor U7823 (N_7823,N_5483,N_5555);
nand U7824 (N_7824,N_5604,N_5396);
nor U7825 (N_7825,N_5414,N_5220);
nand U7826 (N_7826,N_5147,N_4768);
nand U7827 (N_7827,N_5557,N_5694);
or U7828 (N_7828,N_5348,N_4868);
nor U7829 (N_7829,N_5121,N_4085);
nor U7830 (N_7830,N_5454,N_5489);
nor U7831 (N_7831,N_5757,N_5931);
xnor U7832 (N_7832,N_4792,N_5163);
or U7833 (N_7833,N_5555,N_5919);
and U7834 (N_7834,N_4099,N_5893);
nand U7835 (N_7835,N_4812,N_5076);
nand U7836 (N_7836,N_4130,N_4564);
xnor U7837 (N_7837,N_5944,N_5678);
nand U7838 (N_7838,N_5776,N_4242);
xnor U7839 (N_7839,N_5763,N_4261);
and U7840 (N_7840,N_5162,N_5497);
and U7841 (N_7841,N_4247,N_5092);
xnor U7842 (N_7842,N_5984,N_4118);
and U7843 (N_7843,N_4496,N_4715);
nor U7844 (N_7844,N_4140,N_5692);
nor U7845 (N_7845,N_4571,N_4551);
and U7846 (N_7846,N_4706,N_4027);
or U7847 (N_7847,N_5260,N_4930);
nor U7848 (N_7848,N_5822,N_5473);
or U7849 (N_7849,N_4232,N_4284);
nand U7850 (N_7850,N_4491,N_4972);
nand U7851 (N_7851,N_4291,N_4790);
nand U7852 (N_7852,N_4984,N_4778);
xnor U7853 (N_7853,N_4479,N_5072);
nand U7854 (N_7854,N_4011,N_5308);
or U7855 (N_7855,N_5656,N_4675);
and U7856 (N_7856,N_4354,N_4045);
and U7857 (N_7857,N_5048,N_4994);
nand U7858 (N_7858,N_4886,N_4783);
and U7859 (N_7859,N_4214,N_5253);
nand U7860 (N_7860,N_4466,N_5671);
nand U7861 (N_7861,N_5414,N_5823);
nand U7862 (N_7862,N_4646,N_5782);
nand U7863 (N_7863,N_5963,N_5695);
or U7864 (N_7864,N_4051,N_4266);
nor U7865 (N_7865,N_5926,N_4676);
nor U7866 (N_7866,N_4581,N_5137);
nor U7867 (N_7867,N_4261,N_4047);
xor U7868 (N_7868,N_4523,N_4250);
nor U7869 (N_7869,N_4807,N_5779);
or U7870 (N_7870,N_4971,N_5086);
and U7871 (N_7871,N_5834,N_5849);
nor U7872 (N_7872,N_5250,N_5028);
nand U7873 (N_7873,N_4239,N_5155);
nor U7874 (N_7874,N_4426,N_4742);
nand U7875 (N_7875,N_4487,N_5948);
or U7876 (N_7876,N_4542,N_4337);
and U7877 (N_7877,N_5171,N_5480);
or U7878 (N_7878,N_5978,N_4283);
and U7879 (N_7879,N_5896,N_4571);
nor U7880 (N_7880,N_4362,N_4520);
nor U7881 (N_7881,N_5162,N_4247);
nand U7882 (N_7882,N_5283,N_5259);
nand U7883 (N_7883,N_5734,N_4878);
or U7884 (N_7884,N_5340,N_4155);
xnor U7885 (N_7885,N_4743,N_5104);
or U7886 (N_7886,N_5243,N_4555);
or U7887 (N_7887,N_4708,N_4552);
and U7888 (N_7888,N_5094,N_5846);
and U7889 (N_7889,N_4024,N_4374);
and U7890 (N_7890,N_4075,N_4586);
or U7891 (N_7891,N_5208,N_4882);
or U7892 (N_7892,N_4259,N_5113);
xor U7893 (N_7893,N_4302,N_5925);
xor U7894 (N_7894,N_5228,N_4727);
or U7895 (N_7895,N_5263,N_5526);
nand U7896 (N_7896,N_4093,N_4464);
nand U7897 (N_7897,N_5675,N_4421);
nand U7898 (N_7898,N_5969,N_5537);
and U7899 (N_7899,N_5995,N_5198);
nor U7900 (N_7900,N_4121,N_4422);
nor U7901 (N_7901,N_5590,N_4677);
nand U7902 (N_7902,N_4276,N_5753);
or U7903 (N_7903,N_5573,N_5853);
and U7904 (N_7904,N_4440,N_4363);
or U7905 (N_7905,N_5177,N_5669);
nor U7906 (N_7906,N_4662,N_5634);
xor U7907 (N_7907,N_4373,N_4270);
nand U7908 (N_7908,N_5099,N_5012);
or U7909 (N_7909,N_4653,N_5791);
or U7910 (N_7910,N_4410,N_4630);
nor U7911 (N_7911,N_5454,N_5266);
nor U7912 (N_7912,N_4045,N_5556);
or U7913 (N_7913,N_5527,N_4467);
nand U7914 (N_7914,N_5615,N_5937);
nor U7915 (N_7915,N_4867,N_4076);
nand U7916 (N_7916,N_4258,N_4433);
nor U7917 (N_7917,N_4082,N_4222);
or U7918 (N_7918,N_5824,N_4149);
or U7919 (N_7919,N_4190,N_4076);
xor U7920 (N_7920,N_4201,N_4446);
or U7921 (N_7921,N_4853,N_5465);
xor U7922 (N_7922,N_4491,N_5466);
and U7923 (N_7923,N_4471,N_4522);
nor U7924 (N_7924,N_4092,N_5730);
or U7925 (N_7925,N_5759,N_4631);
nand U7926 (N_7926,N_5348,N_4217);
nand U7927 (N_7927,N_4407,N_4239);
or U7928 (N_7928,N_5986,N_4445);
or U7929 (N_7929,N_5223,N_5700);
or U7930 (N_7930,N_4645,N_5740);
nor U7931 (N_7931,N_5124,N_4189);
xor U7932 (N_7932,N_5179,N_5318);
nor U7933 (N_7933,N_4581,N_5739);
or U7934 (N_7934,N_5475,N_5683);
nor U7935 (N_7935,N_5778,N_5499);
nand U7936 (N_7936,N_5850,N_4646);
xor U7937 (N_7937,N_4028,N_4251);
and U7938 (N_7938,N_5386,N_5237);
nor U7939 (N_7939,N_5681,N_5765);
or U7940 (N_7940,N_4673,N_5768);
and U7941 (N_7941,N_4355,N_5650);
or U7942 (N_7942,N_5399,N_4312);
and U7943 (N_7943,N_4653,N_4347);
nor U7944 (N_7944,N_5585,N_4033);
and U7945 (N_7945,N_5812,N_4716);
or U7946 (N_7946,N_4362,N_4941);
and U7947 (N_7947,N_5709,N_5066);
nor U7948 (N_7948,N_4656,N_5262);
or U7949 (N_7949,N_4998,N_4436);
or U7950 (N_7950,N_5121,N_5814);
nor U7951 (N_7951,N_4648,N_4027);
or U7952 (N_7952,N_5569,N_5344);
xnor U7953 (N_7953,N_5848,N_5102);
or U7954 (N_7954,N_5648,N_5302);
and U7955 (N_7955,N_5130,N_5558);
nor U7956 (N_7956,N_4945,N_5779);
or U7957 (N_7957,N_4349,N_4572);
nand U7958 (N_7958,N_4041,N_4974);
nand U7959 (N_7959,N_5826,N_4614);
nor U7960 (N_7960,N_4332,N_4759);
nand U7961 (N_7961,N_4648,N_4402);
or U7962 (N_7962,N_5565,N_5984);
xnor U7963 (N_7963,N_4151,N_4297);
or U7964 (N_7964,N_4442,N_5955);
or U7965 (N_7965,N_4281,N_4487);
nand U7966 (N_7966,N_5446,N_5756);
and U7967 (N_7967,N_4270,N_5860);
and U7968 (N_7968,N_5245,N_5784);
or U7969 (N_7969,N_4557,N_5757);
nand U7970 (N_7970,N_5564,N_5955);
nor U7971 (N_7971,N_5632,N_5846);
or U7972 (N_7972,N_5726,N_4765);
and U7973 (N_7973,N_4413,N_5423);
and U7974 (N_7974,N_5201,N_4121);
or U7975 (N_7975,N_4661,N_5936);
nand U7976 (N_7976,N_5025,N_4486);
and U7977 (N_7977,N_5376,N_5017);
and U7978 (N_7978,N_4380,N_4388);
and U7979 (N_7979,N_5300,N_5349);
and U7980 (N_7980,N_5106,N_5478);
and U7981 (N_7981,N_4454,N_4317);
nor U7982 (N_7982,N_4405,N_4486);
or U7983 (N_7983,N_5232,N_5408);
nor U7984 (N_7984,N_5667,N_5581);
or U7985 (N_7985,N_5782,N_4104);
or U7986 (N_7986,N_4486,N_5856);
xnor U7987 (N_7987,N_4248,N_4149);
or U7988 (N_7988,N_4209,N_4736);
nor U7989 (N_7989,N_5239,N_4176);
nor U7990 (N_7990,N_5003,N_4714);
nand U7991 (N_7991,N_4876,N_4435);
or U7992 (N_7992,N_4597,N_5783);
or U7993 (N_7993,N_4208,N_4936);
and U7994 (N_7994,N_5769,N_4692);
xor U7995 (N_7995,N_5116,N_5961);
nor U7996 (N_7996,N_5873,N_4215);
or U7997 (N_7997,N_5193,N_4390);
nor U7998 (N_7998,N_5168,N_4565);
nand U7999 (N_7999,N_5337,N_4356);
nor U8000 (N_8000,N_7144,N_7713);
and U8001 (N_8001,N_7671,N_6907);
nand U8002 (N_8002,N_6023,N_6870);
and U8003 (N_8003,N_6046,N_6917);
and U8004 (N_8004,N_7841,N_6122);
xnor U8005 (N_8005,N_7892,N_6876);
and U8006 (N_8006,N_6016,N_6922);
nor U8007 (N_8007,N_7706,N_6366);
nor U8008 (N_8008,N_7999,N_6019);
or U8009 (N_8009,N_7285,N_7712);
and U8010 (N_8010,N_6437,N_7330);
or U8011 (N_8011,N_7836,N_6164);
and U8012 (N_8012,N_7755,N_7690);
xnor U8013 (N_8013,N_6483,N_6012);
or U8014 (N_8014,N_7694,N_6079);
nor U8015 (N_8015,N_7499,N_7821);
nor U8016 (N_8016,N_7984,N_6142);
and U8017 (N_8017,N_7398,N_7414);
xor U8018 (N_8018,N_7155,N_7923);
or U8019 (N_8019,N_6027,N_6172);
or U8020 (N_8020,N_6432,N_6977);
nor U8021 (N_8021,N_6487,N_6825);
or U8022 (N_8022,N_6317,N_7983);
and U8023 (N_8023,N_6175,N_7786);
xnor U8024 (N_8024,N_6123,N_6227);
or U8025 (N_8025,N_7185,N_7753);
xor U8026 (N_8026,N_6065,N_6213);
and U8027 (N_8027,N_6404,N_7040);
and U8028 (N_8028,N_6346,N_7976);
or U8029 (N_8029,N_7463,N_6297);
or U8030 (N_8030,N_7909,N_6200);
or U8031 (N_8031,N_6996,N_6493);
and U8032 (N_8032,N_6217,N_6704);
nor U8033 (N_8033,N_6008,N_7558);
nand U8034 (N_8034,N_6764,N_7922);
or U8035 (N_8035,N_6176,N_7241);
and U8036 (N_8036,N_6522,N_6068);
nand U8037 (N_8037,N_7661,N_6697);
nand U8038 (N_8038,N_6341,N_7708);
nor U8039 (N_8039,N_6191,N_6475);
and U8040 (N_8040,N_6334,N_7691);
or U8041 (N_8041,N_7579,N_6375);
nor U8042 (N_8042,N_6116,N_6596);
nor U8043 (N_8043,N_6295,N_7848);
and U8044 (N_8044,N_6115,N_7098);
nand U8045 (N_8045,N_6731,N_7050);
and U8046 (N_8046,N_7022,N_6231);
nor U8047 (N_8047,N_6458,N_7964);
xor U8048 (N_8048,N_6258,N_7352);
nand U8049 (N_8049,N_6809,N_6787);
nor U8050 (N_8050,N_6574,N_6770);
nand U8051 (N_8051,N_7798,N_6933);
nand U8052 (N_8052,N_6170,N_6415);
nor U8053 (N_8053,N_7944,N_7948);
xnor U8054 (N_8054,N_7177,N_6920);
nand U8055 (N_8055,N_6670,N_7009);
nor U8056 (N_8056,N_6815,N_7262);
nand U8057 (N_8057,N_6009,N_6496);
nand U8058 (N_8058,N_7292,N_7271);
and U8059 (N_8059,N_7108,N_7598);
xor U8060 (N_8060,N_7683,N_6740);
nand U8061 (N_8061,N_7876,N_7316);
or U8062 (N_8062,N_7808,N_6605);
xnor U8063 (N_8063,N_6700,N_7510);
or U8064 (N_8064,N_6193,N_7843);
xnor U8065 (N_8065,N_6249,N_7846);
nor U8066 (N_8066,N_7505,N_6843);
nand U8067 (N_8067,N_7387,N_6197);
or U8068 (N_8068,N_6204,N_7130);
nand U8069 (N_8069,N_6344,N_6822);
and U8070 (N_8070,N_6136,N_6631);
and U8071 (N_8071,N_7719,N_6005);
and U8072 (N_8072,N_7560,N_7589);
nand U8073 (N_8073,N_6665,N_6382);
nand U8074 (N_8074,N_7592,N_6951);
or U8075 (N_8075,N_7196,N_7617);
and U8076 (N_8076,N_6167,N_7915);
nor U8077 (N_8077,N_6128,N_6099);
or U8078 (N_8078,N_6971,N_7913);
or U8079 (N_8079,N_7202,N_6982);
or U8080 (N_8080,N_7195,N_6883);
or U8081 (N_8081,N_7379,N_6474);
nand U8082 (N_8082,N_7587,N_6328);
and U8083 (N_8083,N_7498,N_7406);
nand U8084 (N_8084,N_7260,N_7384);
nor U8085 (N_8085,N_7267,N_6538);
or U8086 (N_8086,N_7056,N_7497);
xor U8087 (N_8087,N_7942,N_7169);
nand U8088 (N_8088,N_7917,N_6385);
or U8089 (N_8089,N_7367,N_6096);
nand U8090 (N_8090,N_7862,N_6272);
and U8091 (N_8091,N_7064,N_7404);
and U8092 (N_8092,N_7501,N_6025);
nand U8093 (N_8093,N_6285,N_6148);
nand U8094 (N_8094,N_7326,N_6205);
and U8095 (N_8095,N_6091,N_7466);
nand U8096 (N_8096,N_7073,N_7614);
and U8097 (N_8097,N_6979,N_7817);
and U8098 (N_8098,N_7973,N_6035);
nor U8099 (N_8099,N_6466,N_7464);
nand U8100 (N_8100,N_7325,N_6677);
nand U8101 (N_8101,N_7960,N_6717);
and U8102 (N_8102,N_7628,N_6515);
and U8103 (N_8103,N_6491,N_7420);
nand U8104 (N_8104,N_6645,N_6831);
nor U8105 (N_8105,N_6743,N_6662);
or U8106 (N_8106,N_7572,N_7238);
or U8107 (N_8107,N_6699,N_7904);
or U8108 (N_8108,N_6101,N_7128);
nor U8109 (N_8109,N_6503,N_7882);
and U8110 (N_8110,N_6058,N_7465);
nor U8111 (N_8111,N_6048,N_6462);
and U8112 (N_8112,N_6575,N_6226);
and U8113 (N_8113,N_7473,N_6674);
xor U8114 (N_8114,N_6756,N_6924);
nand U8115 (N_8115,N_7556,N_6439);
and U8116 (N_8116,N_7150,N_7599);
nor U8117 (N_8117,N_6931,N_6838);
and U8118 (N_8118,N_6810,N_7596);
nand U8119 (N_8119,N_7072,N_7375);
xnor U8120 (N_8120,N_6082,N_7158);
or U8121 (N_8121,N_7865,N_7602);
or U8122 (N_8122,N_6848,N_7554);
and U8123 (N_8123,N_7969,N_6429);
or U8124 (N_8124,N_7776,N_7553);
and U8125 (N_8125,N_7941,N_6519);
nand U8126 (N_8126,N_7345,N_7622);
and U8127 (N_8127,N_7322,N_7688);
nand U8128 (N_8128,N_7747,N_7203);
nand U8129 (N_8129,N_7259,N_6311);
or U8130 (N_8130,N_6727,N_6964);
and U8131 (N_8131,N_7548,N_7640);
nand U8132 (N_8132,N_6448,N_7320);
xor U8133 (N_8133,N_7933,N_7122);
nor U8134 (N_8134,N_6780,N_6853);
nor U8135 (N_8135,N_6248,N_6929);
and U8136 (N_8136,N_7716,N_6927);
nor U8137 (N_8137,N_6688,N_7257);
or U8138 (N_8138,N_7936,N_7784);
xor U8139 (N_8139,N_6441,N_6761);
or U8140 (N_8140,N_6478,N_7378);
xnor U8141 (N_8141,N_7791,N_7439);
nor U8142 (N_8142,N_7745,N_7343);
or U8143 (N_8143,N_7675,N_7047);
nand U8144 (N_8144,N_7023,N_7903);
or U8145 (N_8145,N_6088,N_6908);
or U8146 (N_8146,N_7512,N_6266);
nand U8147 (N_8147,N_6653,N_6267);
nand U8148 (N_8148,N_6381,N_7232);
or U8149 (N_8149,N_6215,N_6952);
and U8150 (N_8150,N_7878,N_7492);
or U8151 (N_8151,N_7153,N_7114);
and U8152 (N_8152,N_6552,N_6518);
and U8153 (N_8153,N_6826,N_6513);
xnor U8154 (N_8154,N_6919,N_7718);
or U8155 (N_8155,N_7168,N_7361);
nor U8156 (N_8156,N_6134,N_7243);
nor U8157 (N_8157,N_7568,N_6753);
xnor U8158 (N_8158,N_6582,N_6002);
nand U8159 (N_8159,N_6935,N_7340);
nor U8160 (N_8160,N_6453,N_6257);
xnor U8161 (N_8161,N_6161,N_7118);
xor U8162 (N_8162,N_6560,N_6978);
nand U8163 (N_8163,N_6154,N_6564);
nand U8164 (N_8164,N_7365,N_7523);
nor U8165 (N_8165,N_6943,N_6856);
nand U8166 (N_8166,N_7240,N_7458);
or U8167 (N_8167,N_6472,N_6465);
xor U8168 (N_8168,N_7785,N_6658);
or U8169 (N_8169,N_6018,N_7820);
or U8170 (N_8170,N_6910,N_6745);
nand U8171 (N_8171,N_6421,N_6001);
nor U8172 (N_8172,N_7364,N_6501);
nor U8173 (N_8173,N_6223,N_7571);
or U8174 (N_8174,N_7468,N_6551);
or U8175 (N_8175,N_6335,N_7666);
and U8176 (N_8176,N_7724,N_7715);
or U8177 (N_8177,N_7738,N_6572);
and U8178 (N_8178,N_7812,N_7974);
nor U8179 (N_8179,N_6879,N_7918);
nor U8180 (N_8180,N_7453,N_6313);
nor U8181 (N_8181,N_6999,N_7522);
and U8182 (N_8182,N_6893,N_6064);
nand U8183 (N_8183,N_7729,N_7597);
nand U8184 (N_8184,N_7629,N_7607);
nor U8185 (N_8185,N_6736,N_6632);
xor U8186 (N_8186,N_6681,N_7570);
xnor U8187 (N_8187,N_7758,N_6319);
nand U8188 (N_8188,N_7005,N_7831);
nand U8189 (N_8189,N_7350,N_7231);
and U8190 (N_8190,N_6788,N_7653);
or U8191 (N_8191,N_6782,N_6849);
nand U8192 (N_8192,N_7957,N_6365);
or U8193 (N_8193,N_7462,N_6994);
nor U8194 (N_8194,N_7654,N_7225);
and U8195 (N_8195,N_6647,N_7315);
nand U8196 (N_8196,N_6536,N_6739);
or U8197 (N_8197,N_6891,N_7164);
nor U8198 (N_8198,N_7583,N_6639);
or U8199 (N_8199,N_6377,N_6316);
nor U8200 (N_8200,N_7689,N_6679);
and U8201 (N_8201,N_7682,N_7383);
nor U8202 (N_8202,N_6837,N_7481);
and U8203 (N_8203,N_7778,N_6436);
nor U8204 (N_8204,N_6349,N_7947);
and U8205 (N_8205,N_7437,N_6246);
nor U8206 (N_8206,N_7054,N_7972);
or U8207 (N_8207,N_7392,N_7057);
nor U8208 (N_8208,N_7714,N_6540);
and U8209 (N_8209,N_6000,N_6409);
and U8210 (N_8210,N_6746,N_7020);
nand U8211 (N_8211,N_6062,N_6989);
or U8212 (N_8212,N_6430,N_7783);
nor U8213 (N_8213,N_6203,N_6701);
or U8214 (N_8214,N_6998,N_7276);
nor U8215 (N_8215,N_7170,N_6566);
nand U8216 (N_8216,N_7199,N_6671);
nor U8217 (N_8217,N_7389,N_6767);
nor U8218 (N_8218,N_6616,N_7218);
xnor U8219 (N_8219,N_7066,N_6823);
and U8220 (N_8220,N_7686,N_6238);
and U8221 (N_8221,N_7163,N_7060);
nor U8222 (N_8222,N_7509,N_7253);
or U8223 (N_8223,N_7403,N_7102);
xnor U8224 (N_8224,N_7447,N_6781);
nand U8225 (N_8225,N_6661,N_7584);
nand U8226 (N_8226,N_7782,N_6981);
nand U8227 (N_8227,N_6839,N_7258);
or U8228 (N_8228,N_6155,N_6599);
nor U8229 (N_8229,N_6094,N_7800);
and U8230 (N_8230,N_7669,N_6145);
nor U8231 (N_8231,N_6166,N_7256);
nor U8232 (N_8232,N_7329,N_7857);
or U8233 (N_8233,N_7457,N_7979);
or U8234 (N_8234,N_6043,N_6031);
or U8235 (N_8235,N_7582,N_6629);
or U8236 (N_8236,N_6038,N_7363);
nor U8237 (N_8237,N_7574,N_7989);
and U8238 (N_8238,N_6174,N_6022);
and U8239 (N_8239,N_7312,N_6526);
nand U8240 (N_8240,N_6741,N_6576);
or U8241 (N_8241,N_6709,N_6723);
and U8242 (N_8242,N_6218,N_7519);
and U8243 (N_8243,N_6742,N_7826);
nor U8244 (N_8244,N_6106,N_7588);
nor U8245 (N_8245,N_7143,N_6817);
and U8246 (N_8246,N_6769,N_6725);
nor U8247 (N_8247,N_7112,N_6686);
nand U8248 (N_8248,N_7099,N_6484);
nor U8249 (N_8249,N_6081,N_7513);
nor U8250 (N_8250,N_6874,N_6779);
or U8251 (N_8251,N_6014,N_6733);
xor U8252 (N_8252,N_7393,N_6868);
and U8253 (N_8253,N_7052,N_6798);
or U8254 (N_8254,N_6814,N_6419);
nor U8255 (N_8255,N_7701,N_6512);
or U8256 (N_8256,N_7087,N_7129);
nand U8257 (N_8257,N_7853,N_6221);
xor U8258 (N_8258,N_7905,N_7995);
and U8259 (N_8259,N_6940,N_7699);
nor U8260 (N_8260,N_7968,N_7110);
nor U8261 (N_8261,N_6408,N_7095);
nand U8262 (N_8262,N_6323,N_7839);
or U8263 (N_8263,N_6765,N_7310);
xor U8264 (N_8264,N_7448,N_7665);
and U8265 (N_8265,N_7487,N_7603);
or U8266 (N_8266,N_6942,N_6579);
xor U8267 (N_8267,N_6860,N_7934);
nand U8268 (N_8268,N_7245,N_7667);
nor U8269 (N_8269,N_7673,N_6553);
nor U8270 (N_8270,N_7849,N_7562);
or U8271 (N_8271,N_7946,N_6510);
or U8272 (N_8272,N_7002,N_6143);
or U8273 (N_8273,N_6163,N_7390);
nor U8274 (N_8274,N_7722,N_7593);
nor U8275 (N_8275,N_7609,N_6318);
and U8276 (N_8276,N_6786,N_6293);
or U8277 (N_8277,N_7208,N_6695);
xor U8278 (N_8278,N_7438,N_6973);
nor U8279 (N_8279,N_6525,N_7264);
xnor U8280 (N_8280,N_7024,N_6690);
or U8281 (N_8281,N_6990,N_7070);
or U8282 (N_8282,N_7069,N_7189);
xor U8283 (N_8283,N_7695,N_7741);
nor U8284 (N_8284,N_6102,N_6970);
xor U8285 (N_8285,N_6619,N_6738);
nor U8286 (N_8286,N_7261,N_7772);
nand U8287 (N_8287,N_6077,N_6199);
nand U8288 (N_8288,N_6244,N_7115);
nand U8289 (N_8289,N_6118,N_7482);
and U8290 (N_8290,N_7297,N_6895);
nand U8291 (N_8291,N_7925,N_7080);
and U8292 (N_8292,N_7165,N_6644);
or U8293 (N_8293,N_7612,N_7426);
and U8294 (N_8294,N_7950,N_7250);
nor U8295 (N_8295,N_6824,N_6640);
nor U8296 (N_8296,N_7763,N_7978);
and U8297 (N_8297,N_7266,N_7180);
or U8298 (N_8298,N_7495,N_6991);
nor U8299 (N_8299,N_7637,N_7299);
nor U8300 (N_8300,N_6821,N_6196);
and U8301 (N_8301,N_7304,N_7450);
and U8302 (N_8302,N_6857,N_6771);
and U8303 (N_8303,N_6846,N_6212);
and U8304 (N_8304,N_6300,N_7252);
xnor U8305 (N_8305,N_7802,N_7752);
and U8306 (N_8306,N_6461,N_7930);
or U8307 (N_8307,N_6251,N_7119);
nor U8308 (N_8308,N_7958,N_6371);
and U8309 (N_8309,N_7200,N_7756);
nand U8310 (N_8310,N_7814,N_6353);
nor U8311 (N_8311,N_7415,N_7479);
nor U8312 (N_8312,N_6892,N_6656);
and U8313 (N_8313,N_7425,N_7906);
nand U8314 (N_8314,N_6828,N_7751);
or U8315 (N_8315,N_6953,N_6708);
nor U8316 (N_8316,N_7990,N_7764);
nand U8317 (N_8317,N_6032,N_7178);
nor U8318 (N_8318,N_6119,N_6785);
nand U8319 (N_8319,N_7885,N_7920);
or U8320 (N_8320,N_6378,N_7919);
nand U8321 (N_8321,N_7655,N_6884);
and U8322 (N_8322,N_7212,N_6398);
nand U8323 (N_8323,N_7435,N_6454);
or U8324 (N_8324,N_7334,N_6356);
nor U8325 (N_8325,N_6694,N_7723);
nor U8326 (N_8326,N_7376,N_6889);
nor U8327 (N_8327,N_6277,N_7179);
nor U8328 (N_8328,N_7779,N_6772);
nor U8329 (N_8329,N_7664,N_7027);
nand U8330 (N_8330,N_6948,N_6230);
nor U8331 (N_8331,N_7339,N_6737);
xnor U8332 (N_8332,N_7018,N_6157);
or U8333 (N_8333,N_6726,N_7873);
nand U8334 (N_8334,N_6744,N_6288);
nand U8335 (N_8335,N_6869,N_7059);
nand U8336 (N_8336,N_6958,N_6263);
nor U8337 (N_8337,N_6021,N_7532);
nand U8338 (N_8338,N_6235,N_7391);
and U8339 (N_8339,N_6792,N_6355);
or U8340 (N_8340,N_7140,N_6533);
nor U8341 (N_8341,N_7270,N_6926);
or U8342 (N_8342,N_7549,N_7725);
or U8343 (N_8343,N_6281,N_6125);
nor U8344 (N_8344,N_7046,N_7374);
and U8345 (N_8345,N_7039,N_6053);
and U8346 (N_8346,N_7618,N_7488);
nor U8347 (N_8347,N_7460,N_6292);
and U8348 (N_8348,N_7139,N_6768);
nand U8349 (N_8349,N_6358,N_7636);
nor U8350 (N_8350,N_7818,N_7507);
or U8351 (N_8351,N_6333,N_6185);
nand U8352 (N_8352,N_7840,N_7237);
nand U8353 (N_8353,N_7454,N_7327);
or U8354 (N_8354,N_7044,N_7648);
nand U8355 (N_8355,N_7174,N_7159);
or U8356 (N_8356,N_7141,N_7000);
and U8357 (N_8357,N_6036,N_7182);
xnor U8358 (N_8358,N_6603,N_7564);
or U8359 (N_8359,N_7789,N_6485);
nor U8360 (N_8360,N_7351,N_7888);
or U8361 (N_8361,N_7017,N_6852);
and U8362 (N_8362,N_6243,N_6011);
nand U8363 (N_8363,N_7530,N_7035);
xor U8364 (N_8364,N_7117,N_6443);
nor U8365 (N_8365,N_6312,N_6111);
nor U8366 (N_8366,N_6137,N_6684);
nand U8367 (N_8367,N_6555,N_7992);
nand U8368 (N_8368,N_6992,N_6703);
nor U8369 (N_8369,N_6628,N_7490);
xnor U8370 (N_8370,N_6840,N_6886);
xor U8371 (N_8371,N_6880,N_7216);
nor U8372 (N_8372,N_6370,N_7649);
and U8373 (N_8373,N_6969,N_6354);
nor U8374 (N_8374,N_7824,N_7058);
xnor U8375 (N_8375,N_6711,N_6855);
or U8376 (N_8376,N_7194,N_7739);
nor U8377 (N_8377,N_7434,N_7254);
nor U8378 (N_8378,N_7881,N_7894);
nand U8379 (N_8379,N_6151,N_7503);
xor U8380 (N_8380,N_6626,N_7381);
nand U8381 (N_8381,N_7053,N_7227);
xnor U8382 (N_8382,N_7301,N_7161);
nand U8383 (N_8383,N_6184,N_6417);
or U8384 (N_8384,N_6897,N_6187);
and U8385 (N_8385,N_6804,N_7951);
and U8386 (N_8386,N_7324,N_6539);
or U8387 (N_8387,N_7590,N_6294);
xnor U8388 (N_8388,N_7176,N_6245);
nand U8389 (N_8389,N_6080,N_6988);
nand U8390 (N_8390,N_7470,N_6597);
nand U8391 (N_8391,N_7823,N_7547);
and U8392 (N_8392,N_6265,N_6655);
xnor U8393 (N_8393,N_7284,N_7581);
nand U8394 (N_8394,N_7369,N_6369);
xnor U8395 (N_8395,N_6511,N_7215);
xor U8396 (N_8396,N_7293,N_6577);
nand U8397 (N_8397,N_7015,N_6342);
or U8398 (N_8398,N_6712,N_6449);
or U8399 (N_8399,N_7348,N_7485);
or U8400 (N_8400,N_6286,N_6620);
or U8401 (N_8401,N_6851,N_6089);
nand U8402 (N_8402,N_7737,N_6867);
and U8403 (N_8403,N_7852,N_6055);
nand U8404 (N_8404,N_7138,N_6467);
nand U8405 (N_8405,N_7401,N_6797);
or U8406 (N_8406,N_6207,N_6950);
or U8407 (N_8407,N_6219,N_7962);
or U8408 (N_8408,N_6394,N_7996);
xnor U8409 (N_8409,N_6534,N_6702);
nand U8410 (N_8410,N_6098,N_7405);
and U8411 (N_8411,N_6391,N_7550);
or U8412 (N_8412,N_6178,N_7635);
nor U8413 (N_8413,N_6095,N_7157);
or U8414 (N_8414,N_7956,N_7908);
or U8415 (N_8415,N_7514,N_6007);
nand U8416 (N_8416,N_7480,N_6020);
and U8417 (N_8417,N_6259,N_7754);
nor U8418 (N_8418,N_6216,N_6052);
and U8419 (N_8419,N_6060,N_6627);
and U8420 (N_8420,N_7967,N_7864);
and U8421 (N_8421,N_6451,N_6452);
nand U8422 (N_8422,N_6321,N_6320);
nand U8423 (N_8423,N_6169,N_6918);
or U8424 (N_8424,N_7427,N_6132);
and U8425 (N_8425,N_6121,N_7860);
or U8426 (N_8426,N_6400,N_7703);
nor U8427 (N_8427,N_7489,N_7828);
nand U8428 (N_8428,N_7385,N_6865);
nand U8429 (N_8429,N_6672,N_6913);
nand U8430 (N_8430,N_6944,N_6325);
or U8431 (N_8431,N_7566,N_6808);
nand U8432 (N_8432,N_6914,N_7100);
and U8433 (N_8433,N_7407,N_7736);
xnor U8434 (N_8434,N_6130,N_7028);
nor U8435 (N_8435,N_7806,N_7083);
xor U8436 (N_8436,N_6648,N_6482);
nand U8437 (N_8437,N_7993,N_6070);
or U8438 (N_8438,N_6364,N_6747);
nor U8439 (N_8439,N_7889,N_7127);
nand U8440 (N_8440,N_7181,N_6389);
or U8441 (N_8441,N_6571,N_6410);
xor U8442 (N_8442,N_6026,N_6270);
and U8443 (N_8443,N_6608,N_7837);
or U8444 (N_8444,N_6802,N_7145);
nor U8445 (N_8445,N_7982,N_7604);
nor U8446 (N_8446,N_6149,N_7441);
or U8447 (N_8447,N_7032,N_6006);
or U8448 (N_8448,N_6687,N_7132);
nor U8449 (N_8449,N_6847,N_7937);
and U8450 (N_8450,N_7638,N_6882);
nand U8451 (N_8451,N_7162,N_6179);
and U8452 (N_8452,N_7410,N_6600);
nor U8453 (N_8453,N_6508,N_6524);
and U8454 (N_8454,N_7707,N_6411);
nor U8455 (N_8455,N_7049,N_6315);
or U8456 (N_8456,N_7045,N_6836);
nor U8457 (N_8457,N_7236,N_7085);
nor U8458 (N_8458,N_7875,N_7409);
nand U8459 (N_8459,N_7323,N_6634);
or U8460 (N_8460,N_6446,N_7545);
and U8461 (N_8461,N_7680,N_6562);
or U8462 (N_8462,N_7031,N_6468);
nor U8463 (N_8463,N_7309,N_6287);
nand U8464 (N_8464,N_7190,N_6037);
nor U8465 (N_8465,N_6796,N_6489);
or U8466 (N_8466,N_6435,N_7021);
or U8467 (N_8467,N_7493,N_6282);
and U8468 (N_8468,N_6384,N_6983);
and U8469 (N_8469,N_7220,N_6621);
nor U8470 (N_8470,N_7525,N_6376);
nand U8471 (N_8471,N_6784,N_7014);
and U8472 (N_8472,N_7887,N_6201);
and U8473 (N_8473,N_6220,N_6590);
nor U8474 (N_8474,N_7940,N_6233);
nand U8475 (N_8475,N_6017,N_7280);
and U8476 (N_8476,N_6158,N_6190);
nand U8477 (N_8477,N_6598,N_7016);
xnor U8478 (N_8478,N_7765,N_7611);
and U8479 (N_8479,N_6530,N_7477);
nor U8480 (N_8480,N_7959,N_7953);
nor U8481 (N_8481,N_6256,N_7418);
and U8482 (N_8482,N_6829,N_7825);
or U8483 (N_8483,N_6794,N_6659);
nand U8484 (N_8484,N_6594,N_7034);
xnor U8485 (N_8485,N_7402,N_6844);
or U8486 (N_8486,N_6177,N_7349);
or U8487 (N_8487,N_7198,N_6063);
xnor U8488 (N_8488,N_6673,N_6759);
nor U8489 (N_8489,N_6450,N_7899);
xor U8490 (N_8490,N_7247,N_6329);
and U8491 (N_8491,N_6431,N_7397);
nor U8492 (N_8492,N_6863,N_6271);
and U8493 (N_8493,N_6581,N_6275);
nand U8494 (N_8494,N_6949,N_7921);
and U8495 (N_8495,N_6957,N_7900);
or U8496 (N_8496,N_6873,N_6100);
nand U8497 (N_8497,N_6912,N_7803);
nor U8498 (N_8498,N_7469,N_7214);
nand U8499 (N_8499,N_7832,N_6492);
nor U8500 (N_8500,N_7123,N_6229);
or U8501 (N_8501,N_6010,N_6298);
nor U8502 (N_8502,N_6517,N_7711);
and U8503 (N_8503,N_7205,N_7795);
nand U8504 (N_8504,N_6760,N_7585);
xor U8505 (N_8505,N_7970,N_7134);
or U8506 (N_8506,N_6833,N_6660);
and U8507 (N_8507,N_6202,N_6159);
and U8508 (N_8508,N_6327,N_7943);
nand U8509 (N_8509,N_7676,N_6972);
or U8510 (N_8510,N_7626,N_7125);
xor U8511 (N_8511,N_6514,N_7412);
and U8512 (N_8512,N_6795,N_7281);
xnor U8513 (N_8513,N_6749,N_6405);
nor U8514 (N_8514,N_6611,N_7662);
xor U8515 (N_8515,N_7290,N_6336);
nand U8516 (N_8516,N_7858,N_6545);
and U8517 (N_8517,N_6962,N_7787);
nand U8518 (N_8518,N_6580,N_6801);
nand U8519 (N_8519,N_6854,N_7175);
or U8520 (N_8520,N_7606,N_7985);
nand U8521 (N_8521,N_7358,N_7702);
nor U8522 (N_8522,N_6509,N_6250);
xor U8523 (N_8523,N_6811,N_7030);
and U8524 (N_8524,N_6350,N_7101);
nor U8525 (N_8525,N_7907,N_7424);
nor U8526 (N_8526,N_6586,N_7926);
nand U8527 (N_8527,N_6641,N_6584);
nand U8528 (N_8528,N_7877,N_6013);
nand U8529 (N_8529,N_7632,N_6967);
or U8530 (N_8530,N_7494,N_6162);
xor U8531 (N_8531,N_6718,N_7055);
nor U8532 (N_8532,N_7074,N_7734);
nand U8533 (N_8533,N_7861,N_7478);
and U8534 (N_8534,N_6615,N_7067);
nor U8535 (N_8535,N_7089,N_7952);
nand U8536 (N_8536,N_7167,N_6140);
nand U8537 (N_8537,N_6683,N_6463);
and U8538 (N_8538,N_6338,N_6965);
or U8539 (N_8539,N_6343,N_6234);
or U8540 (N_8540,N_6040,N_7347);
or U8541 (N_8541,N_6752,N_6986);
nor U8542 (N_8542,N_6693,N_6289);
nand U8543 (N_8543,N_6108,N_7377);
nor U8544 (N_8544,N_6563,N_6438);
or U8545 (N_8545,N_6689,N_6516);
nand U8546 (N_8546,N_6393,N_7368);
nand U8547 (N_8547,N_7201,N_6832);
or U8548 (N_8548,N_7273,N_7244);
nand U8549 (N_8549,N_6732,N_6806);
and U8550 (N_8550,N_6520,N_7235);
or U8551 (N_8551,N_6707,N_6956);
and U8552 (N_8552,N_6710,N_7645);
nand U8553 (N_8553,N_6434,N_7961);
and U8554 (N_8554,N_6900,N_7142);
nor U8555 (N_8555,N_7206,N_7173);
and U8556 (N_8556,N_6915,N_7430);
xor U8557 (N_8557,N_7627,N_6047);
and U8558 (N_8558,N_7413,N_7869);
or U8559 (N_8559,N_7605,N_6380);
nor U8560 (N_8560,N_7625,N_7476);
and U8561 (N_8561,N_7762,N_7721);
nand U8562 (N_8562,N_6721,N_6076);
xnor U8563 (N_8563,N_7533,N_7197);
xnor U8564 (N_8564,N_7997,N_7428);
nor U8565 (N_8565,N_6909,N_7234);
nand U8566 (N_8566,N_6505,N_7994);
or U8567 (N_8567,N_7643,N_6131);
and U8568 (N_8568,N_6093,N_6936);
or U8569 (N_8569,N_7126,N_7148);
nor U8570 (N_8570,N_6606,N_6614);
nor U8571 (N_8571,N_6146,N_7090);
and U8572 (N_8572,N_6232,N_7291);
or U8573 (N_8573,N_6367,N_7003);
and U8574 (N_8574,N_7744,N_6604);
nor U8575 (N_8575,N_7193,N_7366);
xor U8576 (N_8576,N_6390,N_6073);
nor U8577 (N_8577,N_7880,N_7517);
nor U8578 (N_8578,N_6691,N_6324);
and U8579 (N_8579,N_6322,N_6253);
xnor U8580 (N_8580,N_7538,N_6887);
and U8581 (N_8581,N_7012,N_7696);
and U8582 (N_8582,N_7578,N_6652);
nand U8583 (N_8583,N_6774,N_6960);
or U8584 (N_8584,N_7573,N_7308);
nor U8585 (N_8585,N_7471,N_7644);
and U8586 (N_8586,N_6024,N_6362);
nand U8587 (N_8587,N_7255,N_6778);
and U8588 (N_8588,N_7467,N_6858);
xor U8589 (N_8589,N_7660,N_6402);
nor U8590 (N_8590,N_6550,N_6276);
nand U8591 (N_8591,N_7986,N_6888);
and U8592 (N_8592,N_7091,N_7455);
and U8593 (N_8593,N_6301,N_6028);
and U8594 (N_8594,N_6859,N_7166);
or U8595 (N_8595,N_6816,N_7188);
and U8596 (N_8596,N_7230,N_7542);
or U8597 (N_8597,N_7767,N_6387);
xor U8598 (N_8598,N_6827,N_6569);
nor U8599 (N_8599,N_6416,N_7980);
or U8600 (N_8600,N_6401,N_7774);
or U8601 (N_8601,N_6442,N_6224);
xnor U8602 (N_8602,N_7433,N_6117);
and U8603 (N_8603,N_6617,N_6547);
nor U8604 (N_8604,N_7272,N_7373);
xnor U8605 (N_8605,N_6045,N_6527);
nor U8606 (N_8606,N_7019,N_6916);
nand U8607 (N_8607,N_7001,N_6934);
nand U8608 (N_8608,N_7884,N_6938);
and U8609 (N_8609,N_6728,N_6034);
nand U8610 (N_8610,N_6049,N_6141);
nor U8611 (N_8611,N_6976,N_7537);
xnor U8612 (N_8612,N_7318,N_7362);
and U8613 (N_8613,N_7354,N_6351);
nand U8614 (N_8614,N_7897,N_6059);
nor U8615 (N_8615,N_6460,N_7440);
nor U8616 (N_8616,N_6383,N_7286);
or U8617 (N_8617,N_7154,N_7082);
nand U8618 (N_8618,N_7740,N_6881);
xor U8619 (N_8619,N_6543,N_6872);
nand U8620 (N_8620,N_7954,N_7328);
and U8621 (N_8621,N_7988,N_6103);
or U8622 (N_8622,N_6374,N_7966);
or U8623 (N_8623,N_7419,N_6585);
and U8624 (N_8624,N_7484,N_6072);
and U8625 (N_8625,N_7071,N_6529);
and U8626 (N_8626,N_7730,N_6799);
or U8627 (N_8627,N_7600,N_6133);
or U8628 (N_8628,N_6422,N_6015);
nor U8629 (N_8629,N_6372,N_7709);
and U8630 (N_8630,N_7631,N_6813);
or U8631 (N_8631,N_6583,N_6735);
or U8632 (N_8632,N_6791,N_7731);
and U8633 (N_8633,N_6871,N_6147);
and U8634 (N_8634,N_7845,N_7491);
nor U8635 (N_8635,N_6878,N_7829);
and U8636 (N_8636,N_6587,N_7360);
xnor U8637 (N_8637,N_6208,N_7621);
nor U8638 (N_8638,N_6192,N_7657);
nor U8639 (N_8639,N_7029,N_7229);
nor U8640 (N_8640,N_7171,N_6896);
and U8641 (N_8641,N_7586,N_7561);
nor U8642 (N_8642,N_7750,N_7781);
nand U8643 (N_8643,N_6623,N_7955);
nand U8644 (N_8644,N_7191,N_6633);
or U8645 (N_8645,N_7251,N_7431);
or U8646 (N_8646,N_6225,N_7449);
and U8647 (N_8647,N_6642,N_6033);
nor U8648 (N_8648,N_6420,N_6650);
and U8649 (N_8649,N_6864,N_6766);
or U8650 (N_8650,N_6899,N_6247);
and U8651 (N_8651,N_7357,N_7679);
nand U8652 (N_8652,N_6835,N_7726);
nor U8653 (N_8653,N_6993,N_7886);
or U8654 (N_8654,N_7697,N_7770);
and U8655 (N_8655,N_6261,N_6963);
nand U8656 (N_8656,N_7868,N_6610);
nor U8657 (N_8657,N_7222,N_6075);
and U8658 (N_8658,N_6601,N_7788);
nand U8659 (N_8659,N_6306,N_6120);
nand U8660 (N_8660,N_6706,N_7451);
nand U8661 (N_8661,N_6589,N_7565);
or U8662 (N_8662,N_7394,N_6473);
xnor U8663 (N_8663,N_7294,N_7735);
or U8664 (N_8664,N_6407,N_6618);
nor U8665 (N_8665,N_6537,N_6083);
nor U8666 (N_8666,N_7816,N_6557);
or U8667 (N_8667,N_7233,N_6546);
xor U8668 (N_8668,N_6819,N_7856);
or U8669 (N_8669,N_6720,N_7076);
and U8670 (N_8670,N_6386,N_7692);
nand U8671 (N_8671,N_7079,N_7486);
or U8672 (N_8672,N_6194,N_7452);
nand U8673 (N_8673,N_6609,N_7678);
nand U8674 (N_8674,N_6310,N_7061);
and U8675 (N_8675,N_7278,N_7337);
and U8676 (N_8676,N_7819,N_7444);
and U8677 (N_8677,N_7442,N_7766);
or U8678 (N_8678,N_6424,N_6729);
nand U8679 (N_8679,N_7146,N_6906);
xor U8680 (N_8680,N_7135,N_7388);
or U8681 (N_8681,N_7036,N_7051);
nand U8682 (N_8682,N_7396,N_6254);
or U8683 (N_8683,N_7249,N_7531);
and U8684 (N_8684,N_6056,N_6637);
or U8685 (N_8685,N_7248,N_7277);
xor U8686 (N_8686,N_6502,N_6129);
nor U8687 (N_8687,N_6591,N_6041);
or U8688 (N_8688,N_6181,N_6189);
nand U8689 (N_8689,N_7835,N_6790);
nor U8690 (N_8690,N_6361,N_6057);
nand U8691 (N_8691,N_6086,N_7239);
and U8692 (N_8692,N_7221,N_6961);
xor U8693 (N_8693,N_7395,N_7528);
or U8694 (N_8694,N_6845,N_7656);
nand U8695 (N_8695,N_6160,N_7551);
or U8696 (N_8696,N_7927,N_7540);
nand U8697 (N_8697,N_7759,N_6470);
nor U8698 (N_8698,N_7105,N_6004);
and U8699 (N_8699,N_7658,N_7775);
nand U8700 (N_8700,N_7382,N_6667);
nand U8701 (N_8701,N_6812,N_7555);
xor U8702 (N_8702,N_6360,N_7502);
nor U8703 (N_8703,N_6715,N_7319);
nor U8704 (N_8704,N_7062,N_6433);
xor U8705 (N_8705,N_7408,N_6127);
or U8706 (N_8706,N_6186,N_7041);
nor U8707 (N_8707,N_7932,N_6211);
xnor U8708 (N_8708,N_7331,N_6758);
nand U8709 (N_8709,N_6395,N_6966);
xor U8710 (N_8710,N_7557,N_7912);
nand U8711 (N_8711,N_7624,N_7777);
or U8712 (N_8712,N_6347,N_7156);
nor U8713 (N_8713,N_7863,N_6528);
or U8714 (N_8714,N_6379,N_7871);
nor U8715 (N_8715,N_7386,N_7620);
and U8716 (N_8716,N_6440,N_6444);
nor U8717 (N_8717,N_6255,N_7133);
nand U8718 (N_8718,N_7793,N_7541);
and U8719 (N_8719,N_7780,N_6156);
nor U8720 (N_8720,N_6299,N_6399);
nand U8721 (N_8721,N_7192,N_7639);
nand U8722 (N_8722,N_7527,N_6901);
nand U8723 (N_8723,N_7577,N_7333);
and U8724 (N_8724,N_7152,N_6800);
nor U8725 (N_8725,N_6283,N_6447);
nand U8726 (N_8726,N_6676,N_7870);
or U8727 (N_8727,N_6932,N_6923);
nand U8728 (N_8728,N_6850,N_7833);
or U8729 (N_8729,N_7681,N_6304);
nand U8730 (N_8730,N_7511,N_7043);
and U8731 (N_8731,N_6426,N_6087);
nor U8732 (N_8732,N_7088,N_7790);
and U8733 (N_8733,N_7268,N_6180);
or U8734 (N_8734,N_6866,N_7822);
nand U8735 (N_8735,N_7077,N_7704);
nor U8736 (N_8736,N_7616,N_7732);
nor U8737 (N_8737,N_6188,N_7223);
and U8738 (N_8738,N_7288,N_7204);
nand U8739 (N_8739,N_6173,N_7663);
or U8740 (N_8740,N_6624,N_7063);
and U8741 (N_8741,N_6559,N_6531);
nor U8742 (N_8742,N_7116,N_6396);
and U8743 (N_8743,N_6066,N_7945);
nor U8744 (N_8744,N_6423,N_6198);
or U8745 (N_8745,N_7275,N_7500);
or U8746 (N_8746,N_7601,N_7417);
and U8747 (N_8747,N_7539,N_6793);
nor U8748 (N_8748,N_7650,N_7526);
nor U8749 (N_8749,N_7757,N_7874);
nor U8750 (N_8750,N_7187,N_7113);
xor U8751 (N_8751,N_7279,N_6085);
or U8752 (N_8752,N_6069,N_6722);
and U8753 (N_8753,N_6937,N_6980);
nor U8754 (N_8754,N_6071,N_7850);
xor U8755 (N_8755,N_6413,N_7844);
and U8756 (N_8756,N_6113,N_6499);
nor U8757 (N_8757,N_7025,N_6947);
nand U8758 (N_8758,N_6968,N_6042);
and U8759 (N_8759,N_7506,N_6570);
nor U8760 (N_8760,N_6209,N_6214);
or U8761 (N_8761,N_7610,N_6168);
nor U8762 (N_8762,N_6521,N_6602);
and U8763 (N_8763,N_7815,N_7896);
nor U8764 (N_8764,N_7684,N_7137);
nor U8765 (N_8765,N_6222,N_7445);
nand U8766 (N_8766,N_6820,N_7949);
nand U8767 (N_8767,N_7619,N_6206);
xor U8768 (N_8768,N_7026,N_6078);
nand U8769 (N_8769,N_6666,N_7630);
nor U8770 (N_8770,N_6783,N_6763);
and U8771 (N_8771,N_7416,N_7372);
and U8772 (N_8772,N_7096,N_6775);
xor U8773 (N_8773,N_7827,N_6340);
or U8774 (N_8774,N_7559,N_7591);
and U8775 (N_8775,N_7981,N_6588);
nor U8776 (N_8776,N_7086,N_6556);
and U8777 (N_8777,N_6719,N_6139);
nand U8778 (N_8778,N_7459,N_7520);
nand U8779 (N_8779,N_6506,N_6029);
and U8780 (N_8780,N_7131,N_6573);
xnor U8781 (N_8781,N_6675,N_7842);
nand U8782 (N_8782,N_6818,N_6930);
nor U8783 (N_8783,N_7033,N_7987);
and U8784 (N_8784,N_7432,N_7421);
and U8785 (N_8785,N_6273,N_6890);
nor U8786 (N_8786,N_7893,N_6481);
nand U8787 (N_8787,N_6630,N_6112);
or U8788 (N_8788,N_7013,N_6308);
and U8789 (N_8789,N_7226,N_7797);
nor U8790 (N_8790,N_7355,N_6373);
nand U8791 (N_8791,N_6544,N_7274);
and U8792 (N_8792,N_7065,N_7544);
nor U8793 (N_8793,N_7567,N_7742);
and U8794 (N_8794,N_7282,N_7109);
or U8795 (N_8795,N_6730,N_6138);
nor U8796 (N_8796,N_6097,N_7647);
or U8797 (N_8797,N_6490,N_7147);
nand U8798 (N_8798,N_6236,N_6326);
nor U8799 (N_8799,N_6997,N_7300);
nor U8800 (N_8800,N_7810,N_6428);
nand U8801 (N_8801,N_6762,N_6260);
or U8802 (N_8802,N_6050,N_6084);
nand U8803 (N_8803,N_7895,N_6696);
and U8804 (N_8804,N_6945,N_6044);
nor U8805 (N_8805,N_6668,N_7346);
xnor U8806 (N_8806,N_7151,N_7120);
nand U8807 (N_8807,N_6269,N_7456);
nand U8808 (N_8808,N_6755,N_6397);
nand U8809 (N_8809,N_7916,N_6337);
and U8810 (N_8810,N_6716,N_6636);
or U8811 (N_8811,N_6114,N_6657);
and U8812 (N_8812,N_7771,N_7124);
xor U8813 (N_8813,N_6183,N_6303);
nand U8814 (N_8814,N_7496,N_6542);
xor U8815 (N_8815,N_7160,N_7094);
nor U8816 (N_8816,N_6182,N_7269);
xnor U8817 (N_8817,N_7575,N_7359);
nor U8818 (N_8818,N_6445,N_6150);
or U8819 (N_8819,N_6469,N_6954);
nand U8820 (N_8820,N_6941,N_7075);
xnor U8821 (N_8821,N_7693,N_6457);
and U8822 (N_8822,N_7353,N_7623);
nor U8823 (N_8823,N_6987,N_7641);
and U8824 (N_8824,N_7149,N_7720);
or U8825 (N_8825,N_6622,N_6664);
or U8826 (N_8826,N_6359,N_7518);
nand U8827 (N_8827,N_6567,N_7855);
nor U8828 (N_8828,N_7768,N_6911);
and U8829 (N_8829,N_7633,N_7975);
nand U8830 (N_8830,N_7939,N_7302);
or U8831 (N_8831,N_7104,N_6669);
nand U8832 (N_8832,N_7891,N_6239);
or U8833 (N_8833,N_7443,N_7859);
nand U8834 (N_8834,N_6898,N_6171);
or U8835 (N_8835,N_6284,N_7400);
xnor U8836 (N_8836,N_7338,N_6925);
and U8837 (N_8837,N_7700,N_6003);
and U8838 (N_8838,N_6984,N_7552);
and U8839 (N_8839,N_7371,N_6507);
nor U8840 (N_8840,N_6296,N_7011);
nand U8841 (N_8841,N_7422,N_7743);
or U8842 (N_8842,N_7314,N_7642);
nor U8843 (N_8843,N_6339,N_7615);
or U8844 (N_8844,N_6471,N_6643);
nand U8845 (N_8845,N_6126,N_7068);
or U8846 (N_8846,N_6504,N_7901);
and U8847 (N_8847,N_7298,N_7461);
and U8848 (N_8848,N_7106,N_6842);
nor U8849 (N_8849,N_6332,N_7048);
and U8850 (N_8850,N_6476,N_6532);
and U8851 (N_8851,N_7809,N_7436);
and U8852 (N_8852,N_6262,N_7306);
nand U8853 (N_8853,N_7830,N_6985);
xor U8854 (N_8854,N_7898,N_6105);
nand U8855 (N_8855,N_6278,N_6144);
nor U8856 (N_8856,N_7038,N_7183);
and U8857 (N_8857,N_6464,N_7006);
and U8858 (N_8858,N_6734,N_7084);
nand U8859 (N_8859,N_7097,N_7710);
or U8860 (N_8860,N_6680,N_7728);
xor U8861 (N_8861,N_7854,N_7515);
nand U8862 (N_8862,N_7792,N_7004);
and U8863 (N_8863,N_6995,N_6523);
nor U8864 (N_8864,N_6549,N_6841);
and U8865 (N_8865,N_7335,N_7529);
and U8866 (N_8866,N_7938,N_6456);
nand U8867 (N_8867,N_6363,N_7242);
or U8868 (N_8868,N_7651,N_7685);
and U8869 (N_8869,N_7677,N_6307);
nor U8870 (N_8870,N_6757,N_7399);
nor U8871 (N_8871,N_6875,N_7332);
and U8872 (N_8872,N_6427,N_6678);
or U8873 (N_8873,N_6698,N_7121);
or U8874 (N_8874,N_7760,N_6290);
or U8875 (N_8875,N_6279,N_7563);
and U8876 (N_8876,N_6252,N_7344);
and U8877 (N_8877,N_6773,N_6921);
or U8878 (N_8878,N_6039,N_7546);
nor U8879 (N_8879,N_7429,N_6830);
or U8880 (N_8880,N_6861,N_7172);
and U8881 (N_8881,N_7042,N_7749);
nand U8882 (N_8882,N_7483,N_7093);
nand U8883 (N_8883,N_7078,N_7674);
nor U8884 (N_8884,N_6314,N_6885);
or U8885 (N_8885,N_6903,N_6455);
nand U8886 (N_8886,N_6280,N_7761);
nor U8887 (N_8887,N_7910,N_6498);
nor U8888 (N_8888,N_6877,N_6124);
xnor U8889 (N_8889,N_6904,N_6345);
or U8890 (N_8890,N_6682,N_7924);
nand U8891 (N_8891,N_7991,N_7305);
xnor U8892 (N_8892,N_7446,N_7283);
and U8893 (N_8893,N_6862,N_7543);
or U8894 (N_8894,N_7769,N_6646);
nand U8895 (N_8895,N_7210,N_7576);
nand U8896 (N_8896,N_7037,N_7963);
nand U8897 (N_8897,N_7475,N_6092);
and U8898 (N_8898,N_7228,N_7883);
or U8899 (N_8899,N_6418,N_6135);
and U8900 (N_8900,N_6625,N_7872);
and U8901 (N_8901,N_6649,N_6939);
nor U8902 (N_8902,N_7521,N_7524);
nand U8903 (N_8903,N_7580,N_7209);
nand U8904 (N_8904,N_7672,N_6241);
nor U8905 (N_8905,N_7652,N_6612);
or U8906 (N_8906,N_6240,N_7534);
xor U8907 (N_8907,N_6486,N_7186);
and U8908 (N_8908,N_6955,N_7008);
nor U8909 (N_8909,N_6685,N_7717);
xor U8910 (N_8910,N_7608,N_6974);
or U8911 (N_8911,N_6651,N_6348);
nor U8912 (N_8912,N_6210,N_6479);
nand U8913 (N_8913,N_7317,N_6928);
and U8914 (N_8914,N_7727,N_6352);
and U8915 (N_8915,N_6305,N_7296);
nand U8916 (N_8916,N_6750,N_6654);
xnor U8917 (N_8917,N_6357,N_7536);
nand U8918 (N_8918,N_7289,N_6607);
nor U8919 (N_8919,N_6565,N_6500);
nor U8920 (N_8920,N_6777,N_6568);
xor U8921 (N_8921,N_7370,N_6494);
or U8922 (N_8922,N_7569,N_6803);
nor U8923 (N_8923,N_6067,N_7796);
xor U8924 (N_8924,N_7773,N_6638);
nor U8925 (N_8925,N_6705,N_7902);
nand U8926 (N_8926,N_6414,N_7807);
or U8927 (N_8927,N_7380,N_6153);
or U8928 (N_8928,N_6165,N_6834);
nor U8929 (N_8929,N_6237,N_7295);
or U8930 (N_8930,N_7804,N_7341);
nor U8931 (N_8931,N_7613,N_7217);
xor U8932 (N_8932,N_6090,N_6495);
xor U8933 (N_8933,N_7668,N_6030);
or U8934 (N_8934,N_6548,N_6074);
nand U8935 (N_8935,N_7010,N_7313);
or U8936 (N_8936,N_6635,N_7698);
and U8937 (N_8937,N_7935,N_7834);
or U8938 (N_8938,N_7670,N_6331);
nand U8939 (N_8939,N_7303,N_7007);
and U8940 (N_8940,N_7847,N_7646);
and U8941 (N_8941,N_7336,N_7965);
nand U8942 (N_8942,N_7411,N_6392);
nand U8943 (N_8943,N_7911,N_6497);
and U8944 (N_8944,N_6291,N_7263);
or U8945 (N_8945,N_6195,N_7851);
nand U8946 (N_8946,N_7929,N_6535);
and U8947 (N_8947,N_7307,N_7092);
or U8948 (N_8948,N_6751,N_6805);
and U8949 (N_8949,N_7866,N_6558);
and U8950 (N_8950,N_6425,N_7111);
or U8951 (N_8951,N_6754,N_6902);
nand U8952 (N_8952,N_6692,N_6807);
nand U8953 (N_8953,N_6242,N_6302);
nand U8954 (N_8954,N_6264,N_6613);
nand U8955 (N_8955,N_6109,N_7659);
or U8956 (N_8956,N_7805,N_7311);
and U8957 (N_8957,N_6776,N_7504);
or U8958 (N_8958,N_6403,N_7081);
xnor U8959 (N_8959,N_6054,N_7746);
or U8960 (N_8960,N_7356,N_6946);
and U8961 (N_8961,N_6477,N_7136);
xnor U8962 (N_8962,N_7811,N_6789);
xor U8963 (N_8963,N_6554,N_6714);
and U8964 (N_8964,N_7867,N_7971);
nor U8965 (N_8965,N_7516,N_6110);
or U8966 (N_8966,N_6592,N_6051);
nand U8967 (N_8967,N_7184,N_6748);
nand U8968 (N_8968,N_7321,N_6480);
nor U8969 (N_8969,N_6959,N_6713);
nand U8970 (N_8970,N_7246,N_6061);
or U8971 (N_8971,N_7733,N_6578);
nor U8972 (N_8972,N_6388,N_6368);
and U8973 (N_8973,N_6459,N_7219);
xor U8974 (N_8974,N_6268,N_7342);
xnor U8975 (N_8975,N_7265,N_6905);
and U8976 (N_8976,N_7207,N_7687);
or U8977 (N_8977,N_7107,N_7838);
nor U8978 (N_8978,N_7287,N_7508);
nand U8979 (N_8979,N_6228,N_7213);
nand U8980 (N_8980,N_7103,N_6107);
nor U8981 (N_8981,N_6541,N_6330);
xor U8982 (N_8982,N_6406,N_7890);
nand U8983 (N_8983,N_7931,N_6412);
nor U8984 (N_8984,N_7794,N_7928);
or U8985 (N_8985,N_7879,N_7595);
xor U8986 (N_8986,N_7474,N_7535);
and U8987 (N_8987,N_7224,N_7914);
or U8988 (N_8988,N_6595,N_6724);
nor U8989 (N_8989,N_7998,N_7211);
or U8990 (N_8990,N_7801,N_6975);
xor U8991 (N_8991,N_6593,N_7813);
nor U8992 (N_8992,N_6488,N_7594);
nor U8993 (N_8993,N_6104,N_7748);
or U8994 (N_8994,N_6561,N_6894);
nand U8995 (N_8995,N_6663,N_7472);
nor U8996 (N_8996,N_7423,N_6274);
and U8997 (N_8997,N_7799,N_6309);
and U8998 (N_8998,N_7705,N_6152);
nor U8999 (N_8999,N_7634,N_7977);
or U9000 (N_9000,N_7242,N_6734);
or U9001 (N_9001,N_6063,N_7491);
nand U9002 (N_9002,N_6857,N_6682);
and U9003 (N_9003,N_7944,N_6944);
nand U9004 (N_9004,N_7103,N_6183);
and U9005 (N_9005,N_7860,N_7981);
nand U9006 (N_9006,N_6365,N_7060);
nand U9007 (N_9007,N_6010,N_7633);
nor U9008 (N_9008,N_6753,N_6418);
or U9009 (N_9009,N_6057,N_7537);
nand U9010 (N_9010,N_7340,N_6062);
nor U9011 (N_9011,N_7697,N_6112);
nand U9012 (N_9012,N_7297,N_6306);
and U9013 (N_9013,N_6375,N_6614);
nand U9014 (N_9014,N_7445,N_7263);
nand U9015 (N_9015,N_7276,N_6234);
nand U9016 (N_9016,N_6065,N_6838);
or U9017 (N_9017,N_7856,N_7371);
nand U9018 (N_9018,N_6125,N_7142);
or U9019 (N_9019,N_6674,N_7516);
nor U9020 (N_9020,N_6397,N_6453);
or U9021 (N_9021,N_6672,N_7017);
xnor U9022 (N_9022,N_7963,N_6773);
or U9023 (N_9023,N_6941,N_6790);
or U9024 (N_9024,N_7533,N_6086);
and U9025 (N_9025,N_7626,N_7226);
nand U9026 (N_9026,N_6469,N_6241);
xor U9027 (N_9027,N_6187,N_7754);
nor U9028 (N_9028,N_7123,N_6902);
nor U9029 (N_9029,N_7150,N_7031);
and U9030 (N_9030,N_6395,N_6634);
or U9031 (N_9031,N_7584,N_6815);
nor U9032 (N_9032,N_6530,N_6907);
or U9033 (N_9033,N_7076,N_6944);
and U9034 (N_9034,N_6450,N_6863);
nand U9035 (N_9035,N_6786,N_6402);
or U9036 (N_9036,N_6443,N_7949);
nand U9037 (N_9037,N_6195,N_7100);
nor U9038 (N_9038,N_7378,N_6475);
and U9039 (N_9039,N_6190,N_6831);
or U9040 (N_9040,N_6623,N_7349);
nor U9041 (N_9041,N_7316,N_6906);
xor U9042 (N_9042,N_6465,N_7392);
nor U9043 (N_9043,N_6458,N_7560);
or U9044 (N_9044,N_7619,N_6719);
nor U9045 (N_9045,N_7768,N_7659);
nand U9046 (N_9046,N_7289,N_7326);
and U9047 (N_9047,N_6136,N_6183);
nor U9048 (N_9048,N_6392,N_6833);
nor U9049 (N_9049,N_7625,N_6525);
or U9050 (N_9050,N_6187,N_7024);
and U9051 (N_9051,N_6664,N_6579);
or U9052 (N_9052,N_6049,N_6517);
or U9053 (N_9053,N_6424,N_6655);
xnor U9054 (N_9054,N_6653,N_6162);
or U9055 (N_9055,N_6550,N_6425);
nor U9056 (N_9056,N_7818,N_6562);
xor U9057 (N_9057,N_7443,N_6839);
or U9058 (N_9058,N_6815,N_6640);
and U9059 (N_9059,N_6587,N_7582);
or U9060 (N_9060,N_6603,N_6501);
nor U9061 (N_9061,N_6587,N_6743);
nor U9062 (N_9062,N_6811,N_6596);
nor U9063 (N_9063,N_6723,N_7915);
nor U9064 (N_9064,N_7954,N_7167);
and U9065 (N_9065,N_7886,N_7571);
nand U9066 (N_9066,N_7278,N_7676);
nor U9067 (N_9067,N_6845,N_6933);
nor U9068 (N_9068,N_7648,N_6853);
and U9069 (N_9069,N_7180,N_6857);
and U9070 (N_9070,N_6494,N_6842);
or U9071 (N_9071,N_7663,N_7405);
and U9072 (N_9072,N_7952,N_7765);
nor U9073 (N_9073,N_7993,N_6016);
nor U9074 (N_9074,N_7355,N_6923);
or U9075 (N_9075,N_7871,N_6640);
and U9076 (N_9076,N_6743,N_6464);
and U9077 (N_9077,N_6771,N_7634);
nor U9078 (N_9078,N_6260,N_7965);
nand U9079 (N_9079,N_6663,N_7338);
nand U9080 (N_9080,N_6194,N_7875);
or U9081 (N_9081,N_7980,N_6573);
nand U9082 (N_9082,N_6359,N_6731);
and U9083 (N_9083,N_7416,N_6749);
and U9084 (N_9084,N_6375,N_7381);
nor U9085 (N_9085,N_7688,N_7623);
or U9086 (N_9086,N_7364,N_7377);
and U9087 (N_9087,N_6105,N_7767);
nor U9088 (N_9088,N_6241,N_7902);
nand U9089 (N_9089,N_6609,N_6697);
or U9090 (N_9090,N_6768,N_6467);
nand U9091 (N_9091,N_6388,N_7809);
nor U9092 (N_9092,N_6601,N_7905);
xor U9093 (N_9093,N_6474,N_7852);
or U9094 (N_9094,N_6645,N_7623);
or U9095 (N_9095,N_7723,N_7300);
and U9096 (N_9096,N_6565,N_6632);
nor U9097 (N_9097,N_6560,N_6512);
nor U9098 (N_9098,N_6238,N_6916);
and U9099 (N_9099,N_7057,N_7960);
or U9100 (N_9100,N_7222,N_7084);
xnor U9101 (N_9101,N_7401,N_6580);
xor U9102 (N_9102,N_7543,N_6367);
nand U9103 (N_9103,N_7412,N_6851);
or U9104 (N_9104,N_6342,N_7763);
nand U9105 (N_9105,N_6290,N_6554);
nor U9106 (N_9106,N_6010,N_6348);
xnor U9107 (N_9107,N_7936,N_6227);
or U9108 (N_9108,N_7395,N_7916);
nor U9109 (N_9109,N_6994,N_7187);
nor U9110 (N_9110,N_6108,N_6478);
nand U9111 (N_9111,N_7903,N_7445);
xor U9112 (N_9112,N_6747,N_6741);
nand U9113 (N_9113,N_7395,N_7660);
or U9114 (N_9114,N_6055,N_6620);
and U9115 (N_9115,N_7256,N_6101);
and U9116 (N_9116,N_7036,N_7422);
nor U9117 (N_9117,N_6037,N_7062);
xnor U9118 (N_9118,N_7194,N_7856);
and U9119 (N_9119,N_6327,N_6480);
nand U9120 (N_9120,N_7365,N_7922);
and U9121 (N_9121,N_7396,N_6034);
nand U9122 (N_9122,N_7092,N_7783);
nor U9123 (N_9123,N_6223,N_7216);
or U9124 (N_9124,N_6860,N_6563);
xnor U9125 (N_9125,N_6699,N_6874);
and U9126 (N_9126,N_7639,N_6353);
nand U9127 (N_9127,N_7889,N_6560);
and U9128 (N_9128,N_6486,N_7317);
xnor U9129 (N_9129,N_6653,N_6431);
nand U9130 (N_9130,N_6856,N_6172);
nor U9131 (N_9131,N_6539,N_6278);
or U9132 (N_9132,N_7716,N_6632);
or U9133 (N_9133,N_7810,N_6550);
xor U9134 (N_9134,N_7479,N_6508);
xor U9135 (N_9135,N_6862,N_7443);
and U9136 (N_9136,N_7498,N_7890);
nand U9137 (N_9137,N_6776,N_6654);
xor U9138 (N_9138,N_6195,N_6775);
nand U9139 (N_9139,N_6694,N_6760);
nand U9140 (N_9140,N_7165,N_7185);
nand U9141 (N_9141,N_6842,N_7905);
nand U9142 (N_9142,N_6655,N_6323);
nor U9143 (N_9143,N_7400,N_7064);
or U9144 (N_9144,N_6176,N_7483);
nand U9145 (N_9145,N_7338,N_7494);
and U9146 (N_9146,N_6557,N_7314);
or U9147 (N_9147,N_7377,N_7903);
nor U9148 (N_9148,N_6844,N_6825);
nand U9149 (N_9149,N_7379,N_6122);
or U9150 (N_9150,N_7506,N_7522);
nor U9151 (N_9151,N_6435,N_7819);
nand U9152 (N_9152,N_7527,N_7335);
nor U9153 (N_9153,N_6309,N_7835);
or U9154 (N_9154,N_7359,N_7881);
nand U9155 (N_9155,N_7574,N_7043);
nand U9156 (N_9156,N_7097,N_6483);
and U9157 (N_9157,N_6250,N_7313);
or U9158 (N_9158,N_7190,N_6121);
or U9159 (N_9159,N_6038,N_6899);
and U9160 (N_9160,N_6477,N_6733);
or U9161 (N_9161,N_6889,N_7227);
nor U9162 (N_9162,N_7402,N_6671);
nor U9163 (N_9163,N_6884,N_7082);
xor U9164 (N_9164,N_6851,N_6948);
or U9165 (N_9165,N_6144,N_6868);
nor U9166 (N_9166,N_7890,N_7952);
nor U9167 (N_9167,N_7660,N_6893);
and U9168 (N_9168,N_6285,N_6764);
or U9169 (N_9169,N_6528,N_7014);
or U9170 (N_9170,N_7906,N_7522);
or U9171 (N_9171,N_7265,N_6134);
and U9172 (N_9172,N_7896,N_7865);
nor U9173 (N_9173,N_7979,N_7706);
or U9174 (N_9174,N_7001,N_7129);
nor U9175 (N_9175,N_7951,N_6815);
and U9176 (N_9176,N_7872,N_7209);
nand U9177 (N_9177,N_6159,N_7335);
nor U9178 (N_9178,N_6922,N_6166);
nor U9179 (N_9179,N_7816,N_6903);
nand U9180 (N_9180,N_6439,N_6651);
nor U9181 (N_9181,N_7874,N_7679);
nor U9182 (N_9182,N_7118,N_7879);
or U9183 (N_9183,N_7965,N_6437);
nor U9184 (N_9184,N_7288,N_6300);
or U9185 (N_9185,N_6493,N_6580);
nand U9186 (N_9186,N_6196,N_6142);
or U9187 (N_9187,N_7688,N_7572);
and U9188 (N_9188,N_6247,N_6413);
and U9189 (N_9189,N_7016,N_7272);
nand U9190 (N_9190,N_7497,N_7294);
nand U9191 (N_9191,N_6399,N_6440);
or U9192 (N_9192,N_6701,N_7043);
xor U9193 (N_9193,N_7847,N_6730);
nor U9194 (N_9194,N_6240,N_6975);
xor U9195 (N_9195,N_7144,N_6395);
nand U9196 (N_9196,N_7343,N_7099);
and U9197 (N_9197,N_7777,N_6441);
or U9198 (N_9198,N_7356,N_7599);
nor U9199 (N_9199,N_7892,N_7674);
and U9200 (N_9200,N_6835,N_6723);
and U9201 (N_9201,N_6791,N_7940);
xor U9202 (N_9202,N_6776,N_6999);
and U9203 (N_9203,N_7331,N_7417);
nor U9204 (N_9204,N_6996,N_6468);
xnor U9205 (N_9205,N_7132,N_6566);
nor U9206 (N_9206,N_7875,N_6415);
nand U9207 (N_9207,N_7218,N_7244);
nand U9208 (N_9208,N_7600,N_6360);
nand U9209 (N_9209,N_7710,N_7548);
nor U9210 (N_9210,N_7145,N_6803);
nor U9211 (N_9211,N_7677,N_7484);
nor U9212 (N_9212,N_7071,N_6439);
nor U9213 (N_9213,N_7138,N_7454);
nand U9214 (N_9214,N_7849,N_6704);
and U9215 (N_9215,N_7737,N_7443);
xnor U9216 (N_9216,N_6486,N_6141);
or U9217 (N_9217,N_7206,N_6989);
nand U9218 (N_9218,N_6869,N_6312);
nor U9219 (N_9219,N_6939,N_6775);
and U9220 (N_9220,N_7480,N_6946);
nand U9221 (N_9221,N_7432,N_6166);
or U9222 (N_9222,N_7845,N_6682);
nor U9223 (N_9223,N_7616,N_6362);
nor U9224 (N_9224,N_7970,N_7738);
nand U9225 (N_9225,N_6574,N_6367);
nor U9226 (N_9226,N_6302,N_6944);
or U9227 (N_9227,N_7373,N_6625);
nor U9228 (N_9228,N_6839,N_6017);
nor U9229 (N_9229,N_7970,N_7002);
or U9230 (N_9230,N_6178,N_6025);
xnor U9231 (N_9231,N_7755,N_6122);
nand U9232 (N_9232,N_6361,N_6598);
and U9233 (N_9233,N_6916,N_6072);
nor U9234 (N_9234,N_7736,N_6592);
or U9235 (N_9235,N_7685,N_6024);
and U9236 (N_9236,N_7472,N_6178);
nand U9237 (N_9237,N_6334,N_7565);
nor U9238 (N_9238,N_6992,N_7948);
and U9239 (N_9239,N_7829,N_6409);
nand U9240 (N_9240,N_6060,N_6281);
and U9241 (N_9241,N_7574,N_6098);
nand U9242 (N_9242,N_7816,N_7346);
or U9243 (N_9243,N_6906,N_6581);
and U9244 (N_9244,N_6604,N_7790);
and U9245 (N_9245,N_7963,N_7992);
or U9246 (N_9246,N_7192,N_6666);
nor U9247 (N_9247,N_6370,N_6189);
or U9248 (N_9248,N_7756,N_7120);
or U9249 (N_9249,N_7357,N_7110);
xnor U9250 (N_9250,N_6661,N_6974);
xnor U9251 (N_9251,N_6858,N_7153);
nor U9252 (N_9252,N_6539,N_7830);
nand U9253 (N_9253,N_6777,N_6805);
and U9254 (N_9254,N_7615,N_7113);
nand U9255 (N_9255,N_7565,N_7924);
or U9256 (N_9256,N_7042,N_7502);
xnor U9257 (N_9257,N_7464,N_6421);
or U9258 (N_9258,N_7203,N_6554);
and U9259 (N_9259,N_7827,N_7189);
or U9260 (N_9260,N_6833,N_7115);
nor U9261 (N_9261,N_6877,N_7533);
nand U9262 (N_9262,N_6606,N_6245);
nand U9263 (N_9263,N_6492,N_6570);
xnor U9264 (N_9264,N_7243,N_6829);
or U9265 (N_9265,N_6741,N_7349);
or U9266 (N_9266,N_7226,N_7910);
and U9267 (N_9267,N_7681,N_6156);
and U9268 (N_9268,N_6574,N_6072);
or U9269 (N_9269,N_6670,N_6007);
nand U9270 (N_9270,N_6912,N_6131);
and U9271 (N_9271,N_7857,N_7591);
nor U9272 (N_9272,N_6678,N_7840);
nand U9273 (N_9273,N_6601,N_6299);
or U9274 (N_9274,N_6143,N_6523);
or U9275 (N_9275,N_7335,N_7008);
and U9276 (N_9276,N_6281,N_7619);
xnor U9277 (N_9277,N_7642,N_6181);
and U9278 (N_9278,N_6787,N_6808);
or U9279 (N_9279,N_6877,N_7765);
nand U9280 (N_9280,N_6839,N_6910);
and U9281 (N_9281,N_6009,N_6000);
nand U9282 (N_9282,N_6932,N_6415);
nor U9283 (N_9283,N_6015,N_7554);
nor U9284 (N_9284,N_7175,N_6152);
and U9285 (N_9285,N_6845,N_6549);
or U9286 (N_9286,N_7590,N_6553);
and U9287 (N_9287,N_7722,N_7024);
nor U9288 (N_9288,N_6887,N_6260);
and U9289 (N_9289,N_7513,N_7790);
and U9290 (N_9290,N_7238,N_6065);
nor U9291 (N_9291,N_7077,N_6484);
nand U9292 (N_9292,N_6128,N_6392);
or U9293 (N_9293,N_7629,N_6662);
xnor U9294 (N_9294,N_6940,N_7323);
nor U9295 (N_9295,N_6830,N_6286);
nand U9296 (N_9296,N_6420,N_6128);
and U9297 (N_9297,N_6283,N_7866);
and U9298 (N_9298,N_7064,N_7300);
nor U9299 (N_9299,N_6676,N_7284);
and U9300 (N_9300,N_7647,N_6742);
nor U9301 (N_9301,N_7000,N_7657);
nor U9302 (N_9302,N_6569,N_6055);
xnor U9303 (N_9303,N_7184,N_6935);
or U9304 (N_9304,N_6989,N_7544);
or U9305 (N_9305,N_7811,N_6945);
or U9306 (N_9306,N_6034,N_6892);
or U9307 (N_9307,N_7418,N_7542);
and U9308 (N_9308,N_7388,N_7776);
and U9309 (N_9309,N_6414,N_7774);
and U9310 (N_9310,N_6369,N_7938);
nand U9311 (N_9311,N_6730,N_6459);
and U9312 (N_9312,N_7909,N_6902);
nand U9313 (N_9313,N_6031,N_6483);
nor U9314 (N_9314,N_6912,N_6481);
or U9315 (N_9315,N_7198,N_6203);
nand U9316 (N_9316,N_6303,N_6810);
nor U9317 (N_9317,N_7740,N_7773);
nand U9318 (N_9318,N_7360,N_6090);
nor U9319 (N_9319,N_7954,N_6274);
xnor U9320 (N_9320,N_7297,N_7964);
and U9321 (N_9321,N_6284,N_7243);
nor U9322 (N_9322,N_6969,N_7565);
nor U9323 (N_9323,N_7860,N_7498);
nand U9324 (N_9324,N_6920,N_6219);
nand U9325 (N_9325,N_6856,N_6779);
and U9326 (N_9326,N_6196,N_6673);
and U9327 (N_9327,N_6612,N_6159);
or U9328 (N_9328,N_6550,N_7899);
xor U9329 (N_9329,N_7806,N_6197);
and U9330 (N_9330,N_6654,N_7851);
or U9331 (N_9331,N_7191,N_7825);
or U9332 (N_9332,N_7207,N_6770);
or U9333 (N_9333,N_7331,N_7948);
xnor U9334 (N_9334,N_6570,N_6506);
xnor U9335 (N_9335,N_7518,N_7887);
nor U9336 (N_9336,N_7476,N_7528);
or U9337 (N_9337,N_7591,N_6975);
nor U9338 (N_9338,N_7631,N_6369);
nand U9339 (N_9339,N_6619,N_7689);
xnor U9340 (N_9340,N_6059,N_6727);
nand U9341 (N_9341,N_7127,N_7024);
nand U9342 (N_9342,N_7856,N_7000);
nand U9343 (N_9343,N_6520,N_6074);
xor U9344 (N_9344,N_7432,N_7651);
and U9345 (N_9345,N_6014,N_7999);
or U9346 (N_9346,N_7903,N_6495);
or U9347 (N_9347,N_7500,N_6868);
or U9348 (N_9348,N_6198,N_7661);
and U9349 (N_9349,N_7430,N_7660);
or U9350 (N_9350,N_7284,N_6030);
and U9351 (N_9351,N_6020,N_6795);
or U9352 (N_9352,N_7027,N_7067);
xnor U9353 (N_9353,N_6662,N_6614);
or U9354 (N_9354,N_6722,N_6547);
xnor U9355 (N_9355,N_6154,N_7983);
and U9356 (N_9356,N_6914,N_6308);
or U9357 (N_9357,N_6710,N_7840);
nor U9358 (N_9358,N_7187,N_7564);
or U9359 (N_9359,N_7757,N_7979);
and U9360 (N_9360,N_7906,N_7014);
xnor U9361 (N_9361,N_7958,N_6223);
or U9362 (N_9362,N_6243,N_7709);
and U9363 (N_9363,N_6746,N_6266);
or U9364 (N_9364,N_6831,N_6070);
nand U9365 (N_9365,N_6628,N_6252);
nor U9366 (N_9366,N_7190,N_7890);
nor U9367 (N_9367,N_7603,N_7540);
xnor U9368 (N_9368,N_7260,N_6898);
and U9369 (N_9369,N_7802,N_6598);
and U9370 (N_9370,N_7753,N_6279);
or U9371 (N_9371,N_6995,N_6412);
nand U9372 (N_9372,N_7329,N_7330);
nor U9373 (N_9373,N_7649,N_6444);
nand U9374 (N_9374,N_7617,N_7294);
xor U9375 (N_9375,N_6906,N_6754);
and U9376 (N_9376,N_6390,N_6951);
nand U9377 (N_9377,N_7203,N_7271);
nor U9378 (N_9378,N_7270,N_7081);
and U9379 (N_9379,N_6767,N_6210);
or U9380 (N_9380,N_6596,N_7320);
nor U9381 (N_9381,N_6892,N_7964);
or U9382 (N_9382,N_6303,N_6377);
or U9383 (N_9383,N_6692,N_6505);
nand U9384 (N_9384,N_6758,N_6667);
and U9385 (N_9385,N_7957,N_7075);
xor U9386 (N_9386,N_7726,N_7336);
nand U9387 (N_9387,N_7359,N_6189);
or U9388 (N_9388,N_6338,N_6733);
nor U9389 (N_9389,N_7045,N_6131);
or U9390 (N_9390,N_6875,N_6038);
and U9391 (N_9391,N_6622,N_6738);
nand U9392 (N_9392,N_7627,N_6213);
nand U9393 (N_9393,N_7404,N_7666);
and U9394 (N_9394,N_6507,N_7643);
or U9395 (N_9395,N_6122,N_6161);
nand U9396 (N_9396,N_6089,N_7944);
and U9397 (N_9397,N_7470,N_7511);
nor U9398 (N_9398,N_7448,N_6618);
nand U9399 (N_9399,N_7393,N_6125);
and U9400 (N_9400,N_6469,N_6294);
and U9401 (N_9401,N_7746,N_7802);
nand U9402 (N_9402,N_6102,N_7061);
nor U9403 (N_9403,N_7079,N_7455);
nor U9404 (N_9404,N_6615,N_7501);
and U9405 (N_9405,N_7677,N_6072);
nor U9406 (N_9406,N_7970,N_7047);
and U9407 (N_9407,N_6529,N_6837);
and U9408 (N_9408,N_7638,N_6600);
and U9409 (N_9409,N_6242,N_6067);
and U9410 (N_9410,N_7827,N_7927);
and U9411 (N_9411,N_6952,N_7945);
and U9412 (N_9412,N_6163,N_6169);
nand U9413 (N_9413,N_7819,N_6677);
xnor U9414 (N_9414,N_7510,N_6447);
or U9415 (N_9415,N_6591,N_6977);
and U9416 (N_9416,N_6309,N_7072);
nand U9417 (N_9417,N_7853,N_6027);
nand U9418 (N_9418,N_7249,N_7796);
and U9419 (N_9419,N_6509,N_6364);
nand U9420 (N_9420,N_7872,N_6120);
or U9421 (N_9421,N_7116,N_6382);
nand U9422 (N_9422,N_7910,N_6078);
or U9423 (N_9423,N_7899,N_6050);
nor U9424 (N_9424,N_7256,N_7400);
nor U9425 (N_9425,N_7007,N_6735);
and U9426 (N_9426,N_6062,N_7608);
and U9427 (N_9427,N_6858,N_7076);
nand U9428 (N_9428,N_7336,N_6339);
nand U9429 (N_9429,N_7213,N_6565);
and U9430 (N_9430,N_7773,N_7006);
or U9431 (N_9431,N_6541,N_7041);
and U9432 (N_9432,N_6329,N_6167);
or U9433 (N_9433,N_6610,N_7742);
or U9434 (N_9434,N_7997,N_7195);
or U9435 (N_9435,N_6512,N_7844);
or U9436 (N_9436,N_6188,N_7133);
nor U9437 (N_9437,N_7484,N_7794);
nor U9438 (N_9438,N_7874,N_6125);
nor U9439 (N_9439,N_6865,N_7342);
nand U9440 (N_9440,N_7201,N_6106);
and U9441 (N_9441,N_6168,N_7465);
nand U9442 (N_9442,N_7806,N_7589);
and U9443 (N_9443,N_7766,N_6841);
xnor U9444 (N_9444,N_7849,N_6435);
nand U9445 (N_9445,N_7562,N_7055);
or U9446 (N_9446,N_7470,N_7711);
nand U9447 (N_9447,N_6114,N_6191);
or U9448 (N_9448,N_7430,N_7906);
and U9449 (N_9449,N_7649,N_6196);
nor U9450 (N_9450,N_7480,N_7519);
nand U9451 (N_9451,N_7994,N_6055);
nand U9452 (N_9452,N_7165,N_7040);
and U9453 (N_9453,N_7036,N_7847);
or U9454 (N_9454,N_6710,N_7506);
nor U9455 (N_9455,N_7064,N_6030);
or U9456 (N_9456,N_7920,N_7772);
and U9457 (N_9457,N_7064,N_7915);
nor U9458 (N_9458,N_7858,N_6498);
nor U9459 (N_9459,N_6718,N_6037);
nand U9460 (N_9460,N_6500,N_6615);
nand U9461 (N_9461,N_6966,N_7948);
or U9462 (N_9462,N_7385,N_6834);
and U9463 (N_9463,N_6930,N_6775);
nor U9464 (N_9464,N_6284,N_7618);
or U9465 (N_9465,N_7494,N_6002);
and U9466 (N_9466,N_6191,N_6233);
and U9467 (N_9467,N_6214,N_6943);
nand U9468 (N_9468,N_7960,N_7514);
xor U9469 (N_9469,N_6265,N_7791);
nand U9470 (N_9470,N_7255,N_6544);
or U9471 (N_9471,N_7246,N_7348);
and U9472 (N_9472,N_7232,N_6513);
xor U9473 (N_9473,N_7127,N_6952);
or U9474 (N_9474,N_6427,N_7215);
nand U9475 (N_9475,N_7182,N_6975);
or U9476 (N_9476,N_6357,N_7170);
nand U9477 (N_9477,N_7240,N_7931);
and U9478 (N_9478,N_7396,N_6965);
or U9479 (N_9479,N_6604,N_7138);
xnor U9480 (N_9480,N_7329,N_7867);
and U9481 (N_9481,N_6623,N_7492);
nor U9482 (N_9482,N_6209,N_6676);
and U9483 (N_9483,N_6301,N_7548);
nor U9484 (N_9484,N_6917,N_6086);
xor U9485 (N_9485,N_7778,N_7427);
nand U9486 (N_9486,N_6648,N_7684);
nor U9487 (N_9487,N_6977,N_7766);
nand U9488 (N_9488,N_7686,N_6019);
xor U9489 (N_9489,N_6372,N_7001);
and U9490 (N_9490,N_7455,N_6129);
or U9491 (N_9491,N_7721,N_6405);
and U9492 (N_9492,N_7741,N_6247);
nand U9493 (N_9493,N_6799,N_7655);
xnor U9494 (N_9494,N_6801,N_6994);
and U9495 (N_9495,N_6679,N_6259);
or U9496 (N_9496,N_7410,N_6853);
nand U9497 (N_9497,N_7972,N_7641);
xnor U9498 (N_9498,N_6248,N_7049);
xnor U9499 (N_9499,N_7402,N_7789);
or U9500 (N_9500,N_7782,N_6582);
or U9501 (N_9501,N_6827,N_6608);
and U9502 (N_9502,N_7445,N_6640);
nand U9503 (N_9503,N_6976,N_6772);
nand U9504 (N_9504,N_6544,N_7957);
or U9505 (N_9505,N_7973,N_6816);
nand U9506 (N_9506,N_6029,N_7513);
nand U9507 (N_9507,N_7728,N_6397);
nand U9508 (N_9508,N_7978,N_6171);
or U9509 (N_9509,N_7602,N_7440);
nand U9510 (N_9510,N_6194,N_7361);
and U9511 (N_9511,N_7565,N_6320);
or U9512 (N_9512,N_6858,N_6203);
or U9513 (N_9513,N_6582,N_7879);
nor U9514 (N_9514,N_7304,N_7022);
nand U9515 (N_9515,N_6163,N_7587);
or U9516 (N_9516,N_6267,N_6921);
or U9517 (N_9517,N_7715,N_6807);
and U9518 (N_9518,N_6357,N_6112);
xor U9519 (N_9519,N_6355,N_7857);
or U9520 (N_9520,N_7441,N_6772);
nand U9521 (N_9521,N_7617,N_6131);
nor U9522 (N_9522,N_6111,N_6804);
xnor U9523 (N_9523,N_7549,N_7879);
and U9524 (N_9524,N_6854,N_6639);
or U9525 (N_9525,N_7825,N_7335);
xnor U9526 (N_9526,N_6485,N_6012);
nand U9527 (N_9527,N_7114,N_7451);
or U9528 (N_9528,N_7599,N_6810);
and U9529 (N_9529,N_7043,N_6099);
or U9530 (N_9530,N_7032,N_6079);
nor U9531 (N_9531,N_6562,N_7111);
or U9532 (N_9532,N_6700,N_6324);
nand U9533 (N_9533,N_7353,N_7120);
nand U9534 (N_9534,N_7143,N_7955);
and U9535 (N_9535,N_7248,N_6272);
nand U9536 (N_9536,N_7480,N_7475);
and U9537 (N_9537,N_7608,N_6921);
nor U9538 (N_9538,N_6380,N_7386);
nor U9539 (N_9539,N_7817,N_6872);
nor U9540 (N_9540,N_6344,N_6465);
and U9541 (N_9541,N_6012,N_6898);
nor U9542 (N_9542,N_7925,N_6138);
nand U9543 (N_9543,N_6697,N_7016);
nor U9544 (N_9544,N_6777,N_6170);
and U9545 (N_9545,N_6425,N_7267);
or U9546 (N_9546,N_6953,N_7299);
or U9547 (N_9547,N_7955,N_7791);
and U9548 (N_9548,N_6081,N_6942);
and U9549 (N_9549,N_7319,N_6737);
or U9550 (N_9550,N_6491,N_6725);
or U9551 (N_9551,N_7812,N_7760);
or U9552 (N_9552,N_6316,N_7415);
nor U9553 (N_9553,N_7574,N_6734);
and U9554 (N_9554,N_7422,N_6957);
and U9555 (N_9555,N_6490,N_7577);
or U9556 (N_9556,N_6284,N_6647);
nor U9557 (N_9557,N_7928,N_6130);
nor U9558 (N_9558,N_7836,N_6539);
or U9559 (N_9559,N_6409,N_6442);
nor U9560 (N_9560,N_7414,N_7278);
nor U9561 (N_9561,N_6641,N_6248);
or U9562 (N_9562,N_7845,N_7850);
nand U9563 (N_9563,N_6432,N_7562);
nor U9564 (N_9564,N_6366,N_7378);
and U9565 (N_9565,N_7036,N_6741);
nand U9566 (N_9566,N_6764,N_6810);
nor U9567 (N_9567,N_7135,N_6236);
nor U9568 (N_9568,N_7429,N_7632);
nor U9569 (N_9569,N_7918,N_7122);
and U9570 (N_9570,N_6377,N_6738);
nand U9571 (N_9571,N_7012,N_7619);
nor U9572 (N_9572,N_7600,N_7084);
nor U9573 (N_9573,N_6150,N_7382);
nor U9574 (N_9574,N_6907,N_7884);
and U9575 (N_9575,N_7269,N_6246);
nor U9576 (N_9576,N_7565,N_6492);
nand U9577 (N_9577,N_6469,N_7128);
nand U9578 (N_9578,N_6406,N_7465);
or U9579 (N_9579,N_7321,N_6087);
nand U9580 (N_9580,N_6323,N_6796);
and U9581 (N_9581,N_7759,N_7972);
and U9582 (N_9582,N_6991,N_7942);
nand U9583 (N_9583,N_6290,N_6937);
xnor U9584 (N_9584,N_7952,N_7625);
and U9585 (N_9585,N_6805,N_7307);
nand U9586 (N_9586,N_7361,N_6999);
nand U9587 (N_9587,N_6757,N_6806);
and U9588 (N_9588,N_7721,N_6959);
and U9589 (N_9589,N_7624,N_7661);
and U9590 (N_9590,N_7061,N_6238);
nand U9591 (N_9591,N_6893,N_7291);
nand U9592 (N_9592,N_6609,N_6340);
nand U9593 (N_9593,N_7267,N_7376);
and U9594 (N_9594,N_7518,N_7306);
nor U9595 (N_9595,N_6464,N_7534);
xor U9596 (N_9596,N_7778,N_6688);
or U9597 (N_9597,N_7423,N_7739);
nor U9598 (N_9598,N_6297,N_7547);
and U9599 (N_9599,N_6610,N_7446);
nand U9600 (N_9600,N_6649,N_6551);
nand U9601 (N_9601,N_7089,N_6370);
and U9602 (N_9602,N_7064,N_6804);
xnor U9603 (N_9603,N_7288,N_6096);
or U9604 (N_9604,N_6701,N_6819);
nor U9605 (N_9605,N_7269,N_6476);
or U9606 (N_9606,N_6323,N_6355);
and U9607 (N_9607,N_7357,N_7947);
and U9608 (N_9608,N_7366,N_7446);
nor U9609 (N_9609,N_7852,N_6305);
nor U9610 (N_9610,N_6588,N_7894);
nor U9611 (N_9611,N_7905,N_7533);
nor U9612 (N_9612,N_6060,N_7919);
xnor U9613 (N_9613,N_7994,N_6554);
and U9614 (N_9614,N_7430,N_6587);
xnor U9615 (N_9615,N_7323,N_7983);
and U9616 (N_9616,N_6641,N_6903);
nor U9617 (N_9617,N_6159,N_7397);
and U9618 (N_9618,N_7303,N_7023);
nor U9619 (N_9619,N_7826,N_7722);
and U9620 (N_9620,N_6490,N_7279);
nand U9621 (N_9621,N_7211,N_7195);
or U9622 (N_9622,N_6531,N_6351);
nor U9623 (N_9623,N_7152,N_6826);
or U9624 (N_9624,N_6258,N_7621);
nand U9625 (N_9625,N_7243,N_6845);
xnor U9626 (N_9626,N_6475,N_6688);
nor U9627 (N_9627,N_6895,N_6954);
nand U9628 (N_9628,N_6009,N_6861);
and U9629 (N_9629,N_7332,N_6047);
nor U9630 (N_9630,N_6219,N_6315);
nand U9631 (N_9631,N_7866,N_7152);
xor U9632 (N_9632,N_6905,N_7849);
nand U9633 (N_9633,N_7473,N_7055);
nor U9634 (N_9634,N_6067,N_7235);
or U9635 (N_9635,N_6041,N_7974);
and U9636 (N_9636,N_6269,N_6836);
or U9637 (N_9637,N_6212,N_7515);
nor U9638 (N_9638,N_7944,N_7679);
or U9639 (N_9639,N_6244,N_7305);
or U9640 (N_9640,N_6175,N_6286);
or U9641 (N_9641,N_6481,N_7977);
nand U9642 (N_9642,N_7696,N_7179);
nor U9643 (N_9643,N_6825,N_6247);
or U9644 (N_9644,N_7986,N_6668);
and U9645 (N_9645,N_6869,N_6007);
nor U9646 (N_9646,N_6567,N_6310);
or U9647 (N_9647,N_7238,N_7112);
nor U9648 (N_9648,N_7241,N_6756);
or U9649 (N_9649,N_6465,N_6778);
nand U9650 (N_9650,N_6375,N_7757);
or U9651 (N_9651,N_7341,N_6747);
or U9652 (N_9652,N_6642,N_6276);
or U9653 (N_9653,N_7493,N_7717);
and U9654 (N_9654,N_6443,N_6358);
nand U9655 (N_9655,N_6175,N_6458);
nor U9656 (N_9656,N_7288,N_7135);
nand U9657 (N_9657,N_7515,N_7712);
and U9658 (N_9658,N_7105,N_6285);
or U9659 (N_9659,N_6568,N_7515);
nor U9660 (N_9660,N_6971,N_6701);
nor U9661 (N_9661,N_6521,N_6579);
xnor U9662 (N_9662,N_6758,N_7399);
xnor U9663 (N_9663,N_7676,N_7790);
xnor U9664 (N_9664,N_7575,N_7555);
nor U9665 (N_9665,N_6345,N_6973);
xor U9666 (N_9666,N_6426,N_6119);
and U9667 (N_9667,N_6657,N_6945);
or U9668 (N_9668,N_7789,N_7523);
or U9669 (N_9669,N_6000,N_7690);
or U9670 (N_9670,N_6260,N_6775);
nand U9671 (N_9671,N_6449,N_7639);
and U9672 (N_9672,N_6107,N_7881);
nor U9673 (N_9673,N_7263,N_7760);
and U9674 (N_9674,N_6928,N_6431);
nand U9675 (N_9675,N_6498,N_6624);
nand U9676 (N_9676,N_6084,N_6626);
xor U9677 (N_9677,N_7258,N_6756);
xnor U9678 (N_9678,N_7218,N_7620);
and U9679 (N_9679,N_6583,N_7885);
or U9680 (N_9680,N_6472,N_7444);
nand U9681 (N_9681,N_7077,N_7835);
xnor U9682 (N_9682,N_7659,N_6601);
nor U9683 (N_9683,N_6096,N_7175);
or U9684 (N_9684,N_6863,N_6059);
nor U9685 (N_9685,N_7614,N_7520);
and U9686 (N_9686,N_6599,N_6410);
nor U9687 (N_9687,N_6216,N_6325);
or U9688 (N_9688,N_7795,N_6174);
nor U9689 (N_9689,N_7011,N_7481);
nor U9690 (N_9690,N_7876,N_7926);
nor U9691 (N_9691,N_7238,N_7650);
xor U9692 (N_9692,N_6583,N_7821);
and U9693 (N_9693,N_7028,N_6908);
and U9694 (N_9694,N_7493,N_7696);
nand U9695 (N_9695,N_7824,N_6077);
or U9696 (N_9696,N_7509,N_6073);
nor U9697 (N_9697,N_7678,N_7339);
xor U9698 (N_9698,N_7370,N_7888);
and U9699 (N_9699,N_6664,N_6767);
or U9700 (N_9700,N_6868,N_6303);
or U9701 (N_9701,N_7989,N_7861);
and U9702 (N_9702,N_7060,N_7369);
nor U9703 (N_9703,N_6408,N_7441);
nand U9704 (N_9704,N_6366,N_7161);
nand U9705 (N_9705,N_6840,N_7073);
xor U9706 (N_9706,N_6848,N_7170);
nor U9707 (N_9707,N_7310,N_7927);
or U9708 (N_9708,N_7038,N_7019);
xor U9709 (N_9709,N_7674,N_7104);
nand U9710 (N_9710,N_6285,N_6981);
or U9711 (N_9711,N_7238,N_7316);
or U9712 (N_9712,N_7605,N_6361);
nor U9713 (N_9713,N_6695,N_7128);
and U9714 (N_9714,N_6356,N_7277);
or U9715 (N_9715,N_6986,N_7429);
nand U9716 (N_9716,N_7943,N_6017);
nand U9717 (N_9717,N_7119,N_7567);
xor U9718 (N_9718,N_6396,N_6552);
nor U9719 (N_9719,N_6261,N_7205);
xor U9720 (N_9720,N_6738,N_7984);
or U9721 (N_9721,N_7704,N_7823);
nand U9722 (N_9722,N_6197,N_7519);
nand U9723 (N_9723,N_7701,N_7476);
nor U9724 (N_9724,N_7105,N_7803);
xnor U9725 (N_9725,N_7422,N_7590);
nand U9726 (N_9726,N_6081,N_7753);
or U9727 (N_9727,N_6198,N_7653);
nor U9728 (N_9728,N_7751,N_6460);
and U9729 (N_9729,N_6797,N_6541);
nand U9730 (N_9730,N_7843,N_7423);
nand U9731 (N_9731,N_7593,N_6461);
and U9732 (N_9732,N_7723,N_6313);
and U9733 (N_9733,N_7644,N_6303);
nor U9734 (N_9734,N_7092,N_6288);
or U9735 (N_9735,N_6707,N_6536);
nand U9736 (N_9736,N_7070,N_6512);
nor U9737 (N_9737,N_6974,N_6301);
xnor U9738 (N_9738,N_7836,N_6763);
or U9739 (N_9739,N_6032,N_7953);
xnor U9740 (N_9740,N_6733,N_6349);
and U9741 (N_9741,N_7581,N_6203);
xor U9742 (N_9742,N_6982,N_7953);
or U9743 (N_9743,N_6251,N_6019);
nor U9744 (N_9744,N_6085,N_7212);
nand U9745 (N_9745,N_7565,N_6780);
nand U9746 (N_9746,N_6022,N_6163);
and U9747 (N_9747,N_6201,N_7447);
nand U9748 (N_9748,N_6186,N_7144);
and U9749 (N_9749,N_6893,N_7843);
and U9750 (N_9750,N_6456,N_7977);
and U9751 (N_9751,N_6870,N_7001);
xor U9752 (N_9752,N_7795,N_6099);
or U9753 (N_9753,N_6695,N_7444);
nor U9754 (N_9754,N_6073,N_6915);
and U9755 (N_9755,N_6889,N_7448);
or U9756 (N_9756,N_6715,N_6884);
nor U9757 (N_9757,N_6542,N_6590);
nor U9758 (N_9758,N_6049,N_7949);
or U9759 (N_9759,N_6866,N_7343);
and U9760 (N_9760,N_6144,N_6570);
nand U9761 (N_9761,N_7326,N_7494);
nor U9762 (N_9762,N_7233,N_7163);
nor U9763 (N_9763,N_7754,N_6698);
nor U9764 (N_9764,N_6814,N_7418);
and U9765 (N_9765,N_7216,N_7021);
and U9766 (N_9766,N_6385,N_6812);
or U9767 (N_9767,N_7319,N_7262);
nor U9768 (N_9768,N_6409,N_7778);
nand U9769 (N_9769,N_7813,N_6694);
nor U9770 (N_9770,N_7276,N_7047);
and U9771 (N_9771,N_7743,N_7070);
nand U9772 (N_9772,N_7833,N_7934);
or U9773 (N_9773,N_7126,N_7067);
nand U9774 (N_9774,N_7038,N_6228);
nor U9775 (N_9775,N_7839,N_6595);
nor U9776 (N_9776,N_7018,N_7424);
nor U9777 (N_9777,N_6149,N_7985);
nor U9778 (N_9778,N_7964,N_7043);
or U9779 (N_9779,N_6448,N_6450);
nand U9780 (N_9780,N_6893,N_6283);
nor U9781 (N_9781,N_6815,N_7005);
nand U9782 (N_9782,N_7694,N_6905);
xor U9783 (N_9783,N_7960,N_6909);
or U9784 (N_9784,N_7267,N_7606);
nor U9785 (N_9785,N_7354,N_6306);
and U9786 (N_9786,N_7883,N_6261);
or U9787 (N_9787,N_6411,N_7231);
nor U9788 (N_9788,N_7564,N_7373);
xnor U9789 (N_9789,N_7594,N_6585);
nor U9790 (N_9790,N_6048,N_6414);
nand U9791 (N_9791,N_7601,N_6702);
or U9792 (N_9792,N_6849,N_6193);
nand U9793 (N_9793,N_6094,N_6734);
nor U9794 (N_9794,N_7281,N_6658);
and U9795 (N_9795,N_6164,N_6104);
xor U9796 (N_9796,N_7090,N_6170);
nand U9797 (N_9797,N_6546,N_6595);
xnor U9798 (N_9798,N_6102,N_7198);
and U9799 (N_9799,N_6398,N_6970);
or U9800 (N_9800,N_7376,N_6990);
nand U9801 (N_9801,N_6423,N_6497);
and U9802 (N_9802,N_6433,N_6519);
xnor U9803 (N_9803,N_6011,N_6429);
nand U9804 (N_9804,N_7379,N_6669);
xor U9805 (N_9805,N_7429,N_6567);
or U9806 (N_9806,N_6308,N_7703);
nor U9807 (N_9807,N_7848,N_6386);
or U9808 (N_9808,N_6883,N_6089);
nand U9809 (N_9809,N_6696,N_7641);
xnor U9810 (N_9810,N_7891,N_7818);
nand U9811 (N_9811,N_7057,N_6812);
and U9812 (N_9812,N_7994,N_7627);
xnor U9813 (N_9813,N_6148,N_7811);
or U9814 (N_9814,N_6180,N_6957);
or U9815 (N_9815,N_6710,N_6957);
or U9816 (N_9816,N_6033,N_6551);
nor U9817 (N_9817,N_7611,N_6256);
or U9818 (N_9818,N_6248,N_6512);
nand U9819 (N_9819,N_7354,N_7937);
and U9820 (N_9820,N_7445,N_7793);
xnor U9821 (N_9821,N_6761,N_6609);
and U9822 (N_9822,N_7303,N_6700);
xor U9823 (N_9823,N_6689,N_6049);
and U9824 (N_9824,N_6082,N_6004);
nand U9825 (N_9825,N_6006,N_7621);
nor U9826 (N_9826,N_7918,N_7524);
or U9827 (N_9827,N_7181,N_7067);
and U9828 (N_9828,N_7556,N_7438);
nor U9829 (N_9829,N_7148,N_6109);
or U9830 (N_9830,N_7268,N_6156);
nand U9831 (N_9831,N_7454,N_7117);
and U9832 (N_9832,N_6538,N_6928);
or U9833 (N_9833,N_6886,N_7928);
and U9834 (N_9834,N_7442,N_6894);
and U9835 (N_9835,N_7917,N_6279);
nand U9836 (N_9836,N_6663,N_7010);
and U9837 (N_9837,N_6430,N_7885);
and U9838 (N_9838,N_7017,N_7903);
nor U9839 (N_9839,N_7208,N_7976);
and U9840 (N_9840,N_7024,N_6491);
nor U9841 (N_9841,N_6940,N_7980);
nor U9842 (N_9842,N_6791,N_7273);
or U9843 (N_9843,N_6435,N_6117);
and U9844 (N_9844,N_6189,N_6936);
nand U9845 (N_9845,N_6534,N_6294);
nor U9846 (N_9846,N_6128,N_7780);
nand U9847 (N_9847,N_7725,N_6460);
or U9848 (N_9848,N_7464,N_7072);
nand U9849 (N_9849,N_7213,N_6116);
and U9850 (N_9850,N_6721,N_6653);
or U9851 (N_9851,N_6774,N_7767);
or U9852 (N_9852,N_6109,N_7732);
nand U9853 (N_9853,N_6305,N_7460);
nand U9854 (N_9854,N_7015,N_7193);
nor U9855 (N_9855,N_7687,N_6889);
and U9856 (N_9856,N_6959,N_6060);
nor U9857 (N_9857,N_7901,N_7838);
nor U9858 (N_9858,N_7081,N_6659);
xor U9859 (N_9859,N_7945,N_7834);
or U9860 (N_9860,N_7206,N_6212);
and U9861 (N_9861,N_7327,N_7061);
nor U9862 (N_9862,N_6275,N_7046);
and U9863 (N_9863,N_6382,N_7315);
or U9864 (N_9864,N_6652,N_7907);
nor U9865 (N_9865,N_7417,N_7707);
nor U9866 (N_9866,N_7684,N_7308);
nor U9867 (N_9867,N_7333,N_7419);
or U9868 (N_9868,N_7412,N_7645);
xnor U9869 (N_9869,N_6633,N_6521);
nand U9870 (N_9870,N_6199,N_7019);
or U9871 (N_9871,N_6537,N_6221);
or U9872 (N_9872,N_6759,N_6923);
nand U9873 (N_9873,N_6746,N_6273);
or U9874 (N_9874,N_6730,N_6808);
xnor U9875 (N_9875,N_6991,N_6106);
nor U9876 (N_9876,N_6131,N_6892);
nand U9877 (N_9877,N_6428,N_7542);
nor U9878 (N_9878,N_7238,N_6691);
and U9879 (N_9879,N_7805,N_7314);
nand U9880 (N_9880,N_6132,N_7019);
or U9881 (N_9881,N_6467,N_7135);
nand U9882 (N_9882,N_7009,N_7875);
nor U9883 (N_9883,N_7193,N_7174);
nor U9884 (N_9884,N_6451,N_6154);
xnor U9885 (N_9885,N_6323,N_6819);
or U9886 (N_9886,N_6644,N_6079);
xor U9887 (N_9887,N_6951,N_6922);
nand U9888 (N_9888,N_7827,N_6344);
xor U9889 (N_9889,N_7224,N_7050);
and U9890 (N_9890,N_6956,N_7611);
nand U9891 (N_9891,N_7327,N_7573);
or U9892 (N_9892,N_7918,N_6528);
nand U9893 (N_9893,N_7196,N_6304);
or U9894 (N_9894,N_6726,N_7017);
and U9895 (N_9895,N_6312,N_7457);
nor U9896 (N_9896,N_6510,N_7616);
and U9897 (N_9897,N_7401,N_6182);
nor U9898 (N_9898,N_6231,N_7088);
or U9899 (N_9899,N_6449,N_7695);
nand U9900 (N_9900,N_7807,N_7566);
and U9901 (N_9901,N_6727,N_6640);
and U9902 (N_9902,N_6731,N_7371);
nor U9903 (N_9903,N_7194,N_7832);
nor U9904 (N_9904,N_6213,N_6323);
nand U9905 (N_9905,N_7655,N_7976);
or U9906 (N_9906,N_7384,N_6326);
nor U9907 (N_9907,N_7874,N_6148);
or U9908 (N_9908,N_7422,N_6202);
and U9909 (N_9909,N_7428,N_7813);
nand U9910 (N_9910,N_7740,N_6938);
and U9911 (N_9911,N_6474,N_6221);
xor U9912 (N_9912,N_7778,N_7818);
or U9913 (N_9913,N_7192,N_7470);
nor U9914 (N_9914,N_7313,N_7781);
xor U9915 (N_9915,N_7348,N_7116);
and U9916 (N_9916,N_7809,N_7574);
or U9917 (N_9917,N_6877,N_6112);
xnor U9918 (N_9918,N_6536,N_7934);
nor U9919 (N_9919,N_6135,N_6232);
nor U9920 (N_9920,N_7697,N_6139);
nand U9921 (N_9921,N_7267,N_6457);
or U9922 (N_9922,N_6120,N_6486);
xnor U9923 (N_9923,N_7364,N_6292);
xnor U9924 (N_9924,N_6725,N_7233);
and U9925 (N_9925,N_6150,N_7536);
nand U9926 (N_9926,N_7313,N_6575);
nor U9927 (N_9927,N_7507,N_6359);
nand U9928 (N_9928,N_7882,N_6554);
nand U9929 (N_9929,N_6980,N_7789);
and U9930 (N_9930,N_6095,N_7631);
nor U9931 (N_9931,N_6894,N_7514);
and U9932 (N_9932,N_7589,N_6255);
nor U9933 (N_9933,N_6383,N_7060);
nand U9934 (N_9934,N_6769,N_7219);
and U9935 (N_9935,N_6848,N_6138);
xnor U9936 (N_9936,N_7501,N_6214);
nand U9937 (N_9937,N_7257,N_6632);
xnor U9938 (N_9938,N_6374,N_6460);
or U9939 (N_9939,N_6569,N_7342);
or U9940 (N_9940,N_7410,N_6234);
nor U9941 (N_9941,N_6742,N_6391);
or U9942 (N_9942,N_7922,N_7047);
nand U9943 (N_9943,N_6716,N_7484);
or U9944 (N_9944,N_7921,N_6790);
and U9945 (N_9945,N_7707,N_7388);
nor U9946 (N_9946,N_6768,N_7114);
and U9947 (N_9947,N_7869,N_7800);
nand U9948 (N_9948,N_6498,N_6679);
nor U9949 (N_9949,N_6768,N_7428);
and U9950 (N_9950,N_6865,N_7555);
or U9951 (N_9951,N_7361,N_6852);
and U9952 (N_9952,N_6842,N_7166);
and U9953 (N_9953,N_6733,N_6970);
nand U9954 (N_9954,N_7353,N_6879);
nand U9955 (N_9955,N_6445,N_6410);
nand U9956 (N_9956,N_6799,N_7004);
and U9957 (N_9957,N_7774,N_7490);
and U9958 (N_9958,N_7283,N_6884);
and U9959 (N_9959,N_6081,N_7100);
nand U9960 (N_9960,N_6653,N_6999);
and U9961 (N_9961,N_6168,N_6396);
or U9962 (N_9962,N_7981,N_7177);
and U9963 (N_9963,N_7509,N_7280);
nand U9964 (N_9964,N_6411,N_6315);
nor U9965 (N_9965,N_6456,N_6860);
xor U9966 (N_9966,N_7766,N_7384);
and U9967 (N_9967,N_6659,N_6737);
or U9968 (N_9968,N_7303,N_6513);
nand U9969 (N_9969,N_7574,N_6603);
nand U9970 (N_9970,N_6721,N_6341);
xor U9971 (N_9971,N_7143,N_6048);
or U9972 (N_9972,N_6932,N_6934);
xnor U9973 (N_9973,N_7500,N_7719);
nor U9974 (N_9974,N_6628,N_6456);
nand U9975 (N_9975,N_6584,N_7574);
nor U9976 (N_9976,N_7707,N_6353);
and U9977 (N_9977,N_6028,N_7771);
or U9978 (N_9978,N_7861,N_6871);
and U9979 (N_9979,N_7180,N_7646);
nor U9980 (N_9980,N_6807,N_6215);
or U9981 (N_9981,N_6844,N_7354);
xnor U9982 (N_9982,N_7925,N_6842);
nor U9983 (N_9983,N_7915,N_6031);
nand U9984 (N_9984,N_6262,N_6550);
nor U9985 (N_9985,N_7856,N_7395);
nor U9986 (N_9986,N_6993,N_7910);
xnor U9987 (N_9987,N_6254,N_7630);
or U9988 (N_9988,N_7323,N_7828);
nand U9989 (N_9989,N_7155,N_6703);
nand U9990 (N_9990,N_6704,N_7262);
and U9991 (N_9991,N_6475,N_7329);
or U9992 (N_9992,N_7792,N_7046);
and U9993 (N_9993,N_6403,N_6736);
nor U9994 (N_9994,N_7464,N_7102);
nand U9995 (N_9995,N_7354,N_7434);
and U9996 (N_9996,N_7694,N_7644);
nor U9997 (N_9997,N_7121,N_7878);
or U9998 (N_9998,N_7745,N_7219);
or U9999 (N_9999,N_6889,N_7338);
nand U10000 (N_10000,N_8490,N_8169);
nand U10001 (N_10001,N_9905,N_9924);
nand U10002 (N_10002,N_8144,N_9000);
and U10003 (N_10003,N_8964,N_9080);
and U10004 (N_10004,N_8422,N_8041);
and U10005 (N_10005,N_9726,N_9003);
nor U10006 (N_10006,N_9558,N_9465);
nor U10007 (N_10007,N_8638,N_8627);
nand U10008 (N_10008,N_8056,N_9881);
and U10009 (N_10009,N_8544,N_8680);
and U10010 (N_10010,N_9838,N_8877);
and U10011 (N_10011,N_8613,N_9024);
or U10012 (N_10012,N_9565,N_9746);
nand U10013 (N_10013,N_8579,N_9248);
nor U10014 (N_10014,N_8929,N_9595);
nand U10015 (N_10015,N_8678,N_9666);
nor U10016 (N_10016,N_9758,N_9743);
or U10017 (N_10017,N_8377,N_8453);
or U10018 (N_10018,N_9522,N_9963);
nor U10019 (N_10019,N_8717,N_9115);
nand U10020 (N_10020,N_9395,N_9362);
or U10021 (N_10021,N_8020,N_8458);
and U10022 (N_10022,N_8094,N_8405);
or U10023 (N_10023,N_9480,N_8112);
nand U10024 (N_10024,N_9437,N_8322);
and U10025 (N_10025,N_8679,N_9373);
xnor U10026 (N_10026,N_8858,N_9897);
or U10027 (N_10027,N_8383,N_9875);
nand U10028 (N_10028,N_8419,N_8621);
nand U10029 (N_10029,N_8974,N_8539);
and U10030 (N_10030,N_8291,N_8015);
nor U10031 (N_10031,N_9671,N_9640);
or U10032 (N_10032,N_8750,N_8861);
nand U10033 (N_10033,N_8372,N_9898);
nand U10034 (N_10034,N_8868,N_8022);
nor U10035 (N_10035,N_9561,N_9956);
and U10036 (N_10036,N_9001,N_8543);
or U10037 (N_10037,N_9074,N_8198);
nand U10038 (N_10038,N_8299,N_8168);
nor U10039 (N_10039,N_8801,N_8618);
nor U10040 (N_10040,N_9809,N_9108);
and U10041 (N_10041,N_8784,N_9686);
xnor U10042 (N_10042,N_9654,N_8869);
or U10043 (N_10043,N_9864,N_9773);
xnor U10044 (N_10044,N_9976,N_9767);
nor U10045 (N_10045,N_9874,N_9774);
or U10046 (N_10046,N_8503,N_8746);
nand U10047 (N_10047,N_8770,N_9338);
nor U10048 (N_10048,N_9668,N_8567);
xor U10049 (N_10049,N_8317,N_8741);
xnor U10050 (N_10050,N_8161,N_9962);
nand U10051 (N_10051,N_9837,N_9946);
xnor U10052 (N_10052,N_8674,N_8077);
and U10053 (N_10053,N_9701,N_9820);
or U10054 (N_10054,N_9321,N_9681);
xnor U10055 (N_10055,N_9759,N_9981);
or U10056 (N_10056,N_9243,N_9698);
nand U10057 (N_10057,N_9256,N_8608);
xor U10058 (N_10058,N_9691,N_8673);
and U10059 (N_10059,N_8334,N_8559);
and U10060 (N_10060,N_9084,N_8612);
xor U10061 (N_10061,N_8259,N_9221);
or U10062 (N_10062,N_8061,N_9078);
nand U10063 (N_10063,N_8229,N_9851);
and U10064 (N_10064,N_8464,N_9937);
xor U10065 (N_10065,N_8328,N_8906);
nor U10066 (N_10066,N_8595,N_8462);
and U10067 (N_10067,N_8472,N_9993);
and U10068 (N_10068,N_8250,N_8243);
nand U10069 (N_10069,N_9061,N_9066);
xnor U10070 (N_10070,N_8517,N_8375);
and U10071 (N_10071,N_9152,N_9232);
or U10072 (N_10072,N_9415,N_8727);
nand U10073 (N_10073,N_8799,N_8658);
nor U10074 (N_10074,N_9380,N_8188);
or U10075 (N_10075,N_8954,N_8211);
and U10076 (N_10076,N_9229,N_8406);
xor U10077 (N_10077,N_9068,N_8930);
nand U10078 (N_10078,N_8786,N_9617);
nand U10079 (N_10079,N_8730,N_8696);
xor U10080 (N_10080,N_8631,N_9740);
nand U10081 (N_10081,N_9130,N_9775);
nand U10082 (N_10082,N_9877,N_8392);
nor U10083 (N_10083,N_9205,N_8755);
and U10084 (N_10084,N_9871,N_8356);
nand U10085 (N_10085,N_8442,N_9970);
and U10086 (N_10086,N_9376,N_9289);
nor U10087 (N_10087,N_9272,N_9992);
nor U10088 (N_10088,N_8586,N_9330);
and U10089 (N_10089,N_9960,N_8451);
xor U10090 (N_10090,N_9233,N_9995);
nor U10091 (N_10091,N_9337,N_9984);
or U10092 (N_10092,N_9927,N_9231);
or U10093 (N_10093,N_9916,N_9163);
nand U10094 (N_10094,N_9323,N_8220);
nand U10095 (N_10095,N_9463,N_9719);
and U10096 (N_10096,N_9386,N_9624);
nor U10097 (N_10097,N_9786,N_9936);
nand U10098 (N_10098,N_9636,N_8561);
or U10099 (N_10099,N_9751,N_9725);
or U10100 (N_10100,N_9270,N_9365);
or U10101 (N_10101,N_8216,N_8558);
and U10102 (N_10102,N_8598,N_8305);
nand U10103 (N_10103,N_8652,N_8626);
xor U10104 (N_10104,N_9684,N_9915);
xor U10105 (N_10105,N_8668,N_8528);
or U10106 (N_10106,N_8689,N_9138);
and U10107 (N_10107,N_9201,N_9326);
nand U10108 (N_10108,N_8206,N_8684);
or U10109 (N_10109,N_9812,N_8183);
and U10110 (N_10110,N_8540,N_8635);
nor U10111 (N_10111,N_8564,N_8908);
or U10112 (N_10112,N_9127,N_9085);
nor U10113 (N_10113,N_9805,N_8478);
and U10114 (N_10114,N_8466,N_8705);
xnor U10115 (N_10115,N_8956,N_9917);
and U10116 (N_10116,N_8002,N_8817);
and U10117 (N_10117,N_8411,N_9510);
nor U10118 (N_10118,N_9649,N_9979);
or U10119 (N_10119,N_9333,N_8060);
or U10120 (N_10120,N_9925,N_9642);
and U10121 (N_10121,N_9996,N_8095);
nor U10122 (N_10122,N_8959,N_8457);
nand U10123 (N_10123,N_8532,N_9884);
or U10124 (N_10124,N_8104,N_9448);
nand U10125 (N_10125,N_9919,N_8504);
or U10126 (N_10126,N_9643,N_8656);
or U10127 (N_10127,N_8233,N_9606);
or U10128 (N_10128,N_9511,N_9034);
nand U10129 (N_10129,N_9801,N_9446);
xor U10130 (N_10130,N_8498,N_9219);
nor U10131 (N_10131,N_8990,N_8475);
or U10132 (N_10132,N_9204,N_9890);
nor U10133 (N_10133,N_9264,N_8890);
or U10134 (N_10134,N_8019,N_9142);
nand U10135 (N_10135,N_9417,N_9348);
nor U10136 (N_10136,N_9542,N_9458);
nand U10137 (N_10137,N_9261,N_9795);
nor U10138 (N_10138,N_9986,N_8366);
and U10139 (N_10139,N_8807,N_8046);
or U10140 (N_10140,N_8506,N_9782);
nor U10141 (N_10141,N_8382,N_9860);
or U10142 (N_10142,N_9361,N_8024);
and U10143 (N_10143,N_8816,N_9468);
xnor U10144 (N_10144,N_8167,N_8724);
nand U10145 (N_10145,N_9699,N_9126);
or U10146 (N_10146,N_9293,N_8887);
and U10147 (N_10147,N_9814,N_9790);
nand U10148 (N_10148,N_8455,N_9299);
nor U10149 (N_10149,N_8833,N_9083);
nand U10150 (N_10150,N_8281,N_8634);
or U10151 (N_10151,N_9182,N_8938);
nor U10152 (N_10152,N_9259,N_8685);
xnor U10153 (N_10153,N_9639,N_8379);
or U10154 (N_10154,N_9501,N_9183);
or U10155 (N_10155,N_8950,N_8324);
and U10156 (N_10156,N_8027,N_9045);
or U10157 (N_10157,N_8201,N_9492);
nand U10158 (N_10158,N_8249,N_9283);
and U10159 (N_10159,N_9096,N_9263);
nor U10160 (N_10160,N_9721,N_8905);
nor U10161 (N_10161,N_9482,N_9736);
nor U10162 (N_10162,N_9474,N_8417);
nor U10163 (N_10163,N_9778,N_8628);
nor U10164 (N_10164,N_8496,N_9077);
or U10165 (N_10165,N_8510,N_8278);
and U10166 (N_10166,N_9102,N_9267);
nand U10167 (N_10167,N_9434,N_9529);
or U10168 (N_10168,N_8686,N_8934);
nor U10169 (N_10169,N_8436,N_9495);
or U10170 (N_10170,N_8309,N_9978);
or U10171 (N_10171,N_9225,N_9822);
nor U10172 (N_10172,N_8428,N_8253);
and U10173 (N_10173,N_8106,N_8482);
nor U10174 (N_10174,N_8163,N_9626);
or U10175 (N_10175,N_9194,N_8092);
nand U10176 (N_10176,N_8234,N_9009);
and U10177 (N_10177,N_9368,N_9803);
nor U10178 (N_10178,N_8697,N_9300);
nand U10179 (N_10179,N_8109,N_9167);
nand U10180 (N_10180,N_8074,N_9297);
nor U10181 (N_10181,N_8891,N_8107);
nand U10182 (N_10182,N_8174,N_8726);
nand U10183 (N_10183,N_9041,N_8194);
or U10184 (N_10184,N_8541,N_8214);
nand U10185 (N_10185,N_9857,N_9889);
nor U10186 (N_10186,N_9982,N_9964);
nor U10187 (N_10187,N_8017,N_9252);
and U10188 (N_10188,N_9548,N_9967);
and U10189 (N_10189,N_9718,N_9763);
nor U10190 (N_10190,N_8399,N_8552);
or U10191 (N_10191,N_9693,N_8512);
or U10192 (N_10192,N_9042,N_8571);
nor U10193 (N_10193,N_8568,N_9650);
xnor U10194 (N_10194,N_9489,N_9904);
nand U10195 (N_10195,N_8763,N_8360);
or U10196 (N_10196,N_8189,N_8976);
nor U10197 (N_10197,N_9900,N_9538);
or U10198 (N_10198,N_8283,N_8912);
or U10199 (N_10199,N_9702,N_9032);
and U10200 (N_10200,N_8308,N_8225);
or U10201 (N_10201,N_8994,N_8669);
or U10202 (N_10202,N_8640,N_9371);
nand U10203 (N_10203,N_8067,N_9662);
nor U10204 (N_10204,N_9239,N_9447);
or U10205 (N_10205,N_8866,N_8344);
nand U10206 (N_10206,N_8639,N_8236);
or U10207 (N_10207,N_9100,N_9597);
or U10208 (N_10208,N_9408,N_9170);
nor U10209 (N_10209,N_8527,N_9113);
or U10210 (N_10210,N_8348,N_9709);
xnor U10211 (N_10211,N_9679,N_9950);
or U10212 (N_10212,N_8748,N_9584);
nand U10213 (N_10213,N_8919,N_9282);
or U10214 (N_10214,N_9532,N_9262);
xnor U10215 (N_10215,N_8747,N_8038);
and U10216 (N_10216,N_8581,N_9724);
and U10217 (N_10217,N_9816,N_8099);
nand U10218 (N_10218,N_9470,N_9572);
nor U10219 (N_10219,N_9485,N_9393);
xor U10220 (N_10220,N_9375,N_8148);
and U10221 (N_10221,N_9294,N_9153);
nor U10222 (N_10222,N_8176,N_9880);
xor U10223 (N_10223,N_8865,N_8511);
xor U10224 (N_10224,N_9585,N_8327);
nand U10225 (N_10225,N_9846,N_9535);
nor U10226 (N_10226,N_8205,N_8819);
and U10227 (N_10227,N_8365,N_9622);
or U10228 (N_10228,N_9352,N_9530);
nor U10229 (N_10229,N_9848,N_9057);
or U10230 (N_10230,N_9332,N_9940);
and U10231 (N_10231,N_8670,N_9493);
and U10232 (N_10232,N_8145,N_9519);
nor U10233 (N_10233,N_8153,N_9443);
or U10234 (N_10234,N_9481,N_8903);
nand U10235 (N_10235,N_8520,N_9451);
nand U10236 (N_10236,N_9308,N_8516);
and U10237 (N_10237,N_9257,N_9603);
and U10238 (N_10238,N_9018,N_8803);
nand U10239 (N_10239,N_9344,N_8850);
nor U10240 (N_10240,N_9133,N_8494);
nor U10241 (N_10241,N_8739,N_9055);
nand U10242 (N_10242,N_8909,N_8393);
and U10243 (N_10243,N_8232,N_9364);
nand U10244 (N_10244,N_9628,N_8863);
nand U10245 (N_10245,N_8218,N_8445);
and U10246 (N_10246,N_9806,N_8603);
nor U10247 (N_10247,N_9214,N_8132);
xor U10248 (N_10248,N_9621,N_9985);
or U10249 (N_10249,N_8646,N_8049);
nor U10250 (N_10250,N_9341,N_8054);
nor U10251 (N_10251,N_8949,N_8040);
or U10252 (N_10252,N_9191,N_9840);
xnor U10253 (N_10253,N_8815,N_9052);
nor U10254 (N_10254,N_8184,N_9112);
nand U10255 (N_10255,N_9385,N_8790);
nor U10256 (N_10256,N_8493,N_8433);
nor U10257 (N_10257,N_8400,N_8387);
nand U10258 (N_10258,N_9712,N_8212);
and U10259 (N_10259,N_9487,N_9253);
and U10260 (N_10260,N_9328,N_8265);
nand U10261 (N_10261,N_9390,N_8333);
nand U10262 (N_10262,N_9195,N_8335);
nor U10263 (N_10263,N_9598,N_8548);
and U10264 (N_10264,N_9619,N_8108);
or U10265 (N_10265,N_9974,N_8072);
or U10266 (N_10266,N_9335,N_9659);
or U10267 (N_10267,N_8809,N_8783);
or U10268 (N_10268,N_8264,N_9502);
nor U10269 (N_10269,N_9957,N_9757);
nor U10270 (N_10270,N_9277,N_9312);
xor U10271 (N_10271,N_9780,N_9159);
or U10272 (N_10272,N_8113,N_8862);
xor U10273 (N_10273,N_9409,N_9952);
or U10274 (N_10274,N_8881,N_8776);
nand U10275 (N_10275,N_9863,N_9768);
nand U10276 (N_10276,N_9644,N_8005);
xnor U10277 (N_10277,N_8509,N_9752);
nor U10278 (N_10278,N_8984,N_9469);
nand U10279 (N_10279,N_8155,N_8350);
nand U10280 (N_10280,N_9665,N_9435);
nor U10281 (N_10281,N_8675,N_9477);
and U10282 (N_10282,N_8172,N_8070);
or U10283 (N_10283,N_9620,N_9947);
and U10284 (N_10284,N_9206,N_9452);
nor U10285 (N_10285,N_9506,N_9955);
nor U10286 (N_10286,N_9802,N_9030);
and U10287 (N_10287,N_9852,N_8032);
nor U10288 (N_10288,N_8916,N_8298);
nor U10289 (N_10289,N_9181,N_9973);
or U10290 (N_10290,N_8483,N_8319);
nor U10291 (N_10291,N_8204,N_9868);
nand U10292 (N_10292,N_9141,N_9761);
or U10293 (N_10293,N_9013,N_9035);
or U10294 (N_10294,N_9902,N_8362);
or U10295 (N_10295,N_9888,N_8449);
or U10296 (N_10296,N_8742,N_9178);
and U10297 (N_10297,N_8058,N_8339);
nor U10298 (N_10298,N_8485,N_8810);
nand U10299 (N_10299,N_9922,N_9179);
or U10300 (N_10300,N_8068,N_8177);
and U10301 (N_10301,N_8376,N_9534);
nand U10302 (N_10302,N_8688,N_9526);
nor U10303 (N_10303,N_8459,N_9841);
nor U10304 (N_10304,N_9872,N_8128);
or U10305 (N_10305,N_8147,N_8057);
nor U10306 (N_10306,N_9989,N_8292);
nand U10307 (N_10307,N_9280,N_8170);
or U10308 (N_10308,N_9524,N_8468);
and U10309 (N_10309,N_9242,N_8467);
or U10310 (N_10310,N_9311,N_8590);
and U10311 (N_10311,N_9680,N_9564);
or U10312 (N_10312,N_8047,N_9954);
nor U10313 (N_10313,N_8471,N_9713);
nand U10314 (N_10314,N_8152,N_8190);
or U10315 (N_10315,N_9056,N_9063);
nor U10316 (N_10316,N_9611,N_9714);
xor U10317 (N_10317,N_9010,N_8515);
and U10318 (N_10318,N_8408,N_9069);
and U10319 (N_10319,N_8732,N_9516);
xor U10320 (N_10320,N_8843,N_9739);
and U10321 (N_10321,N_9423,N_9478);
and U10322 (N_10322,N_9125,N_9291);
or U10323 (N_10323,N_8323,N_8706);
nor U10324 (N_10324,N_9318,N_8708);
or U10325 (N_10325,N_9403,N_9807);
or U10326 (N_10326,N_8270,N_9400);
nand U10327 (N_10327,N_8637,N_8371);
or U10328 (N_10328,N_8910,N_9844);
nor U10329 (N_10329,N_8846,N_8423);
and U10330 (N_10330,N_8332,N_9111);
nor U10331 (N_10331,N_8915,N_9298);
nor U10332 (N_10332,N_9173,N_9991);
nor U10333 (N_10333,N_8712,N_9486);
nor U10334 (N_10334,N_9427,N_8285);
and U10335 (N_10335,N_9655,N_8655);
or U10336 (N_10336,N_9059,N_9137);
and U10337 (N_10337,N_9210,N_8945);
nor U10338 (N_10338,N_9071,N_8569);
and U10339 (N_10339,N_9410,N_8844);
and U10340 (N_10340,N_8968,N_9792);
nor U10341 (N_10341,N_8042,N_9994);
or U10342 (N_10342,N_8349,N_8962);
nor U10343 (N_10343,N_9934,N_8600);
or U10344 (N_10344,N_8606,N_8191);
nand U10345 (N_10345,N_9303,N_8280);
or U10346 (N_10346,N_9116,N_8576);
nor U10347 (N_10347,N_8363,N_8386);
nand U10348 (N_10348,N_8963,N_9131);
nand U10349 (N_10349,N_9945,N_9520);
nor U10350 (N_10350,N_8272,N_9284);
and U10351 (N_10351,N_9836,N_9488);
and U10352 (N_10352,N_9893,N_8760);
nand U10353 (N_10353,N_8083,N_9479);
nor U10354 (N_10354,N_9556,N_9260);
nor U10355 (N_10355,N_9087,N_9869);
nand U10356 (N_10356,N_8140,N_8087);
nand U10357 (N_10357,N_8514,N_8447);
or U10358 (N_10358,N_8583,N_8045);
nand U10359 (N_10359,N_8131,N_8050);
and U10360 (N_10360,N_9454,N_9398);
or U10361 (N_10361,N_8622,N_8538);
and U10362 (N_10362,N_8774,N_8311);
nor U10363 (N_10363,N_8125,N_9760);
and U10364 (N_10364,N_9406,N_9028);
and U10365 (N_10365,N_8031,N_8713);
nor U10366 (N_10366,N_8927,N_8756);
and U10367 (N_10367,N_9855,N_9278);
or U10368 (N_10368,N_8443,N_8217);
and U10369 (N_10369,N_8499,N_9005);
nor U10370 (N_10370,N_9528,N_8325);
or U10371 (N_10371,N_8922,N_9177);
nor U10372 (N_10372,N_8313,N_9865);
and U10373 (N_10373,N_8267,N_9696);
or U10374 (N_10374,N_8480,N_9586);
and U10375 (N_10375,N_8529,N_8864);
xnor U10376 (N_10376,N_9106,N_8254);
or U10377 (N_10377,N_9094,N_9514);
nand U10378 (N_10378,N_9667,N_8980);
nand U10379 (N_10379,N_8704,N_9459);
xor U10380 (N_10380,N_8505,N_8192);
nor U10381 (N_10381,N_9896,N_9811);
nor U10382 (N_10382,N_9324,N_8765);
and U10383 (N_10383,N_8178,N_9237);
nand U10384 (N_10384,N_9779,N_9271);
or U10385 (N_10385,N_9081,N_8316);
nor U10386 (N_10386,N_9673,N_9582);
and U10387 (N_10387,N_8545,N_8772);
or U10388 (N_10388,N_8018,N_8946);
and U10389 (N_10389,N_9789,N_9669);
nor U10390 (N_10390,N_8463,N_9247);
and U10391 (N_10391,N_8737,N_8832);
or U10392 (N_10392,N_8834,N_9793);
and U10393 (N_10393,N_9334,N_9301);
or U10394 (N_10394,N_8744,N_9037);
nor U10395 (N_10395,N_9166,N_9707);
nor U10396 (N_10396,N_9099,N_8166);
nand U10397 (N_10397,N_9347,N_9202);
and U10398 (N_10398,N_9455,N_8754);
or U10399 (N_10399,N_9697,N_8952);
and U10400 (N_10400,N_8597,N_8136);
nor U10401 (N_10401,N_8666,N_9165);
nand U10402 (N_10402,N_8872,N_8897);
nand U10403 (N_10403,N_9966,N_9583);
and U10404 (N_10404,N_9472,N_8694);
nor U10405 (N_10405,N_9791,N_8037);
or U10406 (N_10406,N_8775,N_9154);
nor U10407 (N_10407,N_8312,N_9749);
and U10408 (N_10408,N_9442,N_9464);
and U10409 (N_10409,N_8893,N_9646);
nand U10410 (N_10410,N_9550,N_9571);
and U10411 (N_10411,N_8461,N_9633);
and U10412 (N_10412,N_8196,N_8290);
xnor U10413 (N_10413,N_9764,N_9316);
or U10414 (N_10414,N_8295,N_9124);
nand U10415 (N_10415,N_9145,N_9122);
nand U10416 (N_10416,N_8578,N_9911);
nand U10417 (N_10417,N_9193,N_8830);
nor U10418 (N_10418,N_9290,N_8500);
nor U10419 (N_10419,N_9186,N_8894);
nor U10420 (N_10420,N_8416,N_8841);
or U10421 (N_10421,N_8570,N_8556);
xnor U10422 (N_10422,N_8632,N_9438);
nand U10423 (N_10423,N_8450,N_8481);
xor U10424 (N_10424,N_8209,N_8840);
or U10425 (N_10425,N_8647,N_8553);
nor U10426 (N_10426,N_9211,N_9637);
nor U10427 (N_10427,N_9238,N_8397);
nor U10428 (N_10428,N_9023,N_9616);
nand U10429 (N_10429,N_9008,N_8215);
or U10430 (N_10430,N_8358,N_8016);
and U10431 (N_10431,N_9172,N_8530);
xnor U10432 (N_10432,N_8101,N_8502);
nand U10433 (N_10433,N_9935,N_8663);
nand U10434 (N_10434,N_9717,N_8195);
nor U10435 (N_10435,N_8151,N_8860);
and U10436 (N_10436,N_8121,N_8695);
or U10437 (N_10437,N_8993,N_8849);
or U10438 (N_10438,N_8743,N_9706);
and U10439 (N_10439,N_9545,N_9426);
nor U10440 (N_10440,N_8219,N_9224);
nand U10441 (N_10441,N_8820,N_9079);
and U10442 (N_10442,N_9969,N_8129);
xor U10443 (N_10443,N_8710,N_8624);
and U10444 (N_10444,N_8029,N_9040);
nand U10445 (N_10445,N_9971,N_9515);
nand U10446 (N_10446,N_9351,N_8575);
nand U10447 (N_10447,N_9980,N_9613);
and U10448 (N_10448,N_8226,N_8097);
or U10449 (N_10449,N_8434,N_9439);
and U10450 (N_10450,N_9305,N_9491);
nand U10451 (N_10451,N_8395,N_9310);
nor U10452 (N_10452,N_9887,N_8917);
nor U10453 (N_10453,N_8342,N_9433);
nand U10454 (N_10454,N_8781,N_9494);
nor U10455 (N_10455,N_8895,N_9209);
and U10456 (N_10456,N_8286,N_9110);
nor U10457 (N_10457,N_8800,N_8105);
and U10458 (N_10458,N_9086,N_8115);
nor U10459 (N_10459,N_9072,N_9449);
nor U10460 (N_10460,N_8030,N_8355);
and U10461 (N_10461,N_9218,N_9174);
nand U10462 (N_10462,N_8989,N_9416);
or U10463 (N_10463,N_8645,N_8914);
nor U10464 (N_10464,N_8341,N_9136);
nor U10465 (N_10465,N_8273,N_9070);
xor U10466 (N_10466,N_9878,N_8001);
nor U10467 (N_10467,N_8347,N_8263);
or U10468 (N_10468,N_9536,N_9245);
nand U10469 (N_10469,N_8759,N_8421);
or U10470 (N_10470,N_8431,N_9641);
nor U10471 (N_10471,N_9581,N_9314);
and U10472 (N_10472,N_8315,N_8244);
nor U10473 (N_10473,N_9675,N_9025);
nor U10474 (N_10474,N_9160,N_9678);
and U10475 (N_10475,N_9600,N_9627);
or U10476 (N_10476,N_9876,N_8758);
nand U10477 (N_10477,N_8282,N_8734);
and U10478 (N_10478,N_8958,N_8329);
and U10479 (N_10479,N_8654,N_9064);
nor U10480 (N_10480,N_9733,N_8751);
nand U10481 (N_10481,N_9944,N_8549);
or U10482 (N_10482,N_8373,N_8823);
or U10483 (N_10483,N_8582,N_9207);
nand U10484 (N_10484,N_8470,N_9391);
xnor U10485 (N_10485,N_9512,N_9441);
nand U10486 (N_10486,N_9977,N_8011);
or U10487 (N_10487,N_9928,N_9033);
nor U10488 (N_10488,N_8616,N_9144);
and U10489 (N_10489,N_8983,N_8227);
nand U10490 (N_10490,N_8944,N_8722);
nor U10491 (N_10491,N_8357,N_8479);
nor U10492 (N_10492,N_9862,N_9689);
nor U10493 (N_10493,N_8048,N_9129);
nor U10494 (N_10494,N_9302,N_9527);
or U10495 (N_10495,N_8247,N_9228);
nand U10496 (N_10496,N_9929,N_8789);
nor U10497 (N_10497,N_9533,N_8352);
or U10498 (N_10498,N_8008,N_9043);
xor U10499 (N_10499,N_8223,N_8004);
nand U10500 (N_10500,N_9054,N_9222);
and U10501 (N_10501,N_9453,N_9462);
nor U10502 (N_10502,N_8565,N_8130);
nand U10503 (N_10503,N_8935,N_9101);
or U10504 (N_10504,N_8788,N_9199);
or U10505 (N_10505,N_9569,N_8370);
or U10506 (N_10506,N_8762,N_9720);
and U10507 (N_10507,N_8301,N_9710);
or U10508 (N_10508,N_8023,N_8901);
xor U10509 (N_10509,N_9213,N_8369);
nor U10510 (N_10510,N_8207,N_9358);
nand U10511 (N_10511,N_8477,N_9615);
nand U10512 (N_10512,N_9951,N_9601);
and U10513 (N_10513,N_9483,N_9588);
nand U10514 (N_10514,N_9103,N_8614);
nand U10515 (N_10515,N_9220,N_9687);
and U10516 (N_10516,N_9653,N_8157);
nand U10517 (N_10517,N_8141,N_8767);
or U10518 (N_10518,N_8615,N_8404);
nand U10519 (N_10519,N_8307,N_9176);
and U10520 (N_10520,N_8721,N_9151);
or U10521 (N_10521,N_8435,N_8797);
or U10522 (N_10522,N_8996,N_9563);
nand U10523 (N_10523,N_8051,N_8580);
or U10524 (N_10524,N_8300,N_9562);
nor U10525 (N_10525,N_8562,N_9885);
nand U10526 (N_10526,N_8534,N_8154);
or U10527 (N_10527,N_8142,N_8764);
nor U10528 (N_10528,N_8599,N_8508);
and U10529 (N_10529,N_8066,N_8592);
xnor U10530 (N_10530,N_8454,N_8975);
or U10531 (N_10531,N_9765,N_8547);
nand U10532 (N_10532,N_8648,N_9766);
nor U10533 (N_10533,N_9105,N_9304);
or U10534 (N_10534,N_9109,N_9959);
and U10535 (N_10535,N_9854,N_8409);
nor U10536 (N_10536,N_9799,N_8971);
and U10537 (N_10537,N_8262,N_8257);
nor U10538 (N_10538,N_9346,N_9288);
and U10539 (N_10539,N_9651,N_8651);
nand U10540 (N_10540,N_8021,N_8179);
nand U10541 (N_10541,N_9322,N_9394);
nand U10542 (N_10542,N_9549,N_8855);
nand U10543 (N_10543,N_8792,N_9747);
or U10544 (N_10544,N_8531,N_8098);
or U10545 (N_10545,N_8883,N_8665);
or U10546 (N_10546,N_8641,N_9053);
xor U10547 (N_10547,N_8224,N_8275);
nor U10548 (N_10548,N_9755,N_9060);
and U10549 (N_10549,N_8197,N_8702);
nor U10550 (N_10550,N_9517,N_9313);
and U10551 (N_10551,N_9939,N_9090);
nand U10552 (N_10552,N_8818,N_9217);
or U10553 (N_10553,N_8203,N_8920);
or U10554 (N_10554,N_9589,N_9384);
and U10555 (N_10555,N_9602,N_8081);
xor U10556 (N_10556,N_8884,N_9208);
or U10557 (N_10557,N_8693,N_8972);
nand U10558 (N_10558,N_8013,N_8802);
xnor U10559 (N_10559,N_8714,N_8736);
nand U10560 (N_10560,N_8193,N_8438);
and U10561 (N_10561,N_8252,N_8425);
nor U10562 (N_10562,N_9547,N_8650);
nor U10563 (N_10563,N_8605,N_9728);
nand U10564 (N_10564,N_8969,N_9920);
xnor U10565 (N_10565,N_8856,N_9212);
or U10566 (N_10566,N_8287,N_9796);
nor U10567 (N_10567,N_9551,N_9104);
xnor U10568 (N_10568,N_9397,N_8418);
and U10569 (N_10569,N_8353,N_8682);
or U10570 (N_10570,N_8609,N_8069);
nor U10571 (N_10571,N_9645,N_8034);
nand U10572 (N_10572,N_9785,N_8133);
nor U10573 (N_10573,N_9342,N_9498);
or U10574 (N_10574,N_8374,N_8923);
nand U10575 (N_10575,N_9560,N_8711);
or U10576 (N_10576,N_8119,N_8700);
xnor U10577 (N_10577,N_8831,N_9411);
or U10578 (N_10578,N_8487,N_8258);
xor U10579 (N_10579,N_8926,N_9044);
or U10580 (N_10580,N_8795,N_9509);
nor U10581 (N_10581,N_9508,N_9420);
xnor U10582 (N_10582,N_8488,N_8078);
and U10583 (N_10583,N_8134,N_8279);
nand U10584 (N_10584,N_9748,N_9192);
or U10585 (N_10585,N_9132,N_8314);
nand U10586 (N_10586,N_9810,N_9873);
nand U10587 (N_10587,N_9578,N_8749);
or U10588 (N_10588,N_8997,N_9867);
nor U10589 (N_10589,N_9647,N_8102);
nand U10590 (N_10590,N_8396,N_8063);
nor U10591 (N_10591,N_8228,N_8033);
or U10592 (N_10592,N_9031,N_9396);
nand U10593 (N_10593,N_8966,N_8899);
nor U10594 (N_10594,N_9577,N_9121);
nand U10595 (N_10595,N_8941,N_8302);
or U10596 (N_10596,N_9309,N_8465);
nor U10597 (N_10597,N_8391,N_9664);
and U10598 (N_10598,N_8636,N_8304);
nand U10599 (N_10599,N_8484,N_9531);
nor U10600 (N_10600,N_8123,N_9856);
and U10601 (N_10601,N_8707,N_8537);
nand U10602 (N_10602,N_9389,N_8533);
nor U10603 (N_10603,N_9700,N_9377);
nand U10604 (N_10604,N_9128,N_8321);
nand U10605 (N_10605,N_9387,N_8361);
nand U10606 (N_10606,N_9567,N_8907);
xnor U10607 (N_10607,N_9440,N_9048);
or U10608 (N_10608,N_8630,N_8740);
xnor U10609 (N_10609,N_8091,N_9961);
nor U10610 (N_10610,N_9648,N_8604);
nand U10611 (N_10611,N_8368,N_9244);
nor U10612 (N_10612,N_8084,N_9682);
and U10613 (N_10613,N_9499,N_8591);
nor U10614 (N_10614,N_9591,N_8185);
nor U10615 (N_10615,N_9894,N_9539);
xor U10616 (N_10616,N_9735,N_8839);
or U10617 (N_10617,N_9026,N_9892);
nand U10618 (N_10618,N_9343,N_9788);
nand U10619 (N_10619,N_9184,N_9418);
nor U10620 (N_10620,N_8497,N_8320);
and U10621 (N_10621,N_9910,N_9355);
nor U10622 (N_10622,N_9703,N_9432);
or U10623 (N_10623,N_8981,N_8010);
nand U10624 (N_10624,N_9826,N_8725);
nor U10625 (N_10625,N_8390,N_8035);
nor U10626 (N_10626,N_8126,N_8960);
nor U10627 (N_10627,N_9049,N_9098);
nand U10628 (N_10628,N_8771,N_8936);
nor U10629 (N_10629,N_9038,N_9246);
nand U10630 (N_10630,N_8796,N_8555);
or U10631 (N_10631,N_8085,N_9180);
nand U10632 (N_10632,N_9901,N_8495);
nor U10633 (N_10633,N_8892,N_8943);
xor U10634 (N_10634,N_8703,N_9088);
and U10635 (N_10635,N_9350,N_9457);
or U10636 (N_10636,N_9197,N_9821);
nor U10637 (N_10637,N_8874,N_9235);
nand U10638 (N_10638,N_8213,N_8336);
nor U10639 (N_10639,N_8221,N_9413);
and U10640 (N_10640,N_8940,N_9576);
and U10641 (N_10641,N_8814,N_9381);
or U10642 (N_10642,N_8076,N_9295);
nor U10643 (N_10643,N_8269,N_8554);
or U10644 (N_10644,N_9450,N_9676);
nor U10645 (N_10645,N_9594,N_8080);
or U10646 (N_10646,N_9732,N_9067);
nor U10647 (N_10647,N_9203,N_9990);
xor U10648 (N_10648,N_8879,N_9471);
nand U10649 (N_10649,N_8210,N_8239);
nor U10650 (N_10650,N_9027,N_8127);
or U10651 (N_10651,N_8683,N_9266);
nor U10652 (N_10652,N_9134,N_9842);
xnor U10653 (N_10653,N_9909,N_9949);
xor U10654 (N_10654,N_9198,N_8719);
or U10655 (N_10655,N_8384,N_8043);
or U10656 (N_10656,N_9273,N_9421);
xor U10657 (N_10657,N_9711,N_9555);
nand U10658 (N_10658,N_9593,N_8643);
nand U10659 (N_10659,N_8088,N_8354);
nor U10660 (N_10660,N_9012,N_8753);
nand U10661 (N_10661,N_8979,N_9926);
and U10662 (N_10662,N_8402,N_8296);
nand U10663 (N_10663,N_9336,N_9866);
and U10664 (N_10664,N_9843,N_9570);
nor U10665 (N_10665,N_8306,N_8364);
and U10666 (N_10666,N_8117,N_8310);
and U10667 (N_10667,N_8898,N_8692);
nand U10668 (N_10668,N_8492,N_8426);
nor U10669 (N_10669,N_8441,N_9392);
and U10670 (N_10670,N_8143,N_9605);
xor U10671 (N_10671,N_9399,N_9276);
nand U10672 (N_10672,N_8672,N_8662);
nand U10673 (N_10673,N_9938,N_8560);
and U10674 (N_10674,N_9708,N_9097);
nor U10675 (N_10675,N_8852,N_9882);
and U10676 (N_10676,N_9366,N_9544);
nor U10677 (N_10677,N_9467,N_8165);
and U10678 (N_10678,N_8995,N_8992);
nand U10679 (N_10679,N_8857,N_9824);
or U10680 (N_10680,N_8988,N_8389);
and U10681 (N_10681,N_8222,N_8718);
nor U10682 (N_10682,N_9798,N_8991);
nor U10683 (N_10683,N_9155,N_8367);
nor U10684 (N_10684,N_9674,N_8427);
nand U10685 (N_10685,N_8729,N_9249);
or U10686 (N_10686,N_9073,N_8162);
and U10687 (N_10687,N_8507,N_8978);
and U10688 (N_10688,N_8644,N_8659);
and U10689 (N_10689,N_9744,N_9523);
nand U10690 (N_10690,N_8875,N_9657);
xor U10691 (N_10691,N_8821,N_9445);
xnor U10692 (N_10692,N_9610,N_9340);
nand U10693 (N_10693,N_9419,N_9307);
or U10694 (N_10694,N_9819,N_9424);
nor U10695 (N_10695,N_9729,N_8288);
and U10696 (N_10696,N_9475,N_8235);
xnor U10697 (N_10697,N_8987,N_9635);
or U10698 (N_10698,N_9306,N_8953);
nand U10699 (N_10699,N_9496,N_8836);
and U10700 (N_10700,N_8932,N_8055);
nor U10701 (N_10701,N_8779,N_9158);
xor U10702 (N_10702,N_9147,N_9281);
and U10703 (N_10703,N_8661,N_8585);
nor U10704 (N_10704,N_9828,N_9835);
xor U10705 (N_10705,N_8947,N_8551);
xnor U10706 (N_10706,N_9754,N_8642);
or U10707 (N_10707,N_8733,N_9521);
or U10708 (N_10708,N_9891,N_8574);
and U10709 (N_10709,N_8691,N_8842);
nor U10710 (N_10710,N_8837,N_8782);
nor U10711 (N_10711,N_9972,N_9632);
and U10712 (N_10712,N_8064,N_9240);
and U10713 (N_10713,N_8266,N_9879);
or U10714 (N_10714,N_8410,N_8998);
nor U10715 (N_10715,N_9771,N_8653);
nor U10716 (N_10716,N_9609,N_8625);
nand U10717 (N_10717,N_9552,N_9546);
nand U10718 (N_10718,N_8326,N_9215);
or U10719 (N_10719,N_8246,N_9331);
and U10720 (N_10720,N_8885,N_8274);
nand U10721 (N_10721,N_9829,N_8876);
or U10722 (N_10722,N_9076,N_9171);
and U10723 (N_10723,N_8200,N_8473);
and U10724 (N_10724,N_9850,N_9932);
and U10725 (N_10725,N_8120,N_8676);
or U10726 (N_10726,N_9353,N_9004);
and U10727 (N_10727,N_8671,N_9505);
xnor U10728 (N_10728,N_8942,N_8000);
and U10729 (N_10729,N_9407,N_9379);
or U10730 (N_10730,N_9093,N_8986);
and U10731 (N_10731,N_9853,N_8318);
nor U10732 (N_10732,N_8900,N_9745);
and U10733 (N_10733,N_9075,N_9185);
nand U10734 (N_10734,N_8231,N_9265);
xor U10735 (N_10735,N_9847,N_9705);
nor U10736 (N_10736,N_8059,N_9694);
or U10737 (N_10737,N_8854,N_8619);
or U10738 (N_10738,N_8294,N_9188);
nor U10739 (N_10739,N_8403,N_9658);
nor U10740 (N_10740,N_8999,N_9858);
nand U10741 (N_10741,N_9608,N_9372);
and U10742 (N_10742,N_9625,N_8937);
nand U10743 (N_10743,N_8681,N_9692);
xnor U10744 (N_10744,N_9456,N_8199);
or U10745 (N_10745,N_8090,N_9914);
nand U10746 (N_10746,N_9315,N_9404);
xnor U10747 (N_10747,N_9428,N_8523);
nor U10748 (N_10748,N_8886,N_9356);
xnor U10749 (N_10749,N_8486,N_9861);
xor U10750 (N_10750,N_8256,N_8925);
nand U10751 (N_10751,N_8873,N_8731);
nand U10752 (N_10752,N_8052,N_9808);
or U10753 (N_10753,N_9425,N_9020);
nand U10754 (N_10754,N_9405,N_9663);
and U10755 (N_10755,N_9135,N_8735);
xnor U10756 (N_10756,N_9942,N_8752);
nand U10757 (N_10757,N_9825,N_9827);
nor U10758 (N_10758,N_8521,N_9630);
nor U10759 (N_10759,N_8082,N_8429);
or U10760 (N_10760,N_9899,N_9886);
nor U10761 (N_10761,N_8985,N_8012);
nand U10762 (N_10762,N_8967,N_8446);
and U10763 (N_10763,N_9139,N_9772);
nor U10764 (N_10764,N_9742,N_8768);
nand U10765 (N_10765,N_9383,N_8182);
nand U10766 (N_10766,N_9401,N_9118);
nand U10767 (N_10767,N_9975,N_8277);
nand U10768 (N_10768,N_8584,N_8062);
and U10769 (N_10769,N_8698,N_8566);
xor U10770 (N_10770,N_8769,N_8827);
and U10771 (N_10771,N_9002,N_8838);
and U10772 (N_10772,N_8928,N_9226);
or U10773 (N_10773,N_9817,N_9834);
and U10774 (N_10774,N_9815,N_9367);
xor U10775 (N_10775,N_9363,N_9339);
nand U10776 (N_10776,N_8137,N_8587);
nor U10777 (N_10777,N_8951,N_9412);
or U10778 (N_10778,N_8026,N_9832);
xor U10779 (N_10779,N_9148,N_8240);
nand U10780 (N_10780,N_9414,N_8948);
and U10781 (N_10781,N_9490,N_9422);
nor U10782 (N_10782,N_8828,N_8444);
nor U10783 (N_10783,N_8973,N_9559);
or U10784 (N_10784,N_8778,N_9525);
nand U10785 (N_10785,N_8079,N_8738);
or U10786 (N_10786,N_9573,N_8476);
or U10787 (N_10787,N_8378,N_8878);
or U10788 (N_10788,N_9784,N_8617);
and U10789 (N_10789,N_9091,N_8601);
nor U10790 (N_10790,N_9320,N_9429);
xor U10791 (N_10791,N_8757,N_9968);
nor U10792 (N_10792,N_9870,N_8811);
and U10793 (N_10793,N_9797,N_8573);
xor U10794 (N_10794,N_9107,N_9730);
nor U10795 (N_10795,N_8687,N_8791);
nor U10796 (N_10796,N_8664,N_9965);
nand U10797 (N_10797,N_9022,N_8006);
nor U10798 (N_10798,N_8745,N_9553);
nor U10799 (N_10799,N_8826,N_8171);
nor U10800 (N_10800,N_9236,N_8180);
xnor U10801 (N_10801,N_8825,N_9319);
xnor U10802 (N_10802,N_9285,N_9430);
nor U10803 (N_10803,N_9690,N_9599);
nor U10804 (N_10804,N_8096,N_9476);
xor U10805 (N_10805,N_9286,N_8118);
xnor U10806 (N_10806,N_9164,N_9140);
and U10807 (N_10807,N_9918,N_9958);
or U10808 (N_10808,N_8522,N_8793);
and U10809 (N_10809,N_9444,N_9150);
and U10810 (N_10810,N_8709,N_9015);
and U10811 (N_10811,N_9794,N_8089);
nor U10812 (N_10812,N_9660,N_8785);
or U10813 (N_10813,N_9513,N_9921);
or U10814 (N_10814,N_9695,N_9431);
and U10815 (N_10815,N_8420,N_9933);
or U10816 (N_10816,N_8542,N_9987);
xor U10817 (N_10817,N_8824,N_9999);
and U10818 (N_10818,N_8913,N_8911);
nand U10819 (N_10819,N_9607,N_9382);
nor U10820 (N_10820,N_9762,N_9255);
and U10821 (N_10821,N_8139,N_9737);
nor U10822 (N_10822,N_9541,N_9047);
or U10823 (N_10823,N_9200,N_9777);
nand U10824 (N_10824,N_8805,N_8337);
and U10825 (N_10825,N_8888,N_8039);
nor U10826 (N_10826,N_8557,N_9988);
or U10827 (N_10827,N_9783,N_9036);
xnor U10828 (N_10828,N_8330,N_8394);
or U10829 (N_10829,N_9813,N_9461);
xnor U10830 (N_10830,N_8593,N_8965);
xor U10831 (N_10831,N_8777,N_9251);
and U10832 (N_10832,N_9169,N_9941);
and U10833 (N_10833,N_9162,N_8808);
nand U10834 (N_10834,N_8491,N_8623);
nor U10835 (N_10835,N_9500,N_9903);
xor U10836 (N_10836,N_9016,N_9913);
nand U10837 (N_10837,N_9787,N_8620);
nand U10838 (N_10838,N_9943,N_8343);
nor U10839 (N_10839,N_9058,N_8977);
nand U10840 (N_10840,N_9329,N_9046);
and U10841 (N_10841,N_9359,N_9722);
and U10842 (N_10842,N_8773,N_8340);
and U10843 (N_10843,N_9250,N_8359);
nand U10844 (N_10844,N_8103,N_9317);
xor U10845 (N_10845,N_8902,N_9652);
nand U10846 (N_10846,N_9168,N_8701);
and U10847 (N_10847,N_9274,N_9566);
or U10848 (N_10848,N_9634,N_9738);
or U10849 (N_10849,N_9021,N_9279);
or U10850 (N_10850,N_9287,N_8699);
and U10851 (N_10851,N_8474,N_9234);
nor U10852 (N_10852,N_8122,N_9146);
nor U10853 (N_10853,N_8677,N_9983);
xnor U10854 (N_10854,N_8439,N_8241);
nor U10855 (N_10855,N_9656,N_9540);
and U10856 (N_10856,N_8413,N_9117);
nand U10857 (N_10857,N_9484,N_8164);
nor U10858 (N_10858,N_9360,N_9268);
nor U10859 (N_10859,N_9631,N_8293);
and U10860 (N_10860,N_9883,N_8025);
nor U10861 (N_10861,N_8255,N_9436);
nor U10862 (N_10862,N_9275,N_8181);
or U10863 (N_10863,N_8546,N_8110);
nor U10864 (N_10864,N_9756,N_9189);
nand U10865 (N_10865,N_9592,N_8889);
nor U10866 (N_10866,N_9216,N_9349);
nor U10867 (N_10867,N_8871,N_9504);
and U10868 (N_10868,N_8939,N_8813);
xor U10869 (N_10869,N_9906,N_8381);
nor U10870 (N_10870,N_8111,N_8248);
or U10871 (N_10871,N_8904,N_8931);
xor U10872 (N_10872,N_8660,N_8268);
nor U10873 (N_10873,N_8135,N_9800);
and U10874 (N_10874,N_9683,N_8187);
nor U10875 (N_10875,N_9823,N_8150);
and U10876 (N_10876,N_9354,N_8611);
xnor U10877 (N_10877,N_9614,N_8629);
nor U10878 (N_10878,N_8346,N_9254);
nand U10879 (N_10879,N_9715,N_8116);
nor U10880 (N_10880,N_9612,N_8550);
nand U10881 (N_10881,N_8572,N_8957);
or U10882 (N_10882,N_8563,N_9818);
nor U10883 (N_10883,N_8535,N_8237);
nor U10884 (N_10884,N_8173,N_8093);
nor U10885 (N_10885,N_9388,N_8456);
nor U10886 (N_10886,N_9327,N_8003);
nor U10887 (N_10887,N_9685,N_9912);
nand U10888 (N_10888,N_9830,N_9507);
or U10889 (N_10889,N_9196,N_8053);
nand U10890 (N_10890,N_9503,N_9402);
and U10891 (N_10891,N_8202,N_8242);
and U10892 (N_10892,N_9557,N_9014);
and U10893 (N_10893,N_8345,N_8014);
and U10894 (N_10894,N_9157,N_9849);
or U10895 (N_10895,N_8607,N_9050);
nor U10896 (N_10896,N_9473,N_8822);
or U10897 (N_10897,N_9731,N_8766);
nand U10898 (N_10898,N_9187,N_9143);
nor U10899 (N_10899,N_9670,N_8289);
nor U10900 (N_10900,N_9497,N_9753);
nor U10901 (N_10901,N_9618,N_8156);
and U10902 (N_10902,N_8009,N_9704);
nand U10903 (N_10903,N_8761,N_9241);
nand U10904 (N_10904,N_9859,N_8924);
or U10905 (N_10905,N_8867,N_8602);
xor U10906 (N_10906,N_9998,N_8970);
and U10907 (N_10907,N_8338,N_9269);
or U10908 (N_10908,N_9629,N_8160);
or U10909 (N_10909,N_8848,N_9019);
and U10910 (N_10910,N_9227,N_9006);
or U10911 (N_10911,N_8186,N_9953);
nor U10912 (N_10912,N_8437,N_9575);
nor U10913 (N_10913,N_8804,N_8432);
nand U10914 (N_10914,N_9095,N_8414);
and U10915 (N_10915,N_9930,N_8073);
and U10916 (N_10916,N_9230,N_9923);
and U10917 (N_10917,N_9623,N_8297);
and U10918 (N_10918,N_8424,N_8513);
nor U10919 (N_10919,N_8276,N_8469);
nor U10920 (N_10920,N_8245,N_9190);
or U10921 (N_10921,N_8138,N_8489);
or U10922 (N_10922,N_8007,N_9345);
and U10923 (N_10923,N_8415,N_9568);
nand U10924 (N_10924,N_8075,N_8028);
and U10925 (N_10925,N_8859,N_8526);
or U10926 (N_10926,N_9039,N_8238);
xnor U10927 (N_10927,N_9029,N_8596);
nor U10928 (N_10928,N_8723,N_8071);
nor U10929 (N_10929,N_8251,N_9727);
nor U10930 (N_10930,N_8847,N_8896);
nor U10931 (N_10931,N_9089,N_9466);
nand U10932 (N_10932,N_8452,N_8982);
or U10933 (N_10933,N_8525,N_8385);
nand U10934 (N_10934,N_8780,N_8284);
or U10935 (N_10935,N_8149,N_8460);
or U10936 (N_10936,N_9017,N_8260);
xnor U10937 (N_10937,N_8870,N_9661);
nor U10938 (N_10938,N_8853,N_9839);
or U10939 (N_10939,N_9156,N_8331);
nor U10940 (N_10940,N_9948,N_9223);
or U10941 (N_10941,N_8518,N_9831);
or U10942 (N_10942,N_8086,N_9845);
nand U10943 (N_10943,N_9460,N_9161);
or U10944 (N_10944,N_8955,N_8398);
nor U10945 (N_10945,N_8835,N_9062);
nor U10946 (N_10946,N_9007,N_8594);
and U10947 (N_10947,N_8159,N_9750);
nand U10948 (N_10948,N_9114,N_8589);
and U10949 (N_10949,N_9677,N_8351);
nor U10950 (N_10950,N_8728,N_8829);
or U10951 (N_10951,N_8690,N_9325);
or U10952 (N_10952,N_8208,N_8845);
nand U10953 (N_10953,N_9804,N_9596);
or U10954 (N_10954,N_9378,N_9258);
and U10955 (N_10955,N_8918,N_9833);
xnor U10956 (N_10956,N_8933,N_8230);
or U10957 (N_10957,N_8812,N_8880);
and U10958 (N_10958,N_8158,N_8036);
xnor U10959 (N_10959,N_9537,N_8787);
or U10960 (N_10960,N_8806,N_8114);
nor U10961 (N_10961,N_9065,N_8524);
or U10962 (N_10962,N_8175,N_9716);
or U10963 (N_10963,N_9051,N_8657);
nor U10964 (N_10964,N_9638,N_8440);
xor U10965 (N_10965,N_8882,N_9776);
and U10966 (N_10966,N_9997,N_9574);
xor U10967 (N_10967,N_8588,N_9590);
or U10968 (N_10968,N_8401,N_8610);
and U10969 (N_10969,N_8720,N_8716);
or U10970 (N_10970,N_8065,N_9734);
or U10971 (N_10971,N_8303,N_8715);
or U10972 (N_10972,N_8851,N_9781);
nand U10973 (N_10973,N_9149,N_9587);
or U10974 (N_10974,N_8961,N_9604);
nor U10975 (N_10975,N_8501,N_8412);
and U10976 (N_10976,N_9769,N_9374);
and U10977 (N_10977,N_9688,N_9120);
nor U10978 (N_10978,N_9554,N_8794);
or U10979 (N_10979,N_8448,N_8380);
or U10980 (N_10980,N_8798,N_9580);
and U10981 (N_10981,N_9369,N_9292);
or U10982 (N_10982,N_8388,N_9741);
and U10983 (N_10983,N_8146,N_9895);
or U10984 (N_10984,N_9672,N_9357);
xnor U10985 (N_10985,N_8261,N_9175);
or U10986 (N_10986,N_8430,N_8100);
nand U10987 (N_10987,N_9082,N_8633);
or U10988 (N_10988,N_9543,N_8124);
nand U10989 (N_10989,N_8271,N_8921);
nand U10990 (N_10990,N_9723,N_9296);
nand U10991 (N_10991,N_8649,N_9931);
nor U10992 (N_10992,N_8044,N_8577);
nor U10993 (N_10993,N_9123,N_9908);
nor U10994 (N_10994,N_9770,N_8519);
nor U10995 (N_10995,N_8536,N_8667);
nor U10996 (N_10996,N_9579,N_9370);
nor U10997 (N_10997,N_9518,N_9011);
and U10998 (N_10998,N_8407,N_9907);
xor U10999 (N_10999,N_9119,N_9092);
nor U11000 (N_11000,N_9239,N_9015);
or U11001 (N_11001,N_9714,N_9975);
and U11002 (N_11002,N_9490,N_8469);
nor U11003 (N_11003,N_8634,N_9740);
nand U11004 (N_11004,N_8856,N_8190);
nor U11005 (N_11005,N_8196,N_9990);
nor U11006 (N_11006,N_8068,N_8561);
nand U11007 (N_11007,N_8593,N_8300);
and U11008 (N_11008,N_8996,N_8478);
nor U11009 (N_11009,N_8512,N_8896);
nand U11010 (N_11010,N_8782,N_9239);
or U11011 (N_11011,N_9476,N_9776);
or U11012 (N_11012,N_9859,N_8321);
nor U11013 (N_11013,N_8788,N_8879);
or U11014 (N_11014,N_9020,N_9481);
and U11015 (N_11015,N_9748,N_8899);
nor U11016 (N_11016,N_9302,N_9593);
or U11017 (N_11017,N_8314,N_8014);
and U11018 (N_11018,N_9924,N_9223);
xnor U11019 (N_11019,N_8118,N_9935);
or U11020 (N_11020,N_9104,N_8521);
or U11021 (N_11021,N_8902,N_9026);
nor U11022 (N_11022,N_8602,N_9646);
or U11023 (N_11023,N_8002,N_9621);
nand U11024 (N_11024,N_9379,N_9722);
nor U11025 (N_11025,N_9765,N_9389);
nor U11026 (N_11026,N_9853,N_9686);
nand U11027 (N_11027,N_9584,N_9264);
or U11028 (N_11028,N_8321,N_9842);
xnor U11029 (N_11029,N_8718,N_8332);
and U11030 (N_11030,N_9358,N_9122);
and U11031 (N_11031,N_8161,N_8982);
or U11032 (N_11032,N_8618,N_8077);
nand U11033 (N_11033,N_8205,N_9119);
or U11034 (N_11034,N_8859,N_9559);
nor U11035 (N_11035,N_9012,N_8680);
and U11036 (N_11036,N_9936,N_9812);
and U11037 (N_11037,N_8892,N_8472);
and U11038 (N_11038,N_8504,N_8962);
and U11039 (N_11039,N_9209,N_8704);
xor U11040 (N_11040,N_8988,N_9877);
nand U11041 (N_11041,N_9264,N_9657);
or U11042 (N_11042,N_9555,N_8965);
and U11043 (N_11043,N_9251,N_8868);
or U11044 (N_11044,N_8170,N_9845);
and U11045 (N_11045,N_8565,N_8072);
xor U11046 (N_11046,N_9746,N_9530);
xnor U11047 (N_11047,N_9992,N_8564);
nand U11048 (N_11048,N_8488,N_9918);
and U11049 (N_11049,N_8268,N_9312);
nand U11050 (N_11050,N_8201,N_9429);
nand U11051 (N_11051,N_9172,N_9693);
and U11052 (N_11052,N_8128,N_8108);
nand U11053 (N_11053,N_9073,N_9467);
or U11054 (N_11054,N_8060,N_8121);
nand U11055 (N_11055,N_8809,N_9672);
and U11056 (N_11056,N_9475,N_8116);
xnor U11057 (N_11057,N_8469,N_8789);
nor U11058 (N_11058,N_9036,N_9878);
nor U11059 (N_11059,N_8840,N_9815);
nand U11060 (N_11060,N_8847,N_9510);
nor U11061 (N_11061,N_8956,N_8428);
nand U11062 (N_11062,N_8449,N_8494);
and U11063 (N_11063,N_8112,N_8896);
and U11064 (N_11064,N_8920,N_9752);
xor U11065 (N_11065,N_9725,N_8703);
nand U11066 (N_11066,N_8142,N_9609);
and U11067 (N_11067,N_9497,N_9737);
nand U11068 (N_11068,N_8047,N_9647);
or U11069 (N_11069,N_8866,N_8413);
or U11070 (N_11070,N_9543,N_8428);
and U11071 (N_11071,N_9427,N_8789);
and U11072 (N_11072,N_8352,N_9418);
or U11073 (N_11073,N_8013,N_8525);
or U11074 (N_11074,N_8352,N_8814);
or U11075 (N_11075,N_8421,N_8452);
or U11076 (N_11076,N_9903,N_8512);
or U11077 (N_11077,N_9335,N_8650);
and U11078 (N_11078,N_8036,N_8550);
and U11079 (N_11079,N_8416,N_8650);
xor U11080 (N_11080,N_9140,N_8871);
nor U11081 (N_11081,N_8638,N_9484);
or U11082 (N_11082,N_9016,N_9204);
and U11083 (N_11083,N_9338,N_8288);
nand U11084 (N_11084,N_8952,N_8415);
nor U11085 (N_11085,N_9643,N_8501);
or U11086 (N_11086,N_9169,N_9322);
or U11087 (N_11087,N_8771,N_8129);
xnor U11088 (N_11088,N_9198,N_9879);
and U11089 (N_11089,N_8777,N_9944);
or U11090 (N_11090,N_9154,N_8185);
and U11091 (N_11091,N_8707,N_8367);
nand U11092 (N_11092,N_8983,N_8259);
nand U11093 (N_11093,N_9893,N_8671);
nor U11094 (N_11094,N_8482,N_9700);
or U11095 (N_11095,N_9232,N_9944);
nor U11096 (N_11096,N_9538,N_9272);
nand U11097 (N_11097,N_9106,N_9688);
and U11098 (N_11098,N_8277,N_9727);
xor U11099 (N_11099,N_8191,N_8313);
nor U11100 (N_11100,N_9828,N_8477);
and U11101 (N_11101,N_8560,N_9504);
and U11102 (N_11102,N_8387,N_8126);
xnor U11103 (N_11103,N_8288,N_8881);
xor U11104 (N_11104,N_8770,N_8927);
or U11105 (N_11105,N_8183,N_9736);
or U11106 (N_11106,N_8306,N_8518);
nor U11107 (N_11107,N_8600,N_8524);
and U11108 (N_11108,N_9864,N_8686);
or U11109 (N_11109,N_8723,N_9555);
nand U11110 (N_11110,N_9612,N_8713);
or U11111 (N_11111,N_8080,N_8737);
xnor U11112 (N_11112,N_8799,N_8581);
nand U11113 (N_11113,N_8410,N_8336);
xor U11114 (N_11114,N_8266,N_9535);
xnor U11115 (N_11115,N_8643,N_8195);
nor U11116 (N_11116,N_8171,N_8218);
nor U11117 (N_11117,N_8122,N_8974);
and U11118 (N_11118,N_9363,N_8212);
or U11119 (N_11119,N_9075,N_9424);
and U11120 (N_11120,N_9424,N_9711);
or U11121 (N_11121,N_9326,N_9315);
xor U11122 (N_11122,N_8927,N_8332);
and U11123 (N_11123,N_9375,N_9887);
and U11124 (N_11124,N_9803,N_9485);
and U11125 (N_11125,N_8383,N_9624);
nor U11126 (N_11126,N_9706,N_9696);
nand U11127 (N_11127,N_8307,N_8383);
and U11128 (N_11128,N_8563,N_8413);
xor U11129 (N_11129,N_9285,N_8029);
nand U11130 (N_11130,N_9040,N_9421);
xnor U11131 (N_11131,N_8400,N_8248);
nand U11132 (N_11132,N_9967,N_8059);
xor U11133 (N_11133,N_9385,N_8535);
nand U11134 (N_11134,N_9720,N_8066);
or U11135 (N_11135,N_8972,N_9285);
nand U11136 (N_11136,N_8047,N_9433);
and U11137 (N_11137,N_9903,N_9824);
xor U11138 (N_11138,N_8639,N_8994);
or U11139 (N_11139,N_9544,N_8608);
nand U11140 (N_11140,N_9997,N_8213);
nor U11141 (N_11141,N_9078,N_9516);
and U11142 (N_11142,N_9221,N_9102);
nor U11143 (N_11143,N_8287,N_8808);
and U11144 (N_11144,N_8269,N_8738);
nand U11145 (N_11145,N_8565,N_9745);
and U11146 (N_11146,N_8064,N_9868);
and U11147 (N_11147,N_9686,N_9728);
nor U11148 (N_11148,N_8595,N_8358);
nand U11149 (N_11149,N_8739,N_9740);
and U11150 (N_11150,N_8497,N_9982);
or U11151 (N_11151,N_8548,N_9723);
or U11152 (N_11152,N_9983,N_8681);
or U11153 (N_11153,N_9008,N_8343);
and U11154 (N_11154,N_9882,N_8141);
nor U11155 (N_11155,N_8894,N_8122);
xor U11156 (N_11156,N_8272,N_9249);
nor U11157 (N_11157,N_9993,N_9926);
xnor U11158 (N_11158,N_8617,N_9081);
and U11159 (N_11159,N_9148,N_9671);
and U11160 (N_11160,N_9903,N_8943);
nand U11161 (N_11161,N_8591,N_8206);
and U11162 (N_11162,N_9758,N_8098);
or U11163 (N_11163,N_8782,N_9670);
or U11164 (N_11164,N_9680,N_9069);
xnor U11165 (N_11165,N_9274,N_9511);
or U11166 (N_11166,N_9812,N_9120);
and U11167 (N_11167,N_8913,N_8624);
nor U11168 (N_11168,N_8537,N_9976);
xor U11169 (N_11169,N_8617,N_9777);
nor U11170 (N_11170,N_8064,N_9252);
and U11171 (N_11171,N_8903,N_8643);
nor U11172 (N_11172,N_9138,N_8676);
nand U11173 (N_11173,N_8576,N_9693);
or U11174 (N_11174,N_8712,N_8553);
and U11175 (N_11175,N_8536,N_8275);
nor U11176 (N_11176,N_9051,N_8166);
or U11177 (N_11177,N_8748,N_8545);
and U11178 (N_11178,N_9786,N_9533);
xnor U11179 (N_11179,N_8868,N_9131);
nor U11180 (N_11180,N_9901,N_8112);
xor U11181 (N_11181,N_8741,N_9216);
and U11182 (N_11182,N_9819,N_9540);
or U11183 (N_11183,N_9362,N_9457);
and U11184 (N_11184,N_8846,N_8652);
and U11185 (N_11185,N_9495,N_9412);
or U11186 (N_11186,N_8591,N_9275);
nand U11187 (N_11187,N_8721,N_9460);
nand U11188 (N_11188,N_8322,N_8818);
nand U11189 (N_11189,N_8904,N_8529);
or U11190 (N_11190,N_9596,N_8954);
nand U11191 (N_11191,N_8293,N_9144);
nor U11192 (N_11192,N_8578,N_8301);
nand U11193 (N_11193,N_9215,N_8023);
xnor U11194 (N_11194,N_9886,N_9820);
nor U11195 (N_11195,N_9852,N_8323);
or U11196 (N_11196,N_9747,N_9738);
and U11197 (N_11197,N_9053,N_8536);
and U11198 (N_11198,N_8405,N_8851);
nand U11199 (N_11199,N_8852,N_8771);
nor U11200 (N_11200,N_9768,N_9146);
or U11201 (N_11201,N_9088,N_8834);
nor U11202 (N_11202,N_9404,N_8456);
nand U11203 (N_11203,N_8117,N_9299);
nand U11204 (N_11204,N_8327,N_9596);
nor U11205 (N_11205,N_9598,N_9836);
nand U11206 (N_11206,N_8525,N_8928);
and U11207 (N_11207,N_8047,N_9133);
nor U11208 (N_11208,N_8465,N_8460);
nor U11209 (N_11209,N_8348,N_9650);
nand U11210 (N_11210,N_8849,N_9410);
nand U11211 (N_11211,N_8842,N_9821);
nand U11212 (N_11212,N_8875,N_9091);
nor U11213 (N_11213,N_9018,N_8041);
xnor U11214 (N_11214,N_9344,N_9855);
nand U11215 (N_11215,N_8664,N_8818);
nand U11216 (N_11216,N_9235,N_8389);
and U11217 (N_11217,N_9266,N_9345);
nor U11218 (N_11218,N_9755,N_9229);
nand U11219 (N_11219,N_8253,N_9625);
xnor U11220 (N_11220,N_8642,N_8509);
xor U11221 (N_11221,N_9460,N_9874);
nand U11222 (N_11222,N_8311,N_8792);
nor U11223 (N_11223,N_9406,N_8517);
nand U11224 (N_11224,N_9931,N_8173);
and U11225 (N_11225,N_9931,N_9809);
or U11226 (N_11226,N_8991,N_9197);
nor U11227 (N_11227,N_8606,N_9547);
and U11228 (N_11228,N_9660,N_9041);
and U11229 (N_11229,N_8159,N_8669);
nor U11230 (N_11230,N_9303,N_8249);
and U11231 (N_11231,N_8471,N_9845);
and U11232 (N_11232,N_9422,N_8854);
and U11233 (N_11233,N_8288,N_9891);
nand U11234 (N_11234,N_9406,N_9951);
xnor U11235 (N_11235,N_8895,N_9975);
nor U11236 (N_11236,N_9062,N_9072);
nand U11237 (N_11237,N_9134,N_9130);
xnor U11238 (N_11238,N_8084,N_9020);
or U11239 (N_11239,N_8865,N_8491);
and U11240 (N_11240,N_8368,N_9309);
nand U11241 (N_11241,N_8961,N_9914);
or U11242 (N_11242,N_8628,N_9864);
nor U11243 (N_11243,N_9781,N_8089);
and U11244 (N_11244,N_9788,N_9034);
nand U11245 (N_11245,N_9410,N_9986);
or U11246 (N_11246,N_8994,N_8268);
nand U11247 (N_11247,N_8637,N_8990);
xor U11248 (N_11248,N_8474,N_8895);
and U11249 (N_11249,N_9544,N_8634);
nor U11250 (N_11250,N_9643,N_9749);
and U11251 (N_11251,N_9915,N_9008);
nor U11252 (N_11252,N_9325,N_8039);
xnor U11253 (N_11253,N_9243,N_9529);
and U11254 (N_11254,N_8698,N_8991);
and U11255 (N_11255,N_8550,N_8730);
or U11256 (N_11256,N_8403,N_9710);
nand U11257 (N_11257,N_9314,N_8239);
nand U11258 (N_11258,N_8668,N_8844);
or U11259 (N_11259,N_8652,N_9395);
nand U11260 (N_11260,N_8393,N_9863);
nor U11261 (N_11261,N_8987,N_8153);
nor U11262 (N_11262,N_9575,N_9035);
or U11263 (N_11263,N_8100,N_9331);
nor U11264 (N_11264,N_9493,N_9370);
nor U11265 (N_11265,N_8300,N_9656);
nand U11266 (N_11266,N_8030,N_9306);
nand U11267 (N_11267,N_8895,N_9014);
nand U11268 (N_11268,N_9974,N_8634);
nand U11269 (N_11269,N_8910,N_8959);
nand U11270 (N_11270,N_9465,N_9006);
and U11271 (N_11271,N_8372,N_8487);
and U11272 (N_11272,N_9368,N_9227);
nor U11273 (N_11273,N_9875,N_9480);
and U11274 (N_11274,N_8911,N_9128);
nand U11275 (N_11275,N_8616,N_8409);
or U11276 (N_11276,N_8101,N_9287);
and U11277 (N_11277,N_9512,N_9816);
xnor U11278 (N_11278,N_9535,N_9766);
or U11279 (N_11279,N_9235,N_9159);
nand U11280 (N_11280,N_8904,N_9493);
xnor U11281 (N_11281,N_9414,N_9547);
or U11282 (N_11282,N_9606,N_9333);
and U11283 (N_11283,N_9917,N_8563);
nor U11284 (N_11284,N_9428,N_8828);
xnor U11285 (N_11285,N_8188,N_9361);
and U11286 (N_11286,N_8463,N_9053);
nand U11287 (N_11287,N_8465,N_9332);
or U11288 (N_11288,N_8349,N_8772);
xnor U11289 (N_11289,N_9746,N_8252);
nor U11290 (N_11290,N_9629,N_9214);
and U11291 (N_11291,N_8180,N_8695);
xnor U11292 (N_11292,N_9581,N_9033);
or U11293 (N_11293,N_9673,N_8257);
or U11294 (N_11294,N_9576,N_8793);
nor U11295 (N_11295,N_9145,N_9580);
and U11296 (N_11296,N_9346,N_8039);
nor U11297 (N_11297,N_8495,N_8614);
or U11298 (N_11298,N_8650,N_8212);
nand U11299 (N_11299,N_9565,N_8656);
nor U11300 (N_11300,N_8963,N_8522);
nand U11301 (N_11301,N_9205,N_8734);
or U11302 (N_11302,N_8978,N_8244);
and U11303 (N_11303,N_9990,N_8872);
nor U11304 (N_11304,N_8490,N_8024);
and U11305 (N_11305,N_8392,N_8673);
nor U11306 (N_11306,N_9315,N_9361);
nor U11307 (N_11307,N_8740,N_8304);
nor U11308 (N_11308,N_8556,N_9049);
nor U11309 (N_11309,N_8553,N_9631);
nor U11310 (N_11310,N_9051,N_9516);
nand U11311 (N_11311,N_8458,N_8763);
xnor U11312 (N_11312,N_9995,N_8090);
and U11313 (N_11313,N_9928,N_8052);
or U11314 (N_11314,N_9958,N_8521);
or U11315 (N_11315,N_8786,N_9678);
and U11316 (N_11316,N_8352,N_8204);
and U11317 (N_11317,N_9196,N_8017);
nor U11318 (N_11318,N_9395,N_9977);
nand U11319 (N_11319,N_9954,N_8533);
nor U11320 (N_11320,N_9017,N_9763);
and U11321 (N_11321,N_8735,N_9537);
nor U11322 (N_11322,N_8567,N_9834);
nand U11323 (N_11323,N_9911,N_8611);
or U11324 (N_11324,N_9105,N_9750);
or U11325 (N_11325,N_9270,N_8883);
or U11326 (N_11326,N_8375,N_9666);
nand U11327 (N_11327,N_9698,N_9433);
or U11328 (N_11328,N_9371,N_8597);
and U11329 (N_11329,N_9583,N_9065);
nand U11330 (N_11330,N_9303,N_8722);
nor U11331 (N_11331,N_8587,N_8048);
nor U11332 (N_11332,N_9939,N_8272);
nand U11333 (N_11333,N_9747,N_8148);
or U11334 (N_11334,N_9526,N_9133);
or U11335 (N_11335,N_9164,N_9778);
nand U11336 (N_11336,N_9905,N_9666);
nand U11337 (N_11337,N_8657,N_9318);
nor U11338 (N_11338,N_9973,N_9722);
nor U11339 (N_11339,N_8994,N_8944);
xor U11340 (N_11340,N_9607,N_8302);
nand U11341 (N_11341,N_9067,N_9387);
and U11342 (N_11342,N_8898,N_9472);
or U11343 (N_11343,N_8099,N_9314);
and U11344 (N_11344,N_9501,N_9623);
nor U11345 (N_11345,N_9182,N_8161);
or U11346 (N_11346,N_9731,N_8385);
and U11347 (N_11347,N_9029,N_9773);
xnor U11348 (N_11348,N_9488,N_9556);
nand U11349 (N_11349,N_9190,N_9162);
xor U11350 (N_11350,N_9310,N_8072);
nand U11351 (N_11351,N_9022,N_8358);
or U11352 (N_11352,N_9436,N_8673);
and U11353 (N_11353,N_9588,N_8728);
nor U11354 (N_11354,N_8310,N_8078);
nor U11355 (N_11355,N_8016,N_9600);
nor U11356 (N_11356,N_9329,N_8303);
or U11357 (N_11357,N_8266,N_9222);
xnor U11358 (N_11358,N_8988,N_8871);
or U11359 (N_11359,N_9264,N_9543);
or U11360 (N_11360,N_8771,N_9238);
or U11361 (N_11361,N_9984,N_8366);
nand U11362 (N_11362,N_8012,N_9476);
nand U11363 (N_11363,N_9905,N_8371);
nor U11364 (N_11364,N_9627,N_9692);
or U11365 (N_11365,N_8935,N_9588);
nor U11366 (N_11366,N_8299,N_9189);
and U11367 (N_11367,N_9203,N_9679);
and U11368 (N_11368,N_9804,N_9781);
nor U11369 (N_11369,N_9133,N_8771);
nor U11370 (N_11370,N_9535,N_8397);
or U11371 (N_11371,N_9649,N_8886);
and U11372 (N_11372,N_8761,N_8727);
nor U11373 (N_11373,N_8185,N_8574);
nand U11374 (N_11374,N_8327,N_8663);
and U11375 (N_11375,N_9839,N_8308);
nand U11376 (N_11376,N_8600,N_9378);
and U11377 (N_11377,N_9303,N_9680);
nand U11378 (N_11378,N_9327,N_8610);
nand U11379 (N_11379,N_8125,N_8757);
or U11380 (N_11380,N_8117,N_9076);
nor U11381 (N_11381,N_8920,N_9345);
or U11382 (N_11382,N_9890,N_8336);
nor U11383 (N_11383,N_8001,N_8271);
xnor U11384 (N_11384,N_9335,N_9021);
or U11385 (N_11385,N_9363,N_8749);
nand U11386 (N_11386,N_9775,N_8693);
nand U11387 (N_11387,N_8558,N_8889);
or U11388 (N_11388,N_8082,N_8042);
nand U11389 (N_11389,N_8214,N_8610);
and U11390 (N_11390,N_8863,N_8285);
or U11391 (N_11391,N_8262,N_9286);
or U11392 (N_11392,N_8276,N_8705);
nor U11393 (N_11393,N_9430,N_8015);
and U11394 (N_11394,N_8936,N_8111);
and U11395 (N_11395,N_9031,N_9921);
and U11396 (N_11396,N_8332,N_9014);
or U11397 (N_11397,N_9993,N_9334);
or U11398 (N_11398,N_8576,N_8904);
or U11399 (N_11399,N_9176,N_9873);
nor U11400 (N_11400,N_9394,N_9773);
nor U11401 (N_11401,N_8759,N_9080);
nand U11402 (N_11402,N_9119,N_8089);
nand U11403 (N_11403,N_9391,N_9225);
nor U11404 (N_11404,N_9262,N_8913);
xor U11405 (N_11405,N_9394,N_8519);
and U11406 (N_11406,N_8535,N_8101);
or U11407 (N_11407,N_8477,N_8764);
nor U11408 (N_11408,N_8570,N_9748);
or U11409 (N_11409,N_9786,N_9424);
nand U11410 (N_11410,N_9719,N_8769);
or U11411 (N_11411,N_8002,N_8912);
or U11412 (N_11412,N_9282,N_9700);
xnor U11413 (N_11413,N_9776,N_8269);
xor U11414 (N_11414,N_9562,N_8559);
or U11415 (N_11415,N_9133,N_9666);
or U11416 (N_11416,N_8987,N_9567);
nor U11417 (N_11417,N_9572,N_9320);
nand U11418 (N_11418,N_8940,N_9979);
and U11419 (N_11419,N_9503,N_9107);
nand U11420 (N_11420,N_9593,N_8256);
nor U11421 (N_11421,N_9936,N_8327);
and U11422 (N_11422,N_9634,N_8344);
and U11423 (N_11423,N_9753,N_9738);
xor U11424 (N_11424,N_9167,N_8950);
or U11425 (N_11425,N_9489,N_8912);
or U11426 (N_11426,N_9407,N_8994);
nand U11427 (N_11427,N_9832,N_9154);
or U11428 (N_11428,N_9976,N_9400);
or U11429 (N_11429,N_8970,N_9587);
nand U11430 (N_11430,N_9899,N_8744);
xor U11431 (N_11431,N_9050,N_9506);
or U11432 (N_11432,N_8854,N_8254);
or U11433 (N_11433,N_8414,N_9595);
nor U11434 (N_11434,N_8426,N_8057);
nand U11435 (N_11435,N_8398,N_9955);
and U11436 (N_11436,N_9312,N_9254);
nor U11437 (N_11437,N_9696,N_9904);
or U11438 (N_11438,N_9149,N_9740);
nand U11439 (N_11439,N_9039,N_9228);
nand U11440 (N_11440,N_9220,N_8226);
nand U11441 (N_11441,N_9644,N_9498);
xnor U11442 (N_11442,N_8877,N_8677);
or U11443 (N_11443,N_9557,N_8297);
nor U11444 (N_11444,N_9252,N_9924);
nor U11445 (N_11445,N_8075,N_9213);
xnor U11446 (N_11446,N_8234,N_8579);
nor U11447 (N_11447,N_8434,N_8234);
nor U11448 (N_11448,N_8841,N_8479);
nor U11449 (N_11449,N_8488,N_9322);
nand U11450 (N_11450,N_8626,N_8322);
or U11451 (N_11451,N_8017,N_9787);
nor U11452 (N_11452,N_8315,N_9157);
xor U11453 (N_11453,N_9580,N_9688);
nor U11454 (N_11454,N_9267,N_8308);
nor U11455 (N_11455,N_8974,N_8491);
or U11456 (N_11456,N_8444,N_9614);
and U11457 (N_11457,N_9804,N_9294);
or U11458 (N_11458,N_9863,N_9939);
and U11459 (N_11459,N_9362,N_8973);
nor U11460 (N_11460,N_8805,N_9961);
and U11461 (N_11461,N_8021,N_9672);
nand U11462 (N_11462,N_8482,N_9766);
and U11463 (N_11463,N_9410,N_9850);
nand U11464 (N_11464,N_8387,N_8609);
nand U11465 (N_11465,N_8793,N_9981);
or U11466 (N_11466,N_9541,N_9780);
or U11467 (N_11467,N_8792,N_8863);
nor U11468 (N_11468,N_9988,N_9752);
nor U11469 (N_11469,N_9226,N_9353);
nand U11470 (N_11470,N_9912,N_9905);
nand U11471 (N_11471,N_9046,N_9537);
nand U11472 (N_11472,N_8216,N_9884);
nand U11473 (N_11473,N_8322,N_9582);
or U11474 (N_11474,N_9629,N_8476);
or U11475 (N_11475,N_8362,N_8123);
or U11476 (N_11476,N_8680,N_9125);
xnor U11477 (N_11477,N_8063,N_8453);
xnor U11478 (N_11478,N_8812,N_9563);
nand U11479 (N_11479,N_9848,N_8641);
and U11480 (N_11480,N_8451,N_8268);
nand U11481 (N_11481,N_8152,N_8817);
and U11482 (N_11482,N_8945,N_9908);
xnor U11483 (N_11483,N_8937,N_8244);
and U11484 (N_11484,N_9469,N_8395);
or U11485 (N_11485,N_9290,N_9905);
xor U11486 (N_11486,N_8406,N_9813);
and U11487 (N_11487,N_9875,N_9865);
and U11488 (N_11488,N_9912,N_8249);
nand U11489 (N_11489,N_8551,N_8544);
nand U11490 (N_11490,N_8729,N_9634);
or U11491 (N_11491,N_9368,N_8175);
and U11492 (N_11492,N_9955,N_8152);
nor U11493 (N_11493,N_9791,N_9230);
and U11494 (N_11494,N_8981,N_8736);
nand U11495 (N_11495,N_8596,N_8541);
nor U11496 (N_11496,N_9838,N_9589);
or U11497 (N_11497,N_8985,N_8271);
and U11498 (N_11498,N_8234,N_9953);
nor U11499 (N_11499,N_8072,N_9101);
xnor U11500 (N_11500,N_9906,N_9534);
and U11501 (N_11501,N_9242,N_8275);
nor U11502 (N_11502,N_8727,N_8911);
nand U11503 (N_11503,N_8280,N_8689);
and U11504 (N_11504,N_8235,N_9765);
or U11505 (N_11505,N_8300,N_8109);
and U11506 (N_11506,N_8706,N_9092);
or U11507 (N_11507,N_8092,N_9717);
nor U11508 (N_11508,N_8249,N_8926);
nand U11509 (N_11509,N_8943,N_9213);
or U11510 (N_11510,N_9898,N_9583);
nand U11511 (N_11511,N_8677,N_9408);
nor U11512 (N_11512,N_9571,N_9348);
nor U11513 (N_11513,N_9850,N_8135);
xnor U11514 (N_11514,N_8242,N_9008);
and U11515 (N_11515,N_9948,N_9791);
nor U11516 (N_11516,N_9184,N_8020);
nor U11517 (N_11517,N_9644,N_9798);
nor U11518 (N_11518,N_9593,N_8625);
xor U11519 (N_11519,N_8814,N_9638);
or U11520 (N_11520,N_8708,N_8509);
nor U11521 (N_11521,N_8113,N_9335);
or U11522 (N_11522,N_9017,N_9467);
or U11523 (N_11523,N_8749,N_9835);
or U11524 (N_11524,N_9539,N_9108);
nand U11525 (N_11525,N_9781,N_9420);
and U11526 (N_11526,N_9688,N_8539);
nand U11527 (N_11527,N_9650,N_9881);
nand U11528 (N_11528,N_9115,N_8629);
and U11529 (N_11529,N_8837,N_8645);
nand U11530 (N_11530,N_9860,N_8948);
or U11531 (N_11531,N_9650,N_9217);
and U11532 (N_11532,N_8318,N_8425);
xor U11533 (N_11533,N_9891,N_9819);
xor U11534 (N_11534,N_9154,N_8640);
nand U11535 (N_11535,N_9154,N_8132);
xor U11536 (N_11536,N_8815,N_8231);
xor U11537 (N_11537,N_8799,N_8823);
and U11538 (N_11538,N_8219,N_9769);
or U11539 (N_11539,N_9566,N_9285);
or U11540 (N_11540,N_9271,N_8657);
or U11541 (N_11541,N_9468,N_8624);
nor U11542 (N_11542,N_8716,N_9619);
nor U11543 (N_11543,N_8478,N_8608);
and U11544 (N_11544,N_8665,N_8577);
and U11545 (N_11545,N_9582,N_9822);
nor U11546 (N_11546,N_9488,N_8766);
nor U11547 (N_11547,N_8123,N_8782);
nor U11548 (N_11548,N_8402,N_9200);
and U11549 (N_11549,N_8843,N_8393);
nor U11550 (N_11550,N_9761,N_9750);
or U11551 (N_11551,N_9055,N_9625);
xnor U11552 (N_11552,N_9425,N_8365);
nand U11553 (N_11553,N_8240,N_8520);
nand U11554 (N_11554,N_8575,N_9517);
or U11555 (N_11555,N_8361,N_9465);
and U11556 (N_11556,N_9516,N_9276);
and U11557 (N_11557,N_9314,N_8217);
nor U11558 (N_11558,N_8997,N_9297);
xor U11559 (N_11559,N_8950,N_9925);
or U11560 (N_11560,N_8179,N_9532);
nand U11561 (N_11561,N_9489,N_9369);
nand U11562 (N_11562,N_9800,N_8797);
nand U11563 (N_11563,N_8151,N_9444);
xnor U11564 (N_11564,N_9970,N_9552);
and U11565 (N_11565,N_8394,N_9334);
xnor U11566 (N_11566,N_8132,N_8877);
nor U11567 (N_11567,N_8837,N_8877);
or U11568 (N_11568,N_8464,N_8626);
or U11569 (N_11569,N_8873,N_9537);
or U11570 (N_11570,N_9885,N_8048);
xor U11571 (N_11571,N_9366,N_8011);
or U11572 (N_11572,N_8678,N_9801);
nand U11573 (N_11573,N_8349,N_9482);
nor U11574 (N_11574,N_8382,N_8440);
nor U11575 (N_11575,N_8045,N_9246);
nand U11576 (N_11576,N_9020,N_9395);
nor U11577 (N_11577,N_8171,N_9980);
nand U11578 (N_11578,N_8773,N_8015);
or U11579 (N_11579,N_9362,N_8700);
nor U11580 (N_11580,N_8627,N_9036);
nor U11581 (N_11581,N_9452,N_9301);
nor U11582 (N_11582,N_8079,N_8808);
nand U11583 (N_11583,N_9877,N_9808);
nor U11584 (N_11584,N_9594,N_9094);
xor U11585 (N_11585,N_9132,N_8731);
and U11586 (N_11586,N_8017,N_8855);
nor U11587 (N_11587,N_9675,N_9964);
nor U11588 (N_11588,N_9565,N_8851);
and U11589 (N_11589,N_9262,N_9901);
or U11590 (N_11590,N_8011,N_8981);
nor U11591 (N_11591,N_8054,N_9563);
nand U11592 (N_11592,N_9126,N_9919);
nor U11593 (N_11593,N_8602,N_9579);
and U11594 (N_11594,N_9262,N_9916);
nor U11595 (N_11595,N_9328,N_8743);
and U11596 (N_11596,N_9313,N_9791);
nand U11597 (N_11597,N_8196,N_8950);
or U11598 (N_11598,N_8655,N_8270);
nor U11599 (N_11599,N_8508,N_9776);
or U11600 (N_11600,N_8087,N_9201);
xnor U11601 (N_11601,N_9018,N_9683);
nand U11602 (N_11602,N_9944,N_8991);
and U11603 (N_11603,N_9527,N_8866);
xor U11604 (N_11604,N_9215,N_8699);
and U11605 (N_11605,N_9246,N_8913);
or U11606 (N_11606,N_8570,N_8585);
nand U11607 (N_11607,N_9454,N_9669);
xor U11608 (N_11608,N_9260,N_8389);
or U11609 (N_11609,N_8522,N_8792);
and U11610 (N_11610,N_8702,N_9470);
nand U11611 (N_11611,N_9993,N_9675);
or U11612 (N_11612,N_8734,N_9605);
or U11613 (N_11613,N_9942,N_8497);
nand U11614 (N_11614,N_8401,N_9789);
nand U11615 (N_11615,N_9051,N_8552);
nand U11616 (N_11616,N_9081,N_9785);
nor U11617 (N_11617,N_9987,N_8071);
or U11618 (N_11618,N_8262,N_9949);
and U11619 (N_11619,N_9146,N_8725);
nand U11620 (N_11620,N_8462,N_8709);
nand U11621 (N_11621,N_8772,N_8489);
or U11622 (N_11622,N_9068,N_9662);
and U11623 (N_11623,N_8736,N_9863);
and U11624 (N_11624,N_8284,N_9578);
nand U11625 (N_11625,N_9155,N_8644);
or U11626 (N_11626,N_8285,N_9827);
or U11627 (N_11627,N_8860,N_9252);
nor U11628 (N_11628,N_9896,N_9547);
or U11629 (N_11629,N_8295,N_9901);
nor U11630 (N_11630,N_9733,N_8325);
nand U11631 (N_11631,N_8491,N_9581);
or U11632 (N_11632,N_8257,N_9815);
and U11633 (N_11633,N_8168,N_8639);
or U11634 (N_11634,N_9879,N_9552);
and U11635 (N_11635,N_8175,N_8675);
nor U11636 (N_11636,N_8242,N_9292);
nor U11637 (N_11637,N_9792,N_9764);
xnor U11638 (N_11638,N_8342,N_9903);
nor U11639 (N_11639,N_8146,N_9783);
xnor U11640 (N_11640,N_9625,N_9029);
and U11641 (N_11641,N_8259,N_8724);
and U11642 (N_11642,N_9112,N_9281);
or U11643 (N_11643,N_9655,N_8027);
nand U11644 (N_11644,N_8328,N_8627);
and U11645 (N_11645,N_9710,N_9089);
or U11646 (N_11646,N_9437,N_9372);
or U11647 (N_11647,N_8670,N_8529);
and U11648 (N_11648,N_8734,N_9581);
or U11649 (N_11649,N_8228,N_8729);
and U11650 (N_11650,N_8585,N_8966);
nand U11651 (N_11651,N_9592,N_9394);
nor U11652 (N_11652,N_9681,N_8576);
or U11653 (N_11653,N_8919,N_9090);
nor U11654 (N_11654,N_8856,N_9195);
or U11655 (N_11655,N_8408,N_8773);
or U11656 (N_11656,N_9314,N_8128);
nor U11657 (N_11657,N_8171,N_8934);
nor U11658 (N_11658,N_8109,N_8485);
or U11659 (N_11659,N_8005,N_9145);
or U11660 (N_11660,N_8405,N_9331);
and U11661 (N_11661,N_8031,N_9745);
nor U11662 (N_11662,N_9203,N_8358);
nand U11663 (N_11663,N_8530,N_9066);
and U11664 (N_11664,N_8940,N_9071);
nor U11665 (N_11665,N_9575,N_9065);
and U11666 (N_11666,N_9507,N_9471);
and U11667 (N_11667,N_8634,N_8235);
nand U11668 (N_11668,N_8952,N_8373);
nor U11669 (N_11669,N_8261,N_9319);
nand U11670 (N_11670,N_9638,N_8130);
nor U11671 (N_11671,N_8145,N_9533);
nand U11672 (N_11672,N_9647,N_9202);
nor U11673 (N_11673,N_9375,N_8253);
nor U11674 (N_11674,N_8681,N_8367);
and U11675 (N_11675,N_9094,N_9753);
and U11676 (N_11676,N_8068,N_9948);
or U11677 (N_11677,N_8833,N_9306);
or U11678 (N_11678,N_9093,N_8504);
or U11679 (N_11679,N_9952,N_9558);
or U11680 (N_11680,N_8139,N_9653);
xnor U11681 (N_11681,N_8966,N_9504);
or U11682 (N_11682,N_8798,N_9819);
nand U11683 (N_11683,N_8911,N_8323);
or U11684 (N_11684,N_9768,N_8180);
nor U11685 (N_11685,N_9249,N_8061);
xnor U11686 (N_11686,N_9301,N_9335);
xnor U11687 (N_11687,N_9604,N_9612);
and U11688 (N_11688,N_8942,N_9023);
or U11689 (N_11689,N_8834,N_9744);
and U11690 (N_11690,N_8508,N_9871);
xnor U11691 (N_11691,N_8574,N_9525);
nand U11692 (N_11692,N_8258,N_9725);
nand U11693 (N_11693,N_9387,N_8468);
and U11694 (N_11694,N_8176,N_8571);
xnor U11695 (N_11695,N_8619,N_8746);
or U11696 (N_11696,N_9729,N_9255);
nor U11697 (N_11697,N_9624,N_8072);
and U11698 (N_11698,N_8420,N_9148);
and U11699 (N_11699,N_9057,N_8151);
nand U11700 (N_11700,N_8370,N_9408);
and U11701 (N_11701,N_8053,N_8300);
and U11702 (N_11702,N_9075,N_8880);
nor U11703 (N_11703,N_9443,N_8882);
nor U11704 (N_11704,N_9325,N_9770);
nand U11705 (N_11705,N_8684,N_8353);
and U11706 (N_11706,N_9368,N_8310);
nor U11707 (N_11707,N_8006,N_9379);
and U11708 (N_11708,N_9816,N_9617);
nand U11709 (N_11709,N_9296,N_9756);
xnor U11710 (N_11710,N_9288,N_8603);
xor U11711 (N_11711,N_9995,N_9251);
nor U11712 (N_11712,N_9541,N_9789);
and U11713 (N_11713,N_8927,N_9569);
xnor U11714 (N_11714,N_8848,N_9321);
nor U11715 (N_11715,N_8496,N_9144);
and U11716 (N_11716,N_9458,N_9054);
nor U11717 (N_11717,N_8238,N_9041);
nand U11718 (N_11718,N_8151,N_9074);
and U11719 (N_11719,N_8036,N_8097);
nand U11720 (N_11720,N_8727,N_9741);
or U11721 (N_11721,N_9230,N_8495);
nor U11722 (N_11722,N_8815,N_8070);
and U11723 (N_11723,N_9839,N_9143);
nand U11724 (N_11724,N_8178,N_9542);
and U11725 (N_11725,N_9811,N_9861);
nand U11726 (N_11726,N_8947,N_8838);
or U11727 (N_11727,N_9233,N_9045);
or U11728 (N_11728,N_9353,N_8607);
and U11729 (N_11729,N_8843,N_9410);
xnor U11730 (N_11730,N_9770,N_9913);
and U11731 (N_11731,N_8455,N_8076);
or U11732 (N_11732,N_9464,N_8176);
xnor U11733 (N_11733,N_8139,N_8841);
nor U11734 (N_11734,N_8710,N_8640);
nor U11735 (N_11735,N_9098,N_8143);
nor U11736 (N_11736,N_8344,N_8032);
and U11737 (N_11737,N_8857,N_8993);
xnor U11738 (N_11738,N_8487,N_8795);
nand U11739 (N_11739,N_8649,N_8338);
and U11740 (N_11740,N_8802,N_8963);
nor U11741 (N_11741,N_9463,N_9041);
nor U11742 (N_11742,N_8275,N_8257);
and U11743 (N_11743,N_9275,N_9269);
nand U11744 (N_11744,N_8134,N_9351);
or U11745 (N_11745,N_9576,N_8667);
nor U11746 (N_11746,N_8465,N_9220);
and U11747 (N_11747,N_9584,N_8282);
nor U11748 (N_11748,N_9997,N_9130);
nand U11749 (N_11749,N_9825,N_9250);
xor U11750 (N_11750,N_9773,N_8053);
or U11751 (N_11751,N_9074,N_9536);
and U11752 (N_11752,N_9388,N_9962);
and U11753 (N_11753,N_8535,N_9864);
nand U11754 (N_11754,N_8533,N_9494);
and U11755 (N_11755,N_9827,N_8053);
xnor U11756 (N_11756,N_9836,N_9458);
xor U11757 (N_11757,N_8850,N_9360);
nand U11758 (N_11758,N_8268,N_9092);
nand U11759 (N_11759,N_9945,N_9309);
nand U11760 (N_11760,N_8173,N_8530);
xnor U11761 (N_11761,N_9748,N_9106);
or U11762 (N_11762,N_9265,N_9113);
nand U11763 (N_11763,N_9433,N_8670);
or U11764 (N_11764,N_9950,N_8141);
nand U11765 (N_11765,N_8920,N_8312);
or U11766 (N_11766,N_9582,N_9997);
nor U11767 (N_11767,N_8250,N_8110);
nor U11768 (N_11768,N_9676,N_8092);
nor U11769 (N_11769,N_8683,N_9292);
nor U11770 (N_11770,N_9714,N_9492);
and U11771 (N_11771,N_9461,N_9891);
nand U11772 (N_11772,N_9900,N_8120);
nand U11773 (N_11773,N_8524,N_9547);
or U11774 (N_11774,N_8794,N_9711);
and U11775 (N_11775,N_9650,N_8119);
nor U11776 (N_11776,N_8536,N_9015);
and U11777 (N_11777,N_9303,N_8222);
and U11778 (N_11778,N_8874,N_8356);
nor U11779 (N_11779,N_8184,N_8732);
nand U11780 (N_11780,N_8109,N_8292);
or U11781 (N_11781,N_9027,N_9014);
and U11782 (N_11782,N_9853,N_9753);
nor U11783 (N_11783,N_8046,N_8990);
nand U11784 (N_11784,N_9239,N_8270);
nand U11785 (N_11785,N_8109,N_8611);
nor U11786 (N_11786,N_9175,N_8369);
and U11787 (N_11787,N_9003,N_8319);
or U11788 (N_11788,N_9805,N_8220);
and U11789 (N_11789,N_8555,N_8766);
or U11790 (N_11790,N_9813,N_9057);
nor U11791 (N_11791,N_8690,N_8306);
nor U11792 (N_11792,N_9344,N_8605);
and U11793 (N_11793,N_8507,N_9559);
or U11794 (N_11794,N_8634,N_9669);
and U11795 (N_11795,N_8337,N_9801);
and U11796 (N_11796,N_9706,N_9837);
and U11797 (N_11797,N_9884,N_8839);
or U11798 (N_11798,N_8962,N_9093);
and U11799 (N_11799,N_8398,N_9741);
nand U11800 (N_11800,N_9740,N_9048);
or U11801 (N_11801,N_9441,N_9958);
and U11802 (N_11802,N_8570,N_8670);
and U11803 (N_11803,N_9096,N_8195);
and U11804 (N_11804,N_8214,N_9257);
nor U11805 (N_11805,N_8298,N_9139);
and U11806 (N_11806,N_9673,N_8768);
and U11807 (N_11807,N_9615,N_8783);
or U11808 (N_11808,N_8854,N_9075);
nand U11809 (N_11809,N_8823,N_8484);
or U11810 (N_11810,N_9469,N_8244);
xnor U11811 (N_11811,N_8007,N_9650);
nor U11812 (N_11812,N_8449,N_8513);
nand U11813 (N_11813,N_9761,N_9826);
nor U11814 (N_11814,N_8982,N_8163);
nor U11815 (N_11815,N_8985,N_8046);
nor U11816 (N_11816,N_8595,N_9338);
and U11817 (N_11817,N_9833,N_9563);
xor U11818 (N_11818,N_8139,N_9661);
or U11819 (N_11819,N_9127,N_8121);
or U11820 (N_11820,N_9512,N_9938);
nor U11821 (N_11821,N_8084,N_8170);
and U11822 (N_11822,N_8921,N_9292);
and U11823 (N_11823,N_9202,N_9982);
nor U11824 (N_11824,N_9561,N_9030);
and U11825 (N_11825,N_8157,N_8456);
or U11826 (N_11826,N_9366,N_9913);
nand U11827 (N_11827,N_8623,N_8273);
or U11828 (N_11828,N_9106,N_9025);
nor U11829 (N_11829,N_9889,N_9226);
nand U11830 (N_11830,N_9204,N_8114);
nor U11831 (N_11831,N_8469,N_8594);
xor U11832 (N_11832,N_9162,N_9181);
or U11833 (N_11833,N_9357,N_9146);
xor U11834 (N_11834,N_8968,N_8278);
nor U11835 (N_11835,N_9506,N_8374);
or U11836 (N_11836,N_8991,N_9360);
nor U11837 (N_11837,N_9356,N_8650);
or U11838 (N_11838,N_8446,N_9664);
and U11839 (N_11839,N_8280,N_8406);
nor U11840 (N_11840,N_9020,N_8247);
or U11841 (N_11841,N_8143,N_9850);
or U11842 (N_11842,N_9470,N_9150);
and U11843 (N_11843,N_8680,N_9867);
nor U11844 (N_11844,N_9673,N_9571);
nand U11845 (N_11845,N_8549,N_8026);
nor U11846 (N_11846,N_9168,N_9204);
nor U11847 (N_11847,N_9145,N_8423);
xnor U11848 (N_11848,N_9394,N_8465);
xnor U11849 (N_11849,N_9056,N_9100);
or U11850 (N_11850,N_8318,N_8186);
nand U11851 (N_11851,N_8379,N_9031);
or U11852 (N_11852,N_8628,N_8950);
or U11853 (N_11853,N_9970,N_8140);
and U11854 (N_11854,N_9516,N_9126);
xor U11855 (N_11855,N_8929,N_8931);
nor U11856 (N_11856,N_8874,N_8240);
xor U11857 (N_11857,N_8917,N_9267);
xnor U11858 (N_11858,N_8768,N_8296);
xor U11859 (N_11859,N_8202,N_9991);
nor U11860 (N_11860,N_8981,N_8645);
nor U11861 (N_11861,N_8269,N_8401);
nor U11862 (N_11862,N_9674,N_9144);
or U11863 (N_11863,N_9162,N_8593);
nand U11864 (N_11864,N_8615,N_9710);
nor U11865 (N_11865,N_9006,N_8539);
or U11866 (N_11866,N_8068,N_8538);
or U11867 (N_11867,N_9031,N_8753);
nand U11868 (N_11868,N_8593,N_9046);
and U11869 (N_11869,N_8989,N_9348);
nand U11870 (N_11870,N_8518,N_8827);
nor U11871 (N_11871,N_8251,N_9242);
or U11872 (N_11872,N_8014,N_8622);
nor U11873 (N_11873,N_8456,N_8010);
or U11874 (N_11874,N_8293,N_9822);
nor U11875 (N_11875,N_8334,N_8836);
nor U11876 (N_11876,N_9344,N_9299);
nand U11877 (N_11877,N_8772,N_8761);
nor U11878 (N_11878,N_9435,N_9521);
nor U11879 (N_11879,N_9463,N_8967);
nor U11880 (N_11880,N_9624,N_9148);
nor U11881 (N_11881,N_8011,N_8701);
or U11882 (N_11882,N_8762,N_8838);
nor U11883 (N_11883,N_9757,N_8424);
or U11884 (N_11884,N_8287,N_9906);
nor U11885 (N_11885,N_9197,N_9132);
nand U11886 (N_11886,N_8415,N_8020);
nor U11887 (N_11887,N_9887,N_9218);
xnor U11888 (N_11888,N_9632,N_8316);
nand U11889 (N_11889,N_8791,N_9817);
nor U11890 (N_11890,N_8402,N_9691);
or U11891 (N_11891,N_9521,N_8263);
xnor U11892 (N_11892,N_9154,N_8179);
nor U11893 (N_11893,N_8411,N_8010);
xor U11894 (N_11894,N_9691,N_8299);
nand U11895 (N_11895,N_8106,N_9951);
or U11896 (N_11896,N_9648,N_9855);
and U11897 (N_11897,N_8140,N_9489);
nand U11898 (N_11898,N_8966,N_8670);
and U11899 (N_11899,N_9062,N_8512);
or U11900 (N_11900,N_8029,N_8075);
or U11901 (N_11901,N_8270,N_8076);
nor U11902 (N_11902,N_8304,N_8709);
nand U11903 (N_11903,N_8869,N_8362);
nor U11904 (N_11904,N_8610,N_9206);
and U11905 (N_11905,N_8861,N_9650);
or U11906 (N_11906,N_8398,N_8378);
or U11907 (N_11907,N_8506,N_8443);
or U11908 (N_11908,N_9756,N_9281);
nand U11909 (N_11909,N_8349,N_9448);
nand U11910 (N_11910,N_9055,N_8999);
or U11911 (N_11911,N_9446,N_8212);
or U11912 (N_11912,N_9842,N_8095);
nor U11913 (N_11913,N_9895,N_8112);
or U11914 (N_11914,N_8573,N_9246);
nor U11915 (N_11915,N_9861,N_8778);
or U11916 (N_11916,N_9226,N_8406);
nand U11917 (N_11917,N_9864,N_8027);
xor U11918 (N_11918,N_9517,N_9792);
nand U11919 (N_11919,N_8379,N_9840);
nand U11920 (N_11920,N_8879,N_9999);
or U11921 (N_11921,N_8065,N_9089);
and U11922 (N_11922,N_9994,N_9246);
or U11923 (N_11923,N_8573,N_9328);
nor U11924 (N_11924,N_9753,N_9929);
and U11925 (N_11925,N_9529,N_8613);
or U11926 (N_11926,N_8191,N_9849);
and U11927 (N_11927,N_8495,N_9374);
or U11928 (N_11928,N_9746,N_8085);
and U11929 (N_11929,N_8073,N_9479);
and U11930 (N_11930,N_9075,N_8051);
or U11931 (N_11931,N_8799,N_9715);
or U11932 (N_11932,N_9216,N_8232);
nor U11933 (N_11933,N_9579,N_9253);
or U11934 (N_11934,N_9940,N_9915);
and U11935 (N_11935,N_9883,N_9017);
and U11936 (N_11936,N_9810,N_8267);
xor U11937 (N_11937,N_8932,N_9816);
nand U11938 (N_11938,N_9646,N_9366);
nor U11939 (N_11939,N_8616,N_9167);
nor U11940 (N_11940,N_8836,N_9038);
nor U11941 (N_11941,N_8870,N_8413);
or U11942 (N_11942,N_8806,N_8735);
xor U11943 (N_11943,N_9846,N_8986);
nand U11944 (N_11944,N_8451,N_8751);
and U11945 (N_11945,N_9955,N_9530);
nor U11946 (N_11946,N_9907,N_8540);
nor U11947 (N_11947,N_8678,N_9753);
or U11948 (N_11948,N_8794,N_9262);
nor U11949 (N_11949,N_8318,N_8505);
nand U11950 (N_11950,N_9005,N_9768);
nor U11951 (N_11951,N_9092,N_9837);
and U11952 (N_11952,N_9918,N_9228);
nand U11953 (N_11953,N_8831,N_9788);
or U11954 (N_11954,N_8919,N_9998);
nor U11955 (N_11955,N_9423,N_8789);
nand U11956 (N_11956,N_8454,N_8762);
nand U11957 (N_11957,N_8345,N_8580);
nor U11958 (N_11958,N_8797,N_9089);
nand U11959 (N_11959,N_8883,N_9544);
nor U11960 (N_11960,N_9127,N_9509);
or U11961 (N_11961,N_8479,N_8471);
or U11962 (N_11962,N_8690,N_8709);
and U11963 (N_11963,N_8808,N_8881);
and U11964 (N_11964,N_8904,N_8450);
and U11965 (N_11965,N_8267,N_9132);
nand U11966 (N_11966,N_9298,N_9329);
nor U11967 (N_11967,N_9343,N_9055);
or U11968 (N_11968,N_9459,N_8829);
and U11969 (N_11969,N_9166,N_9242);
or U11970 (N_11970,N_9803,N_9088);
nor U11971 (N_11971,N_9041,N_9195);
nand U11972 (N_11972,N_8785,N_8057);
and U11973 (N_11973,N_9134,N_8476);
nor U11974 (N_11974,N_9095,N_8427);
nor U11975 (N_11975,N_9314,N_9147);
nand U11976 (N_11976,N_9614,N_9619);
or U11977 (N_11977,N_8636,N_8433);
nor U11978 (N_11978,N_9959,N_8566);
nand U11979 (N_11979,N_8573,N_9145);
nor U11980 (N_11980,N_8147,N_8589);
and U11981 (N_11981,N_8987,N_9295);
or U11982 (N_11982,N_8964,N_9346);
and U11983 (N_11983,N_8782,N_9944);
or U11984 (N_11984,N_9283,N_9846);
nor U11985 (N_11985,N_8217,N_8721);
or U11986 (N_11986,N_8883,N_8519);
nor U11987 (N_11987,N_8238,N_8279);
nand U11988 (N_11988,N_9849,N_9480);
and U11989 (N_11989,N_9357,N_8799);
and U11990 (N_11990,N_9484,N_8906);
xor U11991 (N_11991,N_8665,N_8572);
xor U11992 (N_11992,N_9134,N_8524);
and U11993 (N_11993,N_8747,N_9981);
and U11994 (N_11994,N_8263,N_9781);
nand U11995 (N_11995,N_8388,N_9319);
or U11996 (N_11996,N_8666,N_9567);
xnor U11997 (N_11997,N_8634,N_9604);
and U11998 (N_11998,N_9273,N_8346);
or U11999 (N_11999,N_8531,N_9080);
nor U12000 (N_12000,N_11399,N_10989);
and U12001 (N_12001,N_10067,N_10970);
and U12002 (N_12002,N_10541,N_11895);
nor U12003 (N_12003,N_11742,N_11928);
nand U12004 (N_12004,N_11770,N_10048);
or U12005 (N_12005,N_10618,N_11595);
or U12006 (N_12006,N_11534,N_11792);
nand U12007 (N_12007,N_10775,N_11855);
nor U12008 (N_12008,N_11275,N_10333);
and U12009 (N_12009,N_11035,N_11495);
nor U12010 (N_12010,N_10241,N_10218);
nand U12011 (N_12011,N_10927,N_10044);
or U12012 (N_12012,N_11507,N_10813);
xor U12013 (N_12013,N_11550,N_11262);
or U12014 (N_12014,N_10306,N_10599);
or U12015 (N_12015,N_11930,N_11631);
nor U12016 (N_12016,N_10356,N_10191);
and U12017 (N_12017,N_10072,N_11911);
or U12018 (N_12018,N_11562,N_10730);
or U12019 (N_12019,N_11775,N_10979);
xnor U12020 (N_12020,N_10961,N_11776);
and U12021 (N_12021,N_10697,N_10152);
xnor U12022 (N_12022,N_11238,N_10947);
nor U12023 (N_12023,N_10509,N_10153);
or U12024 (N_12024,N_11006,N_11863);
or U12025 (N_12025,N_11810,N_10199);
or U12026 (N_12026,N_11762,N_10227);
nand U12027 (N_12027,N_10861,N_11292);
nor U12028 (N_12028,N_10539,N_11492);
xor U12029 (N_12029,N_11548,N_10843);
nand U12030 (N_12030,N_10787,N_10830);
or U12031 (N_12031,N_10980,N_11710);
or U12032 (N_12032,N_10906,N_10936);
nand U12033 (N_12033,N_10563,N_11878);
xor U12034 (N_12034,N_11535,N_11365);
xor U12035 (N_12035,N_11152,N_10010);
nand U12036 (N_12036,N_11433,N_11981);
and U12037 (N_12037,N_10086,N_10404);
and U12038 (N_12038,N_11840,N_11621);
nor U12039 (N_12039,N_11763,N_10497);
nand U12040 (N_12040,N_10885,N_10726);
or U12041 (N_12041,N_11627,N_11479);
and U12042 (N_12042,N_10869,N_11857);
nand U12043 (N_12043,N_10000,N_11943);
and U12044 (N_12044,N_11564,N_11191);
nor U12045 (N_12045,N_11439,N_11545);
or U12046 (N_12046,N_10949,N_11740);
nor U12047 (N_12047,N_10374,N_11558);
nand U12048 (N_12048,N_11676,N_11636);
or U12049 (N_12049,N_10874,N_11226);
nand U12050 (N_12050,N_10265,N_11644);
and U12051 (N_12051,N_11526,N_11777);
and U12052 (N_12052,N_10997,N_10889);
xor U12053 (N_12053,N_11120,N_10682);
or U12054 (N_12054,N_11056,N_10308);
and U12055 (N_12055,N_11251,N_11092);
nor U12056 (N_12056,N_11711,N_10104);
and U12057 (N_12057,N_10822,N_10430);
nor U12058 (N_12058,N_10942,N_10130);
or U12059 (N_12059,N_11303,N_10346);
and U12060 (N_12060,N_10420,N_11835);
nand U12061 (N_12061,N_10077,N_11187);
nand U12062 (N_12062,N_10425,N_11037);
nand U12063 (N_12063,N_11925,N_11483);
nand U12064 (N_12064,N_10683,N_10564);
nand U12065 (N_12065,N_11880,N_11582);
and U12066 (N_12066,N_10619,N_11811);
nand U12067 (N_12067,N_10606,N_11693);
nor U12068 (N_12068,N_11194,N_10432);
nor U12069 (N_12069,N_10477,N_11899);
nand U12070 (N_12070,N_11195,N_11622);
nand U12071 (N_12071,N_10230,N_10485);
xor U12072 (N_12072,N_10659,N_11235);
and U12073 (N_12073,N_11877,N_10231);
xnor U12074 (N_12074,N_11699,N_11616);
or U12075 (N_12075,N_10609,N_11632);
or U12076 (N_12076,N_10800,N_10455);
nor U12077 (N_12077,N_11975,N_11889);
xor U12078 (N_12078,N_10418,N_11720);
and U12079 (N_12079,N_11718,N_11691);
nor U12080 (N_12080,N_10168,N_10002);
xor U12081 (N_12081,N_11020,N_10003);
nand U12082 (N_12082,N_11665,N_10288);
xor U12083 (N_12083,N_11746,N_10845);
nor U12084 (N_12084,N_11153,N_11480);
nand U12085 (N_12085,N_10728,N_11013);
or U12086 (N_12086,N_11842,N_11858);
nand U12087 (N_12087,N_11108,N_11279);
or U12088 (N_12088,N_10854,N_10272);
nand U12089 (N_12089,N_11966,N_11253);
nand U12090 (N_12090,N_10508,N_10850);
nor U12091 (N_12091,N_10504,N_10267);
or U12092 (N_12092,N_11247,N_11730);
and U12093 (N_12093,N_11313,N_11050);
nand U12094 (N_12094,N_10318,N_10832);
and U12095 (N_12095,N_11908,N_11786);
or U12096 (N_12096,N_11384,N_11087);
xor U12097 (N_12097,N_11172,N_10208);
or U12098 (N_12098,N_11931,N_10116);
nor U12099 (N_12099,N_11128,N_11230);
nor U12100 (N_12100,N_10219,N_11655);
nand U12101 (N_12101,N_11814,N_10762);
xor U12102 (N_12102,N_10157,N_11276);
nor U12103 (N_12103,N_10801,N_10027);
nand U12104 (N_12104,N_10484,N_11596);
or U12105 (N_12105,N_10918,N_10555);
or U12106 (N_12106,N_11530,N_10164);
and U12107 (N_12107,N_10159,N_11354);
xor U12108 (N_12108,N_10953,N_11156);
nand U12109 (N_12109,N_11511,N_11204);
nor U12110 (N_12110,N_10446,N_11097);
nor U12111 (N_12111,N_11683,N_11151);
nor U12112 (N_12112,N_10828,N_11881);
or U12113 (N_12113,N_10693,N_10444);
or U12114 (N_12114,N_11989,N_11353);
nand U12115 (N_12115,N_10323,N_10932);
and U12116 (N_12116,N_10115,N_11910);
nor U12117 (N_12117,N_11465,N_11256);
nand U12118 (N_12118,N_11452,N_11377);
and U12119 (N_12119,N_11958,N_10627);
nor U12120 (N_12120,N_11382,N_11255);
and U12121 (N_12121,N_10424,N_11038);
or U12122 (N_12122,N_11510,N_11263);
xnor U12123 (N_12123,N_11994,N_11915);
nor U12124 (N_12124,N_11397,N_10975);
nor U12125 (N_12125,N_10126,N_10771);
or U12126 (N_12126,N_11117,N_11779);
nand U12127 (N_12127,N_10470,N_11192);
xnor U12128 (N_12128,N_11995,N_10460);
or U12129 (N_12129,N_10160,N_11688);
or U12130 (N_12130,N_10778,N_11054);
nor U12131 (N_12131,N_10400,N_10808);
or U12132 (N_12132,N_10973,N_10417);
or U12133 (N_12133,N_10088,N_10169);
and U12134 (N_12134,N_10053,N_11298);
and U12135 (N_12135,N_10641,N_11268);
nor U12136 (N_12136,N_11017,N_10668);
or U12137 (N_12137,N_10137,N_11307);
xnor U12138 (N_12138,N_10279,N_10748);
xor U12139 (N_12139,N_11150,N_11280);
and U12140 (N_12140,N_11458,N_10638);
or U12141 (N_12141,N_11434,N_11010);
nor U12142 (N_12142,N_10349,N_11062);
nand U12143 (N_12143,N_11233,N_11415);
nand U12144 (N_12144,N_10055,N_11392);
nand U12145 (N_12145,N_10211,N_10473);
nand U12146 (N_12146,N_11012,N_10271);
nor U12147 (N_12147,N_11248,N_10329);
and U12148 (N_12148,N_11768,N_11674);
and U12149 (N_12149,N_10026,N_11780);
or U12150 (N_12150,N_10803,N_10548);
or U12151 (N_12151,N_11847,N_10805);
nand U12152 (N_12152,N_10838,N_10297);
and U12153 (N_12153,N_10738,N_11435);
nand U12154 (N_12154,N_11907,N_10715);
and U12155 (N_12155,N_11305,N_10457);
and U12156 (N_12156,N_11127,N_10671);
or U12157 (N_12157,N_10569,N_11119);
nor U12158 (N_12158,N_11372,N_10145);
or U12159 (N_12159,N_11823,N_10395);
nand U12160 (N_12160,N_10955,N_10507);
nand U12161 (N_12161,N_10930,N_11628);
or U12162 (N_12162,N_10605,N_10025);
nand U12163 (N_12163,N_11756,N_10733);
nand U12164 (N_12164,N_10920,N_11278);
or U12165 (N_12165,N_11019,N_10516);
nor U12166 (N_12166,N_11283,N_11084);
nor U12167 (N_12167,N_11257,N_11888);
xnor U12168 (N_12168,N_10052,N_11497);
nor U12169 (N_12169,N_10431,N_10965);
nor U12170 (N_12170,N_11824,N_11684);
or U12171 (N_12171,N_11031,N_10766);
and U12172 (N_12172,N_10774,N_11042);
and U12173 (N_12173,N_10956,N_11294);
and U12174 (N_12174,N_11373,N_10750);
and U12175 (N_12175,N_10795,N_10944);
nor U12176 (N_12176,N_11991,N_11281);
nand U12177 (N_12177,N_10383,N_11585);
or U12178 (N_12178,N_11099,N_10372);
nand U12179 (N_12179,N_10855,N_11623);
nor U12180 (N_12180,N_10651,N_10253);
nor U12181 (N_12181,N_11242,N_10596);
and U12182 (N_12182,N_11098,N_10338);
xor U12183 (N_12183,N_11629,N_10487);
nand U12184 (N_12184,N_11892,N_10342);
or U12185 (N_12185,N_11520,N_10799);
nand U12186 (N_12186,N_10684,N_10633);
nor U12187 (N_12187,N_11809,N_10001);
nor U12188 (N_12188,N_10071,N_10405);
xnor U12189 (N_12189,N_10696,N_11906);
nand U12190 (N_12190,N_11778,N_10657);
xnor U12191 (N_12191,N_10134,N_10817);
and U12192 (N_12192,N_11515,N_10574);
and U12193 (N_12193,N_11410,N_10197);
or U12194 (N_12194,N_10046,N_11182);
nor U12195 (N_12195,N_11443,N_10571);
or U12196 (N_12196,N_10464,N_10558);
nand U12197 (N_12197,N_10796,N_10471);
or U12198 (N_12198,N_10644,N_11446);
or U12199 (N_12199,N_10380,N_10459);
nor U12200 (N_12200,N_10670,N_10216);
or U12201 (N_12201,N_10552,N_10061);
and U12202 (N_12202,N_11387,N_10519);
and U12203 (N_12203,N_10503,N_10406);
or U12204 (N_12204,N_10587,N_10736);
xnor U12205 (N_12205,N_10623,N_11649);
xnor U12206 (N_12206,N_10802,N_10339);
nand U12207 (N_12207,N_10158,N_10196);
nor U12208 (N_12208,N_11047,N_10794);
nand U12209 (N_12209,N_10387,N_10835);
nand U12210 (N_12210,N_11220,N_10829);
nand U12211 (N_12211,N_10707,N_10362);
nor U12212 (N_12212,N_11146,N_10540);
nor U12213 (N_12213,N_11648,N_11170);
nand U12214 (N_12214,N_11210,N_11867);
and U12215 (N_12215,N_10864,N_11751);
and U12216 (N_12216,N_10994,N_11553);
and U12217 (N_12217,N_10190,N_11816);
and U12218 (N_12218,N_10751,N_10322);
or U12219 (N_12219,N_10089,N_10546);
nand U12220 (N_12220,N_10041,N_11987);
nand U12221 (N_12221,N_11979,N_10185);
or U12222 (N_12222,N_10462,N_10188);
and U12223 (N_12223,N_11694,N_10140);
xor U12224 (N_12224,N_10579,N_11732);
or U12225 (N_12225,N_10852,N_11815);
and U12226 (N_12226,N_11234,N_11190);
nor U12227 (N_12227,N_11971,N_11716);
nand U12228 (N_12228,N_10493,N_11396);
nand U12229 (N_12229,N_11274,N_11707);
or U12230 (N_12230,N_11296,N_10319);
nand U12231 (N_12231,N_10213,N_11455);
or U12232 (N_12232,N_11659,N_11726);
nand U12233 (N_12233,N_10836,N_10447);
and U12234 (N_12234,N_11083,N_11096);
or U12235 (N_12235,N_11747,N_10268);
nand U12236 (N_12236,N_10103,N_11882);
nor U12237 (N_12237,N_10538,N_11838);
and U12238 (N_12238,N_11996,N_11125);
xor U12239 (N_12239,N_10679,N_10243);
nor U12240 (N_12240,N_10959,N_11287);
and U12241 (N_12241,N_10228,N_11528);
nor U12242 (N_12242,N_10857,N_11390);
and U12243 (N_12243,N_11134,N_11609);
and U12244 (N_12244,N_10068,N_10391);
and U12245 (N_12245,N_11884,N_10646);
nand U12246 (N_12246,N_10175,N_11865);
nor U12247 (N_12247,N_10883,N_10968);
and U12248 (N_12248,N_11025,N_10653);
nor U12249 (N_12249,N_11115,N_10441);
nand U12250 (N_12250,N_10226,N_10414);
and U12251 (N_12251,N_10871,N_11918);
and U12252 (N_12252,N_11482,N_10712);
or U12253 (N_12253,N_11589,N_11791);
nor U12254 (N_12254,N_10719,N_10704);
nand U12255 (N_12255,N_11034,N_11527);
and U12256 (N_12256,N_10345,N_11348);
nor U12257 (N_12257,N_11949,N_11522);
xor U12258 (N_12258,N_10809,N_11171);
nand U12259 (N_12259,N_10776,N_10217);
nand U12260 (N_12260,N_11757,N_10937);
xnor U12261 (N_12261,N_11267,N_11846);
nor U12262 (N_12262,N_11708,N_10142);
nor U12263 (N_12263,N_11309,N_10512);
xnor U12264 (N_12264,N_11505,N_11744);
and U12265 (N_12265,N_10903,N_10298);
nand U12266 (N_12266,N_10992,N_11324);
xnor U12267 (N_12267,N_11990,N_10028);
or U12268 (N_12268,N_10030,N_10422);
nand U12269 (N_12269,N_10790,N_11544);
nand U12270 (N_12270,N_11625,N_11848);
or U12271 (N_12271,N_11978,N_11932);
nand U12272 (N_12272,N_11602,N_11784);
nor U12273 (N_12273,N_11972,N_11613);
and U12274 (N_12274,N_11346,N_11349);
and U12275 (N_12275,N_11845,N_10669);
nand U12276 (N_12276,N_10798,N_10632);
xor U12277 (N_12277,N_11921,N_11678);
and U12278 (N_12278,N_11894,N_11651);
nor U12279 (N_12279,N_11597,N_10629);
and U12280 (N_12280,N_11069,N_11124);
or U12281 (N_12281,N_11243,N_10007);
nor U12282 (N_12282,N_11774,N_10437);
nor U12283 (N_12283,N_11870,N_11362);
nor U12284 (N_12284,N_11417,N_10634);
or U12285 (N_12285,N_10106,N_11273);
or U12286 (N_12286,N_10963,N_11359);
nor U12287 (N_12287,N_11566,N_10337);
or U12288 (N_12288,N_10610,N_11706);
nand U12289 (N_12289,N_11232,N_10962);
or U12290 (N_12290,N_11430,N_10643);
or U12291 (N_12291,N_11481,N_11183);
or U12292 (N_12292,N_10550,N_10222);
or U12293 (N_12293,N_10532,N_10084);
and U12294 (N_12294,N_11539,N_11939);
or U12295 (N_12295,N_10178,N_10282);
or U12296 (N_12296,N_11041,N_11941);
or U12297 (N_12297,N_10179,N_10823);
nand U12298 (N_12298,N_10156,N_10662);
nand U12299 (N_12299,N_10545,N_10148);
xnor U12300 (N_12300,N_11942,N_10124);
nor U12301 (N_12301,N_11113,N_11366);
or U12302 (N_12302,N_10045,N_10583);
and U12303 (N_12303,N_10018,N_10549);
and U12304 (N_12304,N_11647,N_10872);
nor U12305 (N_12305,N_10902,N_11022);
nand U12306 (N_12306,N_10011,N_11656);
or U12307 (N_12307,N_10394,N_10515);
or U12308 (N_12308,N_10248,N_11252);
and U12309 (N_12309,N_10370,N_10990);
nor U12310 (N_12310,N_11612,N_10878);
nand U12311 (N_12311,N_10209,N_11619);
xnor U12312 (N_12312,N_10529,N_10278);
or U12313 (N_12313,N_11618,N_10703);
and U12314 (N_12314,N_10720,N_11004);
nand U12315 (N_12315,N_10097,N_11681);
or U12316 (N_12316,N_11211,N_11560);
and U12317 (N_12317,N_11834,N_11578);
xnor U12318 (N_12318,N_11781,N_10811);
and U12319 (N_12319,N_10429,N_11736);
nor U12320 (N_12320,N_11961,N_10511);
nand U12321 (N_12321,N_10492,N_10525);
nand U12322 (N_12322,N_11168,N_11935);
and U12323 (N_12323,N_10702,N_10004);
nor U12324 (N_12324,N_10969,N_11212);
nor U12325 (N_12325,N_10143,N_11999);
or U12326 (N_12326,N_10685,N_11322);
nor U12327 (N_12327,N_10737,N_11166);
and U12328 (N_12328,N_11159,N_11854);
or U12329 (N_12329,N_10138,N_10582);
nor U12330 (N_12330,N_10531,N_10238);
or U12331 (N_12331,N_10352,N_11040);
nor U12332 (N_12332,N_11849,N_11327);
nor U12333 (N_12333,N_11643,N_11690);
nand U12334 (N_12334,N_10310,N_10626);
nor U12335 (N_12335,N_11873,N_11551);
and U12336 (N_12336,N_11788,N_10163);
nand U12337 (N_12337,N_11715,N_10500);
and U12338 (N_12338,N_10987,N_10264);
nor U12339 (N_12339,N_10354,N_10938);
and U12340 (N_12340,N_10166,N_10656);
nand U12341 (N_12341,N_10654,N_10616);
and U12342 (N_12342,N_10882,N_10093);
or U12343 (N_12343,N_11702,N_11689);
or U12344 (N_12344,N_11580,N_11464);
nand U12345 (N_12345,N_10220,N_11594);
or U12346 (N_12346,N_10758,N_11502);
and U12347 (N_12347,N_10933,N_11135);
nand U12348 (N_12348,N_11357,N_10954);
or U12349 (N_12349,N_11800,N_11375);
or U12350 (N_12350,N_11229,N_11451);
nor U12351 (N_12351,N_10313,N_10999);
nand U12352 (N_12352,N_11328,N_11293);
or U12353 (N_12353,N_10221,N_11998);
and U12354 (N_12354,N_10674,N_11103);
nor U12355 (N_12355,N_10409,N_11790);
nor U12356 (N_12356,N_11896,N_11940);
or U12357 (N_12357,N_10886,N_11335);
or U12358 (N_12358,N_10875,N_11922);
or U12359 (N_12359,N_11462,N_11959);
nor U12360 (N_12360,N_10788,N_11246);
and U12361 (N_12361,N_11330,N_10355);
nand U12362 (N_12362,N_10330,N_10357);
nand U12363 (N_12363,N_10824,N_11734);
nor U12364 (N_12364,N_11927,N_10649);
or U12365 (N_12365,N_11723,N_11200);
nor U12366 (N_12366,N_10266,N_10578);
or U12367 (N_12367,N_10698,N_10401);
or U12368 (N_12368,N_11670,N_10478);
or U12369 (N_12369,N_11533,N_10642);
or U12370 (N_12370,N_11011,N_11389);
or U12371 (N_12371,N_11523,N_10063);
and U12372 (N_12372,N_10486,N_10365);
nor U12373 (N_12373,N_11116,N_11599);
nor U12374 (N_12374,N_11667,N_11432);
or U12375 (N_12375,N_11828,N_10204);
nand U12376 (N_12376,N_10128,N_10381);
or U12377 (N_12377,N_11486,N_10263);
or U12378 (N_12378,N_10551,N_11080);
xor U12379 (N_12379,N_11965,N_11109);
or U12380 (N_12380,N_11409,N_11713);
and U12381 (N_12381,N_10735,N_11604);
nand U12382 (N_12382,N_11671,N_11340);
and U12383 (N_12383,N_11291,N_11750);
or U12384 (N_12384,N_11974,N_11078);
or U12385 (N_12385,N_10423,N_10588);
and U12386 (N_12386,N_10699,N_11009);
and U12387 (N_12387,N_11143,N_11323);
nor U12388 (N_12388,N_10786,N_10518);
or U12389 (N_12389,N_11695,N_10522);
or U12390 (N_12390,N_11532,N_11570);
nand U12391 (N_12391,N_10328,N_11219);
nor U12392 (N_12392,N_10326,N_11095);
nor U12393 (N_12393,N_11350,N_11576);
nor U12394 (N_12394,N_10170,N_10589);
and U12395 (N_12395,N_10347,N_11188);
nor U12396 (N_12396,N_10755,N_10759);
and U12397 (N_12397,N_10307,N_11361);
xnor U12398 (N_12398,N_11426,N_10099);
nor U12399 (N_12399,N_11333,N_10373);
nor U12400 (N_12400,N_11852,N_11831);
and U12401 (N_12401,N_11240,N_11712);
nand U12402 (N_12402,N_11586,N_10520);
nor U12403 (N_12403,N_10490,N_11381);
nand U12404 (N_12404,N_11002,N_10946);
and U12405 (N_12405,N_11442,N_10210);
nor U12406 (N_12406,N_11652,N_11202);
and U12407 (N_12407,N_11295,N_11901);
xnor U12408 (N_12408,N_10785,N_10960);
xor U12409 (N_12409,N_11174,N_11717);
nor U12410 (N_12410,N_10392,N_11048);
nor U12411 (N_12411,N_11310,N_11075);
nor U12412 (N_12412,N_10594,N_10098);
and U12413 (N_12413,N_10524,N_10309);
or U12414 (N_12414,N_11951,N_10284);
nand U12415 (N_12415,N_10998,N_10521);
and U12416 (N_12416,N_10314,N_10144);
nor U12417 (N_12417,N_10840,N_11765);
xor U12418 (N_12418,N_11091,N_11752);
xnor U12419 (N_12419,N_11249,N_11351);
nand U12420 (N_12420,N_11661,N_10453);
and U12421 (N_12421,N_10768,N_10122);
nor U12422 (N_12422,N_11224,N_10568);
nor U12423 (N_12423,N_11850,N_11236);
nor U12424 (N_12424,N_10689,N_10252);
or U12425 (N_12425,N_11569,N_11261);
nand U12426 (N_12426,N_11259,N_10870);
and U12427 (N_12427,N_11077,N_10761);
nand U12428 (N_12428,N_10734,N_10691);
nand U12429 (N_12429,N_10593,N_11821);
and U12430 (N_12430,N_10976,N_11079);
and U12431 (N_12431,N_11739,N_10259);
or U12432 (N_12432,N_11587,N_11565);
nand U12433 (N_12433,N_10783,N_11076);
nor U12434 (N_12434,N_10119,N_11748);
and U12435 (N_12435,N_10488,N_11697);
nor U12436 (N_12436,N_11731,N_10951);
and U12437 (N_12437,N_10247,N_11856);
or U12438 (N_12438,N_11937,N_10176);
nor U12439 (N_12439,N_10376,N_11057);
and U12440 (N_12440,N_10701,N_10971);
and U12441 (N_12441,N_11735,N_10398);
nor U12442 (N_12442,N_10631,N_10615);
or U12443 (N_12443,N_11605,N_11008);
nand U12444 (N_12444,N_10335,N_11501);
nor U12445 (N_12445,N_10331,N_10841);
xor U12446 (N_12446,N_11891,N_10502);
nor U12447 (N_12447,N_10483,N_10233);
and U12448 (N_12448,N_11369,N_10544);
or U12449 (N_12449,N_11488,N_11902);
nor U12450 (N_12450,N_11271,N_11461);
and U12451 (N_12451,N_11724,N_10913);
or U12452 (N_12452,N_10262,N_10673);
or U12453 (N_12453,N_10863,N_11064);
nor U12454 (N_12454,N_11641,N_10107);
and U12455 (N_12455,N_10753,N_11663);
nor U12456 (N_12456,N_10127,N_11547);
nand U12457 (N_12457,N_10369,N_11646);
xnor U12458 (N_12458,N_10022,N_11798);
nor U12459 (N_12459,N_10993,N_11913);
and U12460 (N_12460,N_11339,N_11832);
nand U12461 (N_12461,N_10250,N_10637);
and U12462 (N_12462,N_11014,N_11427);
nor U12463 (N_12463,N_10640,N_10079);
and U12464 (N_12464,N_11423,N_11318);
and U12465 (N_12465,N_10203,N_10948);
nand U12466 (N_12466,N_11217,N_10706);
nor U12467 (N_12467,N_11315,N_11887);
nand U12468 (N_12468,N_10407,N_11967);
and U12469 (N_12469,N_11568,N_10815);
nand U12470 (N_12470,N_10060,N_10677);
nor U12471 (N_12471,N_11221,N_10914);
nand U12472 (N_12472,N_10700,N_10344);
or U12473 (N_12473,N_11139,N_10672);
or U12474 (N_12474,N_11537,N_10315);
nor U12475 (N_12475,N_10350,N_11438);
nor U12476 (N_12476,N_10240,N_11543);
and U12477 (N_12477,N_11700,N_10110);
and U12478 (N_12478,N_11938,N_11177);
or U12479 (N_12479,N_10324,N_11411);
nand U12480 (N_12480,N_10879,N_11371);
or U12481 (N_12481,N_10862,N_10109);
nand U12482 (N_12482,N_11015,N_11573);
or U12483 (N_12483,N_10514,N_11874);
or U12484 (N_12484,N_11929,N_10566);
nand U12485 (N_12485,N_11866,N_11196);
and U12486 (N_12486,N_10584,N_11270);
nor U12487 (N_12487,N_10403,N_11806);
and U12488 (N_12488,N_11680,N_10040);
nand U12489 (N_12489,N_11819,N_11985);
and U12490 (N_12490,N_11241,N_11403);
or U12491 (N_12491,N_11957,N_10198);
nand U12492 (N_12492,N_10146,N_10675);
or U12493 (N_12493,N_11123,N_10301);
nand U12494 (N_12494,N_10729,N_10635);
and U12495 (N_12495,N_10245,N_10172);
nor U12496 (N_12496,N_10235,N_11393);
or U12497 (N_12497,N_10784,N_10364);
or U12498 (N_12498,N_11107,N_11679);
nand U12499 (N_12499,N_10066,N_10032);
xnor U12500 (N_12500,N_11755,N_11948);
nor U12501 (N_12501,N_11861,N_11312);
nand U12502 (N_12502,N_11503,N_11175);
or U12503 (N_12503,N_11475,N_10639);
xor U12504 (N_12504,N_11051,N_11905);
or U12505 (N_12505,N_10911,N_10108);
nand U12506 (N_12506,N_11818,N_10173);
or U12507 (N_12507,N_10705,N_11424);
or U12508 (N_12508,N_10988,N_10708);
nor U12509 (N_12509,N_11003,N_10454);
or U12510 (N_12510,N_10244,N_10501);
or U12511 (N_12511,N_11822,N_10873);
nand U12512 (N_12512,N_10924,N_10399);
or U12513 (N_12513,N_11363,N_11634);
or U12514 (N_12514,N_10408,N_11588);
nor U12515 (N_12515,N_10727,N_10206);
nand U12516 (N_12516,N_10258,N_11529);
and U12517 (N_12517,N_10056,N_11685);
and U12518 (N_12518,N_10202,N_10760);
and U12519 (N_12519,N_10562,N_11540);
nor U12520 (N_12520,N_10062,N_11142);
nor U12521 (N_12521,N_11345,N_11584);
nand U12522 (N_12522,N_10663,N_10661);
nor U12523 (N_12523,N_10360,N_11977);
nand U12524 (N_12524,N_10325,N_11620);
nor U12525 (N_12525,N_10411,N_11336);
nor U12526 (N_12526,N_10866,N_10831);
nor U12527 (N_12527,N_11039,N_11431);
nand U12528 (N_12528,N_10385,N_11071);
nand U12529 (N_12529,N_10806,N_10416);
and U12530 (N_12530,N_10754,N_10974);
nand U12531 (N_12531,N_11745,N_10985);
xor U12532 (N_12532,N_11138,N_10556);
or U12533 (N_12533,N_11179,N_10419);
or U12534 (N_12534,N_10591,N_10358);
and U12535 (N_12535,N_11059,N_11759);
nand U12536 (N_12536,N_11478,N_11402);
nor U12537 (N_12537,N_11260,N_10005);
nand U12538 (N_12538,N_11169,N_11288);
or U12539 (N_12539,N_11356,N_10941);
and U12540 (N_12540,N_10928,N_10724);
and U12541 (N_12541,N_10133,N_10161);
nand U12542 (N_12542,N_10839,N_11598);
or U12543 (N_12543,N_10676,N_11841);
nor U12544 (N_12544,N_11986,N_10986);
or U12545 (N_12545,N_11158,N_11945);
or U12546 (N_12546,N_11637,N_10908);
nand U12547 (N_12547,N_10931,N_10260);
nand U12548 (N_12548,N_11112,N_10223);
or U12549 (N_12549,N_11556,N_10523);
nor U12550 (N_12550,N_10327,N_10681);
or U12551 (N_12551,N_11454,N_11474);
nand U12552 (N_12552,N_10334,N_10386);
nand U12553 (N_12553,N_10600,N_10162);
and U12554 (N_12554,N_11795,N_11916);
and U12555 (N_12555,N_10261,N_10665);
and U12556 (N_12556,N_10090,N_10491);
or U12557 (N_12557,N_10842,N_10939);
and U12558 (N_12558,N_10900,N_10016);
nand U12559 (N_12559,N_10859,N_11208);
and U12560 (N_12560,N_10570,N_10592);
and U12561 (N_12561,N_10780,N_11302);
or U12562 (N_12562,N_10825,N_11485);
nand U12563 (N_12563,N_10714,N_10366);
nor U12564 (N_12564,N_11807,N_10721);
or U12565 (N_12565,N_10526,N_11101);
nor U12566 (N_12566,N_10495,N_10481);
nor U12567 (N_12567,N_11980,N_10080);
nand U12568 (N_12568,N_11068,N_11920);
and U12569 (N_12569,N_11147,N_11799);
nor U12570 (N_12570,N_10613,N_10388);
xor U12571 (N_12571,N_11043,N_10978);
xor U12572 (N_12572,N_10543,N_10229);
nor U12573 (N_12573,N_10292,N_11245);
nor U12574 (N_12574,N_10595,N_11764);
nor U12575 (N_12575,N_11924,N_11163);
or U12576 (N_12576,N_11368,N_10576);
or U12577 (N_12577,N_10876,N_10070);
or U12578 (N_12578,N_10853,N_11714);
nand U12579 (N_12579,N_11796,N_10510);
and U12580 (N_12580,N_10332,N_10082);
nand U12581 (N_12581,N_11919,N_11803);
nand U12582 (N_12582,N_10237,N_11385);
nor U12583 (N_12583,N_10402,N_11698);
nor U12584 (N_12584,N_11864,N_11437);
nand U12585 (N_12585,N_11088,N_11131);
nor U12586 (N_12586,N_10135,N_10186);
or U12587 (N_12587,N_10770,N_11808);
nor U12588 (N_12588,N_10201,N_11089);
and U12589 (N_12589,N_11121,N_11074);
and U12590 (N_12590,N_11378,N_11738);
xnor U12591 (N_12591,N_11872,N_11639);
or U12592 (N_12592,N_11216,N_10494);
nor U12593 (N_12593,N_11760,N_10743);
or U12594 (N_12594,N_10440,N_11893);
nand U12595 (N_12595,N_11370,N_10389);
or U12596 (N_12596,N_11319,N_11829);
or U12597 (N_12597,N_10312,N_10996);
xnor U12598 (N_12598,N_11883,N_11962);
or U12599 (N_12599,N_11063,N_11885);
and U12600 (N_12600,N_10896,N_10031);
and U12601 (N_12601,N_10368,N_11286);
nand U12602 (N_12602,N_11269,N_11111);
nand U12603 (N_12603,N_10014,N_11561);
nand U12604 (N_12604,N_10275,N_10645);
or U12605 (N_12605,N_10958,N_11130);
and U12606 (N_12606,N_10246,N_11701);
and U12607 (N_12607,N_10772,N_10287);
nor U12608 (N_12608,N_10075,N_10120);
or U12609 (N_12609,N_10565,N_11463);
or U12610 (N_12610,N_10710,N_11044);
and U12611 (N_12611,N_10111,N_11299);
or U12612 (N_12612,N_11391,N_11186);
nor U12613 (N_12613,N_11218,N_11898);
and U12614 (N_12614,N_11900,N_11843);
nor U12615 (N_12615,N_10943,N_11926);
nand U12616 (N_12616,N_10982,N_10023);
nand U12617 (N_12617,N_11126,N_11859);
nand U12618 (N_12618,N_11093,N_10269);
nor U12619 (N_12619,N_10039,N_11733);
or U12620 (N_12620,N_11072,N_11027);
or U12621 (N_12621,N_11476,N_10575);
nor U12622 (N_12622,N_10482,N_10628);
and U12623 (N_12623,N_10101,N_10899);
and U12624 (N_12624,N_11473,N_11982);
or U12625 (N_12625,N_10709,N_10125);
or U12626 (N_12626,N_11950,N_11316);
nor U12627 (N_12627,N_11376,N_10147);
nand U12628 (N_12628,N_11909,N_10891);
nand U12629 (N_12629,N_10165,N_10224);
nand U12630 (N_12630,N_10461,N_11555);
nand U12631 (N_12631,N_10834,N_10274);
nand U12632 (N_12632,N_11386,N_10012);
and U12633 (N_12633,N_10867,N_11703);
and U12634 (N_12634,N_11797,N_11772);
nand U12635 (N_12635,N_11673,N_11444);
nand U12636 (N_12636,N_10655,N_10586);
and U12637 (N_12637,N_11603,N_10412);
or U12638 (N_12638,N_11090,N_10688);
nand U12639 (N_12639,N_11804,N_11610);
nand U12640 (N_12640,N_11983,N_11988);
nor U12641 (N_12641,N_11468,N_10905);
and U12642 (N_12642,N_10468,N_11028);
and U12643 (N_12643,N_11400,N_10880);
or U12644 (N_12644,N_11519,N_11521);
or U12645 (N_12645,N_10236,N_11936);
and U12646 (N_12646,N_11728,N_11239);
xor U12647 (N_12647,N_11398,N_10458);
nand U12648 (N_12648,N_10764,N_10415);
nor U12649 (N_12649,N_11635,N_11164);
xor U12650 (N_12650,N_10239,N_10438);
nor U12651 (N_12651,N_10456,N_10530);
nand U12652 (N_12652,N_10856,N_10141);
nor U12653 (N_12653,N_11869,N_10187);
nand U12654 (N_12654,N_10057,N_11106);
nand U12655 (N_12655,N_10463,N_10096);
xnor U12656 (N_12656,N_11049,N_11231);
xor U12657 (N_12657,N_10320,N_10752);
xnor U12658 (N_12658,N_11662,N_11203);
xnor U12659 (N_12659,N_10435,N_11489);
or U12660 (N_12660,N_10923,N_11517);
nor U12661 (N_12661,N_10742,N_10851);
nand U12662 (N_12662,N_11871,N_11794);
nor U12663 (N_12663,N_11460,N_10054);
nor U12664 (N_12664,N_10083,N_11145);
nor U12665 (N_12665,N_10316,N_10718);
nor U12666 (N_12666,N_10475,N_10150);
nor U12667 (N_12667,N_10981,N_10397);
nand U12668 (N_12668,N_11167,N_10050);
or U12669 (N_12669,N_11395,N_11360);
and U12670 (N_12670,N_11104,N_10034);
and U12671 (N_12671,N_11923,N_11601);
nor U12672 (N_12672,N_11914,N_10439);
nand U12673 (N_12673,N_10451,N_11367);
or U12674 (N_12674,N_11704,N_11903);
and U12675 (N_12675,N_11934,N_11518);
nand U12676 (N_12676,N_11559,N_11467);
nor U12677 (N_12677,N_10256,N_10181);
nand U12678 (N_12678,N_11577,N_10756);
nor U12679 (N_12679,N_11244,N_10304);
nand U12680 (N_12680,N_10912,N_11450);
nor U12681 (N_12681,N_10741,N_10427);
and U12682 (N_12682,N_11058,N_10371);
nor U12683 (N_12683,N_11955,N_10648);
nor U12684 (N_12684,N_11082,N_11549);
xnor U12685 (N_12685,N_10249,N_10255);
or U12686 (N_12686,N_11338,N_10095);
or U12687 (N_12687,N_10270,N_10877);
nand U12688 (N_12688,N_11758,N_10047);
nand U12689 (N_12689,N_10073,N_10926);
or U12690 (N_12690,N_10744,N_11817);
nand U12691 (N_12691,N_10844,N_10991);
nand U12692 (N_12692,N_11470,N_11141);
or U12693 (N_12693,N_10995,N_10881);
or U12694 (N_12694,N_10773,N_11193);
and U12695 (N_12695,N_11401,N_10952);
nand U12696 (N_12696,N_10580,N_10611);
nor U12697 (N_12697,N_10622,N_11070);
or U12698 (N_12698,N_10597,N_10984);
or U12699 (N_12699,N_10636,N_11615);
nand U12700 (N_12700,N_11970,N_10534);
nand U12701 (N_12701,N_11325,N_11579);
nand U12702 (N_12702,N_11657,N_10105);
nand U12703 (N_12703,N_11314,N_11692);
nand U12704 (N_12704,N_10506,N_10895);
or U12705 (N_12705,N_11836,N_11132);
nand U12706 (N_12706,N_10184,N_11879);
nand U12707 (N_12707,N_11436,N_10608);
nand U12708 (N_12708,N_11388,N_11624);
nor U12709 (N_12709,N_10915,N_11992);
or U12710 (N_12710,N_11542,N_10849);
or U12711 (N_12711,N_11060,N_10723);
or U12712 (N_12712,N_10200,N_11413);
and U12713 (N_12713,N_11277,N_10536);
nand U12714 (N_12714,N_11178,N_10625);
or U12715 (N_12715,N_10858,N_11073);
nand U12716 (N_12716,N_10740,N_11000);
and U12717 (N_12717,N_10295,N_10667);
or U12718 (N_12718,N_11993,N_10299);
nor U12719 (N_12719,N_11741,N_11272);
nand U12720 (N_12720,N_11149,N_10069);
or U12721 (N_12721,N_10029,N_11189);
or U12722 (N_12722,N_11223,N_11046);
nand U12723 (N_12723,N_10687,N_10317);
and U12724 (N_12724,N_10283,N_11984);
nand U12725 (N_12725,N_10607,N_10620);
xnor U12726 (N_12726,N_10804,N_11284);
and U12727 (N_12727,N_11973,N_11331);
nor U12728 (N_12728,N_11484,N_10658);
and U12729 (N_12729,N_11494,N_10983);
nor U12730 (N_12730,N_10666,N_10183);
nand U12731 (N_12731,N_11144,N_10466);
or U12732 (N_12732,N_11137,N_11265);
nor U12733 (N_12733,N_11005,N_11133);
and U12734 (N_12734,N_10294,N_10572);
or U12735 (N_12735,N_11653,N_11421);
nor U12736 (N_12736,N_10901,N_11630);
or U12737 (N_12737,N_10042,N_11459);
xor U12738 (N_12738,N_11352,N_11557);
and U12739 (N_12739,N_11749,N_10006);
nor U12740 (N_12740,N_10281,N_11767);
nor U12741 (N_12741,N_11469,N_11053);
or U12742 (N_12742,N_11161,N_10887);
and U12743 (N_12743,N_11514,N_11007);
or U12744 (N_12744,N_11952,N_11538);
and U12745 (N_12745,N_10035,N_11709);
nor U12746 (N_12746,N_10359,N_11513);
nand U12747 (N_12747,N_10935,N_11118);
nor U12748 (N_12748,N_10782,N_11477);
nor U12749 (N_12749,N_11320,N_10305);
or U12750 (N_12750,N_10174,N_11290);
or U12751 (N_12751,N_11304,N_10449);
nor U12752 (N_12752,N_11045,N_10257);
and U12753 (N_12753,N_11456,N_11525);
xor U12754 (N_12754,N_10212,N_11853);
and U12755 (N_12755,N_10442,N_11769);
and U12756 (N_12756,N_10791,N_11308);
nor U12757 (N_12757,N_11065,N_11614);
and U12758 (N_12758,N_11500,N_10024);
nand U12759 (N_12759,N_11946,N_10537);
and U12760 (N_12760,N_11030,N_10745);
or U12761 (N_12761,N_11412,N_10746);
and U12762 (N_12762,N_10277,N_10136);
and U12763 (N_12763,N_10321,N_11642);
or U12764 (N_12764,N_10302,N_11682);
and U12765 (N_12765,N_11783,N_11055);
and U12766 (N_12766,N_10732,N_10390);
or U12767 (N_12767,N_10517,N_10396);
nor U12768 (N_12768,N_10448,N_10792);
nand U12769 (N_12769,N_11258,N_11813);
xor U12770 (N_12770,N_11787,N_10472);
nor U12771 (N_12771,N_10957,N_10285);
xnor U12772 (N_12772,N_10155,N_11498);
xnor U12773 (N_12773,N_10121,N_10008);
xor U12774 (N_12774,N_11626,N_11801);
nand U12775 (N_12775,N_10092,N_10436);
or U12776 (N_12776,N_10059,N_11677);
and U12777 (N_12777,N_10341,N_11496);
nor U12778 (N_12778,N_10789,N_11719);
xor U12779 (N_12779,N_10076,N_10467);
nor U12780 (N_12780,N_10922,N_10757);
nand U12781 (N_12781,N_10377,N_11033);
or U12782 (N_12782,N_10215,N_11201);
nor U12783 (N_12783,N_11509,N_11789);
nor U12784 (N_12784,N_11890,N_10557);
and U12785 (N_12785,N_10303,N_11675);
nor U12786 (N_12786,N_11499,N_11508);
and U12787 (N_12787,N_10779,N_10884);
nor U12788 (N_12788,N_11198,N_11581);
and U12789 (N_12789,N_11199,N_10711);
or U12790 (N_12790,N_11453,N_11729);
or U12791 (N_12791,N_11771,N_11114);
xnor U12792 (N_12792,N_10038,N_11032);
nand U12793 (N_12793,N_11546,N_11094);
xor U12794 (N_12794,N_11206,N_10289);
or U12795 (N_12795,N_10528,N_10276);
nand U12796 (N_12796,N_10604,N_11827);
or U12797 (N_12797,N_11214,N_11933);
and U12798 (N_12798,N_10716,N_11160);
nand U12799 (N_12799,N_11471,N_10311);
nand U12800 (N_12800,N_10131,N_10722);
xnor U12801 (N_12801,N_11592,N_10680);
nand U12802 (N_12802,N_11440,N_10818);
xnor U12803 (N_12803,N_10351,N_11552);
nor U12804 (N_12804,N_11705,N_10123);
nor U12805 (N_12805,N_11404,N_11686);
nor U12806 (N_12806,N_10559,N_10547);
xnor U12807 (N_12807,N_10826,N_10036);
nand U12808 (N_12808,N_11964,N_11876);
and U12809 (N_12809,N_11687,N_10797);
and U12810 (N_12810,N_11337,N_10967);
nor U12811 (N_12811,N_11289,N_11213);
nand U12812 (N_12812,N_11347,N_10021);
and U12813 (N_12813,N_11136,N_10037);
nand U12814 (N_12814,N_11100,N_10149);
and U12815 (N_12815,N_11868,N_11052);
nand U12816 (N_12816,N_11418,N_11491);
or U12817 (N_12817,N_11960,N_11737);
and U12818 (N_12818,N_10113,N_11374);
nand U12819 (N_12819,N_11591,N_10367);
or U12820 (N_12820,N_11773,N_10382);
nor U12821 (N_12821,N_11617,N_10043);
and U12822 (N_12822,N_11608,N_10498);
and U12823 (N_12823,N_10573,N_10731);
or U12824 (N_12824,N_10821,N_11897);
and U12825 (N_12825,N_11422,N_10650);
nor U12826 (N_12826,N_11176,N_11026);
and U12827 (N_12827,N_11173,N_11785);
and U12828 (N_12828,N_11493,N_11722);
and U12829 (N_12829,N_11184,N_11567);
nand U12830 (N_12830,N_11018,N_11721);
and U12831 (N_12831,N_11001,N_11839);
or U12832 (N_12832,N_10819,N_11633);
nand U12833 (N_12833,N_11638,N_11102);
nand U12834 (N_12834,N_10496,N_10837);
nor U12835 (N_12835,N_11311,N_10019);
nor U12836 (N_12836,N_10180,N_10132);
nor U12837 (N_12837,N_11105,N_10340);
nor U12838 (N_12838,N_11541,N_10296);
nand U12839 (N_12839,N_11326,N_11466);
nor U12840 (N_12840,N_10242,N_11668);
xnor U12841 (N_12841,N_11851,N_11227);
and U12842 (N_12842,N_10612,N_10860);
nand U12843 (N_12843,N_10102,N_10807);
xnor U12844 (N_12844,N_10614,N_10865);
nand U12845 (N_12845,N_10601,N_11254);
or U12846 (N_12846,N_10581,N_10847);
or U12847 (N_12847,N_10972,N_10909);
xor U12848 (N_12848,N_10814,N_11086);
nand U12849 (N_12849,N_10384,N_11449);
and U12850 (N_12850,N_10450,N_11524);
nor U12851 (N_12851,N_10033,N_10527);
nor U12852 (N_12852,N_11862,N_10348);
nand U12853 (N_12853,N_11282,N_11358);
or U12854 (N_12854,N_10554,N_11968);
or U12855 (N_12855,N_11441,N_11571);
and U12856 (N_12856,N_10480,N_11406);
nor U12857 (N_12857,N_10747,N_10290);
and U12858 (N_12858,N_11917,N_10917);
or U12859 (N_12859,N_11572,N_11696);
xor U12860 (N_12860,N_10513,N_11383);
nor U12861 (N_12861,N_10690,N_11654);
nand U12862 (N_12862,N_11207,N_10827);
or U12863 (N_12863,N_10553,N_10065);
or U12864 (N_12864,N_11516,N_10567);
nor U12865 (N_12865,N_10535,N_11956);
nor U12866 (N_12866,N_10009,N_10192);
and U12867 (N_12867,N_10793,N_11754);
and U12868 (N_12868,N_11820,N_10848);
nand U12869 (N_12869,N_10617,N_10934);
or U12870 (N_12870,N_10765,N_10426);
and U12871 (N_12871,N_11394,N_10207);
nor U12872 (N_12872,N_11457,N_11944);
and U12873 (N_12873,N_10251,N_10129);
and U12874 (N_12874,N_11237,N_10177);
and U12875 (N_12875,N_11575,N_11021);
or U12876 (N_12876,N_10898,N_11036);
nor U12877 (N_12877,N_11969,N_10194);
xnor U12878 (N_12878,N_11185,N_10064);
nand U12879 (N_12879,N_11660,N_11408);
nor U12880 (N_12880,N_10379,N_11611);
or U12881 (N_12881,N_11181,N_10560);
and U12882 (N_12882,N_11110,N_11766);
nand U12883 (N_12883,N_10892,N_10603);
xor U12884 (N_12884,N_11600,N_10254);
nor U12885 (N_12885,N_10894,N_10421);
nand U12886 (N_12886,N_11886,N_11997);
and U12887 (N_12887,N_10378,N_11067);
nand U12888 (N_12888,N_11812,N_11490);
or U12889 (N_12889,N_11157,N_11419);
nand U12890 (N_12890,N_11300,N_11574);
nand U12891 (N_12891,N_11761,N_10489);
nor U12892 (N_12892,N_10234,N_11162);
nand U12893 (N_12893,N_11355,N_10049);
nor U12894 (N_12894,N_10916,N_10476);
and U12895 (N_12895,N_10945,N_11205);
or U12896 (N_12896,N_11342,N_11666);
or U12897 (N_12897,N_10100,N_11285);
or U12898 (N_12898,N_11512,N_11029);
or U12899 (N_12899,N_10336,N_11953);
nand U12900 (N_12900,N_10816,N_10621);
nand U12901 (N_12901,N_10888,N_10678);
and U12902 (N_12902,N_10694,N_11583);
and U12903 (N_12903,N_11448,N_10291);
nor U12904 (N_12904,N_10118,N_11061);
nor U12905 (N_12905,N_10343,N_11782);
nand U12906 (N_12906,N_11343,N_11590);
and U12907 (N_12907,N_10094,N_10445);
nand U12908 (N_12908,N_11563,N_10781);
or U12909 (N_12909,N_10193,N_11165);
and U12910 (N_12910,N_10479,N_11180);
and U12911 (N_12911,N_10051,N_11264);
and U12912 (N_12912,N_10081,N_11301);
nand U12913 (N_12913,N_11727,N_11830);
nor U12914 (N_12914,N_10114,N_10273);
nor U12915 (N_12915,N_10117,N_11317);
and U12916 (N_12916,N_11445,N_10919);
or U12917 (N_12917,N_11472,N_10664);
or U12918 (N_12918,N_11407,N_11793);
and U12919 (N_12919,N_11669,N_11844);
nand U12920 (N_12920,N_10907,N_11344);
and U12921 (N_12921,N_10017,N_10232);
and U12922 (N_12922,N_10893,N_11664);
nor U12923 (N_12923,N_10195,N_11912);
xor U12924 (N_12924,N_10868,N_11420);
and U12925 (N_12925,N_10846,N_10074);
nand U12926 (N_12926,N_10393,N_11753);
nor U12927 (N_12927,N_11976,N_11536);
xor U12928 (N_12928,N_10167,N_10205);
or U12929 (N_12929,N_10361,N_11860);
or U12930 (N_12930,N_11947,N_10929);
nor U12931 (N_12931,N_10725,N_10810);
and U12932 (N_12932,N_11122,N_11197);
nor U12933 (N_12933,N_10363,N_10112);
and U12934 (N_12934,N_11023,N_10434);
nor U12935 (N_12935,N_10533,N_10465);
or U12936 (N_12936,N_10977,N_11066);
or U12937 (N_12937,N_11321,N_10505);
and U12938 (N_12938,N_11334,N_11954);
nor U12939 (N_12939,N_10624,N_11024);
nor U12940 (N_12940,N_11379,N_10013);
nor U12941 (N_12941,N_10833,N_10078);
nand U12942 (N_12942,N_10375,N_10921);
and U12943 (N_12943,N_10897,N_10433);
or U12944 (N_12944,N_10015,N_10225);
nand U12945 (N_12945,N_10577,N_11875);
nor U12946 (N_12946,N_11364,N_10739);
and U12947 (N_12947,N_11140,N_10469);
and U12948 (N_12948,N_11225,N_11743);
xnor U12949 (N_12949,N_10964,N_10713);
nor U12950 (N_12950,N_10058,N_10598);
or U12951 (N_12951,N_11904,N_10151);
or U12952 (N_12952,N_10602,N_11725);
and U12953 (N_12953,N_11607,N_11672);
nor U12954 (N_12954,N_10585,N_10091);
nand U12955 (N_12955,N_10692,N_10966);
and U12956 (N_12956,N_10171,N_11425);
nor U12957 (N_12957,N_10474,N_11429);
xnor U12958 (N_12958,N_11825,N_11416);
and U12959 (N_12959,N_11833,N_11085);
nor U12960 (N_12960,N_11414,N_10717);
nor U12961 (N_12961,N_10499,N_11506);
or U12962 (N_12962,N_10214,N_11306);
xnor U12963 (N_12963,N_10749,N_11645);
nand U12964 (N_12964,N_10763,N_11266);
nand U12965 (N_12965,N_10561,N_11332);
xnor U12966 (N_12966,N_11531,N_10767);
and U12967 (N_12967,N_11802,N_11826);
or U12968 (N_12968,N_10300,N_10280);
nor U12969 (N_12969,N_10452,N_11650);
and U12970 (N_12970,N_11297,N_11405);
or U12971 (N_12971,N_11148,N_10139);
nor U12972 (N_12972,N_10910,N_10890);
or U12973 (N_12973,N_10020,N_10950);
and U12974 (N_12974,N_11250,N_11380);
nor U12975 (N_12975,N_10085,N_10652);
nor U12976 (N_12976,N_10925,N_10353);
and U12977 (N_12977,N_11329,N_10769);
and U12978 (N_12978,N_10542,N_10189);
or U12979 (N_12979,N_10410,N_10087);
nand U12980 (N_12980,N_10686,N_11081);
nand U12981 (N_12981,N_10820,N_10293);
nor U12982 (N_12982,N_11658,N_10154);
nand U12983 (N_12983,N_11215,N_10590);
nor U12984 (N_12984,N_11154,N_10647);
nand U12985 (N_12985,N_11228,N_11209);
and U12986 (N_12986,N_10812,N_11155);
or U12987 (N_12987,N_10443,N_11447);
nor U12988 (N_12988,N_11129,N_11963);
nand U12989 (N_12989,N_11016,N_10695);
and U12990 (N_12990,N_11554,N_10904);
nor U12991 (N_12991,N_10286,N_10182);
nand U12992 (N_12992,N_10777,N_11222);
nand U12993 (N_12993,N_11640,N_11837);
nor U12994 (N_12994,N_11341,N_10413);
or U12995 (N_12995,N_11805,N_11606);
xnor U12996 (N_12996,N_11428,N_11593);
and U12997 (N_12997,N_10428,N_11504);
nand U12998 (N_12998,N_11487,N_10660);
and U12999 (N_12999,N_10940,N_10630);
and U13000 (N_13000,N_10340,N_10984);
nor U13001 (N_13001,N_11756,N_10285);
or U13002 (N_13002,N_10944,N_11300);
nand U13003 (N_13003,N_11719,N_11464);
or U13004 (N_13004,N_11057,N_11378);
xnor U13005 (N_13005,N_11296,N_11838);
or U13006 (N_13006,N_11608,N_10236);
and U13007 (N_13007,N_10664,N_11995);
xor U13008 (N_13008,N_10189,N_10362);
or U13009 (N_13009,N_11357,N_11983);
nand U13010 (N_13010,N_11006,N_10583);
and U13011 (N_13011,N_11474,N_11040);
and U13012 (N_13012,N_10711,N_10649);
nand U13013 (N_13013,N_10814,N_10640);
and U13014 (N_13014,N_10863,N_10787);
nor U13015 (N_13015,N_10791,N_10050);
and U13016 (N_13016,N_10943,N_11815);
nand U13017 (N_13017,N_11608,N_11372);
and U13018 (N_13018,N_11848,N_10326);
nor U13019 (N_13019,N_11797,N_11873);
nand U13020 (N_13020,N_10434,N_10896);
nand U13021 (N_13021,N_10965,N_10433);
nor U13022 (N_13022,N_11730,N_11311);
and U13023 (N_13023,N_11446,N_10960);
nor U13024 (N_13024,N_11141,N_10434);
or U13025 (N_13025,N_11935,N_10454);
nand U13026 (N_13026,N_10783,N_10093);
or U13027 (N_13027,N_11281,N_11206);
and U13028 (N_13028,N_11118,N_11236);
nand U13029 (N_13029,N_11428,N_11247);
xnor U13030 (N_13030,N_11596,N_10176);
xnor U13031 (N_13031,N_11669,N_10425);
nand U13032 (N_13032,N_11782,N_10667);
or U13033 (N_13033,N_11171,N_10991);
xnor U13034 (N_13034,N_10737,N_10704);
and U13035 (N_13035,N_11065,N_11550);
nor U13036 (N_13036,N_10637,N_10153);
and U13037 (N_13037,N_11794,N_11013);
nand U13038 (N_13038,N_10766,N_10360);
nand U13039 (N_13039,N_11356,N_11629);
nor U13040 (N_13040,N_11874,N_11993);
xor U13041 (N_13041,N_10633,N_10720);
nand U13042 (N_13042,N_11901,N_10714);
and U13043 (N_13043,N_10031,N_10587);
nand U13044 (N_13044,N_10318,N_10186);
nor U13045 (N_13045,N_10554,N_11721);
nor U13046 (N_13046,N_11580,N_11298);
nor U13047 (N_13047,N_11587,N_10998);
or U13048 (N_13048,N_10263,N_11358);
or U13049 (N_13049,N_11116,N_10771);
or U13050 (N_13050,N_11444,N_10153);
nor U13051 (N_13051,N_10042,N_10014);
or U13052 (N_13052,N_11180,N_11962);
and U13053 (N_13053,N_10029,N_10443);
nand U13054 (N_13054,N_10294,N_10528);
nand U13055 (N_13055,N_10018,N_10562);
and U13056 (N_13056,N_11165,N_11671);
and U13057 (N_13057,N_11224,N_11821);
nor U13058 (N_13058,N_10051,N_10588);
and U13059 (N_13059,N_11885,N_11389);
nand U13060 (N_13060,N_10232,N_10185);
nor U13061 (N_13061,N_11339,N_11490);
or U13062 (N_13062,N_10395,N_10388);
nor U13063 (N_13063,N_11071,N_11225);
nor U13064 (N_13064,N_11465,N_10087);
nand U13065 (N_13065,N_11581,N_11641);
nand U13066 (N_13066,N_10249,N_11136);
and U13067 (N_13067,N_10514,N_10518);
xnor U13068 (N_13068,N_11824,N_11209);
or U13069 (N_13069,N_10535,N_11762);
nand U13070 (N_13070,N_10489,N_10564);
xnor U13071 (N_13071,N_11119,N_11416);
nand U13072 (N_13072,N_10211,N_11940);
nor U13073 (N_13073,N_10418,N_11753);
nor U13074 (N_13074,N_11137,N_11414);
nor U13075 (N_13075,N_11942,N_10951);
nand U13076 (N_13076,N_11314,N_11052);
nand U13077 (N_13077,N_10903,N_11484);
and U13078 (N_13078,N_10746,N_10484);
and U13079 (N_13079,N_11042,N_11898);
or U13080 (N_13080,N_10548,N_11122);
and U13081 (N_13081,N_11620,N_10786);
nand U13082 (N_13082,N_11865,N_11081);
nor U13083 (N_13083,N_10014,N_10346);
nand U13084 (N_13084,N_10434,N_10127);
nor U13085 (N_13085,N_10449,N_10855);
nor U13086 (N_13086,N_11852,N_10776);
or U13087 (N_13087,N_11034,N_11789);
or U13088 (N_13088,N_10100,N_10966);
nand U13089 (N_13089,N_11369,N_10426);
or U13090 (N_13090,N_11883,N_11767);
and U13091 (N_13091,N_10045,N_10003);
and U13092 (N_13092,N_11989,N_10781);
or U13093 (N_13093,N_10492,N_10835);
or U13094 (N_13094,N_11212,N_11555);
nor U13095 (N_13095,N_11700,N_11529);
xnor U13096 (N_13096,N_10978,N_11660);
nand U13097 (N_13097,N_10122,N_10635);
and U13098 (N_13098,N_10130,N_11534);
and U13099 (N_13099,N_10281,N_10556);
nand U13100 (N_13100,N_11791,N_10689);
and U13101 (N_13101,N_11772,N_10136);
xor U13102 (N_13102,N_11431,N_11425);
nor U13103 (N_13103,N_10591,N_10534);
nor U13104 (N_13104,N_10878,N_10970);
xor U13105 (N_13105,N_10138,N_11931);
xor U13106 (N_13106,N_10216,N_11210);
nand U13107 (N_13107,N_10024,N_11063);
or U13108 (N_13108,N_11242,N_10485);
or U13109 (N_13109,N_11815,N_11768);
nor U13110 (N_13110,N_10933,N_10589);
and U13111 (N_13111,N_10268,N_11525);
nand U13112 (N_13112,N_10581,N_11376);
xor U13113 (N_13113,N_10753,N_11358);
nor U13114 (N_13114,N_11871,N_11893);
or U13115 (N_13115,N_10296,N_11187);
xnor U13116 (N_13116,N_10804,N_10401);
or U13117 (N_13117,N_11113,N_11843);
nand U13118 (N_13118,N_11462,N_10458);
nor U13119 (N_13119,N_11933,N_10587);
and U13120 (N_13120,N_10133,N_11849);
or U13121 (N_13121,N_10044,N_10172);
and U13122 (N_13122,N_11708,N_10957);
nand U13123 (N_13123,N_10035,N_10412);
nand U13124 (N_13124,N_11758,N_11741);
and U13125 (N_13125,N_11587,N_11570);
xnor U13126 (N_13126,N_11757,N_10027);
and U13127 (N_13127,N_11517,N_11287);
xnor U13128 (N_13128,N_10792,N_11398);
nand U13129 (N_13129,N_10749,N_10864);
nor U13130 (N_13130,N_11168,N_10543);
and U13131 (N_13131,N_10776,N_10212);
and U13132 (N_13132,N_11249,N_10727);
nor U13133 (N_13133,N_11999,N_10405);
or U13134 (N_13134,N_11758,N_10711);
nand U13135 (N_13135,N_11272,N_10755);
xnor U13136 (N_13136,N_10276,N_11993);
nor U13137 (N_13137,N_10653,N_10026);
nor U13138 (N_13138,N_10168,N_10317);
or U13139 (N_13139,N_10042,N_10513);
and U13140 (N_13140,N_11418,N_10689);
and U13141 (N_13141,N_10095,N_11737);
nor U13142 (N_13142,N_11002,N_11448);
and U13143 (N_13143,N_11833,N_10421);
and U13144 (N_13144,N_11592,N_10180);
xnor U13145 (N_13145,N_11655,N_11872);
and U13146 (N_13146,N_10654,N_10636);
xor U13147 (N_13147,N_11699,N_10572);
and U13148 (N_13148,N_11053,N_10717);
or U13149 (N_13149,N_11375,N_11116);
xnor U13150 (N_13150,N_11831,N_11567);
nand U13151 (N_13151,N_10107,N_10416);
and U13152 (N_13152,N_10069,N_11632);
or U13153 (N_13153,N_10023,N_11244);
nand U13154 (N_13154,N_11573,N_10577);
nor U13155 (N_13155,N_10346,N_10581);
and U13156 (N_13156,N_10693,N_10451);
or U13157 (N_13157,N_10439,N_11072);
and U13158 (N_13158,N_10333,N_11246);
or U13159 (N_13159,N_11427,N_10722);
nor U13160 (N_13160,N_11763,N_10749);
xor U13161 (N_13161,N_11409,N_11004);
nand U13162 (N_13162,N_10230,N_10327);
nand U13163 (N_13163,N_10042,N_10244);
nor U13164 (N_13164,N_10527,N_11503);
nor U13165 (N_13165,N_11431,N_10187);
xor U13166 (N_13166,N_11008,N_10573);
nand U13167 (N_13167,N_11227,N_11610);
nand U13168 (N_13168,N_10130,N_10090);
and U13169 (N_13169,N_10673,N_11651);
or U13170 (N_13170,N_10136,N_11347);
nand U13171 (N_13171,N_10762,N_10389);
nand U13172 (N_13172,N_10384,N_11569);
nand U13173 (N_13173,N_11100,N_10367);
and U13174 (N_13174,N_10989,N_10397);
and U13175 (N_13175,N_10307,N_10264);
or U13176 (N_13176,N_11259,N_11265);
and U13177 (N_13177,N_10708,N_11050);
nor U13178 (N_13178,N_10611,N_10170);
and U13179 (N_13179,N_10650,N_10786);
nor U13180 (N_13180,N_10457,N_11370);
or U13181 (N_13181,N_10430,N_10469);
and U13182 (N_13182,N_11585,N_10870);
or U13183 (N_13183,N_10959,N_10324);
or U13184 (N_13184,N_10548,N_11532);
nor U13185 (N_13185,N_10122,N_11911);
nand U13186 (N_13186,N_10366,N_10846);
and U13187 (N_13187,N_11224,N_10767);
nor U13188 (N_13188,N_11876,N_10394);
xnor U13189 (N_13189,N_10850,N_11819);
or U13190 (N_13190,N_11870,N_10757);
and U13191 (N_13191,N_10679,N_10541);
nor U13192 (N_13192,N_10130,N_11602);
and U13193 (N_13193,N_11423,N_10246);
and U13194 (N_13194,N_11885,N_11630);
nand U13195 (N_13195,N_10152,N_11865);
nand U13196 (N_13196,N_11590,N_11779);
or U13197 (N_13197,N_11280,N_11947);
nand U13198 (N_13198,N_11407,N_10251);
nor U13199 (N_13199,N_11339,N_11623);
nand U13200 (N_13200,N_11152,N_10708);
or U13201 (N_13201,N_11051,N_10700);
nor U13202 (N_13202,N_10005,N_10687);
and U13203 (N_13203,N_11989,N_10624);
or U13204 (N_13204,N_11718,N_10222);
and U13205 (N_13205,N_11517,N_10910);
xnor U13206 (N_13206,N_10962,N_11354);
nand U13207 (N_13207,N_10581,N_11865);
nand U13208 (N_13208,N_10047,N_11931);
or U13209 (N_13209,N_11824,N_11845);
nor U13210 (N_13210,N_11527,N_10342);
and U13211 (N_13211,N_11580,N_11982);
and U13212 (N_13212,N_11231,N_11811);
xnor U13213 (N_13213,N_10205,N_10565);
nand U13214 (N_13214,N_11870,N_11939);
nand U13215 (N_13215,N_11679,N_10268);
xnor U13216 (N_13216,N_10871,N_10002);
nand U13217 (N_13217,N_11179,N_10003);
and U13218 (N_13218,N_11272,N_11856);
nand U13219 (N_13219,N_10406,N_11009);
nand U13220 (N_13220,N_11343,N_10369);
nor U13221 (N_13221,N_11505,N_11356);
and U13222 (N_13222,N_10606,N_11282);
or U13223 (N_13223,N_11125,N_11262);
nand U13224 (N_13224,N_11856,N_10932);
or U13225 (N_13225,N_11275,N_10249);
nor U13226 (N_13226,N_11737,N_11065);
nor U13227 (N_13227,N_10647,N_10222);
nor U13228 (N_13228,N_10574,N_11219);
nand U13229 (N_13229,N_11259,N_10458);
or U13230 (N_13230,N_10283,N_11873);
nand U13231 (N_13231,N_10794,N_11897);
nor U13232 (N_13232,N_10854,N_11813);
and U13233 (N_13233,N_10912,N_11487);
or U13234 (N_13234,N_11080,N_11241);
nand U13235 (N_13235,N_11711,N_11415);
or U13236 (N_13236,N_11306,N_10060);
and U13237 (N_13237,N_11886,N_10801);
nor U13238 (N_13238,N_11582,N_10364);
and U13239 (N_13239,N_11487,N_10563);
and U13240 (N_13240,N_10249,N_10420);
nand U13241 (N_13241,N_11160,N_10199);
or U13242 (N_13242,N_10369,N_10711);
and U13243 (N_13243,N_11705,N_10276);
and U13244 (N_13244,N_11961,N_10394);
xnor U13245 (N_13245,N_10261,N_10050);
nand U13246 (N_13246,N_11331,N_11330);
and U13247 (N_13247,N_11823,N_10823);
and U13248 (N_13248,N_11181,N_11208);
nand U13249 (N_13249,N_10212,N_11607);
or U13250 (N_13250,N_11643,N_11414);
and U13251 (N_13251,N_10528,N_10959);
xor U13252 (N_13252,N_11596,N_10809);
nand U13253 (N_13253,N_10193,N_11624);
or U13254 (N_13254,N_11214,N_11008);
or U13255 (N_13255,N_10726,N_11326);
nand U13256 (N_13256,N_10507,N_10760);
xor U13257 (N_13257,N_11658,N_11927);
and U13258 (N_13258,N_11405,N_10885);
or U13259 (N_13259,N_10151,N_11555);
nor U13260 (N_13260,N_10807,N_11770);
nor U13261 (N_13261,N_11978,N_10139);
and U13262 (N_13262,N_11609,N_10720);
and U13263 (N_13263,N_11514,N_11276);
nor U13264 (N_13264,N_11250,N_10632);
or U13265 (N_13265,N_10429,N_11781);
and U13266 (N_13266,N_11586,N_10632);
or U13267 (N_13267,N_11059,N_11926);
nor U13268 (N_13268,N_10913,N_10701);
or U13269 (N_13269,N_11856,N_11720);
and U13270 (N_13270,N_11093,N_11895);
xor U13271 (N_13271,N_11710,N_11941);
or U13272 (N_13272,N_10349,N_10173);
nand U13273 (N_13273,N_10883,N_11827);
nor U13274 (N_13274,N_11212,N_11973);
or U13275 (N_13275,N_10362,N_11100);
and U13276 (N_13276,N_10450,N_11451);
nand U13277 (N_13277,N_11861,N_11386);
and U13278 (N_13278,N_11200,N_11538);
or U13279 (N_13279,N_10718,N_11406);
nand U13280 (N_13280,N_11158,N_11737);
and U13281 (N_13281,N_10027,N_10177);
and U13282 (N_13282,N_10560,N_10939);
nand U13283 (N_13283,N_10443,N_11883);
or U13284 (N_13284,N_11018,N_11105);
or U13285 (N_13285,N_10927,N_10813);
or U13286 (N_13286,N_10706,N_11384);
nor U13287 (N_13287,N_11504,N_10725);
nand U13288 (N_13288,N_10886,N_10372);
xor U13289 (N_13289,N_10646,N_10684);
nand U13290 (N_13290,N_10574,N_11132);
or U13291 (N_13291,N_11061,N_10617);
nand U13292 (N_13292,N_10145,N_11050);
and U13293 (N_13293,N_10499,N_11552);
nor U13294 (N_13294,N_10153,N_10025);
nand U13295 (N_13295,N_11565,N_10540);
and U13296 (N_13296,N_10503,N_10007);
and U13297 (N_13297,N_10041,N_10561);
or U13298 (N_13298,N_10108,N_10457);
and U13299 (N_13299,N_10489,N_10646);
nand U13300 (N_13300,N_11864,N_11143);
xnor U13301 (N_13301,N_10151,N_11847);
nor U13302 (N_13302,N_11508,N_11200);
and U13303 (N_13303,N_10861,N_10119);
nand U13304 (N_13304,N_10303,N_11240);
nand U13305 (N_13305,N_11538,N_10704);
nand U13306 (N_13306,N_11360,N_11560);
and U13307 (N_13307,N_11449,N_11762);
nor U13308 (N_13308,N_11483,N_10433);
nand U13309 (N_13309,N_10511,N_11719);
or U13310 (N_13310,N_11241,N_10179);
nor U13311 (N_13311,N_11596,N_11500);
nand U13312 (N_13312,N_10257,N_10126);
xnor U13313 (N_13313,N_10313,N_10672);
xor U13314 (N_13314,N_11412,N_10660);
nor U13315 (N_13315,N_11545,N_11767);
nor U13316 (N_13316,N_11017,N_11208);
xnor U13317 (N_13317,N_11400,N_11841);
nand U13318 (N_13318,N_10906,N_11015);
nand U13319 (N_13319,N_10517,N_11942);
or U13320 (N_13320,N_11237,N_10873);
nor U13321 (N_13321,N_10556,N_11209);
xor U13322 (N_13322,N_11433,N_10425);
and U13323 (N_13323,N_10915,N_10790);
or U13324 (N_13324,N_10262,N_10685);
nor U13325 (N_13325,N_10844,N_10266);
nor U13326 (N_13326,N_10469,N_11615);
or U13327 (N_13327,N_11563,N_10600);
nor U13328 (N_13328,N_11912,N_10972);
and U13329 (N_13329,N_10916,N_11784);
nor U13330 (N_13330,N_10639,N_10938);
xnor U13331 (N_13331,N_10672,N_11525);
or U13332 (N_13332,N_11452,N_10969);
or U13333 (N_13333,N_10330,N_11942);
and U13334 (N_13334,N_11541,N_11646);
xnor U13335 (N_13335,N_11618,N_11095);
or U13336 (N_13336,N_10662,N_11875);
nand U13337 (N_13337,N_10920,N_10861);
or U13338 (N_13338,N_11910,N_11278);
and U13339 (N_13339,N_11461,N_10150);
or U13340 (N_13340,N_11978,N_11532);
nor U13341 (N_13341,N_11293,N_10454);
nor U13342 (N_13342,N_11388,N_11104);
nor U13343 (N_13343,N_10735,N_10526);
nand U13344 (N_13344,N_10884,N_10413);
xnor U13345 (N_13345,N_10607,N_10059);
or U13346 (N_13346,N_11988,N_10015);
and U13347 (N_13347,N_11723,N_11607);
and U13348 (N_13348,N_10930,N_10109);
or U13349 (N_13349,N_10851,N_11360);
and U13350 (N_13350,N_11897,N_10602);
nor U13351 (N_13351,N_11653,N_11008);
and U13352 (N_13352,N_11567,N_11803);
xor U13353 (N_13353,N_11565,N_11117);
or U13354 (N_13354,N_10754,N_11970);
or U13355 (N_13355,N_10328,N_10958);
and U13356 (N_13356,N_11201,N_10391);
and U13357 (N_13357,N_10534,N_11488);
or U13358 (N_13358,N_11115,N_10677);
nand U13359 (N_13359,N_10963,N_11275);
nand U13360 (N_13360,N_10226,N_10842);
nand U13361 (N_13361,N_11990,N_11300);
nor U13362 (N_13362,N_11931,N_10858);
nor U13363 (N_13363,N_10549,N_10170);
or U13364 (N_13364,N_11769,N_11758);
nor U13365 (N_13365,N_11222,N_11790);
nand U13366 (N_13366,N_11079,N_11279);
nand U13367 (N_13367,N_11553,N_10372);
nand U13368 (N_13368,N_11968,N_11430);
and U13369 (N_13369,N_11283,N_10662);
nand U13370 (N_13370,N_10911,N_10117);
nor U13371 (N_13371,N_10898,N_10382);
nor U13372 (N_13372,N_10441,N_11007);
and U13373 (N_13373,N_11255,N_10972);
or U13374 (N_13374,N_10258,N_11401);
xnor U13375 (N_13375,N_10417,N_11555);
and U13376 (N_13376,N_11542,N_11228);
nor U13377 (N_13377,N_10418,N_11960);
and U13378 (N_13378,N_11836,N_10716);
xor U13379 (N_13379,N_11414,N_10039);
nor U13380 (N_13380,N_11266,N_11072);
nor U13381 (N_13381,N_11072,N_10661);
or U13382 (N_13382,N_10366,N_11159);
xor U13383 (N_13383,N_10187,N_10071);
and U13384 (N_13384,N_11928,N_10358);
nor U13385 (N_13385,N_10770,N_10634);
and U13386 (N_13386,N_11105,N_11914);
or U13387 (N_13387,N_10206,N_10637);
and U13388 (N_13388,N_10281,N_10036);
nor U13389 (N_13389,N_11536,N_11402);
nor U13390 (N_13390,N_11718,N_11148);
nand U13391 (N_13391,N_10081,N_10808);
nor U13392 (N_13392,N_10138,N_11158);
and U13393 (N_13393,N_11904,N_11053);
nor U13394 (N_13394,N_10176,N_11561);
xnor U13395 (N_13395,N_11102,N_10721);
xor U13396 (N_13396,N_11932,N_10394);
or U13397 (N_13397,N_11026,N_10547);
nand U13398 (N_13398,N_10660,N_10041);
nand U13399 (N_13399,N_11624,N_10530);
and U13400 (N_13400,N_10518,N_10266);
nor U13401 (N_13401,N_11783,N_11678);
and U13402 (N_13402,N_10431,N_10510);
nand U13403 (N_13403,N_11680,N_11354);
nor U13404 (N_13404,N_11135,N_11257);
and U13405 (N_13405,N_11068,N_10353);
or U13406 (N_13406,N_11501,N_11636);
and U13407 (N_13407,N_11447,N_10835);
and U13408 (N_13408,N_10346,N_10365);
or U13409 (N_13409,N_11434,N_11870);
nor U13410 (N_13410,N_11930,N_10957);
or U13411 (N_13411,N_10972,N_11973);
and U13412 (N_13412,N_10332,N_10017);
nor U13413 (N_13413,N_10361,N_11249);
nand U13414 (N_13414,N_10349,N_10069);
nand U13415 (N_13415,N_11715,N_11541);
or U13416 (N_13416,N_11023,N_11557);
nand U13417 (N_13417,N_11359,N_10406);
nor U13418 (N_13418,N_10981,N_11059);
nand U13419 (N_13419,N_10500,N_11768);
and U13420 (N_13420,N_11815,N_10515);
and U13421 (N_13421,N_10774,N_10363);
nor U13422 (N_13422,N_10158,N_11875);
nor U13423 (N_13423,N_10655,N_11399);
or U13424 (N_13424,N_11143,N_11558);
or U13425 (N_13425,N_11292,N_11780);
nor U13426 (N_13426,N_10451,N_11006);
and U13427 (N_13427,N_11700,N_10938);
or U13428 (N_13428,N_11148,N_11668);
nor U13429 (N_13429,N_11437,N_11188);
nor U13430 (N_13430,N_10829,N_11653);
nand U13431 (N_13431,N_11836,N_10050);
nor U13432 (N_13432,N_11413,N_11543);
xnor U13433 (N_13433,N_11898,N_10451);
nor U13434 (N_13434,N_10699,N_11801);
or U13435 (N_13435,N_11326,N_11509);
and U13436 (N_13436,N_10006,N_11872);
and U13437 (N_13437,N_11157,N_10902);
xnor U13438 (N_13438,N_10801,N_11523);
nand U13439 (N_13439,N_11710,N_11171);
xnor U13440 (N_13440,N_11806,N_10473);
nor U13441 (N_13441,N_10278,N_11406);
or U13442 (N_13442,N_11008,N_10177);
nand U13443 (N_13443,N_10720,N_11241);
nor U13444 (N_13444,N_10957,N_11923);
or U13445 (N_13445,N_11639,N_11082);
nor U13446 (N_13446,N_11191,N_11643);
xor U13447 (N_13447,N_10557,N_11473);
nor U13448 (N_13448,N_11279,N_11375);
nor U13449 (N_13449,N_10038,N_10434);
xor U13450 (N_13450,N_11333,N_10824);
nor U13451 (N_13451,N_11640,N_10485);
and U13452 (N_13452,N_11812,N_10645);
nand U13453 (N_13453,N_10025,N_10981);
nor U13454 (N_13454,N_11810,N_11687);
nor U13455 (N_13455,N_10081,N_11172);
or U13456 (N_13456,N_11300,N_11507);
and U13457 (N_13457,N_11360,N_10859);
nand U13458 (N_13458,N_10496,N_11663);
nand U13459 (N_13459,N_11916,N_10302);
or U13460 (N_13460,N_10016,N_10653);
and U13461 (N_13461,N_10240,N_11859);
nor U13462 (N_13462,N_11912,N_10408);
nor U13463 (N_13463,N_11371,N_11329);
and U13464 (N_13464,N_10644,N_11463);
or U13465 (N_13465,N_11770,N_10989);
and U13466 (N_13466,N_10943,N_10433);
and U13467 (N_13467,N_11544,N_11409);
and U13468 (N_13468,N_10015,N_11808);
or U13469 (N_13469,N_10898,N_11644);
nor U13470 (N_13470,N_11167,N_10874);
and U13471 (N_13471,N_10587,N_10253);
nand U13472 (N_13472,N_10108,N_10628);
and U13473 (N_13473,N_11746,N_11647);
nor U13474 (N_13474,N_11645,N_10376);
and U13475 (N_13475,N_10420,N_10806);
or U13476 (N_13476,N_11399,N_10428);
or U13477 (N_13477,N_10539,N_10988);
or U13478 (N_13478,N_11870,N_10006);
or U13479 (N_13479,N_10511,N_11249);
and U13480 (N_13480,N_10010,N_11214);
and U13481 (N_13481,N_10367,N_11286);
or U13482 (N_13482,N_10633,N_10074);
or U13483 (N_13483,N_11689,N_11570);
nand U13484 (N_13484,N_11713,N_10942);
nor U13485 (N_13485,N_10657,N_10330);
xor U13486 (N_13486,N_11072,N_10894);
nand U13487 (N_13487,N_10565,N_11810);
nand U13488 (N_13488,N_11920,N_10645);
and U13489 (N_13489,N_10012,N_11252);
xnor U13490 (N_13490,N_11135,N_10858);
and U13491 (N_13491,N_11521,N_10736);
or U13492 (N_13492,N_10892,N_11943);
or U13493 (N_13493,N_11915,N_11416);
and U13494 (N_13494,N_11945,N_11139);
xnor U13495 (N_13495,N_10156,N_11781);
and U13496 (N_13496,N_11211,N_11075);
nand U13497 (N_13497,N_11935,N_11470);
and U13498 (N_13498,N_11074,N_10293);
nand U13499 (N_13499,N_10839,N_10212);
nor U13500 (N_13500,N_10570,N_11031);
and U13501 (N_13501,N_10073,N_11438);
or U13502 (N_13502,N_11542,N_10150);
nand U13503 (N_13503,N_11198,N_10505);
and U13504 (N_13504,N_10099,N_10724);
nand U13505 (N_13505,N_11583,N_10006);
xor U13506 (N_13506,N_10399,N_11919);
and U13507 (N_13507,N_10893,N_11698);
nand U13508 (N_13508,N_10931,N_10559);
nor U13509 (N_13509,N_11701,N_11342);
and U13510 (N_13510,N_11597,N_10518);
nand U13511 (N_13511,N_11036,N_11924);
nor U13512 (N_13512,N_10772,N_11745);
nor U13513 (N_13513,N_10312,N_10793);
or U13514 (N_13514,N_10983,N_10612);
xnor U13515 (N_13515,N_11059,N_10356);
nor U13516 (N_13516,N_11909,N_10790);
or U13517 (N_13517,N_10336,N_11130);
or U13518 (N_13518,N_10221,N_10850);
or U13519 (N_13519,N_10175,N_10836);
and U13520 (N_13520,N_10647,N_10681);
nor U13521 (N_13521,N_11904,N_11934);
or U13522 (N_13522,N_11345,N_10118);
nor U13523 (N_13523,N_11262,N_10620);
nand U13524 (N_13524,N_11521,N_11223);
or U13525 (N_13525,N_11245,N_11616);
nand U13526 (N_13526,N_10950,N_11041);
and U13527 (N_13527,N_10948,N_10764);
nand U13528 (N_13528,N_11314,N_10414);
or U13529 (N_13529,N_11582,N_11877);
and U13530 (N_13530,N_10417,N_11940);
or U13531 (N_13531,N_10995,N_10104);
nand U13532 (N_13532,N_11366,N_11332);
xor U13533 (N_13533,N_11657,N_10717);
or U13534 (N_13534,N_11441,N_11592);
nand U13535 (N_13535,N_10408,N_10420);
nor U13536 (N_13536,N_10151,N_11462);
nor U13537 (N_13537,N_11519,N_11591);
nand U13538 (N_13538,N_10961,N_10270);
nand U13539 (N_13539,N_11584,N_11297);
nor U13540 (N_13540,N_11452,N_11216);
or U13541 (N_13541,N_11837,N_11072);
nand U13542 (N_13542,N_11062,N_10685);
xnor U13543 (N_13543,N_11828,N_10428);
or U13544 (N_13544,N_10906,N_10385);
nor U13545 (N_13545,N_11642,N_10767);
or U13546 (N_13546,N_11283,N_10504);
nand U13547 (N_13547,N_10360,N_10449);
and U13548 (N_13548,N_11448,N_11805);
or U13549 (N_13549,N_11621,N_10628);
nor U13550 (N_13550,N_11162,N_11748);
nand U13551 (N_13551,N_10411,N_11830);
nand U13552 (N_13552,N_11124,N_11917);
or U13553 (N_13553,N_11378,N_11564);
xor U13554 (N_13554,N_10923,N_11970);
and U13555 (N_13555,N_11670,N_10424);
nand U13556 (N_13556,N_11130,N_10512);
nor U13557 (N_13557,N_10868,N_11203);
and U13558 (N_13558,N_10539,N_10225);
and U13559 (N_13559,N_10990,N_10427);
or U13560 (N_13560,N_11622,N_10292);
or U13561 (N_13561,N_11099,N_11689);
xor U13562 (N_13562,N_11333,N_10775);
xor U13563 (N_13563,N_10946,N_11144);
nor U13564 (N_13564,N_10859,N_11831);
and U13565 (N_13565,N_11481,N_11320);
nor U13566 (N_13566,N_11913,N_10021);
or U13567 (N_13567,N_10534,N_10776);
nor U13568 (N_13568,N_11643,N_11145);
or U13569 (N_13569,N_11479,N_11941);
nand U13570 (N_13570,N_10861,N_10469);
and U13571 (N_13571,N_11750,N_11464);
nand U13572 (N_13572,N_10664,N_10149);
nand U13573 (N_13573,N_10435,N_11936);
xor U13574 (N_13574,N_11066,N_11207);
nand U13575 (N_13575,N_11113,N_11752);
nor U13576 (N_13576,N_10857,N_10416);
nor U13577 (N_13577,N_11855,N_10309);
nor U13578 (N_13578,N_10690,N_11792);
nand U13579 (N_13579,N_10576,N_11276);
or U13580 (N_13580,N_11211,N_10646);
and U13581 (N_13581,N_10830,N_11296);
and U13582 (N_13582,N_11226,N_10824);
nand U13583 (N_13583,N_11109,N_11439);
and U13584 (N_13584,N_10137,N_11476);
xor U13585 (N_13585,N_10636,N_10196);
and U13586 (N_13586,N_10536,N_10501);
nand U13587 (N_13587,N_10831,N_10073);
and U13588 (N_13588,N_10131,N_11313);
and U13589 (N_13589,N_10235,N_10438);
or U13590 (N_13590,N_10579,N_10128);
nor U13591 (N_13591,N_10857,N_11934);
nor U13592 (N_13592,N_10940,N_11041);
and U13593 (N_13593,N_10327,N_10529);
or U13594 (N_13594,N_11880,N_10482);
and U13595 (N_13595,N_11449,N_11700);
nor U13596 (N_13596,N_11667,N_11315);
and U13597 (N_13597,N_11010,N_10044);
and U13598 (N_13598,N_11941,N_11652);
nand U13599 (N_13599,N_11685,N_11208);
nor U13600 (N_13600,N_10363,N_10277);
nor U13601 (N_13601,N_11003,N_11166);
or U13602 (N_13602,N_10730,N_10241);
and U13603 (N_13603,N_10734,N_10153);
nor U13604 (N_13604,N_10499,N_10831);
nor U13605 (N_13605,N_10959,N_10220);
or U13606 (N_13606,N_10366,N_10939);
nand U13607 (N_13607,N_10925,N_10709);
nor U13608 (N_13608,N_11214,N_10847);
or U13609 (N_13609,N_11595,N_11329);
or U13610 (N_13610,N_11962,N_10772);
or U13611 (N_13611,N_11812,N_10211);
or U13612 (N_13612,N_10645,N_11981);
nor U13613 (N_13613,N_10035,N_11635);
nor U13614 (N_13614,N_10790,N_10236);
nand U13615 (N_13615,N_10591,N_10001);
or U13616 (N_13616,N_11211,N_11418);
nor U13617 (N_13617,N_11786,N_11102);
nor U13618 (N_13618,N_11598,N_11928);
nand U13619 (N_13619,N_10574,N_10247);
or U13620 (N_13620,N_10548,N_10984);
xor U13621 (N_13621,N_11317,N_10137);
and U13622 (N_13622,N_10620,N_10154);
and U13623 (N_13623,N_10384,N_11121);
or U13624 (N_13624,N_10766,N_10045);
and U13625 (N_13625,N_10937,N_10157);
or U13626 (N_13626,N_10603,N_10291);
nor U13627 (N_13627,N_11278,N_10098);
nor U13628 (N_13628,N_11589,N_11268);
nor U13629 (N_13629,N_10472,N_10479);
or U13630 (N_13630,N_11555,N_11822);
and U13631 (N_13631,N_10784,N_10800);
nor U13632 (N_13632,N_11647,N_10058);
nand U13633 (N_13633,N_11937,N_10403);
nor U13634 (N_13634,N_10648,N_10965);
nand U13635 (N_13635,N_11775,N_10371);
xor U13636 (N_13636,N_10475,N_10012);
nand U13637 (N_13637,N_10859,N_11431);
and U13638 (N_13638,N_11061,N_10229);
nor U13639 (N_13639,N_11689,N_10743);
nor U13640 (N_13640,N_10728,N_11339);
and U13641 (N_13641,N_10351,N_11946);
and U13642 (N_13642,N_11138,N_11999);
nor U13643 (N_13643,N_10193,N_10826);
nor U13644 (N_13644,N_10065,N_11372);
and U13645 (N_13645,N_11173,N_10704);
and U13646 (N_13646,N_11757,N_10047);
and U13647 (N_13647,N_10758,N_11010);
xor U13648 (N_13648,N_11560,N_11898);
nor U13649 (N_13649,N_10326,N_11795);
nor U13650 (N_13650,N_10471,N_10778);
nor U13651 (N_13651,N_10336,N_11150);
nor U13652 (N_13652,N_11433,N_11720);
and U13653 (N_13653,N_11178,N_11089);
nor U13654 (N_13654,N_11282,N_10753);
and U13655 (N_13655,N_11976,N_10478);
and U13656 (N_13656,N_10369,N_10659);
or U13657 (N_13657,N_11410,N_10782);
nand U13658 (N_13658,N_10580,N_11245);
nand U13659 (N_13659,N_11765,N_10904);
or U13660 (N_13660,N_11445,N_10563);
nand U13661 (N_13661,N_10205,N_10432);
nand U13662 (N_13662,N_11791,N_10669);
nand U13663 (N_13663,N_11444,N_10438);
and U13664 (N_13664,N_11388,N_10414);
or U13665 (N_13665,N_10073,N_10504);
nor U13666 (N_13666,N_11771,N_11723);
and U13667 (N_13667,N_11823,N_11298);
nor U13668 (N_13668,N_11979,N_11626);
nor U13669 (N_13669,N_10028,N_11354);
or U13670 (N_13670,N_10584,N_11034);
and U13671 (N_13671,N_11143,N_10827);
or U13672 (N_13672,N_10453,N_11689);
nor U13673 (N_13673,N_11477,N_11153);
or U13674 (N_13674,N_11855,N_11635);
or U13675 (N_13675,N_11004,N_11173);
and U13676 (N_13676,N_11814,N_10009);
nand U13677 (N_13677,N_10970,N_10351);
or U13678 (N_13678,N_11110,N_10008);
or U13679 (N_13679,N_11507,N_11019);
or U13680 (N_13680,N_10968,N_11691);
or U13681 (N_13681,N_10418,N_11855);
or U13682 (N_13682,N_11884,N_10691);
or U13683 (N_13683,N_11201,N_10896);
and U13684 (N_13684,N_11791,N_10745);
or U13685 (N_13685,N_10486,N_11627);
nor U13686 (N_13686,N_10389,N_11203);
or U13687 (N_13687,N_11560,N_10189);
and U13688 (N_13688,N_11695,N_10413);
or U13689 (N_13689,N_10363,N_11435);
or U13690 (N_13690,N_11467,N_11698);
nand U13691 (N_13691,N_10978,N_10672);
xnor U13692 (N_13692,N_10847,N_11075);
or U13693 (N_13693,N_10606,N_11753);
or U13694 (N_13694,N_10296,N_11366);
nand U13695 (N_13695,N_10467,N_11525);
or U13696 (N_13696,N_10780,N_11693);
nor U13697 (N_13697,N_10979,N_11560);
or U13698 (N_13698,N_11259,N_10702);
nor U13699 (N_13699,N_10468,N_11149);
and U13700 (N_13700,N_11829,N_11702);
and U13701 (N_13701,N_10438,N_11419);
nand U13702 (N_13702,N_11142,N_11895);
nand U13703 (N_13703,N_11863,N_10625);
nor U13704 (N_13704,N_11785,N_11788);
nor U13705 (N_13705,N_10019,N_11492);
and U13706 (N_13706,N_11494,N_11853);
nand U13707 (N_13707,N_11719,N_11249);
and U13708 (N_13708,N_10019,N_11965);
and U13709 (N_13709,N_10389,N_10736);
xor U13710 (N_13710,N_10947,N_11477);
or U13711 (N_13711,N_10205,N_11478);
or U13712 (N_13712,N_10516,N_10423);
and U13713 (N_13713,N_10420,N_10202);
or U13714 (N_13714,N_11719,N_11113);
nor U13715 (N_13715,N_11718,N_11772);
and U13716 (N_13716,N_11893,N_10423);
nor U13717 (N_13717,N_10115,N_10863);
nor U13718 (N_13718,N_11920,N_11140);
and U13719 (N_13719,N_11029,N_10979);
or U13720 (N_13720,N_10111,N_10822);
and U13721 (N_13721,N_10550,N_11221);
nand U13722 (N_13722,N_10574,N_11014);
or U13723 (N_13723,N_11293,N_11699);
nand U13724 (N_13724,N_11191,N_11739);
and U13725 (N_13725,N_10830,N_11192);
and U13726 (N_13726,N_10831,N_11078);
nand U13727 (N_13727,N_10985,N_10007);
or U13728 (N_13728,N_11882,N_10083);
or U13729 (N_13729,N_11325,N_10220);
or U13730 (N_13730,N_11551,N_10544);
or U13731 (N_13731,N_11938,N_10821);
nor U13732 (N_13732,N_10991,N_10288);
nand U13733 (N_13733,N_11843,N_11882);
nor U13734 (N_13734,N_10520,N_11217);
and U13735 (N_13735,N_10937,N_10480);
and U13736 (N_13736,N_11458,N_10779);
or U13737 (N_13737,N_10797,N_11951);
and U13738 (N_13738,N_11830,N_10624);
nor U13739 (N_13739,N_10947,N_10137);
nor U13740 (N_13740,N_10899,N_10529);
nand U13741 (N_13741,N_11496,N_10813);
and U13742 (N_13742,N_11915,N_11872);
nor U13743 (N_13743,N_11589,N_10178);
nand U13744 (N_13744,N_10996,N_10232);
nand U13745 (N_13745,N_10426,N_11001);
or U13746 (N_13746,N_11446,N_11997);
nor U13747 (N_13747,N_10876,N_10626);
and U13748 (N_13748,N_10714,N_11574);
or U13749 (N_13749,N_10434,N_10617);
and U13750 (N_13750,N_10028,N_11649);
nand U13751 (N_13751,N_11190,N_11708);
nor U13752 (N_13752,N_11125,N_10633);
and U13753 (N_13753,N_10619,N_11177);
nand U13754 (N_13754,N_10492,N_10959);
nand U13755 (N_13755,N_11108,N_11971);
nand U13756 (N_13756,N_10061,N_10998);
xor U13757 (N_13757,N_11277,N_10869);
nand U13758 (N_13758,N_10708,N_11475);
or U13759 (N_13759,N_10663,N_11797);
nor U13760 (N_13760,N_10976,N_10058);
nor U13761 (N_13761,N_10642,N_10751);
xnor U13762 (N_13762,N_10184,N_10781);
and U13763 (N_13763,N_11305,N_10612);
or U13764 (N_13764,N_10608,N_11565);
or U13765 (N_13765,N_11349,N_10630);
xnor U13766 (N_13766,N_10294,N_10095);
nand U13767 (N_13767,N_10362,N_11868);
nand U13768 (N_13768,N_10172,N_11474);
nand U13769 (N_13769,N_10696,N_11082);
or U13770 (N_13770,N_10198,N_11587);
nor U13771 (N_13771,N_10976,N_10695);
or U13772 (N_13772,N_11376,N_11479);
or U13773 (N_13773,N_11230,N_11568);
nor U13774 (N_13774,N_11625,N_10195);
nand U13775 (N_13775,N_10716,N_11679);
and U13776 (N_13776,N_10645,N_10793);
nor U13777 (N_13777,N_11475,N_10391);
and U13778 (N_13778,N_10527,N_10396);
or U13779 (N_13779,N_11367,N_11040);
nor U13780 (N_13780,N_11442,N_10762);
nor U13781 (N_13781,N_11420,N_11780);
nor U13782 (N_13782,N_10111,N_10776);
nor U13783 (N_13783,N_10993,N_10500);
nor U13784 (N_13784,N_11704,N_11137);
xor U13785 (N_13785,N_10484,N_10513);
nand U13786 (N_13786,N_11378,N_10372);
and U13787 (N_13787,N_10493,N_11635);
or U13788 (N_13788,N_10425,N_10818);
nand U13789 (N_13789,N_10902,N_10489);
or U13790 (N_13790,N_11572,N_11273);
nand U13791 (N_13791,N_10052,N_11180);
nor U13792 (N_13792,N_11419,N_11528);
or U13793 (N_13793,N_10734,N_10454);
or U13794 (N_13794,N_10976,N_11504);
nor U13795 (N_13795,N_11848,N_10592);
nand U13796 (N_13796,N_11226,N_10183);
nand U13797 (N_13797,N_10519,N_11786);
or U13798 (N_13798,N_11701,N_10509);
xor U13799 (N_13799,N_10539,N_11786);
nor U13800 (N_13800,N_10454,N_11081);
nor U13801 (N_13801,N_11906,N_11440);
and U13802 (N_13802,N_10625,N_10233);
nand U13803 (N_13803,N_10835,N_10647);
nor U13804 (N_13804,N_10956,N_10171);
or U13805 (N_13805,N_10710,N_10062);
or U13806 (N_13806,N_10354,N_11526);
nand U13807 (N_13807,N_10813,N_10038);
and U13808 (N_13808,N_10946,N_11696);
and U13809 (N_13809,N_10750,N_10878);
nand U13810 (N_13810,N_10311,N_11416);
or U13811 (N_13811,N_10805,N_11750);
nand U13812 (N_13812,N_11044,N_10050);
nand U13813 (N_13813,N_10159,N_10815);
and U13814 (N_13814,N_11990,N_10389);
and U13815 (N_13815,N_11179,N_10106);
nand U13816 (N_13816,N_11931,N_11085);
and U13817 (N_13817,N_10856,N_11399);
or U13818 (N_13818,N_11402,N_10213);
nand U13819 (N_13819,N_10194,N_11391);
nor U13820 (N_13820,N_10232,N_10222);
nor U13821 (N_13821,N_11881,N_11267);
xnor U13822 (N_13822,N_11631,N_10607);
nor U13823 (N_13823,N_10836,N_11738);
xnor U13824 (N_13824,N_11948,N_10153);
and U13825 (N_13825,N_10157,N_11319);
or U13826 (N_13826,N_11975,N_11197);
xor U13827 (N_13827,N_10169,N_10667);
and U13828 (N_13828,N_10859,N_11456);
nor U13829 (N_13829,N_11592,N_11000);
xor U13830 (N_13830,N_10244,N_11593);
nor U13831 (N_13831,N_10906,N_11754);
or U13832 (N_13832,N_10017,N_11149);
nor U13833 (N_13833,N_11812,N_10608);
or U13834 (N_13834,N_10074,N_11647);
xor U13835 (N_13835,N_10628,N_10830);
nand U13836 (N_13836,N_11935,N_10142);
or U13837 (N_13837,N_11699,N_10345);
or U13838 (N_13838,N_11407,N_11785);
and U13839 (N_13839,N_10305,N_10355);
xor U13840 (N_13840,N_11761,N_11913);
nand U13841 (N_13841,N_11248,N_11906);
nor U13842 (N_13842,N_11710,N_10587);
or U13843 (N_13843,N_10124,N_10165);
nand U13844 (N_13844,N_11492,N_10975);
or U13845 (N_13845,N_11747,N_11980);
nor U13846 (N_13846,N_11780,N_10101);
and U13847 (N_13847,N_10359,N_10695);
or U13848 (N_13848,N_11071,N_11847);
nor U13849 (N_13849,N_10122,N_10873);
nor U13850 (N_13850,N_11228,N_11809);
and U13851 (N_13851,N_10313,N_11193);
nor U13852 (N_13852,N_11077,N_10590);
xor U13853 (N_13853,N_11450,N_11265);
nor U13854 (N_13854,N_11275,N_10861);
and U13855 (N_13855,N_11162,N_10433);
nor U13856 (N_13856,N_10962,N_10336);
nor U13857 (N_13857,N_11870,N_10555);
and U13858 (N_13858,N_10441,N_11419);
nand U13859 (N_13859,N_11987,N_10028);
and U13860 (N_13860,N_11127,N_10790);
and U13861 (N_13861,N_10208,N_10296);
nor U13862 (N_13862,N_11892,N_10241);
nor U13863 (N_13863,N_10713,N_11485);
or U13864 (N_13864,N_11320,N_11814);
nand U13865 (N_13865,N_10137,N_10665);
and U13866 (N_13866,N_10638,N_11817);
or U13867 (N_13867,N_11580,N_10485);
xor U13868 (N_13868,N_10322,N_10614);
nand U13869 (N_13869,N_10184,N_11311);
nand U13870 (N_13870,N_10526,N_10581);
and U13871 (N_13871,N_10475,N_10252);
nor U13872 (N_13872,N_11426,N_10709);
nor U13873 (N_13873,N_11251,N_11970);
or U13874 (N_13874,N_11276,N_11680);
or U13875 (N_13875,N_10193,N_10922);
nor U13876 (N_13876,N_10438,N_10071);
nor U13877 (N_13877,N_11794,N_10898);
nand U13878 (N_13878,N_11222,N_10524);
nor U13879 (N_13879,N_11089,N_10074);
nor U13880 (N_13880,N_11835,N_10660);
and U13881 (N_13881,N_11858,N_11126);
and U13882 (N_13882,N_10761,N_10675);
xor U13883 (N_13883,N_11696,N_10544);
or U13884 (N_13884,N_11886,N_11109);
nand U13885 (N_13885,N_11380,N_11932);
or U13886 (N_13886,N_10791,N_10214);
nor U13887 (N_13887,N_10541,N_11909);
or U13888 (N_13888,N_10669,N_10203);
nor U13889 (N_13889,N_10622,N_10012);
or U13890 (N_13890,N_10584,N_10860);
nand U13891 (N_13891,N_11448,N_10388);
or U13892 (N_13892,N_10031,N_10857);
nor U13893 (N_13893,N_11491,N_10000);
xor U13894 (N_13894,N_10533,N_11137);
xor U13895 (N_13895,N_10286,N_11820);
nor U13896 (N_13896,N_10089,N_11752);
nor U13897 (N_13897,N_10327,N_10924);
nand U13898 (N_13898,N_10488,N_11277);
or U13899 (N_13899,N_10184,N_11901);
or U13900 (N_13900,N_11872,N_10883);
nand U13901 (N_13901,N_10238,N_10984);
or U13902 (N_13902,N_10420,N_10590);
nor U13903 (N_13903,N_11688,N_10782);
and U13904 (N_13904,N_11764,N_11902);
or U13905 (N_13905,N_10493,N_11050);
nor U13906 (N_13906,N_11566,N_10269);
or U13907 (N_13907,N_11884,N_11111);
and U13908 (N_13908,N_10679,N_10749);
and U13909 (N_13909,N_11330,N_11791);
nor U13910 (N_13910,N_10124,N_10297);
or U13911 (N_13911,N_11841,N_10207);
nor U13912 (N_13912,N_11337,N_11895);
and U13913 (N_13913,N_10758,N_11297);
xnor U13914 (N_13914,N_10842,N_10748);
nor U13915 (N_13915,N_10748,N_10847);
and U13916 (N_13916,N_10916,N_11736);
and U13917 (N_13917,N_11655,N_11790);
nor U13918 (N_13918,N_11272,N_10691);
nand U13919 (N_13919,N_11282,N_11768);
nor U13920 (N_13920,N_10589,N_11691);
or U13921 (N_13921,N_10200,N_11934);
nand U13922 (N_13922,N_11501,N_10932);
and U13923 (N_13923,N_10285,N_11564);
and U13924 (N_13924,N_10898,N_11400);
nor U13925 (N_13925,N_11212,N_11508);
nand U13926 (N_13926,N_10182,N_11929);
and U13927 (N_13927,N_10423,N_11195);
nand U13928 (N_13928,N_10919,N_11018);
and U13929 (N_13929,N_10780,N_10729);
xor U13930 (N_13930,N_10086,N_11076);
nor U13931 (N_13931,N_11456,N_10594);
or U13932 (N_13932,N_10735,N_10059);
or U13933 (N_13933,N_10275,N_11993);
nor U13934 (N_13934,N_11281,N_10557);
and U13935 (N_13935,N_10828,N_10825);
and U13936 (N_13936,N_10119,N_10175);
or U13937 (N_13937,N_10556,N_10655);
and U13938 (N_13938,N_11922,N_10358);
nor U13939 (N_13939,N_11050,N_10826);
nand U13940 (N_13940,N_10057,N_10049);
and U13941 (N_13941,N_10911,N_10676);
and U13942 (N_13942,N_11296,N_11628);
xnor U13943 (N_13943,N_10511,N_10680);
nor U13944 (N_13944,N_10520,N_11906);
or U13945 (N_13945,N_11358,N_11355);
or U13946 (N_13946,N_10228,N_10049);
nand U13947 (N_13947,N_10222,N_11677);
or U13948 (N_13948,N_10797,N_10912);
or U13949 (N_13949,N_10868,N_10783);
and U13950 (N_13950,N_10676,N_10463);
xnor U13951 (N_13951,N_11286,N_11936);
nand U13952 (N_13952,N_11668,N_11916);
or U13953 (N_13953,N_10025,N_11540);
xor U13954 (N_13954,N_11911,N_11734);
nor U13955 (N_13955,N_10073,N_11764);
nand U13956 (N_13956,N_11676,N_10463);
and U13957 (N_13957,N_11447,N_11725);
or U13958 (N_13958,N_10593,N_11668);
or U13959 (N_13959,N_11008,N_10564);
nand U13960 (N_13960,N_11365,N_10640);
nor U13961 (N_13961,N_10072,N_11951);
nand U13962 (N_13962,N_11419,N_10775);
nor U13963 (N_13963,N_10291,N_10354);
and U13964 (N_13964,N_11860,N_11421);
nor U13965 (N_13965,N_11206,N_10067);
or U13966 (N_13966,N_10492,N_11258);
nor U13967 (N_13967,N_10078,N_10357);
nor U13968 (N_13968,N_10423,N_11095);
and U13969 (N_13969,N_11389,N_11925);
nand U13970 (N_13970,N_11660,N_10230);
nor U13971 (N_13971,N_10877,N_11306);
nand U13972 (N_13972,N_10684,N_11766);
or U13973 (N_13973,N_11407,N_11960);
nand U13974 (N_13974,N_11223,N_10005);
nand U13975 (N_13975,N_11985,N_10813);
nand U13976 (N_13976,N_10259,N_10569);
or U13977 (N_13977,N_10746,N_10792);
nor U13978 (N_13978,N_11936,N_11677);
nand U13979 (N_13979,N_10950,N_11440);
and U13980 (N_13980,N_10981,N_10634);
xor U13981 (N_13981,N_11298,N_10207);
nand U13982 (N_13982,N_10828,N_10354);
nor U13983 (N_13983,N_10259,N_10581);
and U13984 (N_13984,N_10989,N_10657);
nand U13985 (N_13985,N_10239,N_11272);
nor U13986 (N_13986,N_11500,N_10118);
nor U13987 (N_13987,N_10978,N_10902);
nor U13988 (N_13988,N_11633,N_10500);
nand U13989 (N_13989,N_10664,N_10728);
nor U13990 (N_13990,N_11554,N_10146);
and U13991 (N_13991,N_10474,N_11511);
or U13992 (N_13992,N_10509,N_11924);
or U13993 (N_13993,N_11125,N_10881);
nand U13994 (N_13994,N_10358,N_11032);
and U13995 (N_13995,N_11091,N_10884);
nor U13996 (N_13996,N_10769,N_11312);
and U13997 (N_13997,N_11916,N_11535);
and U13998 (N_13998,N_11041,N_10714);
nor U13999 (N_13999,N_10570,N_10074);
nand U14000 (N_14000,N_13968,N_12510);
and U14001 (N_14001,N_12044,N_12597);
nand U14002 (N_14002,N_13352,N_13676);
nor U14003 (N_14003,N_12015,N_12012);
nand U14004 (N_14004,N_13430,N_13511);
xnor U14005 (N_14005,N_13632,N_12698);
and U14006 (N_14006,N_13603,N_13645);
xor U14007 (N_14007,N_12455,N_12789);
and U14008 (N_14008,N_12134,N_12443);
nand U14009 (N_14009,N_12096,N_13719);
nand U14010 (N_14010,N_13784,N_12562);
and U14011 (N_14011,N_13677,N_13131);
nand U14012 (N_14012,N_13786,N_12231);
nand U14013 (N_14013,N_12953,N_13366);
and U14014 (N_14014,N_12552,N_13897);
or U14015 (N_14015,N_13622,N_12794);
nor U14016 (N_14016,N_12971,N_13429);
nand U14017 (N_14017,N_13130,N_13240);
nor U14018 (N_14018,N_13295,N_13580);
or U14019 (N_14019,N_12501,N_13926);
nor U14020 (N_14020,N_13656,N_12200);
nor U14021 (N_14021,N_12331,N_13783);
and U14022 (N_14022,N_12996,N_13252);
or U14023 (N_14023,N_13762,N_12683);
and U14024 (N_14024,N_12762,N_12380);
or U14025 (N_14025,N_13041,N_12082);
nand U14026 (N_14026,N_12129,N_13170);
nor U14027 (N_14027,N_13161,N_12578);
xnor U14028 (N_14028,N_12214,N_13198);
nor U14029 (N_14029,N_13563,N_13909);
nand U14030 (N_14030,N_12828,N_13433);
nand U14031 (N_14031,N_13700,N_13290);
nor U14032 (N_14032,N_13848,N_12041);
nor U14033 (N_14033,N_13435,N_13886);
and U14034 (N_14034,N_12737,N_12717);
and U14035 (N_14035,N_13687,N_13851);
nor U14036 (N_14036,N_12132,N_12829);
or U14037 (N_14037,N_12963,N_12230);
xnor U14038 (N_14038,N_13036,N_13809);
and U14039 (N_14039,N_12368,N_13098);
and U14040 (N_14040,N_13401,N_13501);
nand U14041 (N_14041,N_13265,N_12427);
xnor U14042 (N_14042,N_13094,N_12805);
nor U14043 (N_14043,N_13031,N_13110);
and U14044 (N_14044,N_13797,N_12263);
and U14045 (N_14045,N_13086,N_12732);
and U14046 (N_14046,N_12258,N_12574);
or U14047 (N_14047,N_13468,N_13473);
xnor U14048 (N_14048,N_13422,N_12018);
and U14049 (N_14049,N_13074,N_12111);
nand U14050 (N_14050,N_12915,N_13947);
nand U14051 (N_14051,N_12716,N_12268);
or U14052 (N_14052,N_12658,N_12685);
and U14053 (N_14053,N_12172,N_12912);
nand U14054 (N_14054,N_12988,N_12186);
nor U14055 (N_14055,N_13724,N_12809);
and U14056 (N_14056,N_13770,N_13698);
nand U14057 (N_14057,N_13141,N_12959);
and U14058 (N_14058,N_12367,N_12130);
xor U14059 (N_14059,N_13489,N_12792);
or U14060 (N_14060,N_13906,N_13843);
or U14061 (N_14061,N_13990,N_12588);
xnor U14062 (N_14062,N_12495,N_13027);
nor U14063 (N_14063,N_13158,N_13377);
nand U14064 (N_14064,N_12487,N_12972);
nand U14065 (N_14065,N_12317,N_13369);
and U14066 (N_14066,N_13930,N_12970);
nand U14067 (N_14067,N_13046,N_13210);
xnor U14068 (N_14068,N_12902,N_12749);
and U14069 (N_14069,N_12766,N_12121);
and U14070 (N_14070,N_12690,N_12341);
or U14071 (N_14071,N_13703,N_13938);
xnor U14072 (N_14072,N_13845,N_12124);
or U14073 (N_14073,N_13218,N_12918);
or U14074 (N_14074,N_12948,N_13075);
and U14075 (N_14075,N_12118,N_13072);
and U14076 (N_14076,N_13514,N_13313);
and U14077 (N_14077,N_12070,N_12465);
xnor U14078 (N_14078,N_13597,N_12378);
xor U14079 (N_14079,N_13873,N_12966);
and U14080 (N_14080,N_12093,N_12120);
nand U14081 (N_14081,N_13949,N_12933);
or U14082 (N_14082,N_12307,N_12763);
or U14083 (N_14083,N_13494,N_12225);
and U14084 (N_14084,N_12114,N_13378);
or U14085 (N_14085,N_12822,N_12257);
or U14086 (N_14086,N_13385,N_13693);
and U14087 (N_14087,N_13876,N_13100);
nand U14088 (N_14088,N_13894,N_13806);
xor U14089 (N_14089,N_12951,N_13414);
nor U14090 (N_14090,N_12435,N_12388);
and U14091 (N_14091,N_12632,N_12899);
nand U14092 (N_14092,N_13858,N_13743);
or U14093 (N_14093,N_12934,N_12603);
xnor U14094 (N_14094,N_12808,N_13436);
nor U14095 (N_14095,N_13208,N_13345);
or U14096 (N_14096,N_12224,N_12719);
nor U14097 (N_14097,N_13291,N_13531);
and U14098 (N_14098,N_12025,N_12653);
xor U14099 (N_14099,N_12589,N_12673);
or U14100 (N_14100,N_12538,N_12638);
xnor U14101 (N_14101,N_13870,N_12384);
or U14102 (N_14102,N_12927,N_13266);
and U14103 (N_14103,N_12035,N_13201);
or U14104 (N_14104,N_12941,N_13179);
nor U14105 (N_14105,N_12804,N_13103);
or U14106 (N_14106,N_13277,N_13140);
and U14107 (N_14107,N_13661,N_13000);
and U14108 (N_14108,N_13504,N_12730);
nand U14109 (N_14109,N_13863,N_12739);
nand U14110 (N_14110,N_12206,N_12101);
xnor U14111 (N_14111,N_13944,N_13912);
or U14112 (N_14112,N_12440,N_13317);
nor U14113 (N_14113,N_13936,N_13620);
xnor U14114 (N_14114,N_12919,N_12875);
and U14115 (N_14115,N_13409,N_12004);
xnor U14116 (N_14116,N_13890,N_12848);
and U14117 (N_14117,N_12277,N_13296);
nand U14118 (N_14118,N_13079,N_13398);
nor U14119 (N_14119,N_12831,N_13776);
or U14120 (N_14120,N_13824,N_13424);
nor U14121 (N_14121,N_12300,N_13801);
or U14122 (N_14122,N_13678,N_12994);
xor U14123 (N_14123,N_13482,N_13005);
xnor U14124 (N_14124,N_13852,N_13297);
nor U14125 (N_14125,N_13380,N_12938);
nor U14126 (N_14126,N_12787,N_12895);
and U14127 (N_14127,N_12855,N_13310);
nand U14128 (N_14128,N_13284,N_13556);
nor U14129 (N_14129,N_13411,N_12974);
and U14130 (N_14130,N_13211,N_12256);
and U14131 (N_14131,N_12131,N_13749);
nor U14132 (N_14132,N_12694,N_13988);
and U14133 (N_14133,N_13443,N_13434);
or U14134 (N_14134,N_12480,N_13121);
and U14135 (N_14135,N_13815,N_13490);
nand U14136 (N_14136,N_12901,N_13878);
nand U14137 (N_14137,N_13042,N_13493);
and U14138 (N_14138,N_13097,N_12677);
nor U14139 (N_14139,N_13465,N_12850);
and U14140 (N_14140,N_13530,N_13623);
or U14141 (N_14141,N_13523,N_12626);
or U14142 (N_14142,N_13426,N_12086);
and U14143 (N_14143,N_12336,N_13219);
nand U14144 (N_14144,N_12464,N_13699);
nand U14145 (N_14145,N_12356,N_13197);
nand U14146 (N_14146,N_12823,N_12873);
nand U14147 (N_14147,N_12610,N_13246);
or U14148 (N_14148,N_13119,N_12079);
xnor U14149 (N_14149,N_13101,N_12784);
or U14150 (N_14150,N_12559,N_12339);
and U14151 (N_14151,N_13125,N_13441);
and U14152 (N_14152,N_12293,N_13250);
and U14153 (N_14153,N_13710,N_12398);
nor U14154 (N_14154,N_13903,N_13194);
and U14155 (N_14155,N_13804,N_13127);
xor U14156 (N_14156,N_13063,N_12611);
nand U14157 (N_14157,N_13518,N_13664);
or U14158 (N_14158,N_13541,N_12409);
or U14159 (N_14159,N_12984,N_13136);
or U14160 (N_14160,N_13451,N_12387);
nor U14161 (N_14161,N_12615,N_12568);
xor U14162 (N_14162,N_12886,N_12904);
nor U14163 (N_14163,N_13639,N_12099);
or U14164 (N_14164,N_13823,N_13457);
and U14165 (N_14165,N_13108,N_12459);
or U14166 (N_14166,N_12773,N_12279);
nor U14167 (N_14167,N_12602,N_12081);
and U14168 (N_14168,N_13633,N_12014);
nor U14169 (N_14169,N_13260,N_12456);
and U14170 (N_14170,N_13383,N_13793);
or U14171 (N_14171,N_12976,N_13662);
or U14172 (N_14172,N_12532,N_13343);
nand U14173 (N_14173,N_12830,N_13498);
nor U14174 (N_14174,N_13545,N_12500);
and U14175 (N_14175,N_12067,N_12570);
xor U14176 (N_14176,N_12511,N_13828);
or U14177 (N_14177,N_12010,N_12365);
or U14178 (N_14178,N_13006,N_12229);
nor U14179 (N_14179,N_12373,N_13358);
or U14180 (N_14180,N_12674,N_13495);
and U14181 (N_14181,N_13860,N_12346);
or U14182 (N_14182,N_12797,N_13571);
and U14183 (N_14183,N_13855,N_13500);
and U14184 (N_14184,N_13593,N_13765);
and U14185 (N_14185,N_13740,N_12803);
nor U14186 (N_14186,N_12165,N_13900);
nor U14187 (N_14187,N_12546,N_12745);
nand U14188 (N_14188,N_12747,N_13535);
nand U14189 (N_14189,N_12858,N_13348);
or U14190 (N_14190,N_12502,N_12059);
or U14191 (N_14191,N_12275,N_13483);
or U14192 (N_14192,N_12340,N_13349);
nand U14193 (N_14193,N_12844,N_13373);
and U14194 (N_14194,N_13285,N_12218);
nor U14195 (N_14195,N_13355,N_12354);
and U14196 (N_14196,N_13774,N_13539);
xor U14197 (N_14197,N_12498,N_12494);
xnor U14198 (N_14198,N_12631,N_12003);
or U14199 (N_14199,N_13235,N_12028);
xnor U14200 (N_14200,N_13918,N_12452);
or U14201 (N_14201,N_12176,N_12980);
or U14202 (N_14202,N_12859,N_13242);
or U14203 (N_14203,N_13399,N_13659);
nor U14204 (N_14204,N_12285,N_13200);
nor U14205 (N_14205,N_12879,N_12355);
and U14206 (N_14206,N_12592,N_12343);
nand U14207 (N_14207,N_13095,N_13487);
and U14208 (N_14208,N_13566,N_13096);
nor U14209 (N_14209,N_13302,N_12347);
or U14210 (N_14210,N_13526,N_13512);
xnor U14211 (N_14211,N_13185,N_13665);
nor U14212 (N_14212,N_13604,N_12178);
nor U14213 (N_14213,N_13346,N_13163);
or U14214 (N_14214,N_13013,N_12376);
and U14215 (N_14215,N_13969,N_12672);
nand U14216 (N_14216,N_12519,N_12290);
or U14217 (N_14217,N_13800,N_13068);
nor U14218 (N_14218,N_12509,N_12119);
and U14219 (N_14219,N_13596,N_13139);
or U14220 (N_14220,N_13552,N_13789);
nand U14221 (N_14221,N_12900,N_12743);
nand U14222 (N_14222,N_13206,N_12315);
nor U14223 (N_14223,N_12585,N_12168);
and U14224 (N_14224,N_13084,N_13371);
and U14225 (N_14225,N_12582,N_12961);
nor U14226 (N_14226,N_12320,N_12103);
and U14227 (N_14227,N_13015,N_12163);
and U14228 (N_14228,N_13022,N_13254);
nor U14229 (N_14229,N_12945,N_12314);
nand U14230 (N_14230,N_13821,N_12188);
or U14231 (N_14231,N_13256,N_13697);
nand U14232 (N_14232,N_12906,N_13802);
nand U14233 (N_14233,N_12995,N_12389);
nor U14234 (N_14234,N_12569,N_12817);
nor U14235 (N_14235,N_13421,N_13683);
xnor U14236 (N_14236,N_12669,N_12874);
and U14237 (N_14237,N_12397,N_13636);
and U14238 (N_14238,N_12319,N_13869);
nand U14239 (N_14239,N_12105,N_13347);
nor U14240 (N_14240,N_12598,N_12782);
nand U14241 (N_14241,N_12201,N_12534);
or U14242 (N_14242,N_12425,N_12125);
xor U14243 (N_14243,N_12063,N_12508);
nand U14244 (N_14244,N_12174,N_13745);
xor U14245 (N_14245,N_12728,N_13372);
and U14246 (N_14246,N_13065,N_12246);
or U14247 (N_14247,N_12066,N_13638);
or U14248 (N_14248,N_12418,N_13548);
and U14249 (N_14249,N_13502,N_12783);
nor U14250 (N_14250,N_13334,N_13415);
nor U14251 (N_14251,N_13390,N_13294);
and U14252 (N_14252,N_13230,N_13055);
and U14253 (N_14253,N_12234,N_12662);
nor U14254 (N_14254,N_13054,N_12775);
nor U14255 (N_14255,N_13048,N_12548);
or U14256 (N_14256,N_12964,N_12338);
nand U14257 (N_14257,N_13157,N_12575);
and U14258 (N_14258,N_12090,N_13222);
or U14259 (N_14259,N_13529,N_12838);
nand U14260 (N_14260,N_12818,N_13680);
and U14261 (N_14261,N_13268,N_13064);
or U14262 (N_14262,N_13914,N_12055);
nand U14263 (N_14263,N_12664,N_13744);
nor U14264 (N_14264,N_13016,N_13247);
nor U14265 (N_14265,N_12451,N_13367);
or U14266 (N_14266,N_13035,N_13961);
and U14267 (N_14267,N_13326,N_12753);
nand U14268 (N_14268,N_12390,N_12344);
and U14269 (N_14269,N_12239,N_12057);
or U14270 (N_14270,N_13842,N_13261);
and U14271 (N_14271,N_12944,N_13951);
or U14272 (N_14272,N_13788,N_13520);
and U14273 (N_14273,N_13787,N_12557);
nand U14274 (N_14274,N_12637,N_12852);
or U14275 (N_14275,N_13365,N_12386);
xor U14276 (N_14276,N_12774,N_12840);
or U14277 (N_14277,N_13544,N_13572);
nand U14278 (N_14278,N_13827,N_13389);
nand U14279 (N_14279,N_12065,N_13833);
or U14280 (N_14280,N_13454,N_13599);
and U14281 (N_14281,N_12470,N_12499);
and U14282 (N_14282,N_13085,N_13558);
nand U14283 (N_14283,N_13922,N_13705);
and U14284 (N_14284,N_13905,N_13503);
nand U14285 (N_14285,N_13216,N_12094);
xnor U14286 (N_14286,N_12890,N_12713);
nor U14287 (N_14287,N_13120,N_13713);
and U14288 (N_14288,N_13980,N_13318);
nand U14289 (N_14289,N_13109,N_12005);
nand U14290 (N_14290,N_12872,N_12930);
and U14291 (N_14291,N_12553,N_13152);
nor U14292 (N_14292,N_13182,N_13621);
nor U14293 (N_14293,N_13350,N_12238);
nand U14294 (N_14294,N_12244,N_12267);
or U14295 (N_14295,N_12671,N_12247);
nor U14296 (N_14296,N_12997,N_13610);
nor U14297 (N_14297,N_13816,N_12146);
nand U14298 (N_14298,N_12466,N_12411);
nand U14299 (N_14299,N_13320,N_12522);
xnor U14300 (N_14300,N_12143,N_13278);
nor U14301 (N_14301,N_12987,N_12030);
and U14302 (N_14302,N_13183,N_12967);
and U14303 (N_14303,N_13173,N_12929);
and U14304 (N_14304,N_12271,N_12064);
nor U14305 (N_14305,N_13073,N_13416);
nor U14306 (N_14306,N_13344,N_13273);
and U14307 (N_14307,N_13581,N_13998);
nand U14308 (N_14308,N_12819,N_13887);
or U14309 (N_14309,N_13506,N_12740);
or U14310 (N_14310,N_12469,N_12196);
and U14311 (N_14311,N_12911,N_12250);
nor U14312 (N_14312,N_13463,N_12265);
xor U14313 (N_14313,N_12240,N_12222);
and U14314 (N_14314,N_12642,N_13213);
and U14315 (N_14315,N_12017,N_13226);
or U14316 (N_14316,N_13329,N_12609);
nand U14317 (N_14317,N_13948,N_12863);
xnor U14318 (N_14318,N_13805,N_12540);
nand U14319 (N_14319,N_13467,N_12092);
xnor U14320 (N_14320,N_13137,N_13650);
nand U14321 (N_14321,N_12123,N_13631);
nor U14322 (N_14322,N_13117,N_12601);
nor U14323 (N_14323,N_12416,N_12357);
nand U14324 (N_14324,N_13929,N_13898);
nor U14325 (N_14325,N_12233,N_12350);
or U14326 (N_14326,N_13047,N_13794);
and U14327 (N_14327,N_12791,N_13715);
nor U14328 (N_14328,N_12462,N_12243);
nand U14329 (N_14329,N_12016,N_12490);
or U14330 (N_14330,N_12019,N_13202);
or U14331 (N_14331,N_13111,N_13524);
and U14332 (N_14332,N_12274,N_12479);
nor U14333 (N_14333,N_12164,N_12920);
nand U14334 (N_14334,N_13464,N_13673);
and U14335 (N_14335,N_12549,N_13123);
nand U14336 (N_14336,N_12441,N_13505);
or U14337 (N_14337,N_12968,N_13831);
or U14338 (N_14338,N_13830,N_13128);
or U14339 (N_14339,N_13475,N_12680);
nand U14340 (N_14340,N_12748,N_12359);
and U14341 (N_14341,N_13287,N_12369);
nand U14342 (N_14342,N_13655,N_13420);
nor U14343 (N_14343,N_12000,N_12781);
or U14344 (N_14344,N_12696,N_12554);
and U14345 (N_14345,N_12910,N_13303);
or U14346 (N_14346,N_13839,N_12613);
xnor U14347 (N_14347,N_12193,N_13485);
nand U14348 (N_14348,N_12983,N_13327);
nand U14349 (N_14349,N_12663,N_12986);
nor U14350 (N_14350,N_13062,N_13736);
or U14351 (N_14351,N_13452,N_13193);
and U14352 (N_14352,N_12034,N_12127);
and U14353 (N_14353,N_13993,N_12727);
or U14354 (N_14354,N_13895,N_12604);
nor U14355 (N_14355,N_13153,N_12181);
and U14356 (N_14356,N_13053,N_12507);
xor U14357 (N_14357,N_13089,N_12112);
nand U14358 (N_14358,N_12699,N_12149);
nor U14359 (N_14359,N_13057,N_13986);
or U14360 (N_14360,N_12042,N_13133);
nand U14361 (N_14361,N_13829,N_13799);
nor U14362 (N_14362,N_13322,N_13649);
xnor U14363 (N_14363,N_12083,N_12687);
or U14364 (N_14364,N_13160,N_12447);
and U14365 (N_14365,N_12682,N_13551);
or U14366 (N_14366,N_13281,N_12741);
nor U14367 (N_14367,N_12001,N_12349);
and U14368 (N_14368,N_12029,N_12932);
nand U14369 (N_14369,N_13381,N_13722);
nand U14370 (N_14370,N_13825,N_12755);
nand U14371 (N_14371,N_12241,N_12142);
nor U14372 (N_14372,N_13576,N_12162);
nor U14373 (N_14373,N_13204,N_13374);
nor U14374 (N_14374,N_13155,N_12558);
nand U14375 (N_14375,N_12614,N_13438);
nor U14376 (N_14376,N_13975,N_12478);
or U14377 (N_14377,N_12391,N_12923);
or U14378 (N_14378,N_12882,N_13835);
nand U14379 (N_14379,N_13614,N_13868);
nand U14380 (N_14380,N_12047,N_13889);
or U14381 (N_14381,N_13413,N_13175);
nor U14382 (N_14382,N_12095,N_12516);
xnor U14383 (N_14383,N_12584,N_13407);
nor U14384 (N_14384,N_13654,N_13682);
nand U14385 (N_14385,N_13923,N_12991);
and U14386 (N_14386,N_13049,N_12109);
nand U14387 (N_14387,N_12720,N_13461);
or U14388 (N_14388,N_13203,N_13718);
nor U14389 (N_14389,N_12463,N_13024);
or U14390 (N_14390,N_12395,N_12217);
nand U14391 (N_14391,N_12723,N_12272);
or U14392 (N_14392,N_12657,N_12659);
or U14393 (N_14393,N_12641,N_12264);
and U14394 (N_14394,N_13814,N_12969);
xor U14395 (N_14395,N_13028,N_13856);
nor U14396 (N_14396,N_13192,N_12306);
or U14397 (N_14397,N_12947,N_12321);
nor U14398 (N_14398,N_12482,N_12814);
and U14399 (N_14399,N_13190,N_13509);
nor U14400 (N_14400,N_13195,N_12835);
nor U14401 (N_14401,N_12255,N_12556);
nand U14402 (N_14402,N_12885,N_13692);
or U14403 (N_14403,N_12550,N_13129);
and U14404 (N_14404,N_12607,N_12113);
nand U14405 (N_14405,N_12504,N_13428);
nand U14406 (N_14406,N_13453,N_12429);
nor U14407 (N_14407,N_13893,N_13393);
or U14408 (N_14408,N_12594,N_13519);
nor U14409 (N_14409,N_12371,N_13400);
and U14410 (N_14410,N_12156,N_13225);
or U14411 (N_14411,N_12555,N_12541);
and U14412 (N_14412,N_12535,N_12843);
or U14413 (N_14413,N_12424,N_13773);
or U14414 (N_14414,N_12913,N_12399);
nor U14415 (N_14415,N_13602,N_13300);
nand U14416 (N_14416,N_13395,N_13314);
and U14417 (N_14417,N_13323,N_12939);
nor U14418 (N_14418,N_13686,N_13025);
nor U14419 (N_14419,N_12304,N_13819);
or U14420 (N_14420,N_13214,N_13274);
or U14421 (N_14421,N_12209,N_12097);
nor U14422 (N_14422,N_13542,N_12821);
or U14423 (N_14423,N_13528,N_13165);
and U14424 (N_14424,N_13156,N_13249);
nor U14425 (N_14425,N_12058,N_12684);
nor U14426 (N_14426,N_13648,N_13255);
or U14427 (N_14427,N_12496,N_12667);
or U14428 (N_14428,N_13880,N_12757);
or U14429 (N_14429,N_13746,N_13712);
nor U14430 (N_14430,N_12020,N_12517);
nor U14431 (N_14431,N_12135,N_13640);
and U14432 (N_14432,N_12419,N_12643);
or U14433 (N_14433,N_12197,N_13574);
nand U14434 (N_14434,N_13138,N_12571);
nor U14435 (N_14435,N_13594,N_12891);
or U14436 (N_14436,N_12779,N_12975);
nor U14437 (N_14437,N_13769,N_13388);
or U14438 (N_14438,N_13588,N_13641);
or U14439 (N_14439,N_12074,N_12177);
xor U14440 (N_14440,N_12434,N_13124);
and U14441 (N_14441,N_12078,N_13507);
nor U14442 (N_14442,N_12666,N_12711);
nand U14443 (N_14443,N_13231,N_12645);
nor U14444 (N_14444,N_12153,N_13361);
and U14445 (N_14445,N_12316,N_12878);
or U14446 (N_14446,N_13462,N_12223);
nand U14447 (N_14447,N_12288,N_12426);
or U14448 (N_14448,N_12007,N_13764);
or U14449 (N_14449,N_13711,N_12366);
nand U14450 (N_14450,N_13166,N_13704);
nor U14451 (N_14451,N_13033,N_12630);
nor U14452 (N_14452,N_12253,N_13168);
xor U14453 (N_14453,N_13044,N_13570);
nand U14454 (N_14454,N_13293,N_12518);
nor U14455 (N_14455,N_13849,N_12857);
nor U14456 (N_14456,N_12721,N_13392);
or U14457 (N_14457,N_12914,N_12978);
or U14458 (N_14458,N_12006,N_13405);
or U14459 (N_14459,N_12989,N_13853);
xor U14460 (N_14460,N_13331,N_13959);
or U14461 (N_14461,N_13644,N_12039);
and U14462 (N_14462,N_12865,N_12227);
nor U14463 (N_14463,N_13149,N_13761);
xnor U14464 (N_14464,N_12022,N_13642);
nand U14465 (N_14465,N_12259,N_13984);
nand U14466 (N_14466,N_12846,N_12691);
nand U14467 (N_14467,N_13902,N_12203);
xor U14468 (N_14468,N_12318,N_13312);
nand U14469 (N_14469,N_13899,N_13061);
and U14470 (N_14470,N_13971,N_12291);
nor U14471 (N_14471,N_12563,N_12506);
nor U14472 (N_14472,N_12248,N_13589);
or U14473 (N_14473,N_13460,N_13223);
nand U14474 (N_14474,N_13669,N_13978);
xnor U14475 (N_14475,N_13756,N_12351);
and U14476 (N_14476,N_13282,N_12707);
xnor U14477 (N_14477,N_13973,N_13958);
nand U14478 (N_14478,N_12704,N_13080);
xnor U14479 (N_14479,N_13418,N_13229);
or U14480 (N_14480,N_13979,N_13941);
nor U14481 (N_14481,N_13272,N_13534);
nand U14482 (N_14482,N_12798,N_13854);
nand U14483 (N_14483,N_13543,N_13289);
xnor U14484 (N_14484,N_12567,N_13981);
nand U14485 (N_14485,N_12993,N_13215);
nand U14486 (N_14486,N_13444,N_13488);
xnor U14487 (N_14487,N_13002,N_12952);
nor U14488 (N_14488,N_13607,N_13956);
or U14489 (N_14489,N_12646,N_12173);
or U14490 (N_14490,N_12445,N_13099);
nand U14491 (N_14491,N_13217,N_12370);
nor U14492 (N_14492,N_13595,N_12405);
and U14493 (N_14493,N_13364,N_13657);
and U14494 (N_14494,N_12752,N_13147);
or U14495 (N_14495,N_12692,N_13737);
xnor U14496 (N_14496,N_13536,N_13466);
and U14497 (N_14497,N_12527,N_13731);
or U14498 (N_14498,N_12330,N_12046);
or U14499 (N_14499,N_12849,N_13449);
nand U14500 (N_14500,N_12871,N_12688);
nand U14501 (N_14501,N_13663,N_13875);
or U14502 (N_14502,N_12166,N_12954);
or U14503 (N_14503,N_12077,N_12883);
and U14504 (N_14504,N_12790,N_13651);
and U14505 (N_14505,N_13510,N_13283);
and U14506 (N_14506,N_12280,N_13243);
nand U14507 (N_14507,N_13134,N_12363);
nand U14508 (N_14508,N_12295,N_12139);
nor U14509 (N_14509,N_12842,N_13730);
and U14510 (N_14510,N_12219,N_12887);
nor U14511 (N_14511,N_13338,N_13353);
xor U14512 (N_14512,N_12513,N_12284);
xor U14513 (N_14513,N_12374,N_12002);
and U14514 (N_14514,N_13583,N_12523);
or U14515 (N_14515,N_12893,N_12724);
nor U14516 (N_14516,N_13159,N_13037);
and U14517 (N_14517,N_12897,N_12492);
or U14518 (N_14518,N_13600,N_13336);
and U14519 (N_14519,N_13619,N_12618);
xor U14520 (N_14520,N_12061,N_13115);
and U14521 (N_14521,N_12515,N_13591);
nor U14522 (N_14522,N_13921,N_12185);
or U14523 (N_14523,N_12881,N_13850);
nand U14524 (N_14524,N_12403,N_12428);
xor U14525 (N_14525,N_13051,N_13627);
nor U14526 (N_14526,N_12962,N_12420);
xor U14527 (N_14527,N_13716,N_12254);
nand U14528 (N_14528,N_12327,N_13360);
nor U14529 (N_14529,N_13796,N_13379);
and U14530 (N_14530,N_13191,N_13459);
or U14531 (N_14531,N_12652,N_12894);
nor U14532 (N_14532,N_13568,N_13038);
xor U14533 (N_14533,N_13026,N_12936);
nor U14534 (N_14534,N_12211,N_12364);
xor U14535 (N_14535,N_13102,N_13976);
nor U14536 (N_14536,N_13952,N_12335);
and U14537 (N_14537,N_13605,N_12973);
or U14538 (N_14538,N_12215,N_13083);
nand U14539 (N_14539,N_13910,N_13750);
nand U14540 (N_14540,N_12325,N_13245);
nand U14541 (N_14541,N_13859,N_13319);
xnor U14542 (N_14542,N_13394,N_12788);
xnor U14543 (N_14543,N_13069,N_12472);
or U14544 (N_14544,N_12242,N_13725);
xnor U14545 (N_14545,N_12107,N_12213);
or U14546 (N_14546,N_12087,N_13382);
nor U14547 (N_14547,N_13258,N_13728);
nand U14548 (N_14548,N_13009,N_13832);
nand U14549 (N_14549,N_13565,N_13292);
nand U14550 (N_14550,N_12140,N_12693);
nor U14551 (N_14551,N_12474,N_12251);
nor U14552 (N_14552,N_12296,N_13643);
nand U14553 (N_14553,N_13987,N_13935);
xor U14554 (N_14554,N_13408,N_12746);
and U14555 (N_14555,N_12530,N_12815);
xnor U14556 (N_14556,N_13332,N_13232);
and U14557 (N_14557,N_13142,N_12856);
xnor U14558 (N_14558,N_13647,N_12167);
or U14559 (N_14559,N_12430,N_12060);
or U14560 (N_14560,N_12072,N_12080);
or U14561 (N_14561,N_12681,N_12825);
nand U14562 (N_14562,N_12627,N_12750);
xor U14563 (N_14563,N_13945,N_13325);
nor U14564 (N_14564,N_13943,N_12260);
and U14565 (N_14565,N_13671,N_12286);
nand U14566 (N_14566,N_12220,N_13007);
and U14567 (N_14567,N_12665,N_12262);
nor U14568 (N_14568,N_13585,N_12922);
nor U14569 (N_14569,N_13304,N_12308);
and U14570 (N_14570,N_12382,N_13940);
nor U14571 (N_14571,N_12348,N_13919);
or U14572 (N_14572,N_12826,N_13472);
or U14573 (N_14573,N_12867,N_12599);
and U14574 (N_14574,N_12154,N_12361);
nand U14575 (N_14575,N_13513,N_12189);
xnor U14576 (N_14576,N_12269,N_12038);
nor U14577 (N_14577,N_13431,N_13577);
and U14578 (N_14578,N_13135,N_13729);
and U14579 (N_14579,N_13342,N_13606);
nand U14580 (N_14580,N_12612,N_12660);
nand U14581 (N_14581,N_13792,N_12812);
xor U14582 (N_14582,N_13670,N_13363);
nand U14583 (N_14583,N_12770,N_12811);
nand U14584 (N_14584,N_13864,N_13795);
nand U14585 (N_14585,N_13143,N_12407);
nand U14586 (N_14586,N_12888,N_12916);
nand U14587 (N_14587,N_12536,N_13706);
nand U14588 (N_14588,N_12537,N_13913);
and U14589 (N_14589,N_13695,N_12088);
or U14590 (N_14590,N_13751,N_13004);
or U14591 (N_14591,N_13537,N_13782);
nor U14592 (N_14592,N_12198,N_13871);
nand U14593 (N_14593,N_13625,N_12236);
and U14594 (N_14594,N_13113,N_13763);
nand U14595 (N_14595,N_12950,N_12128);
nand U14596 (N_14596,N_13176,N_13020);
nor U14597 (N_14597,N_13066,N_13359);
and U14598 (N_14598,N_12204,N_13931);
and U14599 (N_14599,N_13397,N_12049);
nor U14600 (N_14600,N_13298,N_13634);
nor U14601 (N_14601,N_13748,N_13920);
or U14602 (N_14602,N_13491,N_13780);
nand U14603 (N_14603,N_12309,N_12860);
or U14604 (N_14604,N_13582,N_13368);
nand U14605 (N_14605,N_12232,N_12400);
and U14606 (N_14606,N_13067,N_13227);
xnor U14607 (N_14607,N_12937,N_13148);
nor U14608 (N_14608,N_12311,N_12990);
nand U14609 (N_14609,N_13082,N_13209);
xor U14610 (N_14610,N_13515,N_13456);
nand U14611 (N_14611,N_12138,N_12751);
and U14612 (N_14612,N_13957,N_12422);
nand U14613 (N_14613,N_12328,N_13305);
or U14614 (N_14614,N_12905,N_13807);
and U14615 (N_14615,N_12718,N_13983);
nor U14616 (N_14616,N_13018,N_13116);
or U14617 (N_14617,N_12471,N_12593);
nor U14618 (N_14618,N_12949,N_13154);
and U14619 (N_14619,N_12273,N_12137);
or U14620 (N_14620,N_13275,N_13091);
or U14621 (N_14621,N_13029,N_13070);
and U14622 (N_14622,N_12520,N_13872);
nand U14623 (N_14623,N_12483,N_12841);
and U14624 (N_14624,N_12982,N_13356);
xnor U14625 (N_14625,N_13950,N_12036);
nand U14626 (N_14626,N_12581,N_13540);
and U14627 (N_14627,N_13132,N_12437);
and U14628 (N_14628,N_12449,N_12738);
and U14629 (N_14629,N_12312,N_13045);
or U14630 (N_14630,N_13532,N_13030);
nand U14631 (N_14631,N_13734,N_12226);
or U14632 (N_14632,N_12170,N_13486);
nand U14633 (N_14633,N_13181,N_12158);
nand U14634 (N_14634,N_12362,N_13307);
nand U14635 (N_14635,N_13308,N_12908);
nand U14636 (N_14636,N_12834,N_12412);
nor U14637 (N_14637,N_12071,N_13162);
nor U14638 (N_14638,N_13752,N_13996);
nor U14639 (N_14639,N_12027,N_13077);
nand U14640 (N_14640,N_12266,N_13674);
nand U14641 (N_14641,N_12491,N_13199);
or U14642 (N_14642,N_13630,N_13928);
nand U14643 (N_14643,N_12169,N_12759);
nand U14644 (N_14644,N_13679,N_13933);
and U14645 (N_14645,N_12884,N_13546);
nor U14646 (N_14646,N_13417,N_12085);
or U14647 (N_14647,N_13427,N_13492);
and U14648 (N_14648,N_13781,N_12705);
and U14649 (N_14649,N_12413,N_13241);
and U14650 (N_14650,N_13212,N_13387);
or U14651 (N_14651,N_12147,N_13522);
and U14652 (N_14652,N_12476,N_12182);
and U14653 (N_14653,N_13982,N_13754);
nor U14654 (N_14654,N_13146,N_12207);
and U14655 (N_14655,N_13653,N_13335);
nand U14656 (N_14656,N_13960,N_13471);
nand U14657 (N_14657,N_12326,N_13812);
or U14658 (N_14658,N_12591,N_12675);
or U14659 (N_14659,N_13965,N_13885);
and U14660 (N_14660,N_12377,N_13017);
xor U14661 (N_14661,N_12467,N_13288);
nand U14662 (N_14662,N_12276,N_13977);
nor U14663 (N_14663,N_12337,N_12629);
or U14664 (N_14664,N_13841,N_13060);
or U14665 (N_14665,N_12360,N_13626);
nor U14666 (N_14666,N_13884,N_13997);
and U14667 (N_14667,N_13771,N_13573);
nand U14668 (N_14668,N_13613,N_12722);
or U14669 (N_14669,N_13549,N_13236);
nand U14670 (N_14670,N_13052,N_12421);
xor U14671 (N_14671,N_12493,N_12503);
xnor U14672 (N_14672,N_12458,N_13690);
or U14673 (N_14673,N_12486,N_13263);
or U14674 (N_14674,N_13187,N_12801);
and U14675 (N_14675,N_12621,N_12768);
xor U14676 (N_14676,N_13078,N_13779);
and U14677 (N_14677,N_12634,N_13862);
xor U14678 (N_14678,N_12221,N_12051);
or U14679 (N_14679,N_12283,N_13688);
nand U14680 (N_14680,N_13666,N_12793);
and U14681 (N_14681,N_12414,N_13579);
nand U14682 (N_14682,N_12816,N_12157);
or U14683 (N_14683,N_12301,N_12136);
nand U14684 (N_14684,N_13315,N_13425);
and U14685 (N_14685,N_12216,N_13271);
and U14686 (N_14686,N_12461,N_13942);
or U14687 (N_14687,N_12587,N_12786);
or U14688 (N_14688,N_13758,N_12032);
and U14689 (N_14689,N_13081,N_12622);
xnor U14690 (N_14690,N_12999,N_12709);
and U14691 (N_14691,N_13557,N_13270);
nand U14692 (N_14692,N_13684,N_12931);
nor U14693 (N_14693,N_12237,N_12543);
nor U14694 (N_14694,N_13857,N_12053);
nor U14695 (N_14695,N_13259,N_12332);
nand U14696 (N_14696,N_12289,N_13609);
or U14697 (N_14697,N_13628,N_13708);
or U14698 (N_14698,N_12870,N_13087);
nand U14699 (N_14699,N_12761,N_12514);
or U14700 (N_14700,N_13442,N_12381);
or U14701 (N_14701,N_12026,N_12122);
or U14702 (N_14702,N_13445,N_12926);
nor U14703 (N_14703,N_13629,N_13184);
nor U14704 (N_14704,N_13257,N_12780);
nor U14705 (N_14705,N_13714,N_13008);
or U14706 (N_14706,N_13811,N_13090);
and U14707 (N_14707,N_13904,N_12702);
nor U14708 (N_14708,N_12512,N_13014);
and U14709 (N_14709,N_12639,N_13637);
and U14710 (N_14710,N_12401,N_13207);
or U14711 (N_14711,N_12396,N_13233);
nor U14712 (N_14712,N_13847,N_13733);
nand U14713 (N_14713,N_13333,N_12917);
or U14714 (N_14714,N_13186,N_13755);
nor U14715 (N_14715,N_12521,N_12731);
nor U14716 (N_14716,N_13446,N_13970);
nor U14717 (N_14717,N_13301,N_12037);
nor U14718 (N_14718,N_12833,N_13476);
xnor U14719 (N_14719,N_12068,N_13337);
and U14720 (N_14720,N_13791,N_13822);
or U14721 (N_14721,N_12342,N_13767);
nand U14722 (N_14722,N_13759,N_12676);
nand U14723 (N_14723,N_12892,N_12195);
or U14724 (N_14724,N_12754,N_13114);
or U14725 (N_14725,N_12021,N_13560);
nor U14726 (N_14726,N_13991,N_12485);
or U14727 (N_14727,N_13469,N_13766);
and U14728 (N_14728,N_13553,N_12651);
or U14729 (N_14729,N_13618,N_13790);
or U14730 (N_14730,N_13357,N_12444);
and U14731 (N_14731,N_12345,N_13224);
or U14732 (N_14732,N_13521,N_12827);
or U14733 (N_14733,N_12547,N_13221);
nand U14734 (N_14734,N_13508,N_12800);
or U14735 (N_14735,N_12473,N_12785);
nand U14736 (N_14736,N_12180,N_12205);
nand U14737 (N_14737,N_13228,N_12992);
xor U14738 (N_14738,N_12323,N_12372);
and U14739 (N_14739,N_12628,N_12686);
nand U14740 (N_14740,N_12644,N_12701);
or U14741 (N_14741,N_13757,N_13406);
nand U14742 (N_14742,N_12448,N_13883);
or U14743 (N_14743,N_13550,N_12439);
xnor U14744 (N_14744,N_13598,N_12689);
and U14745 (N_14745,N_12054,N_13911);
nor U14746 (N_14746,N_12551,N_13616);
nor U14747 (N_14747,N_13837,N_13820);
and U14748 (N_14748,N_13396,N_12352);
or U14749 (N_14749,N_13559,N_13188);
xor U14750 (N_14750,N_12322,N_12141);
nand U14751 (N_14751,N_12305,N_13180);
and U14752 (N_14752,N_12110,N_12252);
nor U14753 (N_14753,N_12526,N_12040);
or U14754 (N_14754,N_13299,N_13039);
or U14755 (N_14755,N_13484,N_12624);
and U14756 (N_14756,N_13803,N_13813);
xor U14757 (N_14757,N_12861,N_13244);
xor U14758 (N_14758,N_12235,N_12656);
or U14759 (N_14759,N_13478,N_13901);
nand U14760 (N_14760,N_12617,N_12650);
nand U14761 (N_14761,N_13126,N_12700);
nor U14762 (N_14762,N_13122,N_12261);
and U14763 (N_14763,N_12697,N_12880);
or U14764 (N_14764,N_13735,N_12104);
nand U14765 (N_14765,N_12033,N_12560);
xnor U14766 (N_14766,N_12531,N_13527);
nor U14767 (N_14767,N_12839,N_13059);
nand U14768 (N_14768,N_12334,N_13093);
or U14769 (N_14769,N_13262,N_12943);
or U14770 (N_14770,N_13145,N_13985);
and U14771 (N_14771,N_13760,N_13808);
or U14772 (N_14772,N_13189,N_13169);
and U14773 (N_14773,N_12270,N_13838);
xor U14774 (N_14774,N_12303,N_13689);
xor U14775 (N_14775,N_12778,N_12620);
and U14776 (N_14776,N_13932,N_12869);
and U14777 (N_14777,N_12310,N_12776);
and U14778 (N_14778,N_13567,N_13768);
and U14779 (N_14779,N_13269,N_13892);
nor U14780 (N_14780,N_13384,N_13924);
or U14781 (N_14781,N_13865,N_12729);
and U14782 (N_14782,N_12742,N_13569);
and U14783 (N_14783,N_13286,N_12298);
or U14784 (N_14784,N_12052,N_12889);
nor U14785 (N_14785,N_12126,N_12955);
nand U14786 (N_14786,N_12212,N_12744);
nor U14787 (N_14787,N_13309,N_13328);
or U14788 (N_14788,N_12998,N_12960);
and U14789 (N_14789,N_13071,N_13846);
or U14790 (N_14790,N_13840,N_13056);
and U14791 (N_14791,N_13701,N_12561);
nand U14792 (N_14792,N_12191,N_13351);
and U14793 (N_14793,N_13601,N_12734);
nor U14794 (N_14794,N_13995,N_12771);
nor U14795 (N_14795,N_12654,N_13691);
and U14796 (N_14796,N_12481,N_13034);
nor U14797 (N_14797,N_12866,N_13844);
or U14798 (N_14798,N_13050,N_13474);
nor U14799 (N_14799,N_13178,N_12488);
or U14800 (N_14800,N_12608,N_12358);
or U14801 (N_14801,N_12590,N_13962);
or U14802 (N_14802,N_12117,N_13172);
nor U14803 (N_14803,N_13341,N_12958);
nor U14804 (N_14804,N_12736,N_13578);
xor U14805 (N_14805,N_13974,N_13707);
xor U14806 (N_14806,N_13882,N_13496);
or U14807 (N_14807,N_12460,N_13836);
xor U14808 (N_14808,N_12545,N_13925);
nor U14809 (N_14809,N_12299,N_12655);
and U14810 (N_14810,N_13538,N_12076);
and U14811 (N_14811,N_13220,N_12806);
nor U14812 (N_14812,N_13742,N_12925);
and U14813 (N_14813,N_12600,N_12392);
or U14814 (N_14814,N_12715,N_12100);
or U14815 (N_14815,N_13112,N_13375);
and U14816 (N_14816,N_12009,N_12171);
or U14817 (N_14817,N_13321,N_12877);
nor U14818 (N_14818,N_13455,N_12706);
xor U14819 (N_14819,N_12907,N_12533);
nor U14820 (N_14820,N_12851,N_12565);
and U14821 (N_14821,N_12194,N_13963);
and U14822 (N_14822,N_13753,N_13448);
nor U14823 (N_14823,N_12965,N_13043);
and U14824 (N_14824,N_12832,N_13739);
or U14825 (N_14825,N_12160,N_12324);
nor U14826 (N_14826,N_12847,N_12807);
or U14827 (N_14827,N_12564,N_13672);
and U14828 (N_14828,N_12725,N_12249);
or U14829 (N_14829,N_12796,N_13867);
or U14830 (N_14830,N_13306,N_12183);
nand U14831 (N_14831,N_13003,N_12477);
xor U14832 (N_14832,N_13966,N_12896);
nor U14833 (N_14833,N_12586,N_13877);
and U14834 (N_14834,N_13861,N_13660);
or U14835 (N_14835,N_12404,N_13709);
nand U14836 (N_14836,N_12670,N_12647);
nor U14837 (N_14837,N_12069,N_12089);
and U14838 (N_14838,N_13946,N_12769);
xor U14839 (N_14839,N_13934,N_12442);
nor U14840 (N_14840,N_12606,N_12765);
xor U14841 (N_14841,N_12383,N_12184);
nor U14842 (N_14842,N_12144,N_13964);
and U14843 (N_14843,N_12921,N_13525);
nor U14844 (N_14844,N_12073,N_13205);
and U14845 (N_14845,N_12583,N_12935);
nand U14846 (N_14846,N_12292,N_12408);
and U14847 (N_14847,N_13817,N_13144);
and U14848 (N_14848,N_12756,N_12876);
nand U14849 (N_14849,N_13785,N_12544);
nor U14850 (N_14850,N_13907,N_12145);
xor U14851 (N_14851,N_13177,N_12813);
and U14852 (N_14852,N_12640,N_12940);
xor U14853 (N_14853,N_13032,N_13727);
nor U14854 (N_14854,N_13908,N_12758);
and U14855 (N_14855,N_12159,N_12056);
or U14856 (N_14856,N_12048,N_12155);
or U14857 (N_14857,N_13104,N_13989);
and U14858 (N_14858,N_12580,N_12577);
or U14859 (N_14859,N_12484,N_12977);
nand U14860 (N_14860,N_13419,N_12525);
nor U14861 (N_14861,N_12108,N_12457);
nand U14862 (N_14862,N_13586,N_12854);
nor U14863 (N_14863,N_12179,N_12098);
or U14864 (N_14864,N_13747,N_12375);
nand U14865 (N_14865,N_12605,N_12313);
and U14866 (N_14866,N_13866,N_12023);
or U14867 (N_14867,N_12278,N_13021);
nor U14868 (N_14868,N_13479,N_12772);
nand U14869 (N_14869,N_13818,N_12695);
xor U14870 (N_14870,N_12062,N_12733);
or U14871 (N_14871,N_13423,N_13723);
or U14872 (N_14872,N_13276,N_13955);
and U14873 (N_14873,N_12294,N_12379);
xor U14874 (N_14874,N_13370,N_13076);
nor U14875 (N_14875,N_13279,N_13432);
nor U14876 (N_14876,N_13516,N_13340);
or U14877 (N_14877,N_12795,N_13658);
xor U14878 (N_14878,N_13972,N_12031);
nor U14879 (N_14879,N_12661,N_13010);
nor U14880 (N_14880,N_13391,N_13635);
nor U14881 (N_14881,N_13732,N_12431);
nand U14882 (N_14882,N_12648,N_12572);
nand U14883 (N_14883,N_12712,N_12635);
or U14884 (N_14884,N_13561,N_13592);
nand U14885 (N_14885,N_12287,N_12576);
or U14886 (N_14886,N_13330,N_13376);
nand U14887 (N_14887,N_12824,N_13251);
nand U14888 (N_14888,N_13410,N_12106);
nand U14889 (N_14889,N_13896,N_12764);
nor U14890 (N_14890,N_12864,N_13915);
or U14891 (N_14891,N_12410,N_12497);
xnor U14892 (N_14892,N_12579,N_12528);
nand U14893 (N_14893,N_13440,N_13324);
or U14894 (N_14894,N_13497,N_12957);
or U14895 (N_14895,N_13447,N_13775);
nand U14896 (N_14896,N_13681,N_12726);
xnor U14897 (N_14897,N_12281,N_12385);
nand U14898 (N_14898,N_12187,N_13554);
nand U14899 (N_14899,N_13001,N_13412);
xnor U14900 (N_14900,N_13999,N_12573);
nand U14901 (N_14901,N_13311,N_12845);
xor U14902 (N_14902,N_13954,N_12678);
and U14903 (N_14903,N_12102,N_13881);
nor U14904 (N_14904,N_13011,N_13106);
nand U14905 (N_14905,N_13118,N_13646);
nand U14906 (N_14906,N_13437,N_13917);
xnor U14907 (N_14907,N_12133,N_12438);
and U14908 (N_14908,N_13354,N_12152);
xnor U14909 (N_14909,N_12475,N_13888);
or U14910 (N_14910,N_13624,N_13721);
and U14911 (N_14911,N_13386,N_13772);
or U14912 (N_14912,N_13012,N_12735);
or U14913 (N_14913,N_13652,N_12228);
and U14914 (N_14914,N_12714,N_12636);
and U14915 (N_14915,N_13668,N_13088);
and U14916 (N_14916,N_12956,N_13151);
nor U14917 (N_14917,N_13685,N_13810);
or U14918 (N_14918,N_13264,N_13992);
nor U14919 (N_14919,N_12616,N_13798);
and U14920 (N_14920,N_13477,N_12091);
xor U14921 (N_14921,N_12767,N_12423);
or U14922 (N_14922,N_12417,N_12566);
and U14923 (N_14923,N_12199,N_12013);
nor U14924 (N_14924,N_13196,N_12524);
or U14925 (N_14925,N_13105,N_13499);
nor U14926 (N_14926,N_12208,N_12862);
nor U14927 (N_14927,N_12192,N_12760);
or U14928 (N_14928,N_13150,N_13517);
or U14929 (N_14929,N_12453,N_13874);
nand U14930 (N_14930,N_12353,N_12150);
nand U14931 (N_14931,N_13450,N_12837);
or U14932 (N_14932,N_12777,N_12649);
or U14933 (N_14933,N_12045,N_12668);
or U14934 (N_14934,N_12297,N_13953);
and U14935 (N_14935,N_12539,N_12008);
nor U14936 (N_14936,N_13402,N_12084);
nor U14937 (N_14937,N_12393,N_12802);
and U14938 (N_14938,N_13696,N_12679);
nand U14939 (N_14939,N_12432,N_12799);
and U14940 (N_14940,N_13608,N_13403);
nand U14941 (N_14941,N_13939,N_13107);
nor U14942 (N_14942,N_12406,N_13058);
and U14943 (N_14943,N_12024,N_13937);
nand U14944 (N_14944,N_12190,N_13564);
nor U14945 (N_14945,N_12898,N_13092);
nor U14946 (N_14946,N_13994,N_13547);
and U14947 (N_14947,N_12542,N_12868);
nand U14948 (N_14948,N_13470,N_13777);
nand U14949 (N_14949,N_13967,N_12924);
and U14950 (N_14950,N_13280,N_13738);
nor U14951 (N_14951,N_13590,N_13238);
xor U14952 (N_14952,N_13555,N_13480);
nor U14953 (N_14953,N_12202,N_12011);
and U14954 (N_14954,N_12633,N_12619);
and U14955 (N_14955,N_12810,N_12302);
nor U14956 (N_14956,N_12903,N_13174);
and U14957 (N_14957,N_12450,N_12489);
or U14958 (N_14958,N_13040,N_13675);
nand U14959 (N_14959,N_13617,N_12115);
nand U14960 (N_14960,N_13726,N_12708);
nand U14961 (N_14961,N_12942,N_12175);
nand U14962 (N_14962,N_13171,N_13702);
nand U14963 (N_14963,N_12625,N_13239);
nor U14964 (N_14964,N_12595,N_12853);
nor U14965 (N_14965,N_12282,N_13164);
nor U14966 (N_14966,N_13826,N_13717);
nor U14967 (N_14967,N_12116,N_12415);
nor U14968 (N_14968,N_12446,N_12333);
and U14969 (N_14969,N_13253,N_12161);
nand U14970 (N_14970,N_12454,N_13584);
nor U14971 (N_14971,N_13439,N_13316);
xnor U14972 (N_14972,N_12703,N_12436);
and U14973 (N_14973,N_13234,N_13404);
nor U14974 (N_14974,N_12710,N_13927);
or U14975 (N_14975,N_13248,N_12402);
nor U14976 (N_14976,N_12210,N_12151);
nand U14977 (N_14977,N_13362,N_13916);
nor U14978 (N_14978,N_13562,N_12433);
nor U14979 (N_14979,N_13587,N_13023);
nor U14980 (N_14980,N_13237,N_13481);
nor U14981 (N_14981,N_12981,N_13533);
and U14982 (N_14982,N_13720,N_13834);
or U14983 (N_14983,N_13891,N_13458);
xor U14984 (N_14984,N_13741,N_12623);
or U14985 (N_14985,N_13019,N_12820);
nand U14986 (N_14986,N_12394,N_12946);
nand U14987 (N_14987,N_12245,N_12909);
nor U14988 (N_14988,N_13615,N_12050);
or U14989 (N_14989,N_13575,N_12329);
xnor U14990 (N_14990,N_12928,N_13667);
and U14991 (N_14991,N_13879,N_12596);
and U14992 (N_14992,N_12043,N_13267);
and U14993 (N_14993,N_12075,N_12468);
nor U14994 (N_14994,N_13339,N_13694);
xnor U14995 (N_14995,N_13611,N_13778);
nor U14996 (N_14996,N_13612,N_12529);
or U14997 (N_14997,N_12505,N_12148);
or U14998 (N_14998,N_12985,N_12979);
nor U14999 (N_14999,N_13167,N_12836);
or U15000 (N_15000,N_13563,N_12213);
and U15001 (N_15001,N_13334,N_13508);
or U15002 (N_15002,N_13901,N_12050);
nand U15003 (N_15003,N_12989,N_13192);
nor U15004 (N_15004,N_13760,N_13867);
nor U15005 (N_15005,N_12181,N_13958);
nand U15006 (N_15006,N_12720,N_12384);
xnor U15007 (N_15007,N_13341,N_12762);
nor U15008 (N_15008,N_13210,N_12044);
nor U15009 (N_15009,N_13056,N_12966);
and U15010 (N_15010,N_12815,N_12858);
nor U15011 (N_15011,N_12629,N_12205);
and U15012 (N_15012,N_13947,N_12910);
nand U15013 (N_15013,N_13780,N_12341);
nand U15014 (N_15014,N_12325,N_12831);
and U15015 (N_15015,N_12171,N_12099);
nor U15016 (N_15016,N_12673,N_12126);
nand U15017 (N_15017,N_13972,N_13372);
nand U15018 (N_15018,N_12834,N_13669);
xnor U15019 (N_15019,N_13748,N_12759);
nand U15020 (N_15020,N_12846,N_12483);
nand U15021 (N_15021,N_13843,N_13985);
nor U15022 (N_15022,N_13504,N_13314);
and U15023 (N_15023,N_13825,N_13440);
nand U15024 (N_15024,N_12499,N_13583);
or U15025 (N_15025,N_12390,N_13384);
and U15026 (N_15026,N_13236,N_13425);
nor U15027 (N_15027,N_13386,N_12224);
nor U15028 (N_15028,N_13779,N_12238);
and U15029 (N_15029,N_13024,N_13537);
and U15030 (N_15030,N_13368,N_12751);
and U15031 (N_15031,N_13901,N_12775);
nand U15032 (N_15032,N_13681,N_12112);
nand U15033 (N_15033,N_13311,N_12240);
or U15034 (N_15034,N_13233,N_13333);
nand U15035 (N_15035,N_13765,N_13307);
xor U15036 (N_15036,N_13934,N_13732);
nand U15037 (N_15037,N_12190,N_12840);
or U15038 (N_15038,N_12852,N_13530);
nand U15039 (N_15039,N_13804,N_12062);
nor U15040 (N_15040,N_13797,N_13638);
and U15041 (N_15041,N_12041,N_12388);
nand U15042 (N_15042,N_12470,N_13399);
nand U15043 (N_15043,N_12087,N_12408);
xor U15044 (N_15044,N_12428,N_13011);
and U15045 (N_15045,N_13852,N_12912);
and U15046 (N_15046,N_13257,N_13432);
nor U15047 (N_15047,N_13515,N_13150);
and U15048 (N_15048,N_12242,N_12253);
nand U15049 (N_15049,N_12418,N_13590);
nor U15050 (N_15050,N_13725,N_13510);
or U15051 (N_15051,N_13561,N_13657);
nand U15052 (N_15052,N_12736,N_13906);
and U15053 (N_15053,N_13393,N_13429);
and U15054 (N_15054,N_12281,N_12571);
or U15055 (N_15055,N_13530,N_12977);
and U15056 (N_15056,N_12135,N_13409);
nand U15057 (N_15057,N_12880,N_13342);
or U15058 (N_15058,N_13323,N_13263);
xnor U15059 (N_15059,N_12310,N_12915);
nor U15060 (N_15060,N_12745,N_13598);
or U15061 (N_15061,N_12535,N_13361);
nand U15062 (N_15062,N_13743,N_12387);
nor U15063 (N_15063,N_13563,N_12010);
nor U15064 (N_15064,N_13518,N_13187);
or U15065 (N_15065,N_13228,N_13999);
nor U15066 (N_15066,N_13798,N_13692);
xor U15067 (N_15067,N_13779,N_12326);
xnor U15068 (N_15068,N_12250,N_12357);
and U15069 (N_15069,N_12746,N_12786);
xor U15070 (N_15070,N_13337,N_13638);
nor U15071 (N_15071,N_12995,N_12969);
and U15072 (N_15072,N_12202,N_12829);
and U15073 (N_15073,N_13334,N_12372);
nor U15074 (N_15074,N_13983,N_13376);
xor U15075 (N_15075,N_12309,N_13285);
and U15076 (N_15076,N_12802,N_13930);
or U15077 (N_15077,N_13149,N_13381);
and U15078 (N_15078,N_12626,N_13092);
xnor U15079 (N_15079,N_12399,N_13035);
nor U15080 (N_15080,N_12882,N_12672);
and U15081 (N_15081,N_13414,N_13415);
and U15082 (N_15082,N_12977,N_13414);
or U15083 (N_15083,N_13204,N_13060);
nor U15084 (N_15084,N_13243,N_12501);
nand U15085 (N_15085,N_13451,N_12276);
nor U15086 (N_15086,N_12898,N_13704);
or U15087 (N_15087,N_13650,N_13531);
xor U15088 (N_15088,N_12980,N_13144);
or U15089 (N_15089,N_12575,N_13004);
nand U15090 (N_15090,N_13318,N_13917);
or U15091 (N_15091,N_13269,N_12098);
nand U15092 (N_15092,N_12721,N_12250);
xor U15093 (N_15093,N_13040,N_12134);
nand U15094 (N_15094,N_13982,N_12738);
or U15095 (N_15095,N_13593,N_13892);
nand U15096 (N_15096,N_13700,N_13037);
and U15097 (N_15097,N_13712,N_13488);
or U15098 (N_15098,N_13480,N_12357);
and U15099 (N_15099,N_13787,N_12795);
or U15100 (N_15100,N_12207,N_12719);
and U15101 (N_15101,N_12023,N_13532);
and U15102 (N_15102,N_13196,N_12772);
nand U15103 (N_15103,N_13885,N_12834);
and U15104 (N_15104,N_12630,N_12763);
and U15105 (N_15105,N_12157,N_12486);
or U15106 (N_15106,N_13657,N_12978);
and U15107 (N_15107,N_13061,N_12245);
or U15108 (N_15108,N_13388,N_13299);
nand U15109 (N_15109,N_12381,N_12590);
or U15110 (N_15110,N_12088,N_13585);
nand U15111 (N_15111,N_13871,N_13136);
and U15112 (N_15112,N_13408,N_12385);
and U15113 (N_15113,N_12754,N_12357);
and U15114 (N_15114,N_12769,N_13702);
and U15115 (N_15115,N_13814,N_12022);
xor U15116 (N_15116,N_12670,N_12725);
and U15117 (N_15117,N_13085,N_12464);
nand U15118 (N_15118,N_13631,N_13299);
or U15119 (N_15119,N_13900,N_13747);
and U15120 (N_15120,N_13176,N_12230);
nand U15121 (N_15121,N_12987,N_13906);
or U15122 (N_15122,N_12783,N_13007);
nand U15123 (N_15123,N_13477,N_13795);
and U15124 (N_15124,N_12759,N_13415);
or U15125 (N_15125,N_12625,N_12833);
nand U15126 (N_15126,N_13479,N_12146);
nor U15127 (N_15127,N_12910,N_12675);
nand U15128 (N_15128,N_12752,N_13442);
nor U15129 (N_15129,N_13424,N_13393);
nor U15130 (N_15130,N_13021,N_13807);
and U15131 (N_15131,N_12659,N_12541);
nor U15132 (N_15132,N_13683,N_12698);
xor U15133 (N_15133,N_13382,N_12499);
xor U15134 (N_15134,N_12331,N_12816);
nand U15135 (N_15135,N_13163,N_13711);
nand U15136 (N_15136,N_12032,N_13665);
and U15137 (N_15137,N_12510,N_13327);
nor U15138 (N_15138,N_12544,N_13341);
and U15139 (N_15139,N_13854,N_13602);
nor U15140 (N_15140,N_13937,N_13389);
nor U15141 (N_15141,N_13515,N_12254);
or U15142 (N_15142,N_12942,N_13449);
xor U15143 (N_15143,N_12755,N_12865);
nand U15144 (N_15144,N_12050,N_12542);
nand U15145 (N_15145,N_13134,N_13162);
nor U15146 (N_15146,N_12811,N_12195);
nor U15147 (N_15147,N_13231,N_12741);
or U15148 (N_15148,N_12426,N_13253);
and U15149 (N_15149,N_12792,N_12439);
and U15150 (N_15150,N_13433,N_13799);
nand U15151 (N_15151,N_12912,N_13472);
nand U15152 (N_15152,N_13225,N_12741);
nor U15153 (N_15153,N_12712,N_13584);
or U15154 (N_15154,N_12346,N_13906);
and U15155 (N_15155,N_12656,N_13697);
xnor U15156 (N_15156,N_12717,N_13288);
nor U15157 (N_15157,N_12783,N_12299);
xor U15158 (N_15158,N_13832,N_13393);
or U15159 (N_15159,N_13220,N_13787);
or U15160 (N_15160,N_13217,N_12668);
nand U15161 (N_15161,N_12892,N_13861);
or U15162 (N_15162,N_12313,N_12820);
or U15163 (N_15163,N_12520,N_12271);
xnor U15164 (N_15164,N_12651,N_13035);
and U15165 (N_15165,N_12341,N_12140);
nand U15166 (N_15166,N_12949,N_13367);
and U15167 (N_15167,N_12397,N_12256);
and U15168 (N_15168,N_13651,N_13628);
nor U15169 (N_15169,N_13979,N_13479);
nor U15170 (N_15170,N_12457,N_12550);
or U15171 (N_15171,N_12513,N_12404);
and U15172 (N_15172,N_13916,N_12823);
and U15173 (N_15173,N_12751,N_12936);
nand U15174 (N_15174,N_12805,N_12230);
nand U15175 (N_15175,N_13285,N_13539);
nor U15176 (N_15176,N_12101,N_12487);
nor U15177 (N_15177,N_13347,N_12386);
or U15178 (N_15178,N_13607,N_12063);
nand U15179 (N_15179,N_13744,N_13960);
nor U15180 (N_15180,N_13972,N_13690);
and U15181 (N_15181,N_13167,N_13542);
xnor U15182 (N_15182,N_13595,N_13100);
and U15183 (N_15183,N_12590,N_13905);
nand U15184 (N_15184,N_13767,N_12335);
or U15185 (N_15185,N_13528,N_13318);
nand U15186 (N_15186,N_13820,N_13826);
nand U15187 (N_15187,N_12344,N_13320);
nor U15188 (N_15188,N_13761,N_12222);
nand U15189 (N_15189,N_13483,N_12478);
and U15190 (N_15190,N_13166,N_13635);
nand U15191 (N_15191,N_13033,N_13493);
nand U15192 (N_15192,N_12939,N_13569);
xor U15193 (N_15193,N_13382,N_13927);
or U15194 (N_15194,N_12088,N_12801);
nor U15195 (N_15195,N_13027,N_13181);
nor U15196 (N_15196,N_13275,N_12979);
or U15197 (N_15197,N_13970,N_12943);
nor U15198 (N_15198,N_12431,N_12155);
and U15199 (N_15199,N_12689,N_13304);
and U15200 (N_15200,N_12227,N_13633);
and U15201 (N_15201,N_13563,N_12769);
or U15202 (N_15202,N_13856,N_13004);
nand U15203 (N_15203,N_12621,N_12819);
and U15204 (N_15204,N_13388,N_12397);
nor U15205 (N_15205,N_13741,N_13779);
xnor U15206 (N_15206,N_12416,N_13459);
nand U15207 (N_15207,N_12964,N_12588);
or U15208 (N_15208,N_13611,N_12740);
nor U15209 (N_15209,N_12737,N_12118);
nor U15210 (N_15210,N_13393,N_13609);
nor U15211 (N_15211,N_12501,N_13547);
or U15212 (N_15212,N_12914,N_13958);
or U15213 (N_15213,N_13442,N_12426);
xnor U15214 (N_15214,N_12688,N_12117);
nor U15215 (N_15215,N_13692,N_13750);
and U15216 (N_15216,N_12400,N_13759);
or U15217 (N_15217,N_13297,N_13985);
and U15218 (N_15218,N_13777,N_12094);
nor U15219 (N_15219,N_13212,N_12280);
nor U15220 (N_15220,N_12606,N_12558);
nand U15221 (N_15221,N_12889,N_13223);
and U15222 (N_15222,N_12133,N_12525);
nand U15223 (N_15223,N_13936,N_13781);
nand U15224 (N_15224,N_12849,N_12492);
nand U15225 (N_15225,N_12353,N_13351);
xor U15226 (N_15226,N_12094,N_12475);
nand U15227 (N_15227,N_13325,N_12419);
and U15228 (N_15228,N_12020,N_12372);
and U15229 (N_15229,N_13499,N_13634);
nand U15230 (N_15230,N_13087,N_13449);
nor U15231 (N_15231,N_13102,N_13985);
nand U15232 (N_15232,N_12730,N_13512);
nand U15233 (N_15233,N_12452,N_12561);
or U15234 (N_15234,N_13224,N_13614);
nor U15235 (N_15235,N_13061,N_12800);
nand U15236 (N_15236,N_12602,N_13070);
and U15237 (N_15237,N_13033,N_13278);
nand U15238 (N_15238,N_13145,N_13673);
and U15239 (N_15239,N_12876,N_12037);
and U15240 (N_15240,N_12574,N_13331);
and U15241 (N_15241,N_12511,N_12343);
or U15242 (N_15242,N_13410,N_13089);
nand U15243 (N_15243,N_13985,N_13952);
or U15244 (N_15244,N_12043,N_13548);
nor U15245 (N_15245,N_13170,N_13207);
and U15246 (N_15246,N_13223,N_12903);
or U15247 (N_15247,N_13955,N_12791);
and U15248 (N_15248,N_13508,N_12480);
and U15249 (N_15249,N_12523,N_13818);
xor U15250 (N_15250,N_13814,N_13565);
nor U15251 (N_15251,N_13783,N_12662);
and U15252 (N_15252,N_13926,N_12438);
or U15253 (N_15253,N_13618,N_13164);
or U15254 (N_15254,N_12358,N_13103);
and U15255 (N_15255,N_13095,N_12261);
and U15256 (N_15256,N_12356,N_13357);
or U15257 (N_15257,N_13170,N_12438);
nor U15258 (N_15258,N_12766,N_12139);
nor U15259 (N_15259,N_12148,N_13670);
nand U15260 (N_15260,N_13802,N_12949);
nor U15261 (N_15261,N_13046,N_13404);
and U15262 (N_15262,N_13679,N_12943);
or U15263 (N_15263,N_13354,N_12731);
and U15264 (N_15264,N_13550,N_13607);
and U15265 (N_15265,N_13731,N_13163);
nand U15266 (N_15266,N_13825,N_12279);
and U15267 (N_15267,N_12122,N_12436);
and U15268 (N_15268,N_12380,N_13083);
and U15269 (N_15269,N_13670,N_12918);
xor U15270 (N_15270,N_13021,N_13685);
nand U15271 (N_15271,N_13103,N_12003);
nand U15272 (N_15272,N_12027,N_12399);
nand U15273 (N_15273,N_12638,N_13123);
nor U15274 (N_15274,N_12922,N_13697);
nor U15275 (N_15275,N_12803,N_12821);
or U15276 (N_15276,N_12077,N_13614);
nor U15277 (N_15277,N_13410,N_12734);
nand U15278 (N_15278,N_12737,N_13789);
or U15279 (N_15279,N_13647,N_13079);
nor U15280 (N_15280,N_13069,N_12788);
nor U15281 (N_15281,N_13411,N_13078);
nand U15282 (N_15282,N_12298,N_12114);
and U15283 (N_15283,N_12536,N_13861);
or U15284 (N_15284,N_13680,N_12799);
and U15285 (N_15285,N_12046,N_12555);
or U15286 (N_15286,N_13341,N_12853);
and U15287 (N_15287,N_12512,N_12429);
and U15288 (N_15288,N_12336,N_13099);
and U15289 (N_15289,N_12773,N_12119);
nor U15290 (N_15290,N_13420,N_12392);
xnor U15291 (N_15291,N_12431,N_12517);
nor U15292 (N_15292,N_12251,N_13973);
or U15293 (N_15293,N_12982,N_13280);
nor U15294 (N_15294,N_12731,N_12162);
or U15295 (N_15295,N_12534,N_13055);
nor U15296 (N_15296,N_13153,N_12648);
nor U15297 (N_15297,N_13015,N_12733);
nor U15298 (N_15298,N_12690,N_12071);
nor U15299 (N_15299,N_13264,N_12050);
nand U15300 (N_15300,N_12903,N_13998);
xor U15301 (N_15301,N_12161,N_12183);
and U15302 (N_15302,N_12516,N_13043);
nand U15303 (N_15303,N_12059,N_12733);
nand U15304 (N_15304,N_12263,N_12519);
and U15305 (N_15305,N_12890,N_12937);
and U15306 (N_15306,N_13374,N_13585);
and U15307 (N_15307,N_12916,N_13043);
nand U15308 (N_15308,N_12288,N_12996);
nor U15309 (N_15309,N_12043,N_12717);
nand U15310 (N_15310,N_13902,N_12940);
xor U15311 (N_15311,N_12557,N_12741);
and U15312 (N_15312,N_12015,N_13315);
nand U15313 (N_15313,N_12092,N_12565);
or U15314 (N_15314,N_12811,N_13299);
and U15315 (N_15315,N_13739,N_13823);
or U15316 (N_15316,N_13983,N_13386);
and U15317 (N_15317,N_13400,N_13756);
nor U15318 (N_15318,N_13133,N_13094);
and U15319 (N_15319,N_12744,N_13876);
or U15320 (N_15320,N_12428,N_12082);
nand U15321 (N_15321,N_12368,N_13258);
and U15322 (N_15322,N_13011,N_13077);
nor U15323 (N_15323,N_12703,N_12121);
and U15324 (N_15324,N_12568,N_13742);
nand U15325 (N_15325,N_12401,N_12083);
nor U15326 (N_15326,N_12488,N_13363);
nor U15327 (N_15327,N_12230,N_12496);
and U15328 (N_15328,N_13924,N_12069);
or U15329 (N_15329,N_13506,N_13170);
nand U15330 (N_15330,N_13658,N_12744);
nor U15331 (N_15331,N_13156,N_12013);
nor U15332 (N_15332,N_12909,N_12087);
nor U15333 (N_15333,N_13122,N_12915);
and U15334 (N_15334,N_13395,N_12834);
or U15335 (N_15335,N_13611,N_12172);
nor U15336 (N_15336,N_12323,N_12484);
nor U15337 (N_15337,N_13749,N_12599);
or U15338 (N_15338,N_12065,N_13235);
or U15339 (N_15339,N_13947,N_13972);
nand U15340 (N_15340,N_12508,N_12729);
nand U15341 (N_15341,N_13588,N_13964);
and U15342 (N_15342,N_12008,N_12787);
xor U15343 (N_15343,N_13971,N_12664);
or U15344 (N_15344,N_12203,N_13872);
and U15345 (N_15345,N_12210,N_13369);
or U15346 (N_15346,N_12874,N_12979);
xnor U15347 (N_15347,N_12019,N_12692);
nand U15348 (N_15348,N_13759,N_13575);
or U15349 (N_15349,N_12310,N_13995);
and U15350 (N_15350,N_12717,N_13775);
nand U15351 (N_15351,N_13206,N_12855);
xor U15352 (N_15352,N_13692,N_13557);
nor U15353 (N_15353,N_12490,N_12898);
and U15354 (N_15354,N_13055,N_12845);
or U15355 (N_15355,N_13944,N_12435);
and U15356 (N_15356,N_12212,N_13945);
or U15357 (N_15357,N_13052,N_12572);
xor U15358 (N_15358,N_13539,N_12568);
and U15359 (N_15359,N_12170,N_12121);
and U15360 (N_15360,N_12951,N_13883);
and U15361 (N_15361,N_12162,N_12790);
or U15362 (N_15362,N_13488,N_13847);
nand U15363 (N_15363,N_13457,N_12686);
and U15364 (N_15364,N_12974,N_12001);
xnor U15365 (N_15365,N_13394,N_13753);
nand U15366 (N_15366,N_13410,N_13539);
nor U15367 (N_15367,N_13408,N_13661);
and U15368 (N_15368,N_13257,N_12292);
or U15369 (N_15369,N_13238,N_13848);
or U15370 (N_15370,N_12850,N_12265);
xor U15371 (N_15371,N_13696,N_13325);
or U15372 (N_15372,N_13010,N_12058);
nand U15373 (N_15373,N_13831,N_12671);
nand U15374 (N_15374,N_13913,N_12083);
and U15375 (N_15375,N_13191,N_13621);
xnor U15376 (N_15376,N_13029,N_13989);
nor U15377 (N_15377,N_12482,N_13052);
xnor U15378 (N_15378,N_12917,N_12069);
or U15379 (N_15379,N_12100,N_13461);
nand U15380 (N_15380,N_12110,N_12830);
and U15381 (N_15381,N_12977,N_12450);
nor U15382 (N_15382,N_12262,N_13252);
nor U15383 (N_15383,N_13514,N_12998);
or U15384 (N_15384,N_12945,N_12809);
nand U15385 (N_15385,N_12606,N_13904);
or U15386 (N_15386,N_13221,N_13011);
and U15387 (N_15387,N_12563,N_13363);
and U15388 (N_15388,N_13292,N_12196);
and U15389 (N_15389,N_13076,N_12317);
nor U15390 (N_15390,N_12649,N_12149);
nor U15391 (N_15391,N_12917,N_13063);
nor U15392 (N_15392,N_13026,N_13232);
xnor U15393 (N_15393,N_13099,N_12409);
or U15394 (N_15394,N_13767,N_13383);
nand U15395 (N_15395,N_13943,N_13398);
nand U15396 (N_15396,N_12651,N_13581);
and U15397 (N_15397,N_12899,N_13469);
nand U15398 (N_15398,N_13018,N_12098);
nor U15399 (N_15399,N_12566,N_12191);
xor U15400 (N_15400,N_12868,N_12065);
nand U15401 (N_15401,N_12306,N_12595);
nor U15402 (N_15402,N_12473,N_13215);
nor U15403 (N_15403,N_13473,N_13883);
and U15404 (N_15404,N_13219,N_12874);
nand U15405 (N_15405,N_12875,N_12041);
nor U15406 (N_15406,N_13684,N_12462);
or U15407 (N_15407,N_13313,N_12823);
xor U15408 (N_15408,N_12761,N_13517);
nand U15409 (N_15409,N_12097,N_13989);
nor U15410 (N_15410,N_12470,N_12028);
and U15411 (N_15411,N_12424,N_13567);
or U15412 (N_15412,N_13474,N_13375);
xnor U15413 (N_15413,N_12877,N_13428);
and U15414 (N_15414,N_12655,N_12794);
nand U15415 (N_15415,N_12924,N_12313);
nand U15416 (N_15416,N_13211,N_13914);
nor U15417 (N_15417,N_12810,N_13296);
and U15418 (N_15418,N_13283,N_12718);
xnor U15419 (N_15419,N_12763,N_13479);
or U15420 (N_15420,N_12558,N_13060);
nor U15421 (N_15421,N_12453,N_12157);
nand U15422 (N_15422,N_12135,N_13354);
or U15423 (N_15423,N_13874,N_13233);
or U15424 (N_15424,N_12825,N_13170);
xor U15425 (N_15425,N_12723,N_13011);
xor U15426 (N_15426,N_13875,N_13177);
or U15427 (N_15427,N_12135,N_13322);
and U15428 (N_15428,N_12724,N_13000);
xnor U15429 (N_15429,N_13755,N_13259);
or U15430 (N_15430,N_13611,N_13881);
nand U15431 (N_15431,N_12886,N_13820);
nand U15432 (N_15432,N_12779,N_13077);
and U15433 (N_15433,N_13290,N_12690);
and U15434 (N_15434,N_12407,N_12798);
nor U15435 (N_15435,N_12025,N_12327);
or U15436 (N_15436,N_13834,N_13700);
and U15437 (N_15437,N_13831,N_12712);
nor U15438 (N_15438,N_13904,N_13293);
or U15439 (N_15439,N_13795,N_13076);
and U15440 (N_15440,N_13214,N_12971);
nand U15441 (N_15441,N_12248,N_12033);
or U15442 (N_15442,N_12417,N_12738);
nand U15443 (N_15443,N_13822,N_12238);
nor U15444 (N_15444,N_13865,N_12615);
and U15445 (N_15445,N_13238,N_12016);
and U15446 (N_15446,N_12870,N_12750);
nand U15447 (N_15447,N_12141,N_13115);
nand U15448 (N_15448,N_12200,N_13435);
nor U15449 (N_15449,N_12519,N_12253);
or U15450 (N_15450,N_13923,N_13790);
and U15451 (N_15451,N_12427,N_13310);
nor U15452 (N_15452,N_13159,N_12477);
and U15453 (N_15453,N_13030,N_13930);
nand U15454 (N_15454,N_12484,N_13616);
nor U15455 (N_15455,N_12847,N_12346);
and U15456 (N_15456,N_13690,N_12210);
or U15457 (N_15457,N_13498,N_13431);
nand U15458 (N_15458,N_13058,N_13514);
and U15459 (N_15459,N_13054,N_13381);
nand U15460 (N_15460,N_13231,N_13859);
nor U15461 (N_15461,N_12860,N_12959);
or U15462 (N_15462,N_12140,N_12014);
or U15463 (N_15463,N_13943,N_12279);
and U15464 (N_15464,N_12187,N_12664);
or U15465 (N_15465,N_13054,N_13170);
xnor U15466 (N_15466,N_12287,N_12970);
or U15467 (N_15467,N_12369,N_13461);
nor U15468 (N_15468,N_13317,N_12581);
nand U15469 (N_15469,N_13457,N_12418);
and U15470 (N_15470,N_13209,N_12082);
xnor U15471 (N_15471,N_12303,N_13454);
and U15472 (N_15472,N_12445,N_13848);
and U15473 (N_15473,N_12649,N_13691);
nand U15474 (N_15474,N_13793,N_13155);
xor U15475 (N_15475,N_12382,N_13800);
or U15476 (N_15476,N_12226,N_13737);
nor U15477 (N_15477,N_12069,N_12696);
nand U15478 (N_15478,N_13860,N_12878);
and U15479 (N_15479,N_13279,N_13368);
nand U15480 (N_15480,N_12723,N_13102);
nor U15481 (N_15481,N_13188,N_12515);
nand U15482 (N_15482,N_13133,N_13431);
nand U15483 (N_15483,N_13562,N_12856);
or U15484 (N_15484,N_12221,N_12961);
nand U15485 (N_15485,N_13258,N_12207);
xor U15486 (N_15486,N_12222,N_13083);
nand U15487 (N_15487,N_12684,N_13493);
xnor U15488 (N_15488,N_12328,N_13740);
nand U15489 (N_15489,N_12906,N_13438);
nand U15490 (N_15490,N_12331,N_12315);
and U15491 (N_15491,N_13752,N_13003);
nor U15492 (N_15492,N_12380,N_12599);
nor U15493 (N_15493,N_12623,N_12943);
nor U15494 (N_15494,N_13373,N_13221);
and U15495 (N_15495,N_12834,N_12573);
nor U15496 (N_15496,N_12621,N_12872);
or U15497 (N_15497,N_12436,N_13299);
xor U15498 (N_15498,N_13660,N_12401);
or U15499 (N_15499,N_12942,N_13344);
nor U15500 (N_15500,N_13533,N_12802);
nand U15501 (N_15501,N_12610,N_13447);
or U15502 (N_15502,N_12685,N_13667);
and U15503 (N_15503,N_12642,N_12679);
xnor U15504 (N_15504,N_13652,N_12520);
nor U15505 (N_15505,N_12757,N_12152);
nor U15506 (N_15506,N_12427,N_13956);
or U15507 (N_15507,N_13183,N_12505);
or U15508 (N_15508,N_12869,N_13295);
nor U15509 (N_15509,N_12591,N_13455);
or U15510 (N_15510,N_12711,N_12736);
xnor U15511 (N_15511,N_13476,N_13432);
xnor U15512 (N_15512,N_12916,N_12470);
and U15513 (N_15513,N_13093,N_13915);
and U15514 (N_15514,N_12844,N_13569);
nand U15515 (N_15515,N_13671,N_13237);
nor U15516 (N_15516,N_12453,N_13306);
or U15517 (N_15517,N_13641,N_12515);
nor U15518 (N_15518,N_12942,N_13480);
nand U15519 (N_15519,N_13554,N_12954);
and U15520 (N_15520,N_12612,N_12027);
and U15521 (N_15521,N_12643,N_13197);
and U15522 (N_15522,N_13429,N_12958);
nand U15523 (N_15523,N_12780,N_12345);
nand U15524 (N_15524,N_13085,N_13770);
nand U15525 (N_15525,N_12772,N_13844);
and U15526 (N_15526,N_12153,N_12480);
nor U15527 (N_15527,N_12323,N_13587);
or U15528 (N_15528,N_12082,N_13108);
and U15529 (N_15529,N_13929,N_12609);
or U15530 (N_15530,N_12437,N_12127);
and U15531 (N_15531,N_12247,N_12264);
nor U15532 (N_15532,N_12157,N_13223);
and U15533 (N_15533,N_12633,N_12278);
nand U15534 (N_15534,N_12990,N_12669);
nand U15535 (N_15535,N_13476,N_12224);
nand U15536 (N_15536,N_12220,N_12812);
or U15537 (N_15537,N_12934,N_12957);
and U15538 (N_15538,N_12216,N_12095);
nor U15539 (N_15539,N_13093,N_13639);
nor U15540 (N_15540,N_12604,N_13051);
nand U15541 (N_15541,N_12244,N_13757);
or U15542 (N_15542,N_13982,N_13228);
nand U15543 (N_15543,N_12584,N_13620);
or U15544 (N_15544,N_13807,N_12385);
or U15545 (N_15545,N_12497,N_12056);
nand U15546 (N_15546,N_13280,N_12610);
and U15547 (N_15547,N_13299,N_12051);
or U15548 (N_15548,N_13020,N_12672);
nor U15549 (N_15549,N_13009,N_12939);
or U15550 (N_15550,N_12658,N_13402);
nor U15551 (N_15551,N_12553,N_12120);
and U15552 (N_15552,N_13150,N_13085);
and U15553 (N_15553,N_12525,N_13608);
nor U15554 (N_15554,N_13753,N_12090);
nor U15555 (N_15555,N_13779,N_13392);
nor U15556 (N_15556,N_12309,N_13587);
nor U15557 (N_15557,N_13513,N_13499);
nand U15558 (N_15558,N_12628,N_13148);
nor U15559 (N_15559,N_13272,N_13337);
xnor U15560 (N_15560,N_13990,N_12427);
and U15561 (N_15561,N_12712,N_12627);
nor U15562 (N_15562,N_12585,N_13898);
or U15563 (N_15563,N_13077,N_12445);
nand U15564 (N_15564,N_12195,N_12004);
nand U15565 (N_15565,N_12052,N_13292);
nor U15566 (N_15566,N_13310,N_12827);
xor U15567 (N_15567,N_13222,N_12745);
nor U15568 (N_15568,N_13327,N_13063);
and U15569 (N_15569,N_13973,N_12153);
or U15570 (N_15570,N_13049,N_13088);
or U15571 (N_15571,N_13355,N_12821);
nand U15572 (N_15572,N_13698,N_13760);
nor U15573 (N_15573,N_12349,N_13688);
xor U15574 (N_15574,N_12886,N_13920);
and U15575 (N_15575,N_12769,N_12452);
nand U15576 (N_15576,N_12272,N_13486);
nor U15577 (N_15577,N_12150,N_13644);
and U15578 (N_15578,N_13789,N_12723);
or U15579 (N_15579,N_12130,N_13388);
nor U15580 (N_15580,N_12760,N_12033);
xor U15581 (N_15581,N_13174,N_12749);
nand U15582 (N_15582,N_12970,N_13926);
nor U15583 (N_15583,N_12169,N_12211);
nor U15584 (N_15584,N_13029,N_13515);
or U15585 (N_15585,N_13353,N_13900);
or U15586 (N_15586,N_13649,N_13043);
and U15587 (N_15587,N_13231,N_12096);
nor U15588 (N_15588,N_12751,N_12691);
nand U15589 (N_15589,N_13210,N_12273);
nor U15590 (N_15590,N_12454,N_13814);
nand U15591 (N_15591,N_12338,N_12850);
nor U15592 (N_15592,N_12332,N_12723);
xor U15593 (N_15593,N_13843,N_12231);
xor U15594 (N_15594,N_13116,N_12801);
and U15595 (N_15595,N_12386,N_13086);
nor U15596 (N_15596,N_13341,N_12087);
or U15597 (N_15597,N_13467,N_13063);
and U15598 (N_15598,N_13314,N_12827);
and U15599 (N_15599,N_12967,N_13137);
and U15600 (N_15600,N_13958,N_13441);
or U15601 (N_15601,N_13575,N_13229);
nand U15602 (N_15602,N_13453,N_13161);
and U15603 (N_15603,N_12503,N_13899);
or U15604 (N_15604,N_13401,N_13675);
nor U15605 (N_15605,N_13985,N_13760);
or U15606 (N_15606,N_13848,N_12020);
and U15607 (N_15607,N_12680,N_13452);
and U15608 (N_15608,N_13491,N_12661);
or U15609 (N_15609,N_13662,N_13815);
nor U15610 (N_15610,N_13115,N_12382);
nor U15611 (N_15611,N_12944,N_13411);
or U15612 (N_15612,N_12072,N_12533);
nand U15613 (N_15613,N_12720,N_12222);
nand U15614 (N_15614,N_13834,N_13740);
nand U15615 (N_15615,N_12090,N_13953);
or U15616 (N_15616,N_13425,N_13238);
and U15617 (N_15617,N_13667,N_13412);
and U15618 (N_15618,N_13584,N_12699);
nor U15619 (N_15619,N_12624,N_12190);
and U15620 (N_15620,N_12162,N_13342);
xnor U15621 (N_15621,N_13334,N_12491);
nor U15622 (N_15622,N_12973,N_12392);
nor U15623 (N_15623,N_12605,N_12683);
nor U15624 (N_15624,N_12960,N_13983);
nor U15625 (N_15625,N_12379,N_12866);
and U15626 (N_15626,N_13217,N_13738);
nand U15627 (N_15627,N_12050,N_12858);
or U15628 (N_15628,N_12627,N_13518);
and U15629 (N_15629,N_12639,N_12433);
nor U15630 (N_15630,N_12725,N_12202);
nor U15631 (N_15631,N_13712,N_12970);
and U15632 (N_15632,N_13157,N_12336);
and U15633 (N_15633,N_13598,N_13916);
nand U15634 (N_15634,N_13929,N_13315);
nand U15635 (N_15635,N_13574,N_12264);
and U15636 (N_15636,N_12288,N_12363);
nand U15637 (N_15637,N_13601,N_12276);
or U15638 (N_15638,N_12704,N_13625);
xor U15639 (N_15639,N_13493,N_12495);
xor U15640 (N_15640,N_12615,N_13379);
and U15641 (N_15641,N_12747,N_12051);
nor U15642 (N_15642,N_12951,N_13577);
nand U15643 (N_15643,N_12995,N_13741);
or U15644 (N_15644,N_13483,N_13976);
or U15645 (N_15645,N_12568,N_12242);
nand U15646 (N_15646,N_13740,N_13065);
xor U15647 (N_15647,N_13085,N_13740);
nor U15648 (N_15648,N_12567,N_13968);
or U15649 (N_15649,N_13101,N_13649);
or U15650 (N_15650,N_13686,N_13714);
nand U15651 (N_15651,N_12132,N_13058);
nor U15652 (N_15652,N_13409,N_13690);
nor U15653 (N_15653,N_13268,N_12005);
nand U15654 (N_15654,N_12115,N_12613);
nor U15655 (N_15655,N_12731,N_13537);
nor U15656 (N_15656,N_13747,N_12718);
and U15657 (N_15657,N_13208,N_12203);
and U15658 (N_15658,N_13116,N_13540);
nor U15659 (N_15659,N_13777,N_13072);
and U15660 (N_15660,N_12040,N_13835);
nand U15661 (N_15661,N_12822,N_12810);
xnor U15662 (N_15662,N_13603,N_12048);
nand U15663 (N_15663,N_12322,N_13201);
nand U15664 (N_15664,N_13966,N_12317);
nor U15665 (N_15665,N_13096,N_13518);
or U15666 (N_15666,N_13104,N_12397);
or U15667 (N_15667,N_13149,N_13480);
and U15668 (N_15668,N_12952,N_13586);
and U15669 (N_15669,N_13368,N_12246);
and U15670 (N_15670,N_12607,N_13899);
or U15671 (N_15671,N_13386,N_12338);
nor U15672 (N_15672,N_12655,N_12484);
or U15673 (N_15673,N_12842,N_13407);
and U15674 (N_15674,N_13944,N_12352);
nand U15675 (N_15675,N_13915,N_13713);
xnor U15676 (N_15676,N_13376,N_13721);
or U15677 (N_15677,N_12741,N_13257);
nor U15678 (N_15678,N_12651,N_12205);
and U15679 (N_15679,N_12173,N_13106);
and U15680 (N_15680,N_13023,N_12681);
or U15681 (N_15681,N_12054,N_13104);
nand U15682 (N_15682,N_13486,N_13611);
nand U15683 (N_15683,N_12203,N_12997);
nand U15684 (N_15684,N_12384,N_13032);
nor U15685 (N_15685,N_12535,N_12637);
or U15686 (N_15686,N_13517,N_13601);
nor U15687 (N_15687,N_13373,N_13011);
nand U15688 (N_15688,N_13070,N_13716);
xnor U15689 (N_15689,N_12699,N_12279);
or U15690 (N_15690,N_12947,N_12435);
and U15691 (N_15691,N_13585,N_12228);
and U15692 (N_15692,N_12823,N_13596);
or U15693 (N_15693,N_13175,N_12055);
nand U15694 (N_15694,N_12357,N_12982);
or U15695 (N_15695,N_13255,N_12595);
or U15696 (N_15696,N_12648,N_13134);
and U15697 (N_15697,N_13080,N_12112);
and U15698 (N_15698,N_13939,N_12782);
nor U15699 (N_15699,N_13502,N_12769);
nor U15700 (N_15700,N_13863,N_13351);
nor U15701 (N_15701,N_12380,N_13249);
and U15702 (N_15702,N_12650,N_13141);
xnor U15703 (N_15703,N_12803,N_12189);
nor U15704 (N_15704,N_13268,N_13233);
nand U15705 (N_15705,N_13197,N_13061);
nand U15706 (N_15706,N_13609,N_13784);
or U15707 (N_15707,N_13444,N_13347);
xnor U15708 (N_15708,N_13429,N_12908);
nor U15709 (N_15709,N_12368,N_12382);
nand U15710 (N_15710,N_12423,N_12874);
and U15711 (N_15711,N_12829,N_12008);
nor U15712 (N_15712,N_12515,N_12997);
xnor U15713 (N_15713,N_13714,N_13112);
nor U15714 (N_15714,N_13049,N_13789);
nand U15715 (N_15715,N_12160,N_12810);
and U15716 (N_15716,N_12000,N_13788);
nor U15717 (N_15717,N_13933,N_12115);
nand U15718 (N_15718,N_13029,N_13184);
nand U15719 (N_15719,N_12181,N_12763);
xor U15720 (N_15720,N_12584,N_13282);
and U15721 (N_15721,N_12973,N_12231);
and U15722 (N_15722,N_13903,N_13715);
or U15723 (N_15723,N_13847,N_13347);
nand U15724 (N_15724,N_13578,N_13778);
nand U15725 (N_15725,N_12326,N_12915);
and U15726 (N_15726,N_12937,N_13985);
nand U15727 (N_15727,N_13913,N_13375);
or U15728 (N_15728,N_13738,N_13342);
xor U15729 (N_15729,N_13730,N_13471);
nor U15730 (N_15730,N_12278,N_13001);
nor U15731 (N_15731,N_12626,N_13699);
nand U15732 (N_15732,N_12340,N_12405);
or U15733 (N_15733,N_13905,N_13385);
and U15734 (N_15734,N_12832,N_12044);
nand U15735 (N_15735,N_13456,N_13187);
nand U15736 (N_15736,N_13188,N_13748);
xnor U15737 (N_15737,N_13997,N_13264);
nor U15738 (N_15738,N_13319,N_13087);
xnor U15739 (N_15739,N_13024,N_12593);
nor U15740 (N_15740,N_12492,N_12595);
nand U15741 (N_15741,N_13406,N_13666);
nor U15742 (N_15742,N_13484,N_13786);
or U15743 (N_15743,N_13694,N_12347);
nor U15744 (N_15744,N_13926,N_12137);
nand U15745 (N_15745,N_12120,N_12893);
and U15746 (N_15746,N_12002,N_13850);
and U15747 (N_15747,N_13410,N_12251);
or U15748 (N_15748,N_12204,N_13463);
xor U15749 (N_15749,N_13509,N_13032);
and U15750 (N_15750,N_13428,N_12310);
nand U15751 (N_15751,N_13862,N_12269);
or U15752 (N_15752,N_12022,N_12259);
and U15753 (N_15753,N_12863,N_13723);
or U15754 (N_15754,N_13735,N_12781);
xnor U15755 (N_15755,N_12759,N_12190);
nor U15756 (N_15756,N_13580,N_13458);
nand U15757 (N_15757,N_12014,N_12929);
and U15758 (N_15758,N_12254,N_13795);
nand U15759 (N_15759,N_12509,N_13912);
nor U15760 (N_15760,N_12153,N_13731);
xnor U15761 (N_15761,N_12802,N_13198);
xor U15762 (N_15762,N_13071,N_13537);
or U15763 (N_15763,N_13250,N_12961);
nand U15764 (N_15764,N_13822,N_13595);
nor U15765 (N_15765,N_12241,N_13292);
nor U15766 (N_15766,N_12722,N_12930);
and U15767 (N_15767,N_12841,N_12138);
and U15768 (N_15768,N_13339,N_13455);
and U15769 (N_15769,N_12455,N_13591);
or U15770 (N_15770,N_13042,N_13019);
or U15771 (N_15771,N_13667,N_12647);
nand U15772 (N_15772,N_12987,N_13615);
or U15773 (N_15773,N_12628,N_12934);
and U15774 (N_15774,N_13089,N_13139);
or U15775 (N_15775,N_12139,N_13264);
nor U15776 (N_15776,N_12741,N_13934);
and U15777 (N_15777,N_13975,N_12510);
nor U15778 (N_15778,N_12055,N_12399);
or U15779 (N_15779,N_13347,N_12331);
nand U15780 (N_15780,N_13933,N_13665);
nor U15781 (N_15781,N_13958,N_12289);
nor U15782 (N_15782,N_13978,N_12900);
or U15783 (N_15783,N_12261,N_12030);
nand U15784 (N_15784,N_13904,N_13179);
or U15785 (N_15785,N_12138,N_12578);
nor U15786 (N_15786,N_12957,N_13207);
nor U15787 (N_15787,N_12666,N_13824);
nand U15788 (N_15788,N_12254,N_12735);
or U15789 (N_15789,N_12798,N_13683);
nor U15790 (N_15790,N_12619,N_12104);
and U15791 (N_15791,N_13320,N_12013);
nor U15792 (N_15792,N_13180,N_13282);
or U15793 (N_15793,N_13481,N_13612);
nand U15794 (N_15794,N_12664,N_13648);
nor U15795 (N_15795,N_12119,N_13731);
nor U15796 (N_15796,N_12353,N_12712);
and U15797 (N_15797,N_12368,N_13321);
nand U15798 (N_15798,N_13994,N_13362);
nand U15799 (N_15799,N_12482,N_12808);
or U15800 (N_15800,N_13404,N_13899);
or U15801 (N_15801,N_12559,N_12943);
nor U15802 (N_15802,N_13588,N_12687);
and U15803 (N_15803,N_12529,N_13852);
nor U15804 (N_15804,N_13536,N_12477);
and U15805 (N_15805,N_12118,N_12187);
xnor U15806 (N_15806,N_13960,N_13804);
or U15807 (N_15807,N_13497,N_12746);
or U15808 (N_15808,N_13696,N_12917);
nand U15809 (N_15809,N_12335,N_12820);
nor U15810 (N_15810,N_13832,N_12185);
or U15811 (N_15811,N_12795,N_12778);
nand U15812 (N_15812,N_13026,N_13520);
and U15813 (N_15813,N_12573,N_12256);
and U15814 (N_15814,N_12503,N_12394);
or U15815 (N_15815,N_13576,N_12290);
xnor U15816 (N_15816,N_12948,N_12391);
nand U15817 (N_15817,N_13779,N_12180);
nand U15818 (N_15818,N_12163,N_12563);
nand U15819 (N_15819,N_12319,N_13263);
nand U15820 (N_15820,N_12484,N_12571);
or U15821 (N_15821,N_13243,N_13488);
and U15822 (N_15822,N_12774,N_13704);
nand U15823 (N_15823,N_12425,N_13169);
nand U15824 (N_15824,N_13600,N_13473);
or U15825 (N_15825,N_13114,N_13967);
nand U15826 (N_15826,N_13928,N_12735);
nor U15827 (N_15827,N_13744,N_12882);
nor U15828 (N_15828,N_12467,N_12902);
or U15829 (N_15829,N_13167,N_13505);
and U15830 (N_15830,N_13344,N_13655);
and U15831 (N_15831,N_13104,N_12426);
and U15832 (N_15832,N_13216,N_13541);
and U15833 (N_15833,N_12893,N_12890);
nand U15834 (N_15834,N_12107,N_13831);
or U15835 (N_15835,N_12292,N_13571);
nand U15836 (N_15836,N_13741,N_12693);
nor U15837 (N_15837,N_13695,N_12986);
nand U15838 (N_15838,N_12884,N_13839);
nor U15839 (N_15839,N_13178,N_12372);
or U15840 (N_15840,N_12194,N_13023);
and U15841 (N_15841,N_12429,N_12265);
nor U15842 (N_15842,N_13097,N_13589);
or U15843 (N_15843,N_12851,N_12546);
nand U15844 (N_15844,N_13986,N_12288);
or U15845 (N_15845,N_13925,N_12784);
and U15846 (N_15846,N_12328,N_12253);
or U15847 (N_15847,N_12223,N_12957);
or U15848 (N_15848,N_12352,N_12727);
nand U15849 (N_15849,N_12369,N_13638);
or U15850 (N_15850,N_13706,N_12782);
nor U15851 (N_15851,N_13995,N_12056);
and U15852 (N_15852,N_12498,N_13050);
or U15853 (N_15853,N_12915,N_12849);
and U15854 (N_15854,N_13938,N_12484);
nand U15855 (N_15855,N_12733,N_13980);
nor U15856 (N_15856,N_13299,N_12281);
nor U15857 (N_15857,N_13835,N_13424);
and U15858 (N_15858,N_13528,N_13839);
nor U15859 (N_15859,N_13097,N_13940);
nand U15860 (N_15860,N_12744,N_12773);
or U15861 (N_15861,N_13675,N_12204);
nand U15862 (N_15862,N_12739,N_12946);
nor U15863 (N_15863,N_13747,N_13213);
and U15864 (N_15864,N_12708,N_12554);
nor U15865 (N_15865,N_12956,N_13031);
nor U15866 (N_15866,N_13526,N_13944);
nor U15867 (N_15867,N_13065,N_12253);
or U15868 (N_15868,N_12757,N_13631);
or U15869 (N_15869,N_12301,N_12563);
and U15870 (N_15870,N_12200,N_12261);
and U15871 (N_15871,N_13454,N_13872);
and U15872 (N_15872,N_12001,N_12905);
nor U15873 (N_15873,N_13414,N_13348);
nor U15874 (N_15874,N_13403,N_13853);
and U15875 (N_15875,N_13882,N_13738);
and U15876 (N_15876,N_13288,N_12411);
and U15877 (N_15877,N_13168,N_12923);
and U15878 (N_15878,N_12242,N_13880);
or U15879 (N_15879,N_12806,N_12900);
nor U15880 (N_15880,N_13629,N_13582);
or U15881 (N_15881,N_13090,N_12290);
and U15882 (N_15882,N_12916,N_12095);
and U15883 (N_15883,N_13192,N_13162);
nand U15884 (N_15884,N_12065,N_12502);
nand U15885 (N_15885,N_13670,N_13854);
or U15886 (N_15886,N_13236,N_13774);
and U15887 (N_15887,N_12730,N_13211);
nand U15888 (N_15888,N_12830,N_12065);
nand U15889 (N_15889,N_12048,N_12715);
nor U15890 (N_15890,N_13345,N_12347);
nor U15891 (N_15891,N_12641,N_12204);
and U15892 (N_15892,N_13060,N_13371);
and U15893 (N_15893,N_12907,N_12393);
and U15894 (N_15894,N_13050,N_13300);
nand U15895 (N_15895,N_13382,N_12375);
and U15896 (N_15896,N_13248,N_13745);
nor U15897 (N_15897,N_12541,N_13982);
nand U15898 (N_15898,N_13147,N_13122);
or U15899 (N_15899,N_12827,N_13086);
or U15900 (N_15900,N_13494,N_13713);
nand U15901 (N_15901,N_13827,N_12288);
nor U15902 (N_15902,N_12678,N_13740);
nand U15903 (N_15903,N_12301,N_13796);
nor U15904 (N_15904,N_13622,N_13753);
nand U15905 (N_15905,N_13689,N_13808);
and U15906 (N_15906,N_13002,N_13543);
nor U15907 (N_15907,N_12816,N_12517);
nor U15908 (N_15908,N_13581,N_13634);
and U15909 (N_15909,N_12745,N_13197);
nor U15910 (N_15910,N_12508,N_13535);
or U15911 (N_15911,N_13316,N_12489);
or U15912 (N_15912,N_13001,N_13669);
nand U15913 (N_15913,N_13439,N_12340);
xnor U15914 (N_15914,N_13208,N_13859);
and U15915 (N_15915,N_13744,N_13334);
nand U15916 (N_15916,N_12676,N_12497);
and U15917 (N_15917,N_13531,N_12432);
nand U15918 (N_15918,N_12613,N_12429);
and U15919 (N_15919,N_12709,N_12725);
nor U15920 (N_15920,N_12206,N_13544);
nand U15921 (N_15921,N_13746,N_12575);
and U15922 (N_15922,N_13154,N_13832);
nand U15923 (N_15923,N_12653,N_12976);
and U15924 (N_15924,N_13360,N_12990);
nand U15925 (N_15925,N_12722,N_12406);
nand U15926 (N_15926,N_13709,N_13718);
and U15927 (N_15927,N_12310,N_13986);
xnor U15928 (N_15928,N_13856,N_12847);
nand U15929 (N_15929,N_12342,N_12375);
xor U15930 (N_15930,N_13198,N_12641);
or U15931 (N_15931,N_12934,N_13602);
or U15932 (N_15932,N_12656,N_12617);
xor U15933 (N_15933,N_12395,N_12531);
and U15934 (N_15934,N_12724,N_13925);
or U15935 (N_15935,N_13612,N_13849);
nor U15936 (N_15936,N_12176,N_12099);
nand U15937 (N_15937,N_12240,N_12778);
nor U15938 (N_15938,N_13245,N_12904);
and U15939 (N_15939,N_12192,N_13699);
nand U15940 (N_15940,N_13384,N_12862);
nand U15941 (N_15941,N_13223,N_12983);
and U15942 (N_15942,N_12027,N_12053);
nand U15943 (N_15943,N_13411,N_12968);
nor U15944 (N_15944,N_12420,N_13661);
nand U15945 (N_15945,N_12983,N_12196);
nor U15946 (N_15946,N_13857,N_13183);
nand U15947 (N_15947,N_13957,N_12578);
nand U15948 (N_15948,N_12127,N_13140);
xor U15949 (N_15949,N_13498,N_13357);
or U15950 (N_15950,N_13912,N_12002);
and U15951 (N_15951,N_12167,N_13793);
or U15952 (N_15952,N_12440,N_13993);
or U15953 (N_15953,N_12547,N_12092);
and U15954 (N_15954,N_13312,N_12492);
nor U15955 (N_15955,N_12060,N_12312);
nand U15956 (N_15956,N_13172,N_12791);
nand U15957 (N_15957,N_13018,N_13891);
nand U15958 (N_15958,N_13391,N_12476);
or U15959 (N_15959,N_12249,N_13311);
nand U15960 (N_15960,N_13324,N_13822);
nand U15961 (N_15961,N_12140,N_12428);
and U15962 (N_15962,N_13459,N_12563);
and U15963 (N_15963,N_12472,N_12861);
nor U15964 (N_15964,N_12464,N_13794);
and U15965 (N_15965,N_12572,N_13018);
and U15966 (N_15966,N_13314,N_13628);
and U15967 (N_15967,N_13231,N_12465);
and U15968 (N_15968,N_13987,N_13022);
xnor U15969 (N_15969,N_13260,N_13045);
and U15970 (N_15970,N_13566,N_13226);
nor U15971 (N_15971,N_13057,N_13870);
nor U15972 (N_15972,N_13052,N_12770);
and U15973 (N_15973,N_12602,N_13620);
or U15974 (N_15974,N_12478,N_13589);
and U15975 (N_15975,N_13506,N_12258);
and U15976 (N_15976,N_12305,N_13870);
nor U15977 (N_15977,N_12966,N_13478);
and U15978 (N_15978,N_12124,N_13993);
nand U15979 (N_15979,N_13880,N_13637);
xor U15980 (N_15980,N_12547,N_12568);
nor U15981 (N_15981,N_12245,N_12051);
and U15982 (N_15982,N_13987,N_13613);
and U15983 (N_15983,N_12893,N_12984);
nand U15984 (N_15984,N_12227,N_13267);
and U15985 (N_15985,N_12051,N_12004);
and U15986 (N_15986,N_13018,N_13550);
xor U15987 (N_15987,N_12038,N_12068);
nand U15988 (N_15988,N_13730,N_13425);
or U15989 (N_15989,N_12752,N_12270);
or U15990 (N_15990,N_13850,N_12233);
or U15991 (N_15991,N_13229,N_13762);
or U15992 (N_15992,N_13855,N_13068);
nand U15993 (N_15993,N_12448,N_13262);
nor U15994 (N_15994,N_12504,N_12163);
nand U15995 (N_15995,N_12640,N_13118);
nor U15996 (N_15996,N_13513,N_13114);
nor U15997 (N_15997,N_13498,N_13288);
nor U15998 (N_15998,N_12991,N_13089);
nand U15999 (N_15999,N_12468,N_13618);
or U16000 (N_16000,N_14147,N_15546);
nand U16001 (N_16001,N_15903,N_14214);
or U16002 (N_16002,N_14884,N_14888);
nor U16003 (N_16003,N_14278,N_15327);
or U16004 (N_16004,N_15131,N_15181);
nand U16005 (N_16005,N_15890,N_15739);
xor U16006 (N_16006,N_14657,N_15977);
nor U16007 (N_16007,N_14731,N_15435);
nand U16008 (N_16008,N_15606,N_14634);
nand U16009 (N_16009,N_14937,N_14822);
xnor U16010 (N_16010,N_15270,N_14406);
or U16011 (N_16011,N_15526,N_14067);
and U16012 (N_16012,N_15990,N_14985);
nor U16013 (N_16013,N_14475,N_14956);
nand U16014 (N_16014,N_15792,N_14850);
or U16015 (N_16015,N_14322,N_15169);
nor U16016 (N_16016,N_15483,N_14839);
nor U16017 (N_16017,N_14802,N_14295);
nor U16018 (N_16018,N_14829,N_14766);
nand U16019 (N_16019,N_14751,N_15778);
nor U16020 (N_16020,N_15039,N_15138);
or U16021 (N_16021,N_14800,N_14757);
or U16022 (N_16022,N_14338,N_15186);
nand U16023 (N_16023,N_15204,N_15048);
nand U16024 (N_16024,N_15611,N_15057);
and U16025 (N_16025,N_15948,N_15667);
nor U16026 (N_16026,N_14479,N_14177);
xor U16027 (N_16027,N_14448,N_14717);
nor U16028 (N_16028,N_15498,N_14876);
nor U16029 (N_16029,N_15297,N_15929);
nor U16030 (N_16030,N_15295,N_14249);
or U16031 (N_16031,N_14814,N_15146);
or U16032 (N_16032,N_14105,N_15422);
or U16033 (N_16033,N_15830,N_14698);
xnor U16034 (N_16034,N_15527,N_15097);
and U16035 (N_16035,N_14920,N_15343);
nor U16036 (N_16036,N_14509,N_15868);
or U16037 (N_16037,N_14846,N_15394);
and U16038 (N_16038,N_15877,N_15371);
and U16039 (N_16039,N_15376,N_14723);
and U16040 (N_16040,N_14579,N_15631);
or U16041 (N_16041,N_15214,N_15060);
nand U16042 (N_16042,N_14611,N_14510);
nor U16043 (N_16043,N_14988,N_15587);
nand U16044 (N_16044,N_14117,N_15361);
or U16045 (N_16045,N_14217,N_15025);
xnor U16046 (N_16046,N_14298,N_14445);
nand U16047 (N_16047,N_14020,N_14960);
or U16048 (N_16048,N_15853,N_15370);
nand U16049 (N_16049,N_15628,N_14618);
nand U16050 (N_16050,N_14676,N_14438);
nand U16051 (N_16051,N_15570,N_14423);
and U16052 (N_16052,N_15934,N_15878);
nor U16053 (N_16053,N_14111,N_15659);
and U16054 (N_16054,N_14564,N_15232);
and U16055 (N_16055,N_14941,N_14928);
nand U16056 (N_16056,N_15721,N_14155);
and U16057 (N_16057,N_15734,N_15260);
nor U16058 (N_16058,N_14234,N_15342);
nor U16059 (N_16059,N_15391,N_15231);
xnor U16060 (N_16060,N_14507,N_15378);
nand U16061 (N_16061,N_14193,N_15574);
nor U16062 (N_16062,N_15471,N_14806);
or U16063 (N_16063,N_14545,N_14135);
nand U16064 (N_16064,N_14011,N_14963);
or U16065 (N_16065,N_15530,N_14452);
and U16066 (N_16066,N_14134,N_15261);
xnor U16067 (N_16067,N_14205,N_15512);
nor U16068 (N_16068,N_14550,N_15700);
nand U16069 (N_16069,N_14354,N_15078);
nand U16070 (N_16070,N_14840,N_14774);
nor U16071 (N_16071,N_14022,N_15499);
nand U16072 (N_16072,N_15054,N_15951);
and U16073 (N_16073,N_15363,N_14576);
and U16074 (N_16074,N_14952,N_14054);
nand U16075 (N_16075,N_15180,N_15855);
nand U16076 (N_16076,N_14772,N_14997);
xnor U16077 (N_16077,N_15485,N_14252);
or U16078 (N_16078,N_15461,N_15199);
and U16079 (N_16079,N_15106,N_14262);
or U16080 (N_16080,N_14454,N_14266);
nand U16081 (N_16081,N_15945,N_15018);
or U16082 (N_16082,N_15718,N_15635);
nor U16083 (N_16083,N_15793,N_15848);
nor U16084 (N_16084,N_15589,N_14014);
nor U16085 (N_16085,N_15197,N_15629);
nand U16086 (N_16086,N_15685,N_15641);
nor U16087 (N_16087,N_14531,N_15007);
xnor U16088 (N_16088,N_14444,N_14594);
nor U16089 (N_16089,N_14514,N_15266);
nor U16090 (N_16090,N_15906,N_14484);
and U16091 (N_16091,N_15864,N_15742);
nor U16092 (N_16092,N_14754,N_15531);
nor U16093 (N_16093,N_14967,N_15909);
or U16094 (N_16094,N_15460,N_15006);
nand U16095 (N_16095,N_15768,N_15593);
nand U16096 (N_16096,N_14505,N_15428);
nand U16097 (N_16097,N_15745,N_14572);
and U16098 (N_16098,N_14440,N_14512);
nor U16099 (N_16099,N_15086,N_15744);
or U16100 (N_16100,N_14647,N_15710);
nor U16101 (N_16101,N_15856,N_15735);
or U16102 (N_16102,N_15096,N_14525);
or U16103 (N_16103,N_14144,N_15074);
and U16104 (N_16104,N_14705,N_14108);
and U16105 (N_16105,N_14090,N_15623);
nor U16106 (N_16106,N_14037,N_14598);
and U16107 (N_16107,N_15296,N_15427);
or U16108 (N_16108,N_14778,N_14142);
nor U16109 (N_16109,N_14902,N_15813);
nand U16110 (N_16110,N_14750,N_15646);
and U16111 (N_16111,N_15999,N_14255);
and U16112 (N_16112,N_14974,N_14568);
xnor U16113 (N_16113,N_15365,N_14330);
nand U16114 (N_16114,N_14785,N_15016);
nand U16115 (N_16115,N_14652,N_15368);
or U16116 (N_16116,N_14360,N_15668);
nor U16117 (N_16117,N_14958,N_14442);
and U16118 (N_16118,N_14743,N_15725);
nand U16119 (N_16119,N_15761,N_14752);
nor U16120 (N_16120,N_14885,N_15211);
xor U16121 (N_16121,N_15438,N_14701);
or U16122 (N_16122,N_14028,N_14064);
xnor U16123 (N_16123,N_15382,N_15580);
nand U16124 (N_16124,N_15733,N_14995);
and U16125 (N_16125,N_14461,N_15783);
nand U16126 (N_16126,N_14321,N_14350);
nand U16127 (N_16127,N_15294,N_15695);
nand U16128 (N_16128,N_15669,N_15496);
nand U16129 (N_16129,N_15168,N_14975);
nor U16130 (N_16130,N_15612,N_14399);
nand U16131 (N_16131,N_14110,N_14990);
xor U16132 (N_16132,N_14908,N_14327);
xor U16133 (N_16133,N_14714,N_15504);
nand U16134 (N_16134,N_14502,N_15865);
and U16135 (N_16135,N_15277,N_15741);
and U16136 (N_16136,N_14021,N_14845);
nand U16137 (N_16137,N_14381,N_15189);
nand U16138 (N_16138,N_14793,N_14097);
nand U16139 (N_16139,N_15577,N_15156);
nand U16140 (N_16140,N_15916,N_15280);
nand U16141 (N_16141,N_15300,N_14630);
nor U16142 (N_16142,N_14347,N_15474);
and U16143 (N_16143,N_15366,N_14182);
nand U16144 (N_16144,N_14733,N_15203);
nor U16145 (N_16145,N_14642,N_14194);
nand U16146 (N_16146,N_14981,N_14922);
and U16147 (N_16147,N_15278,N_14398);
or U16148 (N_16148,N_15308,N_15046);
nand U16149 (N_16149,N_15773,N_15448);
and U16150 (N_16150,N_15135,N_15482);
and U16151 (N_16151,N_15047,N_15249);
nand U16152 (N_16152,N_14312,N_14465);
nor U16153 (N_16153,N_15544,N_15900);
nand U16154 (N_16154,N_15979,N_15267);
and U16155 (N_16155,N_14259,N_15652);
nor U16156 (N_16156,N_14878,N_14092);
or U16157 (N_16157,N_14817,N_15055);
nand U16158 (N_16158,N_15080,N_14462);
nor U16159 (N_16159,N_14538,N_14270);
and U16160 (N_16160,N_15191,N_14866);
and U16161 (N_16161,N_15236,N_15320);
nand U16162 (N_16162,N_15235,N_15809);
xnor U16163 (N_16163,N_15633,N_14547);
and U16164 (N_16164,N_15045,N_14362);
nand U16165 (N_16165,N_15289,N_15299);
nand U16166 (N_16166,N_14668,N_14279);
and U16167 (N_16167,N_14719,N_14856);
or U16168 (N_16168,N_15345,N_14775);
and U16169 (N_16169,N_15497,N_14269);
or U16170 (N_16170,N_14086,N_14666);
and U16171 (N_16171,N_14318,N_14732);
or U16172 (N_16172,N_14371,N_14585);
nor U16173 (N_16173,N_14116,N_14424);
or U16174 (N_16174,N_14834,N_15473);
or U16175 (N_16175,N_15147,N_15693);
nor U16176 (N_16176,N_15712,N_14546);
or U16177 (N_16177,N_15584,N_14190);
or U16178 (N_16178,N_14365,N_14250);
nand U16179 (N_16179,N_14632,N_14992);
nand U16180 (N_16180,N_15233,N_15244);
or U16181 (N_16181,N_14284,N_15711);
xor U16182 (N_16182,N_15247,N_15442);
nand U16183 (N_16183,N_15753,N_15804);
nor U16184 (N_16184,N_14175,N_14358);
or U16185 (N_16185,N_15516,N_15901);
and U16186 (N_16186,N_14690,N_14784);
xnor U16187 (N_16187,N_15796,N_14515);
nand U16188 (N_16188,N_14535,N_14712);
and U16189 (N_16189,N_15918,N_14604);
nor U16190 (N_16190,N_15701,N_15409);
nor U16191 (N_16191,N_14374,N_14746);
nand U16192 (N_16192,N_15936,N_14847);
nand U16193 (N_16193,N_14246,N_15515);
nand U16194 (N_16194,N_14953,N_15940);
and U16195 (N_16195,N_15317,N_14897);
nor U16196 (N_16196,N_14661,N_15806);
and U16197 (N_16197,N_14708,N_15256);
nand U16198 (N_16198,N_14835,N_15785);
nor U16199 (N_16199,N_15692,N_15167);
nor U16200 (N_16200,N_14921,N_15784);
and U16201 (N_16201,N_14797,N_14879);
xor U16202 (N_16202,N_15112,N_15756);
or U16203 (N_16203,N_15336,N_15720);
or U16204 (N_16204,N_14987,N_15072);
xor U16205 (N_16205,N_15838,N_15787);
nand U16206 (N_16206,N_14807,N_14313);
or U16207 (N_16207,N_14307,N_14581);
nand U16208 (N_16208,N_15104,N_14859);
and U16209 (N_16209,N_15729,N_14168);
nor U16210 (N_16210,N_14179,N_14304);
or U16211 (N_16211,N_15938,N_15774);
or U16212 (N_16212,N_15942,N_15385);
or U16213 (N_16213,N_15196,N_14449);
nor U16214 (N_16214,N_15538,N_15120);
and U16215 (N_16215,N_15691,N_14289);
nand U16216 (N_16216,N_14286,N_15155);
nor U16217 (N_16217,N_14248,N_15464);
nor U16218 (N_16218,N_14667,N_14201);
and U16219 (N_16219,N_15118,N_15993);
or U16220 (N_16220,N_14123,N_14639);
and U16221 (N_16221,N_14184,N_14133);
or U16222 (N_16222,N_15950,N_14419);
xor U16223 (N_16223,N_15291,N_14889);
nor U16224 (N_16224,N_15061,N_15088);
nand U16225 (N_16225,N_14114,N_15040);
and U16226 (N_16226,N_15549,N_15970);
nor U16227 (N_16227,N_15152,N_14334);
and U16228 (N_16228,N_15535,N_15311);
nor U16229 (N_16229,N_15798,N_15969);
or U16230 (N_16230,N_14715,N_15898);
and U16231 (N_16231,N_15208,N_15707);
or U16232 (N_16232,N_15030,N_14199);
nor U16233 (N_16233,N_15727,N_15367);
nor U16234 (N_16234,N_14272,N_15992);
and U16235 (N_16235,N_15879,N_14385);
or U16236 (N_16236,N_15626,N_15689);
xor U16237 (N_16237,N_14078,N_15273);
and U16238 (N_16238,N_14588,N_15188);
nor U16239 (N_16239,N_15562,N_14606);
xor U16240 (N_16240,N_14240,N_15238);
and U16241 (N_16241,N_15840,N_15899);
xnor U16242 (N_16242,N_15313,N_14687);
or U16243 (N_16243,N_15568,N_14053);
nor U16244 (N_16244,N_14439,N_14287);
nor U16245 (N_16245,N_14738,N_14453);
xor U16246 (N_16246,N_14091,N_15795);
nand U16247 (N_16247,N_14882,N_14023);
and U16248 (N_16248,N_15553,N_14396);
and U16249 (N_16249,N_15965,N_15465);
nand U16250 (N_16250,N_15534,N_15397);
nand U16251 (N_16251,N_14056,N_14210);
and U16252 (N_16252,N_15953,N_15769);
and U16253 (N_16253,N_15800,N_15985);
nand U16254 (N_16254,N_15034,N_15763);
or U16255 (N_16255,N_14010,N_15757);
xnor U16256 (N_16256,N_15750,N_15492);
xor U16257 (N_16257,N_15663,N_15449);
and U16258 (N_16258,N_15713,N_15144);
xnor U16259 (N_16259,N_14700,N_14696);
or U16260 (N_16260,N_15304,N_14962);
xnor U16261 (N_16261,N_15677,N_14597);
and U16262 (N_16262,N_15440,N_15178);
nand U16263 (N_16263,N_14965,N_14570);
nand U16264 (N_16264,N_15392,N_15651);
and U16265 (N_16265,N_15113,N_14183);
nand U16266 (N_16266,N_14624,N_14704);
xor U16267 (N_16267,N_15973,N_15884);
nand U16268 (N_16268,N_15184,N_15158);
and U16269 (N_16269,N_15332,N_14181);
nor U16270 (N_16270,N_15812,N_15837);
xnor U16271 (N_16271,N_15749,N_15066);
or U16272 (N_16272,N_15620,N_15114);
or U16273 (N_16273,N_15049,N_15323);
or U16274 (N_16274,N_14795,N_15662);
and U16275 (N_16275,N_15434,N_14917);
nor U16276 (N_16276,N_14551,N_15615);
and U16277 (N_16277,N_14233,N_14761);
xor U16278 (N_16278,N_14391,N_14103);
and U16279 (N_16279,N_14209,N_14145);
and U16280 (N_16280,N_14041,N_15041);
and U16281 (N_16281,N_14198,N_14034);
and U16282 (N_16282,N_15575,N_15064);
xnor U16283 (N_16283,N_14207,N_14900);
and U16284 (N_16284,N_15312,N_15907);
nand U16285 (N_16285,N_14101,N_14763);
nand U16286 (N_16286,N_15228,N_15073);
or U16287 (N_16287,N_15820,N_15807);
nand U16288 (N_16288,N_15746,N_14934);
nand U16289 (N_16289,N_15145,N_15052);
or U16290 (N_16290,N_14348,N_14109);
xor U16291 (N_16291,N_14609,N_15732);
xnor U16292 (N_16292,N_14710,N_14390);
or U16293 (N_16293,N_15245,N_14837);
nand U16294 (N_16294,N_14858,N_15638);
nand U16295 (N_16295,N_15715,N_15356);
or U16296 (N_16296,N_14855,N_14276);
nor U16297 (N_16297,N_15730,N_14984);
xnor U16298 (N_16298,N_14617,N_14074);
nor U16299 (N_16299,N_14868,N_15076);
or U16300 (N_16300,N_15223,N_14466);
nor U16301 (N_16301,N_14595,N_15415);
or U16302 (N_16302,N_14351,N_14940);
xor U16303 (N_16303,N_15192,N_15021);
or U16304 (N_16304,N_14523,N_15911);
and U16305 (N_16305,N_14359,N_14107);
nor U16306 (N_16306,N_14770,N_15309);
or U16307 (N_16307,N_15198,N_15292);
nor U16308 (N_16308,N_15177,N_14966);
nand U16309 (N_16309,N_14467,N_15697);
or U16310 (N_16310,N_14623,N_14297);
and U16311 (N_16311,N_14015,N_14245);
and U16312 (N_16312,N_15264,N_14281);
and U16313 (N_16313,N_15379,N_15600);
or U16314 (N_16314,N_14842,N_15444);
nand U16315 (N_16315,N_15125,N_15486);
or U16316 (N_16316,N_15596,N_15067);
or U16317 (N_16317,N_15726,N_14747);
or U16318 (N_16318,N_15149,N_15957);
and U16319 (N_16319,N_14228,N_15811);
and U16320 (N_16320,N_14544,N_15904);
and U16321 (N_16321,N_14404,N_15583);
nor U16322 (N_16322,N_14308,N_15673);
xnor U16323 (N_16323,N_15246,N_14560);
nor U16324 (N_16324,N_14559,N_15410);
nor U16325 (N_16325,N_15913,N_15706);
nand U16326 (N_16326,N_14094,N_14748);
nor U16327 (N_16327,N_15329,N_15194);
xor U16328 (N_16328,N_14455,N_14628);
nor U16329 (N_16329,N_14500,N_15595);
nor U16330 (N_16330,N_14783,N_14402);
nor U16331 (N_16331,N_15445,N_15467);
or U16332 (N_16332,N_14202,N_15325);
nor U16333 (N_16333,N_15024,N_15340);
nor U16334 (N_16334,N_15451,N_14978);
nand U16335 (N_16335,N_15998,N_14808);
nand U16336 (N_16336,N_14471,N_14303);
or U16337 (N_16337,N_15609,N_14656);
and U16338 (N_16338,N_14337,N_15050);
xnor U16339 (N_16339,N_15481,N_14843);
and U16340 (N_16340,N_14853,N_15508);
and U16341 (N_16341,N_15251,N_14860);
nand U16342 (N_16342,N_15491,N_15241);
and U16343 (N_16343,N_14936,N_15971);
nand U16344 (N_16344,N_14043,N_14178);
and U16345 (N_16345,N_15839,N_15896);
nor U16346 (N_16346,N_15207,N_15983);
nand U16347 (N_16347,N_14392,N_15153);
nand U16348 (N_16348,N_15013,N_14767);
and U16349 (N_16349,N_15023,N_14818);
xor U16350 (N_16350,N_14411,N_15817);
or U16351 (N_16351,N_14258,N_14019);
nand U16352 (N_16352,N_14039,N_15216);
nor U16353 (N_16353,N_14587,N_15980);
nor U16354 (N_16354,N_15285,N_14857);
nand U16355 (N_16355,N_15829,N_14212);
nand U16356 (N_16356,N_15058,N_15670);
nand U16357 (N_16357,N_15887,N_15699);
or U16358 (N_16358,N_15436,N_15424);
or U16359 (N_16359,N_15963,N_15653);
nand U16360 (N_16360,N_15462,N_14619);
nand U16361 (N_16361,N_14577,N_14300);
or U16362 (N_16362,N_15268,N_15433);
nor U16363 (N_16363,N_14124,N_14169);
or U16364 (N_16364,N_15698,N_14603);
nand U16365 (N_16365,N_14919,N_15500);
xnor U16366 (N_16366,N_15991,N_15869);
xor U16367 (N_16367,N_15824,N_14293);
and U16368 (N_16368,N_14815,N_14457);
nand U16369 (N_16369,N_14283,N_15000);
and U16370 (N_16370,N_14519,N_14345);
nor U16371 (N_16371,N_14734,N_15632);
nand U16372 (N_16372,N_15927,N_15764);
or U16373 (N_16373,N_14115,N_14264);
nand U16374 (N_16374,N_14938,N_15571);
nand U16375 (N_16375,N_14231,N_15946);
and U16376 (N_16376,N_14273,N_14450);
or U16377 (N_16377,N_15919,N_15843);
and U16378 (N_16378,N_15154,N_14993);
and U16379 (N_16379,N_15502,N_14118);
xor U16380 (N_16380,N_15004,N_15318);
nand U16381 (N_16381,N_15897,N_15190);
nor U16382 (N_16382,N_14405,N_15095);
xor U16383 (N_16383,N_14058,N_15123);
and U16384 (N_16384,N_15522,N_15281);
nor U16385 (N_16385,N_14725,N_15601);
nand U16386 (N_16386,N_15551,N_14257);
and U16387 (N_16387,N_15217,N_14582);
or U16388 (N_16388,N_14873,N_14811);
and U16389 (N_16389,N_14513,N_15335);
nor U16390 (N_16390,N_14924,N_15121);
nor U16391 (N_16391,N_15799,N_15234);
and U16392 (N_16392,N_14244,N_14176);
and U16393 (N_16393,N_14063,N_14372);
or U16394 (N_16394,N_15218,N_14660);
xnor U16395 (N_16395,N_14561,N_15351);
nand U16396 (N_16396,N_15852,N_14788);
nor U16397 (N_16397,N_14931,N_15043);
nand U16398 (N_16398,N_14379,N_14006);
and U16399 (N_16399,N_14378,N_14397);
or U16400 (N_16400,N_15437,N_15124);
or U16401 (N_16401,N_15572,N_15565);
nor U16402 (N_16402,N_14481,N_14353);
nand U16403 (N_16403,N_15947,N_14580);
nand U16404 (N_16404,N_15032,N_14989);
nand U16405 (N_16405,N_14291,N_14451);
and U16406 (N_16406,N_14483,N_15107);
nand U16407 (N_16407,N_14607,N_14355);
xor U16408 (N_16408,N_15920,N_14979);
and U16409 (N_16409,N_14164,N_15738);
nand U16410 (N_16410,N_14225,N_14709);
nor U16411 (N_16411,N_15487,N_14574);
or U16412 (N_16412,N_14562,N_14008);
nand U16413 (N_16413,N_14260,N_14641);
or U16414 (N_16414,N_15468,N_14724);
nand U16415 (N_16415,N_14384,N_15282);
nor U16416 (N_16416,N_14222,N_15858);
or U16417 (N_16417,N_14682,N_14415);
and U16418 (N_16418,N_14753,N_14909);
xor U16419 (N_16419,N_15876,N_15910);
and U16420 (N_16420,N_14221,N_14957);
or U16421 (N_16421,N_15166,N_14638);
and U16422 (N_16422,N_14925,N_14740);
nand U16423 (N_16423,N_15027,N_15881);
nand U16424 (N_16424,N_15393,N_14867);
or U16425 (N_16425,N_14068,N_15162);
nand U16426 (N_16426,N_14726,N_14669);
nor U16427 (N_16427,N_14186,N_15413);
nor U16428 (N_16428,N_14605,N_15081);
xor U16429 (N_16429,N_14400,N_14081);
or U16430 (N_16430,N_15116,N_14819);
nor U16431 (N_16431,N_14002,N_14485);
xor U16432 (N_16432,N_14629,N_15794);
nand U16433 (N_16433,N_15867,N_15425);
nor U16434 (N_16434,N_15053,N_15517);
or U16435 (N_16435,N_15529,N_15917);
nor U16436 (N_16436,N_14218,N_14174);
and U16437 (N_16437,N_14739,N_15803);
and U16438 (N_16438,N_14771,N_14803);
nor U16439 (N_16439,N_14171,N_14830);
and U16440 (N_16440,N_14085,N_14776);
nor U16441 (N_16441,N_14227,N_15660);
nor U16442 (N_16442,N_15895,N_15933);
nor U16443 (N_16443,N_14342,N_15954);
or U16444 (N_16444,N_14226,N_15455);
and U16445 (N_16445,N_14389,N_15625);
nor U16446 (N_16446,N_14678,N_14991);
nand U16447 (N_16447,N_14197,N_14048);
and U16448 (N_16448,N_14901,N_14864);
xor U16449 (N_16449,N_15841,N_15298);
or U16450 (N_16450,N_14986,N_15301);
nand U16451 (N_16451,N_14099,N_15219);
nand U16452 (N_16452,N_15805,N_14333);
nor U16453 (N_16453,N_14489,N_15213);
or U16454 (N_16454,N_14472,N_15466);
nand U16455 (N_16455,N_14336,N_15350);
and U16456 (N_16456,N_15224,N_14665);
nor U16457 (N_16457,N_14516,N_14195);
or U16458 (N_16458,N_14238,N_14584);
nor U16459 (N_16459,N_14025,N_15519);
xnor U16460 (N_16460,N_14737,N_15015);
nand U16461 (N_16461,N_14499,N_14159);
and U16462 (N_16462,N_14821,N_15349);
and U16463 (N_16463,N_14120,N_14393);
or U16464 (N_16464,N_15091,N_15303);
nor U16465 (N_16465,N_14395,N_14526);
nand U16466 (N_16466,N_15501,N_14622);
and U16467 (N_16467,N_14670,N_14825);
and U16468 (N_16468,N_14727,N_14129);
nor U16469 (N_16469,N_15010,N_15227);
xnor U16470 (N_16470,N_15344,N_14503);
or U16471 (N_16471,N_15383,N_15560);
nand U16472 (N_16472,N_14779,N_14812);
and U16473 (N_16473,N_14875,N_15362);
or U16474 (N_16474,N_14401,N_14946);
xor U16475 (N_16475,N_15248,N_15275);
or U16476 (N_16476,N_14650,N_15604);
nand U16477 (N_16477,N_15610,N_15480);
and U16478 (N_16478,N_15031,N_15009);
or U16479 (N_16479,N_14612,N_14437);
nand U16480 (N_16480,N_14167,N_14964);
nand U16481 (N_16481,N_15943,N_15863);
and U16482 (N_16482,N_14527,N_15891);
nor U16483 (N_16483,N_15968,N_14944);
xor U16484 (N_16484,N_14229,N_14851);
nand U16485 (N_16485,N_15935,N_14826);
or U16486 (N_16486,N_14764,N_14157);
nand U16487 (N_16487,N_15592,N_15520);
and U16488 (N_16488,N_15831,N_14532);
nor U16489 (N_16489,N_14386,N_15836);
nor U16490 (N_16490,N_15384,N_15771);
or U16491 (N_16491,N_15056,N_15658);
nand U16492 (N_16492,N_14730,N_14403);
xor U16493 (N_16493,N_14435,N_15722);
or U16494 (N_16494,N_14239,N_15597);
nand U16495 (N_16495,N_15286,N_15314);
nor U16496 (N_16496,N_15616,N_15833);
nor U16497 (N_16497,N_14980,N_15459);
nand U16498 (N_16498,N_14113,N_15330);
nand U16499 (N_16499,N_14951,N_15011);
and U16500 (N_16500,N_15821,N_14996);
and U16501 (N_16501,N_15849,N_15014);
or U16502 (N_16502,N_15686,N_14549);
and U16503 (N_16503,N_15952,N_14820);
or U16504 (N_16504,N_14480,N_14636);
nand U16505 (N_16505,N_14805,N_14718);
and U16506 (N_16506,N_14329,N_15185);
nor U16507 (N_16507,N_15215,N_15674);
and U16508 (N_16508,N_14913,N_15569);
nand U16509 (N_16509,N_15226,N_14200);
nand U16510 (N_16510,N_14926,N_14930);
and U16511 (N_16511,N_15931,N_14626);
nor U16512 (N_16512,N_15117,N_14139);
nand U16513 (N_16513,N_15579,N_14416);
nand U16514 (N_16514,N_14804,N_15602);
nor U16515 (N_16515,N_14490,N_15306);
or U16516 (N_16516,N_15212,N_14119);
nand U16517 (N_16517,N_15339,N_14343);
or U16518 (N_16518,N_14935,N_15022);
nand U16519 (N_16519,N_15779,N_15666);
xnor U16520 (N_16520,N_14555,N_15627);
nor U16521 (N_16521,N_15889,N_15272);
and U16522 (N_16522,N_15263,N_15354);
or U16523 (N_16523,N_15622,N_14536);
and U16524 (N_16524,N_15552,N_15767);
or U16525 (N_16525,N_14375,N_15257);
nor U16526 (N_16526,N_14521,N_14948);
nand U16527 (N_16527,N_14241,N_15842);
nand U16528 (N_16528,N_14033,N_14001);
nor U16529 (N_16529,N_15810,N_14789);
nand U16530 (N_16530,N_14080,N_15164);
nor U16531 (N_16531,N_14237,N_15680);
nor U16532 (N_16532,N_14062,N_15456);
or U16533 (N_16533,N_15521,N_14968);
and U16534 (N_16534,N_14914,N_15369);
and U16535 (N_16535,N_15139,N_14904);
nand U16536 (N_16536,N_14760,N_14310);
or U16537 (N_16537,N_14434,N_14204);
or U16538 (N_16538,N_14688,N_14662);
nand U16539 (N_16539,N_15961,N_15637);
xnor U16540 (N_16540,N_14658,N_14602);
nor U16541 (N_16541,N_15374,N_14035);
and U16542 (N_16542,N_15105,N_14185);
or U16543 (N_16543,N_14162,N_14335);
or U16544 (N_16544,N_15923,N_15001);
nand U16545 (N_16545,N_15737,N_15389);
xor U16546 (N_16546,N_14071,N_14050);
or U16547 (N_16547,N_15411,N_14651);
nand U16548 (N_16548,N_15017,N_15924);
nand U16549 (N_16549,N_15822,N_14030);
nor U16550 (N_16550,N_15555,N_15547);
nor U16551 (N_16551,N_15859,N_15274);
nor U16552 (N_16552,N_14433,N_15815);
nor U16553 (N_16553,N_15315,N_14633);
xor U16554 (N_16554,N_14599,N_14616);
xor U16555 (N_16555,N_15850,N_14741);
and U16556 (N_16556,N_14601,N_14161);
nor U16557 (N_16557,N_14863,N_15703);
or U16558 (N_16558,N_15960,N_15558);
nor U16559 (N_16559,N_14150,N_14759);
nand U16560 (N_16560,N_15846,N_14517);
or U16561 (N_16561,N_15989,N_14649);
nor U16562 (N_16562,N_14927,N_14296);
or U16563 (N_16563,N_15523,N_15603);
or U16564 (N_16564,N_14430,N_14254);
xnor U16565 (N_16565,N_14672,N_15069);
xnor U16566 (N_16566,N_15258,N_15696);
nor U16567 (N_16567,N_14801,N_15682);
xnor U16568 (N_16568,N_15414,N_15888);
and U16569 (N_16569,N_15148,N_15545);
and U16570 (N_16570,N_15959,N_14933);
and U16571 (N_16571,N_15926,N_14077);
nor U16572 (N_16572,N_14051,N_14791);
and U16573 (N_16573,N_14976,N_15310);
xnor U16574 (N_16574,N_14299,N_14427);
and U16575 (N_16575,N_15098,N_15134);
nor U16576 (N_16576,N_14331,N_14029);
nor U16577 (N_16577,N_15326,N_15176);
nand U16578 (N_16578,N_14768,N_15477);
nand U16579 (N_16579,N_14729,N_15087);
and U16580 (N_16580,N_15788,N_14098);
and U16581 (N_16581,N_15265,N_14236);
nor U16582 (N_16582,N_14018,N_15752);
nand U16583 (N_16583,N_14075,N_14275);
nor U16584 (N_16584,N_15127,N_15880);
or U16585 (N_16585,N_14065,N_14394);
and U16586 (N_16586,N_15446,N_14943);
nor U16587 (N_16587,N_14596,N_14699);
nor U16588 (N_16588,N_15316,N_14497);
nor U16589 (N_16589,N_15613,N_15457);
and U16590 (N_16590,N_14326,N_15640);
nand U16591 (N_16591,N_14810,N_15488);
nand U16592 (N_16592,N_14268,N_14220);
and U16593 (N_16593,N_15193,N_15834);
xor U16594 (N_16594,N_15518,N_14681);
and U16595 (N_16595,N_15439,N_14954);
and U16596 (N_16596,N_15008,N_15875);
nor U16597 (N_16597,N_14646,N_14892);
xnor U16598 (N_16598,N_15539,N_15678);
or U16599 (N_16599,N_15284,N_15276);
and U16600 (N_16600,N_14648,N_15644);
xnor U16601 (N_16601,N_15775,N_14838);
nand U16602 (N_16602,N_14126,N_14552);
xnor U16603 (N_16603,N_15505,N_14426);
nand U16604 (N_16604,N_14592,N_14414);
or U16605 (N_16605,N_14692,N_15503);
and U16606 (N_16606,N_15594,N_15921);
xor U16607 (N_16607,N_14016,N_15398);
and U16608 (N_16608,N_15743,N_14781);
nand U16609 (N_16609,N_14079,N_15357);
xor U16610 (N_16610,N_14620,N_15566);
and U16611 (N_16611,N_14492,N_15143);
xor U16612 (N_16612,N_15085,N_14961);
nor U16613 (N_16613,N_15914,N_14849);
and U16614 (N_16614,N_15586,N_14456);
or U16615 (N_16615,N_14608,N_15020);
and U16616 (N_16616,N_14880,N_14478);
nand U16617 (N_16617,N_15033,N_15163);
nor U16618 (N_16618,N_15709,N_15723);
or U16619 (N_16619,N_14149,N_15585);
nor U16620 (N_16620,N_14491,N_15528);
and U16621 (N_16621,N_14720,N_15237);
nor U16622 (N_16622,N_14877,N_15099);
or U16623 (N_16623,N_15253,N_14271);
and U16624 (N_16624,N_14823,N_15997);
or U16625 (N_16625,N_15588,N_15654);
xor U16626 (N_16626,N_15765,N_14382);
or U16627 (N_16627,N_14363,N_14755);
nand U16628 (N_16628,N_14643,N_15082);
nand U16629 (N_16629,N_15808,N_14325);
nand U16630 (N_16630,N_15132,N_14932);
nor U16631 (N_16631,N_14076,N_15062);
and U16632 (N_16632,N_15619,N_14977);
and U16633 (N_16633,N_14874,N_15871);
and U16634 (N_16634,N_14436,N_15509);
nand U16635 (N_16635,N_15005,N_15679);
nor U16636 (N_16636,N_14069,N_15542);
nand U16637 (N_16637,N_14973,N_15271);
nand U16638 (N_16638,N_14816,N_14256);
and U16639 (N_16639,N_14663,N_15930);
or U16640 (N_16640,N_15861,N_15476);
and U16641 (N_16641,N_14165,N_15617);
nor U16642 (N_16642,N_15772,N_15634);
and U16643 (N_16643,N_15819,N_14130);
or U16644 (N_16644,N_14625,N_15165);
nor U16645 (N_16645,N_14380,N_15513);
nor U16646 (N_16646,N_15441,N_14073);
and U16647 (N_16647,N_15130,N_14446);
and U16648 (N_16648,N_14132,N_14590);
xor U16649 (N_16649,N_14387,N_15472);
and U16650 (N_16650,N_14591,N_14947);
and U16651 (N_16651,N_15059,N_14045);
or U16652 (N_16652,N_14148,N_15786);
nor U16653 (N_16653,N_15816,N_14196);
nor U16654 (N_16654,N_14615,N_14495);
or U16655 (N_16655,N_14136,N_14422);
or U16656 (N_16656,N_14469,N_14501);
nand U16657 (N_16657,N_14558,N_15093);
nand U16658 (N_16658,N_14945,N_14265);
xnor U16659 (N_16659,N_15665,N_14235);
nand U16660 (N_16660,N_14027,N_14674);
nor U16661 (N_16661,N_14972,N_14024);
and U16662 (N_16662,N_15386,N_15079);
or U16663 (N_16663,N_15832,N_14910);
nand U16664 (N_16664,N_15421,N_15119);
nor U16665 (N_16665,N_14923,N_14736);
xor U16666 (N_16666,N_15353,N_15789);
nand U16667 (N_16667,N_15941,N_14473);
nor U16668 (N_16668,N_15390,N_15418);
or U16669 (N_16669,N_14543,N_14848);
nand U16670 (N_16670,N_15019,N_14417);
and U16671 (N_16671,N_15790,N_15111);
nand U16672 (N_16672,N_15976,N_15430);
xor U16673 (N_16673,N_15037,N_15802);
or U16674 (N_16674,N_15827,N_15347);
or U16675 (N_16675,N_14955,N_14309);
or U16676 (N_16676,N_14998,N_15029);
nand U16677 (N_16677,N_14916,N_15823);
nor U16678 (N_16678,N_15346,N_15719);
nand U16679 (N_16679,N_14072,N_14066);
and U16680 (N_16680,N_14421,N_14418);
and U16681 (N_16681,N_14886,N_15797);
and U16682 (N_16682,N_14154,N_14476);
nand U16683 (N_16683,N_15405,N_14637);
and U16684 (N_16684,N_14140,N_14959);
nand U16685 (N_16685,N_15563,N_14865);
or U16686 (N_16686,N_14049,N_15847);
nor U16687 (N_16687,N_14999,N_15209);
xnor U16688 (N_16688,N_15758,N_14305);
or U16689 (N_16689,N_14745,N_14589);
nand U16690 (N_16690,N_14288,N_15655);
and U16691 (N_16691,N_14339,N_15716);
nand U16692 (N_16692,N_14537,N_14211);
or U16693 (N_16693,N_15187,N_15782);
nand U16694 (N_16694,N_14470,N_14224);
nor U16695 (N_16695,N_15826,N_15242);
and U16696 (N_16696,N_14474,N_15866);
and U16697 (N_16697,N_15642,N_14367);
nand U16698 (N_16698,N_14794,N_15671);
nor U16699 (N_16699,N_14654,N_14861);
nand U16700 (N_16700,N_14773,N_15352);
and U16701 (N_16701,N_14659,N_14315);
nor U16702 (N_16702,N_14383,N_15028);
and U16703 (N_16703,N_15748,N_14833);
nor U16704 (N_16704,N_15159,N_15690);
nand U16705 (N_16705,N_15183,N_14749);
nor U16706 (N_16706,N_14684,N_15341);
nand U16707 (N_16707,N_14143,N_15129);
xnor U16708 (N_16708,N_14125,N_15412);
or U16709 (N_16709,N_15649,N_14429);
or U16710 (N_16710,N_15636,N_15122);
and U16711 (N_16711,N_14290,N_14614);
or U16712 (N_16712,N_15567,N_15250);
nor U16713 (N_16713,N_14610,N_14302);
nand U16714 (N_16714,N_14769,N_15657);
xor U16715 (N_16715,N_15818,N_15801);
nand U16716 (N_16716,N_15550,N_15222);
nor U16717 (N_16717,N_15966,N_14881);
xor U16718 (N_16718,N_14593,N_15676);
or U16719 (N_16719,N_15373,N_15429);
nor U16720 (N_16720,N_14541,N_14655);
or U16721 (N_16721,N_14243,N_15489);
and U16722 (N_16722,N_15038,N_14046);
and U16723 (N_16723,N_15556,N_14042);
nor U16724 (N_16724,N_15605,N_15200);
xor U16725 (N_16725,N_15431,N_14463);
or U16726 (N_16726,N_15664,N_14420);
or U16727 (N_16727,N_15776,N_15288);
nor U16728 (N_16728,N_14758,N_15599);
or U16729 (N_16729,N_14539,N_14377);
nand U16730 (N_16730,N_15978,N_14792);
or U16731 (N_16731,N_15986,N_15102);
and U16732 (N_16732,N_14887,N_14679);
nor U16733 (N_16733,N_14631,N_14799);
and U16734 (N_16734,N_15708,N_14554);
xor U16735 (N_16735,N_14493,N_15239);
or U16736 (N_16736,N_15402,N_15230);
or U16737 (N_16737,N_14870,N_15478);
nor U16738 (N_16738,N_14061,N_14357);
or U16739 (N_16739,N_15229,N_15825);
and U16740 (N_16740,N_15494,N_15944);
nand U16741 (N_16741,N_14929,N_15893);
and U16742 (N_16742,N_14203,N_15860);
nor U16743 (N_16743,N_14036,N_14319);
nand U16744 (N_16744,N_14412,N_15094);
nand U16745 (N_16745,N_14511,N_15259);
nor U16746 (N_16746,N_15220,N_15109);
nor U16747 (N_16747,N_15358,N_14903);
and U16748 (N_16748,N_15128,N_14369);
or U16749 (N_16749,N_14578,N_15608);
nor U16750 (N_16750,N_15688,N_14565);
nand U16751 (N_16751,N_15851,N_14012);
or U16752 (N_16752,N_14366,N_14458);
and U16753 (N_16753,N_14828,N_14172);
or U16754 (N_16754,N_15201,N_14534);
nor U16755 (N_16755,N_14553,N_15777);
and U16756 (N_16756,N_14388,N_14482);
nor U16757 (N_16757,N_14274,N_15598);
or U16758 (N_16758,N_15406,N_14721);
nor U16759 (N_16759,N_15071,N_15495);
nor U16760 (N_16760,N_14689,N_14032);
nand U16761 (N_16761,N_15182,N_14324);
xor U16762 (N_16762,N_14695,N_14112);
and U16763 (N_16763,N_14356,N_14026);
and U16764 (N_16764,N_15770,N_14127);
and U16765 (N_16765,N_14038,N_14082);
and U16766 (N_16766,N_15179,N_15337);
or U16767 (N_16767,N_14600,N_15407);
nor U16768 (N_16768,N_15845,N_15173);
xnor U16769 (N_16769,N_15883,N_15650);
nor U16770 (N_16770,N_14872,N_14530);
nor U16771 (N_16771,N_14088,N_15042);
and U16772 (N_16772,N_14301,N_15533);
and U16773 (N_16773,N_14697,N_15137);
or U16774 (N_16774,N_15754,N_14508);
or U16775 (N_16775,N_14765,N_14832);
nand U16776 (N_16776,N_14796,N_14548);
and U16777 (N_16777,N_14311,N_14529);
and U16778 (N_16778,N_15206,N_14831);
or U16779 (N_16779,N_15844,N_14707);
or U16780 (N_16780,N_15581,N_15404);
or U16781 (N_16781,N_15780,N_14128);
nor U16782 (N_16782,N_15955,N_14232);
or U16783 (N_16783,N_15656,N_15321);
or U16784 (N_16784,N_14899,N_14263);
nand U16785 (N_16785,N_14742,N_14566);
or U16786 (N_16786,N_14216,N_15573);
nor U16787 (N_16787,N_15661,N_15541);
nor U16788 (N_16788,N_14827,N_15100);
or U16789 (N_16789,N_14000,N_15151);
nor U16790 (N_16790,N_15536,N_14282);
and U16791 (N_16791,N_14160,N_14460);
nor U16792 (N_16792,N_15290,N_14328);
and U16793 (N_16793,N_15894,N_14102);
nand U16794 (N_16794,N_14007,N_15012);
and U16795 (N_16795,N_14895,N_14664);
and U16796 (N_16796,N_14428,N_15507);
or U16797 (N_16797,N_15036,N_14586);
or U16798 (N_16798,N_15994,N_15205);
and U16799 (N_16799,N_14059,N_15077);
or U16800 (N_16800,N_14949,N_15885);
and U16801 (N_16801,N_15511,N_14253);
or U16802 (N_16802,N_14141,N_15962);
xor U16803 (N_16803,N_15928,N_15287);
and U16804 (N_16804,N_14557,N_15561);
nor U16805 (N_16805,N_14569,N_14267);
or U16806 (N_16806,N_15814,N_15101);
nand U16807 (N_16807,N_15003,N_15092);
nand U16808 (N_16808,N_15243,N_15387);
nand U16809 (N_16809,N_15639,N_15607);
nor U16810 (N_16810,N_15484,N_15967);
nor U16811 (N_16811,N_14498,N_15870);
nor U16812 (N_16812,N_14106,N_15171);
xor U16813 (N_16813,N_15140,N_15740);
or U16814 (N_16814,N_14017,N_15160);
nand U16815 (N_16815,N_15510,N_15423);
xnor U16816 (N_16816,N_14583,N_14070);
or U16817 (N_16817,N_14982,N_15537);
or U16818 (N_16818,N_15141,N_15035);
nor U16819 (N_16819,N_14912,N_15687);
nor U16820 (N_16820,N_15548,N_15070);
and U16821 (N_16821,N_14716,N_15648);
nand U16822 (N_16822,N_14528,N_15762);
and U16823 (N_16823,N_14970,N_15375);
nand U16824 (N_16824,N_14317,N_15002);
nand U16825 (N_16825,N_14854,N_14563);
xor U16826 (N_16826,N_15279,N_15400);
or U16827 (N_16827,N_14677,N_14575);
nand U16828 (N_16828,N_14138,N_14621);
nand U16829 (N_16829,N_14413,N_15324);
xor U16830 (N_16830,N_15150,N_14223);
and U16831 (N_16831,N_15210,N_15564);
and U16832 (N_16832,N_15908,N_15161);
nor U16833 (N_16833,N_14247,N_14890);
nor U16834 (N_16834,N_15420,N_14242);
or U16835 (N_16835,N_15334,N_15755);
and U16836 (N_16836,N_15681,N_15949);
or U16837 (N_16837,N_15170,N_14251);
or U16838 (N_16838,N_14694,N_14911);
and U16839 (N_16839,N_15355,N_14352);
or U16840 (N_16840,N_14370,N_15417);
nand U16841 (N_16841,N_15493,N_15932);
nor U16842 (N_16842,N_14744,N_14780);
and U16843 (N_16843,N_15254,N_14693);
nor U16844 (N_16844,N_15221,N_15453);
nand U16845 (N_16845,N_14340,N_14344);
and U16846 (N_16846,N_15751,N_14487);
nand U16847 (N_16847,N_15083,N_14052);
nand U16848 (N_16848,N_14488,N_15447);
nand U16849 (N_16849,N_14152,N_15645);
xnor U16850 (N_16850,N_15956,N_14468);
xor U16851 (N_16851,N_15319,N_14121);
and U16852 (N_16852,N_14153,N_14230);
or U16853 (N_16853,N_14756,N_14671);
nor U16854 (N_16854,N_14496,N_14494);
nor U16855 (N_16855,N_15694,N_14191);
nor U16856 (N_16856,N_14907,N_15399);
or U16857 (N_16857,N_14477,N_14044);
nor U16858 (N_16858,N_15939,N_15331);
nor U16859 (N_16859,N_14567,N_15252);
nand U16860 (N_16860,N_15506,N_15925);
nor U16861 (N_16861,N_14683,N_14087);
nor U16862 (N_16862,N_15873,N_14163);
nand U16863 (N_16863,N_14146,N_15240);
and U16864 (N_16864,N_14285,N_14208);
or U16865 (N_16865,N_15759,N_15380);
or U16866 (N_16866,N_14040,N_14180);
nand U16867 (N_16867,N_14060,N_14969);
or U16868 (N_16868,N_14410,N_15902);
or U16869 (N_16869,N_14089,N_14522);
nand U16870 (N_16870,N_15470,N_15396);
nor U16871 (N_16871,N_15090,N_15089);
or U16872 (N_16872,N_14782,N_14376);
xor U16873 (N_16873,N_14504,N_15416);
xor U16874 (N_16874,N_14706,N_14939);
and U16875 (N_16875,N_15403,N_15338);
nand U16876 (N_16876,N_15882,N_14711);
and U16877 (N_16877,N_15490,N_14459);
and U16878 (N_16878,N_15630,N_14407);
nor U16879 (N_16879,N_15458,N_14425);
xnor U16880 (N_16880,N_15915,N_14368);
nand U16881 (N_16881,N_14188,N_14883);
nor U16882 (N_16882,N_14950,N_14653);
xnor U16883 (N_16883,N_15781,N_14323);
nand U16884 (N_16884,N_15322,N_15857);
xnor U16885 (N_16885,N_15675,N_15255);
or U16886 (N_16886,N_15912,N_14762);
nand U16887 (N_16887,N_14187,N_14189);
or U16888 (N_16888,N_15065,N_15618);
nand U16889 (N_16889,N_14813,N_15195);
and U16890 (N_16890,N_14518,N_14685);
and U16891 (N_16891,N_15591,N_14447);
and U16892 (N_16892,N_15328,N_14166);
and U16893 (N_16893,N_14206,N_14777);
nand U16894 (N_16894,N_14906,N_15172);
nand U16895 (N_16895,N_14640,N_14083);
xor U16896 (N_16896,N_15142,N_15590);
and U16897 (N_16897,N_15475,N_14408);
and U16898 (N_16898,N_15452,N_15728);
and U16899 (N_16899,N_14673,N_15401);
and U16900 (N_16900,N_14862,N_14841);
nor U16901 (N_16901,N_14686,N_14314);
or U16902 (N_16902,N_14893,N_15302);
xnor U16903 (N_16903,N_15525,N_14004);
and U16904 (N_16904,N_14009,N_14571);
nand U16905 (N_16905,N_15524,N_14137);
nand U16906 (N_16906,N_15333,N_15377);
and U16907 (N_16907,N_14871,N_14506);
xor U16908 (N_16908,N_14409,N_14787);
nand U16909 (N_16909,N_15075,N_15136);
nand U16910 (N_16910,N_14852,N_14844);
and U16911 (N_16911,N_15225,N_15348);
nor U16912 (N_16912,N_14332,N_15705);
and U16913 (N_16913,N_15828,N_14869);
and U16914 (N_16914,N_14215,N_15202);
nor U16915 (N_16915,N_15269,N_14280);
nor U16916 (N_16916,N_15307,N_15714);
and U16917 (N_16917,N_14786,N_15051);
xnor U16918 (N_16918,N_15996,N_14292);
xor U16919 (N_16919,N_14261,N_14691);
and U16920 (N_16920,N_14994,N_15133);
or U16921 (N_16921,N_15892,N_15576);
nand U16922 (N_16922,N_14055,N_14520);
or U16923 (N_16923,N_15995,N_14533);
nand U16924 (N_16924,N_15293,N_15736);
nand U16925 (N_16925,N_15717,N_15559);
nand U16926 (N_16926,N_15359,N_14790);
xor U16927 (N_16927,N_14824,N_14524);
and U16928 (N_16928,N_14346,N_15044);
or U16929 (N_16929,N_15108,N_15372);
nand U16930 (N_16930,N_15621,N_14798);
nor U16931 (N_16931,N_15704,N_15886);
and U16932 (N_16932,N_15835,N_15958);
nor U16933 (N_16933,N_15388,N_14373);
xor U16934 (N_16934,N_15724,N_15443);
or U16935 (N_16935,N_15981,N_15463);
or U16936 (N_16936,N_15747,N_14971);
nor U16937 (N_16937,N_15582,N_15578);
xor U16938 (N_16938,N_15760,N_14364);
or U16939 (N_16939,N_14349,N_15532);
nor U16940 (N_16940,N_14942,N_15922);
or U16941 (N_16941,N_14627,N_15624);
nor U16942 (N_16942,N_14341,N_14915);
nand U16943 (N_16943,N_15115,N_15974);
or U16944 (N_16944,N_15381,N_14306);
and U16945 (N_16945,N_14047,N_14464);
and U16946 (N_16946,N_15479,N_15905);
nor U16947 (N_16947,N_14100,N_14361);
nor U16948 (N_16948,N_15175,N_15937);
and U16949 (N_16949,N_14096,N_14084);
or U16950 (N_16950,N_14713,N_15103);
nor U16951 (N_16951,N_15872,N_14573);
and U16952 (N_16952,N_14005,N_15683);
or U16953 (N_16953,N_15874,N_14983);
xor U16954 (N_16954,N_14556,N_14894);
nor U16955 (N_16955,N_14095,N_15305);
nand U16956 (N_16956,N_15126,N_14294);
or U16957 (N_16957,N_14093,N_14431);
nor U16958 (N_16958,N_15454,N_15982);
nor U16959 (N_16959,N_15543,N_15174);
xnor U16960 (N_16960,N_14635,N_15469);
xnor U16961 (N_16961,N_14432,N_15364);
nand U16962 (N_16962,N_15988,N_14104);
or U16963 (N_16963,N_14891,N_14680);
nand U16964 (N_16964,N_15987,N_15514);
nor U16965 (N_16965,N_15068,N_14836);
or U16966 (N_16966,N_14703,N_14896);
nand U16967 (N_16967,N_15450,N_14443);
nor U16968 (N_16968,N_14122,N_14898);
nand U16969 (N_16969,N_14722,N_15684);
xnor U16970 (N_16970,N_15554,N_14057);
or U16971 (N_16971,N_15614,N_15731);
nor U16972 (N_16972,N_15408,N_14003);
nor U16973 (N_16973,N_15647,N_14192);
xnor U16974 (N_16974,N_15643,N_15702);
or U16975 (N_16975,N_14905,N_15395);
or U16976 (N_16976,N_15157,N_14151);
nand U16977 (N_16977,N_14316,N_14031);
or U16978 (N_16978,N_15557,N_14486);
and U16979 (N_16979,N_15862,N_15084);
or U16980 (N_16980,N_14170,N_14277);
or U16981 (N_16981,N_15026,N_14675);
nor U16982 (N_16982,N_14613,N_14441);
nand U16983 (N_16983,N_14735,N_14918);
nor U16984 (N_16984,N_14013,N_15063);
or U16985 (N_16985,N_14542,N_14702);
and U16986 (N_16986,N_15262,N_14173);
xnor U16987 (N_16987,N_15964,N_15432);
nor U16988 (N_16988,N_15854,N_15672);
and U16989 (N_16989,N_15419,N_14644);
nor U16990 (N_16990,N_15791,N_15975);
nand U16991 (N_16991,N_14645,N_15766);
and U16992 (N_16992,N_14809,N_15283);
nor U16993 (N_16993,N_14156,N_15972);
or U16994 (N_16994,N_14158,N_15984);
or U16995 (N_16995,N_15360,N_15540);
or U16996 (N_16996,N_14540,N_14728);
nand U16997 (N_16997,N_14131,N_14320);
or U16998 (N_16998,N_14219,N_14213);
and U16999 (N_16999,N_15426,N_15110);
nand U17000 (N_17000,N_14629,N_14226);
or U17001 (N_17001,N_14965,N_14324);
nand U17002 (N_17002,N_14484,N_14424);
nand U17003 (N_17003,N_15562,N_14237);
and U17004 (N_17004,N_14340,N_15826);
nor U17005 (N_17005,N_15396,N_15858);
or U17006 (N_17006,N_15728,N_14030);
xor U17007 (N_17007,N_15859,N_15153);
nor U17008 (N_17008,N_15104,N_14836);
or U17009 (N_17009,N_14018,N_15642);
nand U17010 (N_17010,N_15102,N_14352);
nor U17011 (N_17011,N_15533,N_15297);
nand U17012 (N_17012,N_14990,N_14933);
nor U17013 (N_17013,N_15415,N_15659);
or U17014 (N_17014,N_14545,N_15983);
nand U17015 (N_17015,N_15441,N_14792);
or U17016 (N_17016,N_14247,N_14400);
and U17017 (N_17017,N_14484,N_15316);
and U17018 (N_17018,N_14125,N_14873);
and U17019 (N_17019,N_14106,N_15734);
and U17020 (N_17020,N_15471,N_15448);
nor U17021 (N_17021,N_14407,N_15272);
nor U17022 (N_17022,N_14399,N_14666);
nor U17023 (N_17023,N_15658,N_15717);
nor U17024 (N_17024,N_14770,N_15566);
xor U17025 (N_17025,N_15351,N_15620);
nor U17026 (N_17026,N_15372,N_14579);
nand U17027 (N_17027,N_14477,N_15959);
nor U17028 (N_17028,N_15048,N_15154);
or U17029 (N_17029,N_14179,N_15301);
nor U17030 (N_17030,N_14843,N_14012);
and U17031 (N_17031,N_14017,N_15157);
or U17032 (N_17032,N_14846,N_15385);
nand U17033 (N_17033,N_15139,N_14423);
and U17034 (N_17034,N_15959,N_15400);
nor U17035 (N_17035,N_15906,N_15655);
xor U17036 (N_17036,N_14156,N_15388);
or U17037 (N_17037,N_15735,N_15059);
nand U17038 (N_17038,N_15105,N_15398);
nand U17039 (N_17039,N_14094,N_15360);
and U17040 (N_17040,N_14974,N_15101);
nand U17041 (N_17041,N_14983,N_15903);
nor U17042 (N_17042,N_14241,N_15922);
xor U17043 (N_17043,N_15400,N_14075);
or U17044 (N_17044,N_15224,N_14840);
nor U17045 (N_17045,N_14280,N_15905);
nand U17046 (N_17046,N_14077,N_15371);
or U17047 (N_17047,N_14802,N_15336);
nor U17048 (N_17048,N_15580,N_15772);
or U17049 (N_17049,N_14576,N_15277);
nor U17050 (N_17050,N_14710,N_15857);
and U17051 (N_17051,N_15233,N_15594);
nand U17052 (N_17052,N_15378,N_15322);
nor U17053 (N_17053,N_14440,N_14986);
or U17054 (N_17054,N_15226,N_15640);
and U17055 (N_17055,N_15597,N_15773);
nor U17056 (N_17056,N_15272,N_14133);
nor U17057 (N_17057,N_14014,N_15777);
nand U17058 (N_17058,N_15615,N_15087);
or U17059 (N_17059,N_14553,N_15456);
and U17060 (N_17060,N_15162,N_15295);
or U17061 (N_17061,N_15243,N_14399);
nand U17062 (N_17062,N_14555,N_15337);
xnor U17063 (N_17063,N_15265,N_15893);
or U17064 (N_17064,N_15670,N_14477);
or U17065 (N_17065,N_14291,N_15478);
nand U17066 (N_17066,N_15096,N_15117);
xnor U17067 (N_17067,N_15670,N_15410);
or U17068 (N_17068,N_15302,N_14851);
and U17069 (N_17069,N_14785,N_14249);
nor U17070 (N_17070,N_14641,N_15326);
nor U17071 (N_17071,N_14595,N_15919);
nor U17072 (N_17072,N_14478,N_15692);
and U17073 (N_17073,N_15715,N_15672);
or U17074 (N_17074,N_14864,N_14115);
or U17075 (N_17075,N_15940,N_14227);
or U17076 (N_17076,N_14666,N_15424);
xnor U17077 (N_17077,N_15118,N_14677);
or U17078 (N_17078,N_15039,N_14380);
nand U17079 (N_17079,N_15841,N_15236);
or U17080 (N_17080,N_15256,N_14472);
nand U17081 (N_17081,N_15084,N_14665);
xnor U17082 (N_17082,N_15282,N_14112);
nand U17083 (N_17083,N_15997,N_15611);
and U17084 (N_17084,N_14701,N_14155);
or U17085 (N_17085,N_14420,N_15088);
and U17086 (N_17086,N_14606,N_15554);
nand U17087 (N_17087,N_15434,N_14252);
and U17088 (N_17088,N_14861,N_15839);
or U17089 (N_17089,N_15751,N_15565);
nand U17090 (N_17090,N_15461,N_15952);
nand U17091 (N_17091,N_14332,N_15393);
nor U17092 (N_17092,N_14794,N_14591);
nand U17093 (N_17093,N_14518,N_15307);
nor U17094 (N_17094,N_15331,N_15476);
nor U17095 (N_17095,N_15051,N_15245);
or U17096 (N_17096,N_15281,N_14347);
and U17097 (N_17097,N_14601,N_15423);
or U17098 (N_17098,N_14443,N_14233);
xor U17099 (N_17099,N_15336,N_14180);
nor U17100 (N_17100,N_15217,N_15080);
nand U17101 (N_17101,N_14388,N_15923);
or U17102 (N_17102,N_15406,N_14364);
and U17103 (N_17103,N_15848,N_15280);
and U17104 (N_17104,N_14129,N_14852);
nand U17105 (N_17105,N_15420,N_15869);
xor U17106 (N_17106,N_14738,N_14664);
xor U17107 (N_17107,N_15388,N_15515);
nor U17108 (N_17108,N_15625,N_14660);
nor U17109 (N_17109,N_14480,N_14090);
xnor U17110 (N_17110,N_15360,N_14211);
and U17111 (N_17111,N_15622,N_15642);
nor U17112 (N_17112,N_15825,N_14673);
nor U17113 (N_17113,N_14606,N_14221);
nor U17114 (N_17114,N_15870,N_15984);
nor U17115 (N_17115,N_15478,N_15630);
nand U17116 (N_17116,N_15988,N_14799);
or U17117 (N_17117,N_14386,N_15791);
and U17118 (N_17118,N_14003,N_14449);
nor U17119 (N_17119,N_15451,N_14955);
xor U17120 (N_17120,N_14640,N_15367);
or U17121 (N_17121,N_14026,N_15231);
and U17122 (N_17122,N_15188,N_15487);
and U17123 (N_17123,N_15455,N_14095);
nand U17124 (N_17124,N_14916,N_14874);
or U17125 (N_17125,N_15158,N_14202);
nand U17126 (N_17126,N_14512,N_14528);
and U17127 (N_17127,N_14186,N_14529);
nand U17128 (N_17128,N_15028,N_14017);
nor U17129 (N_17129,N_14119,N_15525);
nor U17130 (N_17130,N_14567,N_15489);
nand U17131 (N_17131,N_14532,N_15358);
nand U17132 (N_17132,N_15190,N_14339);
and U17133 (N_17133,N_15001,N_15420);
and U17134 (N_17134,N_15056,N_14712);
and U17135 (N_17135,N_14520,N_14537);
and U17136 (N_17136,N_15852,N_15261);
nor U17137 (N_17137,N_15033,N_15662);
nor U17138 (N_17138,N_14432,N_15468);
nor U17139 (N_17139,N_15510,N_15154);
nand U17140 (N_17140,N_14198,N_15310);
nor U17141 (N_17141,N_14481,N_14598);
nand U17142 (N_17142,N_15659,N_15711);
and U17143 (N_17143,N_15237,N_14231);
xor U17144 (N_17144,N_15085,N_14962);
and U17145 (N_17145,N_14511,N_14599);
and U17146 (N_17146,N_15182,N_14308);
xnor U17147 (N_17147,N_15098,N_14383);
and U17148 (N_17148,N_15710,N_14969);
nand U17149 (N_17149,N_15415,N_14999);
nand U17150 (N_17150,N_14073,N_15738);
nor U17151 (N_17151,N_14806,N_14153);
nand U17152 (N_17152,N_15893,N_14541);
xnor U17153 (N_17153,N_14973,N_15582);
and U17154 (N_17154,N_14766,N_15907);
nand U17155 (N_17155,N_15081,N_14339);
or U17156 (N_17156,N_15489,N_15068);
nand U17157 (N_17157,N_15347,N_15160);
nor U17158 (N_17158,N_14476,N_15142);
or U17159 (N_17159,N_15497,N_14879);
or U17160 (N_17160,N_14265,N_15797);
or U17161 (N_17161,N_15661,N_15537);
or U17162 (N_17162,N_15919,N_15022);
nand U17163 (N_17163,N_15215,N_15422);
nor U17164 (N_17164,N_14101,N_15493);
xor U17165 (N_17165,N_14910,N_14951);
nand U17166 (N_17166,N_14171,N_15485);
or U17167 (N_17167,N_14189,N_14138);
nor U17168 (N_17168,N_15676,N_14854);
nand U17169 (N_17169,N_14743,N_15512);
xnor U17170 (N_17170,N_14906,N_14515);
xor U17171 (N_17171,N_14636,N_15869);
and U17172 (N_17172,N_15118,N_14439);
or U17173 (N_17173,N_15080,N_14226);
and U17174 (N_17174,N_15555,N_15867);
or U17175 (N_17175,N_15913,N_14015);
or U17176 (N_17176,N_15454,N_14307);
and U17177 (N_17177,N_15367,N_15378);
or U17178 (N_17178,N_15351,N_15906);
nor U17179 (N_17179,N_14668,N_14506);
or U17180 (N_17180,N_14995,N_14041);
nand U17181 (N_17181,N_14852,N_15617);
nand U17182 (N_17182,N_14212,N_15092);
nor U17183 (N_17183,N_14250,N_14966);
or U17184 (N_17184,N_14329,N_14830);
nor U17185 (N_17185,N_14666,N_14749);
and U17186 (N_17186,N_14316,N_14886);
xor U17187 (N_17187,N_15317,N_15392);
nor U17188 (N_17188,N_15272,N_14507);
and U17189 (N_17189,N_14084,N_14995);
nand U17190 (N_17190,N_15603,N_14890);
and U17191 (N_17191,N_14608,N_14221);
nand U17192 (N_17192,N_15789,N_15552);
nor U17193 (N_17193,N_14563,N_15880);
or U17194 (N_17194,N_14968,N_15323);
xor U17195 (N_17195,N_15869,N_15754);
nand U17196 (N_17196,N_15109,N_14902);
nand U17197 (N_17197,N_15324,N_15754);
xor U17198 (N_17198,N_15268,N_15323);
nand U17199 (N_17199,N_15123,N_14881);
or U17200 (N_17200,N_15264,N_15937);
nor U17201 (N_17201,N_15086,N_15199);
nor U17202 (N_17202,N_14056,N_14250);
or U17203 (N_17203,N_15921,N_14639);
or U17204 (N_17204,N_15690,N_15210);
nor U17205 (N_17205,N_14923,N_14173);
nand U17206 (N_17206,N_14776,N_15852);
xnor U17207 (N_17207,N_14929,N_14605);
xor U17208 (N_17208,N_15322,N_14804);
nor U17209 (N_17209,N_15991,N_15190);
xor U17210 (N_17210,N_14726,N_15089);
or U17211 (N_17211,N_14141,N_14821);
or U17212 (N_17212,N_14034,N_14301);
xor U17213 (N_17213,N_15389,N_15465);
xor U17214 (N_17214,N_14986,N_15776);
xnor U17215 (N_17215,N_14650,N_14251);
or U17216 (N_17216,N_14668,N_14257);
xor U17217 (N_17217,N_15901,N_14424);
xnor U17218 (N_17218,N_14183,N_15989);
xor U17219 (N_17219,N_14303,N_14290);
or U17220 (N_17220,N_14275,N_15544);
nor U17221 (N_17221,N_14032,N_14127);
and U17222 (N_17222,N_15939,N_14966);
xor U17223 (N_17223,N_15130,N_15972);
nor U17224 (N_17224,N_14964,N_14684);
nor U17225 (N_17225,N_14725,N_14015);
and U17226 (N_17226,N_15504,N_14270);
or U17227 (N_17227,N_15825,N_15221);
nor U17228 (N_17228,N_14880,N_14242);
or U17229 (N_17229,N_14051,N_15270);
nor U17230 (N_17230,N_14261,N_14314);
nand U17231 (N_17231,N_14361,N_15310);
and U17232 (N_17232,N_14257,N_15996);
or U17233 (N_17233,N_15872,N_14296);
xnor U17234 (N_17234,N_15571,N_15680);
nor U17235 (N_17235,N_15642,N_14231);
and U17236 (N_17236,N_15457,N_14047);
xnor U17237 (N_17237,N_14441,N_15051);
nand U17238 (N_17238,N_14873,N_14672);
nand U17239 (N_17239,N_14025,N_14390);
and U17240 (N_17240,N_14240,N_15256);
nor U17241 (N_17241,N_14452,N_15784);
and U17242 (N_17242,N_14134,N_15144);
xnor U17243 (N_17243,N_14945,N_14809);
nand U17244 (N_17244,N_14620,N_14669);
nand U17245 (N_17245,N_14208,N_15352);
nand U17246 (N_17246,N_15196,N_14545);
and U17247 (N_17247,N_14405,N_15030);
and U17248 (N_17248,N_15449,N_15619);
and U17249 (N_17249,N_15301,N_14542);
nand U17250 (N_17250,N_14605,N_15677);
or U17251 (N_17251,N_15288,N_14598);
and U17252 (N_17252,N_15183,N_15885);
and U17253 (N_17253,N_14947,N_14155);
nand U17254 (N_17254,N_14832,N_15664);
xor U17255 (N_17255,N_15426,N_14894);
and U17256 (N_17256,N_14390,N_15354);
nand U17257 (N_17257,N_14336,N_14939);
nand U17258 (N_17258,N_15233,N_14428);
or U17259 (N_17259,N_14245,N_14698);
or U17260 (N_17260,N_14727,N_15536);
or U17261 (N_17261,N_15545,N_15670);
nand U17262 (N_17262,N_15250,N_15937);
and U17263 (N_17263,N_15978,N_15577);
xor U17264 (N_17264,N_14872,N_14662);
nor U17265 (N_17265,N_14785,N_14596);
xor U17266 (N_17266,N_14518,N_15311);
nor U17267 (N_17267,N_15843,N_15059);
or U17268 (N_17268,N_15519,N_15397);
and U17269 (N_17269,N_14378,N_15563);
nand U17270 (N_17270,N_15652,N_15814);
and U17271 (N_17271,N_14942,N_14420);
nand U17272 (N_17272,N_15730,N_14185);
or U17273 (N_17273,N_14903,N_15823);
nor U17274 (N_17274,N_15711,N_14969);
nor U17275 (N_17275,N_14198,N_14621);
and U17276 (N_17276,N_15306,N_14379);
or U17277 (N_17277,N_14791,N_14467);
or U17278 (N_17278,N_15894,N_15211);
or U17279 (N_17279,N_14156,N_14574);
nand U17280 (N_17280,N_14986,N_14289);
nand U17281 (N_17281,N_15283,N_14301);
or U17282 (N_17282,N_15769,N_14163);
nor U17283 (N_17283,N_14292,N_14022);
xor U17284 (N_17284,N_15400,N_15435);
nand U17285 (N_17285,N_15722,N_15952);
or U17286 (N_17286,N_15967,N_14381);
nor U17287 (N_17287,N_15159,N_14642);
and U17288 (N_17288,N_15559,N_15095);
or U17289 (N_17289,N_14945,N_14376);
or U17290 (N_17290,N_14024,N_15020);
nand U17291 (N_17291,N_15422,N_15693);
nor U17292 (N_17292,N_15690,N_15276);
and U17293 (N_17293,N_15204,N_15102);
and U17294 (N_17294,N_15518,N_14320);
nand U17295 (N_17295,N_14383,N_15492);
and U17296 (N_17296,N_14606,N_14025);
nor U17297 (N_17297,N_15680,N_15324);
nor U17298 (N_17298,N_14056,N_15375);
and U17299 (N_17299,N_15539,N_15833);
or U17300 (N_17300,N_14772,N_14012);
xnor U17301 (N_17301,N_14190,N_15566);
and U17302 (N_17302,N_15019,N_14475);
nor U17303 (N_17303,N_15396,N_14678);
or U17304 (N_17304,N_15141,N_14111);
nor U17305 (N_17305,N_15436,N_14482);
xnor U17306 (N_17306,N_14163,N_14712);
or U17307 (N_17307,N_15422,N_14266);
or U17308 (N_17308,N_15955,N_15616);
nand U17309 (N_17309,N_14235,N_15259);
and U17310 (N_17310,N_14884,N_15143);
nand U17311 (N_17311,N_15003,N_15795);
or U17312 (N_17312,N_15060,N_14187);
or U17313 (N_17313,N_14668,N_15802);
nor U17314 (N_17314,N_15146,N_14586);
nand U17315 (N_17315,N_14898,N_14120);
nor U17316 (N_17316,N_15909,N_14124);
and U17317 (N_17317,N_15858,N_14234);
or U17318 (N_17318,N_14311,N_14426);
and U17319 (N_17319,N_15379,N_14703);
xor U17320 (N_17320,N_15978,N_14970);
and U17321 (N_17321,N_15021,N_14028);
nor U17322 (N_17322,N_14199,N_15900);
xor U17323 (N_17323,N_14221,N_14949);
nand U17324 (N_17324,N_15703,N_14687);
or U17325 (N_17325,N_14640,N_15617);
nand U17326 (N_17326,N_14401,N_15270);
or U17327 (N_17327,N_14739,N_15530);
or U17328 (N_17328,N_14114,N_15661);
nor U17329 (N_17329,N_14482,N_14642);
nor U17330 (N_17330,N_14494,N_15218);
or U17331 (N_17331,N_14686,N_14797);
and U17332 (N_17332,N_14278,N_14977);
xnor U17333 (N_17333,N_14578,N_14261);
xor U17334 (N_17334,N_15772,N_14329);
and U17335 (N_17335,N_14072,N_14332);
nor U17336 (N_17336,N_14573,N_15345);
nor U17337 (N_17337,N_14259,N_15697);
nor U17338 (N_17338,N_15596,N_14812);
nor U17339 (N_17339,N_15780,N_15487);
nand U17340 (N_17340,N_15978,N_14283);
nand U17341 (N_17341,N_14181,N_15285);
nand U17342 (N_17342,N_14480,N_15121);
and U17343 (N_17343,N_14420,N_14336);
xor U17344 (N_17344,N_15724,N_15746);
nand U17345 (N_17345,N_14238,N_14321);
or U17346 (N_17346,N_15794,N_14029);
nor U17347 (N_17347,N_14363,N_15515);
nand U17348 (N_17348,N_15446,N_15767);
nand U17349 (N_17349,N_15372,N_15716);
nand U17350 (N_17350,N_14166,N_15534);
nor U17351 (N_17351,N_14895,N_15197);
nand U17352 (N_17352,N_15115,N_15954);
and U17353 (N_17353,N_15989,N_14531);
and U17354 (N_17354,N_15793,N_15403);
and U17355 (N_17355,N_14565,N_14339);
xor U17356 (N_17356,N_14268,N_15768);
and U17357 (N_17357,N_14046,N_14542);
nor U17358 (N_17358,N_15463,N_15165);
or U17359 (N_17359,N_15112,N_15452);
or U17360 (N_17360,N_14248,N_15222);
or U17361 (N_17361,N_14265,N_15861);
nand U17362 (N_17362,N_14531,N_14947);
and U17363 (N_17363,N_15766,N_15964);
and U17364 (N_17364,N_15691,N_14689);
or U17365 (N_17365,N_15301,N_14749);
and U17366 (N_17366,N_14147,N_14836);
or U17367 (N_17367,N_15519,N_14731);
nor U17368 (N_17368,N_15568,N_15479);
or U17369 (N_17369,N_14455,N_14021);
and U17370 (N_17370,N_14386,N_15080);
or U17371 (N_17371,N_14695,N_14213);
nor U17372 (N_17372,N_15891,N_15365);
nand U17373 (N_17373,N_14135,N_14338);
and U17374 (N_17374,N_15987,N_14497);
or U17375 (N_17375,N_15041,N_15349);
xnor U17376 (N_17376,N_14176,N_14989);
xnor U17377 (N_17377,N_15090,N_14035);
and U17378 (N_17378,N_14518,N_14051);
xnor U17379 (N_17379,N_15645,N_14190);
nor U17380 (N_17380,N_15613,N_15153);
nand U17381 (N_17381,N_14025,N_14824);
and U17382 (N_17382,N_15929,N_14336);
or U17383 (N_17383,N_15357,N_14484);
xnor U17384 (N_17384,N_15559,N_15328);
or U17385 (N_17385,N_15590,N_14814);
nor U17386 (N_17386,N_15113,N_14176);
and U17387 (N_17387,N_15879,N_15405);
or U17388 (N_17388,N_15270,N_15254);
and U17389 (N_17389,N_14737,N_14504);
nand U17390 (N_17390,N_14769,N_14642);
or U17391 (N_17391,N_15121,N_15304);
nand U17392 (N_17392,N_15184,N_14531);
or U17393 (N_17393,N_15339,N_14050);
nand U17394 (N_17394,N_15381,N_14470);
and U17395 (N_17395,N_15737,N_14622);
and U17396 (N_17396,N_14195,N_14587);
xor U17397 (N_17397,N_15621,N_15355);
or U17398 (N_17398,N_15895,N_15006);
nor U17399 (N_17399,N_14478,N_15823);
and U17400 (N_17400,N_14402,N_14762);
nand U17401 (N_17401,N_14077,N_14262);
and U17402 (N_17402,N_14553,N_15538);
or U17403 (N_17403,N_15397,N_15205);
nor U17404 (N_17404,N_14586,N_14239);
and U17405 (N_17405,N_14442,N_15193);
xnor U17406 (N_17406,N_15335,N_14089);
xnor U17407 (N_17407,N_14394,N_14658);
and U17408 (N_17408,N_15540,N_15299);
xor U17409 (N_17409,N_14540,N_15769);
nand U17410 (N_17410,N_14933,N_15025);
and U17411 (N_17411,N_14934,N_14759);
nor U17412 (N_17412,N_14371,N_14199);
nand U17413 (N_17413,N_14945,N_15162);
and U17414 (N_17414,N_14816,N_15233);
nor U17415 (N_17415,N_14371,N_15117);
nor U17416 (N_17416,N_15130,N_14118);
and U17417 (N_17417,N_15779,N_14225);
nand U17418 (N_17418,N_15088,N_15953);
nand U17419 (N_17419,N_14423,N_15440);
nand U17420 (N_17420,N_15900,N_14378);
nor U17421 (N_17421,N_14579,N_15266);
or U17422 (N_17422,N_15682,N_15864);
nor U17423 (N_17423,N_15368,N_15338);
and U17424 (N_17424,N_15591,N_14748);
nor U17425 (N_17425,N_15063,N_15591);
and U17426 (N_17426,N_14238,N_14105);
xnor U17427 (N_17427,N_15426,N_15000);
or U17428 (N_17428,N_14674,N_15627);
xnor U17429 (N_17429,N_15350,N_14422);
and U17430 (N_17430,N_14358,N_14248);
and U17431 (N_17431,N_15035,N_14763);
and U17432 (N_17432,N_15466,N_15857);
nand U17433 (N_17433,N_14874,N_14990);
nand U17434 (N_17434,N_15365,N_14325);
nand U17435 (N_17435,N_14760,N_14548);
nor U17436 (N_17436,N_14031,N_14771);
and U17437 (N_17437,N_15591,N_15012);
and U17438 (N_17438,N_15789,N_15172);
and U17439 (N_17439,N_14206,N_15763);
xnor U17440 (N_17440,N_15544,N_14473);
nor U17441 (N_17441,N_14138,N_15856);
nor U17442 (N_17442,N_14755,N_15336);
nand U17443 (N_17443,N_14631,N_14226);
or U17444 (N_17444,N_14382,N_14341);
or U17445 (N_17445,N_15396,N_14537);
nand U17446 (N_17446,N_15002,N_15279);
nor U17447 (N_17447,N_15346,N_15104);
nor U17448 (N_17448,N_15928,N_14995);
nand U17449 (N_17449,N_15358,N_15066);
nor U17450 (N_17450,N_15054,N_15785);
xor U17451 (N_17451,N_15944,N_14772);
nor U17452 (N_17452,N_14829,N_15002);
nor U17453 (N_17453,N_14558,N_14582);
nor U17454 (N_17454,N_15048,N_15464);
nand U17455 (N_17455,N_14099,N_15466);
xnor U17456 (N_17456,N_15009,N_15520);
xor U17457 (N_17457,N_14999,N_14228);
nor U17458 (N_17458,N_15519,N_15501);
nand U17459 (N_17459,N_14654,N_15113);
nand U17460 (N_17460,N_14024,N_15749);
and U17461 (N_17461,N_14570,N_14035);
or U17462 (N_17462,N_14112,N_14482);
and U17463 (N_17463,N_15104,N_14263);
nand U17464 (N_17464,N_14958,N_14833);
nor U17465 (N_17465,N_14976,N_14219);
nand U17466 (N_17466,N_14236,N_14203);
xnor U17467 (N_17467,N_14018,N_15455);
and U17468 (N_17468,N_15488,N_15911);
nand U17469 (N_17469,N_14057,N_14276);
or U17470 (N_17470,N_15633,N_15110);
nand U17471 (N_17471,N_14209,N_15839);
nand U17472 (N_17472,N_15263,N_14389);
or U17473 (N_17473,N_15416,N_14811);
and U17474 (N_17474,N_14325,N_14802);
nor U17475 (N_17475,N_14938,N_14044);
xnor U17476 (N_17476,N_15955,N_15857);
or U17477 (N_17477,N_14724,N_15819);
and U17478 (N_17478,N_15304,N_15218);
xnor U17479 (N_17479,N_15671,N_14541);
nand U17480 (N_17480,N_15728,N_14896);
nand U17481 (N_17481,N_14602,N_15677);
nor U17482 (N_17482,N_15389,N_14629);
xnor U17483 (N_17483,N_14992,N_15201);
or U17484 (N_17484,N_15768,N_14945);
and U17485 (N_17485,N_14816,N_14863);
nor U17486 (N_17486,N_14111,N_14581);
or U17487 (N_17487,N_14734,N_15747);
and U17488 (N_17488,N_14981,N_14027);
nand U17489 (N_17489,N_15729,N_14246);
nand U17490 (N_17490,N_14514,N_15382);
or U17491 (N_17491,N_14288,N_14510);
or U17492 (N_17492,N_14900,N_15230);
and U17493 (N_17493,N_14890,N_14525);
or U17494 (N_17494,N_14089,N_15246);
nor U17495 (N_17495,N_14675,N_15753);
xnor U17496 (N_17496,N_14966,N_15471);
nor U17497 (N_17497,N_14077,N_15594);
nand U17498 (N_17498,N_15597,N_14490);
xor U17499 (N_17499,N_14727,N_15505);
nor U17500 (N_17500,N_15162,N_15804);
nor U17501 (N_17501,N_15463,N_14571);
and U17502 (N_17502,N_15629,N_15813);
or U17503 (N_17503,N_15070,N_14797);
nor U17504 (N_17504,N_15363,N_15541);
and U17505 (N_17505,N_15349,N_14900);
nand U17506 (N_17506,N_14211,N_15892);
nand U17507 (N_17507,N_14944,N_14914);
or U17508 (N_17508,N_15822,N_15621);
nand U17509 (N_17509,N_14873,N_15829);
or U17510 (N_17510,N_15903,N_15969);
nand U17511 (N_17511,N_14945,N_14627);
and U17512 (N_17512,N_15586,N_15259);
and U17513 (N_17513,N_14684,N_14674);
nor U17514 (N_17514,N_14754,N_15242);
or U17515 (N_17515,N_14019,N_14516);
nand U17516 (N_17516,N_14815,N_14381);
or U17517 (N_17517,N_15302,N_14836);
and U17518 (N_17518,N_14453,N_14078);
or U17519 (N_17519,N_14561,N_14851);
or U17520 (N_17520,N_15428,N_15271);
nor U17521 (N_17521,N_14729,N_15141);
or U17522 (N_17522,N_14591,N_15848);
or U17523 (N_17523,N_14540,N_15714);
nand U17524 (N_17524,N_14275,N_15100);
nor U17525 (N_17525,N_14227,N_14277);
nor U17526 (N_17526,N_14477,N_14536);
nor U17527 (N_17527,N_14846,N_14098);
nor U17528 (N_17528,N_14107,N_15260);
and U17529 (N_17529,N_14791,N_14683);
or U17530 (N_17530,N_14984,N_15731);
nor U17531 (N_17531,N_14167,N_15508);
and U17532 (N_17532,N_14324,N_15304);
nor U17533 (N_17533,N_14749,N_15142);
xor U17534 (N_17534,N_15338,N_14248);
or U17535 (N_17535,N_14637,N_14656);
nand U17536 (N_17536,N_15909,N_15910);
and U17537 (N_17537,N_14664,N_15567);
nor U17538 (N_17538,N_14959,N_15149);
and U17539 (N_17539,N_14028,N_14255);
nand U17540 (N_17540,N_15800,N_14375);
and U17541 (N_17541,N_15496,N_14970);
or U17542 (N_17542,N_15608,N_14398);
xnor U17543 (N_17543,N_15692,N_15821);
and U17544 (N_17544,N_14162,N_15332);
and U17545 (N_17545,N_14512,N_15400);
or U17546 (N_17546,N_15930,N_15233);
nand U17547 (N_17547,N_15002,N_15043);
nor U17548 (N_17548,N_15769,N_15237);
or U17549 (N_17549,N_15692,N_14401);
nor U17550 (N_17550,N_15185,N_15381);
and U17551 (N_17551,N_14561,N_15111);
or U17552 (N_17552,N_15567,N_15982);
nand U17553 (N_17553,N_14495,N_14224);
nor U17554 (N_17554,N_14157,N_15332);
nand U17555 (N_17555,N_15710,N_15629);
or U17556 (N_17556,N_14903,N_15235);
nand U17557 (N_17557,N_14236,N_15057);
xor U17558 (N_17558,N_15890,N_14352);
and U17559 (N_17559,N_15812,N_14961);
nor U17560 (N_17560,N_14684,N_15431);
or U17561 (N_17561,N_14914,N_14950);
or U17562 (N_17562,N_14601,N_14493);
nand U17563 (N_17563,N_15436,N_15094);
or U17564 (N_17564,N_15707,N_15369);
or U17565 (N_17565,N_14388,N_14648);
or U17566 (N_17566,N_14004,N_15905);
nor U17567 (N_17567,N_14582,N_15095);
or U17568 (N_17568,N_14953,N_14598);
and U17569 (N_17569,N_14068,N_14410);
or U17570 (N_17570,N_15937,N_15347);
and U17571 (N_17571,N_14114,N_15205);
or U17572 (N_17572,N_15815,N_15858);
and U17573 (N_17573,N_14877,N_15750);
xnor U17574 (N_17574,N_15631,N_15090);
nand U17575 (N_17575,N_14777,N_15387);
xor U17576 (N_17576,N_14624,N_15706);
xnor U17577 (N_17577,N_14507,N_15740);
or U17578 (N_17578,N_15672,N_14863);
xor U17579 (N_17579,N_15970,N_15825);
nor U17580 (N_17580,N_14675,N_14414);
nand U17581 (N_17581,N_15702,N_14089);
or U17582 (N_17582,N_14375,N_14497);
nor U17583 (N_17583,N_14171,N_15129);
and U17584 (N_17584,N_15006,N_14792);
nand U17585 (N_17585,N_15314,N_14515);
and U17586 (N_17586,N_14907,N_14264);
nor U17587 (N_17587,N_14067,N_15736);
nand U17588 (N_17588,N_15349,N_14631);
nor U17589 (N_17589,N_15276,N_15781);
or U17590 (N_17590,N_15285,N_15166);
nand U17591 (N_17591,N_14432,N_14428);
nor U17592 (N_17592,N_14400,N_14820);
nor U17593 (N_17593,N_14895,N_15556);
nor U17594 (N_17594,N_14936,N_14971);
nor U17595 (N_17595,N_14514,N_15870);
or U17596 (N_17596,N_14832,N_14651);
and U17597 (N_17597,N_14658,N_15110);
and U17598 (N_17598,N_14364,N_15411);
or U17599 (N_17599,N_15220,N_14465);
or U17600 (N_17600,N_14487,N_14593);
nor U17601 (N_17601,N_15100,N_15261);
nand U17602 (N_17602,N_14342,N_15692);
and U17603 (N_17603,N_14273,N_14026);
xnor U17604 (N_17604,N_14420,N_14114);
xnor U17605 (N_17605,N_14005,N_14397);
nand U17606 (N_17606,N_15007,N_15304);
and U17607 (N_17607,N_14681,N_14908);
nor U17608 (N_17608,N_14005,N_15607);
xor U17609 (N_17609,N_15413,N_14849);
nor U17610 (N_17610,N_15700,N_14031);
or U17611 (N_17611,N_14189,N_14057);
nor U17612 (N_17612,N_14651,N_15515);
nor U17613 (N_17613,N_14231,N_15094);
xnor U17614 (N_17614,N_14741,N_14368);
and U17615 (N_17615,N_15281,N_14706);
nand U17616 (N_17616,N_14596,N_15906);
nor U17617 (N_17617,N_15608,N_14067);
nor U17618 (N_17618,N_15478,N_15702);
nand U17619 (N_17619,N_15896,N_15374);
nand U17620 (N_17620,N_14343,N_14219);
nand U17621 (N_17621,N_14594,N_14548);
and U17622 (N_17622,N_15452,N_14334);
and U17623 (N_17623,N_15583,N_15196);
nand U17624 (N_17624,N_14452,N_15181);
and U17625 (N_17625,N_14896,N_15331);
nand U17626 (N_17626,N_15546,N_15420);
xor U17627 (N_17627,N_15945,N_14147);
and U17628 (N_17628,N_14261,N_14232);
or U17629 (N_17629,N_15718,N_15780);
nor U17630 (N_17630,N_14016,N_14102);
or U17631 (N_17631,N_14582,N_15893);
and U17632 (N_17632,N_14541,N_14934);
and U17633 (N_17633,N_15425,N_15915);
nand U17634 (N_17634,N_15518,N_14228);
and U17635 (N_17635,N_14309,N_14609);
nor U17636 (N_17636,N_14632,N_14025);
or U17637 (N_17637,N_15144,N_15017);
and U17638 (N_17638,N_15325,N_15137);
and U17639 (N_17639,N_15688,N_14500);
nor U17640 (N_17640,N_14894,N_14632);
nand U17641 (N_17641,N_14115,N_15910);
and U17642 (N_17642,N_14163,N_14069);
nand U17643 (N_17643,N_14140,N_14235);
or U17644 (N_17644,N_14631,N_14762);
nand U17645 (N_17645,N_14825,N_15467);
or U17646 (N_17646,N_14507,N_14918);
nor U17647 (N_17647,N_15335,N_14763);
and U17648 (N_17648,N_15204,N_15239);
nand U17649 (N_17649,N_15212,N_14283);
xor U17650 (N_17650,N_15670,N_14938);
xor U17651 (N_17651,N_15088,N_14125);
nor U17652 (N_17652,N_15233,N_15940);
or U17653 (N_17653,N_15051,N_15701);
or U17654 (N_17654,N_14535,N_15303);
nor U17655 (N_17655,N_14508,N_14845);
xnor U17656 (N_17656,N_15206,N_15973);
and U17657 (N_17657,N_14433,N_14684);
xor U17658 (N_17658,N_15604,N_14568);
and U17659 (N_17659,N_14633,N_14742);
and U17660 (N_17660,N_15122,N_15762);
nand U17661 (N_17661,N_14012,N_15719);
nor U17662 (N_17662,N_14813,N_14649);
or U17663 (N_17663,N_14391,N_14850);
nand U17664 (N_17664,N_15567,N_15556);
or U17665 (N_17665,N_14912,N_14103);
nand U17666 (N_17666,N_14378,N_15692);
xor U17667 (N_17667,N_14110,N_15241);
nand U17668 (N_17668,N_14166,N_15084);
or U17669 (N_17669,N_14418,N_15204);
nor U17670 (N_17670,N_15305,N_14062);
nand U17671 (N_17671,N_14403,N_14174);
and U17672 (N_17672,N_15294,N_15887);
and U17673 (N_17673,N_14093,N_15943);
or U17674 (N_17674,N_14193,N_15505);
or U17675 (N_17675,N_14565,N_14102);
nor U17676 (N_17676,N_14019,N_15278);
and U17677 (N_17677,N_15816,N_15929);
or U17678 (N_17678,N_14010,N_15127);
nand U17679 (N_17679,N_14185,N_14143);
and U17680 (N_17680,N_14091,N_15329);
or U17681 (N_17681,N_14365,N_15513);
nand U17682 (N_17682,N_15756,N_15093);
or U17683 (N_17683,N_15289,N_15770);
and U17684 (N_17684,N_15104,N_15461);
nor U17685 (N_17685,N_14178,N_15915);
and U17686 (N_17686,N_14343,N_14806);
nor U17687 (N_17687,N_15083,N_15780);
xnor U17688 (N_17688,N_15786,N_14045);
nand U17689 (N_17689,N_14805,N_15514);
or U17690 (N_17690,N_15372,N_15445);
nand U17691 (N_17691,N_15286,N_14901);
or U17692 (N_17692,N_14790,N_14556);
nand U17693 (N_17693,N_14328,N_15749);
and U17694 (N_17694,N_15910,N_15317);
or U17695 (N_17695,N_15200,N_15527);
nand U17696 (N_17696,N_15975,N_15295);
and U17697 (N_17697,N_14069,N_15792);
nand U17698 (N_17698,N_15735,N_14851);
nand U17699 (N_17699,N_14783,N_15619);
and U17700 (N_17700,N_14781,N_15735);
nor U17701 (N_17701,N_14698,N_15057);
or U17702 (N_17702,N_15083,N_15629);
and U17703 (N_17703,N_14228,N_14252);
and U17704 (N_17704,N_15475,N_15397);
and U17705 (N_17705,N_14926,N_15481);
nand U17706 (N_17706,N_14352,N_15636);
nor U17707 (N_17707,N_14266,N_14203);
nand U17708 (N_17708,N_15189,N_15423);
nand U17709 (N_17709,N_14377,N_14684);
nand U17710 (N_17710,N_15172,N_15114);
nor U17711 (N_17711,N_14333,N_15726);
nand U17712 (N_17712,N_14198,N_14097);
nor U17713 (N_17713,N_15882,N_14508);
xnor U17714 (N_17714,N_15025,N_14477);
nor U17715 (N_17715,N_14075,N_14159);
or U17716 (N_17716,N_14967,N_14891);
nand U17717 (N_17717,N_15356,N_14533);
nor U17718 (N_17718,N_15766,N_15260);
nand U17719 (N_17719,N_15014,N_15081);
nor U17720 (N_17720,N_15380,N_14043);
or U17721 (N_17721,N_14832,N_15752);
and U17722 (N_17722,N_14716,N_15233);
or U17723 (N_17723,N_14464,N_15960);
nand U17724 (N_17724,N_14258,N_14213);
xor U17725 (N_17725,N_15034,N_15645);
nor U17726 (N_17726,N_14702,N_15534);
or U17727 (N_17727,N_15367,N_15681);
nor U17728 (N_17728,N_14072,N_14254);
and U17729 (N_17729,N_15227,N_15491);
nor U17730 (N_17730,N_14129,N_15720);
and U17731 (N_17731,N_14813,N_15958);
nand U17732 (N_17732,N_15742,N_15260);
or U17733 (N_17733,N_15241,N_15378);
or U17734 (N_17734,N_15551,N_15026);
nand U17735 (N_17735,N_15275,N_14781);
and U17736 (N_17736,N_14840,N_15526);
or U17737 (N_17737,N_15196,N_15105);
nand U17738 (N_17738,N_15940,N_15784);
and U17739 (N_17739,N_14493,N_14444);
or U17740 (N_17740,N_15044,N_15350);
nand U17741 (N_17741,N_15896,N_14950);
nor U17742 (N_17742,N_14747,N_14586);
and U17743 (N_17743,N_15972,N_14048);
nor U17744 (N_17744,N_15213,N_14072);
nand U17745 (N_17745,N_14173,N_15550);
nor U17746 (N_17746,N_15832,N_15303);
nor U17747 (N_17747,N_14495,N_14571);
or U17748 (N_17748,N_14521,N_14571);
nand U17749 (N_17749,N_14036,N_14689);
nand U17750 (N_17750,N_15270,N_14044);
or U17751 (N_17751,N_15754,N_14566);
xnor U17752 (N_17752,N_15997,N_14026);
nor U17753 (N_17753,N_14063,N_14272);
and U17754 (N_17754,N_14428,N_15158);
or U17755 (N_17755,N_14631,N_15160);
or U17756 (N_17756,N_14699,N_14070);
and U17757 (N_17757,N_14485,N_15807);
nand U17758 (N_17758,N_15310,N_15781);
nand U17759 (N_17759,N_14099,N_15911);
or U17760 (N_17760,N_14907,N_15888);
nand U17761 (N_17761,N_15663,N_15446);
and U17762 (N_17762,N_15364,N_15185);
nor U17763 (N_17763,N_14742,N_14384);
or U17764 (N_17764,N_14843,N_14079);
and U17765 (N_17765,N_14378,N_14459);
nand U17766 (N_17766,N_15814,N_15752);
nand U17767 (N_17767,N_14091,N_14953);
or U17768 (N_17768,N_14455,N_15735);
and U17769 (N_17769,N_14501,N_14641);
nand U17770 (N_17770,N_15523,N_15347);
xnor U17771 (N_17771,N_15813,N_14228);
and U17772 (N_17772,N_14973,N_14931);
xor U17773 (N_17773,N_14500,N_14991);
nor U17774 (N_17774,N_14051,N_14461);
nor U17775 (N_17775,N_15857,N_14839);
nor U17776 (N_17776,N_14333,N_14780);
nor U17777 (N_17777,N_14162,N_14512);
nand U17778 (N_17778,N_14565,N_15258);
or U17779 (N_17779,N_14326,N_15177);
and U17780 (N_17780,N_14431,N_14585);
nor U17781 (N_17781,N_15296,N_14360);
nand U17782 (N_17782,N_15300,N_14961);
xor U17783 (N_17783,N_15089,N_15773);
nor U17784 (N_17784,N_15882,N_14681);
or U17785 (N_17785,N_15238,N_15485);
or U17786 (N_17786,N_15058,N_14294);
and U17787 (N_17787,N_14447,N_14169);
nor U17788 (N_17788,N_14330,N_14158);
or U17789 (N_17789,N_14276,N_14808);
xnor U17790 (N_17790,N_15021,N_15299);
nor U17791 (N_17791,N_15263,N_14940);
nor U17792 (N_17792,N_15294,N_14004);
nand U17793 (N_17793,N_15001,N_14154);
and U17794 (N_17794,N_14945,N_15228);
and U17795 (N_17795,N_15977,N_14486);
nor U17796 (N_17796,N_14071,N_14910);
xnor U17797 (N_17797,N_14101,N_14626);
or U17798 (N_17798,N_14863,N_14326);
and U17799 (N_17799,N_14383,N_14912);
and U17800 (N_17800,N_14873,N_15044);
nand U17801 (N_17801,N_14609,N_15866);
or U17802 (N_17802,N_15478,N_15527);
nand U17803 (N_17803,N_15493,N_15472);
xnor U17804 (N_17804,N_14393,N_14211);
nand U17805 (N_17805,N_14499,N_15099);
and U17806 (N_17806,N_14239,N_14021);
nand U17807 (N_17807,N_14214,N_14327);
xor U17808 (N_17808,N_14439,N_14644);
nand U17809 (N_17809,N_15920,N_15227);
nand U17810 (N_17810,N_14826,N_14073);
and U17811 (N_17811,N_15991,N_14129);
nor U17812 (N_17812,N_14051,N_15091);
and U17813 (N_17813,N_14678,N_15809);
nor U17814 (N_17814,N_14527,N_15349);
or U17815 (N_17815,N_14551,N_14715);
nand U17816 (N_17816,N_15830,N_15784);
and U17817 (N_17817,N_14578,N_15643);
nor U17818 (N_17818,N_15096,N_14864);
nand U17819 (N_17819,N_14331,N_15806);
and U17820 (N_17820,N_14211,N_15897);
xnor U17821 (N_17821,N_14404,N_15884);
nand U17822 (N_17822,N_15837,N_14857);
nand U17823 (N_17823,N_14597,N_15288);
or U17824 (N_17824,N_14414,N_14782);
and U17825 (N_17825,N_15355,N_15180);
or U17826 (N_17826,N_14330,N_15069);
xor U17827 (N_17827,N_15148,N_15851);
nor U17828 (N_17828,N_14809,N_14988);
nor U17829 (N_17829,N_15026,N_14527);
nand U17830 (N_17830,N_14398,N_14085);
nor U17831 (N_17831,N_15740,N_14481);
nand U17832 (N_17832,N_15635,N_15149);
or U17833 (N_17833,N_14888,N_15658);
xnor U17834 (N_17834,N_15007,N_15926);
or U17835 (N_17835,N_15582,N_15293);
nor U17836 (N_17836,N_15503,N_15545);
or U17837 (N_17837,N_14003,N_14351);
and U17838 (N_17838,N_14490,N_14529);
nand U17839 (N_17839,N_15374,N_14289);
nand U17840 (N_17840,N_14964,N_14110);
and U17841 (N_17841,N_15844,N_15747);
nor U17842 (N_17842,N_15807,N_15232);
nand U17843 (N_17843,N_14085,N_15858);
or U17844 (N_17844,N_15363,N_14756);
nand U17845 (N_17845,N_14424,N_15950);
nor U17846 (N_17846,N_14215,N_15857);
and U17847 (N_17847,N_14319,N_15661);
xor U17848 (N_17848,N_15679,N_15783);
or U17849 (N_17849,N_14122,N_15833);
or U17850 (N_17850,N_14885,N_14281);
and U17851 (N_17851,N_15720,N_15373);
or U17852 (N_17852,N_14308,N_15409);
or U17853 (N_17853,N_15080,N_14848);
or U17854 (N_17854,N_15267,N_14546);
and U17855 (N_17855,N_15969,N_14307);
and U17856 (N_17856,N_14221,N_15680);
nand U17857 (N_17857,N_14491,N_14275);
or U17858 (N_17858,N_15818,N_15237);
nand U17859 (N_17859,N_14890,N_14915);
nand U17860 (N_17860,N_14590,N_15608);
nor U17861 (N_17861,N_15617,N_14765);
nor U17862 (N_17862,N_15195,N_14628);
nor U17863 (N_17863,N_15611,N_14326);
and U17864 (N_17864,N_15648,N_15180);
nand U17865 (N_17865,N_14877,N_15422);
nor U17866 (N_17866,N_15335,N_15398);
or U17867 (N_17867,N_15496,N_14893);
nor U17868 (N_17868,N_15048,N_15049);
xnor U17869 (N_17869,N_15617,N_15069);
and U17870 (N_17870,N_15480,N_15385);
nand U17871 (N_17871,N_14562,N_14150);
nor U17872 (N_17872,N_14477,N_14639);
nand U17873 (N_17873,N_14938,N_14226);
and U17874 (N_17874,N_15229,N_15315);
and U17875 (N_17875,N_15928,N_15170);
nor U17876 (N_17876,N_14346,N_15382);
or U17877 (N_17877,N_15853,N_15772);
or U17878 (N_17878,N_15343,N_14440);
nor U17879 (N_17879,N_14468,N_15669);
and U17880 (N_17880,N_14860,N_15520);
nor U17881 (N_17881,N_14953,N_15330);
and U17882 (N_17882,N_15828,N_15789);
nand U17883 (N_17883,N_14887,N_14530);
and U17884 (N_17884,N_15420,N_14309);
nor U17885 (N_17885,N_15088,N_15649);
nand U17886 (N_17886,N_14795,N_14925);
nor U17887 (N_17887,N_14687,N_14839);
and U17888 (N_17888,N_14881,N_15235);
nor U17889 (N_17889,N_15572,N_15083);
or U17890 (N_17890,N_14455,N_15536);
nor U17891 (N_17891,N_15197,N_15069);
or U17892 (N_17892,N_14438,N_14734);
or U17893 (N_17893,N_15950,N_15162);
xor U17894 (N_17894,N_15896,N_14214);
and U17895 (N_17895,N_14221,N_15224);
nor U17896 (N_17896,N_14209,N_14529);
nor U17897 (N_17897,N_15889,N_15036);
nand U17898 (N_17898,N_14408,N_15865);
and U17899 (N_17899,N_15655,N_15657);
or U17900 (N_17900,N_14363,N_15443);
and U17901 (N_17901,N_15973,N_14070);
and U17902 (N_17902,N_15819,N_15625);
and U17903 (N_17903,N_15650,N_14001);
nor U17904 (N_17904,N_14303,N_15267);
xnor U17905 (N_17905,N_15812,N_14610);
or U17906 (N_17906,N_14514,N_14963);
nand U17907 (N_17907,N_14395,N_15725);
nor U17908 (N_17908,N_15187,N_14127);
nand U17909 (N_17909,N_15634,N_15733);
nand U17910 (N_17910,N_14805,N_15572);
and U17911 (N_17911,N_15221,N_14766);
or U17912 (N_17912,N_15962,N_14588);
xor U17913 (N_17913,N_15584,N_14144);
nor U17914 (N_17914,N_14440,N_14848);
xor U17915 (N_17915,N_14768,N_14339);
nand U17916 (N_17916,N_14176,N_15541);
xnor U17917 (N_17917,N_15877,N_15139);
or U17918 (N_17918,N_14395,N_14848);
nor U17919 (N_17919,N_14632,N_14898);
nor U17920 (N_17920,N_15436,N_14674);
and U17921 (N_17921,N_14466,N_14412);
and U17922 (N_17922,N_15968,N_14902);
or U17923 (N_17923,N_14677,N_15974);
and U17924 (N_17924,N_14134,N_15880);
or U17925 (N_17925,N_15586,N_15581);
and U17926 (N_17926,N_14873,N_15095);
xor U17927 (N_17927,N_15960,N_14259);
and U17928 (N_17928,N_15313,N_14540);
or U17929 (N_17929,N_14230,N_14745);
nor U17930 (N_17930,N_15053,N_14578);
nand U17931 (N_17931,N_14533,N_15195);
nor U17932 (N_17932,N_15358,N_15294);
nand U17933 (N_17933,N_14261,N_14041);
and U17934 (N_17934,N_15910,N_14536);
xor U17935 (N_17935,N_15038,N_15071);
nor U17936 (N_17936,N_15731,N_15450);
nor U17937 (N_17937,N_15080,N_15231);
or U17938 (N_17938,N_14344,N_14581);
xnor U17939 (N_17939,N_14532,N_14093);
nand U17940 (N_17940,N_14450,N_14561);
and U17941 (N_17941,N_15143,N_14388);
nand U17942 (N_17942,N_14035,N_15005);
nor U17943 (N_17943,N_15069,N_15692);
xor U17944 (N_17944,N_14612,N_14082);
or U17945 (N_17945,N_15431,N_15571);
and U17946 (N_17946,N_14932,N_14284);
or U17947 (N_17947,N_14066,N_14996);
nor U17948 (N_17948,N_15368,N_15840);
or U17949 (N_17949,N_14492,N_15429);
xor U17950 (N_17950,N_15059,N_14850);
or U17951 (N_17951,N_15588,N_14475);
and U17952 (N_17952,N_14270,N_14676);
or U17953 (N_17953,N_14623,N_15665);
and U17954 (N_17954,N_14604,N_15433);
xnor U17955 (N_17955,N_15175,N_15103);
nor U17956 (N_17956,N_15440,N_14886);
nor U17957 (N_17957,N_14456,N_14569);
and U17958 (N_17958,N_14429,N_15835);
or U17959 (N_17959,N_14358,N_15291);
or U17960 (N_17960,N_15199,N_15321);
nor U17961 (N_17961,N_15073,N_15166);
or U17962 (N_17962,N_14783,N_14009);
nor U17963 (N_17963,N_14095,N_15982);
or U17964 (N_17964,N_14065,N_15217);
nor U17965 (N_17965,N_14446,N_15760);
nand U17966 (N_17966,N_14024,N_15874);
nand U17967 (N_17967,N_14800,N_15781);
or U17968 (N_17968,N_15868,N_14300);
and U17969 (N_17969,N_15715,N_14064);
or U17970 (N_17970,N_15283,N_14940);
nor U17971 (N_17971,N_14109,N_14562);
xnor U17972 (N_17972,N_14560,N_14394);
nor U17973 (N_17973,N_15703,N_14981);
and U17974 (N_17974,N_15689,N_15175);
and U17975 (N_17975,N_14377,N_14300);
and U17976 (N_17976,N_14472,N_15108);
nor U17977 (N_17977,N_15258,N_15105);
nor U17978 (N_17978,N_14420,N_15827);
xnor U17979 (N_17979,N_15754,N_15673);
nand U17980 (N_17980,N_14886,N_15736);
nand U17981 (N_17981,N_14565,N_14431);
nor U17982 (N_17982,N_14838,N_15394);
nand U17983 (N_17983,N_15507,N_15623);
and U17984 (N_17984,N_14467,N_14463);
xnor U17985 (N_17985,N_15446,N_15532);
and U17986 (N_17986,N_15804,N_15625);
nand U17987 (N_17987,N_14440,N_15018);
xor U17988 (N_17988,N_14863,N_15659);
nor U17989 (N_17989,N_15937,N_15982);
nor U17990 (N_17990,N_14013,N_15427);
or U17991 (N_17991,N_15807,N_14245);
or U17992 (N_17992,N_14093,N_15904);
nor U17993 (N_17993,N_14871,N_14876);
or U17994 (N_17994,N_14380,N_15161);
or U17995 (N_17995,N_14814,N_14943);
xor U17996 (N_17996,N_15487,N_15654);
or U17997 (N_17997,N_15214,N_14042);
and U17998 (N_17998,N_15605,N_14557);
xnor U17999 (N_17999,N_15949,N_14957);
nor U18000 (N_18000,N_16089,N_17363);
nand U18001 (N_18001,N_17195,N_17884);
nor U18002 (N_18002,N_16795,N_16568);
nand U18003 (N_18003,N_17590,N_16963);
and U18004 (N_18004,N_16161,N_16815);
and U18005 (N_18005,N_17581,N_16122);
nand U18006 (N_18006,N_16425,N_16358);
or U18007 (N_18007,N_16666,N_16481);
nor U18008 (N_18008,N_17084,N_16810);
or U18009 (N_18009,N_16486,N_16528);
nand U18010 (N_18010,N_17088,N_17587);
nand U18011 (N_18011,N_17068,N_17053);
or U18012 (N_18012,N_17516,N_16171);
nand U18013 (N_18013,N_16411,N_16025);
nand U18014 (N_18014,N_17118,N_17069);
nor U18015 (N_18015,N_17530,N_17675);
or U18016 (N_18016,N_17558,N_17862);
nand U18017 (N_18017,N_17848,N_17751);
nand U18018 (N_18018,N_17125,N_16389);
nor U18019 (N_18019,N_17493,N_17735);
or U18020 (N_18020,N_16067,N_17514);
and U18021 (N_18021,N_17001,N_16013);
and U18022 (N_18022,N_17824,N_17468);
nand U18023 (N_18023,N_16224,N_16840);
or U18024 (N_18024,N_17046,N_17935);
or U18025 (N_18025,N_16729,N_16300);
or U18026 (N_18026,N_17034,N_16146);
nor U18027 (N_18027,N_16539,N_17292);
xnor U18028 (N_18028,N_16355,N_16147);
nand U18029 (N_18029,N_16672,N_17703);
nor U18030 (N_18030,N_17155,N_16827);
nand U18031 (N_18031,N_17537,N_17713);
or U18032 (N_18032,N_16369,N_16833);
or U18033 (N_18033,N_17816,N_16804);
or U18034 (N_18034,N_16599,N_16611);
or U18035 (N_18035,N_17184,N_16744);
or U18036 (N_18036,N_16868,N_16992);
nand U18037 (N_18037,N_17056,N_17305);
nor U18038 (N_18038,N_16386,N_16303);
or U18039 (N_18039,N_16427,N_17905);
xnor U18040 (N_18040,N_16096,N_16091);
or U18041 (N_18041,N_16176,N_17996);
nand U18042 (N_18042,N_17597,N_17762);
nor U18043 (N_18043,N_17176,N_17976);
or U18044 (N_18044,N_17213,N_16726);
and U18045 (N_18045,N_16855,N_16715);
or U18046 (N_18046,N_16601,N_16137);
and U18047 (N_18047,N_16825,N_16768);
nor U18048 (N_18048,N_16033,N_16035);
nand U18049 (N_18049,N_17781,N_17812);
nand U18050 (N_18050,N_16201,N_17523);
and U18051 (N_18051,N_17770,N_17253);
and U18052 (N_18052,N_16724,N_17170);
and U18053 (N_18053,N_17303,N_17027);
nor U18054 (N_18054,N_16969,N_16330);
xor U18055 (N_18055,N_17149,N_17702);
or U18056 (N_18056,N_17786,N_16961);
or U18057 (N_18057,N_16203,N_16124);
nor U18058 (N_18058,N_16291,N_16167);
nor U18059 (N_18059,N_17763,N_17980);
nor U18060 (N_18060,N_17355,N_16678);
and U18061 (N_18061,N_17089,N_16616);
nand U18062 (N_18062,N_17116,N_17028);
nand U18063 (N_18063,N_16749,N_17321);
and U18064 (N_18064,N_16602,N_17851);
xnor U18065 (N_18065,N_16991,N_17758);
or U18066 (N_18066,N_17991,N_16640);
nor U18067 (N_18067,N_17964,N_16354);
and U18068 (N_18068,N_17246,N_17030);
and U18069 (N_18069,N_16445,N_17108);
nor U18070 (N_18070,N_16174,N_17706);
or U18071 (N_18071,N_17014,N_17747);
nor U18072 (N_18072,N_16631,N_16366);
or U18073 (N_18073,N_17994,N_17765);
or U18074 (N_18074,N_17619,N_17110);
nor U18075 (N_18075,N_16928,N_17608);
and U18076 (N_18076,N_17956,N_16456);
and U18077 (N_18077,N_17804,N_16394);
and U18078 (N_18078,N_17111,N_16727);
nor U18079 (N_18079,N_16003,N_17924);
and U18080 (N_18080,N_16641,N_17614);
or U18081 (N_18081,N_16981,N_17696);
nor U18082 (N_18082,N_17230,N_17051);
or U18083 (N_18083,N_17210,N_16031);
or U18084 (N_18084,N_17559,N_16867);
nor U18085 (N_18085,N_16058,N_16865);
and U18086 (N_18086,N_16342,N_16540);
nand U18087 (N_18087,N_16316,N_16114);
nor U18088 (N_18088,N_17607,N_16084);
nand U18089 (N_18089,N_17160,N_17162);
nand U18090 (N_18090,N_17359,N_16069);
nor U18091 (N_18091,N_16955,N_17969);
or U18092 (N_18092,N_16580,N_16413);
or U18093 (N_18093,N_17930,N_16409);
nand U18094 (N_18094,N_16041,N_16883);
xor U18095 (N_18095,N_17265,N_16112);
or U18096 (N_18096,N_17502,N_17031);
xor U18097 (N_18097,N_17333,N_17904);
nor U18098 (N_18098,N_17352,N_17284);
nand U18099 (N_18099,N_17495,N_17868);
and U18100 (N_18100,N_17882,N_17187);
nand U18101 (N_18101,N_17754,N_16449);
or U18102 (N_18102,N_16153,N_16478);
and U18103 (N_18103,N_16095,N_17504);
nand U18104 (N_18104,N_17060,N_17768);
and U18105 (N_18105,N_17551,N_17448);
and U18106 (N_18106,N_17939,N_17256);
xor U18107 (N_18107,N_17165,N_17217);
or U18108 (N_18108,N_17147,N_16260);
nor U18109 (N_18109,N_17711,N_17313);
or U18110 (N_18110,N_17346,N_16982);
and U18111 (N_18111,N_17673,N_16619);
nand U18112 (N_18112,N_16085,N_17995);
xnor U18113 (N_18113,N_17287,N_17311);
or U18114 (N_18114,N_16110,N_16699);
or U18115 (N_18115,N_17278,N_16464);
nor U18116 (N_18116,N_17865,N_16737);
nand U18117 (N_18117,N_17017,N_17986);
nor U18118 (N_18118,N_17442,N_16716);
or U18119 (N_18119,N_16861,N_16107);
nand U18120 (N_18120,N_17387,N_16824);
nand U18121 (N_18121,N_17766,N_17972);
nand U18122 (N_18122,N_16372,N_16617);
xnor U18123 (N_18123,N_17441,N_16663);
nor U18124 (N_18124,N_17745,N_16871);
and U18125 (N_18125,N_17720,N_17693);
or U18126 (N_18126,N_17852,N_16485);
and U18127 (N_18127,N_17338,N_16151);
nor U18128 (N_18128,N_16011,N_17436);
nor U18129 (N_18129,N_17308,N_17827);
or U18130 (N_18130,N_17933,N_17738);
or U18131 (N_18131,N_17512,N_16205);
nand U18132 (N_18132,N_16015,N_16569);
and U18133 (N_18133,N_16392,N_17906);
nand U18134 (N_18134,N_16851,N_17471);
or U18135 (N_18135,N_17499,N_16491);
and U18136 (N_18136,N_16270,N_16063);
or U18137 (N_18137,N_16287,N_17207);
and U18138 (N_18138,N_16071,N_17802);
and U18139 (N_18139,N_17332,N_17074);
and U18140 (N_18140,N_16200,N_16863);
and U18141 (N_18141,N_17261,N_16362);
nand U18142 (N_18142,N_17741,N_17992);
nor U18143 (N_18143,N_16115,N_16162);
and U18144 (N_18144,N_16459,N_16347);
nand U18145 (N_18145,N_16779,N_17534);
nand U18146 (N_18146,N_16022,N_16686);
and U18147 (N_18147,N_17314,N_17909);
or U18148 (N_18148,N_16315,N_16424);
nor U18149 (N_18149,N_17343,N_17266);
nor U18150 (N_18150,N_17339,N_17129);
and U18151 (N_18151,N_17109,N_16391);
nand U18152 (N_18152,N_17055,N_16434);
or U18153 (N_18153,N_16783,N_16059);
and U18154 (N_18154,N_17224,N_16852);
and U18155 (N_18155,N_16074,N_16446);
nand U18156 (N_18156,N_17222,N_16468);
nor U18157 (N_18157,N_17379,N_17592);
and U18158 (N_18158,N_17518,N_17035);
or U18159 (N_18159,N_16739,N_17272);
and U18160 (N_18160,N_16098,N_16971);
or U18161 (N_18161,N_16210,N_16276);
nand U18162 (N_18162,N_17390,N_16769);
nor U18163 (N_18163,N_16809,N_16390);
xor U18164 (N_18164,N_16357,N_17583);
nand U18165 (N_18165,N_16383,N_17076);
or U18166 (N_18166,N_16374,N_16836);
or U18167 (N_18167,N_16562,N_16066);
xnor U18168 (N_18168,N_17669,N_16417);
or U18169 (N_18169,N_17206,N_17179);
nor U18170 (N_18170,N_16054,N_16707);
nand U18171 (N_18171,N_17503,N_16428);
nor U18172 (N_18172,N_16683,N_16521);
and U18173 (N_18173,N_16873,N_16049);
nand U18174 (N_18174,N_16613,N_16719);
nor U18175 (N_18175,N_17895,N_16333);
nand U18176 (N_18176,N_17717,N_16767);
and U18177 (N_18177,N_17524,N_16450);
and U18178 (N_18178,N_16217,N_16322);
or U18179 (N_18179,N_17281,N_17022);
nor U18180 (N_18180,N_16125,N_17778);
or U18181 (N_18181,N_16311,N_17137);
and U18182 (N_18182,N_16692,N_16940);
or U18183 (N_18183,N_17011,N_17984);
and U18184 (N_18184,N_17694,N_16194);
nand U18185 (N_18185,N_17856,N_17624);
nand U18186 (N_18186,N_17844,N_17577);
nor U18187 (N_18187,N_17671,N_16585);
xnor U18188 (N_18188,N_17189,N_16844);
nor U18189 (N_18189,N_17357,N_17626);
nor U18190 (N_18190,N_17200,N_17479);
nand U18191 (N_18191,N_16133,N_17135);
or U18192 (N_18192,N_16774,N_17556);
nand U18193 (N_18193,N_16302,N_17526);
and U18194 (N_18194,N_17948,N_16244);
and U18195 (N_18195,N_17423,N_16312);
xor U18196 (N_18196,N_16475,N_17817);
nor U18197 (N_18197,N_16983,N_16968);
and U18198 (N_18198,N_17231,N_16890);
or U18199 (N_18199,N_16249,N_17609);
xnor U18200 (N_18200,N_16508,N_16495);
or U18201 (N_18201,N_17743,N_16029);
xor U18202 (N_18202,N_16088,N_16627);
or U18203 (N_18203,N_16525,N_17527);
and U18204 (N_18204,N_16423,N_16950);
or U18205 (N_18205,N_17954,N_16297);
nand U18206 (N_18206,N_17212,N_17401);
and U18207 (N_18207,N_16023,N_16913);
nand U18208 (N_18208,N_17150,N_16657);
nand U18209 (N_18209,N_17191,N_16293);
and U18210 (N_18210,N_16835,N_16897);
and U18211 (N_18211,N_16717,N_16236);
nor U18212 (N_18212,N_17121,N_17668);
or U18213 (N_18213,N_16283,N_16043);
nor U18214 (N_18214,N_17368,N_16888);
xor U18215 (N_18215,N_17136,N_17511);
and U18216 (N_18216,N_17012,N_17688);
and U18217 (N_18217,N_16185,N_17329);
nor U18218 (N_18218,N_16172,N_17797);
nand U18219 (N_18219,N_16519,N_16030);
and U18220 (N_18220,N_16473,N_16645);
nand U18221 (N_18221,N_17744,N_17025);
nor U18222 (N_18222,N_17023,N_16170);
nand U18223 (N_18223,N_16944,N_17750);
nor U18224 (N_18224,N_16537,N_16247);
nand U18225 (N_18225,N_16635,N_17925);
and U18226 (N_18226,N_16436,N_16251);
and U18227 (N_18227,N_16614,N_17737);
or U18228 (N_18228,N_17480,N_16404);
or U18229 (N_18229,N_17394,N_17452);
nor U18230 (N_18230,N_17683,N_16552);
nand U18231 (N_18231,N_16917,N_16301);
nand U18232 (N_18232,N_16393,N_17463);
nand U18233 (N_18233,N_16860,N_16024);
and U18234 (N_18234,N_16009,N_16509);
nor U18235 (N_18235,N_17454,N_16880);
and U18236 (N_18236,N_16549,N_17348);
nor U18237 (N_18237,N_17501,N_17845);
or U18238 (N_18238,N_16660,N_17007);
and U18239 (N_18239,N_17400,N_16572);
nor U18240 (N_18240,N_16016,N_17033);
and U18241 (N_18241,N_16820,N_17467);
or U18242 (N_18242,N_17732,N_16040);
or U18243 (N_18243,N_16503,N_17531);
nand U18244 (N_18244,N_16214,N_16144);
and U18245 (N_18245,N_16999,N_16742);
and U18246 (N_18246,N_17126,N_17634);
nor U18247 (N_18247,N_16187,N_16285);
nor U18248 (N_18248,N_17557,N_16255);
xor U18249 (N_18249,N_16697,N_16651);
nand U18250 (N_18250,N_17712,N_17640);
xnor U18251 (N_18251,N_17917,N_16972);
and U18252 (N_18252,N_17815,N_17615);
nand U18253 (N_18253,N_17075,N_17585);
nor U18254 (N_18254,N_17307,N_17044);
nand U18255 (N_18255,N_17918,N_16556);
and U18256 (N_18256,N_17262,N_17795);
xnor U18257 (N_18257,N_16363,N_16269);
and U18258 (N_18258,N_17748,N_16198);
nand U18259 (N_18259,N_17837,N_16988);
and U18260 (N_18260,N_17697,N_16885);
and U18261 (N_18261,N_16329,N_16546);
nand U18262 (N_18262,N_17414,N_17990);
nand U18263 (N_18263,N_16350,N_17013);
nand U18264 (N_18264,N_16228,N_16839);
and U18265 (N_18265,N_17568,N_16348);
and U18266 (N_18266,N_17775,N_17185);
nor U18267 (N_18267,N_16520,N_17029);
nand U18268 (N_18268,N_16507,N_17600);
and U18269 (N_18269,N_16689,N_17296);
or U18270 (N_18270,N_16670,N_16159);
or U18271 (N_18271,N_17532,N_16400);
nand U18272 (N_18272,N_17891,N_16328);
nand U18273 (N_18273,N_17910,N_16952);
nand U18274 (N_18274,N_17753,N_17769);
or U18275 (N_18275,N_17545,N_17081);
or U18276 (N_18276,N_16044,N_16431);
and U18277 (N_18277,N_17999,N_16169);
nor U18278 (N_18278,N_16935,N_16216);
and U18279 (N_18279,N_16684,N_17708);
nor U18280 (N_18280,N_16581,N_17038);
and U18281 (N_18281,N_17490,N_16735);
or U18282 (N_18282,N_17263,N_16643);
or U18283 (N_18283,N_16625,N_17746);
or U18284 (N_18284,N_17090,N_17877);
nand U18285 (N_18285,N_16760,N_17240);
nor U18286 (N_18286,N_17234,N_17628);
nor U18287 (N_18287,N_17589,N_16788);
nand U18288 (N_18288,N_17705,N_17275);
nand U18289 (N_18289,N_17617,N_16649);
or U18290 (N_18290,N_17755,N_17715);
xnor U18291 (N_18291,N_17790,N_16579);
or U18292 (N_18292,N_16131,N_17949);
nand U18293 (N_18293,N_16594,N_16265);
nand U18294 (N_18294,N_17888,N_17131);
xnor U18295 (N_18295,N_16278,N_16837);
nand U18296 (N_18296,N_16946,N_16470);
nand U18297 (N_18297,N_17405,N_17897);
nor U18298 (N_18298,N_17641,N_17546);
nor U18299 (N_18299,N_17959,N_16419);
nor U18300 (N_18300,N_16104,N_17309);
and U18301 (N_18301,N_16762,N_16878);
xor U18302 (N_18302,N_17805,N_17000);
nand U18303 (N_18303,N_17916,N_17470);
nor U18304 (N_18304,N_17039,N_16256);
nor U18305 (N_18305,N_17961,N_17606);
nor U18306 (N_18306,N_16238,N_17901);
or U18307 (N_18307,N_16662,N_17367);
nand U18308 (N_18308,N_17774,N_16081);
xnor U18309 (N_18309,N_17836,N_17465);
nor U18310 (N_18310,N_16910,N_16036);
nor U18311 (N_18311,N_16800,N_17840);
xnor U18312 (N_18312,N_17067,N_16529);
and U18313 (N_18313,N_16032,N_16230);
nor U18314 (N_18314,N_16240,N_17870);
nor U18315 (N_18315,N_17214,N_17937);
or U18316 (N_18316,N_16818,N_16028);
xor U18317 (N_18317,N_17855,N_17473);
or U18318 (N_18318,N_17579,N_16904);
xor U18319 (N_18319,N_16829,N_16489);
nand U18320 (N_18320,N_17105,N_17345);
nor U18321 (N_18321,N_17366,N_16189);
nand U18322 (N_18322,N_17974,N_17298);
xnor U18323 (N_18323,N_17226,N_16179);
and U18324 (N_18324,N_17710,N_16976);
and U18325 (N_18325,N_16834,N_17005);
and U18326 (N_18326,N_16064,N_17325);
nand U18327 (N_18327,N_16932,N_17235);
or U18328 (N_18328,N_17508,N_17404);
or U18329 (N_18329,N_16359,N_16441);
nor U18330 (N_18330,N_16819,N_16243);
and U18331 (N_18331,N_17300,N_16323);
or U18332 (N_18332,N_16722,N_16263);
and U18333 (N_18333,N_17018,N_17466);
or U18334 (N_18334,N_17644,N_16382);
or U18335 (N_18335,N_16026,N_17128);
xor U18336 (N_18336,N_17548,N_17377);
and U18337 (N_18337,N_16547,N_17574);
and U18338 (N_18338,N_17449,N_16466);
or U18339 (N_18339,N_16656,N_16792);
or U18340 (N_18340,N_16889,N_17274);
or U18341 (N_18341,N_16655,N_17497);
nand U18342 (N_18342,N_16894,N_17899);
nor U18343 (N_18343,N_16536,N_16109);
nand U18344 (N_18344,N_16375,N_17138);
or U18345 (N_18345,N_16671,N_16532);
nor U18346 (N_18346,N_17867,N_17413);
nand U18347 (N_18347,N_16268,N_17341);
nand U18348 (N_18348,N_16708,N_16798);
and U18349 (N_18349,N_16801,N_17977);
nand U18350 (N_18350,N_16817,N_17565);
or U18351 (N_18351,N_16242,N_16014);
or U18352 (N_18352,N_16754,N_16195);
nor U18353 (N_18353,N_17861,N_16761);
or U18354 (N_18354,N_16632,N_17113);
xor U18355 (N_18355,N_16918,N_16021);
nand U18356 (N_18356,N_16305,N_17453);
and U18357 (N_18357,N_17885,N_16037);
nor U18358 (N_18358,N_17922,N_17112);
nor U18359 (N_18359,N_17566,N_17426);
and U18360 (N_18360,N_16212,N_17800);
nor U18361 (N_18361,N_16746,N_17876);
and U18362 (N_18362,N_17122,N_17166);
or U18363 (N_18363,N_17674,N_17602);
nand U18364 (N_18364,N_17655,N_16939);
nand U18365 (N_18365,N_17666,N_17312);
xnor U18366 (N_18366,N_17219,N_16004);
nand U18367 (N_18367,N_17047,N_16128);
and U18368 (N_18368,N_17570,N_16092);
and U18369 (N_18369,N_17193,N_17078);
or U18370 (N_18370,N_16196,N_16557);
or U18371 (N_18371,N_17484,N_16186);
and U18372 (N_18372,N_16034,N_17932);
and U18373 (N_18373,N_17835,N_16271);
or U18374 (N_18374,N_17914,N_17215);
nand U18375 (N_18375,N_16558,N_17399);
and U18376 (N_18376,N_17798,N_16083);
and U18377 (N_18377,N_16781,N_16901);
or U18378 (N_18378,N_17236,N_16309);
and U18379 (N_18379,N_16912,N_17979);
and U18380 (N_18380,N_16709,N_17966);
nand U18381 (N_18381,N_16843,N_17544);
nand U18382 (N_18382,N_17180,N_17227);
or U18383 (N_18383,N_16077,N_17794);
and U18384 (N_18384,N_17096,N_16213);
or U18385 (N_18385,N_17662,N_17459);
and U18386 (N_18386,N_16846,N_17392);
and U18387 (N_18387,N_17416,N_16586);
and U18388 (N_18388,N_16636,N_16926);
and U18389 (N_18389,N_17622,N_17494);
nor U18390 (N_18390,N_17659,N_17978);
nand U18391 (N_18391,N_17130,N_17361);
xor U18392 (N_18392,N_17838,N_16590);
nor U18393 (N_18393,N_16296,N_16141);
nand U18394 (N_18394,N_17603,N_16336);
and U18395 (N_18395,N_17646,N_16985);
nor U18396 (N_18396,N_17730,N_16690);
or U18397 (N_18397,N_17211,N_17578);
or U18398 (N_18398,N_17987,N_16094);
xnor U18399 (N_18399,N_16154,N_16515);
and U18400 (N_18400,N_16467,N_17927);
or U18401 (N_18401,N_17550,N_16624);
or U18402 (N_18402,N_16789,N_16956);
nand U18403 (N_18403,N_16560,N_17221);
nor U18404 (N_18404,N_16072,N_17349);
nor U18405 (N_18405,N_17723,N_17943);
nor U18406 (N_18406,N_17555,N_17024);
and U18407 (N_18407,N_16996,N_17811);
nor U18408 (N_18408,N_16506,N_17908);
xnor U18409 (N_18409,N_17639,N_17650);
or U18410 (N_18410,N_17841,N_17456);
or U18411 (N_18411,N_16119,N_16784);
nor U18412 (N_18412,N_16675,N_17391);
nor U18413 (N_18413,N_17684,N_17771);
xnor U18414 (N_18414,N_17015,N_17722);
or U18415 (N_18415,N_17148,N_16753);
nand U18416 (N_18416,N_16637,N_16658);
nand U18417 (N_18417,N_17330,N_16027);
nand U18418 (N_18418,N_17283,N_16480);
xor U18419 (N_18419,N_16451,N_16498);
xor U18420 (N_18420,N_16180,N_17257);
or U18421 (N_18421,N_16219,N_17847);
nand U18422 (N_18422,N_16576,N_17543);
nand U18423 (N_18423,N_17533,N_16062);
nand U18424 (N_18424,N_17601,N_17205);
and U18425 (N_18425,N_17721,N_17302);
or U18426 (N_18426,N_17422,N_16517);
or U18427 (N_18427,N_17920,N_16099);
nand U18428 (N_18428,N_17178,N_16173);
nand U18429 (N_18429,N_17082,N_17567);
and U18430 (N_18430,N_17428,N_16738);
nor U18431 (N_18431,N_17420,N_16121);
and U18432 (N_18432,N_16545,N_16042);
and U18433 (N_18433,N_16494,N_16457);
nor U18434 (N_18434,N_16076,N_16406);
or U18435 (N_18435,N_16875,N_17445);
nand U18436 (N_18436,N_16838,N_16799);
nand U18437 (N_18437,N_17967,N_16785);
nand U18438 (N_18438,N_17340,N_17146);
and U18439 (N_18439,N_17134,N_17407);
and U18440 (N_18440,N_17826,N_16854);
nand U18441 (N_18441,N_17496,N_17049);
nor U18442 (N_18442,N_17699,N_17784);
nand U18443 (N_18443,N_16218,N_17003);
and U18444 (N_18444,N_16945,N_16609);
xor U18445 (N_18445,N_17249,N_16500);
and U18446 (N_18446,N_16250,N_17244);
or U18447 (N_18447,N_16439,N_16566);
or U18448 (N_18448,N_17286,N_16018);
xnor U18449 (N_18449,N_16947,N_16936);
nor U18450 (N_18450,N_17689,N_16421);
and U18451 (N_18451,N_16414,N_17237);
or U18452 (N_18452,N_16523,N_16728);
nand U18453 (N_18453,N_17680,N_17911);
xor U18454 (N_18454,N_16986,N_17692);
nor U18455 (N_18455,N_16280,N_17225);
or U18456 (N_18456,N_16732,N_16156);
nor U18457 (N_18457,N_16765,N_17335);
and U18458 (N_18458,N_16472,N_17799);
and U18459 (N_18459,N_16701,N_17830);
nor U18460 (N_18460,N_17381,N_17194);
or U18461 (N_18461,N_17819,N_17803);
or U18462 (N_18462,N_17782,N_17443);
nand U18463 (N_18463,N_16929,N_17174);
nand U18464 (N_18464,N_16294,N_16319);
xor U18465 (N_18465,N_16188,N_17654);
nand U18466 (N_18466,N_16246,N_16606);
or U18467 (N_18467,N_17337,N_16458);
nand U18468 (N_18468,N_16962,N_17132);
nor U18469 (N_18469,N_16376,N_17757);
nor U18470 (N_18470,N_16262,N_16879);
xor U18471 (N_18471,N_16051,N_16192);
xnor U18472 (N_18472,N_17858,N_16908);
or U18473 (N_18473,N_16984,N_16995);
nor U18474 (N_18474,N_16233,N_16463);
nand U18475 (N_18475,N_17776,N_17432);
nand U18476 (N_18476,N_16454,N_17328);
nand U18477 (N_18477,N_17761,N_16512);
nand U18478 (N_18478,N_16604,N_17760);
or U18479 (N_18479,N_17437,N_17648);
or U18480 (N_18480,N_17740,N_16103);
nand U18481 (N_18481,N_16163,N_16931);
nor U18482 (N_18482,N_17828,N_17395);
nor U18483 (N_18483,N_16654,N_17902);
or U18484 (N_18484,N_16830,N_17822);
and U18485 (N_18485,N_16206,N_17421);
nand U18486 (N_18486,N_16899,N_16629);
nand U18487 (N_18487,N_16775,N_17538);
nand U18488 (N_18488,N_17787,N_16964);
and U18489 (N_18489,N_17663,N_16070);
or U18490 (N_18490,N_17971,N_17808);
and U18491 (N_18491,N_16227,N_17054);
nand U18492 (N_18492,N_16748,N_16320);
and U18493 (N_18493,N_17645,N_16123);
nand U18494 (N_18494,N_17458,N_16087);
or U18495 (N_18495,N_17975,N_17898);
nor U18496 (N_18496,N_17188,N_17104);
and U18497 (N_18497,N_17973,N_16149);
nor U18498 (N_18498,N_17469,N_16620);
and U18499 (N_18499,N_16047,N_16930);
nand U18500 (N_18500,N_17560,N_16065);
nand U18501 (N_18501,N_16866,N_17476);
or U18502 (N_18502,N_17880,N_17792);
or U18503 (N_18503,N_17232,N_16221);
nand U18504 (N_18504,N_17085,N_16239);
nand U18505 (N_18505,N_16395,N_17611);
xnor U18506 (N_18506,N_17970,N_17123);
nor U18507 (N_18507,N_17403,N_16223);
xor U18508 (N_18508,N_16143,N_16561);
and U18509 (N_18509,N_16770,N_17158);
nand U18510 (N_18510,N_17393,N_17915);
xnor U18511 (N_18511,N_17829,N_17728);
nor U18512 (N_18512,N_17216,N_17759);
or U18513 (N_18513,N_17091,N_17059);
and U18514 (N_18514,N_16052,N_17725);
xor U18515 (N_18515,N_17042,N_17549);
and U18516 (N_18516,N_17724,N_17323);
nand U18517 (N_18517,N_17857,N_17520);
or U18518 (N_18518,N_17487,N_16264);
and U18519 (N_18519,N_16461,N_17900);
nand U18520 (N_18520,N_17258,N_17507);
and U18521 (N_18521,N_17429,N_16994);
and U18522 (N_18522,N_16160,N_16847);
xor U18523 (N_18523,N_16685,N_16591);
or U18524 (N_18524,N_16565,N_17052);
or U18525 (N_18525,N_17461,N_17168);
nand U18526 (N_18526,N_17383,N_16324);
nor U18527 (N_18527,N_17686,N_16974);
or U18528 (N_18528,N_17907,N_16416);
and U18529 (N_18529,N_16522,N_17041);
or U18530 (N_18530,N_16352,N_16433);
nand U18531 (N_18531,N_16646,N_17658);
nand U18532 (N_18532,N_17498,N_16960);
and U18533 (N_18533,N_16356,N_16002);
nor U18534 (N_18534,N_17093,N_16061);
and U18535 (N_18535,N_16541,N_16321);
nor U18536 (N_18536,N_17631,N_16207);
nor U18537 (N_18537,N_17637,N_16334);
and U18538 (N_18538,N_17807,N_16339);
nand U18539 (N_18539,N_17163,N_16346);
nor U18540 (N_18540,N_16075,N_16501);
or U18541 (N_18541,N_17953,N_17571);
nand U18542 (N_18542,N_17825,N_16665);
and U18543 (N_18543,N_17719,N_17026);
nor U18544 (N_18544,N_17142,N_16773);
nor U18545 (N_18545,N_16909,N_17623);
nor U18546 (N_18546,N_17415,N_17398);
xnor U18547 (N_18547,N_17955,N_16849);
nand U18548 (N_18548,N_17842,N_16314);
nor U18549 (N_18549,N_16622,N_16777);
or U18550 (N_18550,N_16493,N_17647);
and U18551 (N_18551,N_16272,N_16893);
nor U18552 (N_18552,N_17672,N_17043);
nand U18553 (N_18553,N_16603,N_17373);
xor U18554 (N_18554,N_16380,N_17947);
and U18555 (N_18555,N_17539,N_17903);
nand U18556 (N_18556,N_17167,N_16097);
and U18557 (N_18557,N_16911,N_16644);
xor U18558 (N_18558,N_16437,N_17319);
nand U18559 (N_18559,N_16567,N_17610);
nor U18560 (N_18560,N_17370,N_16377);
xnor U18561 (N_18561,N_16020,N_17440);
or U18562 (N_18562,N_16587,N_16295);
nand U18563 (N_18563,N_17417,N_17460);
nand U18564 (N_18564,N_17772,N_16850);
nor U18565 (N_18565,N_17625,N_16577);
nor U18566 (N_18566,N_17834,N_17813);
nor U18567 (N_18567,N_16634,N_16332);
nor U18568 (N_18568,N_17316,N_17727);
nand U18569 (N_18569,N_16106,N_17952);
nand U18570 (N_18570,N_16120,N_16898);
or U18571 (N_18571,N_17293,N_17981);
nand U18572 (N_18572,N_16668,N_17388);
nor U18573 (N_18573,N_16484,N_16435);
nor U18574 (N_18574,N_16538,N_17097);
or U18575 (N_18575,N_17733,N_17928);
nor U18576 (N_18576,N_17633,N_17951);
and U18577 (N_18577,N_17233,N_17621);
xnor U18578 (N_18578,N_16756,N_17618);
or U18579 (N_18579,N_17950,N_17742);
or U18580 (N_18580,N_16527,N_16808);
and U18581 (N_18581,N_16892,N_17318);
and U18582 (N_18582,N_16667,N_17604);
nor U18583 (N_18583,N_17192,N_17714);
or U18584 (N_18584,N_16674,N_16231);
nand U18585 (N_18585,N_17941,N_16232);
or U18586 (N_18586,N_17505,N_17726);
or U18587 (N_18587,N_16344,N_16415);
nand U18588 (N_18588,N_17541,N_16858);
and U18589 (N_18589,N_17620,N_17500);
or U18590 (N_18590,N_17334,N_17796);
nand U18591 (N_18591,N_16514,N_16856);
nand U18592 (N_18592,N_17106,N_17752);
nor U18593 (N_18593,N_17299,N_16225);
or U18594 (N_18594,N_16712,N_16150);
or U18595 (N_18595,N_16340,N_16401);
and U18596 (N_18596,N_16261,N_16679);
or U18597 (N_18597,N_17285,N_16597);
and U18598 (N_18598,N_16145,N_17374);
nand U18599 (N_18599,N_16008,N_16378);
nand U18600 (N_18600,N_17853,N_16872);
xnor U18601 (N_18601,N_17435,N_17270);
and U18602 (N_18602,N_16530,N_16772);
nor U18603 (N_18603,N_16921,N_17181);
or U18604 (N_18604,N_16183,N_17457);
and U18605 (N_18605,N_17220,N_16621);
xnor U18606 (N_18606,N_17612,N_16693);
or U18607 (N_18607,N_17773,N_17695);
nand U18608 (N_18608,N_16327,N_17186);
nor U18609 (N_18609,N_16082,N_17536);
and U18610 (N_18610,N_17156,N_16998);
and U18611 (N_18611,N_17331,N_17372);
nor U18612 (N_18612,N_17255,N_17154);
or U18613 (N_18613,N_16987,N_16734);
and U18614 (N_18614,N_17777,N_16166);
and U18615 (N_18615,N_17806,N_16274);
xor U18616 (N_18616,N_16307,N_16164);
and U18617 (N_18617,N_16544,N_17965);
nor U18618 (N_18618,N_16736,N_17196);
and U18619 (N_18619,N_16951,N_16105);
or U18620 (N_18620,N_17878,N_16927);
nor U18621 (N_18621,N_16387,N_17653);
nor U18622 (N_18622,N_16368,N_17734);
or U18623 (N_18623,N_17562,N_17040);
and U18624 (N_18624,N_16596,N_16687);
nor U18625 (N_18625,N_16764,N_17576);
and U18626 (N_18626,N_16948,N_16895);
nor U18627 (N_18627,N_16438,N_16139);
xnor U18628 (N_18628,N_16652,N_16924);
xor U18629 (N_18629,N_17810,N_17879);
nor U18630 (N_18630,N_16703,N_16598);
nor U18631 (N_18631,N_17223,N_17942);
or U18632 (N_18632,N_17963,N_16548);
nand U18633 (N_18633,N_17704,N_16148);
and U18634 (N_18634,N_17521,N_16758);
or U18635 (N_18635,N_16471,N_17913);
nand U18636 (N_18636,N_17447,N_17008);
or U18637 (N_18637,N_16286,N_16535);
or U18638 (N_18638,N_16638,N_16298);
xor U18639 (N_18639,N_17100,N_17832);
and U18640 (N_18640,N_17375,N_16563);
and U18641 (N_18641,N_17821,N_17203);
nand U18642 (N_18642,N_17444,N_16526);
xor U18643 (N_18643,N_16197,N_16353);
or U18644 (N_18644,N_16842,N_17912);
nor U18645 (N_18645,N_17140,N_17119);
nor U18646 (N_18646,N_17202,N_16487);
and U18647 (N_18647,N_16900,N_16410);
nand U18648 (N_18648,N_17019,N_17528);
nor U18649 (N_18649,N_16060,N_16570);
or U18650 (N_18650,N_17485,N_17554);
or U18651 (N_18651,N_17268,N_16763);
and U18652 (N_18652,N_16275,N_16182);
nand U18653 (N_18653,N_17642,N_17087);
or U18654 (N_18654,N_16664,N_17242);
nand U18655 (N_18655,N_17120,N_17946);
xor U18656 (N_18656,N_16396,N_16607);
nor U18657 (N_18657,N_16711,N_16288);
and U18658 (N_18658,N_17251,N_17997);
and U18659 (N_18659,N_16136,N_16370);
nand U18660 (N_18660,N_17889,N_16661);
nor U18661 (N_18661,N_16193,N_17665);
or U18662 (N_18662,N_17598,N_16191);
and U18663 (N_18663,N_17580,N_17322);
xnor U18664 (N_18664,N_17785,N_17103);
and U18665 (N_18665,N_17384,N_16648);
nand U18666 (N_18666,N_17164,N_16714);
or U18667 (N_18667,N_17072,N_16745);
nor U18668 (N_18668,N_17783,N_17701);
and U18669 (N_18669,N_16181,N_17936);
nand U18670 (N_18670,N_16553,N_17883);
nand U18671 (N_18671,N_16331,N_16554);
or U18672 (N_18672,N_17960,N_16038);
and U18673 (N_18673,N_16628,N_16177);
xor U18674 (N_18674,N_16497,N_16793);
or U18675 (N_18675,N_17327,N_16290);
or U18676 (N_18676,N_17561,N_17594);
or U18677 (N_18677,N_16292,N_16750);
or U18678 (N_18678,N_17009,N_17010);
nor U18679 (N_18679,N_17718,N_17133);
xnor U18680 (N_18680,N_16673,N_17021);
xor U18681 (N_18681,N_16100,N_16876);
or U18682 (N_18682,N_16005,N_16682);
nand U18683 (N_18683,N_16432,N_17962);
nor U18684 (N_18684,N_16108,N_17157);
and U18685 (N_18685,N_17635,N_17552);
nor U18686 (N_18686,N_17529,N_17145);
and U18687 (N_18687,N_17172,N_16828);
nand U18688 (N_18688,N_16248,N_17006);
or U18689 (N_18689,N_17739,N_16814);
nor U18690 (N_18690,N_16786,N_17894);
nor U18691 (N_18691,N_17651,N_16725);
nor U18692 (N_18692,N_17789,N_16907);
and U18693 (N_18693,N_16919,N_17152);
and U18694 (N_18694,N_16482,N_16412);
nand U18695 (N_18695,N_16053,N_17289);
or U18696 (N_18696,N_17982,N_16573);
or U18697 (N_18697,N_17519,N_17124);
and U18698 (N_18698,N_16234,N_17764);
nand U18699 (N_18699,N_17736,N_17016);
and U18700 (N_18700,N_17182,N_16361);
or U18701 (N_18701,N_17276,N_17814);
nand U18702 (N_18702,N_17050,N_17563);
xor U18703 (N_18703,N_16862,N_16476);
nor U18704 (N_18704,N_16452,N_17114);
or U18705 (N_18705,N_16630,N_16341);
nand U18706 (N_18706,N_17864,N_16720);
or U18707 (N_18707,N_17369,N_17190);
nor U18708 (N_18708,N_16751,N_17887);
or U18709 (N_18709,N_17929,N_17062);
nand U18710 (N_18710,N_16318,N_17491);
or U18711 (N_18711,N_16550,N_17823);
nor U18712 (N_18712,N_17919,N_17873);
or U18713 (N_18713,N_16253,N_17472);
and U18714 (N_18714,N_16965,N_16012);
xor U18715 (N_18715,N_16608,N_16853);
or U18716 (N_18716,N_17342,N_16780);
or U18717 (N_18717,N_17102,N_16702);
or U18718 (N_18718,N_16943,N_17881);
or U18719 (N_18719,N_16388,N_16771);
nand U18720 (N_18720,N_16698,N_17455);
and U18721 (N_18721,N_17756,N_16993);
nand U18722 (N_18722,N_16001,N_16574);
or U18723 (N_18723,N_16721,N_16680);
or U18724 (N_18724,N_17073,N_16277);
or U18725 (N_18725,N_17489,N_17344);
nor U18726 (N_18726,N_16202,N_17767);
nor U18727 (N_18727,N_16046,N_16045);
xor U18728 (N_18728,N_17171,N_16134);
and U18729 (N_18729,N_17716,N_16966);
nand U18730 (N_18730,N_17371,N_16257);
nand U18731 (N_18731,N_16704,N_16282);
nor U18732 (N_18732,N_17218,N_17843);
and U18733 (N_18733,N_17267,N_17643);
nand U18734 (N_18734,N_16050,N_17886);
xor U18735 (N_18735,N_16079,N_17173);
nor U18736 (N_18736,N_17652,N_16351);
nand U18737 (N_18737,N_17070,N_17591);
and U18738 (N_18738,N_17115,N_16571);
xor U18739 (N_18739,N_16267,N_17418);
nor U18740 (N_18740,N_16691,N_16821);
or U18741 (N_18741,N_17117,N_17396);
or U18742 (N_18742,N_16408,N_17153);
nor U18743 (N_18743,N_16385,N_17315);
nand U18744 (N_18744,N_17679,N_17438);
nand U18745 (N_18745,N_17092,N_16582);
nand U18746 (N_18746,N_16811,N_16980);
or U18747 (N_18747,N_16118,N_17896);
nor U18748 (N_18748,N_17066,N_17866);
nor U18749 (N_18749,N_16583,N_16455);
or U18750 (N_18750,N_17380,N_17729);
or U18751 (N_18751,N_16524,N_17356);
xnor U18752 (N_18752,N_17446,N_16791);
nand U18753 (N_18753,N_16575,N_17326);
nor U18754 (N_18754,N_17599,N_16204);
or U18755 (N_18755,N_16959,N_17464);
nand U18756 (N_18756,N_16317,N_16755);
or U18757 (N_18757,N_16610,N_17547);
and U18758 (N_18758,N_17553,N_16006);
or U18759 (N_18759,N_17229,N_17353);
and U18760 (N_18760,N_16891,N_16483);
or U18761 (N_18761,N_16190,N_17793);
nor U18762 (N_18762,N_17522,N_16313);
or U18763 (N_18763,N_17993,N_17586);
nor U18764 (N_18764,N_16010,N_16245);
and U18765 (N_18765,N_17079,N_17360);
or U18766 (N_18766,N_16954,N_17988);
nand U18767 (N_18767,N_17582,N_17107);
or U18768 (N_18768,N_17791,N_16618);
or U18769 (N_18769,N_16258,N_17065);
or U18770 (N_18770,N_17159,N_17890);
nor U18771 (N_18771,N_16848,N_16474);
and U18772 (N_18772,N_17517,N_16308);
nand U18773 (N_18773,N_16896,N_16126);
nor U18774 (N_18774,N_17434,N_16731);
or U18775 (N_18775,N_17280,N_16914);
or U18776 (N_18776,N_16381,N_16759);
nor U18777 (N_18777,N_17569,N_17938);
nor U18778 (N_18778,N_16402,N_16405);
xor U18779 (N_18779,N_17290,N_17324);
or U18780 (N_18780,N_17317,N_16215);
nor U18781 (N_18781,N_16782,N_17032);
or U18782 (N_18782,N_17198,N_17542);
nand U18783 (N_18783,N_16127,N_16967);
nand U18784 (N_18784,N_16499,N_17406);
xnor U18785 (N_18785,N_17593,N_17036);
xor U18786 (N_18786,N_17931,N_17364);
nand U18787 (N_18787,N_17382,N_16531);
nor U18788 (N_18788,N_16266,N_17037);
nand U18789 (N_18789,N_16794,N_17660);
nand U18790 (N_18790,N_17664,N_17451);
nand U18791 (N_18791,N_16695,N_16937);
and U18792 (N_18792,N_16142,N_16226);
nand U18793 (N_18793,N_17080,N_16310);
xnor U18794 (N_18794,N_16642,N_17264);
nand U18795 (N_18795,N_17670,N_16559);
or U18796 (N_18796,N_17064,N_16869);
nor U18797 (N_18797,N_16623,N_16938);
nor U18798 (N_18798,N_17058,N_16845);
nor U18799 (N_18799,N_16403,N_16259);
and U18800 (N_18800,N_17863,N_16325);
and U18801 (N_18801,N_17254,N_17525);
nand U18802 (N_18802,N_16778,N_17063);
xnor U18803 (N_18803,N_16555,N_16740);
nor U18804 (N_18804,N_17801,N_16713);
nand U18805 (N_18805,N_16592,N_17513);
and U18806 (N_18806,N_16949,N_17486);
nand U18807 (N_18807,N_16633,N_16055);
and U18808 (N_18808,N_16933,N_17385);
xor U18809 (N_18809,N_16881,N_16973);
nor U18810 (N_18810,N_16659,N_16504);
xnor U18811 (N_18811,N_16138,N_17573);
and U18812 (N_18812,N_16859,N_17431);
and U18813 (N_18813,N_16743,N_16068);
or U18814 (N_18814,N_17204,N_16903);
nor U18815 (N_18815,N_17127,N_16116);
and U18816 (N_18816,N_16766,N_16102);
or U18817 (N_18817,N_17279,N_17846);
or U18818 (N_18818,N_17944,N_16017);
nand U18819 (N_18819,N_17926,N_16612);
and U18820 (N_18820,N_17004,N_16447);
nor U18821 (N_18821,N_16241,N_16373);
nor U18822 (N_18822,N_16000,N_17575);
or U18823 (N_18823,N_16140,N_16365);
and U18824 (N_18824,N_16857,N_17450);
nand U18825 (N_18825,N_16442,N_16113);
and U18826 (N_18826,N_16934,N_16279);
and U18827 (N_18827,N_17588,N_17248);
nor U18828 (N_18828,N_17661,N_16254);
nor U18829 (N_18829,N_17083,N_17854);
or U18830 (N_18830,N_17310,N_17940);
nor U18831 (N_18831,N_17365,N_17923);
nand U18832 (N_18832,N_17678,N_17071);
or U18833 (N_18833,N_16184,N_17209);
nand U18834 (N_18834,N_17616,N_16056);
or U18835 (N_18835,N_16639,N_16589);
nor U18836 (N_18836,N_16252,N_17860);
nand U18837 (N_18837,N_16922,N_17892);
nand U18838 (N_18838,N_16816,N_16157);
nand U18839 (N_18839,N_16832,N_17419);
nor U18840 (N_18840,N_17201,N_16117);
nand U18841 (N_18841,N_17077,N_16440);
nand U18842 (N_18842,N_16822,N_16477);
and U18843 (N_18843,N_16757,N_16681);
or U18844 (N_18844,N_16806,N_16371);
and U18845 (N_18845,N_17048,N_17408);
and U18846 (N_18846,N_17488,N_17238);
and U18847 (N_18847,N_17336,N_17707);
and U18848 (N_18848,N_17818,N_16886);
or U18849 (N_18849,N_17921,N_17630);
xor U18850 (N_18850,N_17273,N_16543);
nand U18851 (N_18851,N_16803,N_16626);
nand U18852 (N_18852,N_17613,N_17462);
xnor U18853 (N_18853,N_16465,N_16942);
or U18854 (N_18854,N_16430,N_16237);
nand U18855 (N_18855,N_17535,N_17998);
or U18856 (N_18856,N_16379,N_16877);
nand U18857 (N_18857,N_17409,N_16790);
or U18858 (N_18858,N_16542,N_16448);
and U18859 (N_18859,N_16222,N_16496);
nor U18860 (N_18860,N_17378,N_16510);
or U18861 (N_18861,N_17690,N_17020);
nand U18862 (N_18862,N_16677,N_16812);
xnor U18863 (N_18863,N_17430,N_17691);
or U18864 (N_18864,N_16019,N_16584);
or U18865 (N_18865,N_16443,N_16688);
or U18866 (N_18866,N_16429,N_17199);
or U18867 (N_18867,N_16384,N_16360);
and U18868 (N_18868,N_17871,N_17510);
nand U18869 (N_18869,N_16422,N_16831);
or U18870 (N_18870,N_16518,N_17833);
or U18871 (N_18871,N_17269,N_16905);
and U18872 (N_18872,N_17850,N_17101);
and U18873 (N_18873,N_17245,N_17839);
and U18874 (N_18874,N_17306,N_17139);
nor U18875 (N_18875,N_16970,N_17412);
or U18876 (N_18876,N_16979,N_16593);
nand U18877 (N_18877,N_17427,N_16165);
xor U18878 (N_18878,N_16710,N_17477);
and U18879 (N_18879,N_17667,N_17304);
nand U18880 (N_18880,N_17968,N_17301);
nor U18881 (N_18881,N_16367,N_16304);
and U18882 (N_18882,N_17605,N_17506);
xnor U18883 (N_18883,N_16733,N_17045);
nand U18884 (N_18884,N_16101,N_17657);
and U18885 (N_18885,N_17389,N_17595);
xor U18886 (N_18886,N_17681,N_17411);
or U18887 (N_18887,N_17002,N_16902);
nor U18888 (N_18888,N_16462,N_16492);
nor U18889 (N_18889,N_17572,N_17584);
nor U18890 (N_18890,N_17749,N_17945);
xor U18891 (N_18891,N_17831,N_16073);
or U18892 (N_18892,N_16235,N_16479);
or U18893 (N_18893,N_16696,N_17983);
nor U18894 (N_18894,N_17197,N_17320);
nor U18895 (N_18895,N_17288,N_16093);
nand U18896 (N_18896,N_17677,N_16135);
and U18897 (N_18897,N_16653,N_17687);
nand U18898 (N_18898,N_16168,N_17397);
and U18899 (N_18899,N_16407,N_17144);
and U18900 (N_18900,N_16975,N_17875);
and U18901 (N_18901,N_16647,N_16306);
or U18902 (N_18902,N_16864,N_16807);
nand U18903 (N_18903,N_17376,N_17934);
nand U18904 (N_18904,N_16705,N_16997);
and U18905 (N_18905,N_16588,N_16874);
or U18906 (N_18906,N_16595,N_17061);
and U18907 (N_18907,N_16399,N_16923);
nand U18908 (N_18908,N_17859,N_16802);
or U18909 (N_18909,N_17208,N_16229);
xnor U18910 (N_18910,N_16600,N_17402);
nor U18911 (N_18911,N_17869,N_17872);
xnor U18912 (N_18912,N_16220,N_16397);
or U18913 (N_18913,N_16349,N_17989);
nor U18914 (N_18914,N_17492,N_17676);
and U18915 (N_18915,N_17809,N_17239);
nor U18916 (N_18916,N_16741,N_17095);
xor U18917 (N_18917,N_16805,N_17475);
nor U18918 (N_18918,N_17161,N_17893);
and U18919 (N_18919,N_17260,N_17241);
nor U18920 (N_18920,N_16706,N_17874);
nand U18921 (N_18921,N_17700,N_16511);
and U18922 (N_18922,N_17483,N_16796);
nor U18923 (N_18923,N_17629,N_17354);
or U18924 (N_18924,N_16039,N_16426);
and U18925 (N_18925,N_16155,N_16813);
nor U18926 (N_18926,N_17425,N_16915);
and U18927 (N_18927,N_16977,N_16676);
nand U18928 (N_18928,N_17351,N_17709);
nand U18929 (N_18929,N_16048,N_17183);
or U18930 (N_18930,N_17386,N_17780);
and U18931 (N_18931,N_16111,N_16730);
xor U18932 (N_18932,N_16747,N_16211);
and U18933 (N_18933,N_17627,N_16841);
xor U18934 (N_18934,N_17958,N_16718);
xor U18935 (N_18935,N_16953,N_17347);
nand U18936 (N_18936,N_16289,N_16178);
nor U18937 (N_18937,N_16533,N_16418);
and U18938 (N_18938,N_17297,N_17474);
or U18939 (N_18939,N_16209,N_16534);
and U18940 (N_18940,N_16345,N_16090);
nor U18941 (N_18941,N_16199,N_16920);
and U18942 (N_18942,N_16080,N_16605);
and U18943 (N_18943,N_16906,N_16284);
xnor U18944 (N_18944,N_17698,N_17169);
or U18945 (N_18945,N_16364,N_16694);
nor U18946 (N_18946,N_17177,N_17277);
or U18947 (N_18947,N_16957,N_16335);
nand U18948 (N_18948,N_16469,N_17271);
and U18949 (N_18949,N_17515,N_16158);
and U18950 (N_18950,N_17779,N_17985);
and U18951 (N_18951,N_16281,N_16326);
and U18952 (N_18952,N_16130,N_16516);
nor U18953 (N_18953,N_17682,N_16826);
and U18954 (N_18954,N_16453,N_17638);
and U18955 (N_18955,N_16578,N_16882);
nand U18956 (N_18956,N_17175,N_17731);
or U18957 (N_18957,N_16338,N_17509);
or U18958 (N_18958,N_17295,N_17098);
or U18959 (N_18959,N_17685,N_17433);
nand U18960 (N_18960,N_17820,N_16958);
nand U18961 (N_18961,N_17282,N_16989);
and U18962 (N_18962,N_16488,N_17151);
nor U18963 (N_18963,N_16752,N_17350);
nand U18964 (N_18964,N_16398,N_17649);
xnor U18965 (N_18965,N_17636,N_16823);
and U18966 (N_18966,N_16490,N_17849);
nand U18967 (N_18967,N_17259,N_17250);
nand U18968 (N_18968,N_16776,N_16941);
xor U18969 (N_18969,N_17057,N_16299);
and U18970 (N_18970,N_17143,N_16700);
and U18971 (N_18971,N_16551,N_17478);
or U18972 (N_18972,N_16420,N_16444);
nor U18973 (N_18973,N_17141,N_16870);
nor U18974 (N_18974,N_17086,N_16669);
or U18975 (N_18975,N_16132,N_17482);
xor U18976 (N_18976,N_16175,N_16978);
and U18977 (N_18977,N_17632,N_17424);
and U18978 (N_18978,N_16078,N_16502);
and U18979 (N_18979,N_17596,N_16564);
or U18980 (N_18980,N_16887,N_17291);
nor U18981 (N_18981,N_16152,N_16343);
and U18982 (N_18982,N_16884,N_17410);
or U18983 (N_18983,N_17252,N_17094);
or U18984 (N_18984,N_16337,N_17439);
or U18985 (N_18985,N_16273,N_16916);
or U18986 (N_18986,N_16925,N_17362);
or U18987 (N_18987,N_17957,N_17788);
nor U18988 (N_18988,N_17564,N_16208);
nand U18989 (N_18989,N_17540,N_16787);
nand U18990 (N_18990,N_17358,N_17247);
and U18991 (N_18991,N_17243,N_17294);
and U18992 (N_18992,N_16129,N_17099);
nand U18993 (N_18993,N_16505,N_16650);
nor U18994 (N_18994,N_16723,N_16990);
nor U18995 (N_18995,N_16460,N_17481);
and U18996 (N_18996,N_16007,N_16513);
and U18997 (N_18997,N_17228,N_17656);
or U18998 (N_18998,N_16797,N_16086);
nand U18999 (N_18999,N_16057,N_16615);
xor U19000 (N_19000,N_16629,N_16332);
nand U19001 (N_19001,N_16111,N_16144);
and U19002 (N_19002,N_17496,N_16988);
nor U19003 (N_19003,N_17393,N_17854);
or U19004 (N_19004,N_17485,N_17854);
nor U19005 (N_19005,N_16291,N_16944);
nor U19006 (N_19006,N_16888,N_17317);
and U19007 (N_19007,N_16975,N_17707);
nor U19008 (N_19008,N_17770,N_16684);
or U19009 (N_19009,N_17428,N_17859);
xnor U19010 (N_19010,N_16605,N_16436);
nor U19011 (N_19011,N_17223,N_16500);
nand U19012 (N_19012,N_16021,N_17879);
nor U19013 (N_19013,N_16403,N_16836);
xnor U19014 (N_19014,N_17234,N_17461);
or U19015 (N_19015,N_16992,N_16943);
xnor U19016 (N_19016,N_16326,N_16500);
nand U19017 (N_19017,N_16636,N_16689);
or U19018 (N_19018,N_17659,N_16640);
nor U19019 (N_19019,N_16664,N_17827);
or U19020 (N_19020,N_17264,N_17138);
and U19021 (N_19021,N_16391,N_16243);
nand U19022 (N_19022,N_17015,N_16725);
nand U19023 (N_19023,N_17272,N_17791);
nand U19024 (N_19024,N_17105,N_16283);
nor U19025 (N_19025,N_16730,N_17080);
nand U19026 (N_19026,N_17072,N_17550);
nor U19027 (N_19027,N_17518,N_16033);
xnor U19028 (N_19028,N_17516,N_16504);
or U19029 (N_19029,N_16319,N_16058);
nand U19030 (N_19030,N_17378,N_16430);
or U19031 (N_19031,N_16896,N_16003);
and U19032 (N_19032,N_16440,N_16840);
nor U19033 (N_19033,N_17107,N_16766);
nand U19034 (N_19034,N_17352,N_17466);
xnor U19035 (N_19035,N_16660,N_17866);
and U19036 (N_19036,N_16027,N_16289);
nand U19037 (N_19037,N_17015,N_16714);
and U19038 (N_19038,N_16299,N_16903);
nor U19039 (N_19039,N_17064,N_16673);
and U19040 (N_19040,N_17594,N_17718);
and U19041 (N_19041,N_16341,N_16938);
xor U19042 (N_19042,N_16418,N_17878);
xnor U19043 (N_19043,N_16173,N_17088);
or U19044 (N_19044,N_17373,N_17097);
nand U19045 (N_19045,N_16539,N_16110);
nand U19046 (N_19046,N_16828,N_16528);
and U19047 (N_19047,N_17267,N_17260);
xor U19048 (N_19048,N_16729,N_16644);
or U19049 (N_19049,N_16680,N_17127);
nor U19050 (N_19050,N_16065,N_16748);
xor U19051 (N_19051,N_16262,N_16966);
nand U19052 (N_19052,N_16858,N_17961);
xor U19053 (N_19053,N_17699,N_17114);
and U19054 (N_19054,N_17493,N_16440);
nand U19055 (N_19055,N_17171,N_17045);
nor U19056 (N_19056,N_17005,N_16601);
xor U19057 (N_19057,N_16760,N_16259);
nor U19058 (N_19058,N_16131,N_17021);
or U19059 (N_19059,N_16703,N_16108);
xor U19060 (N_19060,N_17185,N_17157);
nor U19061 (N_19061,N_17831,N_17934);
and U19062 (N_19062,N_16191,N_16021);
nor U19063 (N_19063,N_17440,N_17542);
xor U19064 (N_19064,N_17628,N_17640);
or U19065 (N_19065,N_16464,N_17256);
or U19066 (N_19066,N_16552,N_17431);
nand U19067 (N_19067,N_16991,N_16646);
nand U19068 (N_19068,N_16354,N_17558);
nor U19069 (N_19069,N_17956,N_16631);
nand U19070 (N_19070,N_17975,N_16063);
or U19071 (N_19071,N_16138,N_16814);
nor U19072 (N_19072,N_16775,N_16673);
or U19073 (N_19073,N_16143,N_17329);
or U19074 (N_19074,N_17500,N_17106);
nand U19075 (N_19075,N_16248,N_16311);
and U19076 (N_19076,N_16425,N_17268);
nor U19077 (N_19077,N_17971,N_16813);
and U19078 (N_19078,N_17688,N_16743);
or U19079 (N_19079,N_17242,N_17692);
nor U19080 (N_19080,N_16162,N_16890);
nor U19081 (N_19081,N_17692,N_17985);
or U19082 (N_19082,N_17376,N_17115);
or U19083 (N_19083,N_16473,N_17993);
or U19084 (N_19084,N_16326,N_16088);
nand U19085 (N_19085,N_16961,N_16460);
nor U19086 (N_19086,N_16329,N_17155);
nand U19087 (N_19087,N_17166,N_17949);
nand U19088 (N_19088,N_16516,N_16169);
or U19089 (N_19089,N_16388,N_16621);
or U19090 (N_19090,N_17976,N_17747);
nand U19091 (N_19091,N_16981,N_17158);
nand U19092 (N_19092,N_17163,N_17696);
nor U19093 (N_19093,N_16409,N_16780);
xnor U19094 (N_19094,N_16125,N_16221);
and U19095 (N_19095,N_17172,N_16811);
nand U19096 (N_19096,N_16658,N_17976);
or U19097 (N_19097,N_16771,N_17654);
nand U19098 (N_19098,N_16908,N_16137);
or U19099 (N_19099,N_16169,N_16078);
or U19100 (N_19100,N_17986,N_17139);
nor U19101 (N_19101,N_17487,N_17522);
nand U19102 (N_19102,N_17703,N_16940);
nor U19103 (N_19103,N_16268,N_16657);
or U19104 (N_19104,N_17425,N_16518);
or U19105 (N_19105,N_16732,N_17488);
nor U19106 (N_19106,N_17862,N_17087);
and U19107 (N_19107,N_16080,N_17739);
or U19108 (N_19108,N_16541,N_17233);
xnor U19109 (N_19109,N_17508,N_16211);
nor U19110 (N_19110,N_16850,N_16517);
and U19111 (N_19111,N_16898,N_17382);
nor U19112 (N_19112,N_16896,N_16517);
nand U19113 (N_19113,N_16799,N_16806);
nor U19114 (N_19114,N_17517,N_17741);
or U19115 (N_19115,N_16869,N_17468);
or U19116 (N_19116,N_17027,N_16115);
xor U19117 (N_19117,N_17128,N_16213);
or U19118 (N_19118,N_16219,N_16758);
nor U19119 (N_19119,N_17728,N_17834);
nand U19120 (N_19120,N_17682,N_17383);
xnor U19121 (N_19121,N_17986,N_17882);
and U19122 (N_19122,N_16813,N_16088);
nor U19123 (N_19123,N_17152,N_16274);
and U19124 (N_19124,N_16500,N_16350);
nand U19125 (N_19125,N_17980,N_16850);
nor U19126 (N_19126,N_17045,N_17133);
nor U19127 (N_19127,N_16003,N_16795);
or U19128 (N_19128,N_17709,N_17406);
nor U19129 (N_19129,N_16643,N_17735);
or U19130 (N_19130,N_16565,N_16589);
and U19131 (N_19131,N_17704,N_16774);
nand U19132 (N_19132,N_16708,N_17559);
nand U19133 (N_19133,N_16988,N_17897);
xnor U19134 (N_19134,N_16762,N_17254);
or U19135 (N_19135,N_17984,N_17741);
nand U19136 (N_19136,N_17125,N_17985);
or U19137 (N_19137,N_16480,N_16551);
xor U19138 (N_19138,N_17700,N_16439);
and U19139 (N_19139,N_16483,N_16658);
or U19140 (N_19140,N_17523,N_17294);
nand U19141 (N_19141,N_16795,N_16137);
nor U19142 (N_19142,N_17729,N_16296);
nor U19143 (N_19143,N_17940,N_17169);
nor U19144 (N_19144,N_16124,N_16469);
nand U19145 (N_19145,N_16293,N_16677);
nor U19146 (N_19146,N_16127,N_16803);
and U19147 (N_19147,N_16578,N_16896);
nand U19148 (N_19148,N_16598,N_17469);
nor U19149 (N_19149,N_17283,N_17862);
nor U19150 (N_19150,N_17640,N_16163);
and U19151 (N_19151,N_16834,N_16551);
or U19152 (N_19152,N_17449,N_16982);
nand U19153 (N_19153,N_16092,N_16415);
nor U19154 (N_19154,N_17240,N_17442);
nand U19155 (N_19155,N_17519,N_17930);
nor U19156 (N_19156,N_16933,N_17521);
nand U19157 (N_19157,N_17112,N_16874);
nor U19158 (N_19158,N_16211,N_16208);
or U19159 (N_19159,N_16943,N_16672);
nand U19160 (N_19160,N_16777,N_17098);
and U19161 (N_19161,N_17324,N_17296);
nor U19162 (N_19162,N_16480,N_16335);
and U19163 (N_19163,N_16567,N_17318);
and U19164 (N_19164,N_17000,N_17820);
nor U19165 (N_19165,N_17014,N_16837);
nor U19166 (N_19166,N_16455,N_17833);
or U19167 (N_19167,N_17351,N_16741);
nor U19168 (N_19168,N_16989,N_16534);
nor U19169 (N_19169,N_16660,N_17409);
and U19170 (N_19170,N_16249,N_16206);
and U19171 (N_19171,N_17660,N_16105);
nor U19172 (N_19172,N_16712,N_16417);
and U19173 (N_19173,N_17832,N_17872);
and U19174 (N_19174,N_16340,N_17451);
nor U19175 (N_19175,N_17703,N_17666);
nand U19176 (N_19176,N_16807,N_17472);
and U19177 (N_19177,N_17209,N_16688);
xor U19178 (N_19178,N_16410,N_16705);
nand U19179 (N_19179,N_16617,N_16563);
nand U19180 (N_19180,N_16247,N_17753);
nand U19181 (N_19181,N_16851,N_16987);
nand U19182 (N_19182,N_17559,N_16984);
xnor U19183 (N_19183,N_17580,N_16611);
and U19184 (N_19184,N_16478,N_16461);
or U19185 (N_19185,N_17135,N_17855);
xnor U19186 (N_19186,N_17351,N_16023);
or U19187 (N_19187,N_16803,N_17079);
nor U19188 (N_19188,N_17851,N_16689);
or U19189 (N_19189,N_16515,N_16946);
nand U19190 (N_19190,N_17951,N_17725);
xnor U19191 (N_19191,N_16152,N_17613);
or U19192 (N_19192,N_17254,N_16237);
or U19193 (N_19193,N_17168,N_16624);
and U19194 (N_19194,N_17951,N_17940);
nor U19195 (N_19195,N_17255,N_17911);
and U19196 (N_19196,N_16284,N_16626);
or U19197 (N_19197,N_16654,N_17396);
and U19198 (N_19198,N_17356,N_17213);
or U19199 (N_19199,N_16273,N_16970);
nand U19200 (N_19200,N_16103,N_17055);
and U19201 (N_19201,N_16312,N_16938);
and U19202 (N_19202,N_16707,N_16954);
nor U19203 (N_19203,N_16751,N_17890);
nand U19204 (N_19204,N_16046,N_17272);
and U19205 (N_19205,N_17239,N_16281);
and U19206 (N_19206,N_16554,N_16973);
or U19207 (N_19207,N_17046,N_17655);
and U19208 (N_19208,N_17186,N_17258);
or U19209 (N_19209,N_17898,N_17874);
and U19210 (N_19210,N_16300,N_16005);
or U19211 (N_19211,N_17837,N_16748);
nor U19212 (N_19212,N_16627,N_17933);
or U19213 (N_19213,N_17646,N_17496);
and U19214 (N_19214,N_16059,N_17638);
nor U19215 (N_19215,N_17886,N_16364);
nand U19216 (N_19216,N_17495,N_17381);
xnor U19217 (N_19217,N_16453,N_17811);
or U19218 (N_19218,N_17823,N_17886);
and U19219 (N_19219,N_17537,N_16722);
or U19220 (N_19220,N_17180,N_17079);
or U19221 (N_19221,N_17301,N_16407);
nand U19222 (N_19222,N_16068,N_17244);
or U19223 (N_19223,N_16546,N_17656);
xnor U19224 (N_19224,N_16817,N_17398);
and U19225 (N_19225,N_16093,N_17921);
nand U19226 (N_19226,N_16407,N_16499);
nor U19227 (N_19227,N_17162,N_16275);
nor U19228 (N_19228,N_17205,N_16135);
and U19229 (N_19229,N_17707,N_17244);
and U19230 (N_19230,N_16088,N_16567);
and U19231 (N_19231,N_16031,N_17630);
and U19232 (N_19232,N_17058,N_16293);
nor U19233 (N_19233,N_16118,N_16996);
nor U19234 (N_19234,N_16775,N_17536);
or U19235 (N_19235,N_17171,N_17219);
or U19236 (N_19236,N_17320,N_16361);
or U19237 (N_19237,N_16714,N_17455);
nor U19238 (N_19238,N_16573,N_16229);
nor U19239 (N_19239,N_16102,N_16375);
and U19240 (N_19240,N_16621,N_17944);
nor U19241 (N_19241,N_16243,N_16424);
and U19242 (N_19242,N_17405,N_17968);
nand U19243 (N_19243,N_16685,N_16230);
xor U19244 (N_19244,N_17107,N_16535);
nand U19245 (N_19245,N_16017,N_17537);
and U19246 (N_19246,N_16069,N_16243);
or U19247 (N_19247,N_17057,N_16701);
and U19248 (N_19248,N_16084,N_16494);
nand U19249 (N_19249,N_17519,N_16911);
nor U19250 (N_19250,N_17560,N_17281);
or U19251 (N_19251,N_16586,N_17837);
and U19252 (N_19252,N_16860,N_16256);
nor U19253 (N_19253,N_16039,N_16107);
or U19254 (N_19254,N_17789,N_16007);
or U19255 (N_19255,N_16933,N_17337);
and U19256 (N_19256,N_16596,N_17655);
xor U19257 (N_19257,N_16635,N_17060);
xnor U19258 (N_19258,N_16101,N_16036);
or U19259 (N_19259,N_16970,N_16822);
xnor U19260 (N_19260,N_17912,N_16010);
and U19261 (N_19261,N_16706,N_16378);
and U19262 (N_19262,N_16525,N_16609);
nand U19263 (N_19263,N_16383,N_17755);
xnor U19264 (N_19264,N_17271,N_17818);
or U19265 (N_19265,N_16415,N_17022);
nor U19266 (N_19266,N_17596,N_17251);
nor U19267 (N_19267,N_16139,N_17147);
nor U19268 (N_19268,N_17925,N_17606);
or U19269 (N_19269,N_17640,N_16531);
nor U19270 (N_19270,N_16705,N_17297);
and U19271 (N_19271,N_16997,N_16826);
and U19272 (N_19272,N_16624,N_16810);
and U19273 (N_19273,N_17407,N_16646);
nor U19274 (N_19274,N_17259,N_17917);
nand U19275 (N_19275,N_17933,N_16883);
xnor U19276 (N_19276,N_16877,N_16414);
or U19277 (N_19277,N_16206,N_16755);
or U19278 (N_19278,N_17929,N_17289);
or U19279 (N_19279,N_16532,N_16380);
nor U19280 (N_19280,N_16932,N_16516);
nor U19281 (N_19281,N_17664,N_16091);
nand U19282 (N_19282,N_17398,N_17734);
nand U19283 (N_19283,N_17157,N_16345);
xor U19284 (N_19284,N_16330,N_16072);
and U19285 (N_19285,N_16259,N_17244);
nor U19286 (N_19286,N_16786,N_16966);
nand U19287 (N_19287,N_16942,N_17365);
nor U19288 (N_19288,N_17674,N_17416);
nand U19289 (N_19289,N_17634,N_16071);
and U19290 (N_19290,N_16680,N_17138);
nor U19291 (N_19291,N_16716,N_16894);
or U19292 (N_19292,N_17465,N_16726);
nor U19293 (N_19293,N_17873,N_17658);
nor U19294 (N_19294,N_17215,N_16095);
nor U19295 (N_19295,N_17175,N_17548);
nor U19296 (N_19296,N_17796,N_17934);
and U19297 (N_19297,N_17778,N_17267);
or U19298 (N_19298,N_17359,N_16943);
nand U19299 (N_19299,N_17316,N_17688);
nor U19300 (N_19300,N_16499,N_16238);
or U19301 (N_19301,N_16853,N_17073);
xnor U19302 (N_19302,N_17491,N_17362);
and U19303 (N_19303,N_17934,N_16215);
or U19304 (N_19304,N_17550,N_17290);
nand U19305 (N_19305,N_17159,N_17258);
or U19306 (N_19306,N_16973,N_17320);
nand U19307 (N_19307,N_16622,N_16404);
or U19308 (N_19308,N_16542,N_17488);
nand U19309 (N_19309,N_17110,N_17602);
and U19310 (N_19310,N_16953,N_16151);
nand U19311 (N_19311,N_17348,N_16011);
or U19312 (N_19312,N_17792,N_17031);
nand U19313 (N_19313,N_16792,N_17282);
nand U19314 (N_19314,N_16291,N_17067);
xnor U19315 (N_19315,N_16134,N_17917);
nand U19316 (N_19316,N_17240,N_17498);
or U19317 (N_19317,N_16410,N_16157);
nand U19318 (N_19318,N_16701,N_16447);
and U19319 (N_19319,N_16157,N_17302);
or U19320 (N_19320,N_16444,N_16291);
and U19321 (N_19321,N_16074,N_16203);
and U19322 (N_19322,N_16748,N_16087);
nor U19323 (N_19323,N_17502,N_17806);
and U19324 (N_19324,N_16307,N_17633);
nand U19325 (N_19325,N_17210,N_16907);
nand U19326 (N_19326,N_16798,N_17203);
or U19327 (N_19327,N_17625,N_17316);
or U19328 (N_19328,N_16113,N_16670);
nand U19329 (N_19329,N_16966,N_16439);
or U19330 (N_19330,N_17812,N_17950);
nor U19331 (N_19331,N_16806,N_16710);
nor U19332 (N_19332,N_16170,N_16252);
and U19333 (N_19333,N_16915,N_16077);
and U19334 (N_19334,N_16024,N_17712);
xnor U19335 (N_19335,N_16257,N_17415);
xnor U19336 (N_19336,N_17432,N_16792);
or U19337 (N_19337,N_16560,N_16475);
and U19338 (N_19338,N_16698,N_16931);
and U19339 (N_19339,N_16159,N_17021);
nand U19340 (N_19340,N_17970,N_17986);
and U19341 (N_19341,N_16481,N_17986);
nor U19342 (N_19342,N_16943,N_16064);
xor U19343 (N_19343,N_16109,N_17882);
nor U19344 (N_19344,N_17294,N_16076);
or U19345 (N_19345,N_17952,N_16226);
and U19346 (N_19346,N_17902,N_16413);
nand U19347 (N_19347,N_16190,N_16071);
and U19348 (N_19348,N_17189,N_16427);
nor U19349 (N_19349,N_16415,N_16639);
nand U19350 (N_19350,N_16574,N_17735);
nor U19351 (N_19351,N_17945,N_17596);
nor U19352 (N_19352,N_16615,N_17154);
or U19353 (N_19353,N_16038,N_17826);
and U19354 (N_19354,N_17868,N_16392);
and U19355 (N_19355,N_16456,N_17271);
xor U19356 (N_19356,N_16224,N_17324);
and U19357 (N_19357,N_17952,N_17069);
nand U19358 (N_19358,N_16948,N_16970);
nand U19359 (N_19359,N_16385,N_16014);
nand U19360 (N_19360,N_16580,N_17148);
xnor U19361 (N_19361,N_17332,N_17718);
and U19362 (N_19362,N_17164,N_17284);
or U19363 (N_19363,N_17628,N_17501);
nand U19364 (N_19364,N_16227,N_16213);
xor U19365 (N_19365,N_16152,N_17989);
nand U19366 (N_19366,N_16730,N_16404);
and U19367 (N_19367,N_16008,N_16949);
or U19368 (N_19368,N_17587,N_17110);
nand U19369 (N_19369,N_16671,N_17915);
or U19370 (N_19370,N_17355,N_17305);
xnor U19371 (N_19371,N_16856,N_16882);
nor U19372 (N_19372,N_16595,N_17452);
nor U19373 (N_19373,N_16479,N_16861);
nor U19374 (N_19374,N_17538,N_16532);
xor U19375 (N_19375,N_16447,N_17833);
nand U19376 (N_19376,N_16751,N_17971);
nor U19377 (N_19377,N_16960,N_17443);
xor U19378 (N_19378,N_17419,N_17187);
and U19379 (N_19379,N_16574,N_17991);
nor U19380 (N_19380,N_16451,N_17161);
nand U19381 (N_19381,N_16185,N_16146);
nor U19382 (N_19382,N_16184,N_16819);
nor U19383 (N_19383,N_17298,N_17978);
xor U19384 (N_19384,N_16678,N_17308);
nand U19385 (N_19385,N_17079,N_16355);
nand U19386 (N_19386,N_17427,N_16635);
nor U19387 (N_19387,N_16957,N_17572);
and U19388 (N_19388,N_17163,N_16611);
or U19389 (N_19389,N_16701,N_17085);
nor U19390 (N_19390,N_17584,N_17249);
or U19391 (N_19391,N_17479,N_17456);
nand U19392 (N_19392,N_17222,N_17536);
and U19393 (N_19393,N_17777,N_16728);
and U19394 (N_19394,N_17775,N_17506);
xnor U19395 (N_19395,N_16181,N_16010);
and U19396 (N_19396,N_16230,N_17217);
xnor U19397 (N_19397,N_17584,N_16508);
nand U19398 (N_19398,N_17406,N_16158);
nand U19399 (N_19399,N_17257,N_16439);
nand U19400 (N_19400,N_17196,N_17176);
or U19401 (N_19401,N_17335,N_17624);
nor U19402 (N_19402,N_17952,N_17292);
nand U19403 (N_19403,N_17436,N_16091);
and U19404 (N_19404,N_16230,N_17939);
nand U19405 (N_19405,N_16965,N_17065);
or U19406 (N_19406,N_16271,N_16660);
nor U19407 (N_19407,N_16619,N_17378);
nor U19408 (N_19408,N_16164,N_17713);
nand U19409 (N_19409,N_17411,N_16566);
nor U19410 (N_19410,N_17001,N_16762);
or U19411 (N_19411,N_17174,N_17031);
or U19412 (N_19412,N_16415,N_16696);
and U19413 (N_19413,N_17618,N_16602);
nor U19414 (N_19414,N_16118,N_16159);
or U19415 (N_19415,N_16518,N_17012);
and U19416 (N_19416,N_17981,N_17865);
nand U19417 (N_19417,N_16878,N_16627);
and U19418 (N_19418,N_16852,N_16406);
nor U19419 (N_19419,N_16628,N_17780);
nand U19420 (N_19420,N_17259,N_17770);
and U19421 (N_19421,N_16243,N_16421);
and U19422 (N_19422,N_17095,N_17329);
nand U19423 (N_19423,N_16686,N_17083);
and U19424 (N_19424,N_16702,N_17267);
or U19425 (N_19425,N_16218,N_17229);
and U19426 (N_19426,N_16854,N_16869);
and U19427 (N_19427,N_16024,N_16698);
and U19428 (N_19428,N_16585,N_16136);
xor U19429 (N_19429,N_17661,N_17793);
or U19430 (N_19430,N_17101,N_16381);
or U19431 (N_19431,N_16776,N_16925);
nand U19432 (N_19432,N_17318,N_17565);
xor U19433 (N_19433,N_16799,N_16625);
or U19434 (N_19434,N_16822,N_17914);
nand U19435 (N_19435,N_17042,N_16433);
or U19436 (N_19436,N_17597,N_16753);
and U19437 (N_19437,N_16732,N_17097);
and U19438 (N_19438,N_17818,N_17471);
nor U19439 (N_19439,N_16715,N_16535);
or U19440 (N_19440,N_16125,N_17123);
nor U19441 (N_19441,N_17228,N_17379);
or U19442 (N_19442,N_17678,N_16980);
nand U19443 (N_19443,N_16223,N_17378);
nand U19444 (N_19444,N_16275,N_16191);
nand U19445 (N_19445,N_17929,N_17875);
and U19446 (N_19446,N_16087,N_16410);
or U19447 (N_19447,N_17000,N_17681);
or U19448 (N_19448,N_17969,N_16589);
and U19449 (N_19449,N_17220,N_17140);
nand U19450 (N_19450,N_17332,N_16992);
nand U19451 (N_19451,N_17462,N_16167);
nor U19452 (N_19452,N_16899,N_16726);
or U19453 (N_19453,N_16528,N_16273);
nor U19454 (N_19454,N_16623,N_17117);
nand U19455 (N_19455,N_16096,N_16067);
nor U19456 (N_19456,N_17035,N_17713);
and U19457 (N_19457,N_16468,N_17811);
nor U19458 (N_19458,N_17891,N_17703);
nand U19459 (N_19459,N_16738,N_16024);
nand U19460 (N_19460,N_17714,N_17313);
or U19461 (N_19461,N_17796,N_16771);
or U19462 (N_19462,N_16911,N_17958);
or U19463 (N_19463,N_16868,N_16572);
nand U19464 (N_19464,N_17178,N_16748);
nand U19465 (N_19465,N_17145,N_17468);
nand U19466 (N_19466,N_16390,N_16658);
and U19467 (N_19467,N_17095,N_16470);
or U19468 (N_19468,N_17499,N_17950);
and U19469 (N_19469,N_16621,N_17878);
nor U19470 (N_19470,N_16264,N_16342);
nand U19471 (N_19471,N_16047,N_17005);
nor U19472 (N_19472,N_16562,N_16304);
nor U19473 (N_19473,N_17859,N_17377);
or U19474 (N_19474,N_16590,N_17060);
xnor U19475 (N_19475,N_16848,N_16451);
or U19476 (N_19476,N_17464,N_16579);
or U19477 (N_19477,N_16896,N_17695);
and U19478 (N_19478,N_16518,N_17600);
nor U19479 (N_19479,N_16453,N_16632);
nand U19480 (N_19480,N_16880,N_17732);
nand U19481 (N_19481,N_17446,N_16368);
or U19482 (N_19482,N_16236,N_17226);
xnor U19483 (N_19483,N_16156,N_17761);
or U19484 (N_19484,N_17066,N_16285);
xor U19485 (N_19485,N_16301,N_17388);
xor U19486 (N_19486,N_16187,N_17730);
xor U19487 (N_19487,N_16934,N_17753);
or U19488 (N_19488,N_17750,N_16677);
nand U19489 (N_19489,N_16222,N_16963);
and U19490 (N_19490,N_17460,N_17520);
nor U19491 (N_19491,N_17594,N_16518);
and U19492 (N_19492,N_17637,N_17186);
and U19493 (N_19493,N_17315,N_17291);
or U19494 (N_19494,N_16626,N_17636);
nor U19495 (N_19495,N_16008,N_16184);
nand U19496 (N_19496,N_16494,N_17042);
xor U19497 (N_19497,N_16652,N_16425);
nand U19498 (N_19498,N_16427,N_17913);
and U19499 (N_19499,N_17988,N_17891);
nor U19500 (N_19500,N_17349,N_16400);
nand U19501 (N_19501,N_16269,N_17773);
nand U19502 (N_19502,N_16362,N_16108);
nor U19503 (N_19503,N_17721,N_16055);
nand U19504 (N_19504,N_17361,N_17153);
or U19505 (N_19505,N_16558,N_17316);
and U19506 (N_19506,N_17888,N_17887);
and U19507 (N_19507,N_16163,N_17822);
or U19508 (N_19508,N_17763,N_16839);
nor U19509 (N_19509,N_17726,N_16793);
xnor U19510 (N_19510,N_17314,N_16885);
and U19511 (N_19511,N_16906,N_17440);
and U19512 (N_19512,N_16732,N_16244);
nand U19513 (N_19513,N_17625,N_17413);
and U19514 (N_19514,N_16426,N_16841);
and U19515 (N_19515,N_17971,N_16824);
nand U19516 (N_19516,N_16110,N_16525);
nand U19517 (N_19517,N_17047,N_16158);
nor U19518 (N_19518,N_17893,N_16721);
or U19519 (N_19519,N_17867,N_17639);
or U19520 (N_19520,N_16977,N_17986);
and U19521 (N_19521,N_16058,N_17984);
nand U19522 (N_19522,N_16372,N_16494);
xor U19523 (N_19523,N_16218,N_16279);
nor U19524 (N_19524,N_16006,N_17408);
or U19525 (N_19525,N_17696,N_17582);
or U19526 (N_19526,N_16043,N_17969);
and U19527 (N_19527,N_16940,N_17184);
nand U19528 (N_19528,N_16143,N_17702);
or U19529 (N_19529,N_17266,N_16503);
and U19530 (N_19530,N_16910,N_17929);
or U19531 (N_19531,N_16218,N_17426);
or U19532 (N_19532,N_16236,N_17454);
nand U19533 (N_19533,N_16041,N_16093);
or U19534 (N_19534,N_16221,N_17458);
and U19535 (N_19535,N_16544,N_17842);
nor U19536 (N_19536,N_17378,N_17891);
nor U19537 (N_19537,N_17861,N_16956);
or U19538 (N_19538,N_16966,N_17617);
nand U19539 (N_19539,N_17971,N_17004);
xnor U19540 (N_19540,N_17197,N_16982);
nand U19541 (N_19541,N_16721,N_16222);
and U19542 (N_19542,N_17814,N_16055);
and U19543 (N_19543,N_17376,N_17552);
or U19544 (N_19544,N_16408,N_16167);
nor U19545 (N_19545,N_17042,N_16672);
or U19546 (N_19546,N_16240,N_16961);
or U19547 (N_19547,N_16616,N_17065);
nand U19548 (N_19548,N_16253,N_16909);
and U19549 (N_19549,N_16333,N_16560);
nand U19550 (N_19550,N_16720,N_16894);
nand U19551 (N_19551,N_17011,N_16155);
and U19552 (N_19552,N_16661,N_16972);
and U19553 (N_19553,N_17393,N_17534);
nand U19554 (N_19554,N_16769,N_17492);
or U19555 (N_19555,N_17048,N_17036);
nand U19556 (N_19556,N_17123,N_16007);
xor U19557 (N_19557,N_17867,N_17109);
nor U19558 (N_19558,N_17015,N_16277);
or U19559 (N_19559,N_17184,N_17169);
nor U19560 (N_19560,N_16847,N_17592);
or U19561 (N_19561,N_17105,N_16792);
and U19562 (N_19562,N_17042,N_16918);
nor U19563 (N_19563,N_17789,N_16186);
nand U19564 (N_19564,N_17603,N_17269);
and U19565 (N_19565,N_16646,N_16494);
or U19566 (N_19566,N_16635,N_17432);
nand U19567 (N_19567,N_16876,N_16048);
nor U19568 (N_19568,N_16588,N_17968);
nor U19569 (N_19569,N_16326,N_17485);
nand U19570 (N_19570,N_16219,N_16108);
nand U19571 (N_19571,N_17348,N_17875);
xnor U19572 (N_19572,N_16502,N_16048);
and U19573 (N_19573,N_17387,N_16058);
nor U19574 (N_19574,N_16322,N_17404);
or U19575 (N_19575,N_16904,N_17445);
and U19576 (N_19576,N_16079,N_16051);
nor U19577 (N_19577,N_16005,N_17501);
or U19578 (N_19578,N_17262,N_16133);
or U19579 (N_19579,N_16473,N_17994);
or U19580 (N_19580,N_17944,N_16452);
nor U19581 (N_19581,N_17497,N_17289);
xnor U19582 (N_19582,N_17892,N_17913);
and U19583 (N_19583,N_16616,N_17118);
or U19584 (N_19584,N_16494,N_17923);
nor U19585 (N_19585,N_17043,N_17737);
and U19586 (N_19586,N_17480,N_17594);
and U19587 (N_19587,N_16112,N_17231);
nand U19588 (N_19588,N_17717,N_16698);
nor U19589 (N_19589,N_17479,N_16221);
nor U19590 (N_19590,N_17562,N_17316);
or U19591 (N_19591,N_17541,N_16704);
and U19592 (N_19592,N_17210,N_16469);
nor U19593 (N_19593,N_17595,N_17317);
nor U19594 (N_19594,N_16364,N_17957);
or U19595 (N_19595,N_17608,N_16534);
nand U19596 (N_19596,N_17806,N_17908);
or U19597 (N_19597,N_17387,N_16355);
and U19598 (N_19598,N_17467,N_17563);
nor U19599 (N_19599,N_16450,N_16426);
or U19600 (N_19600,N_16288,N_17115);
and U19601 (N_19601,N_17969,N_16033);
and U19602 (N_19602,N_17492,N_17678);
nor U19603 (N_19603,N_16737,N_16928);
nor U19604 (N_19604,N_16623,N_16459);
nand U19605 (N_19605,N_16573,N_16683);
or U19606 (N_19606,N_16389,N_16226);
xnor U19607 (N_19607,N_16835,N_17394);
and U19608 (N_19608,N_17153,N_17574);
and U19609 (N_19609,N_16116,N_16958);
and U19610 (N_19610,N_16579,N_17775);
nor U19611 (N_19611,N_17584,N_16505);
nor U19612 (N_19612,N_17158,N_16747);
nor U19613 (N_19613,N_16464,N_16075);
and U19614 (N_19614,N_17310,N_16320);
xnor U19615 (N_19615,N_17239,N_16024);
nand U19616 (N_19616,N_17207,N_17609);
xnor U19617 (N_19617,N_16900,N_17521);
and U19618 (N_19618,N_16555,N_17809);
nand U19619 (N_19619,N_16801,N_16432);
and U19620 (N_19620,N_16791,N_17449);
and U19621 (N_19621,N_16854,N_16982);
nor U19622 (N_19622,N_16973,N_16100);
nand U19623 (N_19623,N_16409,N_17272);
and U19624 (N_19624,N_16503,N_16910);
nand U19625 (N_19625,N_17466,N_17137);
nand U19626 (N_19626,N_17246,N_16424);
nor U19627 (N_19627,N_16549,N_17308);
and U19628 (N_19628,N_16375,N_17093);
nor U19629 (N_19629,N_17400,N_16315);
or U19630 (N_19630,N_16256,N_17050);
and U19631 (N_19631,N_17666,N_17808);
nor U19632 (N_19632,N_17833,N_16479);
and U19633 (N_19633,N_17498,N_17115);
nor U19634 (N_19634,N_16356,N_17010);
nand U19635 (N_19635,N_16539,N_17461);
nand U19636 (N_19636,N_16899,N_16305);
nand U19637 (N_19637,N_16342,N_16371);
and U19638 (N_19638,N_16756,N_16991);
and U19639 (N_19639,N_16423,N_16275);
nor U19640 (N_19640,N_16704,N_17112);
and U19641 (N_19641,N_17974,N_17095);
nor U19642 (N_19642,N_17586,N_17113);
or U19643 (N_19643,N_16209,N_16532);
nand U19644 (N_19644,N_17119,N_16121);
and U19645 (N_19645,N_17467,N_16588);
nor U19646 (N_19646,N_17790,N_16224);
and U19647 (N_19647,N_17864,N_16455);
or U19648 (N_19648,N_17880,N_16089);
and U19649 (N_19649,N_17046,N_17269);
and U19650 (N_19650,N_17973,N_16891);
and U19651 (N_19651,N_16402,N_17940);
nand U19652 (N_19652,N_16242,N_16749);
or U19653 (N_19653,N_17712,N_16957);
nor U19654 (N_19654,N_16241,N_16726);
or U19655 (N_19655,N_16663,N_17218);
and U19656 (N_19656,N_17614,N_16236);
nand U19657 (N_19657,N_17556,N_17064);
nand U19658 (N_19658,N_17742,N_16600);
nand U19659 (N_19659,N_16677,N_16199);
nor U19660 (N_19660,N_17566,N_16223);
nand U19661 (N_19661,N_16800,N_16413);
or U19662 (N_19662,N_16722,N_17708);
nand U19663 (N_19663,N_16341,N_17398);
xnor U19664 (N_19664,N_16083,N_17640);
and U19665 (N_19665,N_17548,N_16653);
and U19666 (N_19666,N_16927,N_16568);
nand U19667 (N_19667,N_17640,N_17772);
nand U19668 (N_19668,N_17428,N_17122);
or U19669 (N_19669,N_16293,N_17848);
xnor U19670 (N_19670,N_16964,N_16965);
nor U19671 (N_19671,N_16420,N_17668);
and U19672 (N_19672,N_16860,N_16838);
nor U19673 (N_19673,N_17741,N_17627);
xor U19674 (N_19674,N_16380,N_16918);
nor U19675 (N_19675,N_16078,N_17221);
nand U19676 (N_19676,N_16597,N_16088);
or U19677 (N_19677,N_17886,N_16279);
nor U19678 (N_19678,N_16923,N_17413);
nand U19679 (N_19679,N_17661,N_17460);
nor U19680 (N_19680,N_17603,N_17543);
and U19681 (N_19681,N_16580,N_17047);
nor U19682 (N_19682,N_17767,N_16741);
and U19683 (N_19683,N_16687,N_17826);
nor U19684 (N_19684,N_16658,N_17717);
and U19685 (N_19685,N_17583,N_17319);
nor U19686 (N_19686,N_17254,N_16445);
or U19687 (N_19687,N_16527,N_17949);
nand U19688 (N_19688,N_17367,N_17632);
nor U19689 (N_19689,N_16253,N_17512);
and U19690 (N_19690,N_16535,N_16244);
or U19691 (N_19691,N_16806,N_16240);
nand U19692 (N_19692,N_16476,N_17172);
or U19693 (N_19693,N_16350,N_17108);
nor U19694 (N_19694,N_17304,N_16390);
nor U19695 (N_19695,N_16737,N_17975);
nand U19696 (N_19696,N_17439,N_17423);
nor U19697 (N_19697,N_17476,N_17536);
or U19698 (N_19698,N_16041,N_17377);
nor U19699 (N_19699,N_17869,N_17721);
and U19700 (N_19700,N_17319,N_16020);
nand U19701 (N_19701,N_17731,N_16277);
and U19702 (N_19702,N_16634,N_17792);
and U19703 (N_19703,N_17531,N_16363);
nand U19704 (N_19704,N_17292,N_16001);
and U19705 (N_19705,N_16503,N_16034);
nor U19706 (N_19706,N_16754,N_17525);
nand U19707 (N_19707,N_16114,N_16246);
nor U19708 (N_19708,N_16008,N_16416);
and U19709 (N_19709,N_16488,N_16974);
nand U19710 (N_19710,N_16991,N_17587);
or U19711 (N_19711,N_16947,N_16110);
nand U19712 (N_19712,N_16758,N_16622);
and U19713 (N_19713,N_17037,N_16409);
xnor U19714 (N_19714,N_16066,N_17159);
and U19715 (N_19715,N_16455,N_17277);
nor U19716 (N_19716,N_17037,N_17225);
nor U19717 (N_19717,N_17080,N_16684);
nand U19718 (N_19718,N_17136,N_17462);
nand U19719 (N_19719,N_16583,N_17830);
or U19720 (N_19720,N_17889,N_16922);
nand U19721 (N_19721,N_17745,N_16215);
xnor U19722 (N_19722,N_17474,N_16014);
xor U19723 (N_19723,N_16835,N_17952);
xor U19724 (N_19724,N_17140,N_16093);
or U19725 (N_19725,N_16242,N_16576);
nor U19726 (N_19726,N_16352,N_17876);
or U19727 (N_19727,N_17517,N_17332);
and U19728 (N_19728,N_17193,N_16791);
or U19729 (N_19729,N_17991,N_17641);
nand U19730 (N_19730,N_16922,N_17581);
or U19731 (N_19731,N_17327,N_17188);
and U19732 (N_19732,N_16642,N_16346);
nor U19733 (N_19733,N_16875,N_17699);
nand U19734 (N_19734,N_16620,N_17456);
nand U19735 (N_19735,N_16402,N_17120);
or U19736 (N_19736,N_16231,N_17424);
nand U19737 (N_19737,N_17863,N_17521);
nand U19738 (N_19738,N_17231,N_17226);
or U19739 (N_19739,N_16144,N_16864);
and U19740 (N_19740,N_16632,N_16402);
and U19741 (N_19741,N_17752,N_16232);
and U19742 (N_19742,N_16985,N_17120);
and U19743 (N_19743,N_17063,N_16718);
and U19744 (N_19744,N_16559,N_16274);
nand U19745 (N_19745,N_16897,N_16305);
nand U19746 (N_19746,N_16964,N_16306);
nor U19747 (N_19747,N_16846,N_16190);
nand U19748 (N_19748,N_17789,N_17142);
or U19749 (N_19749,N_16687,N_16876);
and U19750 (N_19750,N_17819,N_17514);
nor U19751 (N_19751,N_16925,N_17570);
nand U19752 (N_19752,N_17987,N_16265);
and U19753 (N_19753,N_17036,N_16723);
nor U19754 (N_19754,N_17232,N_17329);
nand U19755 (N_19755,N_16407,N_17290);
xor U19756 (N_19756,N_16000,N_17206);
or U19757 (N_19757,N_17895,N_17293);
or U19758 (N_19758,N_17751,N_17470);
or U19759 (N_19759,N_16703,N_17313);
nor U19760 (N_19760,N_17240,N_16071);
and U19761 (N_19761,N_17711,N_16240);
xnor U19762 (N_19762,N_17714,N_16593);
xnor U19763 (N_19763,N_17703,N_17866);
or U19764 (N_19764,N_16664,N_16523);
nor U19765 (N_19765,N_17051,N_17355);
nand U19766 (N_19766,N_17064,N_17873);
or U19767 (N_19767,N_16258,N_16817);
nor U19768 (N_19768,N_17331,N_17864);
and U19769 (N_19769,N_16629,N_17232);
and U19770 (N_19770,N_16501,N_16372);
or U19771 (N_19771,N_17146,N_16288);
and U19772 (N_19772,N_16078,N_16997);
nand U19773 (N_19773,N_17724,N_16941);
xnor U19774 (N_19774,N_17257,N_17566);
nor U19775 (N_19775,N_17549,N_17457);
and U19776 (N_19776,N_16160,N_17081);
nand U19777 (N_19777,N_17160,N_17279);
nor U19778 (N_19778,N_17313,N_17045);
and U19779 (N_19779,N_16137,N_16692);
or U19780 (N_19780,N_17786,N_17082);
nand U19781 (N_19781,N_17854,N_17269);
and U19782 (N_19782,N_17343,N_17203);
nor U19783 (N_19783,N_16912,N_17578);
and U19784 (N_19784,N_16812,N_16464);
and U19785 (N_19785,N_17104,N_17410);
and U19786 (N_19786,N_16082,N_17531);
xor U19787 (N_19787,N_17521,N_17148);
nor U19788 (N_19788,N_17587,N_17028);
nor U19789 (N_19789,N_17709,N_17463);
nand U19790 (N_19790,N_17152,N_16983);
nor U19791 (N_19791,N_16059,N_17675);
nor U19792 (N_19792,N_16023,N_17147);
or U19793 (N_19793,N_16012,N_17302);
or U19794 (N_19794,N_16645,N_16819);
or U19795 (N_19795,N_16318,N_17882);
xor U19796 (N_19796,N_17832,N_17808);
and U19797 (N_19797,N_16017,N_16859);
and U19798 (N_19798,N_16706,N_17609);
nand U19799 (N_19799,N_16583,N_16513);
nand U19800 (N_19800,N_17972,N_17633);
xor U19801 (N_19801,N_17875,N_16525);
nor U19802 (N_19802,N_17967,N_16820);
or U19803 (N_19803,N_16526,N_16658);
and U19804 (N_19804,N_16856,N_16875);
or U19805 (N_19805,N_17619,N_17065);
nor U19806 (N_19806,N_17224,N_17592);
xnor U19807 (N_19807,N_17267,N_16633);
and U19808 (N_19808,N_17684,N_16656);
nor U19809 (N_19809,N_16815,N_17557);
or U19810 (N_19810,N_17100,N_16421);
nand U19811 (N_19811,N_17641,N_17598);
and U19812 (N_19812,N_16883,N_17889);
and U19813 (N_19813,N_16837,N_16407);
and U19814 (N_19814,N_17440,N_16817);
or U19815 (N_19815,N_16793,N_17102);
or U19816 (N_19816,N_16104,N_16816);
xor U19817 (N_19817,N_16290,N_16903);
nor U19818 (N_19818,N_17454,N_16901);
and U19819 (N_19819,N_17203,N_16871);
or U19820 (N_19820,N_17838,N_17827);
nor U19821 (N_19821,N_16595,N_16298);
or U19822 (N_19822,N_17657,N_16933);
or U19823 (N_19823,N_17082,N_16986);
or U19824 (N_19824,N_17409,N_17365);
or U19825 (N_19825,N_16518,N_16685);
nor U19826 (N_19826,N_17119,N_16938);
or U19827 (N_19827,N_17410,N_16875);
nor U19828 (N_19828,N_16978,N_16118);
xor U19829 (N_19829,N_16325,N_16069);
and U19830 (N_19830,N_17690,N_16024);
and U19831 (N_19831,N_17576,N_16681);
and U19832 (N_19832,N_16961,N_16399);
nand U19833 (N_19833,N_16567,N_17720);
nand U19834 (N_19834,N_17475,N_16521);
nor U19835 (N_19835,N_16062,N_16562);
xor U19836 (N_19836,N_17000,N_16229);
xor U19837 (N_19837,N_16798,N_17035);
xnor U19838 (N_19838,N_16700,N_17886);
nand U19839 (N_19839,N_16191,N_17702);
nor U19840 (N_19840,N_16425,N_16428);
nor U19841 (N_19841,N_16695,N_16543);
nor U19842 (N_19842,N_16114,N_16322);
or U19843 (N_19843,N_16974,N_16772);
and U19844 (N_19844,N_16555,N_16985);
and U19845 (N_19845,N_17441,N_17524);
nor U19846 (N_19846,N_17463,N_17337);
xnor U19847 (N_19847,N_16605,N_16402);
nand U19848 (N_19848,N_17742,N_16208);
nor U19849 (N_19849,N_16586,N_17657);
xor U19850 (N_19850,N_17320,N_16343);
and U19851 (N_19851,N_16939,N_16686);
nand U19852 (N_19852,N_17143,N_17586);
or U19853 (N_19853,N_16541,N_16445);
or U19854 (N_19854,N_17752,N_16004);
nor U19855 (N_19855,N_17234,N_17835);
xnor U19856 (N_19856,N_17187,N_17496);
and U19857 (N_19857,N_17913,N_16896);
nand U19858 (N_19858,N_16726,N_16764);
nand U19859 (N_19859,N_16474,N_17051);
and U19860 (N_19860,N_17443,N_16577);
and U19861 (N_19861,N_17903,N_17948);
and U19862 (N_19862,N_17858,N_16596);
nor U19863 (N_19863,N_16650,N_17917);
nand U19864 (N_19864,N_16059,N_17960);
nand U19865 (N_19865,N_17088,N_16145);
xor U19866 (N_19866,N_16651,N_16626);
nor U19867 (N_19867,N_17722,N_16610);
or U19868 (N_19868,N_16901,N_17614);
nand U19869 (N_19869,N_16971,N_17566);
nor U19870 (N_19870,N_17407,N_17378);
or U19871 (N_19871,N_17449,N_17940);
nor U19872 (N_19872,N_17278,N_17782);
nand U19873 (N_19873,N_16681,N_17942);
and U19874 (N_19874,N_17253,N_17735);
or U19875 (N_19875,N_16246,N_17311);
or U19876 (N_19876,N_17880,N_16420);
xor U19877 (N_19877,N_16262,N_17543);
or U19878 (N_19878,N_16024,N_16248);
nand U19879 (N_19879,N_16259,N_16333);
and U19880 (N_19880,N_16862,N_17976);
nand U19881 (N_19881,N_16145,N_17851);
or U19882 (N_19882,N_16998,N_16343);
nor U19883 (N_19883,N_16732,N_17474);
nand U19884 (N_19884,N_16358,N_17838);
nand U19885 (N_19885,N_16452,N_16827);
nor U19886 (N_19886,N_17877,N_16696);
nand U19887 (N_19887,N_17752,N_17300);
or U19888 (N_19888,N_17831,N_17042);
nand U19889 (N_19889,N_17347,N_17751);
or U19890 (N_19890,N_16454,N_16509);
or U19891 (N_19891,N_17806,N_16663);
and U19892 (N_19892,N_17887,N_16023);
and U19893 (N_19893,N_16009,N_16289);
or U19894 (N_19894,N_16886,N_16960);
nor U19895 (N_19895,N_17288,N_16897);
nor U19896 (N_19896,N_16936,N_16316);
or U19897 (N_19897,N_17220,N_16301);
and U19898 (N_19898,N_17822,N_17220);
nor U19899 (N_19899,N_16841,N_17543);
and U19900 (N_19900,N_17118,N_17244);
nor U19901 (N_19901,N_16666,N_17605);
nor U19902 (N_19902,N_17211,N_17298);
nor U19903 (N_19903,N_17804,N_16393);
nor U19904 (N_19904,N_17446,N_16259);
or U19905 (N_19905,N_16799,N_16431);
or U19906 (N_19906,N_16452,N_16635);
or U19907 (N_19907,N_17808,N_16050);
and U19908 (N_19908,N_16354,N_16120);
xnor U19909 (N_19909,N_17736,N_16574);
nand U19910 (N_19910,N_16510,N_16097);
nor U19911 (N_19911,N_16826,N_17191);
nor U19912 (N_19912,N_16582,N_17462);
nand U19913 (N_19913,N_17646,N_16347);
nand U19914 (N_19914,N_16856,N_16689);
nand U19915 (N_19915,N_16525,N_16817);
or U19916 (N_19916,N_16117,N_16281);
and U19917 (N_19917,N_17777,N_16376);
nand U19918 (N_19918,N_16208,N_17474);
and U19919 (N_19919,N_16662,N_17822);
or U19920 (N_19920,N_16020,N_16999);
and U19921 (N_19921,N_17240,N_17788);
nor U19922 (N_19922,N_16226,N_16310);
and U19923 (N_19923,N_17242,N_17115);
nor U19924 (N_19924,N_16725,N_17618);
nor U19925 (N_19925,N_17762,N_16884);
and U19926 (N_19926,N_16783,N_17635);
nand U19927 (N_19927,N_17135,N_16218);
and U19928 (N_19928,N_16097,N_17777);
and U19929 (N_19929,N_17650,N_17269);
nand U19930 (N_19930,N_16840,N_17888);
and U19931 (N_19931,N_16849,N_16426);
nand U19932 (N_19932,N_17311,N_16984);
nand U19933 (N_19933,N_17304,N_17518);
nand U19934 (N_19934,N_16772,N_16168);
nand U19935 (N_19935,N_17856,N_16423);
xnor U19936 (N_19936,N_16566,N_16438);
nor U19937 (N_19937,N_17081,N_17367);
nand U19938 (N_19938,N_17531,N_17897);
and U19939 (N_19939,N_17419,N_16758);
or U19940 (N_19940,N_16998,N_16291);
and U19941 (N_19941,N_16230,N_16401);
nand U19942 (N_19942,N_16704,N_17260);
nand U19943 (N_19943,N_17467,N_16460);
and U19944 (N_19944,N_17879,N_17863);
nand U19945 (N_19945,N_17827,N_16391);
nor U19946 (N_19946,N_17483,N_16194);
nand U19947 (N_19947,N_16353,N_17439);
or U19948 (N_19948,N_17831,N_17561);
and U19949 (N_19949,N_17376,N_16451);
or U19950 (N_19950,N_17905,N_17772);
or U19951 (N_19951,N_16024,N_17754);
nand U19952 (N_19952,N_17046,N_17167);
nor U19953 (N_19953,N_16069,N_17605);
and U19954 (N_19954,N_17731,N_17703);
xor U19955 (N_19955,N_16667,N_17044);
nor U19956 (N_19956,N_16634,N_16169);
nand U19957 (N_19957,N_16043,N_17851);
and U19958 (N_19958,N_17891,N_16850);
or U19959 (N_19959,N_17364,N_17780);
nand U19960 (N_19960,N_17084,N_16545);
nor U19961 (N_19961,N_16143,N_17020);
nand U19962 (N_19962,N_16440,N_17838);
nand U19963 (N_19963,N_17057,N_17956);
and U19964 (N_19964,N_17181,N_17308);
nor U19965 (N_19965,N_16274,N_17495);
or U19966 (N_19966,N_16809,N_16799);
nand U19967 (N_19967,N_16539,N_17449);
and U19968 (N_19968,N_17061,N_16364);
and U19969 (N_19969,N_17516,N_17816);
and U19970 (N_19970,N_17068,N_16638);
nor U19971 (N_19971,N_16668,N_16685);
xnor U19972 (N_19972,N_16907,N_16570);
and U19973 (N_19973,N_17802,N_17310);
nand U19974 (N_19974,N_16692,N_16388);
nand U19975 (N_19975,N_16306,N_17793);
nand U19976 (N_19976,N_16749,N_17610);
or U19977 (N_19977,N_16353,N_16403);
or U19978 (N_19978,N_17092,N_17535);
nor U19979 (N_19979,N_17964,N_16226);
nor U19980 (N_19980,N_16164,N_17617);
nor U19981 (N_19981,N_16484,N_17861);
xor U19982 (N_19982,N_16588,N_17428);
nand U19983 (N_19983,N_16953,N_17540);
nor U19984 (N_19984,N_16602,N_16733);
nor U19985 (N_19985,N_17056,N_16726);
nor U19986 (N_19986,N_16999,N_16517);
xor U19987 (N_19987,N_17822,N_16755);
nand U19988 (N_19988,N_16843,N_17569);
or U19989 (N_19989,N_17038,N_17127);
and U19990 (N_19990,N_17160,N_17540);
nand U19991 (N_19991,N_16311,N_16625);
nor U19992 (N_19992,N_16667,N_17913);
nor U19993 (N_19993,N_17075,N_17961);
or U19994 (N_19994,N_16229,N_17224);
and U19995 (N_19995,N_17947,N_16270);
nor U19996 (N_19996,N_16299,N_16569);
and U19997 (N_19997,N_16645,N_16087);
xnor U19998 (N_19998,N_16931,N_16137);
nor U19999 (N_19999,N_17300,N_17665);
xor UO_0 (O_0,N_18892,N_18985);
xor UO_1 (O_1,N_18949,N_19552);
nor UO_2 (O_2,N_18282,N_19563);
and UO_3 (O_3,N_19426,N_18764);
xnor UO_4 (O_4,N_18797,N_19770);
nand UO_5 (O_5,N_19903,N_18168);
nor UO_6 (O_6,N_19698,N_19713);
and UO_7 (O_7,N_19099,N_19080);
nor UO_8 (O_8,N_18679,N_18573);
nand UO_9 (O_9,N_19025,N_18906);
nor UO_10 (O_10,N_18186,N_18823);
or UO_11 (O_11,N_19685,N_18898);
nand UO_12 (O_12,N_19854,N_19248);
or UO_13 (O_13,N_18795,N_19406);
nor UO_14 (O_14,N_19879,N_18403);
nor UO_15 (O_15,N_18374,N_19888);
nor UO_16 (O_16,N_18369,N_18059);
nor UO_17 (O_17,N_18836,N_18465);
and UO_18 (O_18,N_19422,N_19533);
or UO_19 (O_19,N_19605,N_19768);
xnor UO_20 (O_20,N_18531,N_18382);
nand UO_21 (O_21,N_18212,N_19776);
or UO_22 (O_22,N_18775,N_19307);
nand UO_23 (O_23,N_19482,N_19984);
nor UO_24 (O_24,N_18504,N_19244);
nand UO_25 (O_25,N_18046,N_19038);
or UO_26 (O_26,N_18884,N_19300);
xnor UO_27 (O_27,N_18452,N_19928);
nor UO_28 (O_28,N_19336,N_19196);
and UO_29 (O_29,N_19208,N_18536);
nor UO_30 (O_30,N_19325,N_18998);
or UO_31 (O_31,N_18239,N_18977);
nor UO_32 (O_32,N_19131,N_18425);
or UO_33 (O_33,N_18125,N_18947);
nor UO_34 (O_34,N_18903,N_19610);
and UO_35 (O_35,N_19716,N_18523);
nand UO_36 (O_36,N_18589,N_18398);
xnor UO_37 (O_37,N_18195,N_19471);
or UO_38 (O_38,N_18311,N_18757);
or UO_39 (O_39,N_19026,N_18596);
nor UO_40 (O_40,N_18097,N_19875);
and UO_41 (O_41,N_18007,N_18950);
or UO_42 (O_42,N_19200,N_19091);
nor UO_43 (O_43,N_18216,N_19214);
or UO_44 (O_44,N_18624,N_18726);
and UO_45 (O_45,N_19298,N_19831);
nand UO_46 (O_46,N_18591,N_18876);
and UO_47 (O_47,N_19855,N_19400);
nand UO_48 (O_48,N_18146,N_19484);
or UO_49 (O_49,N_18151,N_18928);
nor UO_50 (O_50,N_19296,N_19227);
nand UO_51 (O_51,N_18451,N_18184);
and UO_52 (O_52,N_18122,N_18127);
nand UO_53 (O_53,N_19269,N_18912);
nor UO_54 (O_54,N_19281,N_18163);
or UO_55 (O_55,N_19741,N_18552);
xor UO_56 (O_56,N_18063,N_19228);
and UO_57 (O_57,N_19657,N_18684);
nand UO_58 (O_58,N_19184,N_18393);
and UO_59 (O_59,N_18844,N_19806);
or UO_60 (O_60,N_19763,N_18732);
nor UO_61 (O_61,N_18910,N_18780);
xnor UO_62 (O_62,N_18807,N_18816);
xnor UO_63 (O_63,N_19124,N_18991);
nor UO_64 (O_64,N_18677,N_19524);
and UO_65 (O_65,N_19593,N_18032);
nand UO_66 (O_66,N_19149,N_18025);
xnor UO_67 (O_67,N_18133,N_18703);
and UO_68 (O_68,N_18939,N_18649);
nand UO_69 (O_69,N_18568,N_19375);
or UO_70 (O_70,N_18368,N_18326);
and UO_71 (O_71,N_19377,N_18301);
nand UO_72 (O_72,N_19030,N_19122);
nand UO_73 (O_73,N_18512,N_19997);
nand UO_74 (O_74,N_19785,N_18572);
and UO_75 (O_75,N_19931,N_18073);
nor UO_76 (O_76,N_19632,N_18370);
nand UO_77 (O_77,N_19165,N_18197);
xor UO_78 (O_78,N_18538,N_19555);
nand UO_79 (O_79,N_18288,N_19316);
xor UO_80 (O_80,N_19711,N_19311);
xor UO_81 (O_81,N_18938,N_19023);
or UO_82 (O_82,N_19721,N_18148);
nand UO_83 (O_83,N_19364,N_19838);
nor UO_84 (O_84,N_18583,N_19367);
or UO_85 (O_85,N_19541,N_18668);
and UO_86 (O_86,N_19525,N_19852);
and UO_87 (O_87,N_19485,N_18312);
nor UO_88 (O_88,N_18830,N_18238);
and UO_89 (O_89,N_18774,N_19944);
or UO_90 (O_90,N_19608,N_18599);
nor UO_91 (O_91,N_19809,N_19047);
xnor UO_92 (O_92,N_18765,N_19127);
xnor UO_93 (O_93,N_18946,N_18894);
or UO_94 (O_94,N_18350,N_19851);
nand UO_95 (O_95,N_19144,N_18450);
nor UO_96 (O_96,N_19395,N_19386);
xnor UO_97 (O_97,N_18307,N_18172);
and UO_98 (O_98,N_18088,N_19847);
and UO_99 (O_99,N_18592,N_18325);
xnor UO_100 (O_100,N_19897,N_18331);
nand UO_101 (O_101,N_19789,N_19530);
or UO_102 (O_102,N_19719,N_18169);
nor UO_103 (O_103,N_18925,N_19784);
or UO_104 (O_104,N_19992,N_18192);
nor UO_105 (O_105,N_18587,N_18651);
xor UO_106 (O_106,N_18207,N_19217);
and UO_107 (O_107,N_19094,N_19684);
nand UO_108 (O_108,N_19727,N_19696);
xor UO_109 (O_109,N_19166,N_18700);
or UO_110 (O_110,N_18936,N_18029);
or UO_111 (O_111,N_19934,N_19020);
nand UO_112 (O_112,N_18755,N_19927);
xor UO_113 (O_113,N_19117,N_19415);
and UO_114 (O_114,N_19328,N_18824);
or UO_115 (O_115,N_19260,N_18296);
or UO_116 (O_116,N_18497,N_18786);
xnor UO_117 (O_117,N_19376,N_18385);
nor UO_118 (O_118,N_19832,N_18202);
and UO_119 (O_119,N_18174,N_19368);
or UO_120 (O_120,N_19305,N_19310);
and UO_121 (O_121,N_19947,N_18189);
and UO_122 (O_122,N_19141,N_18717);
nor UO_123 (O_123,N_18944,N_19417);
nor UO_124 (O_124,N_19050,N_18935);
or UO_125 (O_125,N_19173,N_18107);
and UO_126 (O_126,N_19892,N_19045);
xor UO_127 (O_127,N_18673,N_18772);
nand UO_128 (O_128,N_19686,N_19955);
and UO_129 (O_129,N_18188,N_18800);
nor UO_130 (O_130,N_19876,N_19858);
and UO_131 (O_131,N_18150,N_18843);
nand UO_132 (O_132,N_19941,N_19098);
and UO_133 (O_133,N_18616,N_18253);
and UO_134 (O_134,N_19546,N_18963);
or UO_135 (O_135,N_19724,N_19004);
nand UO_136 (O_136,N_19322,N_19354);
nand UO_137 (O_137,N_18631,N_18986);
nor UO_138 (O_138,N_19509,N_18476);
nor UO_139 (O_139,N_18295,N_18695);
or UO_140 (O_140,N_18955,N_18655);
xor UO_141 (O_141,N_18085,N_18462);
nand UO_142 (O_142,N_18853,N_19293);
nand UO_143 (O_143,N_18461,N_18023);
xor UO_144 (O_144,N_19407,N_18231);
and UO_145 (O_145,N_19845,N_19948);
xor UO_146 (O_146,N_19700,N_19040);
nor UO_147 (O_147,N_19914,N_18904);
nor UO_148 (O_148,N_19550,N_18094);
or UO_149 (O_149,N_18941,N_18054);
or UO_150 (O_150,N_18870,N_18246);
or UO_151 (O_151,N_18142,N_18579);
nor UO_152 (O_152,N_19528,N_19388);
nor UO_153 (O_153,N_19565,N_18916);
xnor UO_154 (O_154,N_18314,N_19604);
and UO_155 (O_155,N_18850,N_19430);
and UO_156 (O_156,N_19633,N_19839);
xor UO_157 (O_157,N_19522,N_18357);
or UO_158 (O_158,N_18056,N_19647);
nand UO_159 (O_159,N_19844,N_18598);
or UO_160 (O_160,N_18269,N_18068);
xnor UO_161 (O_161,N_19209,N_18584);
nor UO_162 (O_162,N_18860,N_19392);
and UO_163 (O_163,N_19474,N_19637);
nand UO_164 (O_164,N_19121,N_18496);
and UO_165 (O_165,N_19693,N_19722);
or UO_166 (O_166,N_18962,N_19545);
xnor UO_167 (O_167,N_19287,N_19601);
nand UO_168 (O_168,N_19044,N_18617);
nand UO_169 (O_169,N_18835,N_18091);
nor UO_170 (O_170,N_19924,N_19411);
nand UO_171 (O_171,N_19071,N_18447);
and UO_172 (O_172,N_18896,N_19365);
or UO_173 (O_173,N_19114,N_19507);
xnor UO_174 (O_174,N_19429,N_19115);
nand UO_175 (O_175,N_19453,N_18079);
or UO_176 (O_176,N_18338,N_19802);
nand UO_177 (O_177,N_18038,N_18967);
and UO_178 (O_178,N_18284,N_19569);
or UO_179 (O_179,N_18345,N_19245);
nand UO_180 (O_180,N_18981,N_19366);
or UO_181 (O_181,N_18656,N_18152);
nor UO_182 (O_182,N_18402,N_19405);
and UO_183 (O_183,N_18987,N_19884);
nor UO_184 (O_184,N_19046,N_18187);
xnor UO_185 (O_185,N_19495,N_19952);
and UO_186 (O_186,N_19758,N_18535);
and UO_187 (O_187,N_19615,N_18136);
nand UO_188 (O_188,N_18219,N_18638);
nand UO_189 (O_189,N_19451,N_19781);
and UO_190 (O_190,N_18057,N_18653);
nor UO_191 (O_191,N_19126,N_19929);
and UO_192 (O_192,N_19833,N_19480);
or UO_193 (O_193,N_19431,N_19512);
or UO_194 (O_194,N_19349,N_19280);
or UO_195 (O_195,N_19176,N_18305);
nor UO_196 (O_196,N_19382,N_18341);
xor UO_197 (O_197,N_18930,N_18522);
and UO_198 (O_198,N_18711,N_18802);
xor UO_199 (O_199,N_19402,N_19016);
nand UO_200 (O_200,N_19951,N_19194);
and UO_201 (O_201,N_19067,N_18926);
or UO_202 (O_202,N_19962,N_19606);
nor UO_203 (O_203,N_19408,N_19468);
nand UO_204 (O_204,N_19075,N_18490);
nor UO_205 (O_205,N_19666,N_18699);
nor UO_206 (O_206,N_19444,N_19065);
nor UO_207 (O_207,N_18053,N_18798);
xnor UO_208 (O_208,N_18893,N_19456);
nand UO_209 (O_209,N_18760,N_19599);
and UO_210 (O_210,N_18430,N_18229);
and UO_211 (O_211,N_19529,N_19619);
or UO_212 (O_212,N_19745,N_18126);
or UO_213 (O_213,N_19609,N_18316);
and UO_214 (O_214,N_19132,N_19225);
xor UO_215 (O_215,N_19889,N_19794);
and UO_216 (O_216,N_19972,N_18601);
or UO_217 (O_217,N_19500,N_18352);
and UO_218 (O_218,N_19488,N_18931);
nand UO_219 (O_219,N_18759,N_18101);
or UO_220 (O_220,N_18460,N_19201);
xor UO_221 (O_221,N_19345,N_19543);
nor UO_222 (O_222,N_19118,N_18849);
and UO_223 (O_223,N_19486,N_19425);
and UO_224 (O_224,N_19221,N_19873);
nor UO_225 (O_225,N_19380,N_19596);
nand UO_226 (O_226,N_19575,N_19597);
nor UO_227 (O_227,N_18273,N_19805);
xnor UO_228 (O_228,N_19971,N_19896);
nor UO_229 (O_229,N_18457,N_19949);
or UO_230 (O_230,N_18442,N_18173);
nor UO_231 (O_231,N_19714,N_19087);
nand UO_232 (O_232,N_19383,N_18344);
or UO_233 (O_233,N_19238,N_18734);
or UO_234 (O_234,N_19559,N_18483);
nand UO_235 (O_235,N_19229,N_18956);
nand UO_236 (O_236,N_18644,N_18381);
nand UO_237 (O_237,N_18575,N_19549);
nor UO_238 (O_238,N_19462,N_19769);
or UO_239 (O_239,N_18769,N_18562);
and UO_240 (O_240,N_19136,N_19164);
nor UO_241 (O_241,N_18116,N_18218);
nor UO_242 (O_242,N_18156,N_18102);
xor UO_243 (O_243,N_19547,N_18171);
nand UO_244 (O_244,N_18263,N_19317);
and UO_245 (O_245,N_18748,N_18449);
and UO_246 (O_246,N_18153,N_19578);
nand UO_247 (O_247,N_18105,N_18858);
or UO_248 (O_248,N_18399,N_18905);
nand UO_249 (O_249,N_19063,N_19454);
and UO_250 (O_250,N_19048,N_19301);
or UO_251 (O_251,N_19843,N_18020);
xnor UO_252 (O_252,N_19756,N_19133);
nor UO_253 (O_253,N_19906,N_18514);
or UO_254 (O_254,N_18128,N_19146);
nor UO_255 (O_255,N_18002,N_19796);
or UO_256 (O_256,N_19881,N_18782);
nand UO_257 (O_257,N_18328,N_18747);
nor UO_258 (O_258,N_19396,N_18866);
or UO_259 (O_259,N_18373,N_18453);
nor UO_260 (O_260,N_18559,N_18781);
nor UO_261 (O_261,N_18222,N_19324);
and UO_262 (O_262,N_18530,N_19108);
nand UO_263 (O_263,N_19678,N_19314);
xor UO_264 (O_264,N_19147,N_18232);
xnor UO_265 (O_265,N_18542,N_18175);
nor UO_266 (O_266,N_18001,N_19980);
nor UO_267 (O_267,N_19112,N_18294);
nor UO_268 (O_268,N_18489,N_19780);
xnor UO_269 (O_269,N_19557,N_19856);
or UO_270 (O_270,N_18048,N_18890);
and UO_271 (O_271,N_19148,N_19901);
nand UO_272 (O_272,N_18278,N_18570);
or UO_273 (O_273,N_18689,N_18167);
nand UO_274 (O_274,N_18268,N_18958);
nor UO_275 (O_275,N_19813,N_18141);
or UO_276 (O_276,N_19138,N_19640);
and UO_277 (O_277,N_18597,N_18907);
nand UO_278 (O_278,N_18335,N_18245);
and UO_279 (O_279,N_19340,N_18670);
nor UO_280 (O_280,N_18742,N_19007);
nand UO_281 (O_281,N_18756,N_18367);
or UO_282 (O_282,N_18664,N_18050);
nand UO_283 (O_283,N_18550,N_19394);
nor UO_284 (O_284,N_18543,N_19009);
and UO_285 (O_285,N_18193,N_18165);
or UO_286 (O_286,N_18293,N_19102);
nand UO_287 (O_287,N_19682,N_19461);
and UO_288 (O_288,N_18574,N_18793);
nor UO_289 (O_289,N_18720,N_18825);
nor UO_290 (O_290,N_18582,N_18723);
and UO_291 (O_291,N_18468,N_18407);
and UO_292 (O_292,N_19616,N_19241);
nor UO_293 (O_293,N_19932,N_18846);
or UO_294 (O_294,N_18770,N_19373);
nand UO_295 (O_295,N_19765,N_18082);
or UO_296 (O_296,N_18680,N_18934);
xor UO_297 (O_297,N_19926,N_18754);
nand UO_298 (O_298,N_19119,N_18889);
xor UO_299 (O_299,N_19329,N_19808);
or UO_300 (O_300,N_18060,N_19518);
and UO_301 (O_301,N_19819,N_18498);
or UO_302 (O_302,N_18832,N_19679);
or UO_303 (O_303,N_18516,N_18076);
xor UO_304 (O_304,N_19093,N_19441);
and UO_305 (O_305,N_19595,N_19537);
nor UO_306 (O_306,N_19308,N_19922);
and UO_307 (O_307,N_19022,N_18441);
nand UO_308 (O_308,N_18018,N_19729);
or UO_309 (O_309,N_18859,N_19639);
nand UO_310 (O_310,N_18017,N_18581);
xor UO_311 (O_311,N_18833,N_19983);
nand UO_312 (O_312,N_18886,N_19161);
or UO_313 (O_313,N_18940,N_19732);
or UO_314 (O_314,N_18276,N_19742);
and UO_315 (O_315,N_19150,N_19810);
nor UO_316 (O_316,N_19653,N_18267);
nor UO_317 (O_317,N_18790,N_18376);
or UO_318 (O_318,N_19977,N_18454);
nand UO_319 (O_319,N_18283,N_19379);
or UO_320 (O_320,N_19602,N_18387);
and UO_321 (O_321,N_18096,N_19583);
or UO_322 (O_322,N_19612,N_19627);
nand UO_323 (O_323,N_19690,N_19353);
or UO_324 (O_324,N_19899,N_19085);
nor UO_325 (O_325,N_19005,N_19869);
or UO_326 (O_326,N_19861,N_19918);
nand UO_327 (O_327,N_18829,N_18259);
nand UO_328 (O_328,N_18803,N_18157);
nand UO_329 (O_329,N_19982,N_19479);
and UO_330 (O_330,N_18610,N_19291);
xnor UO_331 (O_331,N_19076,N_19222);
and UO_332 (O_332,N_18751,N_18397);
or UO_333 (O_333,N_18473,N_19035);
nor UO_334 (O_334,N_18974,N_19759);
nand UO_335 (O_335,N_18196,N_18515);
xor UO_336 (O_336,N_19672,N_18456);
and UO_337 (O_337,N_18607,N_18084);
nor UO_338 (O_338,N_19830,N_19312);
and UO_339 (O_339,N_19239,N_19240);
nor UO_340 (O_340,N_19703,N_19018);
or UO_341 (O_341,N_18969,N_18628);
or UO_342 (O_342,N_19814,N_18671);
and UO_343 (O_343,N_19446,N_19309);
xor UO_344 (O_344,N_18380,N_18660);
and UO_345 (O_345,N_18182,N_18625);
and UO_346 (O_346,N_18405,N_19677);
xor UO_347 (O_347,N_19370,N_19659);
and UO_348 (O_348,N_18524,N_19634);
nand UO_349 (O_349,N_18036,N_18355);
and UO_350 (O_350,N_19723,N_19853);
nand UO_351 (O_351,N_18090,N_18132);
and UO_352 (O_352,N_18086,N_18459);
or UO_353 (O_353,N_18214,N_19804);
nor UO_354 (O_354,N_19937,N_18224);
and UO_355 (O_355,N_18565,N_18074);
nor UO_356 (O_356,N_18618,N_18155);
nand UO_357 (O_357,N_19074,N_18434);
and UO_358 (O_358,N_18089,N_19416);
nand UO_359 (O_359,N_18556,N_19635);
and UO_360 (O_360,N_18650,N_18724);
and UO_361 (O_361,N_19878,N_19348);
or UO_362 (O_362,N_19728,N_18863);
nor UO_363 (O_363,N_19061,N_19246);
or UO_364 (O_364,N_18736,N_18108);
and UO_365 (O_365,N_18111,N_18880);
xnor UO_366 (O_366,N_18292,N_18008);
or UO_367 (O_367,N_18640,N_19622);
xnor UO_368 (O_368,N_18822,N_19247);
xnor UO_369 (O_369,N_18227,N_19049);
or UO_370 (O_370,N_18487,N_18945);
nor UO_371 (O_371,N_19472,N_18394);
nand UO_372 (O_372,N_18612,N_18665);
or UO_373 (O_373,N_19381,N_18485);
or UO_374 (O_374,N_18069,N_19538);
and UO_375 (O_375,N_19198,N_18470);
nor UO_376 (O_376,N_18033,N_19999);
or UO_377 (O_377,N_19998,N_18594);
and UO_378 (O_378,N_18158,N_19514);
nand UO_379 (O_379,N_18404,N_19010);
or UO_380 (O_380,N_19154,N_18104);
or UO_381 (O_381,N_18633,N_18388);
nor UO_382 (O_382,N_19885,N_18563);
and UO_383 (O_383,N_18554,N_18537);
nand UO_384 (O_384,N_19318,N_18330);
nor UO_385 (O_385,N_19171,N_19687);
and UO_386 (O_386,N_18658,N_19330);
nand UO_387 (O_387,N_18098,N_18217);
or UO_388 (O_388,N_18569,N_18882);
xnor UO_389 (O_389,N_19515,N_19561);
xor UO_390 (O_390,N_19501,N_19335);
or UO_391 (O_391,N_19787,N_19337);
nand UO_392 (O_392,N_18488,N_18809);
xor UO_393 (O_393,N_18979,N_19439);
or UO_394 (O_394,N_18966,N_19420);
and UO_395 (O_395,N_18788,N_19737);
or UO_396 (O_396,N_19458,N_19798);
nor UO_397 (O_397,N_18455,N_19589);
nor UO_398 (O_398,N_19960,N_19865);
xnor UO_399 (O_399,N_18696,N_19907);
and UO_400 (O_400,N_18741,N_18354);
or UO_401 (O_401,N_18364,N_19128);
nand UO_402 (O_402,N_19579,N_19017);
and UO_403 (O_403,N_19333,N_18026);
nor UO_404 (O_404,N_18951,N_19925);
nand UO_405 (O_405,N_18279,N_19116);
nand UO_406 (O_406,N_18274,N_18205);
nand UO_407 (O_407,N_18828,N_19746);
or UO_408 (O_408,N_18315,N_19207);
nand UO_409 (O_409,N_19466,N_18852);
or UO_410 (O_410,N_19470,N_18166);
nand UO_411 (O_411,N_19504,N_18482);
and UO_412 (O_412,N_19827,N_18662);
nand UO_413 (O_413,N_19278,N_18261);
nand UO_414 (O_414,N_19034,N_18177);
and UO_415 (O_415,N_18702,N_18634);
or UO_416 (O_416,N_18719,N_18551);
and UO_417 (O_417,N_19103,N_18440);
and UO_418 (O_418,N_19275,N_18812);
nand UO_419 (O_419,N_19510,N_19398);
nor UO_420 (O_420,N_18810,N_19011);
or UO_421 (O_421,N_18300,N_18704);
and UO_422 (O_422,N_18716,N_19826);
nor UO_423 (O_423,N_19389,N_19674);
nand UO_424 (O_424,N_19232,N_19261);
and UO_425 (O_425,N_19978,N_18847);
xnor UO_426 (O_426,N_18078,N_18324);
xor UO_427 (O_427,N_18978,N_18100);
and UO_428 (O_428,N_19701,N_18766);
nand UO_429 (O_429,N_18045,N_19973);
or UO_430 (O_430,N_18528,N_18686);
xnor UO_431 (O_431,N_18725,N_18303);
nor UO_432 (O_432,N_19452,N_19497);
nand UO_433 (O_433,N_18432,N_18244);
nor UO_434 (O_434,N_18190,N_18281);
xor UO_435 (O_435,N_19641,N_19401);
nor UO_436 (O_436,N_18666,N_19192);
nor UO_437 (O_437,N_19707,N_19027);
xor UO_438 (O_438,N_19015,N_19862);
nor UO_439 (O_439,N_19006,N_19358);
nand UO_440 (O_440,N_19331,N_19863);
xor UO_441 (O_441,N_18873,N_19489);
nor UO_442 (O_442,N_18494,N_18900);
nor UO_443 (O_443,N_18801,N_18423);
and UO_444 (O_444,N_19857,N_18868);
or UO_445 (O_445,N_18710,N_18799);
and UO_446 (O_446,N_19264,N_19399);
or UO_447 (O_447,N_18840,N_18386);
nor UO_448 (O_448,N_19757,N_19848);
nor UO_449 (O_449,N_18749,N_19355);
nor UO_450 (O_450,N_18517,N_18051);
or UO_451 (O_451,N_19113,N_19079);
nand UO_452 (O_452,N_18577,N_19668);
xnor UO_453 (O_453,N_18879,N_19494);
and UO_454 (O_454,N_19777,N_18520);
or UO_455 (O_455,N_19297,N_18505);
and UO_456 (O_456,N_19288,N_18044);
nor UO_457 (O_457,N_19513,N_18871);
and UO_458 (O_458,N_18722,N_19823);
or UO_459 (O_459,N_19152,N_18922);
xor UO_460 (O_460,N_19267,N_19235);
nor UO_461 (O_461,N_18037,N_18285);
xnor UO_462 (O_462,N_19274,N_18917);
nand UO_463 (O_463,N_19553,N_18776);
and UO_464 (O_464,N_18421,N_19134);
nor UO_465 (O_465,N_19252,N_18995);
and UO_466 (O_466,N_19053,N_19302);
nor UO_467 (O_467,N_19012,N_19467);
nor UO_468 (O_468,N_18510,N_19361);
nand UO_469 (O_469,N_18433,N_18491);
and UO_470 (O_470,N_18435,N_19564);
and UO_471 (O_471,N_18789,N_19262);
nand UO_472 (O_472,N_18333,N_19846);
nor UO_473 (O_473,N_19097,N_19202);
nand UO_474 (O_474,N_18134,N_18137);
nand UO_475 (O_475,N_18304,N_19266);
nand UO_476 (O_476,N_18249,N_19059);
and UO_477 (O_477,N_18095,N_19435);
nand UO_478 (O_478,N_18874,N_19123);
nor UO_479 (O_479,N_19084,N_18123);
or UO_480 (O_480,N_18446,N_19705);
nand UO_481 (O_481,N_19570,N_18479);
nand UO_482 (O_482,N_19332,N_19576);
and UO_483 (O_483,N_18478,N_18384);
nand UO_484 (O_484,N_19508,N_19054);
nand UO_485 (O_485,N_19178,N_18061);
nor UO_486 (O_486,N_19111,N_19821);
and UO_487 (O_487,N_18181,N_19709);
and UO_488 (O_488,N_19950,N_19056);
xor UO_489 (O_489,N_18297,N_19975);
nand UO_490 (O_490,N_18558,N_19792);
or UO_491 (O_491,N_19943,N_18047);
nand UO_492 (O_492,N_19574,N_18201);
xnor UO_493 (O_493,N_19779,N_18511);
and UO_494 (O_494,N_18342,N_19391);
nor UO_495 (O_495,N_19195,N_19744);
nor UO_496 (O_496,N_18413,N_19219);
nand UO_497 (O_497,N_18667,N_19442);
nand UO_498 (O_498,N_18738,N_19129);
nor UO_499 (O_499,N_18337,N_19577);
nor UO_500 (O_500,N_18401,N_18897);
nand UO_501 (O_501,N_18444,N_18180);
nand UO_502 (O_502,N_18448,N_19213);
or UO_503 (O_503,N_19255,N_18106);
and UO_504 (O_504,N_18630,N_18340);
nor UO_505 (O_505,N_18529,N_18688);
and UO_506 (O_506,N_18773,N_18643);
or UO_507 (O_507,N_19959,N_18298);
nand UO_508 (O_508,N_18119,N_18021);
and UO_509 (O_509,N_18507,N_19284);
nand UO_510 (O_510,N_18383,N_18692);
and UO_511 (O_511,N_19940,N_18623);
xnor UO_512 (O_512,N_19880,N_18842);
xor UO_513 (O_513,N_18804,N_18299);
and UO_514 (O_514,N_19390,N_18112);
or UO_515 (O_515,N_18994,N_19650);
nand UO_516 (O_516,N_18013,N_18240);
nand UO_517 (O_517,N_19797,N_18428);
nand UO_518 (O_518,N_19180,N_18709);
xnor UO_519 (O_519,N_19938,N_18242);
nand UO_520 (O_520,N_18209,N_18877);
xor UO_521 (O_521,N_19476,N_18179);
nand UO_522 (O_522,N_19384,N_19702);
and UO_523 (O_523,N_18861,N_19321);
nand UO_524 (O_524,N_19460,N_19740);
nor UO_525 (O_525,N_19692,N_18458);
nand UO_526 (O_526,N_18960,N_18016);
nor UO_527 (O_527,N_18778,N_19360);
nor UO_528 (O_528,N_18645,N_18226);
nor UO_529 (O_529,N_18943,N_19436);
nor UO_530 (O_530,N_18302,N_18464);
or UO_531 (O_531,N_18851,N_19211);
or UO_532 (O_532,N_19469,N_19660);
xnor UO_533 (O_533,N_19204,N_19731);
xor UO_534 (O_534,N_18669,N_19694);
nand UO_535 (O_535,N_18415,N_18506);
nor UO_536 (O_536,N_19841,N_19893);
or UO_537 (O_537,N_19276,N_19057);
nor UO_538 (O_538,N_18837,N_19177);
nand UO_539 (O_539,N_18410,N_18009);
nor UO_540 (O_540,N_18614,N_18932);
nor UO_541 (O_541,N_18145,N_19673);
xnor UO_542 (O_542,N_19607,N_18663);
and UO_543 (O_543,N_18379,N_19440);
and UO_544 (O_544,N_18783,N_18595);
and UO_545 (O_545,N_18878,N_18675);
or UO_546 (O_546,N_18901,N_18883);
xnor UO_547 (O_547,N_18838,N_19532);
and UO_548 (O_548,N_19767,N_18888);
or UO_549 (O_549,N_19902,N_18864);
nand UO_550 (O_550,N_18475,N_19242);
nor UO_551 (O_551,N_18973,N_19662);
or UO_552 (O_552,N_19155,N_19945);
nor UO_553 (O_553,N_19062,N_19511);
or UO_554 (O_554,N_18493,N_19726);
nand UO_555 (O_555,N_18990,N_19104);
and UO_556 (O_556,N_18813,N_18919);
nor UO_557 (O_557,N_18211,N_19359);
or UO_558 (O_558,N_18336,N_19736);
nand UO_559 (O_559,N_18323,N_19306);
nor UO_560 (O_560,N_19362,N_19872);
nor UO_561 (O_561,N_18762,N_19226);
nor UO_562 (O_562,N_18289,N_18924);
nor UO_563 (O_563,N_18215,N_19556);
nor UO_564 (O_564,N_18982,N_18767);
or UO_565 (O_565,N_19670,N_18918);
nand UO_566 (O_566,N_18406,N_19378);
nor UO_567 (O_567,N_19755,N_18869);
xnor UO_568 (O_568,N_18080,N_18395);
nor UO_569 (O_569,N_19257,N_18015);
nand UO_570 (O_570,N_18120,N_19220);
and UO_571 (O_571,N_18721,N_19299);
nor UO_572 (O_572,N_18921,N_19712);
and UO_573 (O_573,N_18113,N_19088);
nand UO_574 (O_574,N_19648,N_18027);
and UO_575 (O_575,N_18989,N_19487);
nor UO_576 (O_576,N_18135,N_18234);
and UO_577 (O_577,N_18503,N_19423);
nand UO_578 (O_578,N_18039,N_18549);
and UO_579 (O_579,N_19935,N_18547);
xnor UO_580 (O_580,N_19942,N_19661);
nor UO_581 (O_581,N_19961,N_19969);
nor UO_582 (O_582,N_18431,N_18933);
nor UO_583 (O_583,N_19346,N_18247);
and UO_584 (O_584,N_19966,N_19558);
and UO_585 (O_585,N_19989,N_19542);
nor UO_586 (O_586,N_18280,N_18484);
or UO_587 (O_587,N_18701,N_18635);
nor UO_588 (O_588,N_18525,N_19990);
or UO_589 (O_589,N_18062,N_18971);
nand UO_590 (O_590,N_19140,N_19158);
nand UO_591 (O_591,N_19799,N_19970);
and UO_592 (O_592,N_19623,N_19503);
xnor UO_593 (O_593,N_18287,N_18855);
xor UO_594 (O_594,N_18400,N_19720);
or UO_595 (O_595,N_19531,N_19866);
nand UO_596 (O_596,N_19993,N_18103);
and UO_597 (O_597,N_19414,N_19174);
nand UO_598 (O_598,N_18839,N_19106);
and UO_599 (O_599,N_18541,N_19190);
nor UO_600 (O_600,N_18139,N_19807);
nor UO_601 (O_601,N_19652,N_19315);
nor UO_602 (O_602,N_18414,N_19151);
xor UO_603 (O_603,N_18213,N_19203);
nor UO_604 (O_604,N_19642,N_18983);
or UO_605 (O_605,N_18609,N_18006);
nor UO_606 (O_606,N_19663,N_19859);
and UO_607 (O_607,N_18109,N_18895);
and UO_608 (O_608,N_19828,N_18815);
or UO_609 (O_609,N_19153,N_18887);
and UO_610 (O_610,N_19976,N_18821);
or UO_611 (O_611,N_18463,N_18697);
and UO_612 (O_612,N_18619,N_19427);
or UO_613 (O_613,N_18391,N_18518);
and UO_614 (O_614,N_19762,N_18049);
or UO_615 (O_615,N_18237,N_18739);
xnor UO_616 (O_616,N_19029,N_18953);
nor UO_617 (O_617,N_18785,N_18183);
nand UO_618 (O_618,N_18746,N_19457);
or UO_619 (O_619,N_19582,N_18131);
or UO_620 (O_620,N_18480,N_18019);
nor UO_621 (O_621,N_19028,N_18003);
nor UO_622 (O_622,N_18492,N_19654);
or UO_623 (O_623,N_19667,N_19496);
or UO_624 (O_624,N_18499,N_19083);
nand UO_625 (O_625,N_19078,N_18024);
or UO_626 (O_626,N_18011,N_19372);
and UO_627 (O_627,N_18014,N_19988);
nand UO_628 (O_628,N_19070,N_19573);
or UO_629 (O_629,N_19754,N_18371);
and UO_630 (O_630,N_18262,N_18426);
nor UO_631 (O_631,N_18359,N_18648);
xnor UO_632 (O_632,N_19263,N_19024);
xor UO_633 (O_633,N_19385,N_18603);
and UO_634 (O_634,N_19697,N_19295);
xor UO_635 (O_635,N_19760,N_18272);
nand UO_636 (O_636,N_18392,N_18727);
nor UO_637 (O_637,N_18034,N_19717);
or UO_638 (O_638,N_19551,N_19630);
xnor UO_639 (O_639,N_19996,N_18814);
and UO_640 (O_640,N_18927,N_18681);
nand UO_641 (O_641,N_19793,N_19646);
nand UO_642 (O_642,N_19387,N_19735);
or UO_643 (O_643,N_18418,N_18817);
nor UO_644 (O_644,N_18682,N_19371);
and UO_645 (O_645,N_18412,N_19834);
nor UO_646 (O_646,N_19397,N_18743);
nand UO_647 (O_647,N_18834,N_19304);
nor UO_648 (O_648,N_18712,N_19636);
nor UO_649 (O_649,N_19393,N_19738);
or UO_650 (O_650,N_19064,N_18604);
and UO_651 (O_651,N_19891,N_19568);
and UO_652 (O_652,N_19651,N_18495);
or UO_653 (O_653,N_18143,N_18332);
nor UO_654 (O_654,N_18745,N_19042);
and UO_655 (O_655,N_19824,N_18339);
and UO_656 (O_656,N_19517,N_19268);
nor UO_657 (O_657,N_19739,N_18753);
nor UO_658 (O_658,N_19224,N_18613);
nor UO_659 (O_659,N_18124,N_19628);
nand UO_660 (O_660,N_18360,N_19279);
nand UO_661 (O_661,N_18486,N_18539);
nand UO_662 (O_662,N_19197,N_19188);
nor UO_663 (O_663,N_18540,N_19788);
nor UO_664 (O_664,N_19008,N_19991);
or UO_665 (O_665,N_19688,N_18225);
or UO_666 (O_666,N_19675,N_18993);
nand UO_667 (O_667,N_18768,N_18160);
or UO_668 (O_668,N_18477,N_18144);
and UO_669 (O_669,N_18526,N_18208);
nor UO_670 (O_670,N_18590,N_18358);
nand UO_671 (O_671,N_18417,N_19428);
nor UO_672 (O_672,N_18707,N_18848);
and UO_673 (O_673,N_19618,N_19871);
nor UO_674 (O_674,N_19412,N_18481);
nor UO_675 (O_675,N_19704,N_19052);
nand UO_676 (O_676,N_18257,N_19130);
and UO_677 (O_677,N_19643,N_19908);
nand UO_678 (O_678,N_19540,N_19236);
nand UO_679 (O_679,N_18318,N_19043);
nor UO_680 (O_680,N_18264,N_19464);
or UO_681 (O_681,N_19645,N_18954);
or UO_682 (O_682,N_18622,N_18500);
nand UO_683 (O_683,N_18690,N_19900);
nand UO_684 (O_684,N_19137,N_19905);
or UO_685 (O_685,N_19747,N_19327);
nand UO_686 (O_686,N_18221,N_19786);
nor UO_687 (O_687,N_19979,N_18980);
or UO_688 (O_688,N_18657,N_19560);
or UO_689 (O_689,N_19421,N_19483);
or UO_690 (O_690,N_19107,N_18564);
nand UO_691 (O_691,N_19438,N_18390);
xor UO_692 (O_692,N_19656,N_18715);
nor UO_693 (O_693,N_19303,N_18443);
or UO_694 (O_694,N_18593,N_18911);
or UO_695 (O_695,N_18731,N_19795);
xor UO_696 (O_696,N_18683,N_19058);
and UO_697 (O_697,N_18199,N_19783);
and UO_698 (O_698,N_19566,N_19320);
or UO_699 (O_699,N_18176,N_18642);
nor UO_700 (O_700,N_19644,N_19292);
and UO_701 (O_701,N_18277,N_18794);
and UO_702 (O_702,N_19895,N_18445);
nor UO_703 (O_703,N_19066,N_19521);
nor UO_704 (O_704,N_18066,N_19475);
and UO_705 (O_705,N_18411,N_19790);
nand UO_706 (O_706,N_19764,N_18422);
nor UO_707 (O_707,N_19041,N_18544);
or UO_708 (O_708,N_19586,N_19109);
or UO_709 (O_709,N_19424,N_19277);
or UO_710 (O_710,N_19254,N_18796);
or UO_711 (O_711,N_18820,N_19037);
xnor UO_712 (O_712,N_18698,N_18121);
xnor UO_713 (O_713,N_19933,N_18999);
and UO_714 (O_714,N_18178,N_19986);
nor UO_715 (O_715,N_19801,N_19936);
or UO_716 (O_716,N_18647,N_18586);
and UO_717 (O_717,N_19069,N_19710);
nand UO_718 (O_718,N_19032,N_18792);
nor UO_719 (O_719,N_19156,N_18308);
or UO_720 (O_720,N_18605,N_18959);
nand UO_721 (O_721,N_18872,N_19592);
nor UO_722 (O_722,N_19968,N_19625);
and UO_723 (O_723,N_18857,N_19139);
nor UO_724 (O_724,N_18952,N_19455);
xnor UO_725 (O_725,N_19909,N_18327);
xnor UO_726 (O_726,N_19774,N_19699);
nand UO_727 (O_727,N_19502,N_19708);
nor UO_728 (O_728,N_19974,N_19850);
and UO_729 (O_729,N_18291,N_19205);
nor UO_730 (O_730,N_19981,N_19733);
nor UO_731 (O_731,N_18248,N_19671);
nor UO_732 (O_732,N_19818,N_18845);
nand UO_733 (O_733,N_19752,N_19096);
nor UO_734 (O_734,N_19526,N_19413);
nor UO_735 (O_735,N_18714,N_18735);
nor UO_736 (O_736,N_19815,N_19077);
or UO_737 (O_737,N_18862,N_18317);
nand UO_738 (O_738,N_18972,N_19887);
nand UO_739 (O_739,N_18164,N_18970);
nand UO_740 (O_740,N_19985,N_18576);
nand UO_741 (O_741,N_19749,N_18865);
xnor UO_742 (O_742,N_18818,N_18705);
and UO_743 (O_743,N_18808,N_18022);
nand UO_744 (O_744,N_18042,N_19676);
nor UO_745 (O_745,N_18058,N_19539);
or UO_746 (O_746,N_18913,N_19167);
and UO_747 (O_747,N_18729,N_18161);
and UO_748 (O_748,N_19753,N_19917);
nor UO_749 (O_749,N_18375,N_18639);
nor UO_750 (O_750,N_19829,N_18602);
xor UO_751 (O_751,N_18265,N_18223);
xnor UO_752 (O_752,N_19882,N_19953);
nand UO_753 (O_753,N_18752,N_19168);
nor UO_754 (O_754,N_19505,N_19338);
nor UO_755 (O_755,N_18654,N_18353);
nor UO_756 (O_756,N_19816,N_18466);
xor UO_757 (O_757,N_18071,N_19915);
xnor UO_758 (O_758,N_18436,N_18929);
and UO_759 (O_759,N_19638,N_19344);
nor UO_760 (O_760,N_18637,N_18997);
nor UO_761 (O_761,N_19715,N_19215);
nor UO_762 (O_762,N_18902,N_19680);
nand UO_763 (O_763,N_18546,N_19939);
or UO_764 (O_764,N_18976,N_18320);
nand UO_765 (O_765,N_18310,N_18309);
xor UO_766 (O_766,N_19591,N_18501);
and UO_767 (O_767,N_19233,N_19664);
and UO_768 (O_768,N_19374,N_19230);
and UO_769 (O_769,N_18948,N_19534);
xnor UO_770 (O_770,N_19567,N_19039);
nand UO_771 (O_771,N_18521,N_18114);
xnor UO_772 (O_772,N_18419,N_18055);
nand UO_773 (O_773,N_19073,N_19285);
and UO_774 (O_774,N_19237,N_19342);
nor UO_775 (O_775,N_18676,N_19234);
nor UO_776 (O_776,N_18891,N_19142);
or UO_777 (O_777,N_18915,N_18409);
nand UO_778 (O_778,N_19621,N_19536);
or UO_779 (O_779,N_18129,N_18378);
and UO_780 (O_780,N_19867,N_18147);
nor UO_781 (O_781,N_19289,N_18140);
xnor UO_782 (O_782,N_19216,N_19270);
or UO_783 (O_783,N_18606,N_18138);
nor UO_784 (O_784,N_19181,N_18469);
nor UO_785 (O_785,N_19695,N_18957);
xor UO_786 (O_786,N_18099,N_19493);
xor UO_787 (O_787,N_19965,N_18509);
nand UO_788 (O_788,N_19434,N_19771);
nand UO_789 (O_789,N_19450,N_19210);
and UO_790 (O_790,N_19033,N_19051);
nand UO_791 (O_791,N_19191,N_19265);
nand UO_792 (O_792,N_19649,N_19135);
or UO_793 (O_793,N_19272,N_19437);
and UO_794 (O_794,N_19072,N_19620);
nor UO_795 (O_795,N_18416,N_19491);
nand UO_796 (O_796,N_19182,N_19572);
and UO_797 (O_797,N_18252,N_18854);
nor UO_798 (O_798,N_19223,N_18349);
and UO_799 (O_799,N_19187,N_18347);
nor UO_800 (O_800,N_19669,N_18004);
xnor UO_801 (O_801,N_18117,N_19987);
xor UO_802 (O_802,N_18975,N_19920);
or UO_803 (O_803,N_18693,N_19886);
and UO_804 (O_804,N_18661,N_18204);
nor UO_805 (O_805,N_19967,N_18270);
and UO_806 (O_806,N_18984,N_18322);
xor UO_807 (O_807,N_19842,N_19478);
nand UO_808 (O_808,N_19825,N_19357);
nor UO_809 (O_809,N_19527,N_19193);
and UO_810 (O_810,N_18694,N_18627);
xor UO_811 (O_811,N_19251,N_19750);
nor UO_812 (O_812,N_19002,N_19313);
and UO_813 (O_813,N_18115,N_18321);
and UO_814 (O_814,N_18708,N_18553);
and UO_815 (O_815,N_19773,N_19554);
or UO_816 (O_816,N_19082,N_19614);
nor UO_817 (O_817,N_18356,N_19352);
nor UO_818 (O_818,N_19588,N_19068);
nand UO_819 (O_819,N_19548,N_18787);
nor UO_820 (O_820,N_19145,N_19447);
or UO_821 (O_821,N_19751,N_19218);
or UO_822 (O_822,N_18674,N_19090);
nor UO_823 (O_823,N_18083,N_19913);
nand UO_824 (O_824,N_19160,N_19036);
nor UO_825 (O_825,N_19319,N_19820);
nand UO_826 (O_826,N_19419,N_18615);
xnor UO_827 (O_827,N_18611,N_19499);
and UO_828 (O_828,N_19930,N_19954);
nor UO_829 (O_829,N_19294,N_18149);
and UO_830 (O_830,N_19665,N_19734);
nand UO_831 (O_831,N_18629,N_18713);
nand UO_832 (O_832,N_19535,N_18641);
and UO_833 (O_833,N_19323,N_18233);
or UO_834 (O_834,N_18087,N_18608);
or UO_835 (O_835,N_18408,N_19580);
nor UO_836 (O_836,N_18899,N_18236);
or UO_837 (O_837,N_19590,N_18867);
and UO_838 (O_838,N_19498,N_19519);
and UO_839 (O_839,N_19860,N_19253);
nor UO_840 (O_840,N_18396,N_18361);
xnor UO_841 (O_841,N_19286,N_18365);
or UO_842 (O_842,N_18513,N_18914);
and UO_843 (O_843,N_18996,N_19101);
and UO_844 (O_844,N_18555,N_19271);
nand UO_845 (O_845,N_18621,N_19658);
nor UO_846 (O_846,N_18077,N_18093);
and UO_847 (O_847,N_19100,N_18961);
nor UO_848 (O_848,N_19086,N_19463);
or UO_849 (O_849,N_19350,N_18170);
nand UO_850 (O_850,N_19014,N_19683);
or UO_851 (O_851,N_18377,N_19157);
and UO_852 (O_852,N_19835,N_19243);
or UO_853 (O_853,N_19249,N_18081);
xor UO_854 (O_854,N_19169,N_19433);
nor UO_855 (O_855,N_18064,N_18965);
nor UO_856 (O_856,N_18784,N_18988);
nor UO_857 (O_857,N_19629,N_19912);
and UO_858 (O_858,N_18012,N_19743);
and UO_859 (O_859,N_18730,N_18306);
or UO_860 (O_860,N_19110,N_18652);
nor UO_861 (O_861,N_19778,N_19585);
nand UO_862 (O_862,N_18920,N_19347);
or UO_863 (O_863,N_19163,N_19341);
nand UO_864 (O_864,N_18343,N_18260);
or UO_865 (O_865,N_19811,N_19837);
xor UO_866 (O_866,N_19911,N_18439);
nand UO_867 (O_867,N_18366,N_18937);
or UO_868 (O_868,N_18241,N_19910);
xnor UO_869 (O_869,N_18040,N_18372);
nor UO_870 (O_870,N_19725,N_19766);
xnor UO_871 (O_871,N_18964,N_19631);
nand UO_872 (O_872,N_18256,N_18620);
nor UO_873 (O_873,N_18561,N_18750);
nor UO_874 (O_874,N_19031,N_18626);
and UO_875 (O_875,N_18718,N_18424);
and UO_876 (O_876,N_18758,N_19681);
or UO_877 (O_877,N_19506,N_18811);
or UO_878 (O_878,N_19143,N_18827);
nor UO_879 (O_879,N_19691,N_18243);
nor UO_880 (O_880,N_18043,N_19890);
nor UO_881 (O_881,N_18030,N_18251);
xor UO_882 (O_882,N_19864,N_19782);
nor UO_883 (O_883,N_19175,N_18545);
nor UO_884 (O_884,N_18533,N_18992);
xor UO_885 (O_885,N_18290,N_19125);
nand UO_886 (O_886,N_18075,N_19363);
and UO_887 (O_887,N_18130,N_18881);
nor UO_888 (O_888,N_18659,N_19877);
and UO_889 (O_889,N_18437,N_19520);
nand UO_890 (O_890,N_19105,N_18805);
and UO_891 (O_891,N_18968,N_19001);
nor UO_892 (O_892,N_19448,N_18346);
and UO_893 (O_893,N_19822,N_18200);
or UO_894 (O_894,N_18467,N_19817);
or UO_895 (O_895,N_19523,N_18072);
nor UO_896 (O_896,N_18194,N_19418);
and UO_897 (O_897,N_19339,N_19481);
and UO_898 (O_898,N_19800,N_19212);
and UO_899 (O_899,N_19995,N_19964);
nand UO_900 (O_900,N_18826,N_18052);
xnor UO_901 (O_901,N_18532,N_19730);
nand UO_902 (O_902,N_18438,N_18678);
nand UO_903 (O_903,N_19231,N_19812);
and UO_904 (O_904,N_19092,N_19445);
or UO_905 (O_905,N_19013,N_19273);
nand UO_906 (O_906,N_18571,N_18154);
and UO_907 (O_907,N_19283,N_19089);
nand UO_908 (O_908,N_19898,N_19613);
nor UO_909 (O_909,N_19000,N_19836);
or UO_910 (O_910,N_18031,N_19571);
or UO_911 (O_911,N_19256,N_19956);
xnor UO_912 (O_912,N_19868,N_18363);
and UO_913 (O_913,N_19994,N_18198);
and UO_914 (O_914,N_19410,N_19443);
or UO_915 (O_915,N_19775,N_19206);
nor UO_916 (O_916,N_18588,N_18472);
or UO_917 (O_917,N_18092,N_18389);
and UO_918 (O_918,N_18010,N_18474);
nand UO_919 (O_919,N_19957,N_18831);
nor UO_920 (O_920,N_18258,N_19748);
nand UO_921 (O_921,N_18000,N_19060);
and UO_922 (O_922,N_18908,N_18351);
or UO_923 (O_923,N_18067,N_18585);
or UO_924 (O_924,N_18646,N_19170);
and UO_925 (O_925,N_19334,N_19003);
nand UO_926 (O_926,N_19791,N_19516);
nor UO_927 (O_927,N_18266,N_19581);
nand UO_928 (O_928,N_19958,N_19282);
or UO_929 (O_929,N_19172,N_18471);
nand UO_930 (O_930,N_18744,N_18909);
nor UO_931 (O_931,N_19921,N_19250);
and UO_932 (O_932,N_18737,N_19326);
or UO_933 (O_933,N_18567,N_18041);
nor UO_934 (O_934,N_19021,N_19916);
nor UO_935 (O_935,N_18362,N_18636);
and UO_936 (O_936,N_18220,N_18875);
or UO_937 (O_937,N_18035,N_19803);
nor UO_938 (O_938,N_19562,N_19655);
and UO_939 (O_939,N_18206,N_18527);
nor UO_940 (O_940,N_19840,N_19095);
nand UO_941 (O_941,N_19883,N_18210);
or UO_942 (O_942,N_19598,N_19492);
and UO_943 (O_943,N_18329,N_19923);
or UO_944 (O_944,N_18761,N_18691);
nand UO_945 (O_945,N_19874,N_18763);
xor UO_946 (O_946,N_18508,N_19162);
and UO_947 (O_947,N_18162,N_18519);
or UO_948 (O_948,N_18191,N_19259);
or UO_949 (O_949,N_19189,N_18028);
or UO_950 (O_950,N_18841,N_19459);
nor UO_951 (O_951,N_18856,N_18806);
nand UO_952 (O_952,N_18334,N_19611);
or UO_953 (O_953,N_19477,N_19473);
or UO_954 (O_954,N_18230,N_18771);
and UO_955 (O_955,N_18566,N_18271);
nor UO_956 (O_956,N_19894,N_19544);
xor UO_957 (O_957,N_19179,N_19584);
nor UO_958 (O_958,N_18687,N_18942);
and UO_959 (O_959,N_18255,N_19019);
or UO_960 (O_960,N_19963,N_19403);
and UO_961 (O_961,N_19343,N_19258);
and UO_962 (O_962,N_18502,N_18672);
and UO_963 (O_963,N_19946,N_18728);
and UO_964 (O_964,N_19870,N_19369);
nand UO_965 (O_965,N_18600,N_18275);
nor UO_966 (O_966,N_18534,N_18313);
and UO_967 (O_967,N_19159,N_19055);
and UO_968 (O_968,N_19199,N_19449);
nand UO_969 (O_969,N_18819,N_19626);
nand UO_970 (O_970,N_18427,N_18348);
or UO_971 (O_971,N_18885,N_19183);
nor UO_972 (O_972,N_18923,N_19465);
xor UO_973 (O_973,N_18319,N_19603);
nor UO_974 (O_974,N_18159,N_18557);
or UO_975 (O_975,N_18065,N_19081);
xor UO_976 (O_976,N_18779,N_18733);
or UO_977 (O_977,N_19600,N_18632);
nand UO_978 (O_978,N_18548,N_19689);
and UO_979 (O_979,N_19587,N_18286);
or UO_980 (O_980,N_18560,N_18706);
nand UO_981 (O_981,N_18235,N_18580);
or UO_982 (O_982,N_18250,N_18429);
nor UO_983 (O_983,N_18740,N_19772);
or UO_984 (O_984,N_19351,N_18203);
and UO_985 (O_985,N_19186,N_19904);
and UO_986 (O_986,N_19706,N_19617);
or UO_987 (O_987,N_19761,N_19409);
nand UO_988 (O_988,N_18005,N_18185);
nor UO_989 (O_989,N_19624,N_18420);
or UO_990 (O_990,N_19356,N_18110);
and UO_991 (O_991,N_18254,N_19718);
nand UO_992 (O_992,N_18777,N_19919);
xor UO_993 (O_993,N_18578,N_19594);
or UO_994 (O_994,N_18070,N_19432);
xor UO_995 (O_995,N_19185,N_18228);
nand UO_996 (O_996,N_19490,N_19404);
or UO_997 (O_997,N_18118,N_19120);
nand UO_998 (O_998,N_19849,N_19290);
nor UO_999 (O_999,N_18685,N_18791);
and UO_1000 (O_1000,N_18829,N_19971);
and UO_1001 (O_1001,N_18708,N_19819);
nor UO_1002 (O_1002,N_19429,N_18089);
and UO_1003 (O_1003,N_18511,N_18983);
nor UO_1004 (O_1004,N_18771,N_18799);
and UO_1005 (O_1005,N_18355,N_18571);
xor UO_1006 (O_1006,N_18082,N_19485);
nor UO_1007 (O_1007,N_18481,N_18003);
nand UO_1008 (O_1008,N_18475,N_18655);
nor UO_1009 (O_1009,N_18813,N_18136);
nor UO_1010 (O_1010,N_18416,N_18409);
and UO_1011 (O_1011,N_19616,N_18260);
or UO_1012 (O_1012,N_19274,N_18952);
nand UO_1013 (O_1013,N_18577,N_18743);
and UO_1014 (O_1014,N_19771,N_18724);
and UO_1015 (O_1015,N_19498,N_19915);
nand UO_1016 (O_1016,N_18193,N_19346);
nor UO_1017 (O_1017,N_19021,N_18213);
xor UO_1018 (O_1018,N_18834,N_18370);
or UO_1019 (O_1019,N_18615,N_18007);
nor UO_1020 (O_1020,N_18421,N_18002);
nand UO_1021 (O_1021,N_18813,N_18553);
or UO_1022 (O_1022,N_19541,N_18205);
and UO_1023 (O_1023,N_18197,N_19466);
nor UO_1024 (O_1024,N_19644,N_18499);
nor UO_1025 (O_1025,N_18800,N_19984);
nand UO_1026 (O_1026,N_18401,N_19169);
or UO_1027 (O_1027,N_19538,N_19890);
and UO_1028 (O_1028,N_19893,N_18361);
and UO_1029 (O_1029,N_19915,N_19447);
and UO_1030 (O_1030,N_19491,N_18153);
xnor UO_1031 (O_1031,N_19143,N_18346);
nor UO_1032 (O_1032,N_18816,N_18618);
xor UO_1033 (O_1033,N_18712,N_19020);
and UO_1034 (O_1034,N_19956,N_18914);
or UO_1035 (O_1035,N_19028,N_18840);
or UO_1036 (O_1036,N_19963,N_19336);
nand UO_1037 (O_1037,N_19849,N_19910);
or UO_1038 (O_1038,N_18065,N_18969);
or UO_1039 (O_1039,N_18589,N_19134);
xor UO_1040 (O_1040,N_18827,N_19129);
and UO_1041 (O_1041,N_19496,N_19624);
or UO_1042 (O_1042,N_18885,N_18612);
nand UO_1043 (O_1043,N_19025,N_19612);
nand UO_1044 (O_1044,N_18764,N_18351);
nor UO_1045 (O_1045,N_18576,N_19371);
nand UO_1046 (O_1046,N_18489,N_18409);
or UO_1047 (O_1047,N_18190,N_19835);
nand UO_1048 (O_1048,N_18156,N_18193);
xnor UO_1049 (O_1049,N_19380,N_18530);
or UO_1050 (O_1050,N_18915,N_19128);
xnor UO_1051 (O_1051,N_19882,N_18527);
and UO_1052 (O_1052,N_19769,N_19861);
or UO_1053 (O_1053,N_19913,N_19505);
or UO_1054 (O_1054,N_19073,N_18260);
and UO_1055 (O_1055,N_18292,N_19448);
nand UO_1056 (O_1056,N_19286,N_19720);
and UO_1057 (O_1057,N_19696,N_19058);
and UO_1058 (O_1058,N_19648,N_19045);
nor UO_1059 (O_1059,N_18521,N_19110);
and UO_1060 (O_1060,N_18655,N_19774);
nor UO_1061 (O_1061,N_19107,N_19809);
or UO_1062 (O_1062,N_18011,N_18144);
nor UO_1063 (O_1063,N_19614,N_19172);
nor UO_1064 (O_1064,N_18643,N_19555);
and UO_1065 (O_1065,N_19702,N_19399);
or UO_1066 (O_1066,N_19617,N_18279);
or UO_1067 (O_1067,N_18401,N_19046);
or UO_1068 (O_1068,N_19581,N_18620);
nor UO_1069 (O_1069,N_18816,N_19940);
nand UO_1070 (O_1070,N_19250,N_19070);
and UO_1071 (O_1071,N_18312,N_18355);
xnor UO_1072 (O_1072,N_19170,N_19596);
and UO_1073 (O_1073,N_19080,N_19154);
and UO_1074 (O_1074,N_19733,N_18418);
nor UO_1075 (O_1075,N_18755,N_19797);
nor UO_1076 (O_1076,N_19287,N_18088);
nand UO_1077 (O_1077,N_19825,N_19615);
or UO_1078 (O_1078,N_18174,N_19369);
or UO_1079 (O_1079,N_19150,N_18244);
and UO_1080 (O_1080,N_19488,N_19768);
and UO_1081 (O_1081,N_19156,N_19666);
and UO_1082 (O_1082,N_18032,N_19363);
and UO_1083 (O_1083,N_18405,N_19210);
and UO_1084 (O_1084,N_18606,N_19735);
nand UO_1085 (O_1085,N_18323,N_18980);
nor UO_1086 (O_1086,N_18105,N_19348);
and UO_1087 (O_1087,N_18227,N_18577);
or UO_1088 (O_1088,N_19121,N_18599);
or UO_1089 (O_1089,N_18906,N_19029);
or UO_1090 (O_1090,N_18970,N_18579);
xnor UO_1091 (O_1091,N_18385,N_18209);
nand UO_1092 (O_1092,N_19403,N_19055);
and UO_1093 (O_1093,N_19911,N_18775);
xor UO_1094 (O_1094,N_18985,N_18203);
nor UO_1095 (O_1095,N_19586,N_18098);
nand UO_1096 (O_1096,N_19177,N_19197);
and UO_1097 (O_1097,N_18850,N_18760);
and UO_1098 (O_1098,N_19366,N_18512);
and UO_1099 (O_1099,N_19530,N_19550);
and UO_1100 (O_1100,N_18475,N_19749);
and UO_1101 (O_1101,N_19162,N_18343);
xnor UO_1102 (O_1102,N_19747,N_19676);
and UO_1103 (O_1103,N_19535,N_18358);
nand UO_1104 (O_1104,N_19970,N_18903);
and UO_1105 (O_1105,N_18787,N_18636);
and UO_1106 (O_1106,N_19098,N_18740);
or UO_1107 (O_1107,N_18511,N_19058);
nand UO_1108 (O_1108,N_19001,N_19539);
xor UO_1109 (O_1109,N_18711,N_18693);
nand UO_1110 (O_1110,N_19478,N_19927);
nand UO_1111 (O_1111,N_18920,N_18816);
or UO_1112 (O_1112,N_19414,N_19295);
nor UO_1113 (O_1113,N_19240,N_19248);
nor UO_1114 (O_1114,N_18933,N_19417);
nand UO_1115 (O_1115,N_19848,N_19100);
and UO_1116 (O_1116,N_18477,N_19894);
nand UO_1117 (O_1117,N_18589,N_19818);
nand UO_1118 (O_1118,N_18184,N_19054);
nor UO_1119 (O_1119,N_18345,N_18192);
xor UO_1120 (O_1120,N_19636,N_18818);
nor UO_1121 (O_1121,N_18497,N_18781);
and UO_1122 (O_1122,N_18159,N_18463);
xor UO_1123 (O_1123,N_18309,N_18864);
xnor UO_1124 (O_1124,N_18288,N_18511);
or UO_1125 (O_1125,N_19538,N_19866);
nor UO_1126 (O_1126,N_18791,N_19609);
and UO_1127 (O_1127,N_19339,N_19398);
nor UO_1128 (O_1128,N_18253,N_18026);
nand UO_1129 (O_1129,N_19680,N_19795);
nand UO_1130 (O_1130,N_18996,N_19126);
xor UO_1131 (O_1131,N_18168,N_19245);
nor UO_1132 (O_1132,N_18245,N_18804);
or UO_1133 (O_1133,N_18210,N_18585);
nand UO_1134 (O_1134,N_19039,N_19350);
nand UO_1135 (O_1135,N_18620,N_18343);
nor UO_1136 (O_1136,N_19621,N_19194);
nor UO_1137 (O_1137,N_19052,N_19645);
nor UO_1138 (O_1138,N_18626,N_19684);
and UO_1139 (O_1139,N_19690,N_18073);
or UO_1140 (O_1140,N_18639,N_18463);
and UO_1141 (O_1141,N_19488,N_18428);
and UO_1142 (O_1142,N_18159,N_19422);
and UO_1143 (O_1143,N_19521,N_18438);
and UO_1144 (O_1144,N_18530,N_19193);
nor UO_1145 (O_1145,N_18919,N_18845);
or UO_1146 (O_1146,N_18348,N_18788);
nor UO_1147 (O_1147,N_19977,N_18918);
nand UO_1148 (O_1148,N_18414,N_19015);
nor UO_1149 (O_1149,N_18301,N_18321);
and UO_1150 (O_1150,N_18391,N_19536);
and UO_1151 (O_1151,N_18073,N_18959);
or UO_1152 (O_1152,N_18338,N_18432);
and UO_1153 (O_1153,N_19337,N_19472);
or UO_1154 (O_1154,N_18600,N_19203);
or UO_1155 (O_1155,N_19988,N_19255);
or UO_1156 (O_1156,N_19198,N_18267);
nand UO_1157 (O_1157,N_18190,N_18059);
or UO_1158 (O_1158,N_18220,N_18586);
nand UO_1159 (O_1159,N_18158,N_18525);
and UO_1160 (O_1160,N_19330,N_18264);
xor UO_1161 (O_1161,N_18159,N_19002);
and UO_1162 (O_1162,N_19742,N_18651);
and UO_1163 (O_1163,N_18543,N_19577);
or UO_1164 (O_1164,N_19544,N_19883);
and UO_1165 (O_1165,N_19068,N_19794);
nand UO_1166 (O_1166,N_18203,N_18379);
nor UO_1167 (O_1167,N_18529,N_18860);
nand UO_1168 (O_1168,N_19683,N_18218);
nand UO_1169 (O_1169,N_18676,N_18760);
xor UO_1170 (O_1170,N_19696,N_19085);
and UO_1171 (O_1171,N_18614,N_19549);
or UO_1172 (O_1172,N_19118,N_19444);
xnor UO_1173 (O_1173,N_19578,N_18250);
and UO_1174 (O_1174,N_19284,N_18586);
and UO_1175 (O_1175,N_18410,N_19820);
and UO_1176 (O_1176,N_18856,N_19759);
xor UO_1177 (O_1177,N_19739,N_19389);
and UO_1178 (O_1178,N_18813,N_18817);
nand UO_1179 (O_1179,N_19532,N_19733);
and UO_1180 (O_1180,N_18189,N_18836);
nand UO_1181 (O_1181,N_19299,N_18756);
nor UO_1182 (O_1182,N_19205,N_19120);
and UO_1183 (O_1183,N_18419,N_19907);
nand UO_1184 (O_1184,N_18518,N_19380);
and UO_1185 (O_1185,N_19638,N_18983);
xor UO_1186 (O_1186,N_19598,N_18472);
nor UO_1187 (O_1187,N_18630,N_18171);
and UO_1188 (O_1188,N_18565,N_18443);
nand UO_1189 (O_1189,N_18989,N_18100);
xnor UO_1190 (O_1190,N_18463,N_19351);
nand UO_1191 (O_1191,N_18276,N_18527);
xor UO_1192 (O_1192,N_18465,N_19077);
nand UO_1193 (O_1193,N_18545,N_18231);
nor UO_1194 (O_1194,N_19606,N_19096);
nand UO_1195 (O_1195,N_18077,N_18489);
nor UO_1196 (O_1196,N_19444,N_19143);
xnor UO_1197 (O_1197,N_19834,N_19269);
nor UO_1198 (O_1198,N_18062,N_19398);
nand UO_1199 (O_1199,N_18171,N_19814);
and UO_1200 (O_1200,N_18071,N_19366);
xor UO_1201 (O_1201,N_18893,N_18731);
nor UO_1202 (O_1202,N_19971,N_19863);
xor UO_1203 (O_1203,N_18339,N_18037);
nor UO_1204 (O_1204,N_19206,N_19911);
nor UO_1205 (O_1205,N_18621,N_18480);
or UO_1206 (O_1206,N_18784,N_18889);
and UO_1207 (O_1207,N_19676,N_18541);
xor UO_1208 (O_1208,N_19753,N_19943);
nand UO_1209 (O_1209,N_19328,N_19317);
and UO_1210 (O_1210,N_18292,N_18437);
and UO_1211 (O_1211,N_19179,N_19507);
or UO_1212 (O_1212,N_19296,N_18475);
nor UO_1213 (O_1213,N_19085,N_18632);
xor UO_1214 (O_1214,N_19271,N_19926);
nand UO_1215 (O_1215,N_18471,N_18072);
nor UO_1216 (O_1216,N_18913,N_18984);
nor UO_1217 (O_1217,N_19548,N_19488);
and UO_1218 (O_1218,N_19750,N_19776);
nand UO_1219 (O_1219,N_19860,N_19706);
and UO_1220 (O_1220,N_18095,N_19826);
nand UO_1221 (O_1221,N_19214,N_19737);
nand UO_1222 (O_1222,N_19146,N_18828);
nand UO_1223 (O_1223,N_19661,N_19945);
and UO_1224 (O_1224,N_18272,N_19585);
nand UO_1225 (O_1225,N_19365,N_19097);
nor UO_1226 (O_1226,N_19608,N_19609);
or UO_1227 (O_1227,N_18068,N_18506);
and UO_1228 (O_1228,N_18872,N_18469);
xor UO_1229 (O_1229,N_19637,N_18036);
or UO_1230 (O_1230,N_18630,N_18662);
nand UO_1231 (O_1231,N_18734,N_18839);
and UO_1232 (O_1232,N_19164,N_19607);
or UO_1233 (O_1233,N_19336,N_19401);
nand UO_1234 (O_1234,N_19687,N_18445);
xor UO_1235 (O_1235,N_19571,N_18274);
nor UO_1236 (O_1236,N_19512,N_19160);
and UO_1237 (O_1237,N_18248,N_18454);
and UO_1238 (O_1238,N_19077,N_18080);
or UO_1239 (O_1239,N_19110,N_18796);
nor UO_1240 (O_1240,N_19591,N_18772);
and UO_1241 (O_1241,N_19198,N_19795);
nand UO_1242 (O_1242,N_19161,N_19130);
nand UO_1243 (O_1243,N_18289,N_18162);
nor UO_1244 (O_1244,N_19152,N_19838);
nor UO_1245 (O_1245,N_19846,N_18447);
nor UO_1246 (O_1246,N_18833,N_18158);
and UO_1247 (O_1247,N_19287,N_19106);
nor UO_1248 (O_1248,N_18899,N_19494);
or UO_1249 (O_1249,N_18379,N_18283);
and UO_1250 (O_1250,N_18838,N_19973);
or UO_1251 (O_1251,N_18078,N_18777);
and UO_1252 (O_1252,N_19470,N_19012);
nor UO_1253 (O_1253,N_18413,N_19622);
and UO_1254 (O_1254,N_19471,N_19805);
or UO_1255 (O_1255,N_19374,N_19055);
nand UO_1256 (O_1256,N_18022,N_19573);
or UO_1257 (O_1257,N_18603,N_18030);
nor UO_1258 (O_1258,N_18964,N_19300);
nand UO_1259 (O_1259,N_18388,N_18844);
and UO_1260 (O_1260,N_19969,N_19950);
and UO_1261 (O_1261,N_18253,N_19699);
and UO_1262 (O_1262,N_18752,N_18719);
or UO_1263 (O_1263,N_18984,N_19651);
nor UO_1264 (O_1264,N_19956,N_18998);
nand UO_1265 (O_1265,N_19885,N_18630);
xnor UO_1266 (O_1266,N_18434,N_18157);
or UO_1267 (O_1267,N_19723,N_18723);
and UO_1268 (O_1268,N_19433,N_18607);
nor UO_1269 (O_1269,N_19838,N_19762);
or UO_1270 (O_1270,N_19046,N_18690);
or UO_1271 (O_1271,N_19291,N_19370);
and UO_1272 (O_1272,N_19560,N_18169);
or UO_1273 (O_1273,N_18817,N_18087);
nor UO_1274 (O_1274,N_19745,N_18386);
nor UO_1275 (O_1275,N_18229,N_19974);
or UO_1276 (O_1276,N_18117,N_18145);
or UO_1277 (O_1277,N_18798,N_19593);
nor UO_1278 (O_1278,N_18645,N_18802);
nand UO_1279 (O_1279,N_18800,N_19428);
and UO_1280 (O_1280,N_19245,N_19148);
nand UO_1281 (O_1281,N_18730,N_18806);
and UO_1282 (O_1282,N_19940,N_19001);
xor UO_1283 (O_1283,N_19817,N_18134);
and UO_1284 (O_1284,N_18025,N_18528);
or UO_1285 (O_1285,N_18267,N_19231);
nand UO_1286 (O_1286,N_18799,N_18424);
nor UO_1287 (O_1287,N_18900,N_18341);
nor UO_1288 (O_1288,N_18822,N_19782);
xnor UO_1289 (O_1289,N_18317,N_18527);
and UO_1290 (O_1290,N_18981,N_19441);
nand UO_1291 (O_1291,N_18572,N_18947);
nand UO_1292 (O_1292,N_19072,N_19280);
xor UO_1293 (O_1293,N_19896,N_18761);
nor UO_1294 (O_1294,N_18242,N_18979);
and UO_1295 (O_1295,N_18613,N_19989);
and UO_1296 (O_1296,N_19526,N_18207);
xnor UO_1297 (O_1297,N_19201,N_19241);
nor UO_1298 (O_1298,N_19067,N_18761);
and UO_1299 (O_1299,N_18643,N_18977);
or UO_1300 (O_1300,N_18836,N_19314);
and UO_1301 (O_1301,N_19000,N_18560);
nor UO_1302 (O_1302,N_19468,N_18983);
and UO_1303 (O_1303,N_18122,N_18044);
nor UO_1304 (O_1304,N_18339,N_18025);
nand UO_1305 (O_1305,N_18451,N_18580);
and UO_1306 (O_1306,N_19692,N_19392);
or UO_1307 (O_1307,N_19770,N_19164);
xor UO_1308 (O_1308,N_18145,N_18458);
nand UO_1309 (O_1309,N_19759,N_18610);
or UO_1310 (O_1310,N_19114,N_18054);
and UO_1311 (O_1311,N_19449,N_18587);
nor UO_1312 (O_1312,N_18160,N_19845);
xnor UO_1313 (O_1313,N_18347,N_19894);
nand UO_1314 (O_1314,N_19615,N_19278);
or UO_1315 (O_1315,N_19953,N_18183);
nand UO_1316 (O_1316,N_18483,N_19347);
and UO_1317 (O_1317,N_19513,N_19213);
and UO_1318 (O_1318,N_18552,N_19285);
or UO_1319 (O_1319,N_19605,N_19320);
and UO_1320 (O_1320,N_19791,N_19377);
nand UO_1321 (O_1321,N_19008,N_18416);
nand UO_1322 (O_1322,N_18203,N_19036);
and UO_1323 (O_1323,N_19717,N_18454);
nand UO_1324 (O_1324,N_19393,N_18937);
or UO_1325 (O_1325,N_18135,N_19838);
nor UO_1326 (O_1326,N_18548,N_19782);
or UO_1327 (O_1327,N_19892,N_19862);
and UO_1328 (O_1328,N_18798,N_18254);
xor UO_1329 (O_1329,N_18107,N_18741);
and UO_1330 (O_1330,N_18266,N_19422);
and UO_1331 (O_1331,N_19496,N_19333);
nand UO_1332 (O_1332,N_19952,N_18903);
or UO_1333 (O_1333,N_19217,N_19621);
and UO_1334 (O_1334,N_19814,N_18589);
xor UO_1335 (O_1335,N_18599,N_19082);
nor UO_1336 (O_1336,N_18240,N_18318);
nand UO_1337 (O_1337,N_19819,N_18097);
and UO_1338 (O_1338,N_19001,N_18532);
and UO_1339 (O_1339,N_19697,N_19838);
and UO_1340 (O_1340,N_18156,N_19564);
nand UO_1341 (O_1341,N_18650,N_19507);
or UO_1342 (O_1342,N_18340,N_18310);
nor UO_1343 (O_1343,N_18526,N_18657);
nand UO_1344 (O_1344,N_18524,N_19309);
nor UO_1345 (O_1345,N_19877,N_18385);
or UO_1346 (O_1346,N_19434,N_19574);
or UO_1347 (O_1347,N_19850,N_19130);
or UO_1348 (O_1348,N_19233,N_18807);
and UO_1349 (O_1349,N_19276,N_19125);
nand UO_1350 (O_1350,N_19229,N_19448);
nand UO_1351 (O_1351,N_18404,N_18896);
nand UO_1352 (O_1352,N_18018,N_19442);
nand UO_1353 (O_1353,N_18818,N_19488);
nor UO_1354 (O_1354,N_18032,N_19852);
and UO_1355 (O_1355,N_18017,N_18364);
or UO_1356 (O_1356,N_18337,N_19757);
and UO_1357 (O_1357,N_19483,N_19995);
or UO_1358 (O_1358,N_18014,N_19064);
xnor UO_1359 (O_1359,N_18925,N_19497);
nand UO_1360 (O_1360,N_18286,N_18452);
nand UO_1361 (O_1361,N_19102,N_19560);
or UO_1362 (O_1362,N_18775,N_18392);
nand UO_1363 (O_1363,N_19472,N_18397);
nor UO_1364 (O_1364,N_18548,N_19519);
xor UO_1365 (O_1365,N_18789,N_18424);
and UO_1366 (O_1366,N_19023,N_18041);
or UO_1367 (O_1367,N_18798,N_18761);
or UO_1368 (O_1368,N_18285,N_18200);
and UO_1369 (O_1369,N_19929,N_19726);
nand UO_1370 (O_1370,N_19729,N_19826);
or UO_1371 (O_1371,N_18235,N_18413);
nand UO_1372 (O_1372,N_18165,N_18454);
and UO_1373 (O_1373,N_19126,N_19584);
or UO_1374 (O_1374,N_18506,N_18818);
xor UO_1375 (O_1375,N_18094,N_18212);
nand UO_1376 (O_1376,N_18251,N_18681);
xnor UO_1377 (O_1377,N_19085,N_19808);
nor UO_1378 (O_1378,N_19775,N_19396);
nand UO_1379 (O_1379,N_18086,N_19383);
nand UO_1380 (O_1380,N_19679,N_19590);
xor UO_1381 (O_1381,N_19298,N_18179);
xnor UO_1382 (O_1382,N_19872,N_18992);
nor UO_1383 (O_1383,N_18587,N_19963);
or UO_1384 (O_1384,N_18525,N_18939);
xnor UO_1385 (O_1385,N_19794,N_19502);
nand UO_1386 (O_1386,N_18411,N_19531);
xnor UO_1387 (O_1387,N_18035,N_18761);
nor UO_1388 (O_1388,N_18037,N_18602);
nor UO_1389 (O_1389,N_18748,N_19257);
nor UO_1390 (O_1390,N_18091,N_18505);
or UO_1391 (O_1391,N_19493,N_18196);
or UO_1392 (O_1392,N_18239,N_19975);
nand UO_1393 (O_1393,N_19196,N_18668);
nand UO_1394 (O_1394,N_19060,N_18436);
xnor UO_1395 (O_1395,N_18566,N_19694);
and UO_1396 (O_1396,N_19133,N_19964);
and UO_1397 (O_1397,N_19755,N_18904);
and UO_1398 (O_1398,N_18307,N_19665);
or UO_1399 (O_1399,N_18837,N_19802);
nor UO_1400 (O_1400,N_18729,N_18018);
nand UO_1401 (O_1401,N_19857,N_18534);
or UO_1402 (O_1402,N_18138,N_19860);
nor UO_1403 (O_1403,N_18192,N_18940);
or UO_1404 (O_1404,N_19174,N_19848);
nor UO_1405 (O_1405,N_18876,N_18381);
and UO_1406 (O_1406,N_19489,N_19045);
nor UO_1407 (O_1407,N_18467,N_19022);
and UO_1408 (O_1408,N_19107,N_19313);
or UO_1409 (O_1409,N_18917,N_19020);
nor UO_1410 (O_1410,N_18973,N_18056);
nor UO_1411 (O_1411,N_19466,N_18212);
or UO_1412 (O_1412,N_19030,N_19311);
or UO_1413 (O_1413,N_18873,N_18447);
or UO_1414 (O_1414,N_18072,N_19525);
xnor UO_1415 (O_1415,N_19708,N_19212);
or UO_1416 (O_1416,N_18164,N_18442);
nand UO_1417 (O_1417,N_19552,N_18217);
nand UO_1418 (O_1418,N_19634,N_18484);
or UO_1419 (O_1419,N_18701,N_18372);
nor UO_1420 (O_1420,N_18822,N_19616);
or UO_1421 (O_1421,N_19864,N_18540);
nand UO_1422 (O_1422,N_19911,N_19135);
or UO_1423 (O_1423,N_19119,N_19195);
xnor UO_1424 (O_1424,N_19660,N_19294);
nand UO_1425 (O_1425,N_18942,N_19198);
nand UO_1426 (O_1426,N_19335,N_19539);
or UO_1427 (O_1427,N_19266,N_18484);
and UO_1428 (O_1428,N_18240,N_18699);
nor UO_1429 (O_1429,N_18120,N_19914);
or UO_1430 (O_1430,N_18929,N_18196);
and UO_1431 (O_1431,N_18579,N_18515);
or UO_1432 (O_1432,N_18156,N_18090);
and UO_1433 (O_1433,N_18085,N_18501);
nand UO_1434 (O_1434,N_19720,N_19565);
nand UO_1435 (O_1435,N_18911,N_18975);
nor UO_1436 (O_1436,N_18926,N_18876);
or UO_1437 (O_1437,N_18528,N_19057);
and UO_1438 (O_1438,N_19428,N_19280);
nand UO_1439 (O_1439,N_18991,N_18779);
or UO_1440 (O_1440,N_19920,N_19482);
and UO_1441 (O_1441,N_19581,N_19960);
and UO_1442 (O_1442,N_19462,N_19267);
nor UO_1443 (O_1443,N_19154,N_18626);
nor UO_1444 (O_1444,N_19383,N_19740);
nor UO_1445 (O_1445,N_18502,N_18057);
nor UO_1446 (O_1446,N_19953,N_19218);
nor UO_1447 (O_1447,N_19965,N_18807);
and UO_1448 (O_1448,N_19982,N_19151);
nor UO_1449 (O_1449,N_19041,N_18626);
nor UO_1450 (O_1450,N_19427,N_18196);
nand UO_1451 (O_1451,N_19874,N_19530);
nor UO_1452 (O_1452,N_18810,N_18486);
nor UO_1453 (O_1453,N_18244,N_19770);
or UO_1454 (O_1454,N_18396,N_19417);
or UO_1455 (O_1455,N_18146,N_19989);
and UO_1456 (O_1456,N_19796,N_18156);
nor UO_1457 (O_1457,N_18037,N_18740);
nor UO_1458 (O_1458,N_18660,N_19159);
xnor UO_1459 (O_1459,N_19889,N_18582);
nand UO_1460 (O_1460,N_18203,N_19063);
or UO_1461 (O_1461,N_18098,N_18853);
and UO_1462 (O_1462,N_18420,N_18709);
nand UO_1463 (O_1463,N_18428,N_18974);
nor UO_1464 (O_1464,N_19063,N_18941);
xnor UO_1465 (O_1465,N_18689,N_19413);
nand UO_1466 (O_1466,N_18824,N_18042);
nor UO_1467 (O_1467,N_19971,N_18860);
nand UO_1468 (O_1468,N_19464,N_18093);
nand UO_1469 (O_1469,N_19387,N_18142);
nand UO_1470 (O_1470,N_18272,N_19148);
nor UO_1471 (O_1471,N_18955,N_19637);
nor UO_1472 (O_1472,N_18175,N_18832);
and UO_1473 (O_1473,N_19915,N_19428);
nand UO_1474 (O_1474,N_18075,N_19117);
nor UO_1475 (O_1475,N_18211,N_19023);
and UO_1476 (O_1476,N_18901,N_18532);
or UO_1477 (O_1477,N_19971,N_19093);
xor UO_1478 (O_1478,N_18325,N_19702);
xnor UO_1479 (O_1479,N_18848,N_19126);
and UO_1480 (O_1480,N_19505,N_19701);
and UO_1481 (O_1481,N_18264,N_18393);
xnor UO_1482 (O_1482,N_18216,N_18452);
nor UO_1483 (O_1483,N_19887,N_18517);
or UO_1484 (O_1484,N_18340,N_18306);
nand UO_1485 (O_1485,N_19036,N_19996);
or UO_1486 (O_1486,N_19874,N_18130);
nand UO_1487 (O_1487,N_18164,N_19565);
or UO_1488 (O_1488,N_19775,N_19642);
nor UO_1489 (O_1489,N_19443,N_19523);
and UO_1490 (O_1490,N_19341,N_19481);
or UO_1491 (O_1491,N_18738,N_19558);
xnor UO_1492 (O_1492,N_19556,N_19236);
and UO_1493 (O_1493,N_18642,N_18602);
nand UO_1494 (O_1494,N_19947,N_19684);
or UO_1495 (O_1495,N_18488,N_19318);
and UO_1496 (O_1496,N_19298,N_18869);
or UO_1497 (O_1497,N_18545,N_18102);
xnor UO_1498 (O_1498,N_19802,N_18237);
nand UO_1499 (O_1499,N_18450,N_18683);
nand UO_1500 (O_1500,N_18187,N_19098);
and UO_1501 (O_1501,N_18560,N_19919);
nor UO_1502 (O_1502,N_18303,N_19891);
and UO_1503 (O_1503,N_18833,N_18270);
nand UO_1504 (O_1504,N_18420,N_18703);
or UO_1505 (O_1505,N_18022,N_19090);
xnor UO_1506 (O_1506,N_19924,N_19506);
nor UO_1507 (O_1507,N_18345,N_19620);
and UO_1508 (O_1508,N_18435,N_18555);
or UO_1509 (O_1509,N_19929,N_18389);
and UO_1510 (O_1510,N_18900,N_18579);
and UO_1511 (O_1511,N_19465,N_19934);
or UO_1512 (O_1512,N_18198,N_19675);
nand UO_1513 (O_1513,N_19036,N_19027);
and UO_1514 (O_1514,N_18441,N_19892);
or UO_1515 (O_1515,N_18706,N_19520);
and UO_1516 (O_1516,N_18237,N_18590);
xnor UO_1517 (O_1517,N_19051,N_19826);
nor UO_1518 (O_1518,N_18755,N_19594);
nor UO_1519 (O_1519,N_19791,N_19434);
or UO_1520 (O_1520,N_18978,N_19290);
nand UO_1521 (O_1521,N_18267,N_19405);
nor UO_1522 (O_1522,N_19735,N_18752);
or UO_1523 (O_1523,N_19935,N_18735);
xnor UO_1524 (O_1524,N_18841,N_18734);
nor UO_1525 (O_1525,N_18846,N_18832);
nor UO_1526 (O_1526,N_19994,N_18746);
or UO_1527 (O_1527,N_18157,N_19924);
nor UO_1528 (O_1528,N_19866,N_19751);
and UO_1529 (O_1529,N_19182,N_19536);
nor UO_1530 (O_1530,N_19591,N_18560);
nor UO_1531 (O_1531,N_19643,N_18068);
or UO_1532 (O_1532,N_18705,N_19934);
nand UO_1533 (O_1533,N_19410,N_18586);
or UO_1534 (O_1534,N_18844,N_18411);
nor UO_1535 (O_1535,N_18043,N_19742);
or UO_1536 (O_1536,N_19778,N_18464);
or UO_1537 (O_1537,N_19854,N_18703);
xor UO_1538 (O_1538,N_19156,N_19505);
nor UO_1539 (O_1539,N_19556,N_19940);
nand UO_1540 (O_1540,N_19745,N_18395);
or UO_1541 (O_1541,N_19752,N_18570);
nand UO_1542 (O_1542,N_19041,N_19503);
xor UO_1543 (O_1543,N_18113,N_18192);
and UO_1544 (O_1544,N_19697,N_19176);
and UO_1545 (O_1545,N_18165,N_18732);
nand UO_1546 (O_1546,N_18631,N_19420);
nor UO_1547 (O_1547,N_19264,N_19996);
nor UO_1548 (O_1548,N_19309,N_18835);
or UO_1549 (O_1549,N_19796,N_19146);
nand UO_1550 (O_1550,N_18420,N_18009);
xor UO_1551 (O_1551,N_19268,N_18396);
or UO_1552 (O_1552,N_19249,N_18129);
or UO_1553 (O_1553,N_18824,N_18423);
and UO_1554 (O_1554,N_19816,N_18628);
or UO_1555 (O_1555,N_18627,N_18246);
and UO_1556 (O_1556,N_18315,N_18386);
nor UO_1557 (O_1557,N_19967,N_18731);
or UO_1558 (O_1558,N_19075,N_18060);
nand UO_1559 (O_1559,N_18005,N_19001);
and UO_1560 (O_1560,N_19202,N_19163);
and UO_1561 (O_1561,N_19162,N_19416);
xor UO_1562 (O_1562,N_19543,N_18990);
or UO_1563 (O_1563,N_18511,N_18716);
nor UO_1564 (O_1564,N_18601,N_18815);
and UO_1565 (O_1565,N_18137,N_19127);
and UO_1566 (O_1566,N_18881,N_18010);
and UO_1567 (O_1567,N_18796,N_18730);
nand UO_1568 (O_1568,N_19820,N_18061);
nand UO_1569 (O_1569,N_19889,N_19739);
or UO_1570 (O_1570,N_18077,N_18707);
nor UO_1571 (O_1571,N_19705,N_19280);
or UO_1572 (O_1572,N_19940,N_18829);
nand UO_1573 (O_1573,N_19039,N_18357);
xnor UO_1574 (O_1574,N_18195,N_18456);
nor UO_1575 (O_1575,N_19227,N_19452);
and UO_1576 (O_1576,N_19547,N_19805);
nand UO_1577 (O_1577,N_19981,N_18120);
and UO_1578 (O_1578,N_19308,N_18498);
and UO_1579 (O_1579,N_18801,N_18955);
xor UO_1580 (O_1580,N_18874,N_18384);
nand UO_1581 (O_1581,N_18476,N_18812);
nor UO_1582 (O_1582,N_19806,N_19578);
nor UO_1583 (O_1583,N_18428,N_19801);
nor UO_1584 (O_1584,N_19017,N_19481);
nor UO_1585 (O_1585,N_18044,N_19586);
nand UO_1586 (O_1586,N_18065,N_18551);
and UO_1587 (O_1587,N_19728,N_19587);
and UO_1588 (O_1588,N_19860,N_18474);
nor UO_1589 (O_1589,N_19383,N_19441);
xnor UO_1590 (O_1590,N_18337,N_19559);
and UO_1591 (O_1591,N_18165,N_18498);
nand UO_1592 (O_1592,N_19669,N_18528);
nor UO_1593 (O_1593,N_18836,N_19301);
nand UO_1594 (O_1594,N_19367,N_18477);
nand UO_1595 (O_1595,N_19709,N_19680);
or UO_1596 (O_1596,N_18603,N_19717);
nor UO_1597 (O_1597,N_19524,N_18026);
xnor UO_1598 (O_1598,N_19623,N_19710);
nor UO_1599 (O_1599,N_19935,N_19201);
xnor UO_1600 (O_1600,N_18037,N_18666);
or UO_1601 (O_1601,N_19472,N_19363);
xnor UO_1602 (O_1602,N_18650,N_19757);
nand UO_1603 (O_1603,N_18590,N_19137);
nor UO_1604 (O_1604,N_19533,N_19943);
nor UO_1605 (O_1605,N_18904,N_19469);
or UO_1606 (O_1606,N_18284,N_18918);
or UO_1607 (O_1607,N_19427,N_18493);
xor UO_1608 (O_1608,N_18516,N_19069);
or UO_1609 (O_1609,N_18791,N_19304);
and UO_1610 (O_1610,N_19976,N_19946);
xnor UO_1611 (O_1611,N_19908,N_19251);
nor UO_1612 (O_1612,N_18351,N_18110);
nand UO_1613 (O_1613,N_19175,N_18248);
and UO_1614 (O_1614,N_19157,N_19630);
nor UO_1615 (O_1615,N_19464,N_18120);
nor UO_1616 (O_1616,N_19205,N_19733);
or UO_1617 (O_1617,N_19997,N_18949);
or UO_1618 (O_1618,N_19257,N_19033);
and UO_1619 (O_1619,N_18602,N_19734);
or UO_1620 (O_1620,N_19558,N_19779);
and UO_1621 (O_1621,N_18604,N_18700);
or UO_1622 (O_1622,N_19823,N_19215);
nand UO_1623 (O_1623,N_18394,N_18130);
and UO_1624 (O_1624,N_18290,N_19587);
nand UO_1625 (O_1625,N_19476,N_18774);
or UO_1626 (O_1626,N_18228,N_19395);
or UO_1627 (O_1627,N_18549,N_19359);
nand UO_1628 (O_1628,N_19623,N_19603);
or UO_1629 (O_1629,N_19928,N_19330);
or UO_1630 (O_1630,N_18586,N_19209);
and UO_1631 (O_1631,N_19814,N_18165);
nand UO_1632 (O_1632,N_19348,N_19036);
nor UO_1633 (O_1633,N_19347,N_19691);
nor UO_1634 (O_1634,N_19791,N_18898);
xnor UO_1635 (O_1635,N_19643,N_18097);
or UO_1636 (O_1636,N_19222,N_18534);
nor UO_1637 (O_1637,N_19824,N_19112);
nor UO_1638 (O_1638,N_18887,N_18360);
and UO_1639 (O_1639,N_19184,N_19093);
nand UO_1640 (O_1640,N_19300,N_19670);
and UO_1641 (O_1641,N_18135,N_19776);
nand UO_1642 (O_1642,N_18658,N_18802);
or UO_1643 (O_1643,N_18151,N_18410);
nand UO_1644 (O_1644,N_19359,N_18173);
or UO_1645 (O_1645,N_19314,N_19664);
and UO_1646 (O_1646,N_19931,N_18437);
nand UO_1647 (O_1647,N_18308,N_19246);
and UO_1648 (O_1648,N_19540,N_18581);
nand UO_1649 (O_1649,N_19587,N_19763);
nand UO_1650 (O_1650,N_18755,N_19582);
nor UO_1651 (O_1651,N_19840,N_18806);
xor UO_1652 (O_1652,N_18487,N_19646);
or UO_1653 (O_1653,N_19472,N_19424);
nand UO_1654 (O_1654,N_19347,N_19768);
and UO_1655 (O_1655,N_19501,N_19018);
nor UO_1656 (O_1656,N_19988,N_19752);
or UO_1657 (O_1657,N_19618,N_19468);
nand UO_1658 (O_1658,N_19338,N_18600);
nor UO_1659 (O_1659,N_18142,N_18685);
or UO_1660 (O_1660,N_19742,N_18126);
or UO_1661 (O_1661,N_19721,N_18129);
nor UO_1662 (O_1662,N_18477,N_19746);
or UO_1663 (O_1663,N_18965,N_19540);
or UO_1664 (O_1664,N_18561,N_18928);
xnor UO_1665 (O_1665,N_19570,N_18080);
xor UO_1666 (O_1666,N_19951,N_19894);
nand UO_1667 (O_1667,N_18825,N_19287);
and UO_1668 (O_1668,N_18396,N_19657);
nor UO_1669 (O_1669,N_19410,N_19367);
xor UO_1670 (O_1670,N_18283,N_19530);
or UO_1671 (O_1671,N_18323,N_19266);
nor UO_1672 (O_1672,N_18106,N_19483);
and UO_1673 (O_1673,N_19937,N_19460);
and UO_1674 (O_1674,N_19846,N_18231);
nand UO_1675 (O_1675,N_18075,N_18069);
or UO_1676 (O_1676,N_19038,N_18634);
nor UO_1677 (O_1677,N_18925,N_18589);
nor UO_1678 (O_1678,N_18094,N_19064);
and UO_1679 (O_1679,N_18249,N_19866);
nand UO_1680 (O_1680,N_19188,N_18862);
xnor UO_1681 (O_1681,N_19249,N_19158);
or UO_1682 (O_1682,N_19019,N_18277);
nand UO_1683 (O_1683,N_19427,N_18672);
and UO_1684 (O_1684,N_18444,N_18260);
xnor UO_1685 (O_1685,N_18936,N_18415);
and UO_1686 (O_1686,N_19832,N_18347);
nand UO_1687 (O_1687,N_18297,N_19670);
xor UO_1688 (O_1688,N_18329,N_18986);
and UO_1689 (O_1689,N_18564,N_18413);
and UO_1690 (O_1690,N_18371,N_19716);
and UO_1691 (O_1691,N_18624,N_19749);
nor UO_1692 (O_1692,N_19149,N_19659);
nand UO_1693 (O_1693,N_18980,N_19203);
and UO_1694 (O_1694,N_19532,N_19860);
or UO_1695 (O_1695,N_18023,N_19066);
nand UO_1696 (O_1696,N_19278,N_19325);
and UO_1697 (O_1697,N_18737,N_18481);
and UO_1698 (O_1698,N_19893,N_19930);
nor UO_1699 (O_1699,N_18492,N_18851);
and UO_1700 (O_1700,N_19785,N_19443);
or UO_1701 (O_1701,N_19640,N_18073);
xnor UO_1702 (O_1702,N_19933,N_19182);
or UO_1703 (O_1703,N_19469,N_19607);
nand UO_1704 (O_1704,N_18501,N_19714);
xor UO_1705 (O_1705,N_18845,N_18523);
nand UO_1706 (O_1706,N_18401,N_19687);
nor UO_1707 (O_1707,N_19683,N_19730);
nand UO_1708 (O_1708,N_19345,N_19869);
or UO_1709 (O_1709,N_18118,N_19126);
or UO_1710 (O_1710,N_18864,N_19958);
xnor UO_1711 (O_1711,N_18681,N_18983);
and UO_1712 (O_1712,N_18550,N_19408);
nor UO_1713 (O_1713,N_19778,N_19478);
nor UO_1714 (O_1714,N_19897,N_19426);
nand UO_1715 (O_1715,N_19955,N_19143);
and UO_1716 (O_1716,N_18992,N_19972);
nand UO_1717 (O_1717,N_18434,N_19564);
nor UO_1718 (O_1718,N_19600,N_18132);
xor UO_1719 (O_1719,N_19355,N_18904);
nand UO_1720 (O_1720,N_19382,N_19259);
nor UO_1721 (O_1721,N_18215,N_18289);
or UO_1722 (O_1722,N_19836,N_18459);
and UO_1723 (O_1723,N_18350,N_18487);
and UO_1724 (O_1724,N_19103,N_18545);
and UO_1725 (O_1725,N_19662,N_19764);
and UO_1726 (O_1726,N_19815,N_18332);
nor UO_1727 (O_1727,N_18929,N_19100);
nand UO_1728 (O_1728,N_19186,N_19026);
nor UO_1729 (O_1729,N_18373,N_19551);
or UO_1730 (O_1730,N_18331,N_18122);
nand UO_1731 (O_1731,N_18732,N_19160);
xor UO_1732 (O_1732,N_19146,N_19026);
and UO_1733 (O_1733,N_18302,N_19719);
or UO_1734 (O_1734,N_18044,N_18861);
nand UO_1735 (O_1735,N_19902,N_19897);
or UO_1736 (O_1736,N_18794,N_18025);
nand UO_1737 (O_1737,N_19123,N_18822);
or UO_1738 (O_1738,N_18581,N_19173);
nor UO_1739 (O_1739,N_19380,N_18243);
and UO_1740 (O_1740,N_19640,N_19953);
and UO_1741 (O_1741,N_18037,N_19362);
and UO_1742 (O_1742,N_18076,N_19654);
nor UO_1743 (O_1743,N_18119,N_18178);
and UO_1744 (O_1744,N_19545,N_18561);
nor UO_1745 (O_1745,N_18490,N_18934);
nand UO_1746 (O_1746,N_18853,N_19388);
or UO_1747 (O_1747,N_19994,N_19449);
or UO_1748 (O_1748,N_18667,N_18876);
or UO_1749 (O_1749,N_18257,N_19086);
nor UO_1750 (O_1750,N_19568,N_18420);
nand UO_1751 (O_1751,N_18161,N_18568);
or UO_1752 (O_1752,N_18269,N_19212);
nor UO_1753 (O_1753,N_18822,N_18137);
or UO_1754 (O_1754,N_19465,N_18376);
nand UO_1755 (O_1755,N_19259,N_19161);
and UO_1756 (O_1756,N_19665,N_18292);
or UO_1757 (O_1757,N_19926,N_18763);
and UO_1758 (O_1758,N_19983,N_19239);
or UO_1759 (O_1759,N_19295,N_19588);
xnor UO_1760 (O_1760,N_19954,N_19831);
xnor UO_1761 (O_1761,N_19659,N_19255);
or UO_1762 (O_1762,N_19421,N_18081);
nor UO_1763 (O_1763,N_18682,N_18982);
nor UO_1764 (O_1764,N_19906,N_19689);
nand UO_1765 (O_1765,N_19065,N_19484);
nor UO_1766 (O_1766,N_18087,N_19633);
and UO_1767 (O_1767,N_19549,N_18632);
or UO_1768 (O_1768,N_18619,N_18520);
and UO_1769 (O_1769,N_19824,N_19829);
nor UO_1770 (O_1770,N_18554,N_19133);
nand UO_1771 (O_1771,N_19883,N_19494);
and UO_1772 (O_1772,N_18199,N_18544);
and UO_1773 (O_1773,N_19867,N_19323);
or UO_1774 (O_1774,N_19058,N_18292);
nor UO_1775 (O_1775,N_18179,N_19425);
and UO_1776 (O_1776,N_19283,N_18025);
xor UO_1777 (O_1777,N_18153,N_18462);
nand UO_1778 (O_1778,N_19032,N_19155);
nor UO_1779 (O_1779,N_19158,N_19593);
nand UO_1780 (O_1780,N_18290,N_19209);
or UO_1781 (O_1781,N_19654,N_19671);
and UO_1782 (O_1782,N_18364,N_19111);
and UO_1783 (O_1783,N_18008,N_18789);
nand UO_1784 (O_1784,N_18504,N_18542);
xor UO_1785 (O_1785,N_19367,N_18446);
or UO_1786 (O_1786,N_19982,N_19484);
or UO_1787 (O_1787,N_19012,N_19775);
nand UO_1788 (O_1788,N_18046,N_18290);
xor UO_1789 (O_1789,N_19565,N_18841);
and UO_1790 (O_1790,N_18430,N_19367);
and UO_1791 (O_1791,N_19899,N_18353);
nand UO_1792 (O_1792,N_18296,N_18094);
nand UO_1793 (O_1793,N_19682,N_19709);
or UO_1794 (O_1794,N_19731,N_18864);
nor UO_1795 (O_1795,N_19144,N_18539);
or UO_1796 (O_1796,N_18109,N_18737);
and UO_1797 (O_1797,N_19611,N_19847);
nand UO_1798 (O_1798,N_18017,N_18872);
nand UO_1799 (O_1799,N_18524,N_19893);
or UO_1800 (O_1800,N_18347,N_18323);
and UO_1801 (O_1801,N_19451,N_19975);
or UO_1802 (O_1802,N_19182,N_19787);
nand UO_1803 (O_1803,N_19081,N_19356);
nand UO_1804 (O_1804,N_19263,N_18980);
nor UO_1805 (O_1805,N_18359,N_19292);
or UO_1806 (O_1806,N_18378,N_18907);
and UO_1807 (O_1807,N_18446,N_18663);
nor UO_1808 (O_1808,N_18090,N_19568);
nor UO_1809 (O_1809,N_18602,N_19170);
or UO_1810 (O_1810,N_19509,N_18558);
nand UO_1811 (O_1811,N_19686,N_19849);
or UO_1812 (O_1812,N_18194,N_19185);
or UO_1813 (O_1813,N_18935,N_19233);
nand UO_1814 (O_1814,N_18627,N_19682);
nor UO_1815 (O_1815,N_18701,N_19863);
nand UO_1816 (O_1816,N_19460,N_19279);
xnor UO_1817 (O_1817,N_19065,N_18582);
nor UO_1818 (O_1818,N_19827,N_18115);
xnor UO_1819 (O_1819,N_19375,N_18135);
xnor UO_1820 (O_1820,N_18474,N_18045);
nor UO_1821 (O_1821,N_19196,N_18170);
nand UO_1822 (O_1822,N_19810,N_19280);
and UO_1823 (O_1823,N_18788,N_19236);
or UO_1824 (O_1824,N_19987,N_19393);
nor UO_1825 (O_1825,N_19255,N_19176);
or UO_1826 (O_1826,N_19880,N_19071);
nor UO_1827 (O_1827,N_18439,N_18508);
or UO_1828 (O_1828,N_19246,N_19003);
nand UO_1829 (O_1829,N_18294,N_19270);
nand UO_1830 (O_1830,N_19536,N_19007);
or UO_1831 (O_1831,N_18866,N_19408);
xor UO_1832 (O_1832,N_19872,N_18769);
or UO_1833 (O_1833,N_18979,N_19311);
or UO_1834 (O_1834,N_19477,N_19412);
or UO_1835 (O_1835,N_18297,N_19140);
and UO_1836 (O_1836,N_18624,N_19510);
xor UO_1837 (O_1837,N_19819,N_19869);
nor UO_1838 (O_1838,N_18587,N_18692);
nand UO_1839 (O_1839,N_19745,N_19121);
or UO_1840 (O_1840,N_18235,N_18132);
and UO_1841 (O_1841,N_19918,N_18115);
nor UO_1842 (O_1842,N_18586,N_18825);
nand UO_1843 (O_1843,N_19870,N_18795);
and UO_1844 (O_1844,N_18905,N_19395);
xnor UO_1845 (O_1845,N_19371,N_19341);
or UO_1846 (O_1846,N_18326,N_18239);
nand UO_1847 (O_1847,N_19581,N_19229);
and UO_1848 (O_1848,N_18353,N_19627);
nor UO_1849 (O_1849,N_19707,N_18804);
xor UO_1850 (O_1850,N_19642,N_18637);
and UO_1851 (O_1851,N_19411,N_18290);
nor UO_1852 (O_1852,N_18611,N_18883);
and UO_1853 (O_1853,N_18714,N_19689);
nor UO_1854 (O_1854,N_19180,N_19600);
or UO_1855 (O_1855,N_18325,N_18069);
or UO_1856 (O_1856,N_19364,N_19789);
nor UO_1857 (O_1857,N_19089,N_18575);
and UO_1858 (O_1858,N_19076,N_18352);
nand UO_1859 (O_1859,N_19057,N_19770);
and UO_1860 (O_1860,N_18496,N_18923);
or UO_1861 (O_1861,N_18930,N_19034);
or UO_1862 (O_1862,N_18037,N_18401);
nand UO_1863 (O_1863,N_19267,N_18530);
and UO_1864 (O_1864,N_19623,N_19542);
nand UO_1865 (O_1865,N_19550,N_19904);
and UO_1866 (O_1866,N_18229,N_18080);
nor UO_1867 (O_1867,N_18301,N_19565);
or UO_1868 (O_1868,N_18666,N_18912);
and UO_1869 (O_1869,N_18306,N_19326);
nand UO_1870 (O_1870,N_18663,N_18965);
and UO_1871 (O_1871,N_18931,N_19317);
nand UO_1872 (O_1872,N_19278,N_19928);
nor UO_1873 (O_1873,N_18804,N_19719);
xor UO_1874 (O_1874,N_19088,N_19594);
and UO_1875 (O_1875,N_18679,N_18470);
or UO_1876 (O_1876,N_18102,N_18996);
and UO_1877 (O_1877,N_19650,N_19373);
and UO_1878 (O_1878,N_18888,N_19542);
nor UO_1879 (O_1879,N_19855,N_18853);
and UO_1880 (O_1880,N_18945,N_18397);
or UO_1881 (O_1881,N_19286,N_19594);
and UO_1882 (O_1882,N_18610,N_19128);
xnor UO_1883 (O_1883,N_18626,N_18514);
nand UO_1884 (O_1884,N_19314,N_19953);
or UO_1885 (O_1885,N_18854,N_19967);
or UO_1886 (O_1886,N_18581,N_18776);
xnor UO_1887 (O_1887,N_18336,N_19604);
nor UO_1888 (O_1888,N_18726,N_18697);
nand UO_1889 (O_1889,N_18055,N_19637);
and UO_1890 (O_1890,N_19047,N_19224);
or UO_1891 (O_1891,N_19770,N_18259);
or UO_1892 (O_1892,N_18532,N_19438);
or UO_1893 (O_1893,N_18215,N_18468);
nand UO_1894 (O_1894,N_19401,N_19480);
xnor UO_1895 (O_1895,N_18319,N_19828);
or UO_1896 (O_1896,N_18278,N_19070);
nor UO_1897 (O_1897,N_19555,N_19123);
or UO_1898 (O_1898,N_18769,N_18116);
nand UO_1899 (O_1899,N_18281,N_19990);
nand UO_1900 (O_1900,N_19995,N_19629);
xnor UO_1901 (O_1901,N_19924,N_19788);
and UO_1902 (O_1902,N_19804,N_18252);
or UO_1903 (O_1903,N_18556,N_19055);
or UO_1904 (O_1904,N_19233,N_19706);
xor UO_1905 (O_1905,N_19193,N_19941);
or UO_1906 (O_1906,N_19281,N_18589);
and UO_1907 (O_1907,N_18042,N_19853);
nor UO_1908 (O_1908,N_19465,N_19238);
nand UO_1909 (O_1909,N_19809,N_19372);
nor UO_1910 (O_1910,N_18228,N_19951);
nand UO_1911 (O_1911,N_18299,N_19369);
nor UO_1912 (O_1912,N_18280,N_18420);
and UO_1913 (O_1913,N_19575,N_18639);
nor UO_1914 (O_1914,N_19667,N_18638);
and UO_1915 (O_1915,N_18115,N_18488);
and UO_1916 (O_1916,N_19149,N_18992);
and UO_1917 (O_1917,N_18191,N_18896);
nand UO_1918 (O_1918,N_18199,N_19455);
nand UO_1919 (O_1919,N_19989,N_18273);
nor UO_1920 (O_1920,N_19067,N_18445);
or UO_1921 (O_1921,N_18103,N_18510);
or UO_1922 (O_1922,N_19155,N_19180);
nor UO_1923 (O_1923,N_18256,N_19570);
nor UO_1924 (O_1924,N_18265,N_19393);
nand UO_1925 (O_1925,N_19241,N_19771);
nand UO_1926 (O_1926,N_19367,N_18703);
and UO_1927 (O_1927,N_19719,N_18491);
and UO_1928 (O_1928,N_19452,N_18089);
nand UO_1929 (O_1929,N_19776,N_18315);
and UO_1930 (O_1930,N_18992,N_19884);
nand UO_1931 (O_1931,N_18385,N_18616);
or UO_1932 (O_1932,N_19123,N_19887);
xor UO_1933 (O_1933,N_18468,N_18649);
or UO_1934 (O_1934,N_19040,N_18139);
nand UO_1935 (O_1935,N_18145,N_19183);
and UO_1936 (O_1936,N_19321,N_18134);
nand UO_1937 (O_1937,N_19712,N_19658);
xor UO_1938 (O_1938,N_18533,N_19545);
nor UO_1939 (O_1939,N_18228,N_19554);
nor UO_1940 (O_1940,N_19383,N_19350);
nand UO_1941 (O_1941,N_19816,N_19224);
nor UO_1942 (O_1942,N_19407,N_19672);
nor UO_1943 (O_1943,N_18355,N_18636);
or UO_1944 (O_1944,N_19158,N_19280);
nand UO_1945 (O_1945,N_19675,N_19055);
xor UO_1946 (O_1946,N_19664,N_18774);
xnor UO_1947 (O_1947,N_18040,N_18652);
or UO_1948 (O_1948,N_19390,N_19835);
nand UO_1949 (O_1949,N_18723,N_19209);
xnor UO_1950 (O_1950,N_19838,N_19540);
or UO_1951 (O_1951,N_18238,N_19779);
nor UO_1952 (O_1952,N_19643,N_19359);
xor UO_1953 (O_1953,N_18149,N_19073);
nand UO_1954 (O_1954,N_18756,N_18402);
xnor UO_1955 (O_1955,N_18665,N_19745);
and UO_1956 (O_1956,N_19589,N_18475);
and UO_1957 (O_1957,N_19712,N_19343);
and UO_1958 (O_1958,N_19843,N_19925);
nand UO_1959 (O_1959,N_18578,N_18444);
or UO_1960 (O_1960,N_18856,N_19469);
or UO_1961 (O_1961,N_19945,N_18071);
and UO_1962 (O_1962,N_19727,N_18027);
nand UO_1963 (O_1963,N_18495,N_18176);
or UO_1964 (O_1964,N_19103,N_18995);
and UO_1965 (O_1965,N_18690,N_19535);
and UO_1966 (O_1966,N_19975,N_19763);
nand UO_1967 (O_1967,N_19107,N_19652);
xor UO_1968 (O_1968,N_19677,N_19905);
nand UO_1969 (O_1969,N_18226,N_19414);
and UO_1970 (O_1970,N_19548,N_19471);
nor UO_1971 (O_1971,N_18898,N_19660);
and UO_1972 (O_1972,N_18357,N_18287);
nand UO_1973 (O_1973,N_18774,N_19185);
nand UO_1974 (O_1974,N_18173,N_19564);
nor UO_1975 (O_1975,N_18431,N_18964);
nor UO_1976 (O_1976,N_18759,N_19082);
xor UO_1977 (O_1977,N_18631,N_19098);
and UO_1978 (O_1978,N_19141,N_18694);
xnor UO_1979 (O_1979,N_19836,N_18822);
nand UO_1980 (O_1980,N_19070,N_19105);
and UO_1981 (O_1981,N_19967,N_19033);
or UO_1982 (O_1982,N_18449,N_19676);
nor UO_1983 (O_1983,N_18689,N_19627);
or UO_1984 (O_1984,N_18741,N_18085);
nor UO_1985 (O_1985,N_19546,N_18722);
xnor UO_1986 (O_1986,N_18190,N_19788);
or UO_1987 (O_1987,N_19980,N_19705);
nand UO_1988 (O_1988,N_18091,N_18742);
nand UO_1989 (O_1989,N_18587,N_18272);
nand UO_1990 (O_1990,N_19098,N_19022);
and UO_1991 (O_1991,N_19807,N_19287);
or UO_1992 (O_1992,N_18033,N_19729);
nand UO_1993 (O_1993,N_18910,N_18681);
nor UO_1994 (O_1994,N_18707,N_18039);
or UO_1995 (O_1995,N_19798,N_18402);
nand UO_1996 (O_1996,N_19325,N_19047);
and UO_1997 (O_1997,N_18266,N_18457);
nor UO_1998 (O_1998,N_19910,N_18605);
xor UO_1999 (O_1999,N_18155,N_19413);
nand UO_2000 (O_2000,N_19275,N_19252);
nor UO_2001 (O_2001,N_18209,N_19340);
or UO_2002 (O_2002,N_18259,N_19562);
xor UO_2003 (O_2003,N_18264,N_19050);
nor UO_2004 (O_2004,N_19327,N_19440);
nor UO_2005 (O_2005,N_19029,N_18984);
nand UO_2006 (O_2006,N_18142,N_18128);
and UO_2007 (O_2007,N_18771,N_18159);
nand UO_2008 (O_2008,N_18594,N_18458);
nor UO_2009 (O_2009,N_19682,N_19519);
and UO_2010 (O_2010,N_18783,N_18136);
or UO_2011 (O_2011,N_19526,N_19749);
and UO_2012 (O_2012,N_19697,N_18659);
nand UO_2013 (O_2013,N_18481,N_18556);
or UO_2014 (O_2014,N_18371,N_18386);
or UO_2015 (O_2015,N_18291,N_19237);
and UO_2016 (O_2016,N_19285,N_18814);
and UO_2017 (O_2017,N_18256,N_18517);
nor UO_2018 (O_2018,N_19920,N_18434);
or UO_2019 (O_2019,N_18867,N_18904);
nor UO_2020 (O_2020,N_18236,N_19781);
or UO_2021 (O_2021,N_19599,N_18735);
or UO_2022 (O_2022,N_18990,N_19386);
nand UO_2023 (O_2023,N_19010,N_18595);
or UO_2024 (O_2024,N_18673,N_18326);
or UO_2025 (O_2025,N_19284,N_18217);
nor UO_2026 (O_2026,N_18300,N_19390);
nand UO_2027 (O_2027,N_18089,N_19560);
nand UO_2028 (O_2028,N_19735,N_18208);
nand UO_2029 (O_2029,N_19386,N_19218);
nor UO_2030 (O_2030,N_19824,N_18305);
and UO_2031 (O_2031,N_19677,N_19848);
xor UO_2032 (O_2032,N_19622,N_18358);
nand UO_2033 (O_2033,N_18326,N_19162);
xor UO_2034 (O_2034,N_19455,N_19911);
nand UO_2035 (O_2035,N_19593,N_19012);
and UO_2036 (O_2036,N_19194,N_18188);
and UO_2037 (O_2037,N_18376,N_18738);
nand UO_2038 (O_2038,N_19232,N_19077);
nor UO_2039 (O_2039,N_18014,N_18000);
and UO_2040 (O_2040,N_18301,N_18636);
nor UO_2041 (O_2041,N_19176,N_18095);
nor UO_2042 (O_2042,N_19279,N_18841);
and UO_2043 (O_2043,N_19879,N_19755);
or UO_2044 (O_2044,N_19739,N_19618);
nor UO_2045 (O_2045,N_19351,N_18700);
nor UO_2046 (O_2046,N_18419,N_18971);
and UO_2047 (O_2047,N_18017,N_19809);
nand UO_2048 (O_2048,N_19532,N_18761);
or UO_2049 (O_2049,N_18220,N_18874);
nand UO_2050 (O_2050,N_18060,N_18742);
nor UO_2051 (O_2051,N_19067,N_18336);
or UO_2052 (O_2052,N_18741,N_18420);
and UO_2053 (O_2053,N_18469,N_18410);
or UO_2054 (O_2054,N_19450,N_18520);
and UO_2055 (O_2055,N_19496,N_19298);
and UO_2056 (O_2056,N_19664,N_19235);
nor UO_2057 (O_2057,N_18029,N_19558);
and UO_2058 (O_2058,N_18387,N_19718);
nand UO_2059 (O_2059,N_18256,N_19952);
or UO_2060 (O_2060,N_18223,N_18033);
nand UO_2061 (O_2061,N_19037,N_18557);
or UO_2062 (O_2062,N_19862,N_18793);
nor UO_2063 (O_2063,N_18168,N_19466);
nor UO_2064 (O_2064,N_18181,N_19342);
nor UO_2065 (O_2065,N_19405,N_19336);
and UO_2066 (O_2066,N_18366,N_19006);
or UO_2067 (O_2067,N_19904,N_19545);
nor UO_2068 (O_2068,N_19147,N_18981);
xnor UO_2069 (O_2069,N_18205,N_19545);
and UO_2070 (O_2070,N_18884,N_18117);
or UO_2071 (O_2071,N_18127,N_19303);
nor UO_2072 (O_2072,N_19522,N_19231);
or UO_2073 (O_2073,N_18067,N_19507);
nor UO_2074 (O_2074,N_19520,N_19813);
xor UO_2075 (O_2075,N_19613,N_18536);
nand UO_2076 (O_2076,N_18554,N_18776);
or UO_2077 (O_2077,N_18835,N_19315);
nor UO_2078 (O_2078,N_19304,N_18217);
and UO_2079 (O_2079,N_19135,N_18440);
or UO_2080 (O_2080,N_19853,N_19654);
or UO_2081 (O_2081,N_18731,N_19904);
or UO_2082 (O_2082,N_18644,N_18034);
nor UO_2083 (O_2083,N_19583,N_19565);
and UO_2084 (O_2084,N_18543,N_19151);
nor UO_2085 (O_2085,N_19084,N_19243);
nand UO_2086 (O_2086,N_18658,N_18136);
nand UO_2087 (O_2087,N_19329,N_18753);
nor UO_2088 (O_2088,N_19423,N_18907);
nand UO_2089 (O_2089,N_18808,N_19964);
or UO_2090 (O_2090,N_19846,N_19870);
nor UO_2091 (O_2091,N_18026,N_19856);
nor UO_2092 (O_2092,N_18623,N_19636);
xnor UO_2093 (O_2093,N_18927,N_18917);
or UO_2094 (O_2094,N_18836,N_18716);
nand UO_2095 (O_2095,N_18094,N_18962);
or UO_2096 (O_2096,N_19651,N_19293);
nor UO_2097 (O_2097,N_18125,N_19374);
nor UO_2098 (O_2098,N_18908,N_18633);
or UO_2099 (O_2099,N_18351,N_19291);
or UO_2100 (O_2100,N_19040,N_18115);
nor UO_2101 (O_2101,N_18071,N_19781);
xor UO_2102 (O_2102,N_19286,N_18258);
or UO_2103 (O_2103,N_19953,N_18197);
nor UO_2104 (O_2104,N_18832,N_19652);
nor UO_2105 (O_2105,N_19420,N_18620);
xor UO_2106 (O_2106,N_18175,N_19248);
and UO_2107 (O_2107,N_18669,N_19273);
and UO_2108 (O_2108,N_18863,N_19400);
and UO_2109 (O_2109,N_19730,N_19004);
xnor UO_2110 (O_2110,N_19915,N_18315);
nor UO_2111 (O_2111,N_19151,N_18905);
and UO_2112 (O_2112,N_18234,N_18331);
xor UO_2113 (O_2113,N_18157,N_19464);
nand UO_2114 (O_2114,N_18144,N_18919);
and UO_2115 (O_2115,N_19119,N_19121);
nor UO_2116 (O_2116,N_18984,N_18536);
xnor UO_2117 (O_2117,N_19926,N_18119);
nor UO_2118 (O_2118,N_19081,N_18676);
and UO_2119 (O_2119,N_19286,N_19025);
and UO_2120 (O_2120,N_18540,N_19514);
or UO_2121 (O_2121,N_19906,N_18181);
or UO_2122 (O_2122,N_19691,N_18517);
nand UO_2123 (O_2123,N_18107,N_19519);
and UO_2124 (O_2124,N_19835,N_19993);
nand UO_2125 (O_2125,N_19182,N_19134);
or UO_2126 (O_2126,N_19275,N_18028);
and UO_2127 (O_2127,N_19761,N_19348);
or UO_2128 (O_2128,N_18705,N_19220);
or UO_2129 (O_2129,N_19655,N_18750);
or UO_2130 (O_2130,N_19447,N_19865);
nand UO_2131 (O_2131,N_18744,N_19809);
nand UO_2132 (O_2132,N_18433,N_19522);
nor UO_2133 (O_2133,N_19366,N_19860);
or UO_2134 (O_2134,N_18824,N_18458);
and UO_2135 (O_2135,N_19089,N_18906);
nor UO_2136 (O_2136,N_19346,N_19909);
and UO_2137 (O_2137,N_18654,N_19970);
or UO_2138 (O_2138,N_18174,N_19182);
nor UO_2139 (O_2139,N_18604,N_19759);
or UO_2140 (O_2140,N_18556,N_18643);
nor UO_2141 (O_2141,N_19657,N_18308);
nand UO_2142 (O_2142,N_18422,N_19401);
nand UO_2143 (O_2143,N_19847,N_18067);
or UO_2144 (O_2144,N_18877,N_19966);
and UO_2145 (O_2145,N_18064,N_18474);
or UO_2146 (O_2146,N_19277,N_18255);
or UO_2147 (O_2147,N_19003,N_18571);
or UO_2148 (O_2148,N_18675,N_18742);
nor UO_2149 (O_2149,N_19978,N_19720);
and UO_2150 (O_2150,N_19540,N_19726);
xnor UO_2151 (O_2151,N_19501,N_19575);
xor UO_2152 (O_2152,N_18838,N_18744);
and UO_2153 (O_2153,N_19997,N_18802);
xnor UO_2154 (O_2154,N_18432,N_19379);
nand UO_2155 (O_2155,N_19121,N_19141);
nand UO_2156 (O_2156,N_18513,N_18576);
nor UO_2157 (O_2157,N_19393,N_19802);
and UO_2158 (O_2158,N_18794,N_19186);
nand UO_2159 (O_2159,N_19334,N_18763);
or UO_2160 (O_2160,N_19513,N_18686);
and UO_2161 (O_2161,N_18852,N_19165);
or UO_2162 (O_2162,N_18490,N_19385);
nor UO_2163 (O_2163,N_19103,N_19670);
nor UO_2164 (O_2164,N_19604,N_18893);
xnor UO_2165 (O_2165,N_18971,N_18553);
xnor UO_2166 (O_2166,N_18052,N_19541);
nand UO_2167 (O_2167,N_18807,N_19289);
or UO_2168 (O_2168,N_18411,N_18010);
xnor UO_2169 (O_2169,N_19931,N_18585);
and UO_2170 (O_2170,N_18820,N_19738);
nand UO_2171 (O_2171,N_18496,N_19047);
nor UO_2172 (O_2172,N_18868,N_18576);
nand UO_2173 (O_2173,N_19308,N_19789);
nand UO_2174 (O_2174,N_18562,N_18496);
or UO_2175 (O_2175,N_18945,N_18939);
and UO_2176 (O_2176,N_19106,N_18873);
nand UO_2177 (O_2177,N_19205,N_18328);
xnor UO_2178 (O_2178,N_18795,N_19809);
and UO_2179 (O_2179,N_18611,N_19229);
or UO_2180 (O_2180,N_19532,N_18267);
and UO_2181 (O_2181,N_18987,N_19331);
nor UO_2182 (O_2182,N_18604,N_18675);
and UO_2183 (O_2183,N_18485,N_19350);
xnor UO_2184 (O_2184,N_19175,N_19834);
nand UO_2185 (O_2185,N_19659,N_18872);
or UO_2186 (O_2186,N_19641,N_18135);
and UO_2187 (O_2187,N_18539,N_19760);
nand UO_2188 (O_2188,N_19662,N_19505);
or UO_2189 (O_2189,N_18477,N_19496);
or UO_2190 (O_2190,N_18924,N_18657);
nor UO_2191 (O_2191,N_18773,N_18281);
and UO_2192 (O_2192,N_18342,N_18653);
nand UO_2193 (O_2193,N_18385,N_19776);
and UO_2194 (O_2194,N_19884,N_19368);
and UO_2195 (O_2195,N_19413,N_18772);
nand UO_2196 (O_2196,N_19806,N_18174);
nor UO_2197 (O_2197,N_18555,N_18387);
nand UO_2198 (O_2198,N_18633,N_18079);
nor UO_2199 (O_2199,N_18319,N_19931);
xor UO_2200 (O_2200,N_19427,N_19215);
and UO_2201 (O_2201,N_18692,N_18500);
nand UO_2202 (O_2202,N_18023,N_19121);
and UO_2203 (O_2203,N_19304,N_19363);
nor UO_2204 (O_2204,N_18878,N_19090);
or UO_2205 (O_2205,N_18999,N_18481);
nor UO_2206 (O_2206,N_18761,N_18898);
or UO_2207 (O_2207,N_19870,N_19392);
or UO_2208 (O_2208,N_19220,N_18532);
nand UO_2209 (O_2209,N_19287,N_19702);
nor UO_2210 (O_2210,N_18908,N_18281);
nor UO_2211 (O_2211,N_19549,N_18615);
or UO_2212 (O_2212,N_18281,N_19685);
or UO_2213 (O_2213,N_18443,N_18377);
nor UO_2214 (O_2214,N_19945,N_19752);
nand UO_2215 (O_2215,N_18244,N_19219);
nand UO_2216 (O_2216,N_19753,N_18579);
nor UO_2217 (O_2217,N_18262,N_18705);
nor UO_2218 (O_2218,N_19322,N_19418);
nand UO_2219 (O_2219,N_19993,N_18925);
or UO_2220 (O_2220,N_18883,N_18184);
nor UO_2221 (O_2221,N_18443,N_19322);
and UO_2222 (O_2222,N_19037,N_19052);
and UO_2223 (O_2223,N_18590,N_19026);
and UO_2224 (O_2224,N_18505,N_19097);
or UO_2225 (O_2225,N_18443,N_19228);
nand UO_2226 (O_2226,N_18093,N_19564);
nor UO_2227 (O_2227,N_19425,N_18214);
xor UO_2228 (O_2228,N_19085,N_18440);
or UO_2229 (O_2229,N_18874,N_18741);
or UO_2230 (O_2230,N_18619,N_19723);
or UO_2231 (O_2231,N_19435,N_19097);
or UO_2232 (O_2232,N_18260,N_19033);
nand UO_2233 (O_2233,N_19679,N_18602);
xnor UO_2234 (O_2234,N_19309,N_18785);
nor UO_2235 (O_2235,N_19069,N_19238);
nor UO_2236 (O_2236,N_18519,N_19752);
nand UO_2237 (O_2237,N_19540,N_18778);
xnor UO_2238 (O_2238,N_18745,N_19145);
nand UO_2239 (O_2239,N_19705,N_18310);
and UO_2240 (O_2240,N_18131,N_19688);
nand UO_2241 (O_2241,N_18191,N_18860);
nand UO_2242 (O_2242,N_19972,N_19612);
or UO_2243 (O_2243,N_18027,N_19987);
and UO_2244 (O_2244,N_19988,N_19614);
xnor UO_2245 (O_2245,N_18944,N_18815);
nand UO_2246 (O_2246,N_19120,N_19358);
or UO_2247 (O_2247,N_19943,N_18924);
and UO_2248 (O_2248,N_19828,N_18471);
and UO_2249 (O_2249,N_19523,N_18417);
or UO_2250 (O_2250,N_19006,N_18881);
and UO_2251 (O_2251,N_19938,N_19091);
nand UO_2252 (O_2252,N_18486,N_19899);
and UO_2253 (O_2253,N_19228,N_19081);
and UO_2254 (O_2254,N_18458,N_19961);
and UO_2255 (O_2255,N_19966,N_18803);
xnor UO_2256 (O_2256,N_18432,N_19092);
nor UO_2257 (O_2257,N_18086,N_18983);
nor UO_2258 (O_2258,N_19006,N_19822);
nor UO_2259 (O_2259,N_18047,N_19874);
xor UO_2260 (O_2260,N_19153,N_19277);
and UO_2261 (O_2261,N_19277,N_18300);
nand UO_2262 (O_2262,N_18667,N_19764);
nor UO_2263 (O_2263,N_18710,N_19542);
nor UO_2264 (O_2264,N_18860,N_19624);
and UO_2265 (O_2265,N_18751,N_18661);
nand UO_2266 (O_2266,N_18299,N_19674);
nand UO_2267 (O_2267,N_18837,N_19664);
nand UO_2268 (O_2268,N_18188,N_19610);
nand UO_2269 (O_2269,N_18768,N_19973);
nand UO_2270 (O_2270,N_18663,N_19645);
nor UO_2271 (O_2271,N_19072,N_19113);
xnor UO_2272 (O_2272,N_18661,N_19974);
xor UO_2273 (O_2273,N_18196,N_19249);
nor UO_2274 (O_2274,N_18429,N_18997);
nand UO_2275 (O_2275,N_18881,N_18762);
or UO_2276 (O_2276,N_18635,N_19236);
nand UO_2277 (O_2277,N_18812,N_18210);
or UO_2278 (O_2278,N_19780,N_18195);
or UO_2279 (O_2279,N_18554,N_18831);
nand UO_2280 (O_2280,N_19542,N_18549);
xor UO_2281 (O_2281,N_18979,N_19872);
nor UO_2282 (O_2282,N_18572,N_18262);
and UO_2283 (O_2283,N_19970,N_18311);
or UO_2284 (O_2284,N_18865,N_18896);
nor UO_2285 (O_2285,N_18749,N_18671);
or UO_2286 (O_2286,N_19972,N_18655);
or UO_2287 (O_2287,N_18498,N_18374);
and UO_2288 (O_2288,N_19589,N_19479);
or UO_2289 (O_2289,N_19199,N_19732);
and UO_2290 (O_2290,N_18149,N_19118);
and UO_2291 (O_2291,N_18731,N_19123);
nor UO_2292 (O_2292,N_18945,N_19977);
nor UO_2293 (O_2293,N_18938,N_19288);
and UO_2294 (O_2294,N_18694,N_18046);
and UO_2295 (O_2295,N_18160,N_19265);
nand UO_2296 (O_2296,N_19301,N_19931);
and UO_2297 (O_2297,N_18253,N_19046);
nand UO_2298 (O_2298,N_19018,N_18115);
and UO_2299 (O_2299,N_19875,N_19518);
and UO_2300 (O_2300,N_18677,N_18236);
nand UO_2301 (O_2301,N_18435,N_18199);
or UO_2302 (O_2302,N_19138,N_19006);
nor UO_2303 (O_2303,N_18176,N_18883);
nand UO_2304 (O_2304,N_19745,N_19558);
xnor UO_2305 (O_2305,N_18567,N_19203);
nor UO_2306 (O_2306,N_18306,N_19512);
nor UO_2307 (O_2307,N_18460,N_18634);
xnor UO_2308 (O_2308,N_19518,N_19641);
and UO_2309 (O_2309,N_18339,N_19767);
nor UO_2310 (O_2310,N_19865,N_19039);
nor UO_2311 (O_2311,N_18247,N_18343);
nor UO_2312 (O_2312,N_18654,N_19245);
or UO_2313 (O_2313,N_19299,N_19414);
and UO_2314 (O_2314,N_19149,N_19576);
and UO_2315 (O_2315,N_19110,N_19774);
nand UO_2316 (O_2316,N_19614,N_18669);
and UO_2317 (O_2317,N_18727,N_18698);
or UO_2318 (O_2318,N_18915,N_19770);
and UO_2319 (O_2319,N_19913,N_18719);
nand UO_2320 (O_2320,N_19821,N_18266);
nand UO_2321 (O_2321,N_19637,N_18368);
nand UO_2322 (O_2322,N_18137,N_19095);
nand UO_2323 (O_2323,N_19626,N_18442);
xor UO_2324 (O_2324,N_19036,N_19898);
xnor UO_2325 (O_2325,N_18490,N_18338);
nand UO_2326 (O_2326,N_18128,N_19371);
nor UO_2327 (O_2327,N_19040,N_19032);
nand UO_2328 (O_2328,N_18856,N_19196);
and UO_2329 (O_2329,N_19082,N_19806);
and UO_2330 (O_2330,N_18078,N_19408);
xnor UO_2331 (O_2331,N_19349,N_18321);
xor UO_2332 (O_2332,N_18672,N_19839);
or UO_2333 (O_2333,N_19125,N_18835);
nand UO_2334 (O_2334,N_18775,N_18515);
nand UO_2335 (O_2335,N_18750,N_19877);
nor UO_2336 (O_2336,N_19430,N_18380);
and UO_2337 (O_2337,N_18165,N_19038);
and UO_2338 (O_2338,N_19610,N_19902);
nand UO_2339 (O_2339,N_19010,N_18717);
or UO_2340 (O_2340,N_19265,N_18871);
nor UO_2341 (O_2341,N_18622,N_18707);
nand UO_2342 (O_2342,N_19812,N_18319);
and UO_2343 (O_2343,N_19004,N_19915);
or UO_2344 (O_2344,N_19217,N_19979);
nor UO_2345 (O_2345,N_19775,N_18381);
nand UO_2346 (O_2346,N_19381,N_18920);
or UO_2347 (O_2347,N_18704,N_19252);
nand UO_2348 (O_2348,N_18762,N_18080);
nand UO_2349 (O_2349,N_19613,N_19877);
or UO_2350 (O_2350,N_18394,N_19763);
and UO_2351 (O_2351,N_18791,N_18518);
nand UO_2352 (O_2352,N_18886,N_19338);
nand UO_2353 (O_2353,N_18221,N_18029);
nand UO_2354 (O_2354,N_18993,N_18053);
nor UO_2355 (O_2355,N_19899,N_18314);
or UO_2356 (O_2356,N_19219,N_18260);
and UO_2357 (O_2357,N_18207,N_19366);
nor UO_2358 (O_2358,N_18068,N_19874);
nor UO_2359 (O_2359,N_19231,N_18046);
or UO_2360 (O_2360,N_18876,N_18889);
and UO_2361 (O_2361,N_19941,N_18645);
and UO_2362 (O_2362,N_18391,N_18746);
xor UO_2363 (O_2363,N_19957,N_19293);
xor UO_2364 (O_2364,N_18068,N_19720);
and UO_2365 (O_2365,N_18162,N_19082);
nand UO_2366 (O_2366,N_19761,N_18389);
or UO_2367 (O_2367,N_18724,N_19803);
nand UO_2368 (O_2368,N_18202,N_19915);
nand UO_2369 (O_2369,N_19394,N_19921);
nand UO_2370 (O_2370,N_19112,N_18217);
nand UO_2371 (O_2371,N_19327,N_18593);
nor UO_2372 (O_2372,N_19310,N_18104);
nand UO_2373 (O_2373,N_19045,N_19934);
nand UO_2374 (O_2374,N_18927,N_18510);
nand UO_2375 (O_2375,N_19931,N_19097);
xnor UO_2376 (O_2376,N_19570,N_19322);
xnor UO_2377 (O_2377,N_19815,N_19677);
xor UO_2378 (O_2378,N_19004,N_19385);
nand UO_2379 (O_2379,N_18743,N_18924);
nor UO_2380 (O_2380,N_19537,N_19643);
nand UO_2381 (O_2381,N_18436,N_19982);
nand UO_2382 (O_2382,N_19428,N_19797);
xor UO_2383 (O_2383,N_19503,N_19303);
xor UO_2384 (O_2384,N_19189,N_19670);
or UO_2385 (O_2385,N_18817,N_18914);
nand UO_2386 (O_2386,N_18537,N_19395);
nand UO_2387 (O_2387,N_19065,N_18108);
or UO_2388 (O_2388,N_19915,N_19667);
nor UO_2389 (O_2389,N_18106,N_19539);
nand UO_2390 (O_2390,N_19880,N_18331);
nand UO_2391 (O_2391,N_19820,N_19208);
or UO_2392 (O_2392,N_19048,N_18372);
nor UO_2393 (O_2393,N_18983,N_18679);
nor UO_2394 (O_2394,N_18088,N_18877);
nor UO_2395 (O_2395,N_18111,N_19938);
or UO_2396 (O_2396,N_19452,N_19197);
nand UO_2397 (O_2397,N_18508,N_19444);
nor UO_2398 (O_2398,N_19084,N_18016);
and UO_2399 (O_2399,N_19032,N_18417);
and UO_2400 (O_2400,N_19394,N_19849);
nor UO_2401 (O_2401,N_19304,N_18670);
nor UO_2402 (O_2402,N_19912,N_19456);
nor UO_2403 (O_2403,N_18712,N_18192);
or UO_2404 (O_2404,N_19939,N_19809);
and UO_2405 (O_2405,N_18366,N_19920);
and UO_2406 (O_2406,N_19743,N_19557);
and UO_2407 (O_2407,N_18329,N_18144);
or UO_2408 (O_2408,N_18507,N_19902);
or UO_2409 (O_2409,N_19178,N_18575);
xnor UO_2410 (O_2410,N_18713,N_19206);
or UO_2411 (O_2411,N_18107,N_18853);
or UO_2412 (O_2412,N_19557,N_19671);
xnor UO_2413 (O_2413,N_18738,N_19669);
and UO_2414 (O_2414,N_19198,N_18636);
nor UO_2415 (O_2415,N_19860,N_19075);
and UO_2416 (O_2416,N_19245,N_19111);
or UO_2417 (O_2417,N_18274,N_18006);
or UO_2418 (O_2418,N_19274,N_18842);
nor UO_2419 (O_2419,N_18680,N_18781);
and UO_2420 (O_2420,N_19090,N_18450);
nor UO_2421 (O_2421,N_19779,N_19982);
and UO_2422 (O_2422,N_19079,N_19808);
and UO_2423 (O_2423,N_19746,N_19755);
or UO_2424 (O_2424,N_18035,N_19710);
and UO_2425 (O_2425,N_18764,N_19768);
xnor UO_2426 (O_2426,N_18840,N_19858);
nor UO_2427 (O_2427,N_18745,N_19874);
nor UO_2428 (O_2428,N_18933,N_18039);
and UO_2429 (O_2429,N_19404,N_19407);
nor UO_2430 (O_2430,N_19607,N_18119);
and UO_2431 (O_2431,N_19730,N_18955);
and UO_2432 (O_2432,N_19233,N_19871);
and UO_2433 (O_2433,N_18293,N_19320);
nor UO_2434 (O_2434,N_18782,N_18437);
and UO_2435 (O_2435,N_19521,N_18740);
xor UO_2436 (O_2436,N_19208,N_19641);
nor UO_2437 (O_2437,N_19337,N_18852);
xnor UO_2438 (O_2438,N_18852,N_19117);
and UO_2439 (O_2439,N_19839,N_18179);
and UO_2440 (O_2440,N_19619,N_19062);
or UO_2441 (O_2441,N_18535,N_19648);
nand UO_2442 (O_2442,N_18555,N_18782);
and UO_2443 (O_2443,N_19378,N_18974);
or UO_2444 (O_2444,N_19670,N_19245);
nand UO_2445 (O_2445,N_19729,N_18208);
or UO_2446 (O_2446,N_19903,N_18967);
or UO_2447 (O_2447,N_18055,N_19384);
nand UO_2448 (O_2448,N_19175,N_18002);
nor UO_2449 (O_2449,N_19411,N_19560);
and UO_2450 (O_2450,N_18928,N_19756);
nor UO_2451 (O_2451,N_19539,N_18149);
and UO_2452 (O_2452,N_18785,N_19315);
nor UO_2453 (O_2453,N_19621,N_18332);
and UO_2454 (O_2454,N_19688,N_18476);
nor UO_2455 (O_2455,N_19187,N_19832);
and UO_2456 (O_2456,N_19964,N_18457);
or UO_2457 (O_2457,N_18696,N_18689);
and UO_2458 (O_2458,N_19968,N_18784);
nand UO_2459 (O_2459,N_19279,N_18142);
and UO_2460 (O_2460,N_19495,N_18495);
or UO_2461 (O_2461,N_19277,N_19830);
and UO_2462 (O_2462,N_18096,N_18215);
or UO_2463 (O_2463,N_18392,N_19798);
or UO_2464 (O_2464,N_19200,N_18778);
and UO_2465 (O_2465,N_19560,N_18419);
nand UO_2466 (O_2466,N_19117,N_19444);
or UO_2467 (O_2467,N_19950,N_19584);
nand UO_2468 (O_2468,N_19909,N_18309);
xnor UO_2469 (O_2469,N_19041,N_18939);
nand UO_2470 (O_2470,N_19302,N_18207);
nor UO_2471 (O_2471,N_18202,N_19354);
and UO_2472 (O_2472,N_19808,N_18322);
and UO_2473 (O_2473,N_18300,N_19967);
nor UO_2474 (O_2474,N_19366,N_19229);
nand UO_2475 (O_2475,N_19098,N_18345);
nor UO_2476 (O_2476,N_19974,N_19216);
or UO_2477 (O_2477,N_18331,N_18210);
or UO_2478 (O_2478,N_19782,N_18066);
xnor UO_2479 (O_2479,N_19725,N_19342);
or UO_2480 (O_2480,N_18328,N_19811);
nor UO_2481 (O_2481,N_18310,N_19870);
nand UO_2482 (O_2482,N_19302,N_18426);
xor UO_2483 (O_2483,N_19521,N_19375);
nor UO_2484 (O_2484,N_18146,N_18802);
nand UO_2485 (O_2485,N_18420,N_18317);
and UO_2486 (O_2486,N_18540,N_19057);
or UO_2487 (O_2487,N_18912,N_19918);
xor UO_2488 (O_2488,N_18874,N_18379);
nand UO_2489 (O_2489,N_18932,N_18825);
nor UO_2490 (O_2490,N_18785,N_18577);
nor UO_2491 (O_2491,N_18638,N_18966);
and UO_2492 (O_2492,N_19335,N_19973);
and UO_2493 (O_2493,N_18479,N_18368);
and UO_2494 (O_2494,N_18730,N_19393);
or UO_2495 (O_2495,N_19487,N_18966);
xor UO_2496 (O_2496,N_18736,N_19868);
nor UO_2497 (O_2497,N_18235,N_18192);
xnor UO_2498 (O_2498,N_19530,N_19383);
or UO_2499 (O_2499,N_18687,N_18381);
endmodule