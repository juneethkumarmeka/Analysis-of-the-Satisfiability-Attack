module basic_1500_15000_2000_5_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_716,In_1104);
nor U1 (N_1,In_1055,In_1306);
nand U2 (N_2,In_464,In_854);
or U3 (N_3,In_1033,In_1046);
or U4 (N_4,In_1018,In_863);
nand U5 (N_5,In_64,In_879);
and U6 (N_6,In_1009,In_1166);
or U7 (N_7,In_1290,In_1432);
nor U8 (N_8,In_1224,In_1217);
or U9 (N_9,In_717,In_1404);
or U10 (N_10,In_974,In_189);
and U11 (N_11,In_1322,In_669);
and U12 (N_12,In_1115,In_810);
nor U13 (N_13,In_1072,In_618);
nor U14 (N_14,In_846,In_1434);
nand U15 (N_15,In_921,In_1277);
or U16 (N_16,In_559,In_1351);
nand U17 (N_17,In_88,In_690);
and U18 (N_18,In_606,In_406);
nor U19 (N_19,In_775,In_1303);
nor U20 (N_20,In_1028,In_154);
or U21 (N_21,In_310,In_92);
and U22 (N_22,In_1328,In_144);
nand U23 (N_23,In_1472,In_1423);
and U24 (N_24,In_355,In_434);
or U25 (N_25,In_1263,In_495);
or U26 (N_26,In_897,In_23);
nand U27 (N_27,In_226,In_421);
or U28 (N_28,In_264,In_306);
and U29 (N_29,In_31,In_1309);
nand U30 (N_30,In_886,In_1342);
nor U31 (N_31,In_1395,In_590);
nand U32 (N_32,In_707,In_1268);
and U33 (N_33,In_530,In_165);
and U34 (N_34,In_484,In_54);
or U35 (N_35,In_76,In_311);
nor U36 (N_36,In_1105,In_303);
and U37 (N_37,In_572,In_890);
or U38 (N_38,In_1481,In_1243);
nor U39 (N_39,In_944,In_1120);
xnor U40 (N_40,In_515,In_777);
and U41 (N_41,In_156,In_192);
and U42 (N_42,In_1275,In_1379);
or U43 (N_43,In_754,In_546);
or U44 (N_44,In_528,In_688);
or U45 (N_45,In_1215,In_933);
nor U46 (N_46,In_229,In_1220);
or U47 (N_47,In_1278,In_168);
or U48 (N_48,In_1394,In_809);
nand U49 (N_49,In_969,In_751);
or U50 (N_50,In_1272,In_374);
or U51 (N_51,In_909,In_554);
or U52 (N_52,In_654,In_788);
and U53 (N_53,In_1377,In_1208);
and U54 (N_54,In_170,In_451);
nand U55 (N_55,In_1134,In_230);
nor U56 (N_56,In_1043,In_115);
nand U57 (N_57,In_1386,In_345);
nand U58 (N_58,In_866,In_1122);
and U59 (N_59,In_992,In_384);
and U60 (N_60,In_29,In_1052);
nor U61 (N_61,In_468,In_847);
nor U62 (N_62,In_758,In_638);
or U63 (N_63,In_409,In_1267);
nand U64 (N_64,In_1123,In_1416);
nor U65 (N_65,In_1388,In_1262);
nand U66 (N_66,In_390,In_212);
nand U67 (N_67,In_475,In_242);
and U68 (N_68,In_348,In_919);
nor U69 (N_69,In_161,In_822);
nand U70 (N_70,In_857,In_198);
nand U71 (N_71,In_1013,In_637);
and U72 (N_72,In_146,In_1152);
and U73 (N_73,In_1056,In_1173);
and U74 (N_74,In_131,In_1470);
or U75 (N_75,In_49,In_1171);
or U76 (N_76,In_838,In_1344);
nand U77 (N_77,In_645,In_12);
or U78 (N_78,In_816,In_1227);
or U79 (N_79,In_1437,In_63);
and U80 (N_80,In_429,In_999);
xnor U81 (N_81,In_524,In_650);
or U82 (N_82,In_534,In_153);
nor U83 (N_83,In_947,In_811);
or U84 (N_84,In_1447,In_1069);
or U85 (N_85,In_493,In_1011);
nand U86 (N_86,In_1453,In_61);
or U87 (N_87,In_556,In_1025);
nor U88 (N_88,In_594,In_157);
nand U89 (N_89,In_281,In_480);
nand U90 (N_90,In_730,In_10);
nand U91 (N_91,In_1459,In_128);
and U92 (N_92,In_1298,In_248);
nand U93 (N_93,In_363,In_139);
and U94 (N_94,In_881,In_911);
nor U95 (N_95,In_1064,In_38);
or U96 (N_96,In_727,In_693);
or U97 (N_97,In_1361,In_724);
or U98 (N_98,In_1355,In_1477);
and U99 (N_99,In_85,In_448);
and U100 (N_100,In_1330,In_1476);
nor U101 (N_101,In_603,In_1287);
or U102 (N_102,In_625,In_744);
or U103 (N_103,In_83,In_1381);
or U104 (N_104,In_50,In_353);
nor U105 (N_105,In_623,In_400);
and U106 (N_106,In_1362,In_71);
or U107 (N_107,In_132,In_753);
nand U108 (N_108,In_986,In_1271);
or U109 (N_109,In_1113,In_268);
nor U110 (N_110,In_864,In_507);
nor U111 (N_111,In_75,In_245);
nor U112 (N_112,In_496,In_426);
nand U113 (N_113,In_1027,In_516);
nand U114 (N_114,In_1291,In_1062);
nand U115 (N_115,In_492,In_1185);
or U116 (N_116,In_734,In_1390);
nor U117 (N_117,In_697,In_845);
nor U118 (N_118,In_551,In_652);
or U119 (N_119,In_1392,In_47);
and U120 (N_120,In_917,In_547);
nand U121 (N_121,In_1341,In_494);
nor U122 (N_122,In_955,In_659);
and U123 (N_123,In_438,In_487);
and U124 (N_124,In_685,In_446);
nor U125 (N_125,In_382,In_1418);
or U126 (N_126,In_1373,In_276);
nand U127 (N_127,In_378,In_781);
nor U128 (N_128,In_704,In_371);
nor U129 (N_129,In_179,In_1293);
nor U130 (N_130,In_725,In_1020);
and U131 (N_131,In_1479,In_569);
nor U132 (N_132,In_80,In_1286);
xnor U133 (N_133,In_454,In_483);
nor U134 (N_134,In_315,In_873);
or U135 (N_135,In_65,In_343);
or U136 (N_136,In_792,In_647);
nand U137 (N_137,In_883,In_856);
nor U138 (N_138,In_1308,In_1225);
nor U139 (N_139,In_571,In_583);
nor U140 (N_140,In_931,In_861);
nor U141 (N_141,In_499,In_1022);
or U142 (N_142,In_968,In_970);
nand U143 (N_143,In_591,In_720);
nand U144 (N_144,In_213,In_975);
and U145 (N_145,In_206,In_719);
or U146 (N_146,In_769,In_1250);
nand U147 (N_147,In_280,In_162);
or U148 (N_148,In_1218,In_40);
nor U149 (N_149,In_190,In_870);
nor U150 (N_150,In_477,In_147);
nand U151 (N_151,In_729,In_195);
or U152 (N_152,In_13,In_978);
and U153 (N_153,In_967,In_1247);
nand U154 (N_154,In_985,In_687);
and U155 (N_155,In_1167,In_1354);
and U156 (N_156,In_236,In_635);
and U157 (N_157,In_90,In_1154);
nor U158 (N_158,In_640,In_45);
nor U159 (N_159,In_848,In_296);
or U160 (N_160,In_1079,In_370);
nor U161 (N_161,In_381,In_130);
nand U162 (N_162,In_778,In_436);
or U163 (N_163,In_689,In_747);
nor U164 (N_164,In_895,In_932);
or U165 (N_165,In_842,In_20);
nand U166 (N_166,In_545,In_674);
nand U167 (N_167,In_962,In_627);
xor U168 (N_168,In_207,In_1194);
or U169 (N_169,In_1438,In_37);
nand U170 (N_170,In_1116,In_359);
nand U171 (N_171,In_119,In_1422);
nand U172 (N_172,In_749,In_595);
or U173 (N_173,In_32,In_1106);
or U174 (N_174,In_773,In_1336);
or U175 (N_175,In_101,In_418);
or U176 (N_176,In_562,In_1037);
nor U177 (N_177,In_95,In_755);
nand U178 (N_178,In_1050,In_1029);
and U179 (N_179,In_808,In_631);
nor U180 (N_180,In_314,In_15);
or U181 (N_181,In_1107,In_708);
nor U182 (N_182,In_575,In_185);
nor U183 (N_183,In_1091,In_430);
or U184 (N_184,In_1238,In_24);
and U185 (N_185,In_1260,In_1270);
nor U186 (N_186,In_622,In_1367);
nor U187 (N_187,In_9,In_427);
nand U188 (N_188,In_906,In_1254);
nor U189 (N_189,In_536,In_580);
nor U190 (N_190,In_386,In_899);
nand U191 (N_191,In_684,In_825);
and U192 (N_192,In_424,In_7);
nor U193 (N_193,In_661,In_521);
or U194 (N_194,In_1053,In_450);
nor U195 (N_195,In_1162,In_1436);
or U196 (N_196,In_988,In_1026);
nor U197 (N_197,In_639,In_476);
nor U198 (N_198,In_626,In_174);
nor U199 (N_199,In_1421,In_966);
nand U200 (N_200,In_740,In_1410);
and U201 (N_201,In_1121,In_332);
and U202 (N_202,In_209,In_412);
or U203 (N_203,In_1415,In_203);
or U204 (N_204,In_1021,In_972);
or U205 (N_205,In_1307,In_366);
or U206 (N_206,In_608,In_505);
nand U207 (N_207,In_56,In_794);
or U208 (N_208,In_577,In_1492);
or U209 (N_209,In_250,In_1190);
nor U210 (N_210,In_1389,In_892);
xnor U211 (N_211,In_553,In_105);
nand U212 (N_212,In_1387,In_1199);
or U213 (N_213,In_828,In_287);
nor U214 (N_214,In_963,In_682);
nor U215 (N_215,In_413,In_70);
and U216 (N_216,In_256,In_1200);
nor U217 (N_217,In_1015,In_1337);
xnor U218 (N_218,In_573,In_711);
and U219 (N_219,In_217,In_951);
and U220 (N_220,In_558,In_238);
xor U221 (N_221,In_705,In_1092);
or U222 (N_222,In_1396,In_987);
and U223 (N_223,In_1374,In_1297);
nand U224 (N_224,In_1140,In_1301);
or U225 (N_225,In_48,In_880);
and U226 (N_226,In_352,In_544);
and U227 (N_227,In_321,In_937);
or U228 (N_228,In_1085,In_188);
and U229 (N_229,In_913,In_116);
or U230 (N_230,In_677,In_181);
nor U231 (N_231,In_733,In_908);
nor U232 (N_232,In_316,In_59);
or U233 (N_233,In_914,In_1465);
nand U234 (N_234,In_1172,In_425);
nand U235 (N_235,In_304,In_1032);
xnor U236 (N_236,In_1024,In_776);
and U237 (N_237,In_1360,In_1467);
nor U238 (N_238,In_1102,In_87);
nand U239 (N_239,In_994,In_57);
nor U240 (N_240,In_1371,In_533);
and U241 (N_241,In_764,In_262);
or U242 (N_242,In_411,In_1304);
and U243 (N_243,In_319,In_389);
nor U244 (N_244,In_894,In_803);
or U245 (N_245,In_624,In_643);
or U246 (N_246,In_1160,In_486);
nand U247 (N_247,In_301,In_664);
or U248 (N_248,In_1498,In_959);
xor U249 (N_249,In_1111,In_313);
and U250 (N_250,In_1325,In_472);
and U251 (N_251,In_993,In_1314);
nand U252 (N_252,In_983,In_609);
and U253 (N_253,In_1261,In_841);
nand U254 (N_254,In_743,In_761);
nand U255 (N_255,In_1346,In_200);
or U256 (N_256,In_172,In_586);
or U257 (N_257,In_774,In_1138);
nor U258 (N_258,In_33,In_333);
and U259 (N_259,In_194,In_1443);
and U260 (N_260,In_399,In_884);
or U261 (N_261,In_973,In_117);
xnor U262 (N_262,In_220,In_1357);
nor U263 (N_263,In_122,In_1299);
or U264 (N_264,In_1158,In_709);
nor U265 (N_265,In_1391,In_1364);
or U266 (N_266,In_201,In_435);
or U267 (N_267,In_791,In_349);
and U268 (N_268,In_1001,In_662);
nor U269 (N_269,In_1075,In_1497);
and U270 (N_270,In_663,In_878);
or U271 (N_271,In_1406,In_277);
or U272 (N_272,In_796,In_191);
nand U273 (N_273,In_982,In_814);
or U274 (N_274,In_35,In_829);
or U275 (N_275,In_644,In_578);
and U276 (N_276,In_1445,In_341);
and U277 (N_277,In_42,In_1499);
nand U278 (N_278,In_1066,In_1236);
or U279 (N_279,In_1324,In_286);
and U280 (N_280,In_258,In_489);
or U281 (N_281,In_1030,In_1480);
and U282 (N_282,In_568,In_1216);
nand U283 (N_283,In_1191,In_581);
nand U284 (N_284,In_294,In_1223);
and U285 (N_285,In_1446,In_1284);
and U286 (N_286,In_2,In_1493);
and U287 (N_287,In_785,In_990);
and U288 (N_288,In_282,In_126);
nor U289 (N_289,In_713,In_237);
or U290 (N_290,In_109,In_197);
nor U291 (N_291,In_1397,In_945);
or U292 (N_292,In_1186,In_1078);
and U293 (N_293,In_1407,In_34);
nand U294 (N_294,In_1087,In_766);
or U295 (N_295,In_801,In_169);
and U296 (N_296,In_1041,In_317);
nand U297 (N_297,In_283,In_1449);
nand U298 (N_298,In_1474,In_28);
or U299 (N_299,In_1057,In_1274);
or U300 (N_300,In_1128,In_867);
nand U301 (N_301,In_1189,In_1244);
or U302 (N_302,In_673,In_178);
nand U303 (N_303,In_610,In_96);
and U304 (N_304,In_666,In_1237);
nand U305 (N_305,In_155,In_16);
nor U306 (N_306,In_706,In_1188);
nand U307 (N_307,In_741,In_467);
nand U308 (N_308,In_771,In_111);
nand U309 (N_309,In_592,In_1317);
nor U310 (N_310,In_166,In_617);
nand U311 (N_311,In_138,In_927);
or U312 (N_312,In_53,In_1455);
nor U313 (N_313,In_1210,In_183);
nor U314 (N_314,In_1246,In_1413);
and U315 (N_315,In_1313,In_1295);
and U316 (N_316,In_490,In_428);
nand U317 (N_317,In_1209,In_672);
nor U318 (N_318,In_136,In_364);
and U319 (N_319,In_902,In_453);
nand U320 (N_320,In_636,In_1426);
or U321 (N_321,In_930,In_1097);
or U322 (N_322,In_681,In_1036);
or U323 (N_323,In_1441,In_445);
nor U324 (N_324,In_634,In_208);
or U325 (N_325,In_216,In_1203);
nand U326 (N_326,In_1310,In_1207);
nand U327 (N_327,In_1164,In_1255);
and U328 (N_328,In_68,In_896);
nor U329 (N_329,In_1280,In_731);
nand U330 (N_330,In_347,In_1363);
and U331 (N_331,In_531,In_997);
nor U332 (N_332,In_1311,In_175);
or U333 (N_333,In_550,In_941);
or U334 (N_334,In_106,In_465);
nand U335 (N_335,In_605,In_929);
nand U336 (N_336,In_855,In_588);
nand U337 (N_337,In_599,In_695);
and U338 (N_338,In_679,In_851);
and U339 (N_339,In_658,In_368);
nand U340 (N_340,In_1264,In_1148);
xnor U341 (N_341,In_219,In_538);
and U342 (N_342,In_133,In_478);
or U343 (N_343,In_305,In_1204);
or U344 (N_344,In_1320,In_1181);
nand U345 (N_345,In_1228,In_267);
nor U346 (N_346,In_1233,In_89);
or U347 (N_347,In_312,In_1159);
or U348 (N_348,In_613,In_55);
and U349 (N_349,In_1348,In_529);
or U350 (N_350,In_288,In_649);
nor U351 (N_351,In_539,In_1002);
and U352 (N_352,In_239,In_205);
nor U353 (N_353,In_995,In_653);
nand U354 (N_354,In_632,In_1405);
and U355 (N_355,In_405,In_1383);
and U356 (N_356,In_957,In_1385);
xor U357 (N_357,In_1365,In_699);
nor U358 (N_358,In_25,In_215);
and U359 (N_359,In_173,In_812);
nand U360 (N_360,In_722,In_804);
nor U361 (N_361,In_807,In_920);
or U362 (N_362,In_1496,In_877);
and U363 (N_363,In_6,In_285);
nor U364 (N_364,In_1327,In_112);
or U365 (N_365,In_834,In_555);
or U366 (N_366,In_44,In_1151);
and U367 (N_367,In_420,In_1130);
and U368 (N_368,In_1206,In_77);
or U369 (N_369,In_1067,In_923);
nor U370 (N_370,In_844,In_11);
and U371 (N_371,In_735,In_1408);
or U372 (N_372,In_1401,In_1376);
nor U373 (N_373,In_566,In_1283);
and U374 (N_374,In_900,In_149);
nor U375 (N_375,In_1229,In_971);
nand U376 (N_376,In_1031,In_850);
or U377 (N_377,In_1319,In_84);
nor U378 (N_378,In_269,In_58);
xor U379 (N_379,In_103,In_309);
or U380 (N_380,In_86,In_543);
nand U381 (N_381,In_1071,In_452);
nor U382 (N_382,In_819,In_508);
nand U383 (N_383,In_630,In_441);
or U384 (N_384,In_398,In_67);
nand U385 (N_385,In_542,In_152);
xor U386 (N_386,In_1109,In_872);
nor U387 (N_387,In_1012,In_380);
nor U388 (N_388,In_1175,In_1096);
nand U389 (N_389,In_885,In_1252);
nor U390 (N_390,In_1239,In_1146);
or U391 (N_391,In_1155,In_422);
nand U392 (N_392,In_905,In_271);
nor U393 (N_393,In_651,In_176);
nand U394 (N_394,In_437,In_1051);
nand U395 (N_395,In_73,In_164);
nand U396 (N_396,In_1253,In_943);
or U397 (N_397,In_1084,In_1005);
nor U398 (N_398,In_1452,In_680);
nor U399 (N_399,In_1241,In_797);
and U400 (N_400,In_1393,In_97);
nand U401 (N_401,In_1456,In_893);
nand U402 (N_402,In_259,In_1475);
or U403 (N_403,In_298,In_263);
or U404 (N_404,In_43,In_862);
nand U405 (N_405,In_125,In_1040);
and U406 (N_406,In_1326,In_1073);
nor U407 (N_407,In_1420,In_802);
and U408 (N_408,In_548,In_1478);
nand U409 (N_409,In_1076,In_602);
nor U410 (N_410,In_1494,In_1157);
and U411 (N_411,In_1193,In_1485);
nor U412 (N_412,In_1187,In_1461);
nor U413 (N_413,In_308,In_714);
or U414 (N_414,In_510,In_402);
and U415 (N_415,In_820,In_579);
or U416 (N_416,In_401,In_1147);
nand U417 (N_417,In_501,In_324);
nand U418 (N_418,In_1197,In_836);
or U419 (N_419,In_1177,In_1417);
or U420 (N_420,In_1039,In_1259);
or U421 (N_421,In_1129,In_1192);
or U422 (N_422,In_787,In_1350);
nor U423 (N_423,In_93,In_961);
xor U424 (N_424,In_51,In_396);
nand U425 (N_425,In_646,In_1369);
or U426 (N_426,In_1487,In_419);
nand U427 (N_427,In_1144,In_142);
or U428 (N_428,In_1179,In_752);
or U429 (N_429,In_526,In_789);
or U430 (N_430,In_14,In_1099);
and U431 (N_431,In_222,In_1370);
or U432 (N_432,In_915,In_628);
nor U433 (N_433,In_134,In_757);
and U434 (N_434,In_1141,In_940);
or U435 (N_435,In_1089,In_691);
and U436 (N_436,In_1135,In_981);
nor U437 (N_437,In_196,In_443);
nor U438 (N_438,In_1242,In_858);
nand U439 (N_439,In_1352,In_601);
nor U440 (N_440,In_949,In_439);
or U441 (N_441,In_275,In_124);
and U442 (N_442,In_1294,In_415);
or U443 (N_443,In_1333,In_815);
and U444 (N_444,In_956,In_82);
or U445 (N_445,In_1201,In_1439);
and U446 (N_446,In_261,In_504);
nand U447 (N_447,In_1240,In_1305);
nor U448 (N_448,In_1473,In_148);
or U449 (N_449,In_557,In_291);
nand U450 (N_450,In_1090,In_948);
nand U451 (N_451,In_481,In_696);
nor U452 (N_452,In_1234,In_779);
or U453 (N_453,In_1110,In_447);
nand U454 (N_454,In_471,In_167);
or U455 (N_455,In_1048,In_1004);
or U456 (N_456,In_907,In_233);
or U457 (N_457,In_596,In_795);
and U458 (N_458,In_552,In_840);
and U459 (N_459,In_620,In_742);
and U460 (N_460,In_329,In_1378);
nor U461 (N_461,In_473,In_806);
nand U462 (N_462,In_1489,In_1495);
nand U463 (N_463,In_284,In_252);
or U464 (N_464,In_1419,In_1149);
or U465 (N_465,In_1450,In_793);
nand U466 (N_466,In_395,In_657);
nor U467 (N_467,In_676,In_1488);
nand U468 (N_468,In_537,In_19);
nor U469 (N_469,In_350,In_849);
nand U470 (N_470,In_827,In_293);
nor U471 (N_471,In_351,In_522);
nor U472 (N_472,In_335,In_1316);
or U473 (N_473,In_408,In_938);
nor U474 (N_474,In_1086,In_1318);
nor U475 (N_475,In_567,In_830);
or U476 (N_476,In_171,In_433);
nand U477 (N_477,In_0,In_561);
and U478 (N_478,In_273,In_799);
and U479 (N_479,In_274,In_1482);
and U480 (N_480,In_449,In_81);
nand U481 (N_481,In_1454,In_1070);
and U482 (N_482,In_1226,In_1212);
nor U483 (N_483,In_1323,In_1296);
or U484 (N_484,In_598,In_393);
and U485 (N_485,In_564,In_835);
nor U486 (N_486,In_1368,In_1484);
nor U487 (N_487,In_1249,In_912);
nor U488 (N_488,In_41,In_241);
or U489 (N_489,In_1466,In_800);
or U490 (N_490,In_1161,In_414);
or U491 (N_491,In_678,In_254);
nor U492 (N_492,In_272,In_221);
nor U493 (N_493,In_839,In_8);
nand U494 (N_494,In_290,In_1300);
nand U495 (N_495,In_244,In_466);
or U496 (N_496,In_996,In_249);
or U497 (N_497,In_1196,In_1083);
and U498 (N_498,In_600,In_377);
or U499 (N_499,In_1343,In_876);
or U500 (N_500,In_667,In_376);
or U501 (N_501,In_1184,In_790);
nor U502 (N_502,In_3,In_257);
nor U503 (N_503,In_520,In_1014);
or U504 (N_504,In_1347,In_1007);
or U505 (N_505,In_110,In_1412);
nor U506 (N_506,In_302,In_240);
or U507 (N_507,In_514,In_1178);
nand U508 (N_508,In_589,In_346);
and U509 (N_509,In_266,In_768);
nor U510 (N_510,In_404,In_30);
nor U511 (N_511,In_1430,In_833);
or U512 (N_512,In_1463,In_260);
nand U513 (N_513,In_177,In_1108);
nand U514 (N_514,In_1088,In_1195);
nand U515 (N_515,In_223,In_210);
or U516 (N_516,In_765,In_184);
nor U517 (N_517,In_431,In_925);
nor U518 (N_518,In_107,In_1061);
nor U519 (N_519,In_407,In_1425);
nor U520 (N_520,In_491,In_151);
and U521 (N_521,In_39,In_950);
nor U522 (N_522,In_607,In_1150);
nor U523 (N_523,In_120,In_326);
nor U524 (N_524,In_1490,In_1399);
nor U525 (N_525,In_1276,In_123);
and U526 (N_526,In_954,In_365);
or U527 (N_527,In_1006,In_541);
xor U528 (N_528,In_114,In_1345);
and U529 (N_529,In_91,In_1258);
and U530 (N_530,In_307,In_1431);
or U531 (N_531,In_1038,In_462);
xor U532 (N_532,In_1462,In_1054);
nor U533 (N_533,In_1125,In_1119);
or U534 (N_534,In_442,In_247);
or U535 (N_535,In_745,In_1358);
nand U536 (N_536,In_423,In_576);
nor U537 (N_537,In_1414,In_460);
nor U538 (N_538,In_457,In_22);
or U539 (N_539,In_1339,In_549);
and U540 (N_540,In_202,In_686);
nor U541 (N_541,In_330,In_367);
nand U542 (N_542,In_1137,In_204);
or U543 (N_543,In_979,In_1428);
and U544 (N_544,In_1000,In_503);
nor U545 (N_545,In_512,In_952);
and U546 (N_546,In_612,In_255);
nor U547 (N_547,In_253,In_1356);
and U548 (N_548,In_770,In_98);
and U549 (N_549,In_1429,In_1460);
nor U550 (N_550,In_1251,In_234);
nor U551 (N_551,In_1003,In_1103);
or U552 (N_552,In_1098,In_459);
and U553 (N_553,In_629,In_823);
nand U554 (N_554,In_1359,In_671);
and U555 (N_555,In_701,In_52);
nor U556 (N_556,In_383,In_633);
nand U557 (N_557,In_113,In_479);
and U558 (N_558,In_1273,In_1380);
or U559 (N_559,In_597,In_1180);
and U560 (N_560,In_587,In_1065);
nor U561 (N_561,In_942,In_832);
xnor U562 (N_562,In_540,In_150);
and U563 (N_563,In_1282,In_1366);
or U564 (N_564,In_668,In_66);
or U565 (N_565,In_642,In_193);
xor U566 (N_566,In_325,In_158);
xnor U567 (N_567,In_1168,In_660);
or U568 (N_568,In_648,In_163);
or U569 (N_569,In_763,In_340);
nor U570 (N_570,In_918,In_417);
or U571 (N_571,In_604,In_26);
nand U572 (N_572,In_344,In_891);
and U573 (N_573,In_79,In_852);
and U574 (N_574,In_354,In_1133);
nand U575 (N_575,In_859,In_118);
and U576 (N_576,In_392,In_750);
xnor U577 (N_577,In_1321,In_560);
or U578 (N_578,In_903,In_1023);
nand U579 (N_579,In_535,In_1382);
nor U580 (N_580,In_703,In_403);
nor U581 (N_581,In_243,In_463);
or U582 (N_582,In_1335,In_875);
and U583 (N_583,In_1112,In_563);
nor U584 (N_584,In_712,In_369);
and U585 (N_585,In_375,In_1398);
nor U586 (N_586,In_1045,In_698);
or U587 (N_587,In_748,In_297);
and U588 (N_588,In_187,In_339);
or U589 (N_589,In_1451,In_1219);
or U590 (N_590,In_322,In_888);
and U591 (N_591,In_1008,In_410);
nor U592 (N_592,In_715,In_726);
nand U593 (N_593,In_1288,In_1340);
or U594 (N_594,In_69,In_517);
and U595 (N_595,In_1131,In_251);
and U596 (N_596,In_901,In_62);
and U597 (N_597,In_482,In_1101);
nor U598 (N_598,In_159,In_334);
nand U599 (N_599,In_926,In_211);
and U600 (N_600,In_1302,In_670);
and U601 (N_601,In_1245,In_1256);
nor U602 (N_602,In_532,In_104);
nor U603 (N_603,In_1094,In_379);
and U604 (N_604,In_328,In_1136);
or U605 (N_605,In_278,In_1068);
or U606 (N_606,In_928,In_782);
and U607 (N_607,In_358,In_17);
and U608 (N_608,In_99,In_129);
nand U609 (N_609,In_1034,In_1440);
and U610 (N_610,In_718,In_960);
and U611 (N_611,In_1315,In_498);
nor U612 (N_612,In_485,In_989);
or U613 (N_613,In_300,In_224);
or U614 (N_614,In_78,In_525);
nand U615 (N_615,In_180,In_818);
or U616 (N_616,In_1424,In_182);
and U617 (N_617,In_488,In_519);
nor U618 (N_618,In_1114,In_805);
or U619 (N_619,In_1183,In_882);
nand U620 (N_620,In_1329,In_444);
or U621 (N_621,In_621,In_121);
nand U622 (N_622,In_1142,In_140);
or U623 (N_623,In_1458,In_523);
or U624 (N_624,In_1049,In_1491);
nand U625 (N_625,In_1468,In_511);
nand U626 (N_626,In_1,In_977);
or U627 (N_627,In_721,In_1132);
nor U628 (N_628,In_1232,In_953);
nor U629 (N_629,In_1198,In_1126);
nor U630 (N_630,In_391,In_497);
nor U631 (N_631,In_1060,In_656);
nand U632 (N_632,In_1222,In_853);
or U633 (N_633,In_665,In_1469);
and U634 (N_634,In_738,In_299);
and U635 (N_635,In_1402,In_1269);
nand U636 (N_636,In_141,In_1486);
nand U637 (N_637,In_21,In_1010);
or U638 (N_638,In_619,In_1211);
or U639 (N_639,In_527,In_737);
nor U640 (N_640,In_323,In_1483);
nand U641 (N_641,In_1289,In_1384);
xnor U642 (N_642,In_102,In_675);
nor U643 (N_643,In_338,In_320);
nand U644 (N_644,In_570,In_145);
nand U645 (N_645,In_1176,In_394);
and U646 (N_646,In_74,In_27);
nor U647 (N_647,In_456,In_1163);
or U648 (N_648,In_860,In_1042);
nor U649 (N_649,In_736,In_924);
or U650 (N_650,In_342,In_1080);
nor U651 (N_651,In_1081,In_461);
and U652 (N_652,In_1170,In_1143);
and U653 (N_653,In_585,In_1156);
or U654 (N_654,In_1444,In_1266);
and U655 (N_655,In_732,In_998);
nand U656 (N_656,In_683,In_946);
nor U657 (N_657,In_265,In_874);
and U658 (N_658,In_1292,In_964);
or U659 (N_659,In_1312,In_143);
and U660 (N_660,In_1353,In_1074);
or U661 (N_661,In_1059,In_565);
or U662 (N_662,In_798,In_1213);
and U663 (N_663,In_739,In_1435);
or U664 (N_664,In_710,In_1372);
or U665 (N_665,In_1448,In_1165);
or U666 (N_666,In_1214,In_934);
or U667 (N_667,In_416,In_470);
or U668 (N_668,In_1095,In_865);
nor U669 (N_669,In_373,In_440);
nand U670 (N_670,In_1403,In_922);
nor U671 (N_671,In_357,In_824);
and U672 (N_672,In_1375,In_1139);
or U673 (N_673,In_615,In_432);
nor U674 (N_674,In_46,In_100);
and U675 (N_675,In_235,In_574);
nand U676 (N_676,In_108,In_1153);
or U677 (N_677,In_397,In_94);
nand U678 (N_678,In_1230,In_387);
nand U679 (N_679,In_593,In_474);
and U680 (N_680,In_904,In_616);
nor U681 (N_681,In_1205,In_991);
nand U682 (N_682,In_916,In_18);
and U683 (N_683,In_60,In_388);
or U684 (N_684,In_1349,In_817);
nand U685 (N_685,In_584,In_1338);
nand U686 (N_686,In_958,In_910);
or U687 (N_687,In_4,In_362);
nand U688 (N_688,In_214,In_980);
and U689 (N_689,In_746,In_976);
nand U690 (N_690,In_1427,In_772);
nand U691 (N_691,In_1100,In_1442);
or U692 (N_692,In_1248,In_965);
and U693 (N_693,In_871,In_336);
and U694 (N_694,In_760,In_1331);
and U695 (N_695,In_1285,In_1231);
nor U696 (N_696,In_372,In_1058);
nor U697 (N_697,In_469,In_1117);
and U698 (N_698,In_692,In_318);
and U699 (N_699,In_331,In_458);
nand U700 (N_700,In_500,In_1019);
nor U701 (N_701,In_887,In_270);
nand U702 (N_702,In_821,In_455);
nand U703 (N_703,In_1457,In_1279);
or U704 (N_704,In_641,In_1047);
and U705 (N_705,In_702,In_780);
nor U706 (N_706,In_160,In_292);
or U707 (N_707,In_231,In_228);
nor U708 (N_708,In_1409,In_759);
or U709 (N_709,In_1063,In_1082);
and U710 (N_710,In_1174,In_1464);
and U711 (N_711,In_1471,In_327);
nor U712 (N_712,In_898,In_694);
or U713 (N_713,In_1118,In_502);
nand U714 (N_714,In_1093,In_127);
nor U715 (N_715,In_518,In_1182);
and U716 (N_716,In_135,In_984);
xor U717 (N_717,In_361,In_218);
nand U718 (N_718,In_1016,In_227);
and U719 (N_719,In_385,In_826);
and U720 (N_720,In_869,In_225);
and U721 (N_721,In_1169,In_1281);
or U722 (N_722,In_1433,In_506);
nand U723 (N_723,In_337,In_936);
or U724 (N_724,In_1411,In_728);
or U725 (N_725,In_5,In_767);
and U726 (N_726,In_843,In_831);
or U727 (N_727,In_655,In_1077);
nor U728 (N_728,In_868,In_786);
nand U729 (N_729,In_1221,In_1332);
xnor U730 (N_730,In_1202,In_762);
or U731 (N_731,In_1145,In_137);
nor U732 (N_732,In_289,In_186);
nand U733 (N_733,In_1124,In_232);
or U734 (N_734,In_72,In_279);
or U735 (N_735,In_360,In_582);
and U736 (N_736,In_1400,In_1334);
and U737 (N_737,In_700,In_813);
or U738 (N_738,In_614,In_939);
nand U739 (N_739,In_509,In_1257);
or U740 (N_740,In_1044,In_246);
nand U741 (N_741,In_1235,In_756);
nor U742 (N_742,In_837,In_295);
and U743 (N_743,In_36,In_199);
nor U744 (N_744,In_723,In_1035);
nand U745 (N_745,In_935,In_783);
nand U746 (N_746,In_1017,In_611);
nand U747 (N_747,In_356,In_513);
nand U748 (N_748,In_1265,In_889);
and U749 (N_749,In_1127,In_784);
nor U750 (N_750,In_1172,In_1416);
nor U751 (N_751,In_196,In_1130);
xnor U752 (N_752,In_500,In_662);
nand U753 (N_753,In_1401,In_524);
nor U754 (N_754,In_1224,In_258);
and U755 (N_755,In_569,In_1363);
or U756 (N_756,In_186,In_1335);
nor U757 (N_757,In_798,In_481);
nand U758 (N_758,In_389,In_1495);
nand U759 (N_759,In_677,In_531);
nor U760 (N_760,In_169,In_126);
nor U761 (N_761,In_1237,In_908);
nor U762 (N_762,In_564,In_458);
nand U763 (N_763,In_48,In_1110);
nor U764 (N_764,In_484,In_1031);
or U765 (N_765,In_647,In_491);
or U766 (N_766,In_310,In_176);
and U767 (N_767,In_1479,In_255);
nand U768 (N_768,In_1356,In_1230);
or U769 (N_769,In_815,In_966);
nand U770 (N_770,In_1218,In_218);
nand U771 (N_771,In_592,In_873);
nor U772 (N_772,In_685,In_579);
and U773 (N_773,In_952,In_311);
nor U774 (N_774,In_318,In_862);
or U775 (N_775,In_706,In_1304);
and U776 (N_776,In_844,In_71);
or U777 (N_777,In_353,In_1479);
and U778 (N_778,In_565,In_433);
or U779 (N_779,In_714,In_1171);
nand U780 (N_780,In_343,In_1175);
nor U781 (N_781,In_286,In_40);
or U782 (N_782,In_1417,In_535);
or U783 (N_783,In_1469,In_62);
nor U784 (N_784,In_24,In_433);
and U785 (N_785,In_927,In_57);
nor U786 (N_786,In_874,In_1375);
and U787 (N_787,In_1236,In_1311);
and U788 (N_788,In_1443,In_922);
or U789 (N_789,In_1496,In_883);
nor U790 (N_790,In_787,In_1247);
and U791 (N_791,In_101,In_1210);
nor U792 (N_792,In_669,In_1047);
nand U793 (N_793,In_1493,In_1137);
nand U794 (N_794,In_152,In_659);
and U795 (N_795,In_1196,In_638);
and U796 (N_796,In_1493,In_1167);
and U797 (N_797,In_1320,In_120);
xnor U798 (N_798,In_79,In_584);
nor U799 (N_799,In_0,In_613);
and U800 (N_800,In_1045,In_1334);
xnor U801 (N_801,In_194,In_634);
xnor U802 (N_802,In_1435,In_505);
nor U803 (N_803,In_1197,In_1360);
xor U804 (N_804,In_1144,In_156);
or U805 (N_805,In_1117,In_1156);
nand U806 (N_806,In_684,In_286);
and U807 (N_807,In_630,In_240);
nand U808 (N_808,In_309,In_1201);
or U809 (N_809,In_423,In_1349);
and U810 (N_810,In_395,In_1121);
or U811 (N_811,In_812,In_341);
nand U812 (N_812,In_423,In_1281);
or U813 (N_813,In_237,In_1003);
nor U814 (N_814,In_837,In_505);
or U815 (N_815,In_1123,In_1132);
xor U816 (N_816,In_1457,In_365);
or U817 (N_817,In_156,In_281);
and U818 (N_818,In_14,In_490);
nand U819 (N_819,In_1096,In_83);
or U820 (N_820,In_788,In_98);
and U821 (N_821,In_53,In_377);
or U822 (N_822,In_471,In_1229);
xor U823 (N_823,In_708,In_115);
and U824 (N_824,In_1079,In_760);
or U825 (N_825,In_27,In_1352);
nand U826 (N_826,In_406,In_1271);
or U827 (N_827,In_1444,In_478);
nor U828 (N_828,In_1450,In_1242);
and U829 (N_829,In_347,In_49);
nand U830 (N_830,In_1059,In_845);
nor U831 (N_831,In_1092,In_425);
or U832 (N_832,In_1056,In_206);
or U833 (N_833,In_481,In_765);
nor U834 (N_834,In_1198,In_909);
and U835 (N_835,In_357,In_1353);
nor U836 (N_836,In_1409,In_83);
or U837 (N_837,In_451,In_794);
and U838 (N_838,In_1481,In_548);
nand U839 (N_839,In_32,In_1321);
nand U840 (N_840,In_305,In_1322);
and U841 (N_841,In_533,In_1129);
nand U842 (N_842,In_321,In_1014);
or U843 (N_843,In_537,In_796);
and U844 (N_844,In_436,In_201);
and U845 (N_845,In_1158,In_1182);
nand U846 (N_846,In_1230,In_494);
and U847 (N_847,In_1022,In_341);
nand U848 (N_848,In_1411,In_1369);
nor U849 (N_849,In_132,In_1160);
and U850 (N_850,In_268,In_257);
nand U851 (N_851,In_1039,In_431);
nor U852 (N_852,In_1223,In_1422);
nand U853 (N_853,In_205,In_1077);
nor U854 (N_854,In_1025,In_183);
nand U855 (N_855,In_974,In_1104);
nand U856 (N_856,In_512,In_659);
nor U857 (N_857,In_611,In_1375);
and U858 (N_858,In_33,In_1150);
and U859 (N_859,In_791,In_1399);
nand U860 (N_860,In_548,In_460);
and U861 (N_861,In_909,In_1459);
and U862 (N_862,In_299,In_614);
and U863 (N_863,In_517,In_426);
or U864 (N_864,In_986,In_1364);
or U865 (N_865,In_1305,In_473);
nor U866 (N_866,In_44,In_157);
or U867 (N_867,In_266,In_1429);
nor U868 (N_868,In_561,In_93);
and U869 (N_869,In_1211,In_449);
and U870 (N_870,In_1032,In_1011);
and U871 (N_871,In_1451,In_1311);
or U872 (N_872,In_1031,In_1211);
or U873 (N_873,In_932,In_600);
nand U874 (N_874,In_1461,In_551);
or U875 (N_875,In_86,In_1357);
or U876 (N_876,In_1312,In_817);
or U877 (N_877,In_1099,In_332);
and U878 (N_878,In_1162,In_434);
or U879 (N_879,In_248,In_744);
nor U880 (N_880,In_449,In_477);
and U881 (N_881,In_559,In_75);
or U882 (N_882,In_470,In_944);
nand U883 (N_883,In_975,In_501);
or U884 (N_884,In_1010,In_859);
and U885 (N_885,In_275,In_1049);
and U886 (N_886,In_866,In_1294);
or U887 (N_887,In_131,In_912);
or U888 (N_888,In_681,In_533);
or U889 (N_889,In_673,In_1491);
and U890 (N_890,In_9,In_223);
or U891 (N_891,In_603,In_533);
and U892 (N_892,In_1188,In_955);
nor U893 (N_893,In_1125,In_1366);
nor U894 (N_894,In_784,In_839);
or U895 (N_895,In_205,In_519);
nor U896 (N_896,In_155,In_1016);
or U897 (N_897,In_276,In_58);
or U898 (N_898,In_1027,In_444);
nand U899 (N_899,In_1389,In_865);
and U900 (N_900,In_182,In_1320);
nand U901 (N_901,In_1244,In_703);
or U902 (N_902,In_114,In_71);
or U903 (N_903,In_125,In_996);
and U904 (N_904,In_1183,In_1284);
or U905 (N_905,In_982,In_1470);
nor U906 (N_906,In_334,In_340);
or U907 (N_907,In_763,In_625);
and U908 (N_908,In_1269,In_1192);
nor U909 (N_909,In_400,In_744);
or U910 (N_910,In_852,In_913);
nand U911 (N_911,In_1097,In_278);
and U912 (N_912,In_23,In_445);
nor U913 (N_913,In_1301,In_1059);
or U914 (N_914,In_1170,In_920);
nor U915 (N_915,In_1310,In_809);
nor U916 (N_916,In_188,In_1131);
and U917 (N_917,In_1140,In_1482);
nand U918 (N_918,In_881,In_925);
and U919 (N_919,In_1345,In_1135);
and U920 (N_920,In_249,In_985);
nand U921 (N_921,In_990,In_999);
or U922 (N_922,In_1404,In_306);
and U923 (N_923,In_733,In_1458);
or U924 (N_924,In_862,In_256);
or U925 (N_925,In_461,In_793);
nand U926 (N_926,In_972,In_1181);
nor U927 (N_927,In_549,In_978);
and U928 (N_928,In_207,In_107);
nor U929 (N_929,In_556,In_1259);
and U930 (N_930,In_1121,In_188);
nor U931 (N_931,In_104,In_880);
nor U932 (N_932,In_1490,In_93);
nor U933 (N_933,In_1202,In_1241);
and U934 (N_934,In_889,In_497);
and U935 (N_935,In_333,In_355);
or U936 (N_936,In_421,In_1433);
and U937 (N_937,In_250,In_1217);
nor U938 (N_938,In_1439,In_146);
nor U939 (N_939,In_681,In_904);
nand U940 (N_940,In_20,In_289);
nand U941 (N_941,In_621,In_136);
nor U942 (N_942,In_839,In_1003);
nand U943 (N_943,In_1103,In_1366);
or U944 (N_944,In_1204,In_21);
xnor U945 (N_945,In_10,In_238);
nand U946 (N_946,In_1244,In_556);
or U947 (N_947,In_232,In_583);
nand U948 (N_948,In_488,In_895);
and U949 (N_949,In_566,In_931);
and U950 (N_950,In_117,In_765);
or U951 (N_951,In_278,In_1177);
nand U952 (N_952,In_1258,In_959);
nand U953 (N_953,In_1458,In_464);
nand U954 (N_954,In_1399,In_974);
nor U955 (N_955,In_117,In_1413);
and U956 (N_956,In_244,In_601);
nor U957 (N_957,In_703,In_34);
nand U958 (N_958,In_1028,In_1478);
nor U959 (N_959,In_762,In_259);
nor U960 (N_960,In_1406,In_1354);
or U961 (N_961,In_776,In_386);
nand U962 (N_962,In_1254,In_216);
and U963 (N_963,In_892,In_1117);
or U964 (N_964,In_889,In_1398);
nor U965 (N_965,In_537,In_1020);
nor U966 (N_966,In_644,In_1395);
nor U967 (N_967,In_550,In_1220);
and U968 (N_968,In_1106,In_234);
or U969 (N_969,In_1212,In_1166);
xnor U970 (N_970,In_434,In_1079);
nand U971 (N_971,In_814,In_1359);
nand U972 (N_972,In_283,In_911);
or U973 (N_973,In_78,In_634);
or U974 (N_974,In_158,In_910);
nor U975 (N_975,In_971,In_751);
or U976 (N_976,In_794,In_428);
nor U977 (N_977,In_1294,In_265);
nor U978 (N_978,In_494,In_101);
nand U979 (N_979,In_945,In_30);
nor U980 (N_980,In_264,In_1298);
xnor U981 (N_981,In_216,In_896);
nor U982 (N_982,In_1437,In_455);
nand U983 (N_983,In_272,In_1163);
or U984 (N_984,In_638,In_82);
or U985 (N_985,In_283,In_443);
nand U986 (N_986,In_505,In_1071);
and U987 (N_987,In_564,In_342);
and U988 (N_988,In_787,In_1172);
or U989 (N_989,In_356,In_302);
nand U990 (N_990,In_584,In_883);
nor U991 (N_991,In_314,In_1297);
or U992 (N_992,In_1379,In_503);
or U993 (N_993,In_1453,In_459);
and U994 (N_994,In_534,In_850);
and U995 (N_995,In_1269,In_1479);
and U996 (N_996,In_1421,In_775);
nor U997 (N_997,In_350,In_1326);
nor U998 (N_998,In_781,In_879);
nand U999 (N_999,In_601,In_1295);
nor U1000 (N_1000,In_1284,In_1219);
or U1001 (N_1001,In_368,In_14);
and U1002 (N_1002,In_1116,In_1293);
nor U1003 (N_1003,In_778,In_1129);
and U1004 (N_1004,In_348,In_938);
nand U1005 (N_1005,In_1383,In_373);
or U1006 (N_1006,In_1443,In_1296);
and U1007 (N_1007,In_794,In_1447);
nor U1008 (N_1008,In_1434,In_381);
nor U1009 (N_1009,In_36,In_367);
or U1010 (N_1010,In_1000,In_105);
nand U1011 (N_1011,In_730,In_524);
and U1012 (N_1012,In_977,In_191);
and U1013 (N_1013,In_813,In_344);
nor U1014 (N_1014,In_1118,In_220);
and U1015 (N_1015,In_319,In_979);
and U1016 (N_1016,In_318,In_854);
nor U1017 (N_1017,In_700,In_1268);
or U1018 (N_1018,In_178,In_165);
or U1019 (N_1019,In_1279,In_767);
and U1020 (N_1020,In_1033,In_1067);
nand U1021 (N_1021,In_904,In_536);
or U1022 (N_1022,In_1355,In_1441);
nand U1023 (N_1023,In_1149,In_973);
nand U1024 (N_1024,In_1068,In_346);
or U1025 (N_1025,In_1131,In_1040);
nor U1026 (N_1026,In_902,In_747);
nor U1027 (N_1027,In_307,In_288);
nand U1028 (N_1028,In_646,In_872);
or U1029 (N_1029,In_827,In_780);
and U1030 (N_1030,In_432,In_123);
nand U1031 (N_1031,In_1207,In_1343);
nor U1032 (N_1032,In_237,In_692);
nand U1033 (N_1033,In_721,In_889);
or U1034 (N_1034,In_1156,In_1148);
nand U1035 (N_1035,In_428,In_926);
nand U1036 (N_1036,In_1364,In_1431);
nand U1037 (N_1037,In_1181,In_1485);
or U1038 (N_1038,In_149,In_1024);
nor U1039 (N_1039,In_558,In_232);
xnor U1040 (N_1040,In_256,In_183);
and U1041 (N_1041,In_237,In_814);
nor U1042 (N_1042,In_739,In_1488);
nor U1043 (N_1043,In_711,In_78);
nand U1044 (N_1044,In_78,In_1166);
nand U1045 (N_1045,In_6,In_1227);
and U1046 (N_1046,In_10,In_97);
nand U1047 (N_1047,In_777,In_1113);
nand U1048 (N_1048,In_1240,In_1245);
nor U1049 (N_1049,In_802,In_1064);
and U1050 (N_1050,In_769,In_767);
or U1051 (N_1051,In_27,In_710);
nor U1052 (N_1052,In_224,In_1220);
and U1053 (N_1053,In_311,In_1303);
nor U1054 (N_1054,In_1037,In_716);
nand U1055 (N_1055,In_288,In_550);
nor U1056 (N_1056,In_1295,In_322);
or U1057 (N_1057,In_828,In_1082);
nor U1058 (N_1058,In_1481,In_1103);
nor U1059 (N_1059,In_134,In_1494);
and U1060 (N_1060,In_413,In_539);
nor U1061 (N_1061,In_1096,In_197);
or U1062 (N_1062,In_997,In_263);
nor U1063 (N_1063,In_1023,In_1156);
or U1064 (N_1064,In_669,In_226);
nand U1065 (N_1065,In_375,In_596);
nand U1066 (N_1066,In_1153,In_880);
nor U1067 (N_1067,In_1074,In_60);
nor U1068 (N_1068,In_1100,In_716);
and U1069 (N_1069,In_142,In_897);
and U1070 (N_1070,In_1113,In_1177);
nor U1071 (N_1071,In_445,In_1277);
nor U1072 (N_1072,In_563,In_143);
nand U1073 (N_1073,In_646,In_812);
nor U1074 (N_1074,In_259,In_324);
nand U1075 (N_1075,In_1195,In_30);
and U1076 (N_1076,In_445,In_785);
nor U1077 (N_1077,In_822,In_452);
and U1078 (N_1078,In_1026,In_131);
nand U1079 (N_1079,In_277,In_302);
nand U1080 (N_1080,In_257,In_375);
nand U1081 (N_1081,In_1328,In_1435);
and U1082 (N_1082,In_1186,In_276);
nor U1083 (N_1083,In_1200,In_1115);
nand U1084 (N_1084,In_118,In_1216);
nor U1085 (N_1085,In_760,In_309);
or U1086 (N_1086,In_1442,In_1475);
nand U1087 (N_1087,In_202,In_69);
nor U1088 (N_1088,In_1366,In_631);
nor U1089 (N_1089,In_56,In_1426);
xor U1090 (N_1090,In_1017,In_1499);
or U1091 (N_1091,In_482,In_334);
xor U1092 (N_1092,In_147,In_785);
nor U1093 (N_1093,In_1043,In_1384);
nor U1094 (N_1094,In_1087,In_761);
or U1095 (N_1095,In_446,In_1445);
or U1096 (N_1096,In_967,In_611);
nor U1097 (N_1097,In_383,In_564);
and U1098 (N_1098,In_1120,In_167);
xnor U1099 (N_1099,In_158,In_6);
and U1100 (N_1100,In_1080,In_1271);
or U1101 (N_1101,In_609,In_807);
or U1102 (N_1102,In_906,In_220);
nand U1103 (N_1103,In_173,In_108);
nand U1104 (N_1104,In_997,In_929);
or U1105 (N_1105,In_804,In_1489);
nand U1106 (N_1106,In_1164,In_685);
nor U1107 (N_1107,In_1339,In_222);
or U1108 (N_1108,In_1430,In_810);
nor U1109 (N_1109,In_282,In_1068);
nand U1110 (N_1110,In_1356,In_1413);
nor U1111 (N_1111,In_129,In_862);
and U1112 (N_1112,In_81,In_956);
nor U1113 (N_1113,In_1309,In_151);
and U1114 (N_1114,In_685,In_420);
nor U1115 (N_1115,In_1378,In_1230);
and U1116 (N_1116,In_575,In_1098);
xnor U1117 (N_1117,In_1489,In_1001);
and U1118 (N_1118,In_566,In_898);
nand U1119 (N_1119,In_303,In_1091);
nand U1120 (N_1120,In_638,In_1146);
or U1121 (N_1121,In_885,In_791);
nand U1122 (N_1122,In_586,In_981);
nor U1123 (N_1123,In_666,In_1090);
and U1124 (N_1124,In_745,In_406);
nor U1125 (N_1125,In_503,In_368);
nor U1126 (N_1126,In_1388,In_1413);
xnor U1127 (N_1127,In_1443,In_186);
nor U1128 (N_1128,In_786,In_764);
and U1129 (N_1129,In_1151,In_286);
or U1130 (N_1130,In_1079,In_533);
nand U1131 (N_1131,In_643,In_78);
nand U1132 (N_1132,In_1387,In_328);
nor U1133 (N_1133,In_107,In_1120);
nand U1134 (N_1134,In_725,In_1169);
or U1135 (N_1135,In_1258,In_565);
and U1136 (N_1136,In_654,In_1428);
nor U1137 (N_1137,In_14,In_249);
nor U1138 (N_1138,In_1258,In_1182);
or U1139 (N_1139,In_855,In_445);
or U1140 (N_1140,In_1277,In_795);
or U1141 (N_1141,In_210,In_430);
nand U1142 (N_1142,In_1238,In_832);
or U1143 (N_1143,In_965,In_378);
and U1144 (N_1144,In_1339,In_1332);
and U1145 (N_1145,In_33,In_437);
nor U1146 (N_1146,In_245,In_927);
or U1147 (N_1147,In_1104,In_1024);
and U1148 (N_1148,In_1051,In_1367);
nand U1149 (N_1149,In_231,In_1028);
nor U1150 (N_1150,In_1082,In_580);
nand U1151 (N_1151,In_1003,In_868);
and U1152 (N_1152,In_591,In_1101);
or U1153 (N_1153,In_484,In_1427);
xnor U1154 (N_1154,In_4,In_152);
or U1155 (N_1155,In_1463,In_943);
or U1156 (N_1156,In_723,In_307);
nor U1157 (N_1157,In_102,In_1485);
nand U1158 (N_1158,In_666,In_1344);
and U1159 (N_1159,In_996,In_910);
or U1160 (N_1160,In_297,In_212);
nand U1161 (N_1161,In_746,In_563);
nor U1162 (N_1162,In_479,In_23);
nor U1163 (N_1163,In_215,In_28);
nor U1164 (N_1164,In_1196,In_1067);
nor U1165 (N_1165,In_1180,In_608);
or U1166 (N_1166,In_586,In_227);
nor U1167 (N_1167,In_922,In_404);
or U1168 (N_1168,In_845,In_283);
or U1169 (N_1169,In_456,In_733);
nor U1170 (N_1170,In_945,In_60);
and U1171 (N_1171,In_844,In_148);
nand U1172 (N_1172,In_1454,In_707);
nand U1173 (N_1173,In_1123,In_1205);
and U1174 (N_1174,In_841,In_248);
or U1175 (N_1175,In_1126,In_466);
nand U1176 (N_1176,In_457,In_185);
or U1177 (N_1177,In_1217,In_61);
nor U1178 (N_1178,In_314,In_628);
nor U1179 (N_1179,In_160,In_1077);
and U1180 (N_1180,In_1278,In_864);
and U1181 (N_1181,In_1230,In_26);
and U1182 (N_1182,In_363,In_7);
and U1183 (N_1183,In_650,In_333);
xnor U1184 (N_1184,In_1473,In_1496);
nor U1185 (N_1185,In_1489,In_419);
or U1186 (N_1186,In_1373,In_5);
or U1187 (N_1187,In_84,In_11);
and U1188 (N_1188,In_866,In_1488);
xnor U1189 (N_1189,In_562,In_1250);
nand U1190 (N_1190,In_205,In_367);
nand U1191 (N_1191,In_1103,In_369);
and U1192 (N_1192,In_541,In_523);
nor U1193 (N_1193,In_650,In_1331);
nor U1194 (N_1194,In_969,In_390);
or U1195 (N_1195,In_905,In_1192);
nand U1196 (N_1196,In_111,In_774);
or U1197 (N_1197,In_1499,In_115);
nor U1198 (N_1198,In_791,In_1403);
and U1199 (N_1199,In_85,In_1152);
nand U1200 (N_1200,In_316,In_82);
and U1201 (N_1201,In_1306,In_1434);
and U1202 (N_1202,In_124,In_645);
nand U1203 (N_1203,In_1478,In_434);
or U1204 (N_1204,In_674,In_1319);
nand U1205 (N_1205,In_942,In_1159);
nand U1206 (N_1206,In_1151,In_565);
and U1207 (N_1207,In_1352,In_473);
or U1208 (N_1208,In_546,In_893);
or U1209 (N_1209,In_314,In_1322);
or U1210 (N_1210,In_959,In_475);
and U1211 (N_1211,In_647,In_1104);
nand U1212 (N_1212,In_1039,In_1005);
and U1213 (N_1213,In_784,In_542);
nor U1214 (N_1214,In_281,In_1111);
or U1215 (N_1215,In_633,In_697);
nand U1216 (N_1216,In_1153,In_98);
and U1217 (N_1217,In_1119,In_345);
and U1218 (N_1218,In_701,In_99);
or U1219 (N_1219,In_1447,In_179);
or U1220 (N_1220,In_766,In_914);
and U1221 (N_1221,In_449,In_155);
nor U1222 (N_1222,In_1027,In_1217);
or U1223 (N_1223,In_956,In_1370);
and U1224 (N_1224,In_257,In_816);
and U1225 (N_1225,In_1329,In_1305);
nor U1226 (N_1226,In_444,In_832);
and U1227 (N_1227,In_1451,In_510);
or U1228 (N_1228,In_1035,In_1063);
and U1229 (N_1229,In_427,In_1059);
nor U1230 (N_1230,In_1205,In_1016);
nor U1231 (N_1231,In_575,In_673);
and U1232 (N_1232,In_202,In_453);
nand U1233 (N_1233,In_1457,In_1405);
or U1234 (N_1234,In_1250,In_263);
nand U1235 (N_1235,In_395,In_1273);
nor U1236 (N_1236,In_168,In_1452);
or U1237 (N_1237,In_696,In_547);
and U1238 (N_1238,In_535,In_144);
nand U1239 (N_1239,In_905,In_1010);
and U1240 (N_1240,In_952,In_1372);
nand U1241 (N_1241,In_1491,In_433);
or U1242 (N_1242,In_487,In_1407);
nor U1243 (N_1243,In_751,In_2);
or U1244 (N_1244,In_953,In_222);
and U1245 (N_1245,In_115,In_730);
and U1246 (N_1246,In_1012,In_274);
and U1247 (N_1247,In_1397,In_275);
nand U1248 (N_1248,In_1476,In_1412);
nand U1249 (N_1249,In_990,In_1483);
nor U1250 (N_1250,In_416,In_1246);
and U1251 (N_1251,In_697,In_1346);
and U1252 (N_1252,In_876,In_632);
nor U1253 (N_1253,In_863,In_608);
or U1254 (N_1254,In_685,In_845);
or U1255 (N_1255,In_562,In_1170);
and U1256 (N_1256,In_694,In_84);
nor U1257 (N_1257,In_322,In_645);
nand U1258 (N_1258,In_803,In_964);
and U1259 (N_1259,In_1198,In_26);
nand U1260 (N_1260,In_964,In_540);
or U1261 (N_1261,In_387,In_415);
or U1262 (N_1262,In_1045,In_775);
nand U1263 (N_1263,In_676,In_563);
nor U1264 (N_1264,In_1199,In_352);
or U1265 (N_1265,In_931,In_196);
or U1266 (N_1266,In_32,In_394);
nand U1267 (N_1267,In_277,In_881);
or U1268 (N_1268,In_924,In_1053);
nand U1269 (N_1269,In_190,In_1053);
or U1270 (N_1270,In_649,In_264);
or U1271 (N_1271,In_514,In_1061);
nor U1272 (N_1272,In_1235,In_987);
nor U1273 (N_1273,In_1467,In_1127);
nand U1274 (N_1274,In_1172,In_202);
or U1275 (N_1275,In_983,In_224);
nor U1276 (N_1276,In_848,In_1371);
or U1277 (N_1277,In_1168,In_1491);
nand U1278 (N_1278,In_387,In_109);
nor U1279 (N_1279,In_11,In_1350);
nor U1280 (N_1280,In_988,In_345);
nor U1281 (N_1281,In_73,In_50);
or U1282 (N_1282,In_544,In_448);
nand U1283 (N_1283,In_433,In_1422);
or U1284 (N_1284,In_163,In_1425);
and U1285 (N_1285,In_1406,In_875);
or U1286 (N_1286,In_267,In_607);
nor U1287 (N_1287,In_460,In_517);
and U1288 (N_1288,In_63,In_1111);
and U1289 (N_1289,In_487,In_827);
and U1290 (N_1290,In_96,In_6);
nand U1291 (N_1291,In_294,In_714);
xor U1292 (N_1292,In_1153,In_99);
and U1293 (N_1293,In_1340,In_479);
nor U1294 (N_1294,In_694,In_57);
or U1295 (N_1295,In_643,In_889);
and U1296 (N_1296,In_761,In_1094);
and U1297 (N_1297,In_1281,In_1007);
and U1298 (N_1298,In_1357,In_475);
nor U1299 (N_1299,In_452,In_1105);
nor U1300 (N_1300,In_174,In_343);
and U1301 (N_1301,In_903,In_1001);
or U1302 (N_1302,In_622,In_177);
and U1303 (N_1303,In_200,In_1205);
or U1304 (N_1304,In_824,In_606);
nand U1305 (N_1305,In_1404,In_662);
or U1306 (N_1306,In_1457,In_81);
or U1307 (N_1307,In_344,In_769);
nand U1308 (N_1308,In_200,In_214);
or U1309 (N_1309,In_567,In_117);
and U1310 (N_1310,In_731,In_170);
and U1311 (N_1311,In_632,In_341);
or U1312 (N_1312,In_809,In_355);
nand U1313 (N_1313,In_83,In_405);
and U1314 (N_1314,In_965,In_1455);
and U1315 (N_1315,In_667,In_502);
and U1316 (N_1316,In_491,In_756);
nor U1317 (N_1317,In_993,In_1224);
xor U1318 (N_1318,In_135,In_657);
nand U1319 (N_1319,In_705,In_1478);
and U1320 (N_1320,In_694,In_203);
and U1321 (N_1321,In_1244,In_207);
and U1322 (N_1322,In_506,In_766);
nand U1323 (N_1323,In_814,In_1196);
and U1324 (N_1324,In_608,In_1431);
nor U1325 (N_1325,In_553,In_318);
nand U1326 (N_1326,In_526,In_536);
nor U1327 (N_1327,In_1212,In_912);
nand U1328 (N_1328,In_776,In_49);
or U1329 (N_1329,In_287,In_293);
or U1330 (N_1330,In_386,In_53);
nand U1331 (N_1331,In_1309,In_166);
nand U1332 (N_1332,In_604,In_581);
and U1333 (N_1333,In_163,In_443);
or U1334 (N_1334,In_411,In_715);
nor U1335 (N_1335,In_364,In_902);
nor U1336 (N_1336,In_544,In_939);
nand U1337 (N_1337,In_857,In_513);
and U1338 (N_1338,In_1458,In_1436);
nor U1339 (N_1339,In_1233,In_196);
nor U1340 (N_1340,In_174,In_1132);
or U1341 (N_1341,In_1087,In_376);
and U1342 (N_1342,In_1325,In_945);
nand U1343 (N_1343,In_758,In_1377);
and U1344 (N_1344,In_940,In_351);
nand U1345 (N_1345,In_685,In_317);
and U1346 (N_1346,In_423,In_1254);
or U1347 (N_1347,In_495,In_996);
or U1348 (N_1348,In_588,In_409);
nand U1349 (N_1349,In_1457,In_1379);
nand U1350 (N_1350,In_1377,In_484);
nor U1351 (N_1351,In_13,In_984);
nor U1352 (N_1352,In_859,In_79);
and U1353 (N_1353,In_794,In_733);
nor U1354 (N_1354,In_158,In_878);
nor U1355 (N_1355,In_1490,In_792);
and U1356 (N_1356,In_354,In_805);
or U1357 (N_1357,In_799,In_282);
nand U1358 (N_1358,In_545,In_882);
and U1359 (N_1359,In_481,In_169);
or U1360 (N_1360,In_681,In_19);
and U1361 (N_1361,In_568,In_822);
nor U1362 (N_1362,In_2,In_1455);
nand U1363 (N_1363,In_1462,In_546);
and U1364 (N_1364,In_614,In_822);
nand U1365 (N_1365,In_1193,In_236);
nand U1366 (N_1366,In_69,In_543);
nor U1367 (N_1367,In_1141,In_141);
nand U1368 (N_1368,In_585,In_494);
nand U1369 (N_1369,In_1329,In_733);
or U1370 (N_1370,In_401,In_763);
nor U1371 (N_1371,In_943,In_404);
or U1372 (N_1372,In_185,In_103);
nor U1373 (N_1373,In_817,In_535);
or U1374 (N_1374,In_353,In_606);
and U1375 (N_1375,In_417,In_911);
and U1376 (N_1376,In_965,In_1);
nor U1377 (N_1377,In_863,In_490);
nor U1378 (N_1378,In_389,In_764);
nor U1379 (N_1379,In_113,In_1217);
nor U1380 (N_1380,In_1116,In_1479);
and U1381 (N_1381,In_8,In_284);
nand U1382 (N_1382,In_1459,In_569);
nor U1383 (N_1383,In_1204,In_1184);
and U1384 (N_1384,In_702,In_1285);
nor U1385 (N_1385,In_1370,In_526);
nand U1386 (N_1386,In_1422,In_132);
nor U1387 (N_1387,In_51,In_1147);
nor U1388 (N_1388,In_1163,In_328);
or U1389 (N_1389,In_290,In_1470);
nor U1390 (N_1390,In_642,In_1113);
nand U1391 (N_1391,In_359,In_553);
nor U1392 (N_1392,In_1055,In_689);
or U1393 (N_1393,In_146,In_227);
nor U1394 (N_1394,In_724,In_967);
nand U1395 (N_1395,In_1024,In_710);
and U1396 (N_1396,In_1061,In_710);
nor U1397 (N_1397,In_24,In_1273);
nor U1398 (N_1398,In_1340,In_1358);
nand U1399 (N_1399,In_1309,In_1081);
nor U1400 (N_1400,In_367,In_577);
or U1401 (N_1401,In_166,In_802);
and U1402 (N_1402,In_574,In_1030);
and U1403 (N_1403,In_1159,In_773);
or U1404 (N_1404,In_1054,In_1066);
nand U1405 (N_1405,In_1238,In_765);
nand U1406 (N_1406,In_464,In_418);
and U1407 (N_1407,In_1259,In_328);
nand U1408 (N_1408,In_1226,In_972);
nand U1409 (N_1409,In_178,In_1350);
and U1410 (N_1410,In_862,In_963);
nor U1411 (N_1411,In_1017,In_797);
and U1412 (N_1412,In_1179,In_848);
nand U1413 (N_1413,In_802,In_26);
and U1414 (N_1414,In_173,In_872);
and U1415 (N_1415,In_980,In_616);
or U1416 (N_1416,In_1386,In_443);
nand U1417 (N_1417,In_436,In_961);
or U1418 (N_1418,In_1120,In_461);
nor U1419 (N_1419,In_516,In_1024);
or U1420 (N_1420,In_656,In_1258);
or U1421 (N_1421,In_998,In_320);
nand U1422 (N_1422,In_465,In_482);
nor U1423 (N_1423,In_1255,In_81);
nor U1424 (N_1424,In_1398,In_1347);
or U1425 (N_1425,In_14,In_106);
nor U1426 (N_1426,In_931,In_1436);
nand U1427 (N_1427,In_1109,In_271);
nand U1428 (N_1428,In_88,In_299);
nand U1429 (N_1429,In_1341,In_545);
or U1430 (N_1430,In_395,In_1162);
nor U1431 (N_1431,In_160,In_369);
nand U1432 (N_1432,In_485,In_643);
nand U1433 (N_1433,In_1369,In_751);
and U1434 (N_1434,In_202,In_1040);
nand U1435 (N_1435,In_1253,In_125);
nor U1436 (N_1436,In_637,In_299);
or U1437 (N_1437,In_1496,In_91);
and U1438 (N_1438,In_957,In_202);
and U1439 (N_1439,In_489,In_602);
nor U1440 (N_1440,In_1399,In_899);
and U1441 (N_1441,In_516,In_1272);
or U1442 (N_1442,In_1423,In_43);
or U1443 (N_1443,In_619,In_5);
or U1444 (N_1444,In_694,In_1055);
xnor U1445 (N_1445,In_494,In_964);
and U1446 (N_1446,In_635,In_1131);
and U1447 (N_1447,In_1418,In_820);
nand U1448 (N_1448,In_923,In_366);
nor U1449 (N_1449,In_423,In_50);
nor U1450 (N_1450,In_1203,In_891);
nor U1451 (N_1451,In_1327,In_780);
nand U1452 (N_1452,In_463,In_765);
nand U1453 (N_1453,In_75,In_47);
nand U1454 (N_1454,In_1248,In_1235);
or U1455 (N_1455,In_1231,In_1324);
xnor U1456 (N_1456,In_285,In_563);
nand U1457 (N_1457,In_953,In_368);
or U1458 (N_1458,In_1357,In_287);
or U1459 (N_1459,In_733,In_573);
nand U1460 (N_1460,In_297,In_1227);
nand U1461 (N_1461,In_558,In_1246);
nor U1462 (N_1462,In_120,In_1246);
nor U1463 (N_1463,In_1333,In_881);
or U1464 (N_1464,In_334,In_162);
nand U1465 (N_1465,In_590,In_1494);
nand U1466 (N_1466,In_656,In_1196);
and U1467 (N_1467,In_321,In_474);
and U1468 (N_1468,In_1382,In_594);
and U1469 (N_1469,In_1467,In_1164);
or U1470 (N_1470,In_19,In_1190);
nor U1471 (N_1471,In_823,In_1283);
nand U1472 (N_1472,In_341,In_40);
or U1473 (N_1473,In_56,In_679);
nor U1474 (N_1474,In_988,In_102);
and U1475 (N_1475,In_1304,In_508);
or U1476 (N_1476,In_1031,In_1208);
nand U1477 (N_1477,In_1174,In_593);
and U1478 (N_1478,In_600,In_595);
nand U1479 (N_1479,In_1366,In_211);
and U1480 (N_1480,In_1374,In_143);
nor U1481 (N_1481,In_357,In_856);
nor U1482 (N_1482,In_1005,In_1275);
nand U1483 (N_1483,In_521,In_1486);
or U1484 (N_1484,In_1392,In_1238);
and U1485 (N_1485,In_887,In_1158);
nand U1486 (N_1486,In_1382,In_206);
nand U1487 (N_1487,In_1074,In_1130);
or U1488 (N_1488,In_1316,In_1066);
nor U1489 (N_1489,In_135,In_453);
nand U1490 (N_1490,In_401,In_708);
and U1491 (N_1491,In_449,In_243);
or U1492 (N_1492,In_1226,In_713);
nand U1493 (N_1493,In_1425,In_284);
nor U1494 (N_1494,In_685,In_440);
nand U1495 (N_1495,In_98,In_1264);
nand U1496 (N_1496,In_302,In_1491);
nor U1497 (N_1497,In_761,In_1301);
nand U1498 (N_1498,In_957,In_735);
or U1499 (N_1499,In_954,In_681);
or U1500 (N_1500,In_1483,In_1091);
and U1501 (N_1501,In_60,In_24);
and U1502 (N_1502,In_685,In_1131);
nor U1503 (N_1503,In_1442,In_863);
or U1504 (N_1504,In_123,In_91);
nand U1505 (N_1505,In_1128,In_777);
nand U1506 (N_1506,In_671,In_102);
and U1507 (N_1507,In_1203,In_1003);
or U1508 (N_1508,In_1323,In_1482);
or U1509 (N_1509,In_1016,In_789);
or U1510 (N_1510,In_63,In_977);
xor U1511 (N_1511,In_276,In_349);
nand U1512 (N_1512,In_16,In_102);
and U1513 (N_1513,In_618,In_768);
and U1514 (N_1514,In_458,In_355);
nand U1515 (N_1515,In_543,In_883);
nor U1516 (N_1516,In_224,In_1045);
or U1517 (N_1517,In_201,In_613);
nor U1518 (N_1518,In_602,In_201);
and U1519 (N_1519,In_860,In_753);
nand U1520 (N_1520,In_889,In_60);
nor U1521 (N_1521,In_1067,In_1323);
nand U1522 (N_1522,In_445,In_300);
and U1523 (N_1523,In_451,In_474);
nand U1524 (N_1524,In_1258,In_678);
nand U1525 (N_1525,In_868,In_716);
nand U1526 (N_1526,In_678,In_984);
or U1527 (N_1527,In_1320,In_942);
and U1528 (N_1528,In_924,In_347);
nand U1529 (N_1529,In_920,In_1457);
or U1530 (N_1530,In_55,In_397);
nor U1531 (N_1531,In_1192,In_411);
nor U1532 (N_1532,In_115,In_1113);
nand U1533 (N_1533,In_351,In_5);
nand U1534 (N_1534,In_927,In_1400);
nand U1535 (N_1535,In_572,In_257);
or U1536 (N_1536,In_1062,In_783);
and U1537 (N_1537,In_100,In_105);
nor U1538 (N_1538,In_1067,In_1008);
nor U1539 (N_1539,In_279,In_781);
or U1540 (N_1540,In_529,In_505);
nor U1541 (N_1541,In_936,In_446);
and U1542 (N_1542,In_1378,In_1119);
nand U1543 (N_1543,In_851,In_1268);
or U1544 (N_1544,In_576,In_394);
nor U1545 (N_1545,In_780,In_224);
and U1546 (N_1546,In_1403,In_889);
nand U1547 (N_1547,In_802,In_1419);
or U1548 (N_1548,In_1454,In_84);
nand U1549 (N_1549,In_1041,In_617);
and U1550 (N_1550,In_973,In_378);
nor U1551 (N_1551,In_653,In_1000);
nor U1552 (N_1552,In_509,In_1000);
or U1553 (N_1553,In_446,In_1180);
nor U1554 (N_1554,In_1183,In_1021);
nand U1555 (N_1555,In_1159,In_17);
nor U1556 (N_1556,In_617,In_556);
and U1557 (N_1557,In_27,In_1098);
nand U1558 (N_1558,In_226,In_510);
nand U1559 (N_1559,In_62,In_1000);
or U1560 (N_1560,In_943,In_891);
or U1561 (N_1561,In_627,In_222);
and U1562 (N_1562,In_856,In_794);
or U1563 (N_1563,In_238,In_1135);
or U1564 (N_1564,In_865,In_859);
nand U1565 (N_1565,In_591,In_570);
or U1566 (N_1566,In_1305,In_595);
and U1567 (N_1567,In_579,In_221);
and U1568 (N_1568,In_234,In_1372);
nand U1569 (N_1569,In_658,In_1446);
and U1570 (N_1570,In_891,In_575);
nand U1571 (N_1571,In_411,In_1302);
nand U1572 (N_1572,In_985,In_119);
or U1573 (N_1573,In_70,In_739);
and U1574 (N_1574,In_1315,In_567);
and U1575 (N_1575,In_1304,In_72);
nand U1576 (N_1576,In_635,In_804);
nor U1577 (N_1577,In_910,In_1238);
nand U1578 (N_1578,In_56,In_50);
and U1579 (N_1579,In_1325,In_223);
and U1580 (N_1580,In_201,In_679);
nand U1581 (N_1581,In_477,In_1103);
or U1582 (N_1582,In_808,In_34);
or U1583 (N_1583,In_1442,In_555);
or U1584 (N_1584,In_497,In_138);
nor U1585 (N_1585,In_1419,In_1112);
nor U1586 (N_1586,In_728,In_899);
xor U1587 (N_1587,In_131,In_196);
and U1588 (N_1588,In_994,In_1004);
and U1589 (N_1589,In_953,In_1339);
or U1590 (N_1590,In_1178,In_982);
nand U1591 (N_1591,In_1370,In_251);
or U1592 (N_1592,In_1208,In_1027);
nor U1593 (N_1593,In_910,In_1181);
nor U1594 (N_1594,In_48,In_23);
and U1595 (N_1595,In_242,In_667);
nor U1596 (N_1596,In_1449,In_1496);
or U1597 (N_1597,In_1432,In_308);
nor U1598 (N_1598,In_1239,In_793);
and U1599 (N_1599,In_1193,In_1448);
nor U1600 (N_1600,In_1318,In_1195);
nand U1601 (N_1601,In_53,In_934);
nand U1602 (N_1602,In_121,In_117);
xor U1603 (N_1603,In_118,In_1431);
or U1604 (N_1604,In_1361,In_116);
xnor U1605 (N_1605,In_1479,In_102);
nand U1606 (N_1606,In_989,In_749);
nand U1607 (N_1607,In_312,In_1357);
or U1608 (N_1608,In_459,In_623);
nor U1609 (N_1609,In_1448,In_99);
nand U1610 (N_1610,In_520,In_376);
or U1611 (N_1611,In_1294,In_784);
xor U1612 (N_1612,In_149,In_288);
and U1613 (N_1613,In_1090,In_1239);
nand U1614 (N_1614,In_1217,In_683);
and U1615 (N_1615,In_40,In_816);
nand U1616 (N_1616,In_401,In_694);
nor U1617 (N_1617,In_786,In_1280);
nand U1618 (N_1618,In_1360,In_908);
and U1619 (N_1619,In_527,In_21);
nor U1620 (N_1620,In_1270,In_1210);
nand U1621 (N_1621,In_1156,In_371);
nor U1622 (N_1622,In_900,In_424);
nand U1623 (N_1623,In_184,In_374);
or U1624 (N_1624,In_851,In_27);
nand U1625 (N_1625,In_471,In_697);
nand U1626 (N_1626,In_1458,In_737);
or U1627 (N_1627,In_1351,In_1348);
nor U1628 (N_1628,In_588,In_1003);
nor U1629 (N_1629,In_708,In_263);
nand U1630 (N_1630,In_927,In_184);
or U1631 (N_1631,In_1152,In_1243);
or U1632 (N_1632,In_361,In_1266);
nor U1633 (N_1633,In_688,In_478);
or U1634 (N_1634,In_1404,In_453);
nand U1635 (N_1635,In_330,In_369);
nor U1636 (N_1636,In_447,In_354);
and U1637 (N_1637,In_161,In_447);
nor U1638 (N_1638,In_1422,In_622);
or U1639 (N_1639,In_636,In_80);
and U1640 (N_1640,In_204,In_762);
and U1641 (N_1641,In_920,In_347);
or U1642 (N_1642,In_916,In_1163);
and U1643 (N_1643,In_213,In_997);
or U1644 (N_1644,In_1074,In_417);
nor U1645 (N_1645,In_338,In_831);
nand U1646 (N_1646,In_1318,In_293);
or U1647 (N_1647,In_589,In_1385);
xor U1648 (N_1648,In_963,In_1346);
or U1649 (N_1649,In_526,In_1420);
or U1650 (N_1650,In_943,In_1192);
nor U1651 (N_1651,In_20,In_1424);
or U1652 (N_1652,In_1439,In_197);
nand U1653 (N_1653,In_591,In_1277);
nand U1654 (N_1654,In_1254,In_935);
nor U1655 (N_1655,In_1166,In_739);
and U1656 (N_1656,In_1025,In_484);
nand U1657 (N_1657,In_1046,In_56);
nand U1658 (N_1658,In_458,In_793);
nor U1659 (N_1659,In_175,In_79);
and U1660 (N_1660,In_1011,In_489);
and U1661 (N_1661,In_411,In_300);
and U1662 (N_1662,In_1132,In_193);
and U1663 (N_1663,In_974,In_1090);
or U1664 (N_1664,In_980,In_701);
nand U1665 (N_1665,In_1254,In_191);
or U1666 (N_1666,In_936,In_310);
and U1667 (N_1667,In_1361,In_72);
nor U1668 (N_1668,In_617,In_744);
nor U1669 (N_1669,In_1181,In_639);
or U1670 (N_1670,In_299,In_291);
nor U1671 (N_1671,In_351,In_1191);
or U1672 (N_1672,In_577,In_831);
nand U1673 (N_1673,In_436,In_837);
xnor U1674 (N_1674,In_1163,In_523);
and U1675 (N_1675,In_604,In_309);
or U1676 (N_1676,In_232,In_329);
nor U1677 (N_1677,In_539,In_837);
nor U1678 (N_1678,In_462,In_317);
or U1679 (N_1679,In_1088,In_1379);
nor U1680 (N_1680,In_1343,In_793);
nor U1681 (N_1681,In_305,In_797);
nand U1682 (N_1682,In_407,In_281);
nand U1683 (N_1683,In_823,In_750);
or U1684 (N_1684,In_1283,In_1111);
or U1685 (N_1685,In_623,In_447);
nor U1686 (N_1686,In_212,In_571);
or U1687 (N_1687,In_1489,In_1249);
nand U1688 (N_1688,In_978,In_860);
and U1689 (N_1689,In_1294,In_65);
or U1690 (N_1690,In_183,In_405);
nor U1691 (N_1691,In_307,In_1383);
nand U1692 (N_1692,In_781,In_362);
or U1693 (N_1693,In_300,In_1379);
nor U1694 (N_1694,In_201,In_736);
or U1695 (N_1695,In_511,In_836);
and U1696 (N_1696,In_1296,In_1195);
nor U1697 (N_1697,In_243,In_1389);
nor U1698 (N_1698,In_914,In_20);
and U1699 (N_1699,In_535,In_543);
or U1700 (N_1700,In_684,In_179);
and U1701 (N_1701,In_727,In_920);
nand U1702 (N_1702,In_843,In_365);
or U1703 (N_1703,In_721,In_864);
and U1704 (N_1704,In_1121,In_752);
nand U1705 (N_1705,In_164,In_157);
or U1706 (N_1706,In_1207,In_946);
nand U1707 (N_1707,In_293,In_691);
nor U1708 (N_1708,In_736,In_429);
or U1709 (N_1709,In_1107,In_1389);
nand U1710 (N_1710,In_1055,In_160);
nor U1711 (N_1711,In_21,In_831);
nor U1712 (N_1712,In_1494,In_341);
nor U1713 (N_1713,In_331,In_1185);
and U1714 (N_1714,In_1161,In_535);
nand U1715 (N_1715,In_1061,In_1351);
nand U1716 (N_1716,In_348,In_80);
xnor U1717 (N_1717,In_621,In_1444);
nor U1718 (N_1718,In_1010,In_1357);
or U1719 (N_1719,In_269,In_736);
nand U1720 (N_1720,In_470,In_1336);
nand U1721 (N_1721,In_1082,In_635);
nor U1722 (N_1722,In_612,In_1104);
or U1723 (N_1723,In_1343,In_877);
or U1724 (N_1724,In_1110,In_1206);
nor U1725 (N_1725,In_1480,In_1418);
or U1726 (N_1726,In_713,In_270);
nand U1727 (N_1727,In_235,In_1144);
nand U1728 (N_1728,In_142,In_878);
nor U1729 (N_1729,In_643,In_282);
or U1730 (N_1730,In_146,In_421);
nand U1731 (N_1731,In_1371,In_764);
and U1732 (N_1732,In_1336,In_690);
and U1733 (N_1733,In_536,In_1471);
and U1734 (N_1734,In_387,In_1218);
nand U1735 (N_1735,In_497,In_285);
and U1736 (N_1736,In_146,In_1352);
nor U1737 (N_1737,In_889,In_267);
and U1738 (N_1738,In_832,In_1067);
nand U1739 (N_1739,In_38,In_337);
xor U1740 (N_1740,In_503,In_158);
or U1741 (N_1741,In_645,In_156);
and U1742 (N_1742,In_341,In_912);
nand U1743 (N_1743,In_1399,In_890);
nand U1744 (N_1744,In_1157,In_605);
nor U1745 (N_1745,In_1458,In_1427);
nor U1746 (N_1746,In_1039,In_842);
nand U1747 (N_1747,In_288,In_1383);
nor U1748 (N_1748,In_1436,In_1122);
nand U1749 (N_1749,In_1143,In_442);
or U1750 (N_1750,In_827,In_1162);
nand U1751 (N_1751,In_1012,In_1233);
nor U1752 (N_1752,In_278,In_105);
and U1753 (N_1753,In_748,In_491);
nor U1754 (N_1754,In_543,In_943);
nor U1755 (N_1755,In_1297,In_1339);
xnor U1756 (N_1756,In_46,In_1352);
nand U1757 (N_1757,In_1039,In_1151);
nor U1758 (N_1758,In_828,In_862);
nor U1759 (N_1759,In_1279,In_724);
xnor U1760 (N_1760,In_925,In_1177);
and U1761 (N_1761,In_1437,In_764);
or U1762 (N_1762,In_887,In_1400);
nand U1763 (N_1763,In_864,In_176);
nor U1764 (N_1764,In_1247,In_748);
nand U1765 (N_1765,In_459,In_1082);
and U1766 (N_1766,In_209,In_1038);
or U1767 (N_1767,In_29,In_657);
nor U1768 (N_1768,In_1109,In_593);
or U1769 (N_1769,In_892,In_1369);
nor U1770 (N_1770,In_802,In_443);
or U1771 (N_1771,In_324,In_403);
and U1772 (N_1772,In_539,In_1098);
nor U1773 (N_1773,In_60,In_251);
and U1774 (N_1774,In_1048,In_1249);
or U1775 (N_1775,In_965,In_238);
nor U1776 (N_1776,In_1284,In_932);
or U1777 (N_1777,In_50,In_654);
and U1778 (N_1778,In_931,In_341);
or U1779 (N_1779,In_350,In_526);
or U1780 (N_1780,In_372,In_29);
and U1781 (N_1781,In_277,In_1216);
or U1782 (N_1782,In_171,In_302);
nor U1783 (N_1783,In_1393,In_1246);
and U1784 (N_1784,In_775,In_1132);
or U1785 (N_1785,In_908,In_1407);
nand U1786 (N_1786,In_197,In_1411);
or U1787 (N_1787,In_67,In_1221);
nor U1788 (N_1788,In_1424,In_164);
and U1789 (N_1789,In_449,In_309);
nand U1790 (N_1790,In_840,In_1176);
nor U1791 (N_1791,In_200,In_69);
or U1792 (N_1792,In_173,In_1459);
or U1793 (N_1793,In_232,In_46);
and U1794 (N_1794,In_257,In_284);
nor U1795 (N_1795,In_234,In_823);
nand U1796 (N_1796,In_580,In_131);
and U1797 (N_1797,In_1247,In_829);
nand U1798 (N_1798,In_70,In_616);
or U1799 (N_1799,In_916,In_764);
nor U1800 (N_1800,In_642,In_677);
or U1801 (N_1801,In_825,In_833);
nor U1802 (N_1802,In_718,In_1242);
nand U1803 (N_1803,In_857,In_1389);
and U1804 (N_1804,In_645,In_820);
nand U1805 (N_1805,In_1325,In_1312);
or U1806 (N_1806,In_1281,In_546);
or U1807 (N_1807,In_1210,In_3);
nor U1808 (N_1808,In_806,In_511);
nor U1809 (N_1809,In_508,In_843);
nand U1810 (N_1810,In_584,In_1199);
or U1811 (N_1811,In_1043,In_875);
or U1812 (N_1812,In_360,In_634);
and U1813 (N_1813,In_165,In_308);
nor U1814 (N_1814,In_548,In_1456);
or U1815 (N_1815,In_1093,In_1417);
or U1816 (N_1816,In_525,In_1484);
nand U1817 (N_1817,In_1499,In_752);
nand U1818 (N_1818,In_41,In_814);
xnor U1819 (N_1819,In_1314,In_907);
and U1820 (N_1820,In_896,In_980);
nand U1821 (N_1821,In_477,In_1394);
nand U1822 (N_1822,In_1173,In_1499);
nor U1823 (N_1823,In_507,In_103);
nor U1824 (N_1824,In_1443,In_765);
nor U1825 (N_1825,In_1493,In_917);
xnor U1826 (N_1826,In_276,In_318);
or U1827 (N_1827,In_392,In_1345);
and U1828 (N_1828,In_102,In_150);
and U1829 (N_1829,In_209,In_564);
nand U1830 (N_1830,In_28,In_1451);
xor U1831 (N_1831,In_56,In_628);
nor U1832 (N_1832,In_316,In_440);
nand U1833 (N_1833,In_194,In_782);
nand U1834 (N_1834,In_248,In_344);
nand U1835 (N_1835,In_89,In_1218);
nor U1836 (N_1836,In_420,In_749);
nand U1837 (N_1837,In_1109,In_273);
or U1838 (N_1838,In_860,In_1002);
or U1839 (N_1839,In_1053,In_1275);
or U1840 (N_1840,In_377,In_118);
and U1841 (N_1841,In_101,In_976);
xor U1842 (N_1842,In_831,In_440);
and U1843 (N_1843,In_1249,In_1449);
nor U1844 (N_1844,In_1187,In_1316);
nor U1845 (N_1845,In_647,In_785);
nor U1846 (N_1846,In_1141,In_1459);
or U1847 (N_1847,In_898,In_522);
xnor U1848 (N_1848,In_747,In_218);
nand U1849 (N_1849,In_419,In_567);
and U1850 (N_1850,In_559,In_1161);
and U1851 (N_1851,In_1203,In_837);
nand U1852 (N_1852,In_246,In_906);
and U1853 (N_1853,In_1163,In_650);
nor U1854 (N_1854,In_700,In_1064);
and U1855 (N_1855,In_174,In_175);
nand U1856 (N_1856,In_446,In_7);
or U1857 (N_1857,In_1439,In_685);
nor U1858 (N_1858,In_272,In_149);
nand U1859 (N_1859,In_496,In_471);
nor U1860 (N_1860,In_143,In_1219);
nor U1861 (N_1861,In_1001,In_1301);
and U1862 (N_1862,In_1051,In_1373);
nor U1863 (N_1863,In_31,In_1175);
or U1864 (N_1864,In_456,In_144);
nand U1865 (N_1865,In_1424,In_410);
nor U1866 (N_1866,In_623,In_1187);
or U1867 (N_1867,In_817,In_829);
nor U1868 (N_1868,In_1197,In_531);
and U1869 (N_1869,In_966,In_797);
nor U1870 (N_1870,In_102,In_109);
nand U1871 (N_1871,In_1401,In_90);
and U1872 (N_1872,In_1293,In_244);
nand U1873 (N_1873,In_636,In_946);
nor U1874 (N_1874,In_126,In_1056);
or U1875 (N_1875,In_1235,In_1003);
nor U1876 (N_1876,In_147,In_871);
or U1877 (N_1877,In_352,In_424);
and U1878 (N_1878,In_1245,In_1416);
nor U1879 (N_1879,In_490,In_550);
or U1880 (N_1880,In_1381,In_1346);
nor U1881 (N_1881,In_358,In_241);
nor U1882 (N_1882,In_262,In_980);
and U1883 (N_1883,In_1393,In_94);
and U1884 (N_1884,In_84,In_937);
nor U1885 (N_1885,In_578,In_1402);
and U1886 (N_1886,In_620,In_1230);
nand U1887 (N_1887,In_1277,In_524);
nor U1888 (N_1888,In_604,In_959);
nand U1889 (N_1889,In_819,In_58);
and U1890 (N_1890,In_1143,In_359);
nand U1891 (N_1891,In_1062,In_677);
nand U1892 (N_1892,In_1430,In_681);
nor U1893 (N_1893,In_481,In_914);
and U1894 (N_1894,In_254,In_487);
and U1895 (N_1895,In_1441,In_1143);
xor U1896 (N_1896,In_722,In_1114);
and U1897 (N_1897,In_590,In_804);
nor U1898 (N_1898,In_1367,In_441);
or U1899 (N_1899,In_901,In_585);
nor U1900 (N_1900,In_1459,In_968);
or U1901 (N_1901,In_847,In_13);
xor U1902 (N_1902,In_366,In_23);
nand U1903 (N_1903,In_22,In_1000);
nor U1904 (N_1904,In_72,In_651);
nor U1905 (N_1905,In_972,In_485);
or U1906 (N_1906,In_243,In_200);
and U1907 (N_1907,In_192,In_1479);
or U1908 (N_1908,In_496,In_133);
nand U1909 (N_1909,In_114,In_108);
nand U1910 (N_1910,In_1473,In_1238);
and U1911 (N_1911,In_828,In_1007);
or U1912 (N_1912,In_378,In_320);
or U1913 (N_1913,In_782,In_1069);
or U1914 (N_1914,In_569,In_266);
xor U1915 (N_1915,In_778,In_270);
xor U1916 (N_1916,In_707,In_806);
or U1917 (N_1917,In_150,In_938);
or U1918 (N_1918,In_971,In_1326);
nand U1919 (N_1919,In_348,In_1085);
or U1920 (N_1920,In_957,In_1287);
nor U1921 (N_1921,In_1373,In_1462);
nand U1922 (N_1922,In_176,In_862);
nand U1923 (N_1923,In_1430,In_338);
and U1924 (N_1924,In_1000,In_441);
nor U1925 (N_1925,In_1352,In_349);
and U1926 (N_1926,In_329,In_1144);
and U1927 (N_1927,In_1271,In_43);
and U1928 (N_1928,In_419,In_1250);
nand U1929 (N_1929,In_120,In_532);
nor U1930 (N_1930,In_366,In_1452);
and U1931 (N_1931,In_342,In_139);
nand U1932 (N_1932,In_636,In_748);
nor U1933 (N_1933,In_1346,In_103);
nand U1934 (N_1934,In_281,In_320);
nand U1935 (N_1935,In_379,In_1307);
or U1936 (N_1936,In_24,In_227);
or U1937 (N_1937,In_1074,In_370);
nand U1938 (N_1938,In_654,In_1278);
and U1939 (N_1939,In_607,In_1059);
nor U1940 (N_1940,In_87,In_1172);
or U1941 (N_1941,In_122,In_985);
nor U1942 (N_1942,In_328,In_1146);
and U1943 (N_1943,In_849,In_299);
xor U1944 (N_1944,In_1091,In_1264);
and U1945 (N_1945,In_1181,In_851);
and U1946 (N_1946,In_452,In_493);
or U1947 (N_1947,In_824,In_1278);
or U1948 (N_1948,In_1014,In_600);
nand U1949 (N_1949,In_1458,In_490);
nor U1950 (N_1950,In_1331,In_104);
and U1951 (N_1951,In_145,In_508);
or U1952 (N_1952,In_130,In_765);
and U1953 (N_1953,In_1125,In_1033);
nand U1954 (N_1954,In_1185,In_168);
nand U1955 (N_1955,In_521,In_304);
nand U1956 (N_1956,In_342,In_1396);
or U1957 (N_1957,In_1060,In_583);
nor U1958 (N_1958,In_22,In_504);
and U1959 (N_1959,In_1017,In_1181);
and U1960 (N_1960,In_217,In_419);
nand U1961 (N_1961,In_999,In_178);
and U1962 (N_1962,In_1288,In_864);
nor U1963 (N_1963,In_1385,In_317);
or U1964 (N_1964,In_1355,In_1025);
nor U1965 (N_1965,In_279,In_1074);
and U1966 (N_1966,In_422,In_751);
nor U1967 (N_1967,In_870,In_628);
nor U1968 (N_1968,In_1373,In_744);
or U1969 (N_1969,In_74,In_792);
nand U1970 (N_1970,In_62,In_344);
or U1971 (N_1971,In_1484,In_1239);
and U1972 (N_1972,In_617,In_897);
nand U1973 (N_1973,In_845,In_649);
or U1974 (N_1974,In_623,In_741);
or U1975 (N_1975,In_1326,In_514);
nor U1976 (N_1976,In_83,In_1364);
nand U1977 (N_1977,In_1325,In_411);
or U1978 (N_1978,In_954,In_847);
or U1979 (N_1979,In_736,In_767);
or U1980 (N_1980,In_294,In_138);
nand U1981 (N_1981,In_150,In_1435);
or U1982 (N_1982,In_565,In_422);
nand U1983 (N_1983,In_862,In_193);
nand U1984 (N_1984,In_1002,In_1113);
and U1985 (N_1985,In_650,In_238);
and U1986 (N_1986,In_69,In_493);
nor U1987 (N_1987,In_635,In_225);
or U1988 (N_1988,In_1160,In_1020);
nor U1989 (N_1989,In_1232,In_1248);
nor U1990 (N_1990,In_346,In_257);
nand U1991 (N_1991,In_976,In_723);
nor U1992 (N_1992,In_381,In_891);
or U1993 (N_1993,In_849,In_555);
and U1994 (N_1994,In_970,In_1109);
and U1995 (N_1995,In_238,In_1037);
or U1996 (N_1996,In_693,In_688);
nand U1997 (N_1997,In_832,In_732);
or U1998 (N_1998,In_1466,In_401);
or U1999 (N_1999,In_1384,In_1266);
nand U2000 (N_2000,In_488,In_1383);
nand U2001 (N_2001,In_1352,In_323);
xor U2002 (N_2002,In_713,In_947);
and U2003 (N_2003,In_63,In_1327);
nor U2004 (N_2004,In_1320,In_813);
and U2005 (N_2005,In_480,In_527);
nand U2006 (N_2006,In_48,In_1470);
or U2007 (N_2007,In_200,In_388);
and U2008 (N_2008,In_230,In_1251);
nor U2009 (N_2009,In_364,In_156);
nand U2010 (N_2010,In_304,In_1056);
nand U2011 (N_2011,In_1196,In_923);
or U2012 (N_2012,In_634,In_61);
xor U2013 (N_2013,In_491,In_1280);
nand U2014 (N_2014,In_862,In_491);
nand U2015 (N_2015,In_1134,In_981);
or U2016 (N_2016,In_249,In_598);
and U2017 (N_2017,In_1334,In_36);
nand U2018 (N_2018,In_1127,In_646);
or U2019 (N_2019,In_1209,In_1012);
xnor U2020 (N_2020,In_481,In_237);
nand U2021 (N_2021,In_830,In_257);
nor U2022 (N_2022,In_542,In_1096);
nand U2023 (N_2023,In_188,In_518);
or U2024 (N_2024,In_1217,In_597);
and U2025 (N_2025,In_1442,In_780);
and U2026 (N_2026,In_229,In_1334);
or U2027 (N_2027,In_1458,In_691);
nand U2028 (N_2028,In_912,In_135);
nand U2029 (N_2029,In_583,In_1321);
or U2030 (N_2030,In_1188,In_1176);
xor U2031 (N_2031,In_1271,In_925);
nand U2032 (N_2032,In_721,In_804);
or U2033 (N_2033,In_1206,In_67);
and U2034 (N_2034,In_995,In_1085);
nor U2035 (N_2035,In_1360,In_299);
nor U2036 (N_2036,In_670,In_254);
nor U2037 (N_2037,In_690,In_227);
nor U2038 (N_2038,In_1258,In_204);
and U2039 (N_2039,In_122,In_354);
and U2040 (N_2040,In_457,In_867);
nor U2041 (N_2041,In_694,In_0);
nand U2042 (N_2042,In_33,In_1319);
and U2043 (N_2043,In_119,In_968);
nor U2044 (N_2044,In_1143,In_1478);
nand U2045 (N_2045,In_1073,In_1052);
or U2046 (N_2046,In_346,In_481);
xor U2047 (N_2047,In_294,In_1407);
and U2048 (N_2048,In_1069,In_459);
and U2049 (N_2049,In_584,In_144);
nand U2050 (N_2050,In_918,In_1003);
nor U2051 (N_2051,In_790,In_1329);
nor U2052 (N_2052,In_411,In_650);
or U2053 (N_2053,In_548,In_1041);
nor U2054 (N_2054,In_879,In_1414);
or U2055 (N_2055,In_1093,In_1490);
and U2056 (N_2056,In_577,In_368);
nor U2057 (N_2057,In_790,In_1365);
nand U2058 (N_2058,In_204,In_231);
nor U2059 (N_2059,In_952,In_1229);
nor U2060 (N_2060,In_952,In_237);
nand U2061 (N_2061,In_1476,In_630);
nor U2062 (N_2062,In_1412,In_1042);
nand U2063 (N_2063,In_408,In_1306);
nand U2064 (N_2064,In_443,In_260);
nand U2065 (N_2065,In_667,In_184);
or U2066 (N_2066,In_254,In_378);
or U2067 (N_2067,In_724,In_277);
xnor U2068 (N_2068,In_1421,In_1080);
and U2069 (N_2069,In_73,In_739);
nor U2070 (N_2070,In_1195,In_800);
nor U2071 (N_2071,In_1264,In_477);
and U2072 (N_2072,In_542,In_749);
nor U2073 (N_2073,In_870,In_254);
nand U2074 (N_2074,In_395,In_741);
nand U2075 (N_2075,In_1215,In_1123);
and U2076 (N_2076,In_165,In_1025);
nand U2077 (N_2077,In_41,In_945);
or U2078 (N_2078,In_230,In_882);
nand U2079 (N_2079,In_130,In_1208);
nor U2080 (N_2080,In_16,In_1203);
and U2081 (N_2081,In_276,In_268);
nor U2082 (N_2082,In_199,In_942);
and U2083 (N_2083,In_75,In_175);
nor U2084 (N_2084,In_48,In_507);
nand U2085 (N_2085,In_1235,In_497);
nor U2086 (N_2086,In_1283,In_378);
or U2087 (N_2087,In_240,In_248);
and U2088 (N_2088,In_921,In_664);
or U2089 (N_2089,In_679,In_572);
nor U2090 (N_2090,In_563,In_69);
or U2091 (N_2091,In_1158,In_1078);
nor U2092 (N_2092,In_923,In_998);
and U2093 (N_2093,In_156,In_104);
or U2094 (N_2094,In_18,In_147);
and U2095 (N_2095,In_1245,In_1302);
and U2096 (N_2096,In_1240,In_428);
nor U2097 (N_2097,In_406,In_1492);
or U2098 (N_2098,In_1472,In_416);
xor U2099 (N_2099,In_1106,In_1393);
nand U2100 (N_2100,In_1310,In_536);
xor U2101 (N_2101,In_972,In_303);
and U2102 (N_2102,In_426,In_646);
nor U2103 (N_2103,In_827,In_871);
and U2104 (N_2104,In_572,In_1362);
or U2105 (N_2105,In_613,In_178);
and U2106 (N_2106,In_507,In_1207);
xor U2107 (N_2107,In_314,In_626);
nor U2108 (N_2108,In_934,In_1120);
nor U2109 (N_2109,In_324,In_632);
or U2110 (N_2110,In_970,In_1209);
xor U2111 (N_2111,In_1104,In_558);
nor U2112 (N_2112,In_1476,In_1467);
or U2113 (N_2113,In_1412,In_1107);
xnor U2114 (N_2114,In_857,In_306);
xor U2115 (N_2115,In_728,In_2);
and U2116 (N_2116,In_915,In_299);
and U2117 (N_2117,In_690,In_817);
or U2118 (N_2118,In_326,In_570);
nor U2119 (N_2119,In_890,In_1010);
or U2120 (N_2120,In_266,In_415);
or U2121 (N_2121,In_1118,In_885);
and U2122 (N_2122,In_1107,In_1381);
and U2123 (N_2123,In_840,In_1404);
or U2124 (N_2124,In_803,In_19);
nor U2125 (N_2125,In_1150,In_789);
nand U2126 (N_2126,In_346,In_744);
nand U2127 (N_2127,In_867,In_897);
nand U2128 (N_2128,In_629,In_806);
nand U2129 (N_2129,In_1161,In_78);
or U2130 (N_2130,In_435,In_693);
nor U2131 (N_2131,In_1431,In_1096);
and U2132 (N_2132,In_1029,In_1194);
and U2133 (N_2133,In_132,In_812);
or U2134 (N_2134,In_760,In_1433);
or U2135 (N_2135,In_448,In_1404);
or U2136 (N_2136,In_970,In_1375);
nor U2137 (N_2137,In_453,In_659);
and U2138 (N_2138,In_543,In_267);
nand U2139 (N_2139,In_1138,In_721);
nor U2140 (N_2140,In_1015,In_1179);
or U2141 (N_2141,In_678,In_90);
and U2142 (N_2142,In_1172,In_156);
and U2143 (N_2143,In_945,In_1237);
and U2144 (N_2144,In_742,In_191);
and U2145 (N_2145,In_308,In_1342);
nor U2146 (N_2146,In_725,In_224);
and U2147 (N_2147,In_515,In_981);
nor U2148 (N_2148,In_856,In_1183);
or U2149 (N_2149,In_185,In_3);
or U2150 (N_2150,In_1462,In_1163);
and U2151 (N_2151,In_676,In_493);
and U2152 (N_2152,In_674,In_1249);
or U2153 (N_2153,In_96,In_1162);
or U2154 (N_2154,In_152,In_834);
or U2155 (N_2155,In_1242,In_685);
nor U2156 (N_2156,In_869,In_1292);
or U2157 (N_2157,In_224,In_549);
nor U2158 (N_2158,In_1498,In_1151);
nand U2159 (N_2159,In_1244,In_1260);
and U2160 (N_2160,In_1212,In_1204);
and U2161 (N_2161,In_931,In_438);
xnor U2162 (N_2162,In_1134,In_755);
or U2163 (N_2163,In_1362,In_1303);
or U2164 (N_2164,In_524,In_166);
or U2165 (N_2165,In_745,In_1380);
nor U2166 (N_2166,In_639,In_216);
nor U2167 (N_2167,In_269,In_359);
or U2168 (N_2168,In_866,In_1183);
and U2169 (N_2169,In_469,In_1368);
and U2170 (N_2170,In_505,In_345);
nor U2171 (N_2171,In_1328,In_270);
nor U2172 (N_2172,In_804,In_45);
and U2173 (N_2173,In_803,In_240);
and U2174 (N_2174,In_1291,In_353);
or U2175 (N_2175,In_1359,In_245);
nand U2176 (N_2176,In_224,In_175);
nor U2177 (N_2177,In_419,In_1257);
and U2178 (N_2178,In_918,In_718);
nand U2179 (N_2179,In_992,In_262);
or U2180 (N_2180,In_1323,In_870);
or U2181 (N_2181,In_580,In_1356);
or U2182 (N_2182,In_1316,In_172);
and U2183 (N_2183,In_674,In_830);
or U2184 (N_2184,In_220,In_809);
and U2185 (N_2185,In_686,In_82);
or U2186 (N_2186,In_482,In_1497);
and U2187 (N_2187,In_183,In_958);
nor U2188 (N_2188,In_1189,In_1036);
or U2189 (N_2189,In_1163,In_334);
nor U2190 (N_2190,In_175,In_194);
nor U2191 (N_2191,In_985,In_387);
or U2192 (N_2192,In_180,In_652);
nor U2193 (N_2193,In_807,In_733);
or U2194 (N_2194,In_1238,In_166);
nor U2195 (N_2195,In_111,In_72);
nor U2196 (N_2196,In_819,In_1383);
or U2197 (N_2197,In_168,In_1192);
and U2198 (N_2198,In_666,In_1134);
or U2199 (N_2199,In_905,In_1123);
and U2200 (N_2200,In_8,In_1046);
or U2201 (N_2201,In_48,In_603);
and U2202 (N_2202,In_1499,In_561);
and U2203 (N_2203,In_1306,In_1400);
and U2204 (N_2204,In_814,In_1);
nand U2205 (N_2205,In_1025,In_728);
or U2206 (N_2206,In_754,In_452);
and U2207 (N_2207,In_1335,In_213);
nor U2208 (N_2208,In_558,In_207);
nand U2209 (N_2209,In_453,In_524);
nand U2210 (N_2210,In_938,In_388);
nor U2211 (N_2211,In_190,In_1322);
nor U2212 (N_2212,In_542,In_427);
and U2213 (N_2213,In_514,In_1287);
or U2214 (N_2214,In_1068,In_1043);
or U2215 (N_2215,In_6,In_419);
nor U2216 (N_2216,In_866,In_100);
or U2217 (N_2217,In_616,In_938);
or U2218 (N_2218,In_433,In_1372);
and U2219 (N_2219,In_138,In_764);
nor U2220 (N_2220,In_1246,In_150);
nand U2221 (N_2221,In_156,In_413);
and U2222 (N_2222,In_972,In_1263);
or U2223 (N_2223,In_498,In_50);
and U2224 (N_2224,In_973,In_812);
or U2225 (N_2225,In_1397,In_779);
nand U2226 (N_2226,In_505,In_814);
nand U2227 (N_2227,In_490,In_569);
and U2228 (N_2228,In_401,In_421);
nand U2229 (N_2229,In_297,In_983);
and U2230 (N_2230,In_1178,In_673);
nor U2231 (N_2231,In_1101,In_59);
nand U2232 (N_2232,In_1270,In_952);
or U2233 (N_2233,In_340,In_792);
nand U2234 (N_2234,In_480,In_1114);
xor U2235 (N_2235,In_820,In_585);
and U2236 (N_2236,In_588,In_888);
nand U2237 (N_2237,In_703,In_913);
nand U2238 (N_2238,In_173,In_238);
or U2239 (N_2239,In_11,In_475);
nand U2240 (N_2240,In_686,In_602);
or U2241 (N_2241,In_335,In_855);
nor U2242 (N_2242,In_314,In_967);
nand U2243 (N_2243,In_1283,In_1395);
and U2244 (N_2244,In_952,In_495);
nor U2245 (N_2245,In_1442,In_710);
nor U2246 (N_2246,In_707,In_80);
or U2247 (N_2247,In_1394,In_282);
or U2248 (N_2248,In_1099,In_378);
nor U2249 (N_2249,In_1323,In_839);
nor U2250 (N_2250,In_603,In_619);
nand U2251 (N_2251,In_154,In_1405);
and U2252 (N_2252,In_608,In_1294);
and U2253 (N_2253,In_1167,In_802);
xnor U2254 (N_2254,In_1028,In_1477);
or U2255 (N_2255,In_139,In_410);
or U2256 (N_2256,In_818,In_598);
nand U2257 (N_2257,In_120,In_112);
or U2258 (N_2258,In_872,In_334);
nand U2259 (N_2259,In_62,In_1184);
nor U2260 (N_2260,In_1052,In_1351);
nor U2261 (N_2261,In_1390,In_1035);
and U2262 (N_2262,In_733,In_716);
nor U2263 (N_2263,In_706,In_183);
nand U2264 (N_2264,In_517,In_783);
or U2265 (N_2265,In_768,In_1189);
or U2266 (N_2266,In_536,In_1009);
nor U2267 (N_2267,In_956,In_1166);
or U2268 (N_2268,In_1446,In_407);
or U2269 (N_2269,In_849,In_944);
or U2270 (N_2270,In_353,In_971);
nand U2271 (N_2271,In_802,In_1039);
nor U2272 (N_2272,In_1442,In_1017);
nand U2273 (N_2273,In_660,In_1197);
or U2274 (N_2274,In_1261,In_1016);
and U2275 (N_2275,In_718,In_899);
nand U2276 (N_2276,In_140,In_837);
nand U2277 (N_2277,In_888,In_691);
and U2278 (N_2278,In_917,In_762);
nor U2279 (N_2279,In_978,In_1459);
nand U2280 (N_2280,In_1132,In_369);
nand U2281 (N_2281,In_1378,In_33);
nand U2282 (N_2282,In_165,In_179);
and U2283 (N_2283,In_1274,In_784);
xnor U2284 (N_2284,In_1460,In_1142);
nor U2285 (N_2285,In_63,In_558);
or U2286 (N_2286,In_360,In_106);
nand U2287 (N_2287,In_607,In_32);
and U2288 (N_2288,In_35,In_203);
nor U2289 (N_2289,In_1046,In_1226);
and U2290 (N_2290,In_862,In_353);
and U2291 (N_2291,In_1254,In_715);
nor U2292 (N_2292,In_741,In_274);
or U2293 (N_2293,In_119,In_56);
nand U2294 (N_2294,In_357,In_1028);
nor U2295 (N_2295,In_876,In_67);
nand U2296 (N_2296,In_163,In_632);
and U2297 (N_2297,In_687,In_618);
nor U2298 (N_2298,In_473,In_632);
or U2299 (N_2299,In_225,In_1078);
nand U2300 (N_2300,In_495,In_517);
or U2301 (N_2301,In_968,In_1320);
or U2302 (N_2302,In_503,In_957);
or U2303 (N_2303,In_1324,In_1287);
nand U2304 (N_2304,In_271,In_838);
and U2305 (N_2305,In_1456,In_1110);
and U2306 (N_2306,In_1422,In_1296);
and U2307 (N_2307,In_393,In_911);
and U2308 (N_2308,In_640,In_342);
and U2309 (N_2309,In_124,In_1157);
nor U2310 (N_2310,In_713,In_1037);
nand U2311 (N_2311,In_1034,In_502);
nand U2312 (N_2312,In_681,In_1468);
and U2313 (N_2313,In_1117,In_432);
nand U2314 (N_2314,In_923,In_1491);
and U2315 (N_2315,In_889,In_284);
and U2316 (N_2316,In_396,In_734);
or U2317 (N_2317,In_1230,In_185);
or U2318 (N_2318,In_1301,In_912);
or U2319 (N_2319,In_65,In_1205);
or U2320 (N_2320,In_630,In_589);
and U2321 (N_2321,In_84,In_433);
xnor U2322 (N_2322,In_1425,In_112);
nand U2323 (N_2323,In_108,In_36);
and U2324 (N_2324,In_888,In_833);
nor U2325 (N_2325,In_1400,In_1197);
nand U2326 (N_2326,In_736,In_1374);
and U2327 (N_2327,In_1467,In_468);
nor U2328 (N_2328,In_1175,In_547);
or U2329 (N_2329,In_960,In_1332);
nand U2330 (N_2330,In_161,In_456);
nor U2331 (N_2331,In_224,In_998);
or U2332 (N_2332,In_405,In_549);
nor U2333 (N_2333,In_259,In_230);
nor U2334 (N_2334,In_1175,In_1466);
nand U2335 (N_2335,In_1411,In_793);
or U2336 (N_2336,In_348,In_265);
or U2337 (N_2337,In_1237,In_289);
or U2338 (N_2338,In_979,In_61);
or U2339 (N_2339,In_245,In_139);
or U2340 (N_2340,In_974,In_1433);
nand U2341 (N_2341,In_1009,In_1260);
and U2342 (N_2342,In_368,In_556);
or U2343 (N_2343,In_31,In_259);
nor U2344 (N_2344,In_978,In_1025);
nor U2345 (N_2345,In_1112,In_554);
or U2346 (N_2346,In_639,In_702);
or U2347 (N_2347,In_31,In_1436);
or U2348 (N_2348,In_1304,In_1434);
nand U2349 (N_2349,In_1261,In_284);
nand U2350 (N_2350,In_1263,In_605);
and U2351 (N_2351,In_1284,In_1257);
or U2352 (N_2352,In_1342,In_420);
and U2353 (N_2353,In_943,In_1114);
nor U2354 (N_2354,In_1248,In_157);
nor U2355 (N_2355,In_418,In_60);
xor U2356 (N_2356,In_297,In_577);
or U2357 (N_2357,In_1276,In_1187);
nand U2358 (N_2358,In_1147,In_897);
or U2359 (N_2359,In_922,In_1386);
nand U2360 (N_2360,In_509,In_247);
or U2361 (N_2361,In_506,In_1484);
nor U2362 (N_2362,In_517,In_804);
nor U2363 (N_2363,In_975,In_948);
or U2364 (N_2364,In_637,In_446);
or U2365 (N_2365,In_1121,In_1400);
or U2366 (N_2366,In_1444,In_899);
nor U2367 (N_2367,In_264,In_624);
nand U2368 (N_2368,In_924,In_221);
nor U2369 (N_2369,In_577,In_345);
nand U2370 (N_2370,In_2,In_487);
and U2371 (N_2371,In_77,In_61);
nor U2372 (N_2372,In_703,In_890);
nand U2373 (N_2373,In_831,In_1371);
nand U2374 (N_2374,In_1465,In_560);
nand U2375 (N_2375,In_1429,In_184);
and U2376 (N_2376,In_58,In_128);
and U2377 (N_2377,In_426,In_1414);
nand U2378 (N_2378,In_90,In_1468);
or U2379 (N_2379,In_811,In_1424);
nand U2380 (N_2380,In_1129,In_1478);
and U2381 (N_2381,In_45,In_643);
or U2382 (N_2382,In_503,In_215);
or U2383 (N_2383,In_142,In_218);
or U2384 (N_2384,In_267,In_203);
xnor U2385 (N_2385,In_1347,In_790);
nand U2386 (N_2386,In_60,In_1389);
and U2387 (N_2387,In_489,In_386);
nor U2388 (N_2388,In_910,In_883);
nor U2389 (N_2389,In_933,In_1180);
and U2390 (N_2390,In_1204,In_1497);
nor U2391 (N_2391,In_531,In_1194);
or U2392 (N_2392,In_890,In_959);
xnor U2393 (N_2393,In_380,In_84);
nand U2394 (N_2394,In_913,In_143);
nor U2395 (N_2395,In_483,In_171);
nor U2396 (N_2396,In_537,In_795);
or U2397 (N_2397,In_371,In_445);
nand U2398 (N_2398,In_1227,In_1224);
nand U2399 (N_2399,In_549,In_1207);
or U2400 (N_2400,In_990,In_12);
and U2401 (N_2401,In_1141,In_421);
and U2402 (N_2402,In_424,In_962);
nand U2403 (N_2403,In_657,In_755);
nand U2404 (N_2404,In_532,In_666);
and U2405 (N_2405,In_684,In_247);
or U2406 (N_2406,In_440,In_157);
nor U2407 (N_2407,In_1101,In_313);
and U2408 (N_2408,In_386,In_363);
nand U2409 (N_2409,In_1285,In_524);
or U2410 (N_2410,In_625,In_1482);
or U2411 (N_2411,In_1206,In_217);
nand U2412 (N_2412,In_1249,In_575);
and U2413 (N_2413,In_715,In_521);
nor U2414 (N_2414,In_239,In_271);
nand U2415 (N_2415,In_586,In_78);
or U2416 (N_2416,In_436,In_1399);
and U2417 (N_2417,In_987,In_257);
nor U2418 (N_2418,In_747,In_1035);
nor U2419 (N_2419,In_399,In_816);
and U2420 (N_2420,In_888,In_513);
or U2421 (N_2421,In_314,In_222);
and U2422 (N_2422,In_342,In_112);
nand U2423 (N_2423,In_797,In_1298);
nor U2424 (N_2424,In_696,In_1494);
and U2425 (N_2425,In_152,In_516);
nand U2426 (N_2426,In_1436,In_420);
or U2427 (N_2427,In_925,In_499);
nand U2428 (N_2428,In_1301,In_787);
nand U2429 (N_2429,In_508,In_629);
nand U2430 (N_2430,In_585,In_1032);
and U2431 (N_2431,In_1208,In_686);
nand U2432 (N_2432,In_953,In_770);
and U2433 (N_2433,In_933,In_218);
xor U2434 (N_2434,In_800,In_1079);
and U2435 (N_2435,In_844,In_792);
or U2436 (N_2436,In_377,In_1284);
and U2437 (N_2437,In_548,In_554);
and U2438 (N_2438,In_654,In_753);
nor U2439 (N_2439,In_1490,In_433);
nor U2440 (N_2440,In_393,In_728);
or U2441 (N_2441,In_1315,In_352);
xnor U2442 (N_2442,In_727,In_1021);
nor U2443 (N_2443,In_981,In_1065);
nor U2444 (N_2444,In_1171,In_1406);
or U2445 (N_2445,In_1494,In_244);
nand U2446 (N_2446,In_513,In_643);
and U2447 (N_2447,In_293,In_612);
and U2448 (N_2448,In_325,In_1452);
nor U2449 (N_2449,In_1176,In_943);
nand U2450 (N_2450,In_416,In_403);
or U2451 (N_2451,In_53,In_957);
nand U2452 (N_2452,In_1490,In_789);
or U2453 (N_2453,In_938,In_818);
nand U2454 (N_2454,In_1197,In_799);
nor U2455 (N_2455,In_309,In_72);
nand U2456 (N_2456,In_305,In_724);
nand U2457 (N_2457,In_260,In_1403);
nand U2458 (N_2458,In_980,In_1313);
nand U2459 (N_2459,In_543,In_983);
or U2460 (N_2460,In_535,In_872);
nand U2461 (N_2461,In_104,In_608);
nand U2462 (N_2462,In_1182,In_856);
or U2463 (N_2463,In_333,In_216);
nor U2464 (N_2464,In_431,In_1483);
nand U2465 (N_2465,In_913,In_821);
or U2466 (N_2466,In_1143,In_231);
nor U2467 (N_2467,In_1050,In_204);
and U2468 (N_2468,In_823,In_1040);
and U2469 (N_2469,In_397,In_1246);
and U2470 (N_2470,In_767,In_563);
nand U2471 (N_2471,In_65,In_378);
nor U2472 (N_2472,In_492,In_866);
and U2473 (N_2473,In_990,In_249);
or U2474 (N_2474,In_1292,In_146);
and U2475 (N_2475,In_962,In_366);
and U2476 (N_2476,In_1034,In_313);
nand U2477 (N_2477,In_1242,In_693);
and U2478 (N_2478,In_1076,In_1425);
or U2479 (N_2479,In_153,In_565);
nor U2480 (N_2480,In_452,In_1282);
xnor U2481 (N_2481,In_320,In_803);
nor U2482 (N_2482,In_709,In_557);
nand U2483 (N_2483,In_201,In_1179);
nor U2484 (N_2484,In_93,In_711);
and U2485 (N_2485,In_324,In_328);
and U2486 (N_2486,In_601,In_228);
and U2487 (N_2487,In_848,In_25);
and U2488 (N_2488,In_1066,In_652);
nand U2489 (N_2489,In_768,In_994);
and U2490 (N_2490,In_146,In_1494);
nand U2491 (N_2491,In_233,In_378);
and U2492 (N_2492,In_312,In_454);
nand U2493 (N_2493,In_1172,In_346);
or U2494 (N_2494,In_1291,In_1307);
or U2495 (N_2495,In_598,In_1273);
and U2496 (N_2496,In_1300,In_1461);
and U2497 (N_2497,In_1056,In_185);
or U2498 (N_2498,In_174,In_383);
nor U2499 (N_2499,In_1167,In_1452);
and U2500 (N_2500,In_810,In_64);
nor U2501 (N_2501,In_365,In_1078);
and U2502 (N_2502,In_223,In_198);
and U2503 (N_2503,In_305,In_252);
and U2504 (N_2504,In_410,In_279);
and U2505 (N_2505,In_1096,In_873);
or U2506 (N_2506,In_1373,In_98);
xnor U2507 (N_2507,In_1213,In_229);
nand U2508 (N_2508,In_936,In_1368);
and U2509 (N_2509,In_622,In_1416);
nand U2510 (N_2510,In_977,In_76);
nand U2511 (N_2511,In_936,In_66);
nand U2512 (N_2512,In_730,In_635);
nor U2513 (N_2513,In_220,In_1418);
nand U2514 (N_2514,In_306,In_1006);
or U2515 (N_2515,In_292,In_1049);
or U2516 (N_2516,In_13,In_581);
nand U2517 (N_2517,In_1258,In_947);
nand U2518 (N_2518,In_223,In_1307);
or U2519 (N_2519,In_1424,In_812);
xnor U2520 (N_2520,In_331,In_569);
nor U2521 (N_2521,In_118,In_101);
and U2522 (N_2522,In_268,In_349);
or U2523 (N_2523,In_840,In_1436);
and U2524 (N_2524,In_1268,In_360);
or U2525 (N_2525,In_1344,In_525);
nor U2526 (N_2526,In_1244,In_1375);
and U2527 (N_2527,In_1414,In_627);
nand U2528 (N_2528,In_762,In_1201);
nand U2529 (N_2529,In_1237,In_1008);
or U2530 (N_2530,In_726,In_1273);
or U2531 (N_2531,In_808,In_567);
and U2532 (N_2532,In_418,In_1358);
or U2533 (N_2533,In_1021,In_671);
and U2534 (N_2534,In_1226,In_175);
nor U2535 (N_2535,In_487,In_465);
or U2536 (N_2536,In_654,In_350);
nor U2537 (N_2537,In_816,In_1001);
or U2538 (N_2538,In_318,In_982);
and U2539 (N_2539,In_969,In_187);
or U2540 (N_2540,In_458,In_790);
or U2541 (N_2541,In_1242,In_705);
nand U2542 (N_2542,In_355,In_945);
nand U2543 (N_2543,In_396,In_1342);
nor U2544 (N_2544,In_995,In_203);
or U2545 (N_2545,In_893,In_1249);
or U2546 (N_2546,In_1200,In_436);
or U2547 (N_2547,In_1463,In_633);
or U2548 (N_2548,In_1399,In_1216);
or U2549 (N_2549,In_690,In_899);
and U2550 (N_2550,In_702,In_12);
nand U2551 (N_2551,In_742,In_987);
nand U2552 (N_2552,In_959,In_408);
and U2553 (N_2553,In_813,In_20);
and U2554 (N_2554,In_1408,In_1474);
nand U2555 (N_2555,In_652,In_258);
nor U2556 (N_2556,In_1303,In_763);
nand U2557 (N_2557,In_433,In_647);
nand U2558 (N_2558,In_282,In_376);
and U2559 (N_2559,In_364,In_865);
and U2560 (N_2560,In_1191,In_76);
nor U2561 (N_2561,In_1242,In_291);
and U2562 (N_2562,In_220,In_725);
nor U2563 (N_2563,In_62,In_709);
nand U2564 (N_2564,In_939,In_949);
nand U2565 (N_2565,In_493,In_285);
and U2566 (N_2566,In_1070,In_645);
nand U2567 (N_2567,In_501,In_1245);
and U2568 (N_2568,In_469,In_377);
nand U2569 (N_2569,In_225,In_1417);
nand U2570 (N_2570,In_282,In_1125);
and U2571 (N_2571,In_725,In_919);
and U2572 (N_2572,In_1038,In_1477);
nand U2573 (N_2573,In_543,In_24);
nor U2574 (N_2574,In_1010,In_471);
or U2575 (N_2575,In_33,In_85);
nand U2576 (N_2576,In_866,In_597);
nor U2577 (N_2577,In_1088,In_594);
and U2578 (N_2578,In_886,In_1486);
and U2579 (N_2579,In_1212,In_724);
or U2580 (N_2580,In_1381,In_1321);
and U2581 (N_2581,In_1440,In_349);
or U2582 (N_2582,In_1248,In_1033);
nor U2583 (N_2583,In_147,In_21);
nor U2584 (N_2584,In_1013,In_1095);
nand U2585 (N_2585,In_489,In_838);
nand U2586 (N_2586,In_800,In_5);
nor U2587 (N_2587,In_1174,In_522);
or U2588 (N_2588,In_1377,In_121);
nand U2589 (N_2589,In_332,In_746);
and U2590 (N_2590,In_875,In_1460);
nand U2591 (N_2591,In_639,In_1055);
or U2592 (N_2592,In_423,In_1396);
and U2593 (N_2593,In_962,In_1173);
and U2594 (N_2594,In_413,In_384);
and U2595 (N_2595,In_758,In_173);
or U2596 (N_2596,In_1307,In_1234);
nand U2597 (N_2597,In_1079,In_422);
and U2598 (N_2598,In_87,In_876);
or U2599 (N_2599,In_448,In_697);
or U2600 (N_2600,In_1384,In_146);
or U2601 (N_2601,In_532,In_641);
nand U2602 (N_2602,In_1275,In_1131);
and U2603 (N_2603,In_127,In_208);
and U2604 (N_2604,In_1132,In_498);
nor U2605 (N_2605,In_795,In_602);
nand U2606 (N_2606,In_579,In_1248);
or U2607 (N_2607,In_1040,In_1342);
nor U2608 (N_2608,In_745,In_1423);
nand U2609 (N_2609,In_228,In_525);
and U2610 (N_2610,In_128,In_76);
nor U2611 (N_2611,In_673,In_116);
nand U2612 (N_2612,In_1352,In_1046);
or U2613 (N_2613,In_900,In_24);
nor U2614 (N_2614,In_1017,In_263);
or U2615 (N_2615,In_286,In_1174);
nand U2616 (N_2616,In_1090,In_1134);
or U2617 (N_2617,In_867,In_59);
and U2618 (N_2618,In_1372,In_85);
nand U2619 (N_2619,In_527,In_104);
or U2620 (N_2620,In_1177,In_738);
nand U2621 (N_2621,In_909,In_1226);
xnor U2622 (N_2622,In_1076,In_593);
nor U2623 (N_2623,In_82,In_694);
nand U2624 (N_2624,In_855,In_263);
nand U2625 (N_2625,In_496,In_340);
and U2626 (N_2626,In_285,In_338);
nand U2627 (N_2627,In_461,In_698);
or U2628 (N_2628,In_1065,In_1376);
and U2629 (N_2629,In_1355,In_992);
and U2630 (N_2630,In_549,In_1429);
or U2631 (N_2631,In_1259,In_149);
or U2632 (N_2632,In_1331,In_376);
nor U2633 (N_2633,In_1212,In_644);
nor U2634 (N_2634,In_505,In_1098);
and U2635 (N_2635,In_395,In_933);
nand U2636 (N_2636,In_885,In_402);
nor U2637 (N_2637,In_884,In_621);
or U2638 (N_2638,In_1248,In_867);
nand U2639 (N_2639,In_775,In_157);
nor U2640 (N_2640,In_1183,In_611);
nand U2641 (N_2641,In_1236,In_1370);
or U2642 (N_2642,In_206,In_800);
nand U2643 (N_2643,In_266,In_1201);
nor U2644 (N_2644,In_1139,In_187);
nor U2645 (N_2645,In_16,In_637);
and U2646 (N_2646,In_1207,In_979);
nor U2647 (N_2647,In_146,In_418);
or U2648 (N_2648,In_434,In_383);
nand U2649 (N_2649,In_13,In_144);
or U2650 (N_2650,In_473,In_756);
nand U2651 (N_2651,In_202,In_965);
and U2652 (N_2652,In_1139,In_407);
or U2653 (N_2653,In_771,In_324);
and U2654 (N_2654,In_112,In_848);
and U2655 (N_2655,In_73,In_764);
nor U2656 (N_2656,In_802,In_431);
xnor U2657 (N_2657,In_918,In_1117);
and U2658 (N_2658,In_1208,In_379);
and U2659 (N_2659,In_460,In_182);
or U2660 (N_2660,In_1463,In_295);
or U2661 (N_2661,In_292,In_713);
nand U2662 (N_2662,In_524,In_90);
or U2663 (N_2663,In_784,In_1122);
or U2664 (N_2664,In_676,In_581);
nand U2665 (N_2665,In_547,In_1119);
nand U2666 (N_2666,In_203,In_110);
and U2667 (N_2667,In_694,In_1168);
nor U2668 (N_2668,In_463,In_1209);
or U2669 (N_2669,In_838,In_351);
nand U2670 (N_2670,In_1102,In_1022);
nand U2671 (N_2671,In_965,In_818);
nand U2672 (N_2672,In_1460,In_509);
and U2673 (N_2673,In_1179,In_566);
nand U2674 (N_2674,In_470,In_1082);
and U2675 (N_2675,In_699,In_687);
or U2676 (N_2676,In_1455,In_78);
and U2677 (N_2677,In_992,In_1061);
or U2678 (N_2678,In_1388,In_765);
nand U2679 (N_2679,In_886,In_304);
nand U2680 (N_2680,In_928,In_341);
or U2681 (N_2681,In_454,In_8);
and U2682 (N_2682,In_1008,In_1024);
nand U2683 (N_2683,In_380,In_767);
nand U2684 (N_2684,In_787,In_392);
xor U2685 (N_2685,In_1037,In_273);
nor U2686 (N_2686,In_850,In_845);
and U2687 (N_2687,In_1483,In_1263);
or U2688 (N_2688,In_1407,In_1425);
nand U2689 (N_2689,In_1162,In_605);
nand U2690 (N_2690,In_248,In_867);
and U2691 (N_2691,In_505,In_781);
nand U2692 (N_2692,In_697,In_1083);
nand U2693 (N_2693,In_33,In_603);
and U2694 (N_2694,In_492,In_669);
or U2695 (N_2695,In_1123,In_602);
or U2696 (N_2696,In_1458,In_265);
and U2697 (N_2697,In_1247,In_402);
and U2698 (N_2698,In_32,In_590);
nand U2699 (N_2699,In_471,In_789);
and U2700 (N_2700,In_398,In_1358);
or U2701 (N_2701,In_1040,In_991);
nand U2702 (N_2702,In_1339,In_1210);
and U2703 (N_2703,In_310,In_101);
nand U2704 (N_2704,In_243,In_57);
and U2705 (N_2705,In_263,In_628);
nand U2706 (N_2706,In_1023,In_1429);
or U2707 (N_2707,In_1277,In_1003);
nand U2708 (N_2708,In_350,In_271);
nor U2709 (N_2709,In_1135,In_1306);
nand U2710 (N_2710,In_484,In_124);
nor U2711 (N_2711,In_280,In_236);
nand U2712 (N_2712,In_1163,In_1056);
xor U2713 (N_2713,In_390,In_487);
nor U2714 (N_2714,In_1149,In_1020);
nor U2715 (N_2715,In_665,In_1073);
or U2716 (N_2716,In_492,In_73);
nor U2717 (N_2717,In_114,In_335);
nand U2718 (N_2718,In_600,In_970);
or U2719 (N_2719,In_1118,In_836);
nor U2720 (N_2720,In_520,In_1400);
nor U2721 (N_2721,In_995,In_37);
nand U2722 (N_2722,In_723,In_602);
nor U2723 (N_2723,In_425,In_991);
and U2724 (N_2724,In_1028,In_435);
nand U2725 (N_2725,In_1270,In_480);
and U2726 (N_2726,In_144,In_969);
or U2727 (N_2727,In_1433,In_558);
nor U2728 (N_2728,In_533,In_545);
nor U2729 (N_2729,In_263,In_1255);
nor U2730 (N_2730,In_963,In_151);
nand U2731 (N_2731,In_1053,In_870);
and U2732 (N_2732,In_810,In_1402);
or U2733 (N_2733,In_313,In_1055);
nand U2734 (N_2734,In_495,In_841);
and U2735 (N_2735,In_1279,In_689);
and U2736 (N_2736,In_421,In_1421);
or U2737 (N_2737,In_851,In_1315);
or U2738 (N_2738,In_908,In_527);
nand U2739 (N_2739,In_1064,In_1022);
or U2740 (N_2740,In_1478,In_1441);
and U2741 (N_2741,In_326,In_544);
nand U2742 (N_2742,In_1359,In_863);
nor U2743 (N_2743,In_983,In_1295);
nand U2744 (N_2744,In_1364,In_759);
or U2745 (N_2745,In_1434,In_529);
and U2746 (N_2746,In_481,In_208);
and U2747 (N_2747,In_1237,In_1473);
and U2748 (N_2748,In_6,In_361);
or U2749 (N_2749,In_531,In_1204);
xnor U2750 (N_2750,In_528,In_416);
nand U2751 (N_2751,In_1482,In_487);
or U2752 (N_2752,In_798,In_64);
nor U2753 (N_2753,In_492,In_1189);
nand U2754 (N_2754,In_329,In_447);
nand U2755 (N_2755,In_262,In_325);
nor U2756 (N_2756,In_1365,In_118);
and U2757 (N_2757,In_751,In_652);
nor U2758 (N_2758,In_1449,In_1241);
or U2759 (N_2759,In_326,In_192);
nand U2760 (N_2760,In_3,In_434);
nand U2761 (N_2761,In_1321,In_954);
nand U2762 (N_2762,In_1051,In_1151);
nor U2763 (N_2763,In_1115,In_1326);
or U2764 (N_2764,In_131,In_1326);
nand U2765 (N_2765,In_641,In_806);
or U2766 (N_2766,In_528,In_773);
nor U2767 (N_2767,In_670,In_800);
or U2768 (N_2768,In_308,In_421);
and U2769 (N_2769,In_1495,In_687);
nand U2770 (N_2770,In_545,In_443);
and U2771 (N_2771,In_1173,In_1064);
nor U2772 (N_2772,In_1040,In_300);
nor U2773 (N_2773,In_507,In_575);
nand U2774 (N_2774,In_936,In_327);
nor U2775 (N_2775,In_164,In_842);
xnor U2776 (N_2776,In_1476,In_252);
and U2777 (N_2777,In_717,In_940);
xor U2778 (N_2778,In_1346,In_1007);
xnor U2779 (N_2779,In_701,In_905);
and U2780 (N_2780,In_951,In_511);
nand U2781 (N_2781,In_1008,In_248);
nor U2782 (N_2782,In_711,In_147);
and U2783 (N_2783,In_987,In_1045);
and U2784 (N_2784,In_1350,In_815);
or U2785 (N_2785,In_1212,In_1498);
or U2786 (N_2786,In_1002,In_1010);
xor U2787 (N_2787,In_903,In_736);
nand U2788 (N_2788,In_1461,In_372);
or U2789 (N_2789,In_29,In_1408);
or U2790 (N_2790,In_989,In_856);
nor U2791 (N_2791,In_874,In_855);
or U2792 (N_2792,In_1454,In_269);
and U2793 (N_2793,In_529,In_1237);
nor U2794 (N_2794,In_1329,In_191);
xnor U2795 (N_2795,In_422,In_289);
nor U2796 (N_2796,In_713,In_726);
and U2797 (N_2797,In_722,In_1347);
and U2798 (N_2798,In_704,In_863);
nor U2799 (N_2799,In_639,In_1);
or U2800 (N_2800,In_230,In_1367);
and U2801 (N_2801,In_103,In_960);
or U2802 (N_2802,In_828,In_1012);
nand U2803 (N_2803,In_1332,In_943);
nand U2804 (N_2804,In_776,In_1021);
nor U2805 (N_2805,In_1461,In_1107);
nand U2806 (N_2806,In_658,In_656);
nand U2807 (N_2807,In_715,In_926);
nand U2808 (N_2808,In_1259,In_456);
or U2809 (N_2809,In_114,In_264);
nand U2810 (N_2810,In_716,In_375);
nor U2811 (N_2811,In_728,In_1367);
and U2812 (N_2812,In_934,In_577);
and U2813 (N_2813,In_1497,In_408);
or U2814 (N_2814,In_967,In_143);
nor U2815 (N_2815,In_832,In_811);
nand U2816 (N_2816,In_255,In_1165);
or U2817 (N_2817,In_900,In_711);
nor U2818 (N_2818,In_1410,In_523);
or U2819 (N_2819,In_393,In_1491);
nand U2820 (N_2820,In_906,In_390);
nor U2821 (N_2821,In_1270,In_1004);
and U2822 (N_2822,In_882,In_430);
nor U2823 (N_2823,In_791,In_1348);
and U2824 (N_2824,In_855,In_869);
nand U2825 (N_2825,In_1015,In_197);
and U2826 (N_2826,In_927,In_1227);
or U2827 (N_2827,In_893,In_1304);
or U2828 (N_2828,In_1060,In_735);
nand U2829 (N_2829,In_1387,In_486);
or U2830 (N_2830,In_565,In_1133);
and U2831 (N_2831,In_901,In_455);
nor U2832 (N_2832,In_205,In_240);
and U2833 (N_2833,In_379,In_1442);
nor U2834 (N_2834,In_551,In_1224);
nor U2835 (N_2835,In_1491,In_609);
nor U2836 (N_2836,In_898,In_421);
nand U2837 (N_2837,In_11,In_1416);
or U2838 (N_2838,In_1294,In_1169);
nand U2839 (N_2839,In_1374,In_887);
nor U2840 (N_2840,In_1122,In_589);
and U2841 (N_2841,In_1441,In_453);
or U2842 (N_2842,In_978,In_689);
nand U2843 (N_2843,In_1155,In_833);
or U2844 (N_2844,In_253,In_576);
and U2845 (N_2845,In_485,In_235);
nor U2846 (N_2846,In_1250,In_428);
nand U2847 (N_2847,In_1337,In_995);
or U2848 (N_2848,In_553,In_479);
and U2849 (N_2849,In_993,In_1207);
nor U2850 (N_2850,In_161,In_1003);
nand U2851 (N_2851,In_1400,In_1351);
nor U2852 (N_2852,In_84,In_917);
nor U2853 (N_2853,In_1282,In_594);
or U2854 (N_2854,In_748,In_566);
or U2855 (N_2855,In_1075,In_1214);
nand U2856 (N_2856,In_1303,In_1489);
nand U2857 (N_2857,In_516,In_1094);
nor U2858 (N_2858,In_803,In_387);
and U2859 (N_2859,In_1155,In_1202);
nand U2860 (N_2860,In_1295,In_1427);
nand U2861 (N_2861,In_600,In_544);
nand U2862 (N_2862,In_1302,In_1457);
nor U2863 (N_2863,In_234,In_1331);
or U2864 (N_2864,In_75,In_1168);
or U2865 (N_2865,In_194,In_493);
and U2866 (N_2866,In_1190,In_866);
and U2867 (N_2867,In_1249,In_1377);
and U2868 (N_2868,In_1091,In_22);
and U2869 (N_2869,In_252,In_320);
or U2870 (N_2870,In_968,In_550);
nand U2871 (N_2871,In_1157,In_578);
nand U2872 (N_2872,In_207,In_696);
nand U2873 (N_2873,In_1478,In_1499);
nor U2874 (N_2874,In_252,In_1343);
and U2875 (N_2875,In_345,In_174);
or U2876 (N_2876,In_470,In_1270);
nand U2877 (N_2877,In_809,In_18);
nor U2878 (N_2878,In_11,In_1084);
nor U2879 (N_2879,In_202,In_1287);
or U2880 (N_2880,In_812,In_1436);
xnor U2881 (N_2881,In_1353,In_66);
nand U2882 (N_2882,In_1414,In_377);
nand U2883 (N_2883,In_148,In_628);
nor U2884 (N_2884,In_181,In_427);
or U2885 (N_2885,In_241,In_380);
nor U2886 (N_2886,In_1086,In_954);
nor U2887 (N_2887,In_470,In_596);
or U2888 (N_2888,In_1180,In_1198);
and U2889 (N_2889,In_1269,In_1369);
or U2890 (N_2890,In_868,In_354);
or U2891 (N_2891,In_62,In_1495);
nor U2892 (N_2892,In_647,In_1204);
nand U2893 (N_2893,In_1249,In_1217);
and U2894 (N_2894,In_731,In_543);
nor U2895 (N_2895,In_1367,In_1330);
or U2896 (N_2896,In_1290,In_1474);
or U2897 (N_2897,In_549,In_297);
nand U2898 (N_2898,In_705,In_117);
and U2899 (N_2899,In_35,In_758);
nor U2900 (N_2900,In_500,In_39);
nand U2901 (N_2901,In_868,In_639);
and U2902 (N_2902,In_2,In_990);
nor U2903 (N_2903,In_905,In_586);
or U2904 (N_2904,In_757,In_578);
and U2905 (N_2905,In_648,In_58);
nand U2906 (N_2906,In_1077,In_738);
or U2907 (N_2907,In_1182,In_1430);
nor U2908 (N_2908,In_1128,In_698);
nor U2909 (N_2909,In_848,In_194);
xor U2910 (N_2910,In_726,In_1261);
xnor U2911 (N_2911,In_189,In_824);
nand U2912 (N_2912,In_1124,In_242);
nand U2913 (N_2913,In_931,In_574);
or U2914 (N_2914,In_887,In_1425);
nand U2915 (N_2915,In_926,In_845);
nor U2916 (N_2916,In_1115,In_1130);
and U2917 (N_2917,In_1262,In_621);
or U2918 (N_2918,In_875,In_1034);
nor U2919 (N_2919,In_372,In_868);
nor U2920 (N_2920,In_152,In_96);
nand U2921 (N_2921,In_218,In_1073);
nor U2922 (N_2922,In_1445,In_315);
nor U2923 (N_2923,In_1400,In_1167);
and U2924 (N_2924,In_285,In_220);
nor U2925 (N_2925,In_853,In_826);
nor U2926 (N_2926,In_632,In_435);
or U2927 (N_2927,In_349,In_1185);
xnor U2928 (N_2928,In_819,In_1276);
or U2929 (N_2929,In_1156,In_958);
or U2930 (N_2930,In_941,In_1222);
nor U2931 (N_2931,In_1188,In_1247);
and U2932 (N_2932,In_547,In_762);
and U2933 (N_2933,In_71,In_1192);
nand U2934 (N_2934,In_1384,In_144);
and U2935 (N_2935,In_400,In_29);
nor U2936 (N_2936,In_865,In_783);
or U2937 (N_2937,In_433,In_1090);
nor U2938 (N_2938,In_75,In_10);
and U2939 (N_2939,In_490,In_189);
or U2940 (N_2940,In_9,In_1094);
nand U2941 (N_2941,In_144,In_902);
and U2942 (N_2942,In_1261,In_1250);
nand U2943 (N_2943,In_1089,In_310);
and U2944 (N_2944,In_477,In_798);
and U2945 (N_2945,In_1070,In_1272);
nand U2946 (N_2946,In_313,In_934);
nor U2947 (N_2947,In_1412,In_538);
and U2948 (N_2948,In_1310,In_419);
nor U2949 (N_2949,In_336,In_692);
nor U2950 (N_2950,In_159,In_381);
or U2951 (N_2951,In_1119,In_33);
or U2952 (N_2952,In_1463,In_38);
or U2953 (N_2953,In_1200,In_1047);
or U2954 (N_2954,In_1097,In_157);
nand U2955 (N_2955,In_965,In_354);
and U2956 (N_2956,In_1255,In_384);
and U2957 (N_2957,In_3,In_653);
or U2958 (N_2958,In_841,In_1224);
and U2959 (N_2959,In_576,In_911);
or U2960 (N_2960,In_1450,In_150);
nor U2961 (N_2961,In_1171,In_854);
or U2962 (N_2962,In_671,In_1188);
nand U2963 (N_2963,In_277,In_196);
and U2964 (N_2964,In_623,In_243);
nor U2965 (N_2965,In_408,In_1316);
nand U2966 (N_2966,In_202,In_493);
nand U2967 (N_2967,In_851,In_1266);
xnor U2968 (N_2968,In_811,In_534);
nand U2969 (N_2969,In_855,In_933);
nor U2970 (N_2970,In_469,In_699);
nand U2971 (N_2971,In_1287,In_1464);
or U2972 (N_2972,In_914,In_1434);
or U2973 (N_2973,In_581,In_1335);
nor U2974 (N_2974,In_930,In_380);
or U2975 (N_2975,In_1377,In_1358);
nor U2976 (N_2976,In_682,In_516);
nand U2977 (N_2977,In_377,In_984);
nand U2978 (N_2978,In_967,In_469);
nor U2979 (N_2979,In_1111,In_1282);
xnor U2980 (N_2980,In_860,In_1374);
or U2981 (N_2981,In_276,In_370);
or U2982 (N_2982,In_1038,In_389);
nand U2983 (N_2983,In_1484,In_947);
or U2984 (N_2984,In_472,In_1042);
nor U2985 (N_2985,In_1134,In_412);
nor U2986 (N_2986,In_598,In_956);
nand U2987 (N_2987,In_822,In_1);
and U2988 (N_2988,In_950,In_811);
or U2989 (N_2989,In_1455,In_776);
nor U2990 (N_2990,In_1186,In_818);
nand U2991 (N_2991,In_1340,In_592);
nor U2992 (N_2992,In_19,In_597);
nor U2993 (N_2993,In_1427,In_455);
nor U2994 (N_2994,In_424,In_508);
and U2995 (N_2995,In_1375,In_347);
and U2996 (N_2996,In_1113,In_116);
xnor U2997 (N_2997,In_958,In_735);
nor U2998 (N_2998,In_442,In_900);
nor U2999 (N_2999,In_884,In_425);
and U3000 (N_3000,N_623,N_1758);
xor U3001 (N_3001,N_2612,N_1877);
or U3002 (N_3002,N_2770,N_2055);
and U3003 (N_3003,N_1253,N_1786);
xnor U3004 (N_3004,N_2877,N_2762);
nand U3005 (N_3005,N_2126,N_1885);
nand U3006 (N_3006,N_414,N_2318);
nor U3007 (N_3007,N_1398,N_396);
and U3008 (N_3008,N_2480,N_2385);
and U3009 (N_3009,N_1144,N_1052);
and U3010 (N_3010,N_2304,N_46);
nor U3011 (N_3011,N_2493,N_209);
or U3012 (N_3012,N_2212,N_2758);
nor U3013 (N_3013,N_2907,N_1345);
and U3014 (N_3014,N_326,N_340);
or U3015 (N_3015,N_43,N_2004);
and U3016 (N_3016,N_840,N_2672);
and U3017 (N_3017,N_1826,N_257);
nand U3018 (N_3018,N_410,N_2699);
and U3019 (N_3019,N_188,N_1640);
and U3020 (N_3020,N_1905,N_214);
or U3021 (N_3021,N_1598,N_1392);
xor U3022 (N_3022,N_138,N_1866);
and U3023 (N_3023,N_2873,N_1651);
or U3024 (N_3024,N_1523,N_2765);
nand U3025 (N_3025,N_848,N_2081);
and U3026 (N_3026,N_1634,N_1703);
or U3027 (N_3027,N_1125,N_2157);
nor U3028 (N_3028,N_858,N_1802);
nand U3029 (N_3029,N_1372,N_1024);
and U3030 (N_3030,N_1935,N_2146);
nor U3031 (N_3031,N_2627,N_1136);
or U3032 (N_3032,N_694,N_2373);
nand U3033 (N_3033,N_1113,N_1727);
and U3034 (N_3034,N_2162,N_2987);
nand U3035 (N_3035,N_1278,N_2053);
nor U3036 (N_3036,N_2848,N_722);
and U3037 (N_3037,N_2705,N_1030);
nor U3038 (N_3038,N_85,N_2869);
and U3039 (N_3039,N_1603,N_428);
nor U3040 (N_3040,N_2648,N_1124);
nand U3041 (N_3041,N_1035,N_823);
or U3042 (N_3042,N_2664,N_1776);
nand U3043 (N_3043,N_531,N_2909);
and U3044 (N_3044,N_1536,N_358);
or U3045 (N_3045,N_2076,N_2694);
nand U3046 (N_3046,N_1022,N_1464);
and U3047 (N_3047,N_1586,N_2471);
nand U3048 (N_3048,N_1956,N_853);
nor U3049 (N_3049,N_2125,N_1131);
and U3050 (N_3050,N_1244,N_1314);
nand U3051 (N_3051,N_2851,N_930);
nand U3052 (N_3052,N_966,N_2898);
nor U3053 (N_3053,N_2087,N_1737);
xor U3054 (N_3054,N_1105,N_2271);
or U3055 (N_3055,N_2130,N_1316);
and U3056 (N_3056,N_2936,N_2388);
or U3057 (N_3057,N_2794,N_588);
nor U3058 (N_3058,N_1209,N_913);
and U3059 (N_3059,N_2001,N_2514);
and U3060 (N_3060,N_1752,N_2095);
and U3061 (N_3061,N_305,N_1241);
and U3062 (N_3062,N_2623,N_1694);
or U3063 (N_3063,N_1638,N_1397);
or U3064 (N_3064,N_1978,N_2177);
and U3065 (N_3065,N_2943,N_24);
nor U3066 (N_3066,N_2738,N_2143);
nor U3067 (N_3067,N_9,N_1734);
nor U3068 (N_3068,N_1138,N_141);
and U3069 (N_3069,N_1960,N_2844);
or U3070 (N_3070,N_1225,N_364);
or U3071 (N_3071,N_118,N_468);
nor U3072 (N_3072,N_2719,N_1544);
nor U3073 (N_3073,N_1863,N_2860);
nor U3074 (N_3074,N_1891,N_77);
nand U3075 (N_3075,N_826,N_2656);
or U3076 (N_3076,N_1782,N_816);
or U3077 (N_3077,N_2194,N_516);
or U3078 (N_3078,N_1573,N_1515);
nand U3079 (N_3079,N_543,N_674);
or U3080 (N_3080,N_782,N_986);
nand U3081 (N_3081,N_1516,N_573);
nand U3082 (N_3082,N_1875,N_1331);
or U3083 (N_3083,N_1618,N_746);
nor U3084 (N_3084,N_1182,N_2747);
nor U3085 (N_3085,N_618,N_2599);
nor U3086 (N_3086,N_160,N_2206);
nor U3087 (N_3087,N_453,N_2611);
nor U3088 (N_3088,N_605,N_942);
nor U3089 (N_3089,N_492,N_558);
or U3090 (N_3090,N_2715,N_949);
nor U3091 (N_3091,N_459,N_1981);
and U3092 (N_3092,N_1028,N_1551);
or U3093 (N_3093,N_748,N_1277);
nor U3094 (N_3094,N_830,N_2435);
nand U3095 (N_3095,N_2755,N_1);
nor U3096 (N_3096,N_2215,N_2812);
nor U3097 (N_3097,N_733,N_2193);
nand U3098 (N_3098,N_788,N_524);
and U3099 (N_3099,N_2655,N_2988);
and U3100 (N_3100,N_1477,N_1977);
and U3101 (N_3101,N_2098,N_1655);
or U3102 (N_3102,N_1092,N_2740);
nor U3103 (N_3103,N_2297,N_1221);
or U3104 (N_3104,N_1134,N_1079);
xnor U3105 (N_3105,N_2298,N_520);
or U3106 (N_3106,N_1949,N_1567);
nand U3107 (N_3107,N_477,N_1025);
or U3108 (N_3108,N_1625,N_2264);
nand U3109 (N_3109,N_1993,N_435);
nor U3110 (N_3110,N_2312,N_1728);
nor U3111 (N_3111,N_1608,N_947);
nor U3112 (N_3112,N_1527,N_2827);
or U3113 (N_3113,N_801,N_1165);
nand U3114 (N_3114,N_1672,N_1157);
nor U3115 (N_3115,N_2077,N_1133);
and U3116 (N_3116,N_1502,N_2859);
and U3117 (N_3117,N_2631,N_1713);
or U3118 (N_3118,N_881,N_1961);
nand U3119 (N_3119,N_624,N_344);
or U3120 (N_3120,N_1393,N_756);
and U3121 (N_3121,N_2613,N_415);
nor U3122 (N_3122,N_298,N_2016);
nor U3123 (N_3123,N_2543,N_1274);
and U3124 (N_3124,N_39,N_1000);
or U3125 (N_3125,N_2536,N_1285);
and U3126 (N_3126,N_1389,N_1992);
nand U3127 (N_3127,N_1198,N_81);
nand U3128 (N_3128,N_394,N_370);
nand U3129 (N_3129,N_1499,N_855);
or U3130 (N_3130,N_1853,N_2107);
or U3131 (N_3131,N_646,N_2785);
or U3132 (N_3132,N_2201,N_937);
or U3133 (N_3133,N_1449,N_661);
and U3134 (N_3134,N_2069,N_652);
nor U3135 (N_3135,N_354,N_2695);
and U3136 (N_3136,N_880,N_210);
and U3137 (N_3137,N_925,N_395);
and U3138 (N_3138,N_476,N_2129);
or U3139 (N_3139,N_452,N_556);
or U3140 (N_3140,N_1391,N_2377);
nand U3141 (N_3141,N_1964,N_2176);
nand U3142 (N_3142,N_967,N_1864);
and U3143 (N_3143,N_263,N_248);
and U3144 (N_3144,N_131,N_2414);
nand U3145 (N_3145,N_515,N_1036);
and U3146 (N_3146,N_1078,N_1310);
nand U3147 (N_3147,N_334,N_2403);
nand U3148 (N_3148,N_2222,N_1458);
and U3149 (N_3149,N_1649,N_1809);
and U3150 (N_3150,N_2729,N_332);
or U3151 (N_3151,N_1303,N_1525);
nor U3152 (N_3152,N_1470,N_662);
nor U3153 (N_3153,N_2238,N_1560);
nor U3154 (N_3154,N_1018,N_125);
nor U3155 (N_3155,N_1216,N_1064);
and U3156 (N_3156,N_1266,N_1558);
or U3157 (N_3157,N_2019,N_2432);
nor U3158 (N_3158,N_2818,N_1243);
nand U3159 (N_3159,N_1411,N_2195);
nand U3160 (N_3160,N_2286,N_1942);
nand U3161 (N_3161,N_2856,N_2287);
or U3162 (N_3162,N_1669,N_2587);
and U3163 (N_3163,N_451,N_2398);
and U3164 (N_3164,N_1210,N_953);
nand U3165 (N_3165,N_176,N_383);
or U3166 (N_3166,N_1417,N_1287);
and U3167 (N_3167,N_2996,N_2457);
and U3168 (N_3168,N_1119,N_2084);
and U3169 (N_3169,N_2576,N_362);
and U3170 (N_3170,N_2119,N_1682);
xor U3171 (N_3171,N_2824,N_831);
or U3172 (N_3172,N_2717,N_1980);
nor U3173 (N_3173,N_1947,N_2982);
and U3174 (N_3174,N_962,N_711);
nand U3175 (N_3175,N_551,N_2307);
or U3176 (N_3176,N_2736,N_2905);
nor U3177 (N_3177,N_2014,N_973);
or U3178 (N_3178,N_835,N_2769);
and U3179 (N_3179,N_1091,N_1187);
nand U3180 (N_3180,N_2990,N_2911);
nor U3181 (N_3181,N_1719,N_1653);
nor U3182 (N_3182,N_760,N_2608);
or U3183 (N_3183,N_2440,N_625);
nor U3184 (N_3184,N_1347,N_2497);
nand U3185 (N_3185,N_2991,N_2380);
nor U3186 (N_3186,N_2487,N_1341);
and U3187 (N_3187,N_2746,N_1468);
nor U3188 (N_3188,N_2556,N_1535);
nor U3189 (N_3189,N_282,N_1171);
nor U3190 (N_3190,N_224,N_2293);
xor U3191 (N_3191,N_204,N_2949);
and U3192 (N_3192,N_817,N_235);
or U3193 (N_3193,N_2389,N_2788);
and U3194 (N_3194,N_2914,N_2506);
or U3195 (N_3195,N_1997,N_136);
nand U3196 (N_3196,N_898,N_1858);
nor U3197 (N_3197,N_2775,N_634);
nand U3198 (N_3198,N_2722,N_432);
or U3199 (N_3199,N_1466,N_1821);
nor U3200 (N_3200,N_2867,N_1881);
and U3201 (N_3201,N_2115,N_976);
and U3202 (N_3202,N_1270,N_970);
and U3203 (N_3203,N_498,N_2647);
or U3204 (N_3204,N_1944,N_388);
nand U3205 (N_3205,N_2583,N_750);
nand U3206 (N_3206,N_1365,N_1305);
nand U3207 (N_3207,N_806,N_1869);
xor U3208 (N_3208,N_2463,N_1697);
nor U3209 (N_3209,N_1912,N_91);
or U3210 (N_3210,N_2408,N_314);
and U3211 (N_3211,N_2972,N_1434);
nor U3212 (N_3212,N_959,N_1931);
nor U3213 (N_3213,N_2340,N_265);
nor U3214 (N_3214,N_1808,N_2674);
and U3215 (N_3215,N_2744,N_2650);
and U3216 (N_3216,N_2123,N_83);
nor U3217 (N_3217,N_574,N_1600);
nand U3218 (N_3218,N_54,N_2295);
nor U3219 (N_3219,N_1054,N_1259);
and U3220 (N_3220,N_1780,N_931);
and U3221 (N_3221,N_401,N_495);
and U3222 (N_3222,N_339,N_397);
and U3223 (N_3223,N_1939,N_17);
nor U3224 (N_3224,N_747,N_2690);
nand U3225 (N_3225,N_387,N_1901);
or U3226 (N_3226,N_1862,N_2434);
or U3227 (N_3227,N_2845,N_1907);
and U3228 (N_3228,N_206,N_659);
nand U3229 (N_3229,N_743,N_56);
and U3230 (N_3230,N_1539,N_596);
or U3231 (N_3231,N_96,N_640);
nand U3232 (N_3232,N_940,N_1142);
nor U3233 (N_3233,N_2468,N_599);
nand U3234 (N_3234,N_1899,N_645);
and U3235 (N_3235,N_2742,N_2062);
nor U3236 (N_3236,N_800,N_669);
nor U3237 (N_3237,N_761,N_2154);
and U3238 (N_3238,N_450,N_1557);
nand U3239 (N_3239,N_1888,N_147);
nor U3240 (N_3240,N_2839,N_1548);
and U3241 (N_3241,N_984,N_1192);
nor U3242 (N_3242,N_2394,N_1718);
or U3243 (N_3243,N_2624,N_114);
nor U3244 (N_3244,N_1708,N_2103);
nor U3245 (N_3245,N_1002,N_2444);
xor U3246 (N_3246,N_1685,N_302);
nor U3247 (N_3247,N_1609,N_1246);
and U3248 (N_3248,N_155,N_2396);
or U3249 (N_3249,N_1626,N_827);
nand U3250 (N_3250,N_704,N_2692);
nor U3251 (N_3251,N_208,N_927);
and U3252 (N_3252,N_2605,N_2498);
or U3253 (N_3253,N_1333,N_1771);
and U3254 (N_3254,N_1787,N_2523);
or U3255 (N_3255,N_1568,N_1941);
nor U3256 (N_3256,N_1810,N_1205);
and U3257 (N_3257,N_2252,N_1958);
and U3258 (N_3258,N_1631,N_73);
nand U3259 (N_3259,N_412,N_179);
nor U3260 (N_3260,N_2508,N_2709);
nor U3261 (N_3261,N_371,N_2120);
and U3262 (N_3262,N_923,N_2870);
nand U3263 (N_3263,N_2961,N_1486);
nor U3264 (N_3264,N_169,N_2895);
and U3265 (N_3265,N_2227,N_580);
nand U3266 (N_3266,N_2501,N_903);
nand U3267 (N_3267,N_1596,N_725);
nor U3268 (N_3268,N_2888,N_779);
nand U3269 (N_3269,N_709,N_2622);
nor U3270 (N_3270,N_995,N_2853);
nand U3271 (N_3271,N_1705,N_1739);
and U3272 (N_3272,N_1985,N_977);
nor U3273 (N_3273,N_469,N_2512);
or U3274 (N_3274,N_245,N_442);
and U3275 (N_3275,N_69,N_2537);
and U3276 (N_3276,N_2223,N_2864);
or U3277 (N_3277,N_668,N_509);
nand U3278 (N_3278,N_1433,N_2550);
nand U3279 (N_3279,N_505,N_1431);
nand U3280 (N_3280,N_869,N_1237);
nor U3281 (N_3281,N_1355,N_744);
and U3282 (N_3282,N_1096,N_2447);
nand U3283 (N_3283,N_1623,N_2302);
nor U3284 (N_3284,N_1204,N_2787);
xnor U3285 (N_3285,N_365,N_207);
and U3286 (N_3286,N_1057,N_71);
or U3287 (N_3287,N_1818,N_2181);
or U3288 (N_3288,N_2791,N_1356);
nand U3289 (N_3289,N_1267,N_378);
nor U3290 (N_3290,N_1185,N_534);
and U3291 (N_3291,N_1166,N_1293);
nor U3292 (N_3292,N_2391,N_2980);
or U3293 (N_3293,N_974,N_2525);
and U3294 (N_3294,N_1994,N_281);
and U3295 (N_3295,N_2216,N_2828);
nor U3296 (N_3296,N_856,N_1589);
xor U3297 (N_3297,N_2757,N_10);
nor U3298 (N_3298,N_1349,N_1822);
and U3299 (N_3299,N_2042,N_2721);
and U3300 (N_3300,N_161,N_491);
or U3301 (N_3301,N_1212,N_1473);
and U3302 (N_3302,N_2606,N_1563);
or U3303 (N_3303,N_643,N_1461);
nor U3304 (N_3304,N_2731,N_2561);
or U3305 (N_3305,N_1616,N_2696);
nand U3306 (N_3306,N_764,N_1399);
nor U3307 (N_3307,N_2118,N_2687);
nor U3308 (N_3308,N_1413,N_2494);
or U3309 (N_3309,N_2263,N_297);
and U3310 (N_3310,N_1147,N_2842);
and U3311 (N_3311,N_2110,N_2651);
or U3312 (N_3312,N_778,N_2681);
and U3313 (N_3313,N_2934,N_1450);
nand U3314 (N_3314,N_1579,N_381);
and U3315 (N_3315,N_1690,N_1742);
and U3316 (N_3316,N_1670,N_1480);
nor U3317 (N_3317,N_2575,N_581);
or U3318 (N_3318,N_2832,N_484);
nor U3319 (N_3319,N_2436,N_75);
and U3320 (N_3320,N_299,N_1766);
and U3321 (N_3321,N_240,N_2485);
or U3322 (N_3322,N_620,N_1887);
and U3323 (N_3323,N_324,N_1150);
or U3324 (N_3324,N_258,N_1082);
nand U3325 (N_3325,N_1522,N_1778);
nor U3326 (N_3326,N_184,N_730);
nand U3327 (N_3327,N_568,N_2891);
or U3328 (N_3328,N_1627,N_1763);
or U3329 (N_3329,N_59,N_2899);
or U3330 (N_3330,N_1338,N_318);
nand U3331 (N_3331,N_2983,N_2167);
or U3332 (N_3332,N_2580,N_1843);
and U3333 (N_3333,N_1874,N_2383);
nand U3334 (N_3334,N_2370,N_2108);
nor U3335 (N_3335,N_1575,N_2932);
and U3336 (N_3336,N_2425,N_2831);
and U3337 (N_3337,N_1865,N_2773);
nand U3338 (N_3338,N_252,N_1946);
and U3339 (N_3339,N_1982,N_2962);
nor U3340 (N_3340,N_472,N_647);
nand U3341 (N_3341,N_249,N_797);
and U3342 (N_3342,N_2002,N_818);
and U3343 (N_3343,N_2153,N_1749);
or U3344 (N_3344,N_1779,N_225);
and U3345 (N_3345,N_2031,N_2344);
nand U3346 (N_3346,N_1081,N_2526);
and U3347 (N_3347,N_1803,N_342);
xor U3348 (N_3348,N_1827,N_1842);
and U3349 (N_3349,N_2058,N_550);
and U3350 (N_3350,N_2549,N_2950);
and U3351 (N_3351,N_2813,N_1404);
and U3352 (N_3352,N_1635,N_1224);
nand U3353 (N_3353,N_2815,N_145);
or U3354 (N_3354,N_2106,N_13);
nand U3355 (N_3355,N_681,N_6);
and U3356 (N_3356,N_529,N_2469);
nor U3357 (N_3357,N_1529,N_510);
and U3358 (N_3358,N_1619,N_2347);
nand U3359 (N_3359,N_917,N_1049);
nor U3360 (N_3360,N_672,N_851);
or U3361 (N_3361,N_2771,N_1976);
or U3362 (N_3362,N_166,N_286);
or U3363 (N_3363,N_2951,N_2168);
or U3364 (N_3364,N_30,N_812);
or U3365 (N_3365,N_2784,N_2178);
and U3366 (N_3366,N_72,N_2798);
nor U3367 (N_3367,N_1571,N_2884);
and U3368 (N_3368,N_560,N_1995);
nor U3369 (N_3369,N_2808,N_837);
and U3370 (N_3370,N_843,N_2251);
or U3371 (N_3371,N_352,N_2509);
nand U3372 (N_3372,N_2532,N_975);
nor U3373 (N_3373,N_631,N_2174);
and U3374 (N_3374,N_1870,N_2299);
nand U3375 (N_3375,N_403,N_301);
and U3376 (N_3376,N_673,N_1379);
nor U3377 (N_3377,N_1061,N_663);
or U3378 (N_3378,N_2064,N_2041);
or U3379 (N_3379,N_671,N_2628);
or U3380 (N_3380,N_246,N_1148);
or U3381 (N_3381,N_2244,N_2970);
or U3382 (N_3382,N_1288,N_18);
or U3383 (N_3383,N_2164,N_944);
nor U3384 (N_3384,N_994,N_1855);
or U3385 (N_3385,N_963,N_2979);
or U3386 (N_3386,N_2280,N_1606);
and U3387 (N_3387,N_201,N_2489);
nand U3388 (N_3388,N_2973,N_170);
nor U3389 (N_3389,N_1176,N_1911);
nor U3390 (N_3390,N_2964,N_2882);
nor U3391 (N_3391,N_687,N_1712);
or U3392 (N_3392,N_1711,N_715);
nor U3393 (N_3393,N_1922,N_1933);
and U3394 (N_3394,N_2904,N_2082);
nand U3395 (N_3395,N_2685,N_1731);
nand U3396 (N_3396,N_1066,N_1735);
nor U3397 (N_3397,N_2947,N_1405);
and U3398 (N_3398,N_480,N_1528);
or U3399 (N_3399,N_1040,N_2496);
and U3400 (N_3400,N_713,N_2643);
or U3401 (N_3401,N_1665,N_1280);
or U3402 (N_3402,N_1846,N_346);
nand U3403 (N_3403,N_102,N_682);
or U3404 (N_3404,N_1923,N_794);
nand U3405 (N_3405,N_844,N_2806);
nand U3406 (N_3406,N_1726,N_443);
nand U3407 (N_3407,N_1106,N_1943);
and U3408 (N_3408,N_1010,N_2817);
nor U3409 (N_3409,N_2713,N_1128);
or U3410 (N_3410,N_1403,N_1467);
nand U3411 (N_3411,N_2273,N_1789);
nor U3412 (N_3412,N_611,N_2417);
or U3413 (N_3413,N_2900,N_2505);
nor U3414 (N_3414,N_1820,N_439);
and U3415 (N_3415,N_1326,N_1017);
and U3416 (N_3416,N_1860,N_929);
nor U3417 (N_3417,N_2249,N_805);
nor U3418 (N_3418,N_904,N_1744);
and U3419 (N_3419,N_1298,N_2598);
nand U3420 (N_3420,N_1745,N_1181);
and U3421 (N_3421,N_655,N_2835);
nor U3422 (N_3422,N_2616,N_290);
nand U3423 (N_3423,N_2342,N_2766);
and U3424 (N_3424,N_941,N_1184);
nand U3425 (N_3425,N_1984,N_763);
and U3426 (N_3426,N_463,N_393);
nand U3427 (N_3427,N_2875,N_1746);
nand U3428 (N_3428,N_1353,N_295);
nor U3429 (N_3429,N_1574,N_2405);
nor U3430 (N_3430,N_486,N_8);
nand U3431 (N_3431,N_1765,N_1089);
or U3432 (N_3432,N_92,N_1013);
or U3433 (N_3433,N_628,N_1699);
nand U3434 (N_3434,N_168,N_1945);
or U3435 (N_3435,N_1252,N_2354);
nand U3436 (N_3436,N_727,N_2399);
or U3437 (N_3437,N_2897,N_1503);
nand U3438 (N_3438,N_2449,N_1701);
or U3439 (N_3439,N_667,N_288);
and U3440 (N_3440,N_1952,N_2446);
and U3441 (N_3441,N_1263,N_641);
and U3442 (N_3442,N_819,N_579);
nor U3443 (N_3443,N_2234,N_475);
nand U3444 (N_3444,N_1424,N_1798);
or U3445 (N_3445,N_1773,N_306);
and U3446 (N_3446,N_2574,N_1463);
or U3447 (N_3447,N_1370,N_901);
and U3448 (N_3448,N_2018,N_36);
or U3449 (N_3449,N_2547,N_1597);
and U3450 (N_3450,N_2317,N_1624);
or U3451 (N_3451,N_601,N_260);
nand U3452 (N_3452,N_1876,N_771);
nor U3453 (N_3453,N_2570,N_2915);
or U3454 (N_3454,N_2232,N_1058);
nor U3455 (N_3455,N_2994,N_608);
and U3456 (N_3456,N_813,N_1357);
nor U3457 (N_3457,N_316,N_2998);
nor U3458 (N_3458,N_2197,N_2261);
or U3459 (N_3459,N_2782,N_1979);
nand U3460 (N_3460,N_968,N_1496);
and U3461 (N_3461,N_1955,N_1637);
and U3462 (N_3462,N_312,N_1580);
nand U3463 (N_3463,N_2931,N_197);
nand U3464 (N_3464,N_1657,N_2662);
nand U3465 (N_3465,N_1055,N_1654);
nor U3466 (N_3466,N_2535,N_2700);
or U3467 (N_3467,N_1769,N_1807);
nand U3468 (N_3468,N_1362,N_541);
or U3469 (N_3469,N_1183,N_2241);
and U3470 (N_3470,N_896,N_1260);
nand U3471 (N_3471,N_512,N_2789);
and U3472 (N_3472,N_2341,N_537);
nor U3473 (N_3473,N_2892,N_2418);
nor U3474 (N_3474,N_1967,N_2752);
or U3475 (N_3475,N_1696,N_1774);
nand U3476 (N_3476,N_1561,N_363);
or U3477 (N_3477,N_115,N_2258);
and U3478 (N_3478,N_250,N_1889);
or U3479 (N_3479,N_1792,N_243);
and U3480 (N_3480,N_1479,N_572);
or U3481 (N_3481,N_427,N_2637);
and U3482 (N_3482,N_2268,N_593);
or U3483 (N_3483,N_1710,N_158);
xnor U3484 (N_3484,N_884,N_190);
and U3485 (N_3485,N_2708,N_965);
or U3486 (N_3486,N_728,N_1990);
and U3487 (N_3487,N_470,N_1991);
nor U3488 (N_3488,N_2786,N_2190);
nand U3489 (N_3489,N_985,N_2923);
and U3490 (N_3490,N_770,N_164);
and U3491 (N_3491,N_2763,N_2149);
nor U3492 (N_3492,N_863,N_1959);
nor U3493 (N_3493,N_40,N_1004);
nor U3494 (N_3494,N_1195,N_2428);
or U3495 (N_3495,N_1777,N_1740);
or U3496 (N_3496,N_1008,N_19);
and U3497 (N_3497,N_284,N_2353);
or U3498 (N_3498,N_167,N_2452);
nand U3499 (N_3499,N_1340,N_399);
and U3500 (N_3500,N_2847,N_2569);
nand U3501 (N_3501,N_1408,N_2940);
or U3502 (N_3502,N_726,N_842);
nor U3503 (N_3503,N_2292,N_2114);
nand U3504 (N_3504,N_1077,N_2756);
nor U3505 (N_3505,N_610,N_2416);
nand U3506 (N_3506,N_810,N_2968);
and U3507 (N_3507,N_211,N_2571);
nand U3508 (N_3508,N_1279,N_1736);
and U3509 (N_3509,N_2793,N_850);
nand U3510 (N_3510,N_1918,N_2595);
and U3511 (N_3511,N_523,N_798);
or U3512 (N_3512,N_2739,N_2288);
nor U3513 (N_3513,N_126,N_195);
nor U3514 (N_3514,N_1213,N_1806);
or U3515 (N_3515,N_1076,N_2734);
and U3516 (N_3516,N_497,N_1104);
and U3517 (N_3517,N_1729,N_2138);
or U3518 (N_3518,N_2386,N_50);
nand U3519 (N_3519,N_1973,N_2780);
nand U3520 (N_3520,N_1240,N_1271);
or U3521 (N_3521,N_2723,N_1235);
and U3522 (N_3522,N_1085,N_1633);
or U3523 (N_3523,N_1487,N_1038);
and U3524 (N_3524,N_2333,N_1756);
nand U3525 (N_3525,N_2530,N_2372);
nor U3526 (N_3526,N_2684,N_429);
nor U3527 (N_3527,N_690,N_2602);
nand U3528 (N_3528,N_2443,N_1762);
nor U3529 (N_3529,N_1559,N_1336);
xnor U3530 (N_3530,N_1120,N_2008);
or U3531 (N_3531,N_2275,N_1239);
nand U3532 (N_3532,N_217,N_978);
nor U3533 (N_3533,N_1725,N_1953);
and U3534 (N_3534,N_2688,N_2431);
nand U3535 (N_3535,N_389,N_1541);
nand U3536 (N_3536,N_57,N_2052);
nand U3537 (N_3537,N_292,N_2310);
nor U3538 (N_3538,N_614,N_2686);
or U3539 (N_3539,N_1395,N_1785);
or U3540 (N_3540,N_1903,N_2539);
nor U3541 (N_3541,N_2568,N_2024);
or U3542 (N_3542,N_1033,N_2357);
xnor U3543 (N_3543,N_1110,N_2161);
nor U3544 (N_3544,N_2924,N_1368);
nand U3545 (N_3545,N_795,N_592);
nor U3546 (N_3546,N_1683,N_1109);
and U3547 (N_3547,N_2117,N_1569);
nand U3548 (N_3548,N_327,N_274);
nor U3549 (N_3549,N_1691,N_2374);
nand U3550 (N_3550,N_2906,N_525);
and U3551 (N_3551,N_1193,N_2862);
and U3552 (N_3552,N_1170,N_1519);
and U3553 (N_3553,N_720,N_2617);
nand U3554 (N_3554,N_2226,N_1916);
nand U3555 (N_3555,N_1754,N_2349);
nand U3556 (N_3556,N_2282,N_2035);
and U3557 (N_3557,N_3,N_417);
xor U3558 (N_3558,N_2820,N_2702);
or U3559 (N_3559,N_1229,N_1123);
xor U3560 (N_3560,N_609,N_2984);
or U3561 (N_3561,N_1475,N_1371);
and U3562 (N_3562,N_1673,N_1748);
or U3563 (N_3563,N_1646,N_1186);
and U3564 (N_3564,N_2460,N_1937);
and U3565 (N_3565,N_1972,N_89);
xor U3566 (N_3566,N_1380,N_749);
xor U3567 (N_3567,N_2495,N_1334);
nand U3568 (N_3568,N_822,N_821);
nor U3569 (N_3569,N_251,N_1443);
and U3570 (N_3570,N_656,N_1360);
and U3571 (N_3571,N_2675,N_1476);
nand U3572 (N_3572,N_2479,N_2854);
xnor U3573 (N_3573,N_1840,N_2230);
nor U3574 (N_3574,N_16,N_873);
or U3575 (N_3575,N_1854,N_1400);
or U3576 (N_3576,N_2855,N_594);
or U3577 (N_3577,N_2735,N_409);
and U3578 (N_3578,N_1311,N_1714);
and U3579 (N_3579,N_244,N_1871);
and U3580 (N_3580,N_1543,N_376);
or U3581 (N_3581,N_1056,N_1163);
and U3582 (N_3582,N_1074,N_1100);
nor U3583 (N_3583,N_2669,N_906);
nand U3584 (N_3584,N_1547,N_1275);
nand U3585 (N_3585,N_293,N_2652);
or U3586 (N_3586,N_877,N_2121);
nor U3587 (N_3587,N_718,N_602);
or U3588 (N_3588,N_2781,N_2100);
and U3589 (N_3589,N_2677,N_992);
xor U3590 (N_3590,N_2466,N_1996);
nor U3591 (N_3591,N_1648,N_2426);
nor U3592 (N_3592,N_1327,N_351);
nand U3593 (N_3593,N_307,N_382);
nor U3594 (N_3594,N_1494,N_2659);
and U3595 (N_3595,N_1330,N_650);
nand U3596 (N_3596,N_1894,N_1582);
and U3597 (N_3597,N_242,N_1006);
and U3598 (N_3598,N_2646,N_2156);
and U3599 (N_3599,N_890,N_2422);
nor U3600 (N_3600,N_1612,N_2521);
xnor U3601 (N_3601,N_1793,N_1679);
and U3602 (N_3602,N_1819,N_2472);
and U3603 (N_3603,N_2032,N_338);
nand U3604 (N_3604,N_1908,N_2716);
or U3605 (N_3605,N_2922,N_1498);
or U3606 (N_3606,N_1425,N_1046);
or U3607 (N_3607,N_402,N_1242);
xor U3608 (N_3608,N_876,N_833);
xnor U3609 (N_3609,N_2348,N_2912);
nand U3610 (N_3610,N_127,N_664);
or U3611 (N_3611,N_2937,N_361);
nor U3612 (N_3612,N_445,N_1988);
or U3613 (N_3613,N_1675,N_2941);
and U3614 (N_3614,N_2049,N_1426);
nand U3615 (N_3615,N_422,N_2682);
or U3616 (N_3616,N_2112,N_1435);
nor U3617 (N_3617,N_323,N_1770);
and U3618 (N_3618,N_539,N_1951);
and U3619 (N_3619,N_1751,N_273);
nor U3620 (N_3620,N_2073,N_173);
xnor U3621 (N_3621,N_814,N_336);
and U3622 (N_3622,N_935,N_1965);
nor U3623 (N_3623,N_888,N_2009);
nand U3624 (N_3624,N_1258,N_2630);
nor U3625 (N_3625,N_123,N_1328);
or U3626 (N_3626,N_2136,N_345);
or U3627 (N_3627,N_2645,N_2852);
nor U3628 (N_3628,N_2375,N_111);
nor U3629 (N_3629,N_407,N_2010);
or U3630 (N_3630,N_1513,N_1348);
and U3631 (N_3631,N_2166,N_2581);
nor U3632 (N_3632,N_1135,N_373);
and U3633 (N_3633,N_2423,N_2749);
nand U3634 (N_3634,N_82,N_2477);
and U3635 (N_3635,N_2211,N_261);
or U3636 (N_3636,N_1026,N_2276);
nor U3637 (N_3637,N_533,N_186);
and U3638 (N_3638,N_2451,N_2109);
or U3639 (N_3639,N_1188,N_1364);
or U3640 (N_3640,N_1367,N_1909);
nand U3641 (N_3641,N_1542,N_1788);
or U3642 (N_3642,N_1143,N_1416);
nor U3643 (N_3643,N_1518,N_202);
and U3644 (N_3644,N_1966,N_1692);
and U3645 (N_3645,N_64,N_181);
or U3646 (N_3646,N_1369,N_1462);
nand U3647 (N_3647,N_2559,N_933);
or U3648 (N_3648,N_708,N_499);
nand U3649 (N_3649,N_2332,N_2044);
or U3650 (N_3650,N_1629,N_2603);
nor U3651 (N_3651,N_172,N_2067);
nand U3652 (N_3652,N_1388,N_2247);
nand U3653 (N_3653,N_255,N_612);
and U3654 (N_3654,N_1019,N_129);
xor U3655 (N_3655,N_1873,N_1781);
or U3656 (N_3656,N_2562,N_146);
or U3657 (N_3657,N_2088,N_1509);
nand U3658 (N_3658,N_791,N_2104);
nand U3659 (N_3659,N_175,N_2462);
or U3660 (N_3660,N_1247,N_695);
nor U3661 (N_3661,N_1343,N_2407);
nand U3662 (N_3662,N_2837,N_1111);
nand U3663 (N_3663,N_514,N_2366);
or U3664 (N_3664,N_1358,N_406);
nand U3665 (N_3665,N_1882,N_1783);
nand U3666 (N_3666,N_1437,N_1419);
or U3667 (N_3667,N_315,N_2283);
or U3668 (N_3668,N_2113,N_66);
nand U3669 (N_3669,N_1895,N_2668);
nand U3670 (N_3670,N_1915,N_548);
nand U3671 (N_3671,N_1474,N_1088);
nor U3672 (N_3672,N_107,N_341);
nand U3673 (N_3673,N_866,N_707);
and U3674 (N_3674,N_434,N_1759);
nor U3675 (N_3675,N_256,N_1321);
and U3676 (N_3676,N_462,N_1968);
nor U3677 (N_3677,N_2319,N_1577);
nor U3678 (N_3678,N_264,N_253);
or U3679 (N_3679,N_1162,N_2838);
or U3680 (N_3680,N_2927,N_2455);
nor U3681 (N_3681,N_1309,N_254);
or U3682 (N_3682,N_2720,N_932);
nor U3683 (N_3683,N_212,N_789);
and U3684 (N_3684,N_2626,N_2958);
or U3685 (N_3685,N_619,N_1043);
or U3686 (N_3686,N_2989,N_2849);
nand U3687 (N_3687,N_2102,N_2382);
or U3688 (N_3688,N_1335,N_776);
and U3689 (N_3689,N_2680,N_1505);
nand U3690 (N_3690,N_685,N_200);
or U3691 (N_3691,N_2910,N_2704);
and U3692 (N_3692,N_691,N_2952);
nand U3693 (N_3693,N_2977,N_269);
or U3694 (N_3694,N_784,N_2465);
and U3695 (N_3695,N_2810,N_35);
and U3696 (N_3696,N_2516,N_2640);
nor U3697 (N_3697,N_159,N_1265);
and U3698 (N_3698,N_456,N_945);
nor U3699 (N_3699,N_275,N_2406);
nand U3700 (N_3700,N_981,N_1118);
or U3701 (N_3701,N_2224,N_621);
nor U3702 (N_3702,N_1428,N_1674);
or U3703 (N_3703,N_1130,N_2379);
or U3704 (N_3704,N_1478,N_1484);
nor U3705 (N_3705,N_2339,N_2209);
and U3706 (N_3706,N_2577,N_232);
and U3707 (N_3707,N_2819,N_7);
and U3708 (N_3708,N_1962,N_228);
nand U3709 (N_3709,N_1094,N_792);
nand U3710 (N_3710,N_171,N_377);
nor U3711 (N_3711,N_1441,N_1436);
nand U3712 (N_3712,N_2566,N_2938);
or U3713 (N_3713,N_2097,N_1129);
nand U3714 (N_3714,N_1194,N_657);
xor U3715 (N_3715,N_199,N_897);
and U3716 (N_3716,N_1588,N_1639);
nand U3717 (N_3717,N_2841,N_538);
or U3718 (N_3718,N_921,N_989);
and U3719 (N_3719,N_1755,N_2541);
nor U3720 (N_3720,N_2200,N_1938);
and U3721 (N_3721,N_1684,N_1552);
and U3722 (N_3722,N_1570,N_2778);
and U3723 (N_3723,N_133,N_781);
and U3724 (N_3724,N_777,N_1037);
nor U3725 (N_3725,N_2809,N_1797);
or U3726 (N_3726,N_2410,N_2185);
nand U3727 (N_3727,N_1446,N_2527);
or U3728 (N_3728,N_2392,N_1761);
or U3729 (N_3729,N_1644,N_279);
or U3730 (N_3730,N_2165,N_1934);
nand U3731 (N_3731,N_1615,N_337);
nor U3732 (N_3732,N_1722,N_1359);
or U3733 (N_3733,N_1313,N_1080);
or U3734 (N_3734,N_1132,N_1834);
xor U3735 (N_3735,N_860,N_2754);
nand U3736 (N_3736,N_2657,N_1677);
or U3737 (N_3737,N_2554,N_1913);
or U3738 (N_3738,N_536,N_490);
xor U3739 (N_3739,N_871,N_2667);
or U3740 (N_3740,N_1706,N_267);
nand U3741 (N_3741,N_1585,N_1001);
or U3742 (N_3742,N_2139,N_577);
and U3743 (N_3743,N_2326,N_154);
nand U3744 (N_3744,N_174,N_1906);
nand U3745 (N_3745,N_2865,N_374);
and U3746 (N_3746,N_2303,N_1511);
nor U3747 (N_3747,N_1073,N_1687);
nand U3748 (N_3748,N_2151,N_2942);
and U3749 (N_3749,N_1168,N_865);
nor U3750 (N_3750,N_626,N_2442);
nor U3751 (N_3751,N_2127,N_1202);
and U3752 (N_3752,N_870,N_1723);
and U3753 (N_3753,N_1047,N_889);
nor U3754 (N_3754,N_1501,N_1532);
nand U3755 (N_3755,N_1825,N_2772);
and U3756 (N_3756,N_954,N_5);
nor U3757 (N_3757,N_934,N_68);
xnor U3758 (N_3758,N_2578,N_2930);
nor U3759 (N_3759,N_2706,N_2300);
nor U3760 (N_3760,N_540,N_270);
or U3761 (N_3761,N_1879,N_951);
nand U3762 (N_3762,N_1375,N_2237);
and U3763 (N_3763,N_1268,N_1897);
or U3764 (N_3764,N_79,N_654);
or U3765 (N_3765,N_883,N_2850);
nor U3766 (N_3766,N_436,N_1549);
nor U3767 (N_3767,N_2202,N_2327);
nand U3768 (N_3768,N_2858,N_847);
and U3769 (N_3769,N_2248,N_1892);
or U3770 (N_3770,N_2691,N_982);
and U3771 (N_3771,N_2269,N_570);
and U3772 (N_3772,N_1097,N_1811);
nor U3773 (N_3773,N_426,N_2133);
nor U3774 (N_3774,N_1121,N_1304);
or U3775 (N_3775,N_1051,N_2779);
and U3776 (N_3776,N_878,N_239);
nor U3777 (N_3777,N_2565,N_191);
and U3778 (N_3778,N_411,N_23);
nand U3779 (N_3779,N_391,N_1251);
nand U3780 (N_3780,N_1302,N_180);
or U3781 (N_3781,N_287,N_2822);
or U3782 (N_3782,N_464,N_105);
nand U3783 (N_3783,N_22,N_2198);
nor U3784 (N_3784,N_1601,N_1175);
nand U3785 (N_3785,N_584,N_1611);
nor U3786 (N_3786,N_2879,N_2358);
or U3787 (N_3787,N_2679,N_2714);
nor U3788 (N_3788,N_2011,N_908);
and U3789 (N_3789,N_712,N_576);
nor U3790 (N_3790,N_368,N_2801);
and U3791 (N_3791,N_1554,N_2800);
and U3792 (N_3792,N_1643,N_604);
nand U3793 (N_3793,N_1926,N_2059);
nand U3794 (N_3794,N_205,N_1593);
xnor U3795 (N_3795,N_638,N_706);
nand U3796 (N_3796,N_1126,N_1325);
nand U3797 (N_3797,N_2141,N_1893);
nor U3798 (N_3798,N_2421,N_1299);
nor U3799 (N_3799,N_1660,N_1459);
nor U3800 (N_3800,N_419,N_1189);
nand U3801 (N_3801,N_2502,N_2316);
nor U3802 (N_3802,N_535,N_1254);
and U3803 (N_3803,N_2834,N_1156);
xnor U3804 (N_3804,N_1386,N_157);
nor U3805 (N_3805,N_2350,N_1929);
and U3806 (N_3806,N_575,N_372);
or U3807 (N_3807,N_2593,N_1910);
or U3808 (N_3808,N_2294,N_55);
or U3809 (N_3809,N_1414,N_1521);
or U3810 (N_3810,N_1636,N_2208);
and U3811 (N_3811,N_767,N_2000);
or U3812 (N_3812,N_178,N_2843);
nand U3813 (N_3813,N_1919,N_2171);
nand U3814 (N_3814,N_2093,N_2187);
nand U3815 (N_3815,N_153,N_2308);
and U3816 (N_3816,N_689,N_1664);
nand U3817 (N_3817,N_1384,N_2131);
nand U3818 (N_3818,N_2957,N_2799);
and U3819 (N_3819,N_1339,N_1721);
nand U3820 (N_3820,N_1998,N_1218);
nand U3821 (N_3821,N_723,N_1087);
or U3822 (N_3822,N_2217,N_2250);
or U3823 (N_3823,N_455,N_1986);
and U3824 (N_3824,N_359,N_1329);
nand U3825 (N_3825,N_2397,N_424);
and U3826 (N_3826,N_1472,N_2218);
nor U3827 (N_3827,N_552,N_447);
and U3828 (N_3828,N_2045,N_2322);
and U3829 (N_3829,N_1342,N_1767);
and U3830 (N_3830,N_2795,N_231);
nor U3831 (N_3831,N_993,N_639);
or U3832 (N_3832,N_117,N_2678);
and U3833 (N_3833,N_1412,N_753);
nor U3834 (N_3834,N_1211,N_2607);
nor U3835 (N_3835,N_943,N_493);
or U3836 (N_3836,N_542,N_15);
and U3837 (N_3837,N_914,N_2336);
nand U3838 (N_3838,N_2889,N_972);
and U3839 (N_3839,N_633,N_1500);
and U3840 (N_3840,N_2825,N_1583);
or U3841 (N_3841,N_1197,N_2245);
nor U3842 (N_3842,N_42,N_793);
and U3843 (N_3843,N_2916,N_2967);
nor U3844 (N_3844,N_1954,N_1925);
nand U3845 (N_3845,N_1290,N_2615);
and U3846 (N_3846,N_2563,N_385);
and U3847 (N_3847,N_1506,N_1750);
nand U3848 (N_3848,N_2634,N_2229);
or U3849 (N_3849,N_2954,N_807);
nor U3850 (N_3850,N_94,N_2012);
nand U3851 (N_3851,N_1264,N_1060);
nor U3852 (N_3852,N_1659,N_2037);
and U3853 (N_3853,N_2204,N_1139);
and U3854 (N_3854,N_33,N_360);
and U3855 (N_3855,N_32,N_1069);
nand U3856 (N_3856,N_51,N_230);
nor U3857 (N_3857,N_2207,N_87);
nand U3858 (N_3858,N_2070,N_1103);
nor U3859 (N_3859,N_1666,N_1656);
nor U3860 (N_3860,N_2027,N_1050);
nand U3861 (N_3861,N_902,N_1847);
nand U3862 (N_3862,N_319,N_1083);
nor U3863 (N_3863,N_1378,N_2863);
or U3864 (N_3864,N_892,N_802);
nand U3865 (N_3865,N_2903,N_1071);
or U3866 (N_3866,N_2116,N_1632);
nand U3867 (N_3867,N_2180,N_2124);
and U3868 (N_3868,N_1537,N_2296);
nor U3869 (N_3869,N_2913,N_144);
and U3870 (N_3870,N_780,N_1645);
or U3871 (N_3871,N_1553,N_1141);
nor U3872 (N_3872,N_1114,N_1286);
or U3873 (N_3873,N_2528,N_2225);
and U3874 (N_3874,N_2726,N_1550);
xor U3875 (N_3875,N_1291,N_1351);
nand U3876 (N_3876,N_1753,N_233);
nand U3877 (N_3877,N_2006,N_296);
nand U3878 (N_3878,N_328,N_80);
nand U3879 (N_3879,N_1098,N_2633);
nor U3880 (N_3880,N_1312,N_1297);
nand U3881 (N_3881,N_987,N_1262);
and U3882 (N_3882,N_2311,N_757);
and U3883 (N_3883,N_2140,N_2750);
and U3884 (N_3884,N_1075,N_311);
or U3885 (N_3885,N_2091,N_241);
nor U3886 (N_3886,N_2802,N_948);
nor U3887 (N_3887,N_2255,N_1622);
or U3888 (N_3888,N_754,N_1720);
nand U3889 (N_3889,N_1859,N_2671);
nand U3890 (N_3890,N_2902,N_759);
nor U3891 (N_3891,N_569,N_320);
xor U3892 (N_3892,N_765,N_2661);
nand U3893 (N_3893,N_2066,N_2748);
xor U3894 (N_3894,N_731,N_2056);
nor U3895 (N_3895,N_1799,N_2068);
nor U3896 (N_3896,N_152,N_1471);
nand U3897 (N_3897,N_76,N_606);
nand U3898 (N_3898,N_769,N_140);
nand U3899 (N_3899,N_58,N_2534);
or U3900 (N_3900,N_2476,N_1676);
nand U3901 (N_3901,N_2728,N_1738);
or U3902 (N_3902,N_2995,N_2313);
nand U3903 (N_3903,N_1578,N_1032);
and U3904 (N_3904,N_825,N_1768);
nor U3905 (N_3905,N_2960,N_2427);
and U3906 (N_3906,N_2826,N_808);
or U3907 (N_3907,N_2538,N_86);
nand U3908 (N_3908,N_2579,N_2629);
nand U3909 (N_3909,N_2555,N_1948);
nand U3910 (N_3910,N_1828,N_2101);
or U3911 (N_3911,N_2846,N_2334);
nand U3912 (N_3912,N_2518,N_554);
nand U3913 (N_3913,N_839,N_2925);
or U3914 (N_3914,N_1546,N_1140);
nand U3915 (N_3915,N_12,N_1306);
and U3916 (N_3916,N_2270,N_1117);
nand U3917 (N_3917,N_44,N_998);
or U3918 (N_3918,N_1065,N_590);
or U3919 (N_3919,N_629,N_1497);
nor U3920 (N_3920,N_1178,N_1406);
nor U3921 (N_3921,N_2152,N_163);
or U3922 (N_3922,N_688,N_104);
nor U3923 (N_3923,N_862,N_2220);
and U3924 (N_3924,N_444,N_1861);
nor U3925 (N_3925,N_1872,N_561);
xor U3926 (N_3926,N_1747,N_1289);
nand U3927 (N_3927,N_423,N_1890);
nor U3928 (N_3928,N_2732,N_2040);
or U3929 (N_3929,N_2159,N_1507);
nand U3930 (N_3930,N_2918,N_857);
or U3931 (N_3931,N_2632,N_867);
nor U3932 (N_3932,N_905,N_454);
or U3933 (N_3933,N_2558,N_2880);
nor U3934 (N_3934,N_113,N_1698);
or U3935 (N_3935,N_1829,N_1257);
and U3936 (N_3936,N_2071,N_2878);
or U3937 (N_3937,N_2725,N_803);
nand U3938 (N_3938,N_1896,N_1272);
and U3939 (N_3939,N_2999,N_1249);
or U3940 (N_3940,N_613,N_2278);
or U3941 (N_3941,N_2519,N_964);
and U3942 (N_3942,N_2948,N_142);
nand U3943 (N_3943,N_2448,N_1011);
or U3944 (N_3944,N_2315,N_2438);
or U3945 (N_3945,N_1595,N_139);
and U3946 (N_3946,N_679,N_2033);
and U3947 (N_3947,N_2503,N_1427);
nor U3948 (N_3948,N_97,N_1605);
nor U3949 (N_3949,N_1020,N_2919);
and U3950 (N_3950,N_2965,N_1974);
nor U3951 (N_3951,N_1833,N_1457);
nor U3952 (N_3952,N_696,N_101);
nor U3953 (N_3953,N_2490,N_2364);
nor U3954 (N_3954,N_213,N_227);
or U3955 (N_3955,N_280,N_467);
and U3956 (N_3956,N_2147,N_2458);
nand U3957 (N_3957,N_1686,N_2807);
nand U3958 (N_3958,N_458,N_2361);
and U3959 (N_3959,N_1775,N_0);
nand U3960 (N_3960,N_2301,N_28);
or U3961 (N_3961,N_2840,N_1839);
and U3962 (N_3962,N_271,N_2876);
or U3963 (N_3963,N_1090,N_461);
nand U3964 (N_3964,N_2393,N_1383);
nor U3965 (N_3965,N_1700,N_2395);
and U3966 (N_3966,N_405,N_1390);
nor U3967 (N_3967,N_1323,N_732);
xnor U3968 (N_3968,N_565,N_2063);
or U3969 (N_3969,N_2289,N_2928);
nand U3970 (N_3970,N_2478,N_2387);
or U3971 (N_3971,N_2279,N_2360);
or U3972 (N_3972,N_2169,N_1301);
nor U3973 (N_3973,N_2345,N_1219);
nand U3974 (N_3974,N_2172,N_2510);
and U3975 (N_3975,N_919,N_2243);
xor U3976 (N_3976,N_1531,N_1805);
nor U3977 (N_3977,N_1245,N_595);
nand U3978 (N_3978,N_2644,N_738);
nand U3979 (N_3979,N_300,N_2639);
or U3980 (N_3980,N_132,N_1160);
and U3981 (N_3981,N_27,N_1300);
and U3982 (N_3982,N_330,N_2710);
or U3983 (N_3983,N_1296,N_2981);
or U3984 (N_3984,N_1387,N_2467);
and U3985 (N_3985,N_755,N_1914);
nor U3986 (N_3986,N_1112,N_1856);
or U3987 (N_3987,N_21,N_1223);
xnor U3988 (N_3988,N_2935,N_1493);
nor U3989 (N_3989,N_1607,N_1381);
or U3990 (N_3990,N_2511,N_1837);
or U3991 (N_3991,N_2868,N_1003);
nand U3992 (N_3992,N_2567,N_1836);
nand U3993 (N_3993,N_834,N_2604);
nand U3994 (N_3994,N_1014,N_665);
nand U3995 (N_3995,N_1898,N_2470);
or U3996 (N_3996,N_2355,N_1401);
and U3997 (N_3997,N_957,N_1155);
nor U3998 (N_3998,N_108,N_1693);
or U3999 (N_3999,N_2666,N_2481);
and U4000 (N_4000,N_215,N_2483);
and U4001 (N_4001,N_796,N_1084);
nand U4002 (N_4002,N_946,N_2210);
and U4003 (N_4003,N_1917,N_1167);
or U4004 (N_4004,N_65,N_2367);
nand U4005 (N_4005,N_2281,N_2761);
or U4006 (N_4006,N_522,N_591);
and U4007 (N_4007,N_1250,N_2021);
or U4008 (N_4008,N_2551,N_2917);
and U4009 (N_4009,N_149,N_440);
nand U4010 (N_4010,N_1394,N_1208);
and U4011 (N_4011,N_2926,N_1295);
nand U4012 (N_4012,N_2546,N_1492);
nand U4013 (N_4013,N_2830,N_2075);
nor U4014 (N_4014,N_1154,N_2621);
or U4015 (N_4015,N_2966,N_886);
or U4016 (N_4016,N_266,N_1620);
nand U4017 (N_4017,N_1641,N_466);
nand U4018 (N_4018,N_2272,N_1510);
nor U4019 (N_4019,N_518,N_2233);
or U4020 (N_4020,N_1366,N_1517);
or U4021 (N_4021,N_134,N_1456);
and U4022 (N_4022,N_1950,N_2203);
xor U4023 (N_4023,N_950,N_1231);
nor U4024 (N_4024,N_2256,N_1709);
nand U4025 (N_4025,N_2036,N_294);
nand U4026 (N_4026,N_1063,N_489);
or U4027 (N_4027,N_838,N_366);
nand U4028 (N_4028,N_2072,N_2522);
xor U4029 (N_4029,N_1526,N_1029);
nand U4030 (N_4030,N_578,N_2415);
nor U4031 (N_4031,N_1533,N_1812);
and U4032 (N_4032,N_1173,N_1086);
and U4033 (N_4033,N_2997,N_1282);
and U4034 (N_4034,N_2094,N_2005);
nand U4035 (N_4035,N_481,N_2985);
or U4036 (N_4036,N_740,N_721);
nor U4037 (N_4037,N_2409,N_2945);
nor U4038 (N_4038,N_1373,N_2636);
nand U4039 (N_4039,N_1791,N_939);
or U4040 (N_4040,N_2743,N_2552);
nor U4041 (N_4041,N_1031,N_683);
or U4042 (N_4042,N_20,N_1350);
and U4043 (N_4043,N_2475,N_2507);
and U4044 (N_4044,N_1490,N_1255);
nor U4045 (N_4045,N_143,N_1174);
and U4046 (N_4046,N_88,N_2158);
or U4047 (N_4047,N_1796,N_1179);
nor U4048 (N_4048,N_276,N_321);
and U4049 (N_4049,N_2573,N_1667);
nand U4050 (N_4050,N_1730,N_1485);
or U4051 (N_4051,N_2074,N_1444);
and U4052 (N_4052,N_2461,N_2872);
or U4053 (N_4053,N_2134,N_545);
and U4054 (N_4054,N_2219,N_701);
or U4055 (N_4055,N_907,N_868);
nand U4056 (N_4056,N_120,N_473);
nand U4057 (N_4057,N_2513,N_2883);
or U4058 (N_4058,N_1592,N_1545);
nor U4059 (N_4059,N_702,N_1200);
nand U4060 (N_4060,N_2553,N_2343);
or U4061 (N_4061,N_2492,N_2797);
nand U4062 (N_4062,N_1005,N_203);
xor U4063 (N_4063,N_2020,N_2974);
nor U4064 (N_4064,N_304,N_1228);
nor U4065 (N_4065,N_1220,N_193);
and U4066 (N_4066,N_2083,N_2007);
nor U4067 (N_4067,N_729,N_2887);
or U4068 (N_4068,N_2894,N_2992);
nand U4069 (N_4069,N_2111,N_1867);
and U4070 (N_4070,N_617,N_1963);
and U4071 (N_4071,N_1800,N_2697);
nor U4072 (N_4072,N_1153,N_1191);
nand U4073 (N_4073,N_1382,N_2085);
or U4074 (N_4074,N_936,N_1248);
or U4075 (N_4075,N_1555,N_2148);
nand U4076 (N_4076,N_2625,N_1102);
and U4077 (N_4077,N_918,N_2776);
nand U4078 (N_4078,N_2886,N_448);
nor U4079 (N_4079,N_247,N_1023);
or U4080 (N_4080,N_1207,N_268);
nand U4081 (N_4081,N_2533,N_1784);
or U4082 (N_4082,N_758,N_2356);
and U4083 (N_4083,N_1681,N_2610);
nor U4084 (N_4084,N_2145,N_2515);
or U4085 (N_4085,N_2796,N_1346);
and U4086 (N_4086,N_367,N_2352);
or U4087 (N_4087,N_1447,N_2689);
nor U4088 (N_4088,N_501,N_2529);
or U4089 (N_4089,N_2642,N_2753);
nor U4090 (N_4090,N_1530,N_2594);
and U4091 (N_4091,N_2262,N_446);
and U4092 (N_4092,N_329,N_1453);
and U4093 (N_4093,N_885,N_2137);
or U4094 (N_4094,N_2051,N_1904);
nor U4095 (N_4095,N_1743,N_1238);
nor U4096 (N_4096,N_1320,N_303);
or U4097 (N_4097,N_124,N_355);
xnor U4098 (N_4098,N_1489,N_1883);
nor U4099 (N_4099,N_1276,N_546);
nor U4100 (N_4100,N_2833,N_1418);
nand U4101 (N_4101,N_438,N_2260);
nor U4102 (N_4102,N_1841,N_598);
nor U4103 (N_4103,N_1628,N_1363);
and U4104 (N_4104,N_1172,N_1572);
nand U4105 (N_4105,N_1021,N_2221);
nor U4106 (N_4106,N_2337,N_278);
nand U4107 (N_4107,N_1576,N_658);
or U4108 (N_4108,N_928,N_547);
nor U4109 (N_4109,N_1614,N_1584);
or U4110 (N_4110,N_1878,N_1932);
and U4111 (N_4111,N_1234,N_845);
and U4112 (N_4112,N_916,N_2189);
nand U4113 (N_4113,N_997,N_2257);
and U4114 (N_4114,N_2142,N_2026);
nand U4115 (N_4115,N_1845,N_1201);
or U4116 (N_4116,N_567,N_1757);
nor U4117 (N_4117,N_2419,N_1307);
nand U4118 (N_4118,N_1442,N_2881);
nor U4119 (N_4119,N_95,N_2614);
nand U4120 (N_4120,N_1230,N_2727);
or U4121 (N_4121,N_2184,N_2693);
nand U4122 (N_4122,N_331,N_2971);
nor U4123 (N_4123,N_607,N_1161);
and U4124 (N_4124,N_2641,N_1062);
nor U4125 (N_4125,N_1454,N_990);
and U4126 (N_4126,N_2718,N_2805);
or U4127 (N_4127,N_680,N_2253);
and U4128 (N_4128,N_1376,N_2213);
nand U4129 (N_4129,N_1482,N_700);
or U4130 (N_4130,N_1410,N_1439);
nand U4131 (N_4131,N_527,N_926);
or U4132 (N_4132,N_2430,N_772);
nor U4133 (N_4133,N_2592,N_912);
and U4134 (N_4134,N_1415,N_398);
nor U4135 (N_4135,N_1455,N_2703);
nor U4136 (N_4136,N_724,N_386);
or U4137 (N_4137,N_1420,N_1772);
nor U4138 (N_4138,N_1158,N_603);
and U4139 (N_4139,N_938,N_2986);
and U4140 (N_4140,N_151,N_1816);
or U4141 (N_4141,N_418,N_488);
nand U4142 (N_4142,N_1015,N_2803);
or U4143 (N_4143,N_11,N_262);
nand U4144 (N_4144,N_1508,N_2584);
nand U4145 (N_4145,N_1460,N_2871);
and U4146 (N_4146,N_2025,N_2619);
or U4147 (N_4147,N_60,N_2034);
or U4148 (N_4148,N_735,N_1324);
and U4149 (N_4149,N_78,N_431);
and U4150 (N_4150,N_2572,N_637);
nand U4151 (N_4151,N_1217,N_285);
or U4152 (N_4152,N_2921,N_615);
nor U4153 (N_4153,N_2609,N_347);
nand U4154 (N_4154,N_899,N_2411);
and U4155 (N_4155,N_1012,N_1671);
nor U4156 (N_4156,N_375,N_2638);
or U4157 (N_4157,N_1921,N_1741);
and U4158 (N_4158,N_1630,N_2499);
xor U4159 (N_4159,N_348,N_198);
and U4160 (N_4160,N_2737,N_2155);
nand U4161 (N_4161,N_2823,N_2588);
and U4162 (N_4162,N_1844,N_99);
nor U4163 (N_4163,N_2600,N_1830);
and U4164 (N_4164,N_325,N_2401);
nand U4165 (N_4165,N_2048,N_956);
xnor U4166 (N_4166,N_226,N_1556);
nand U4167 (N_4167,N_2953,N_559);
nor U4168 (N_4168,N_2323,N_441);
or U4169 (N_4169,N_1256,N_2993);
nor U4170 (N_4170,N_2586,N_1101);
nand U4171 (N_4171,N_2654,N_2321);
nand U4172 (N_4172,N_2324,N_1936);
nand U4173 (N_4173,N_2698,N_774);
nand U4174 (N_4174,N_894,N_189);
nor U4175 (N_4175,N_1409,N_1581);
nand U4176 (N_4176,N_586,N_2821);
and U4177 (N_4177,N_1432,N_1146);
or U4178 (N_4178,N_63,N_563);
nand U4179 (N_4179,N_1851,N_2338);
or U4180 (N_4180,N_2596,N_958);
and U4181 (N_4181,N_2517,N_1374);
nor U4182 (N_4182,N_999,N_2266);
nor U4183 (N_4183,N_2090,N_1969);
nor U4184 (N_4184,N_920,N_627);
xnor U4185 (N_4185,N_553,N_1520);
and U4186 (N_4186,N_2192,N_1115);
nand U4187 (N_4187,N_705,N_1196);
or U4188 (N_4188,N_2486,N_1044);
nand U4189 (N_4189,N_333,N_2464);
nor U4190 (N_4190,N_676,N_2454);
and U4191 (N_4191,N_2620,N_2305);
nor U4192 (N_4192,N_234,N_2874);
or U4193 (N_4193,N_1261,N_2441);
nor U4194 (N_4194,N_1647,N_922);
nor U4195 (N_4195,N_642,N_1322);
and U4196 (N_4196,N_2445,N_2015);
and U4197 (N_4197,N_421,N_2929);
or U4198 (N_4198,N_2500,N_130);
nand U4199 (N_4199,N_622,N_1283);
nor U4200 (N_4200,N_587,N_1396);
nand U4201 (N_4201,N_775,N_45);
nand U4202 (N_4202,N_1352,N_2182);
nand U4203 (N_4203,N_135,N_2060);
and U4204 (N_4204,N_508,N_762);
nand U4205 (N_4205,N_2665,N_1016);
nand U4206 (N_4206,N_786,N_2022);
or U4207 (N_4207,N_2601,N_2804);
nor U4208 (N_4208,N_1465,N_1438);
nor U4209 (N_4209,N_1602,N_1817);
or U4210 (N_4210,N_1662,N_2346);
nor U4211 (N_4211,N_308,N_474);
nand U4212 (N_4212,N_2274,N_1957);
nand U4213 (N_4213,N_2267,N_2376);
and U4214 (N_4214,N_2437,N_820);
or U4215 (N_4215,N_221,N_137);
and U4216 (N_4216,N_1902,N_1177);
nand U4217 (N_4217,N_1724,N_566);
nor U4218 (N_4218,N_1199,N_736);
and U4219 (N_4219,N_1009,N_1107);
xor U4220 (N_4220,N_504,N_1149);
nor U4221 (N_4221,N_983,N_61);
or U4222 (N_4222,N_675,N_2047);
nor U4223 (N_4223,N_2975,N_549);
or U4224 (N_4224,N_2046,N_1292);
nand U4225 (N_4225,N_1566,N_2228);
and U4226 (N_4226,N_2866,N_2450);
nor U4227 (N_4227,N_2759,N_2284);
nand U4228 (N_4228,N_2328,N_828);
nand U4229 (N_4229,N_1093,N_893);
nor U4230 (N_4230,N_1695,N_513);
nand U4231 (N_4231,N_2128,N_182);
and U4232 (N_4232,N_2329,N_2920);
and U4233 (N_4233,N_2028,N_103);
or U4234 (N_4234,N_1704,N_2384);
nand U4235 (N_4235,N_1591,N_1663);
or U4236 (N_4236,N_2404,N_915);
and U4237 (N_4237,N_2057,N_2186);
nand U4238 (N_4238,N_1423,N_2542);
nand U4239 (N_4239,N_2163,N_277);
or U4240 (N_4240,N_2767,N_2673);
and U4241 (N_4241,N_2029,N_219);
nor U4242 (N_4242,N_2291,N_2955);
nor U4243 (N_4243,N_1099,N_1920);
nor U4244 (N_4244,N_116,N_37);
or U4245 (N_4245,N_1733,N_2242);
or U4246 (N_4246,N_1702,N_651);
nor U4247 (N_4247,N_1127,N_1661);
or U4248 (N_4248,N_2179,N_425);
nand U4249 (N_4249,N_400,N_2524);
nand U4250 (N_4250,N_121,N_2191);
nor U4251 (N_4251,N_955,N_636);
nand U4252 (N_4252,N_2,N_2188);
or U4253 (N_4253,N_2277,N_2199);
nand U4254 (N_4254,N_1794,N_1824);
or U4255 (N_4255,N_582,N_309);
nor U4256 (N_4256,N_192,N_2381);
and U4257 (N_4257,N_787,N_2054);
or U4258 (N_4258,N_2023,N_507);
or U4259 (N_4259,N_272,N_2122);
or U4260 (N_4260,N_482,N_653);
and U4261 (N_4261,N_220,N_555);
or U4262 (N_4262,N_2484,N_699);
or U4263 (N_4263,N_1232,N_460);
or U4264 (N_4264,N_2764,N_630);
and U4265 (N_4265,N_528,N_1072);
nand U4266 (N_4266,N_1732,N_526);
nand U4267 (N_4267,N_2065,N_737);
nor U4268 (N_4268,N_1233,N_2369);
or U4269 (N_4269,N_521,N_952);
nor U4270 (N_4270,N_836,N_1534);
nand U4271 (N_4271,N_1070,N_532);
nand U4272 (N_4272,N_1402,N_437);
nor U4273 (N_4273,N_2325,N_2751);
nand U4274 (N_4274,N_2663,N_562);
or U4275 (N_4275,N_1924,N_811);
nand U4276 (N_4276,N_1562,N_741);
nor U4277 (N_4277,N_487,N_745);
or U4278 (N_4278,N_785,N_291);
or U4279 (N_4279,N_589,N_2359);
and U4280 (N_4280,N_2946,N_1760);
nand U4281 (N_4281,N_2488,N_2240);
or U4282 (N_4282,N_1971,N_222);
nand U4283 (N_4283,N_1590,N_670);
or U4284 (N_4284,N_283,N_710);
nand U4285 (N_4285,N_2582,N_2331);
nand U4286 (N_4286,N_980,N_1617);
nand U4287 (N_4287,N_1831,N_734);
and U4288 (N_4288,N_1203,N_2078);
nor U4289 (N_4289,N_766,N_2963);
nand U4290 (N_4290,N_1715,N_1801);
nor U4291 (N_4291,N_1987,N_852);
and U4292 (N_4292,N_430,N_2790);
and U4293 (N_4293,N_979,N_2540);
nand U4294 (N_4294,N_1524,N_2811);
nand U4295 (N_4295,N_714,N_909);
nor U4296 (N_4296,N_1068,N_2086);
and U4297 (N_4297,N_1469,N_2320);
or U4298 (N_4298,N_571,N_1159);
xnor U4299 (N_4299,N_678,N_1440);
nor U4300 (N_4300,N_1707,N_2564);
or U4301 (N_4301,N_2235,N_41);
and U4302 (N_4302,N_677,N_2205);
and U4303 (N_4303,N_289,N_1668);
nor U4304 (N_4304,N_449,N_1900);
nor U4305 (N_4305,N_1849,N_1928);
nand U4306 (N_4306,N_313,N_1048);
and U4307 (N_4307,N_2144,N_1689);
or U4308 (N_4308,N_716,N_177);
and U4309 (N_4309,N_1042,N_1429);
and U4310 (N_4310,N_1764,N_1151);
nor U4311 (N_4311,N_2783,N_1613);
or U4312 (N_4312,N_2456,N_824);
and U4313 (N_4313,N_2285,N_783);
nand U4314 (N_4314,N_259,N_2959);
or U4315 (N_4315,N_2092,N_2896);
and U4316 (N_4316,N_2745,N_2585);
nor U4317 (N_4317,N_2670,N_369);
or U4318 (N_4318,N_413,N_2080);
nor U4319 (N_4319,N_1795,N_1621);
nor U4320 (N_4320,N_1034,N_1108);
nor U4321 (N_4321,N_2239,N_2956);
or U4322 (N_4322,N_1868,N_1813);
nor U4323 (N_4323,N_1587,N_1214);
nand U4324 (N_4324,N_502,N_49);
or U4325 (N_4325,N_1227,N_2545);
and U4326 (N_4326,N_911,N_2741);
nand U4327 (N_4327,N_1491,N_2309);
xor U4328 (N_4328,N_1337,N_1319);
nor U4329 (N_4329,N_1045,N_1407);
and U4330 (N_4330,N_832,N_1815);
or U4331 (N_4331,N_1451,N_148);
nor U4332 (N_4332,N_519,N_895);
and U4333 (N_4333,N_122,N_70);
or U4334 (N_4334,N_2660,N_1678);
nand U4335 (N_4335,N_2424,N_1717);
xor U4336 (N_4336,N_1332,N_742);
and U4337 (N_4337,N_752,N_2933);
nand U4338 (N_4338,N_1116,N_2003);
nor U4339 (N_4339,N_1284,N_310);
and U4340 (N_4340,N_2768,N_343);
or U4341 (N_4341,N_408,N_1652);
nor U4342 (N_4342,N_1027,N_67);
or U4343 (N_4343,N_2306,N_62);
or U4344 (N_4344,N_194,N_335);
nand U4345 (N_4345,N_1039,N_2590);
nand U4346 (N_4346,N_1848,N_29);
or U4347 (N_4347,N_2520,N_644);
and U4348 (N_4348,N_1145,N_544);
nor U4349 (N_4349,N_2175,N_47);
and U4350 (N_4350,N_511,N_196);
xnor U4351 (N_4351,N_74,N_517);
xnor U4352 (N_4352,N_1385,N_882);
nor U4353 (N_4353,N_698,N_597);
nand U4354 (N_4354,N_1814,N_433);
and U4355 (N_4355,N_1317,N_1886);
and U4356 (N_4356,N_353,N_1983);
and U4357 (N_4357,N_2439,N_90);
nor U4358 (N_4358,N_1504,N_703);
nand U4359 (N_4359,N_635,N_874);
nand U4360 (N_4360,N_93,N_1850);
or U4361 (N_4361,N_1422,N_2400);
nor U4362 (N_4362,N_465,N_1053);
and U4363 (N_4363,N_2214,N_2733);
nand U4364 (N_4364,N_2246,N_887);
nand U4365 (N_4365,N_2363,N_773);
and U4366 (N_4366,N_496,N_1930);
and U4367 (N_4367,N_112,N_1838);
nand U4368 (N_4368,N_483,N_162);
nor U4369 (N_4369,N_649,N_1041);
or U4370 (N_4370,N_2259,N_991);
nor U4371 (N_4371,N_26,N_2183);
nand U4372 (N_4372,N_2816,N_356);
and U4373 (N_4373,N_846,N_684);
nor U4374 (N_4374,N_2829,N_390);
nand U4375 (N_4375,N_1642,N_183);
and U4376 (N_4376,N_719,N_1318);
and U4377 (N_4377,N_2597,N_2030);
nor U4378 (N_4378,N_1688,N_38);
and U4379 (N_4379,N_1999,N_1680);
or U4380 (N_4380,N_53,N_859);
and U4381 (N_4381,N_996,N_100);
and U4382 (N_4382,N_1067,N_1604);
nor U4383 (N_4383,N_2017,N_1610);
or U4384 (N_4384,N_804,N_2560);
and U4385 (N_4385,N_223,N_799);
nand U4386 (N_4386,N_2474,N_1452);
and U4387 (N_4387,N_1308,N_2420);
nor U4388 (N_4388,N_2173,N_2658);
or U4389 (N_4389,N_156,N_119);
and U4390 (N_4390,N_1377,N_2236);
or U4391 (N_4391,N_2589,N_971);
or U4392 (N_4392,N_379,N_697);
or U4393 (N_4393,N_457,N_2459);
and U4394 (N_4394,N_1927,N_872);
nor U4395 (N_4395,N_2618,N_557);
or U4396 (N_4396,N_2314,N_392);
or U4397 (N_4397,N_1164,N_1565);
nor U4398 (N_4398,N_2160,N_471);
nor U4399 (N_4399,N_1852,N_2150);
and U4400 (N_4400,N_600,N_380);
and U4401 (N_4401,N_2290,N_2730);
or U4402 (N_4402,N_910,N_1059);
or U4403 (N_4403,N_1884,N_1344);
or U4404 (N_4404,N_2676,N_864);
nand U4405 (N_4405,N_1180,N_2038);
or U4406 (N_4406,N_751,N_2196);
and U4407 (N_4407,N_815,N_2724);
and U4408 (N_4408,N_503,N_988);
and U4409 (N_4409,N_1269,N_1832);
or U4410 (N_4410,N_854,N_4);
or U4411 (N_4411,N_2901,N_98);
nor U4412 (N_4412,N_238,N_1514);
xnor U4413 (N_4413,N_2591,N_686);
or U4414 (N_4414,N_861,N_2944);
nand U4415 (N_4415,N_165,N_2433);
and U4416 (N_4416,N_1538,N_1512);
or U4417 (N_4417,N_2774,N_1495);
nor U4418 (N_4418,N_2473,N_2712);
or U4419 (N_4419,N_349,N_1989);
and U4420 (N_4420,N_2429,N_2413);
nand U4421 (N_4421,N_1169,N_790);
nor U4422 (N_4422,N_110,N_1137);
nor U4423 (N_4423,N_187,N_2861);
or U4424 (N_4424,N_34,N_2544);
or U4425 (N_4425,N_2482,N_849);
and U4426 (N_4426,N_216,N_2504);
nand U4427 (N_4427,N_2976,N_583);
and U4428 (N_4428,N_2857,N_2330);
and U4429 (N_4429,N_1488,N_2061);
or U4430 (N_4430,N_2013,N_494);
nor U4431 (N_4431,N_2089,N_2683);
nand U4432 (N_4432,N_357,N_1361);
nand U4433 (N_4433,N_237,N_2978);
nor U4434 (N_4434,N_2390,N_322);
or U4435 (N_4435,N_768,N_2760);
and U4436 (N_4436,N_1236,N_218);
and U4437 (N_4437,N_891,N_1599);
nor U4438 (N_4438,N_2649,N_660);
nand U4439 (N_4439,N_1430,N_31);
and U4440 (N_4440,N_924,N_150);
and U4441 (N_4441,N_2893,N_616);
nand U4442 (N_4442,N_2548,N_1540);
and U4443 (N_4443,N_1315,N_969);
or U4444 (N_4444,N_1007,N_52);
nor U4445 (N_4445,N_2132,N_2453);
nand U4446 (N_4446,N_2939,N_1152);
nor U4447 (N_4447,N_739,N_25);
and U4448 (N_4448,N_1880,N_2653);
or U4449 (N_4449,N_2265,N_1790);
nand U4450 (N_4450,N_692,N_14);
nand U4451 (N_4451,N_350,N_2890);
nor U4452 (N_4452,N_1281,N_384);
nor U4453 (N_4453,N_1448,N_2378);
nor U4454 (N_4454,N_2039,N_1222);
and U4455 (N_4455,N_1445,N_1716);
nor U4456 (N_4456,N_2170,N_1215);
nand U4457 (N_4457,N_2836,N_1294);
nand U4458 (N_4458,N_185,N_1421);
nand U4459 (N_4459,N_1122,N_485);
or U4460 (N_4460,N_2792,N_1658);
nor U4461 (N_4461,N_1975,N_2969);
or U4462 (N_4462,N_1835,N_693);
nand U4463 (N_4463,N_1481,N_2557);
and U4464 (N_4464,N_564,N_809);
and U4465 (N_4465,N_2635,N_1273);
and U4466 (N_4466,N_900,N_1564);
or U4467 (N_4467,N_84,N_1483);
nand U4468 (N_4468,N_506,N_2335);
nand U4469 (N_4469,N_961,N_2491);
or U4470 (N_4470,N_2908,N_2254);
xor U4471 (N_4471,N_1650,N_2099);
or U4472 (N_4472,N_2368,N_1970);
nor U4473 (N_4473,N_2351,N_2402);
nor U4474 (N_4474,N_960,N_2371);
nor U4475 (N_4475,N_2365,N_317);
nand U4476 (N_4476,N_1190,N_2531);
nor U4477 (N_4477,N_530,N_500);
or U4478 (N_4478,N_2885,N_2707);
nand U4479 (N_4479,N_841,N_2050);
nand U4480 (N_4480,N_2814,N_2043);
nor U4481 (N_4481,N_106,N_236);
nor U4482 (N_4482,N_829,N_478);
nand U4483 (N_4483,N_2701,N_1857);
nor U4484 (N_4484,N_2231,N_2412);
and U4485 (N_4485,N_416,N_717);
nor U4486 (N_4486,N_1594,N_2135);
or U4487 (N_4487,N_1354,N_404);
or U4488 (N_4488,N_2096,N_1823);
nor U4489 (N_4489,N_2362,N_2105);
nand U4490 (N_4490,N_128,N_229);
nor U4491 (N_4491,N_48,N_875);
and U4492 (N_4492,N_585,N_1095);
nand U4493 (N_4493,N_420,N_2079);
nand U4494 (N_4494,N_1206,N_1226);
and U4495 (N_4495,N_479,N_879);
and U4496 (N_4496,N_109,N_1940);
or U4497 (N_4497,N_632,N_2711);
nor U4498 (N_4498,N_1804,N_2777);
nand U4499 (N_4499,N_648,N_666);
or U4500 (N_4500,N_399,N_722);
and U4501 (N_4501,N_1036,N_672);
nand U4502 (N_4502,N_791,N_1728);
nand U4503 (N_4503,N_57,N_81);
nor U4504 (N_4504,N_2147,N_55);
or U4505 (N_4505,N_657,N_1586);
and U4506 (N_4506,N_432,N_464);
or U4507 (N_4507,N_1956,N_603);
nor U4508 (N_4508,N_2662,N_200);
xnor U4509 (N_4509,N_2253,N_637);
or U4510 (N_4510,N_2656,N_1335);
and U4511 (N_4511,N_2745,N_649);
nor U4512 (N_4512,N_2445,N_383);
nand U4513 (N_4513,N_1800,N_2508);
and U4514 (N_4514,N_263,N_1124);
and U4515 (N_4515,N_2176,N_2083);
nand U4516 (N_4516,N_895,N_318);
nand U4517 (N_4517,N_1691,N_388);
or U4518 (N_4518,N_1082,N_2212);
and U4519 (N_4519,N_2254,N_874);
nor U4520 (N_4520,N_616,N_36);
nand U4521 (N_4521,N_2703,N_235);
nor U4522 (N_4522,N_880,N_2488);
nor U4523 (N_4523,N_2256,N_580);
nor U4524 (N_4524,N_2470,N_2110);
nor U4525 (N_4525,N_1338,N_2624);
nand U4526 (N_4526,N_1243,N_1090);
or U4527 (N_4527,N_2140,N_1895);
nor U4528 (N_4528,N_1516,N_1831);
and U4529 (N_4529,N_500,N_2351);
and U4530 (N_4530,N_2521,N_1185);
nor U4531 (N_4531,N_2955,N_1049);
xnor U4532 (N_4532,N_2159,N_1332);
nand U4533 (N_4533,N_2987,N_2379);
and U4534 (N_4534,N_2652,N_2011);
nand U4535 (N_4535,N_1879,N_472);
nor U4536 (N_4536,N_1401,N_1568);
nor U4537 (N_4537,N_906,N_2612);
nor U4538 (N_4538,N_2133,N_322);
nand U4539 (N_4539,N_473,N_1812);
and U4540 (N_4540,N_2292,N_2693);
nand U4541 (N_4541,N_627,N_1015);
nand U4542 (N_4542,N_146,N_2537);
nand U4543 (N_4543,N_1858,N_1771);
or U4544 (N_4544,N_1669,N_1895);
nor U4545 (N_4545,N_267,N_2163);
nor U4546 (N_4546,N_698,N_1173);
nor U4547 (N_4547,N_1845,N_1758);
or U4548 (N_4548,N_640,N_1094);
or U4549 (N_4549,N_2803,N_2715);
nor U4550 (N_4550,N_13,N_2001);
nor U4551 (N_4551,N_716,N_2558);
and U4552 (N_4552,N_1565,N_585);
and U4553 (N_4553,N_19,N_2310);
nor U4554 (N_4554,N_1958,N_2625);
and U4555 (N_4555,N_161,N_1473);
nor U4556 (N_4556,N_1307,N_1047);
nand U4557 (N_4557,N_1995,N_2163);
nor U4558 (N_4558,N_1678,N_2392);
or U4559 (N_4559,N_1194,N_1179);
nor U4560 (N_4560,N_2810,N_156);
and U4561 (N_4561,N_968,N_1905);
nand U4562 (N_4562,N_2911,N_595);
nand U4563 (N_4563,N_2476,N_2320);
and U4564 (N_4564,N_937,N_336);
and U4565 (N_4565,N_2285,N_838);
nand U4566 (N_4566,N_395,N_2899);
nand U4567 (N_4567,N_2762,N_2911);
nand U4568 (N_4568,N_609,N_2620);
nand U4569 (N_4569,N_354,N_2312);
nor U4570 (N_4570,N_1734,N_1844);
or U4571 (N_4571,N_2091,N_1958);
nand U4572 (N_4572,N_2404,N_1010);
and U4573 (N_4573,N_2019,N_180);
and U4574 (N_4574,N_593,N_12);
xnor U4575 (N_4575,N_2833,N_429);
nand U4576 (N_4576,N_858,N_795);
nand U4577 (N_4577,N_421,N_1019);
or U4578 (N_4578,N_866,N_1375);
or U4579 (N_4579,N_1280,N_725);
and U4580 (N_4580,N_787,N_1612);
nand U4581 (N_4581,N_799,N_2123);
nor U4582 (N_4582,N_401,N_1992);
and U4583 (N_4583,N_2115,N_1089);
or U4584 (N_4584,N_835,N_545);
and U4585 (N_4585,N_1359,N_23);
and U4586 (N_4586,N_462,N_1389);
nor U4587 (N_4587,N_2269,N_2063);
or U4588 (N_4588,N_2480,N_303);
or U4589 (N_4589,N_2411,N_545);
and U4590 (N_4590,N_410,N_980);
or U4591 (N_4591,N_1708,N_993);
or U4592 (N_4592,N_451,N_405);
and U4593 (N_4593,N_2818,N_1464);
or U4594 (N_4594,N_1334,N_1112);
and U4595 (N_4595,N_2666,N_672);
and U4596 (N_4596,N_1903,N_1321);
and U4597 (N_4597,N_211,N_297);
nand U4598 (N_4598,N_1102,N_64);
and U4599 (N_4599,N_1159,N_1373);
or U4600 (N_4600,N_837,N_1189);
nor U4601 (N_4601,N_1223,N_2047);
nand U4602 (N_4602,N_1978,N_841);
and U4603 (N_4603,N_1723,N_127);
and U4604 (N_4604,N_1653,N_203);
nor U4605 (N_4605,N_1091,N_1978);
nor U4606 (N_4606,N_1580,N_1328);
nand U4607 (N_4607,N_2479,N_1254);
nor U4608 (N_4608,N_1877,N_1786);
nand U4609 (N_4609,N_204,N_248);
nand U4610 (N_4610,N_2717,N_1511);
xnor U4611 (N_4611,N_747,N_187);
or U4612 (N_4612,N_1259,N_280);
and U4613 (N_4613,N_1597,N_2690);
or U4614 (N_4614,N_2750,N_509);
xor U4615 (N_4615,N_2981,N_1400);
or U4616 (N_4616,N_1299,N_1583);
xnor U4617 (N_4617,N_75,N_723);
nand U4618 (N_4618,N_1908,N_1566);
and U4619 (N_4619,N_1231,N_20);
or U4620 (N_4620,N_143,N_381);
nor U4621 (N_4621,N_2671,N_2778);
nand U4622 (N_4622,N_1627,N_1577);
and U4623 (N_4623,N_2656,N_2451);
nand U4624 (N_4624,N_635,N_2167);
nand U4625 (N_4625,N_1923,N_2328);
nor U4626 (N_4626,N_1018,N_2976);
nor U4627 (N_4627,N_2931,N_1943);
nor U4628 (N_4628,N_1179,N_1436);
and U4629 (N_4629,N_2251,N_1130);
nor U4630 (N_4630,N_2034,N_971);
nand U4631 (N_4631,N_2053,N_256);
nand U4632 (N_4632,N_1523,N_992);
and U4633 (N_4633,N_2298,N_2437);
and U4634 (N_4634,N_400,N_1677);
or U4635 (N_4635,N_2519,N_1946);
nor U4636 (N_4636,N_713,N_617);
nand U4637 (N_4637,N_2018,N_2591);
and U4638 (N_4638,N_1754,N_1091);
and U4639 (N_4639,N_2062,N_746);
nor U4640 (N_4640,N_2122,N_1834);
nor U4641 (N_4641,N_511,N_1836);
nor U4642 (N_4642,N_2811,N_2958);
nand U4643 (N_4643,N_192,N_1314);
nor U4644 (N_4644,N_2510,N_178);
nand U4645 (N_4645,N_2269,N_2957);
or U4646 (N_4646,N_2927,N_1926);
nor U4647 (N_4647,N_245,N_1830);
and U4648 (N_4648,N_917,N_2655);
or U4649 (N_4649,N_598,N_1210);
and U4650 (N_4650,N_1971,N_1991);
nor U4651 (N_4651,N_708,N_216);
xnor U4652 (N_4652,N_234,N_1310);
nand U4653 (N_4653,N_1158,N_534);
nand U4654 (N_4654,N_390,N_1999);
nor U4655 (N_4655,N_1328,N_473);
nand U4656 (N_4656,N_674,N_204);
nand U4657 (N_4657,N_2553,N_841);
and U4658 (N_4658,N_2167,N_2851);
and U4659 (N_4659,N_2445,N_1486);
nor U4660 (N_4660,N_2453,N_854);
or U4661 (N_4661,N_2181,N_1563);
nor U4662 (N_4662,N_978,N_2194);
nor U4663 (N_4663,N_1934,N_1266);
nand U4664 (N_4664,N_1979,N_2523);
nand U4665 (N_4665,N_873,N_1972);
and U4666 (N_4666,N_2153,N_706);
xor U4667 (N_4667,N_1992,N_442);
nand U4668 (N_4668,N_917,N_418);
nand U4669 (N_4669,N_2900,N_994);
nand U4670 (N_4670,N_2022,N_27);
and U4671 (N_4671,N_703,N_1831);
xor U4672 (N_4672,N_1906,N_460);
nor U4673 (N_4673,N_2105,N_321);
or U4674 (N_4674,N_2959,N_487);
and U4675 (N_4675,N_2399,N_2528);
nor U4676 (N_4676,N_2064,N_1514);
or U4677 (N_4677,N_2986,N_376);
or U4678 (N_4678,N_1957,N_1882);
and U4679 (N_4679,N_1310,N_2461);
and U4680 (N_4680,N_413,N_1329);
nor U4681 (N_4681,N_165,N_1129);
or U4682 (N_4682,N_1352,N_789);
nand U4683 (N_4683,N_341,N_26);
and U4684 (N_4684,N_125,N_325);
or U4685 (N_4685,N_1512,N_2881);
and U4686 (N_4686,N_1565,N_243);
xnor U4687 (N_4687,N_1479,N_2342);
or U4688 (N_4688,N_2640,N_2197);
and U4689 (N_4689,N_2541,N_968);
and U4690 (N_4690,N_2713,N_2436);
and U4691 (N_4691,N_1351,N_192);
nand U4692 (N_4692,N_968,N_2867);
and U4693 (N_4693,N_94,N_2882);
or U4694 (N_4694,N_2551,N_1964);
nor U4695 (N_4695,N_1659,N_1357);
or U4696 (N_4696,N_399,N_1835);
and U4697 (N_4697,N_1565,N_911);
nor U4698 (N_4698,N_1693,N_2094);
xnor U4699 (N_4699,N_734,N_778);
or U4700 (N_4700,N_2529,N_1378);
or U4701 (N_4701,N_665,N_1125);
and U4702 (N_4702,N_680,N_1023);
and U4703 (N_4703,N_2351,N_1174);
nor U4704 (N_4704,N_445,N_1723);
or U4705 (N_4705,N_241,N_1786);
and U4706 (N_4706,N_782,N_1031);
nand U4707 (N_4707,N_2486,N_2438);
nand U4708 (N_4708,N_323,N_1039);
nor U4709 (N_4709,N_1564,N_2469);
nor U4710 (N_4710,N_2919,N_310);
nor U4711 (N_4711,N_902,N_2057);
nand U4712 (N_4712,N_481,N_2072);
nor U4713 (N_4713,N_519,N_765);
nand U4714 (N_4714,N_31,N_2566);
or U4715 (N_4715,N_1776,N_2439);
or U4716 (N_4716,N_1702,N_2605);
or U4717 (N_4717,N_874,N_735);
or U4718 (N_4718,N_1580,N_2451);
and U4719 (N_4719,N_2824,N_2000);
and U4720 (N_4720,N_2686,N_191);
nor U4721 (N_4721,N_1149,N_378);
nand U4722 (N_4722,N_1215,N_957);
nor U4723 (N_4723,N_658,N_1946);
and U4724 (N_4724,N_2266,N_464);
nor U4725 (N_4725,N_2512,N_2152);
nor U4726 (N_4726,N_386,N_2547);
nor U4727 (N_4727,N_2916,N_2871);
and U4728 (N_4728,N_916,N_34);
nand U4729 (N_4729,N_1641,N_2327);
or U4730 (N_4730,N_1874,N_1273);
nor U4731 (N_4731,N_982,N_2556);
and U4732 (N_4732,N_232,N_593);
nor U4733 (N_4733,N_918,N_2386);
nor U4734 (N_4734,N_1345,N_2283);
nor U4735 (N_4735,N_2827,N_1646);
and U4736 (N_4736,N_1762,N_1705);
nor U4737 (N_4737,N_796,N_2752);
or U4738 (N_4738,N_79,N_1612);
or U4739 (N_4739,N_1548,N_1996);
or U4740 (N_4740,N_2939,N_970);
or U4741 (N_4741,N_1687,N_1690);
and U4742 (N_4742,N_1030,N_2469);
nand U4743 (N_4743,N_2417,N_1496);
or U4744 (N_4744,N_259,N_59);
and U4745 (N_4745,N_1132,N_404);
or U4746 (N_4746,N_725,N_2825);
or U4747 (N_4747,N_1169,N_2573);
nor U4748 (N_4748,N_15,N_2261);
nand U4749 (N_4749,N_983,N_2651);
or U4750 (N_4750,N_2483,N_2463);
nand U4751 (N_4751,N_557,N_1009);
and U4752 (N_4752,N_1471,N_2179);
and U4753 (N_4753,N_1439,N_833);
or U4754 (N_4754,N_2756,N_2099);
or U4755 (N_4755,N_1097,N_2309);
nand U4756 (N_4756,N_2767,N_577);
nor U4757 (N_4757,N_2984,N_1523);
nor U4758 (N_4758,N_1961,N_448);
nor U4759 (N_4759,N_336,N_1153);
and U4760 (N_4760,N_1325,N_854);
or U4761 (N_4761,N_1326,N_80);
nand U4762 (N_4762,N_140,N_818);
and U4763 (N_4763,N_1214,N_2457);
or U4764 (N_4764,N_1302,N_2514);
nand U4765 (N_4765,N_71,N_802);
and U4766 (N_4766,N_2718,N_1947);
nor U4767 (N_4767,N_1461,N_2949);
nand U4768 (N_4768,N_559,N_642);
nor U4769 (N_4769,N_1549,N_1503);
xnor U4770 (N_4770,N_1834,N_220);
and U4771 (N_4771,N_1047,N_969);
or U4772 (N_4772,N_2312,N_1556);
and U4773 (N_4773,N_1547,N_1620);
or U4774 (N_4774,N_1307,N_2685);
xor U4775 (N_4775,N_1628,N_2397);
xnor U4776 (N_4776,N_323,N_884);
nand U4777 (N_4777,N_375,N_2629);
nand U4778 (N_4778,N_836,N_2576);
nor U4779 (N_4779,N_1215,N_2692);
and U4780 (N_4780,N_1657,N_2434);
nor U4781 (N_4781,N_1728,N_778);
nor U4782 (N_4782,N_11,N_1674);
and U4783 (N_4783,N_2676,N_88);
nor U4784 (N_4784,N_222,N_1327);
or U4785 (N_4785,N_2486,N_2039);
or U4786 (N_4786,N_1608,N_697);
or U4787 (N_4787,N_1713,N_1398);
or U4788 (N_4788,N_1432,N_1851);
or U4789 (N_4789,N_2681,N_2167);
or U4790 (N_4790,N_1075,N_2786);
xnor U4791 (N_4791,N_1173,N_2692);
nor U4792 (N_4792,N_1449,N_1507);
or U4793 (N_4793,N_475,N_783);
nand U4794 (N_4794,N_780,N_1918);
nand U4795 (N_4795,N_399,N_2709);
nand U4796 (N_4796,N_726,N_957);
nor U4797 (N_4797,N_2357,N_1439);
and U4798 (N_4798,N_570,N_1492);
nand U4799 (N_4799,N_1511,N_1491);
or U4800 (N_4800,N_1899,N_1707);
and U4801 (N_4801,N_499,N_1608);
or U4802 (N_4802,N_893,N_1776);
and U4803 (N_4803,N_426,N_488);
nand U4804 (N_4804,N_518,N_506);
or U4805 (N_4805,N_2673,N_770);
nor U4806 (N_4806,N_2528,N_2868);
or U4807 (N_4807,N_2066,N_1082);
nor U4808 (N_4808,N_349,N_2890);
or U4809 (N_4809,N_1695,N_2948);
nand U4810 (N_4810,N_1882,N_589);
nand U4811 (N_4811,N_705,N_2591);
nand U4812 (N_4812,N_1629,N_2003);
xor U4813 (N_4813,N_1547,N_43);
or U4814 (N_4814,N_283,N_2101);
nor U4815 (N_4815,N_466,N_1791);
or U4816 (N_4816,N_2318,N_1538);
and U4817 (N_4817,N_2463,N_2838);
nand U4818 (N_4818,N_869,N_2907);
nor U4819 (N_4819,N_887,N_1164);
nand U4820 (N_4820,N_1018,N_2526);
xor U4821 (N_4821,N_461,N_819);
nand U4822 (N_4822,N_1149,N_755);
nor U4823 (N_4823,N_2367,N_1766);
and U4824 (N_4824,N_1247,N_1282);
or U4825 (N_4825,N_2613,N_2160);
or U4826 (N_4826,N_309,N_1606);
nand U4827 (N_4827,N_2978,N_2563);
or U4828 (N_4828,N_1851,N_2941);
or U4829 (N_4829,N_2361,N_2695);
or U4830 (N_4830,N_1078,N_1967);
or U4831 (N_4831,N_646,N_153);
nor U4832 (N_4832,N_849,N_2881);
and U4833 (N_4833,N_1960,N_1579);
and U4834 (N_4834,N_193,N_2562);
or U4835 (N_4835,N_196,N_1104);
or U4836 (N_4836,N_1726,N_1134);
nand U4837 (N_4837,N_2815,N_2906);
and U4838 (N_4838,N_1863,N_2172);
and U4839 (N_4839,N_2033,N_916);
and U4840 (N_4840,N_2187,N_1733);
nor U4841 (N_4841,N_1282,N_808);
nor U4842 (N_4842,N_1209,N_2861);
xor U4843 (N_4843,N_1803,N_2647);
nor U4844 (N_4844,N_1340,N_1990);
nor U4845 (N_4845,N_1919,N_2558);
nor U4846 (N_4846,N_1798,N_2683);
nand U4847 (N_4847,N_222,N_2699);
and U4848 (N_4848,N_469,N_956);
nor U4849 (N_4849,N_1138,N_521);
and U4850 (N_4850,N_1820,N_268);
or U4851 (N_4851,N_2403,N_972);
nor U4852 (N_4852,N_2490,N_545);
nand U4853 (N_4853,N_2684,N_965);
nor U4854 (N_4854,N_1291,N_1928);
and U4855 (N_4855,N_2297,N_2550);
or U4856 (N_4856,N_1300,N_640);
nand U4857 (N_4857,N_1948,N_2855);
and U4858 (N_4858,N_199,N_2876);
or U4859 (N_4859,N_1266,N_1186);
nor U4860 (N_4860,N_2349,N_2239);
nand U4861 (N_4861,N_365,N_1886);
and U4862 (N_4862,N_2305,N_2614);
nand U4863 (N_4863,N_2057,N_673);
and U4864 (N_4864,N_2440,N_524);
nand U4865 (N_4865,N_288,N_1286);
nor U4866 (N_4866,N_1064,N_1454);
xor U4867 (N_4867,N_388,N_1954);
nand U4868 (N_4868,N_1714,N_1574);
or U4869 (N_4869,N_751,N_453);
and U4870 (N_4870,N_1643,N_1762);
and U4871 (N_4871,N_959,N_838);
nand U4872 (N_4872,N_2389,N_1725);
nor U4873 (N_4873,N_2517,N_2768);
and U4874 (N_4874,N_416,N_1480);
and U4875 (N_4875,N_656,N_662);
nand U4876 (N_4876,N_1139,N_443);
or U4877 (N_4877,N_2324,N_771);
nor U4878 (N_4878,N_2783,N_606);
nor U4879 (N_4879,N_1964,N_44);
nand U4880 (N_4880,N_2346,N_612);
xor U4881 (N_4881,N_226,N_2377);
or U4882 (N_4882,N_1006,N_1132);
or U4883 (N_4883,N_352,N_1223);
nand U4884 (N_4884,N_1985,N_2771);
nor U4885 (N_4885,N_2725,N_1111);
nor U4886 (N_4886,N_2052,N_2348);
nor U4887 (N_4887,N_2325,N_1335);
nand U4888 (N_4888,N_2787,N_852);
and U4889 (N_4889,N_2579,N_1168);
or U4890 (N_4890,N_2853,N_860);
nand U4891 (N_4891,N_544,N_82);
nor U4892 (N_4892,N_368,N_2217);
nand U4893 (N_4893,N_59,N_356);
and U4894 (N_4894,N_2601,N_940);
nand U4895 (N_4895,N_716,N_1106);
and U4896 (N_4896,N_690,N_1258);
and U4897 (N_4897,N_2928,N_2460);
nor U4898 (N_4898,N_239,N_332);
or U4899 (N_4899,N_204,N_2782);
and U4900 (N_4900,N_761,N_465);
nor U4901 (N_4901,N_2318,N_989);
or U4902 (N_4902,N_2802,N_2388);
nand U4903 (N_4903,N_1099,N_2909);
or U4904 (N_4904,N_1141,N_2977);
nand U4905 (N_4905,N_1543,N_896);
nor U4906 (N_4906,N_2260,N_149);
and U4907 (N_4907,N_2144,N_1471);
nor U4908 (N_4908,N_2530,N_152);
and U4909 (N_4909,N_1186,N_38);
nor U4910 (N_4910,N_2575,N_488);
nand U4911 (N_4911,N_2574,N_54);
and U4912 (N_4912,N_581,N_1608);
nand U4913 (N_4913,N_212,N_2272);
nor U4914 (N_4914,N_2321,N_2609);
or U4915 (N_4915,N_923,N_430);
nor U4916 (N_4916,N_2227,N_1101);
and U4917 (N_4917,N_2485,N_156);
or U4918 (N_4918,N_673,N_186);
nor U4919 (N_4919,N_574,N_11);
xor U4920 (N_4920,N_1491,N_2180);
nand U4921 (N_4921,N_1857,N_1254);
nor U4922 (N_4922,N_389,N_1774);
nand U4923 (N_4923,N_2958,N_256);
nor U4924 (N_4924,N_2574,N_484);
and U4925 (N_4925,N_1015,N_2739);
and U4926 (N_4926,N_68,N_837);
nand U4927 (N_4927,N_2595,N_1402);
or U4928 (N_4928,N_2646,N_929);
nand U4929 (N_4929,N_789,N_2871);
nor U4930 (N_4930,N_1204,N_474);
nor U4931 (N_4931,N_709,N_1065);
nand U4932 (N_4932,N_2063,N_1035);
nand U4933 (N_4933,N_2522,N_2509);
xor U4934 (N_4934,N_2208,N_976);
and U4935 (N_4935,N_214,N_1599);
nor U4936 (N_4936,N_1329,N_589);
nor U4937 (N_4937,N_1115,N_2183);
nand U4938 (N_4938,N_1389,N_2782);
or U4939 (N_4939,N_2396,N_1113);
nor U4940 (N_4940,N_2044,N_1595);
nand U4941 (N_4941,N_2924,N_2844);
nor U4942 (N_4942,N_2639,N_2266);
nor U4943 (N_4943,N_877,N_2126);
xnor U4944 (N_4944,N_14,N_1958);
and U4945 (N_4945,N_99,N_1781);
nor U4946 (N_4946,N_2803,N_2830);
and U4947 (N_4947,N_1432,N_515);
and U4948 (N_4948,N_2130,N_780);
or U4949 (N_4949,N_507,N_1361);
nand U4950 (N_4950,N_2451,N_1544);
nand U4951 (N_4951,N_434,N_2077);
nor U4952 (N_4952,N_499,N_193);
or U4953 (N_4953,N_2877,N_2337);
or U4954 (N_4954,N_2083,N_1617);
xor U4955 (N_4955,N_352,N_117);
nor U4956 (N_4956,N_2516,N_1655);
nor U4957 (N_4957,N_1419,N_606);
or U4958 (N_4958,N_2432,N_244);
nand U4959 (N_4959,N_804,N_1596);
or U4960 (N_4960,N_2385,N_569);
nor U4961 (N_4961,N_913,N_73);
nand U4962 (N_4962,N_2919,N_1627);
or U4963 (N_4963,N_2162,N_2684);
nand U4964 (N_4964,N_1570,N_1118);
or U4965 (N_4965,N_2442,N_126);
and U4966 (N_4966,N_2702,N_708);
nor U4967 (N_4967,N_83,N_2061);
or U4968 (N_4968,N_1386,N_2841);
nor U4969 (N_4969,N_1416,N_2645);
nor U4970 (N_4970,N_14,N_517);
nand U4971 (N_4971,N_2949,N_85);
nor U4972 (N_4972,N_1663,N_2101);
nor U4973 (N_4973,N_1978,N_576);
or U4974 (N_4974,N_119,N_2200);
nor U4975 (N_4975,N_285,N_330);
nor U4976 (N_4976,N_1797,N_1495);
and U4977 (N_4977,N_2464,N_2981);
or U4978 (N_4978,N_660,N_1151);
nor U4979 (N_4979,N_1609,N_2203);
nor U4980 (N_4980,N_1965,N_863);
nor U4981 (N_4981,N_2362,N_1526);
and U4982 (N_4982,N_341,N_2097);
and U4983 (N_4983,N_2996,N_248);
nor U4984 (N_4984,N_165,N_1610);
nor U4985 (N_4985,N_2257,N_1967);
nor U4986 (N_4986,N_669,N_930);
or U4987 (N_4987,N_2040,N_1627);
nor U4988 (N_4988,N_667,N_2136);
and U4989 (N_4989,N_2741,N_2995);
and U4990 (N_4990,N_2440,N_2227);
nand U4991 (N_4991,N_1649,N_1281);
and U4992 (N_4992,N_805,N_1519);
nand U4993 (N_4993,N_2411,N_920);
or U4994 (N_4994,N_1182,N_967);
nor U4995 (N_4995,N_1774,N_597);
nor U4996 (N_4996,N_1539,N_1598);
and U4997 (N_4997,N_2871,N_1744);
nor U4998 (N_4998,N_1026,N_654);
or U4999 (N_4999,N_2731,N_2966);
or U5000 (N_5000,N_1093,N_1013);
or U5001 (N_5001,N_2046,N_836);
nor U5002 (N_5002,N_668,N_600);
nand U5003 (N_5003,N_2468,N_215);
or U5004 (N_5004,N_466,N_2676);
or U5005 (N_5005,N_2438,N_109);
and U5006 (N_5006,N_2650,N_1593);
or U5007 (N_5007,N_2461,N_53);
nand U5008 (N_5008,N_337,N_2656);
or U5009 (N_5009,N_2872,N_1963);
and U5010 (N_5010,N_2401,N_2118);
and U5011 (N_5011,N_1315,N_867);
nor U5012 (N_5012,N_1021,N_209);
and U5013 (N_5013,N_1855,N_141);
nor U5014 (N_5014,N_2021,N_2983);
or U5015 (N_5015,N_1644,N_246);
nor U5016 (N_5016,N_2669,N_2167);
or U5017 (N_5017,N_2127,N_1870);
nand U5018 (N_5018,N_1483,N_2045);
or U5019 (N_5019,N_2007,N_796);
or U5020 (N_5020,N_832,N_1333);
nand U5021 (N_5021,N_1709,N_686);
nand U5022 (N_5022,N_2922,N_860);
nand U5023 (N_5023,N_870,N_41);
and U5024 (N_5024,N_1260,N_2368);
or U5025 (N_5025,N_439,N_490);
and U5026 (N_5026,N_583,N_1304);
nor U5027 (N_5027,N_1061,N_1611);
and U5028 (N_5028,N_1457,N_214);
nor U5029 (N_5029,N_611,N_2505);
nor U5030 (N_5030,N_2477,N_943);
nand U5031 (N_5031,N_1189,N_343);
and U5032 (N_5032,N_36,N_529);
nand U5033 (N_5033,N_2022,N_1348);
nor U5034 (N_5034,N_871,N_344);
nor U5035 (N_5035,N_1037,N_1496);
and U5036 (N_5036,N_672,N_1586);
or U5037 (N_5037,N_2391,N_1896);
nand U5038 (N_5038,N_2041,N_1584);
or U5039 (N_5039,N_2103,N_765);
nor U5040 (N_5040,N_194,N_1596);
nand U5041 (N_5041,N_1916,N_2562);
and U5042 (N_5042,N_770,N_1798);
nand U5043 (N_5043,N_486,N_1025);
and U5044 (N_5044,N_1818,N_531);
and U5045 (N_5045,N_2960,N_300);
nand U5046 (N_5046,N_325,N_247);
and U5047 (N_5047,N_1202,N_289);
and U5048 (N_5048,N_2861,N_870);
or U5049 (N_5049,N_345,N_216);
nor U5050 (N_5050,N_728,N_1458);
and U5051 (N_5051,N_2621,N_112);
nand U5052 (N_5052,N_2131,N_894);
nand U5053 (N_5053,N_1049,N_81);
nor U5054 (N_5054,N_2107,N_97);
nand U5055 (N_5055,N_2064,N_180);
or U5056 (N_5056,N_2183,N_2538);
or U5057 (N_5057,N_1213,N_680);
nand U5058 (N_5058,N_450,N_1833);
and U5059 (N_5059,N_2906,N_2944);
nor U5060 (N_5060,N_2502,N_2603);
nor U5061 (N_5061,N_2634,N_798);
nor U5062 (N_5062,N_2808,N_1282);
and U5063 (N_5063,N_2252,N_669);
nand U5064 (N_5064,N_36,N_2677);
and U5065 (N_5065,N_1411,N_2708);
nor U5066 (N_5066,N_1236,N_1623);
nand U5067 (N_5067,N_1473,N_2435);
nor U5068 (N_5068,N_1360,N_2377);
or U5069 (N_5069,N_6,N_1436);
nor U5070 (N_5070,N_2374,N_2879);
nor U5071 (N_5071,N_2523,N_2191);
nand U5072 (N_5072,N_1958,N_774);
or U5073 (N_5073,N_870,N_2593);
nor U5074 (N_5074,N_574,N_861);
nor U5075 (N_5075,N_2222,N_686);
nand U5076 (N_5076,N_540,N_546);
nor U5077 (N_5077,N_1961,N_2302);
nand U5078 (N_5078,N_1598,N_1059);
nand U5079 (N_5079,N_1482,N_2279);
nor U5080 (N_5080,N_1406,N_2930);
and U5081 (N_5081,N_1604,N_369);
and U5082 (N_5082,N_2101,N_362);
or U5083 (N_5083,N_1492,N_880);
nor U5084 (N_5084,N_1847,N_146);
nand U5085 (N_5085,N_2383,N_2585);
and U5086 (N_5086,N_1373,N_512);
and U5087 (N_5087,N_1140,N_2077);
nand U5088 (N_5088,N_2682,N_1825);
or U5089 (N_5089,N_1261,N_1693);
nor U5090 (N_5090,N_2062,N_2765);
nand U5091 (N_5091,N_293,N_2724);
nand U5092 (N_5092,N_258,N_721);
nand U5093 (N_5093,N_1596,N_1536);
nand U5094 (N_5094,N_1854,N_2324);
or U5095 (N_5095,N_1738,N_11);
and U5096 (N_5096,N_2442,N_2264);
and U5097 (N_5097,N_2323,N_2241);
and U5098 (N_5098,N_837,N_1758);
or U5099 (N_5099,N_1322,N_1555);
nand U5100 (N_5100,N_2195,N_1965);
or U5101 (N_5101,N_1603,N_551);
and U5102 (N_5102,N_501,N_780);
nand U5103 (N_5103,N_216,N_2092);
or U5104 (N_5104,N_1872,N_1890);
and U5105 (N_5105,N_2881,N_1968);
nand U5106 (N_5106,N_2459,N_1646);
and U5107 (N_5107,N_2305,N_597);
nor U5108 (N_5108,N_142,N_2410);
nor U5109 (N_5109,N_442,N_1148);
xnor U5110 (N_5110,N_2869,N_2543);
nor U5111 (N_5111,N_1973,N_2552);
nor U5112 (N_5112,N_1585,N_656);
nor U5113 (N_5113,N_200,N_1481);
or U5114 (N_5114,N_1636,N_2314);
and U5115 (N_5115,N_1532,N_2897);
nand U5116 (N_5116,N_138,N_1534);
nand U5117 (N_5117,N_2675,N_986);
nor U5118 (N_5118,N_2060,N_1699);
nor U5119 (N_5119,N_2080,N_2010);
and U5120 (N_5120,N_180,N_1585);
or U5121 (N_5121,N_2480,N_973);
nand U5122 (N_5122,N_1318,N_1930);
or U5123 (N_5123,N_1116,N_823);
or U5124 (N_5124,N_783,N_1199);
nor U5125 (N_5125,N_852,N_1988);
nand U5126 (N_5126,N_2040,N_1791);
nor U5127 (N_5127,N_737,N_2212);
nor U5128 (N_5128,N_1819,N_2094);
nor U5129 (N_5129,N_2529,N_1055);
and U5130 (N_5130,N_1264,N_99);
or U5131 (N_5131,N_1211,N_2378);
nor U5132 (N_5132,N_2984,N_1505);
nor U5133 (N_5133,N_2766,N_1385);
nor U5134 (N_5134,N_1516,N_1321);
nand U5135 (N_5135,N_2915,N_70);
nor U5136 (N_5136,N_2574,N_2909);
nand U5137 (N_5137,N_1977,N_272);
and U5138 (N_5138,N_2618,N_2811);
nand U5139 (N_5139,N_685,N_1847);
xnor U5140 (N_5140,N_2109,N_2197);
and U5141 (N_5141,N_2804,N_2235);
or U5142 (N_5142,N_2718,N_2141);
and U5143 (N_5143,N_1021,N_2165);
and U5144 (N_5144,N_717,N_2712);
nor U5145 (N_5145,N_2821,N_13);
and U5146 (N_5146,N_557,N_2445);
nand U5147 (N_5147,N_610,N_909);
nor U5148 (N_5148,N_2163,N_640);
or U5149 (N_5149,N_524,N_2804);
and U5150 (N_5150,N_2406,N_1245);
and U5151 (N_5151,N_1617,N_2356);
and U5152 (N_5152,N_2524,N_168);
and U5153 (N_5153,N_970,N_1365);
nor U5154 (N_5154,N_805,N_330);
xor U5155 (N_5155,N_653,N_826);
or U5156 (N_5156,N_868,N_610);
or U5157 (N_5157,N_1657,N_1849);
and U5158 (N_5158,N_2207,N_535);
and U5159 (N_5159,N_1461,N_947);
or U5160 (N_5160,N_5,N_2768);
or U5161 (N_5161,N_52,N_2747);
nand U5162 (N_5162,N_2632,N_1338);
and U5163 (N_5163,N_2097,N_347);
and U5164 (N_5164,N_2674,N_430);
nand U5165 (N_5165,N_1891,N_2775);
and U5166 (N_5166,N_1669,N_1146);
nand U5167 (N_5167,N_1269,N_525);
and U5168 (N_5168,N_1458,N_2212);
nand U5169 (N_5169,N_2724,N_1687);
or U5170 (N_5170,N_2166,N_1453);
nand U5171 (N_5171,N_558,N_780);
nor U5172 (N_5172,N_963,N_1760);
or U5173 (N_5173,N_1465,N_1471);
nand U5174 (N_5174,N_2024,N_2893);
nor U5175 (N_5175,N_771,N_1417);
or U5176 (N_5176,N_2733,N_2342);
nor U5177 (N_5177,N_1676,N_1080);
or U5178 (N_5178,N_1271,N_682);
nor U5179 (N_5179,N_975,N_161);
and U5180 (N_5180,N_1993,N_2618);
nor U5181 (N_5181,N_2488,N_1647);
nand U5182 (N_5182,N_581,N_1170);
nor U5183 (N_5183,N_1798,N_2540);
or U5184 (N_5184,N_949,N_1533);
or U5185 (N_5185,N_1105,N_1873);
nor U5186 (N_5186,N_2742,N_651);
nor U5187 (N_5187,N_605,N_1226);
nand U5188 (N_5188,N_1889,N_1975);
or U5189 (N_5189,N_2934,N_1254);
and U5190 (N_5190,N_1929,N_1075);
nor U5191 (N_5191,N_1072,N_608);
nor U5192 (N_5192,N_1002,N_1352);
nor U5193 (N_5193,N_224,N_549);
or U5194 (N_5194,N_760,N_1621);
nor U5195 (N_5195,N_1331,N_2624);
nand U5196 (N_5196,N_954,N_2126);
or U5197 (N_5197,N_893,N_1497);
and U5198 (N_5198,N_1488,N_1419);
nand U5199 (N_5199,N_2060,N_1636);
and U5200 (N_5200,N_2671,N_1835);
or U5201 (N_5201,N_12,N_622);
nor U5202 (N_5202,N_132,N_89);
nand U5203 (N_5203,N_1175,N_789);
and U5204 (N_5204,N_1500,N_516);
nor U5205 (N_5205,N_1421,N_1034);
and U5206 (N_5206,N_324,N_1347);
nand U5207 (N_5207,N_1915,N_391);
and U5208 (N_5208,N_2661,N_217);
nor U5209 (N_5209,N_2590,N_133);
or U5210 (N_5210,N_1451,N_2592);
nor U5211 (N_5211,N_22,N_2958);
or U5212 (N_5212,N_1169,N_2968);
nand U5213 (N_5213,N_1917,N_537);
or U5214 (N_5214,N_2823,N_1432);
or U5215 (N_5215,N_1437,N_667);
nor U5216 (N_5216,N_2326,N_2777);
nor U5217 (N_5217,N_1592,N_1835);
nor U5218 (N_5218,N_496,N_2108);
nor U5219 (N_5219,N_2031,N_809);
or U5220 (N_5220,N_228,N_2174);
nor U5221 (N_5221,N_1847,N_644);
or U5222 (N_5222,N_1058,N_289);
xor U5223 (N_5223,N_710,N_2175);
and U5224 (N_5224,N_2812,N_232);
and U5225 (N_5225,N_2375,N_1106);
and U5226 (N_5226,N_1759,N_1883);
nor U5227 (N_5227,N_2783,N_490);
or U5228 (N_5228,N_652,N_379);
nand U5229 (N_5229,N_942,N_2803);
nor U5230 (N_5230,N_855,N_253);
nor U5231 (N_5231,N_1319,N_714);
and U5232 (N_5232,N_755,N_2195);
nand U5233 (N_5233,N_1540,N_126);
or U5234 (N_5234,N_2537,N_1706);
or U5235 (N_5235,N_1257,N_2050);
and U5236 (N_5236,N_2300,N_262);
and U5237 (N_5237,N_2355,N_1127);
and U5238 (N_5238,N_830,N_2646);
nor U5239 (N_5239,N_2223,N_2895);
and U5240 (N_5240,N_651,N_1443);
xnor U5241 (N_5241,N_1785,N_2184);
nand U5242 (N_5242,N_585,N_143);
or U5243 (N_5243,N_2814,N_2272);
or U5244 (N_5244,N_546,N_719);
nor U5245 (N_5245,N_484,N_2483);
or U5246 (N_5246,N_939,N_1324);
nand U5247 (N_5247,N_1867,N_2957);
nand U5248 (N_5248,N_2641,N_2187);
nand U5249 (N_5249,N_595,N_686);
and U5250 (N_5250,N_1587,N_1431);
nand U5251 (N_5251,N_2135,N_2074);
nand U5252 (N_5252,N_2434,N_557);
nor U5253 (N_5253,N_1721,N_687);
nor U5254 (N_5254,N_249,N_157);
nand U5255 (N_5255,N_2078,N_946);
and U5256 (N_5256,N_169,N_2874);
nor U5257 (N_5257,N_375,N_175);
and U5258 (N_5258,N_2960,N_748);
nand U5259 (N_5259,N_2098,N_2671);
and U5260 (N_5260,N_1786,N_1421);
or U5261 (N_5261,N_793,N_388);
or U5262 (N_5262,N_2886,N_2455);
or U5263 (N_5263,N_1163,N_1482);
nor U5264 (N_5264,N_1906,N_891);
nor U5265 (N_5265,N_2328,N_1935);
and U5266 (N_5266,N_993,N_2413);
nor U5267 (N_5267,N_2352,N_84);
and U5268 (N_5268,N_1009,N_2303);
nand U5269 (N_5269,N_617,N_215);
nor U5270 (N_5270,N_90,N_2139);
xor U5271 (N_5271,N_1737,N_509);
or U5272 (N_5272,N_2884,N_505);
nor U5273 (N_5273,N_1046,N_1189);
nor U5274 (N_5274,N_2471,N_1437);
nand U5275 (N_5275,N_30,N_925);
nor U5276 (N_5276,N_2914,N_2166);
or U5277 (N_5277,N_2993,N_2515);
nor U5278 (N_5278,N_111,N_1521);
nor U5279 (N_5279,N_773,N_2033);
and U5280 (N_5280,N_2913,N_694);
nand U5281 (N_5281,N_803,N_1946);
or U5282 (N_5282,N_456,N_2067);
or U5283 (N_5283,N_532,N_581);
and U5284 (N_5284,N_2628,N_2414);
and U5285 (N_5285,N_702,N_1593);
nand U5286 (N_5286,N_1413,N_1601);
xnor U5287 (N_5287,N_2079,N_1376);
and U5288 (N_5288,N_1833,N_157);
and U5289 (N_5289,N_427,N_1882);
and U5290 (N_5290,N_2477,N_320);
and U5291 (N_5291,N_517,N_1644);
nand U5292 (N_5292,N_2265,N_209);
or U5293 (N_5293,N_2115,N_1936);
nand U5294 (N_5294,N_2883,N_1152);
nand U5295 (N_5295,N_2584,N_1792);
nand U5296 (N_5296,N_2497,N_2059);
nand U5297 (N_5297,N_1946,N_934);
nor U5298 (N_5298,N_1841,N_2435);
and U5299 (N_5299,N_2057,N_1521);
nor U5300 (N_5300,N_1056,N_1189);
and U5301 (N_5301,N_2446,N_768);
and U5302 (N_5302,N_1415,N_2077);
nor U5303 (N_5303,N_1382,N_2498);
and U5304 (N_5304,N_156,N_1363);
and U5305 (N_5305,N_1132,N_2195);
or U5306 (N_5306,N_762,N_2085);
or U5307 (N_5307,N_2921,N_342);
or U5308 (N_5308,N_385,N_328);
nand U5309 (N_5309,N_2572,N_1066);
or U5310 (N_5310,N_553,N_590);
nand U5311 (N_5311,N_2861,N_2858);
nand U5312 (N_5312,N_1815,N_1190);
or U5313 (N_5313,N_1789,N_1074);
and U5314 (N_5314,N_2312,N_2517);
nor U5315 (N_5315,N_1191,N_2788);
nand U5316 (N_5316,N_2781,N_1610);
nor U5317 (N_5317,N_470,N_2320);
and U5318 (N_5318,N_1300,N_1033);
nand U5319 (N_5319,N_701,N_815);
nand U5320 (N_5320,N_1849,N_2009);
or U5321 (N_5321,N_2464,N_485);
nand U5322 (N_5322,N_2933,N_22);
nand U5323 (N_5323,N_1366,N_1808);
nor U5324 (N_5324,N_2941,N_1916);
nor U5325 (N_5325,N_815,N_2456);
and U5326 (N_5326,N_1045,N_2771);
or U5327 (N_5327,N_378,N_165);
and U5328 (N_5328,N_399,N_2947);
xnor U5329 (N_5329,N_2511,N_1785);
nand U5330 (N_5330,N_1563,N_2122);
and U5331 (N_5331,N_804,N_2378);
nor U5332 (N_5332,N_726,N_998);
or U5333 (N_5333,N_1616,N_2731);
nand U5334 (N_5334,N_1139,N_864);
and U5335 (N_5335,N_99,N_562);
nor U5336 (N_5336,N_525,N_2976);
nor U5337 (N_5337,N_275,N_571);
or U5338 (N_5338,N_2944,N_1715);
nor U5339 (N_5339,N_2967,N_1042);
or U5340 (N_5340,N_2142,N_436);
and U5341 (N_5341,N_2926,N_530);
nor U5342 (N_5342,N_2493,N_1622);
and U5343 (N_5343,N_2889,N_2529);
or U5344 (N_5344,N_2494,N_639);
nor U5345 (N_5345,N_2923,N_510);
nand U5346 (N_5346,N_1033,N_2405);
nand U5347 (N_5347,N_2486,N_2757);
and U5348 (N_5348,N_753,N_2620);
or U5349 (N_5349,N_162,N_1281);
and U5350 (N_5350,N_331,N_2456);
or U5351 (N_5351,N_54,N_2871);
nor U5352 (N_5352,N_531,N_2721);
and U5353 (N_5353,N_1246,N_966);
nand U5354 (N_5354,N_2020,N_1707);
nand U5355 (N_5355,N_67,N_1413);
or U5356 (N_5356,N_2053,N_2655);
nor U5357 (N_5357,N_2320,N_1683);
xor U5358 (N_5358,N_2741,N_2815);
and U5359 (N_5359,N_110,N_743);
and U5360 (N_5360,N_1004,N_2906);
nor U5361 (N_5361,N_155,N_530);
xor U5362 (N_5362,N_2966,N_1988);
nor U5363 (N_5363,N_2398,N_2548);
and U5364 (N_5364,N_2578,N_902);
or U5365 (N_5365,N_2569,N_1499);
and U5366 (N_5366,N_2336,N_2023);
or U5367 (N_5367,N_170,N_664);
and U5368 (N_5368,N_2328,N_798);
nand U5369 (N_5369,N_1570,N_1023);
nor U5370 (N_5370,N_2126,N_793);
nand U5371 (N_5371,N_2268,N_82);
nand U5372 (N_5372,N_372,N_2901);
nor U5373 (N_5373,N_679,N_1116);
and U5374 (N_5374,N_656,N_2286);
or U5375 (N_5375,N_1116,N_1090);
and U5376 (N_5376,N_1574,N_967);
nand U5377 (N_5377,N_831,N_448);
xnor U5378 (N_5378,N_1618,N_2346);
xor U5379 (N_5379,N_1937,N_1644);
nor U5380 (N_5380,N_76,N_263);
nor U5381 (N_5381,N_897,N_2172);
and U5382 (N_5382,N_1395,N_2235);
and U5383 (N_5383,N_2685,N_2833);
nand U5384 (N_5384,N_2995,N_953);
nor U5385 (N_5385,N_2670,N_2576);
and U5386 (N_5386,N_1034,N_1064);
nand U5387 (N_5387,N_1826,N_1809);
nand U5388 (N_5388,N_1784,N_2982);
nand U5389 (N_5389,N_1021,N_665);
nor U5390 (N_5390,N_169,N_742);
or U5391 (N_5391,N_2343,N_1054);
or U5392 (N_5392,N_1222,N_404);
or U5393 (N_5393,N_281,N_1229);
or U5394 (N_5394,N_1961,N_1852);
and U5395 (N_5395,N_1204,N_2557);
and U5396 (N_5396,N_916,N_2546);
nor U5397 (N_5397,N_595,N_2564);
and U5398 (N_5398,N_2256,N_1000);
nor U5399 (N_5399,N_1205,N_630);
and U5400 (N_5400,N_1761,N_476);
or U5401 (N_5401,N_884,N_109);
xor U5402 (N_5402,N_2070,N_2103);
or U5403 (N_5403,N_2258,N_2974);
and U5404 (N_5404,N_1613,N_810);
and U5405 (N_5405,N_2380,N_2763);
nand U5406 (N_5406,N_968,N_2984);
or U5407 (N_5407,N_1028,N_381);
nand U5408 (N_5408,N_1618,N_181);
nand U5409 (N_5409,N_2918,N_2647);
and U5410 (N_5410,N_1799,N_76);
nand U5411 (N_5411,N_1410,N_17);
nand U5412 (N_5412,N_2165,N_2969);
and U5413 (N_5413,N_1018,N_2009);
and U5414 (N_5414,N_154,N_1732);
or U5415 (N_5415,N_2790,N_2008);
and U5416 (N_5416,N_641,N_1695);
or U5417 (N_5417,N_693,N_1441);
or U5418 (N_5418,N_956,N_1115);
and U5419 (N_5419,N_545,N_1230);
or U5420 (N_5420,N_1785,N_910);
nor U5421 (N_5421,N_1408,N_347);
and U5422 (N_5422,N_1983,N_973);
nor U5423 (N_5423,N_1231,N_1517);
or U5424 (N_5424,N_1604,N_476);
or U5425 (N_5425,N_1186,N_1356);
and U5426 (N_5426,N_1485,N_1887);
or U5427 (N_5427,N_2765,N_382);
or U5428 (N_5428,N_105,N_2637);
and U5429 (N_5429,N_761,N_497);
nand U5430 (N_5430,N_1714,N_408);
nand U5431 (N_5431,N_328,N_529);
xor U5432 (N_5432,N_2976,N_2280);
or U5433 (N_5433,N_2216,N_1031);
nor U5434 (N_5434,N_1829,N_815);
and U5435 (N_5435,N_292,N_1283);
and U5436 (N_5436,N_1306,N_939);
or U5437 (N_5437,N_2770,N_497);
nand U5438 (N_5438,N_2530,N_1106);
or U5439 (N_5439,N_210,N_2781);
or U5440 (N_5440,N_2673,N_444);
nand U5441 (N_5441,N_973,N_1894);
or U5442 (N_5442,N_199,N_1388);
or U5443 (N_5443,N_1000,N_1765);
or U5444 (N_5444,N_603,N_1715);
or U5445 (N_5445,N_2086,N_2107);
nor U5446 (N_5446,N_2231,N_1130);
nor U5447 (N_5447,N_323,N_720);
xnor U5448 (N_5448,N_1946,N_668);
and U5449 (N_5449,N_681,N_2159);
nand U5450 (N_5450,N_2482,N_2901);
or U5451 (N_5451,N_1209,N_1291);
nand U5452 (N_5452,N_1522,N_271);
and U5453 (N_5453,N_345,N_974);
and U5454 (N_5454,N_2692,N_1205);
or U5455 (N_5455,N_553,N_255);
or U5456 (N_5456,N_1664,N_182);
or U5457 (N_5457,N_1035,N_1495);
and U5458 (N_5458,N_2892,N_1508);
or U5459 (N_5459,N_1374,N_1059);
nand U5460 (N_5460,N_497,N_744);
nor U5461 (N_5461,N_46,N_2135);
nand U5462 (N_5462,N_2763,N_22);
or U5463 (N_5463,N_1416,N_410);
nand U5464 (N_5464,N_1367,N_1655);
nor U5465 (N_5465,N_2810,N_2423);
and U5466 (N_5466,N_2342,N_2056);
nand U5467 (N_5467,N_79,N_990);
or U5468 (N_5468,N_1364,N_868);
or U5469 (N_5469,N_940,N_654);
and U5470 (N_5470,N_300,N_612);
nor U5471 (N_5471,N_355,N_140);
and U5472 (N_5472,N_2815,N_1047);
nand U5473 (N_5473,N_1831,N_1112);
and U5474 (N_5474,N_414,N_351);
nor U5475 (N_5475,N_932,N_1353);
or U5476 (N_5476,N_832,N_865);
nor U5477 (N_5477,N_663,N_2474);
and U5478 (N_5478,N_412,N_1684);
xor U5479 (N_5479,N_501,N_1883);
nor U5480 (N_5480,N_452,N_1732);
nor U5481 (N_5481,N_736,N_1109);
nand U5482 (N_5482,N_1773,N_1997);
nor U5483 (N_5483,N_812,N_2340);
or U5484 (N_5484,N_2307,N_1067);
and U5485 (N_5485,N_1376,N_1055);
and U5486 (N_5486,N_351,N_1610);
or U5487 (N_5487,N_1096,N_2509);
nand U5488 (N_5488,N_102,N_773);
nor U5489 (N_5489,N_1823,N_1409);
nor U5490 (N_5490,N_1943,N_104);
nand U5491 (N_5491,N_2525,N_778);
and U5492 (N_5492,N_301,N_1775);
nor U5493 (N_5493,N_1578,N_865);
nor U5494 (N_5494,N_2666,N_2756);
and U5495 (N_5495,N_288,N_153);
nand U5496 (N_5496,N_1481,N_2536);
and U5497 (N_5497,N_2580,N_286);
and U5498 (N_5498,N_1331,N_1703);
and U5499 (N_5499,N_2998,N_2687);
nand U5500 (N_5500,N_18,N_1020);
or U5501 (N_5501,N_819,N_60);
nand U5502 (N_5502,N_2530,N_1622);
and U5503 (N_5503,N_1534,N_2676);
and U5504 (N_5504,N_133,N_129);
and U5505 (N_5505,N_229,N_2481);
or U5506 (N_5506,N_508,N_851);
nor U5507 (N_5507,N_2011,N_842);
and U5508 (N_5508,N_386,N_134);
nand U5509 (N_5509,N_1610,N_2439);
nor U5510 (N_5510,N_2772,N_2175);
nand U5511 (N_5511,N_1100,N_1461);
or U5512 (N_5512,N_1595,N_2983);
or U5513 (N_5513,N_1962,N_1698);
nor U5514 (N_5514,N_90,N_867);
and U5515 (N_5515,N_156,N_1116);
nand U5516 (N_5516,N_2418,N_2585);
nor U5517 (N_5517,N_2665,N_2043);
nand U5518 (N_5518,N_1794,N_206);
nor U5519 (N_5519,N_1829,N_1469);
nand U5520 (N_5520,N_2328,N_411);
or U5521 (N_5521,N_2370,N_1608);
or U5522 (N_5522,N_2851,N_1860);
or U5523 (N_5523,N_578,N_1447);
nor U5524 (N_5524,N_499,N_1809);
nand U5525 (N_5525,N_518,N_52);
nor U5526 (N_5526,N_2186,N_1106);
nor U5527 (N_5527,N_1020,N_2962);
nor U5528 (N_5528,N_2677,N_2894);
nor U5529 (N_5529,N_892,N_2486);
or U5530 (N_5530,N_1485,N_1683);
and U5531 (N_5531,N_1139,N_2400);
or U5532 (N_5532,N_158,N_748);
nand U5533 (N_5533,N_131,N_1335);
nand U5534 (N_5534,N_375,N_613);
nor U5535 (N_5535,N_1925,N_951);
nand U5536 (N_5536,N_2907,N_2669);
or U5537 (N_5537,N_2106,N_2135);
or U5538 (N_5538,N_1493,N_299);
nor U5539 (N_5539,N_2693,N_1460);
nand U5540 (N_5540,N_1655,N_2178);
nor U5541 (N_5541,N_305,N_2220);
xnor U5542 (N_5542,N_800,N_985);
and U5543 (N_5543,N_770,N_1286);
and U5544 (N_5544,N_1455,N_685);
or U5545 (N_5545,N_2222,N_2979);
nor U5546 (N_5546,N_797,N_2465);
nand U5547 (N_5547,N_2581,N_2442);
xnor U5548 (N_5548,N_878,N_2960);
nand U5549 (N_5549,N_2389,N_1152);
nor U5550 (N_5550,N_866,N_1248);
nor U5551 (N_5551,N_1483,N_678);
nand U5552 (N_5552,N_2854,N_132);
and U5553 (N_5553,N_2718,N_2987);
and U5554 (N_5554,N_1882,N_15);
nand U5555 (N_5555,N_2064,N_1925);
or U5556 (N_5556,N_2966,N_1606);
nand U5557 (N_5557,N_717,N_1043);
or U5558 (N_5558,N_2557,N_446);
nor U5559 (N_5559,N_16,N_2418);
and U5560 (N_5560,N_2320,N_1849);
nand U5561 (N_5561,N_436,N_1231);
nand U5562 (N_5562,N_494,N_1970);
and U5563 (N_5563,N_10,N_2965);
nand U5564 (N_5564,N_172,N_2651);
nor U5565 (N_5565,N_2249,N_2750);
nor U5566 (N_5566,N_772,N_725);
nor U5567 (N_5567,N_1732,N_996);
nand U5568 (N_5568,N_2042,N_2541);
nor U5569 (N_5569,N_2202,N_644);
and U5570 (N_5570,N_43,N_2191);
nand U5571 (N_5571,N_2939,N_1249);
nor U5572 (N_5572,N_1588,N_1958);
and U5573 (N_5573,N_2008,N_364);
nand U5574 (N_5574,N_2764,N_894);
or U5575 (N_5575,N_2097,N_163);
and U5576 (N_5576,N_313,N_802);
nor U5577 (N_5577,N_266,N_1891);
and U5578 (N_5578,N_337,N_606);
and U5579 (N_5579,N_804,N_885);
nor U5580 (N_5580,N_2127,N_2302);
or U5581 (N_5581,N_2344,N_2949);
and U5582 (N_5582,N_597,N_2178);
or U5583 (N_5583,N_949,N_1083);
nand U5584 (N_5584,N_1144,N_2326);
nor U5585 (N_5585,N_2262,N_1146);
nor U5586 (N_5586,N_1797,N_1356);
and U5587 (N_5587,N_1114,N_1171);
nor U5588 (N_5588,N_757,N_2553);
xnor U5589 (N_5589,N_2763,N_1751);
or U5590 (N_5590,N_1071,N_2889);
or U5591 (N_5591,N_2479,N_99);
nand U5592 (N_5592,N_513,N_920);
nand U5593 (N_5593,N_1854,N_1123);
nor U5594 (N_5594,N_1123,N_53);
or U5595 (N_5595,N_829,N_908);
nor U5596 (N_5596,N_2642,N_221);
and U5597 (N_5597,N_1713,N_1723);
nor U5598 (N_5598,N_1205,N_2721);
nand U5599 (N_5599,N_1458,N_945);
nor U5600 (N_5600,N_2527,N_2730);
nand U5601 (N_5601,N_2739,N_2580);
or U5602 (N_5602,N_1718,N_95);
nand U5603 (N_5603,N_253,N_250);
and U5604 (N_5604,N_1238,N_1422);
or U5605 (N_5605,N_2229,N_1837);
nor U5606 (N_5606,N_830,N_1159);
and U5607 (N_5607,N_2855,N_1688);
or U5608 (N_5608,N_2293,N_1675);
and U5609 (N_5609,N_2634,N_223);
nor U5610 (N_5610,N_1241,N_1082);
or U5611 (N_5611,N_1786,N_2623);
nor U5612 (N_5612,N_769,N_2763);
nor U5613 (N_5613,N_767,N_2258);
and U5614 (N_5614,N_924,N_348);
nand U5615 (N_5615,N_1284,N_922);
nor U5616 (N_5616,N_1902,N_72);
nand U5617 (N_5617,N_80,N_224);
nand U5618 (N_5618,N_1729,N_2759);
or U5619 (N_5619,N_2821,N_912);
nand U5620 (N_5620,N_2925,N_208);
and U5621 (N_5621,N_2874,N_2199);
nor U5622 (N_5622,N_2981,N_1755);
or U5623 (N_5623,N_2165,N_2383);
and U5624 (N_5624,N_2026,N_101);
nor U5625 (N_5625,N_259,N_1045);
and U5626 (N_5626,N_2692,N_2776);
or U5627 (N_5627,N_2608,N_1832);
and U5628 (N_5628,N_2331,N_563);
or U5629 (N_5629,N_2531,N_2492);
and U5630 (N_5630,N_116,N_2422);
and U5631 (N_5631,N_617,N_2723);
nand U5632 (N_5632,N_655,N_2450);
and U5633 (N_5633,N_895,N_1641);
or U5634 (N_5634,N_2129,N_2645);
nor U5635 (N_5635,N_2703,N_2771);
or U5636 (N_5636,N_2434,N_543);
nor U5637 (N_5637,N_1826,N_633);
nand U5638 (N_5638,N_405,N_595);
or U5639 (N_5639,N_1103,N_151);
nor U5640 (N_5640,N_2763,N_2786);
and U5641 (N_5641,N_2766,N_1854);
xnor U5642 (N_5642,N_547,N_331);
and U5643 (N_5643,N_1865,N_1785);
nand U5644 (N_5644,N_778,N_2385);
and U5645 (N_5645,N_1143,N_2394);
nand U5646 (N_5646,N_1987,N_1864);
or U5647 (N_5647,N_1076,N_2927);
nor U5648 (N_5648,N_1982,N_899);
nor U5649 (N_5649,N_7,N_1375);
nand U5650 (N_5650,N_2425,N_1473);
and U5651 (N_5651,N_2238,N_2235);
and U5652 (N_5652,N_327,N_1538);
nand U5653 (N_5653,N_591,N_999);
nor U5654 (N_5654,N_1466,N_734);
nor U5655 (N_5655,N_2775,N_1568);
nor U5656 (N_5656,N_1488,N_2247);
and U5657 (N_5657,N_509,N_620);
nand U5658 (N_5658,N_780,N_548);
or U5659 (N_5659,N_1136,N_151);
nor U5660 (N_5660,N_2327,N_2864);
xor U5661 (N_5661,N_865,N_1895);
and U5662 (N_5662,N_353,N_1353);
nand U5663 (N_5663,N_2439,N_1227);
or U5664 (N_5664,N_2246,N_2164);
nor U5665 (N_5665,N_342,N_1786);
or U5666 (N_5666,N_506,N_1286);
and U5667 (N_5667,N_1749,N_974);
nor U5668 (N_5668,N_2358,N_1824);
nor U5669 (N_5669,N_2718,N_701);
nor U5670 (N_5670,N_2538,N_127);
and U5671 (N_5671,N_232,N_1092);
nand U5672 (N_5672,N_1156,N_381);
nand U5673 (N_5673,N_2713,N_891);
nand U5674 (N_5674,N_1327,N_2603);
and U5675 (N_5675,N_1911,N_2826);
nor U5676 (N_5676,N_1952,N_52);
nor U5677 (N_5677,N_2739,N_1321);
or U5678 (N_5678,N_284,N_295);
and U5679 (N_5679,N_303,N_2853);
nor U5680 (N_5680,N_357,N_1455);
nand U5681 (N_5681,N_537,N_2533);
nand U5682 (N_5682,N_219,N_747);
nor U5683 (N_5683,N_2347,N_2114);
nand U5684 (N_5684,N_2247,N_2617);
nand U5685 (N_5685,N_1866,N_996);
nand U5686 (N_5686,N_625,N_2151);
nand U5687 (N_5687,N_1692,N_2713);
and U5688 (N_5688,N_2939,N_1980);
or U5689 (N_5689,N_531,N_2404);
or U5690 (N_5690,N_663,N_1752);
nand U5691 (N_5691,N_1157,N_170);
nand U5692 (N_5692,N_2907,N_2477);
nand U5693 (N_5693,N_741,N_2904);
nor U5694 (N_5694,N_574,N_2414);
nor U5695 (N_5695,N_2920,N_298);
or U5696 (N_5696,N_418,N_2366);
nor U5697 (N_5697,N_445,N_1951);
and U5698 (N_5698,N_2297,N_1046);
nand U5699 (N_5699,N_1915,N_1545);
nor U5700 (N_5700,N_2939,N_1858);
nand U5701 (N_5701,N_2937,N_1310);
nor U5702 (N_5702,N_2742,N_2124);
nand U5703 (N_5703,N_1314,N_612);
nor U5704 (N_5704,N_2033,N_2505);
nand U5705 (N_5705,N_49,N_1967);
or U5706 (N_5706,N_113,N_2580);
and U5707 (N_5707,N_2473,N_1038);
or U5708 (N_5708,N_2631,N_2276);
and U5709 (N_5709,N_2749,N_1275);
nand U5710 (N_5710,N_2204,N_833);
and U5711 (N_5711,N_1284,N_1619);
or U5712 (N_5712,N_669,N_2490);
or U5713 (N_5713,N_2753,N_517);
nor U5714 (N_5714,N_1272,N_367);
and U5715 (N_5715,N_368,N_2393);
or U5716 (N_5716,N_884,N_312);
nor U5717 (N_5717,N_1288,N_486);
and U5718 (N_5718,N_1791,N_1356);
nor U5719 (N_5719,N_1085,N_1978);
nand U5720 (N_5720,N_155,N_1568);
nor U5721 (N_5721,N_722,N_1298);
or U5722 (N_5722,N_49,N_1674);
or U5723 (N_5723,N_2135,N_2561);
or U5724 (N_5724,N_1193,N_799);
nor U5725 (N_5725,N_2638,N_683);
nand U5726 (N_5726,N_292,N_739);
nand U5727 (N_5727,N_1443,N_841);
nor U5728 (N_5728,N_1702,N_879);
nor U5729 (N_5729,N_2615,N_1234);
and U5730 (N_5730,N_202,N_1228);
and U5731 (N_5731,N_2568,N_271);
nor U5732 (N_5732,N_2748,N_2654);
nor U5733 (N_5733,N_2747,N_631);
xnor U5734 (N_5734,N_1193,N_203);
or U5735 (N_5735,N_1917,N_250);
and U5736 (N_5736,N_1113,N_1424);
nor U5737 (N_5737,N_996,N_2129);
or U5738 (N_5738,N_1380,N_1593);
or U5739 (N_5739,N_1998,N_1174);
nand U5740 (N_5740,N_1543,N_1479);
nand U5741 (N_5741,N_258,N_70);
and U5742 (N_5742,N_2096,N_905);
or U5743 (N_5743,N_701,N_382);
or U5744 (N_5744,N_1645,N_1614);
and U5745 (N_5745,N_1258,N_539);
or U5746 (N_5746,N_1030,N_833);
and U5747 (N_5747,N_1939,N_2524);
nand U5748 (N_5748,N_985,N_1693);
and U5749 (N_5749,N_2533,N_1962);
or U5750 (N_5750,N_2582,N_2822);
and U5751 (N_5751,N_2623,N_2541);
nor U5752 (N_5752,N_2455,N_53);
nor U5753 (N_5753,N_2544,N_2589);
nor U5754 (N_5754,N_54,N_1217);
or U5755 (N_5755,N_2259,N_1357);
nor U5756 (N_5756,N_2025,N_2752);
nand U5757 (N_5757,N_2663,N_2288);
nor U5758 (N_5758,N_2035,N_2976);
nor U5759 (N_5759,N_606,N_2200);
nor U5760 (N_5760,N_2077,N_682);
or U5761 (N_5761,N_654,N_2774);
nor U5762 (N_5762,N_2768,N_1767);
nand U5763 (N_5763,N_0,N_1082);
nor U5764 (N_5764,N_1083,N_398);
nand U5765 (N_5765,N_422,N_557);
nor U5766 (N_5766,N_2629,N_1611);
or U5767 (N_5767,N_2879,N_1127);
nand U5768 (N_5768,N_1070,N_2409);
nor U5769 (N_5769,N_333,N_2663);
nor U5770 (N_5770,N_687,N_2603);
and U5771 (N_5771,N_1515,N_79);
nand U5772 (N_5772,N_2889,N_1816);
and U5773 (N_5773,N_1807,N_1660);
nand U5774 (N_5774,N_1871,N_1975);
nor U5775 (N_5775,N_852,N_993);
or U5776 (N_5776,N_2241,N_188);
and U5777 (N_5777,N_2457,N_2803);
nand U5778 (N_5778,N_1523,N_1222);
nand U5779 (N_5779,N_650,N_332);
and U5780 (N_5780,N_719,N_620);
xor U5781 (N_5781,N_2697,N_389);
nand U5782 (N_5782,N_1116,N_747);
or U5783 (N_5783,N_1148,N_1177);
nor U5784 (N_5784,N_2032,N_1996);
nor U5785 (N_5785,N_919,N_885);
nor U5786 (N_5786,N_2755,N_253);
and U5787 (N_5787,N_1563,N_1343);
and U5788 (N_5788,N_1034,N_2684);
and U5789 (N_5789,N_2672,N_694);
nand U5790 (N_5790,N_376,N_1261);
nor U5791 (N_5791,N_2232,N_720);
or U5792 (N_5792,N_1573,N_1016);
nand U5793 (N_5793,N_2090,N_2834);
nor U5794 (N_5794,N_1737,N_1333);
nand U5795 (N_5795,N_2920,N_975);
or U5796 (N_5796,N_261,N_1308);
nand U5797 (N_5797,N_2594,N_2619);
nand U5798 (N_5798,N_2301,N_2519);
or U5799 (N_5799,N_2647,N_2184);
nor U5800 (N_5800,N_6,N_1835);
or U5801 (N_5801,N_1002,N_418);
or U5802 (N_5802,N_1660,N_472);
or U5803 (N_5803,N_2918,N_2410);
nor U5804 (N_5804,N_2982,N_2375);
xnor U5805 (N_5805,N_1739,N_1246);
and U5806 (N_5806,N_889,N_1992);
nand U5807 (N_5807,N_1246,N_2769);
nor U5808 (N_5808,N_1966,N_213);
and U5809 (N_5809,N_1914,N_178);
or U5810 (N_5810,N_2014,N_1537);
nand U5811 (N_5811,N_645,N_1015);
and U5812 (N_5812,N_2312,N_2251);
or U5813 (N_5813,N_2518,N_1573);
and U5814 (N_5814,N_615,N_1225);
nand U5815 (N_5815,N_849,N_639);
or U5816 (N_5816,N_2246,N_249);
or U5817 (N_5817,N_170,N_1896);
nand U5818 (N_5818,N_734,N_2350);
and U5819 (N_5819,N_2105,N_2485);
nor U5820 (N_5820,N_2828,N_1217);
or U5821 (N_5821,N_801,N_380);
nor U5822 (N_5822,N_2983,N_1304);
or U5823 (N_5823,N_1466,N_1234);
nor U5824 (N_5824,N_1475,N_608);
nor U5825 (N_5825,N_330,N_2779);
and U5826 (N_5826,N_2384,N_1006);
or U5827 (N_5827,N_2756,N_57);
and U5828 (N_5828,N_2264,N_2285);
and U5829 (N_5829,N_1418,N_1339);
and U5830 (N_5830,N_394,N_1633);
or U5831 (N_5831,N_2843,N_1139);
nand U5832 (N_5832,N_732,N_1944);
or U5833 (N_5833,N_2573,N_1390);
nor U5834 (N_5834,N_2558,N_1914);
nand U5835 (N_5835,N_519,N_2007);
nor U5836 (N_5836,N_1456,N_2121);
and U5837 (N_5837,N_1404,N_418);
nand U5838 (N_5838,N_1133,N_130);
and U5839 (N_5839,N_55,N_2546);
nor U5840 (N_5840,N_2465,N_1409);
and U5841 (N_5841,N_2691,N_908);
or U5842 (N_5842,N_1374,N_2827);
or U5843 (N_5843,N_1070,N_397);
nor U5844 (N_5844,N_278,N_1312);
and U5845 (N_5845,N_2080,N_2899);
or U5846 (N_5846,N_1917,N_1680);
or U5847 (N_5847,N_1253,N_1892);
and U5848 (N_5848,N_2362,N_548);
nand U5849 (N_5849,N_2887,N_406);
and U5850 (N_5850,N_209,N_1318);
nor U5851 (N_5851,N_111,N_2422);
or U5852 (N_5852,N_1563,N_482);
nor U5853 (N_5853,N_2729,N_559);
xor U5854 (N_5854,N_1203,N_1134);
nor U5855 (N_5855,N_347,N_1534);
nand U5856 (N_5856,N_64,N_1113);
or U5857 (N_5857,N_2984,N_994);
or U5858 (N_5858,N_2788,N_1273);
or U5859 (N_5859,N_1691,N_1512);
and U5860 (N_5860,N_357,N_735);
nand U5861 (N_5861,N_940,N_2533);
and U5862 (N_5862,N_369,N_148);
or U5863 (N_5863,N_157,N_1904);
and U5864 (N_5864,N_885,N_2613);
nor U5865 (N_5865,N_1228,N_2816);
nor U5866 (N_5866,N_2845,N_2084);
nand U5867 (N_5867,N_1337,N_536);
and U5868 (N_5868,N_2756,N_2607);
nand U5869 (N_5869,N_2603,N_403);
nor U5870 (N_5870,N_2467,N_987);
or U5871 (N_5871,N_471,N_2437);
or U5872 (N_5872,N_117,N_313);
or U5873 (N_5873,N_2642,N_2169);
nand U5874 (N_5874,N_1190,N_142);
or U5875 (N_5875,N_2823,N_2991);
and U5876 (N_5876,N_2025,N_1516);
or U5877 (N_5877,N_1522,N_1249);
or U5878 (N_5878,N_1597,N_2743);
nor U5879 (N_5879,N_1432,N_1921);
and U5880 (N_5880,N_2263,N_998);
nor U5881 (N_5881,N_996,N_1150);
nand U5882 (N_5882,N_2985,N_1320);
nor U5883 (N_5883,N_152,N_1751);
or U5884 (N_5884,N_1417,N_1001);
nor U5885 (N_5885,N_1687,N_1317);
nor U5886 (N_5886,N_1846,N_1691);
nand U5887 (N_5887,N_1548,N_617);
nor U5888 (N_5888,N_282,N_2323);
and U5889 (N_5889,N_290,N_863);
nor U5890 (N_5890,N_1609,N_1044);
nand U5891 (N_5891,N_1592,N_914);
nand U5892 (N_5892,N_2092,N_2061);
nor U5893 (N_5893,N_630,N_1178);
nor U5894 (N_5894,N_2523,N_1535);
nand U5895 (N_5895,N_136,N_2139);
or U5896 (N_5896,N_930,N_2044);
nor U5897 (N_5897,N_2904,N_2137);
nand U5898 (N_5898,N_2731,N_667);
nor U5899 (N_5899,N_212,N_1852);
and U5900 (N_5900,N_505,N_2203);
nor U5901 (N_5901,N_1338,N_1180);
and U5902 (N_5902,N_2160,N_2023);
nand U5903 (N_5903,N_1520,N_2277);
nand U5904 (N_5904,N_2848,N_483);
nand U5905 (N_5905,N_2548,N_2131);
or U5906 (N_5906,N_1941,N_2235);
nand U5907 (N_5907,N_1209,N_2094);
or U5908 (N_5908,N_1670,N_2391);
and U5909 (N_5909,N_2621,N_1352);
and U5910 (N_5910,N_205,N_881);
and U5911 (N_5911,N_1029,N_2776);
or U5912 (N_5912,N_150,N_2913);
nor U5913 (N_5913,N_629,N_316);
and U5914 (N_5914,N_2647,N_437);
nand U5915 (N_5915,N_1287,N_2028);
nand U5916 (N_5916,N_1114,N_1061);
and U5917 (N_5917,N_1309,N_2625);
nor U5918 (N_5918,N_2665,N_596);
nand U5919 (N_5919,N_2099,N_1341);
nand U5920 (N_5920,N_702,N_2657);
or U5921 (N_5921,N_231,N_592);
nor U5922 (N_5922,N_698,N_2416);
or U5923 (N_5923,N_1356,N_1116);
or U5924 (N_5924,N_577,N_1382);
nor U5925 (N_5925,N_2563,N_174);
nor U5926 (N_5926,N_2689,N_960);
nor U5927 (N_5927,N_2865,N_2035);
or U5928 (N_5928,N_537,N_1887);
nor U5929 (N_5929,N_1252,N_2638);
nor U5930 (N_5930,N_316,N_2871);
and U5931 (N_5931,N_742,N_806);
nand U5932 (N_5932,N_1485,N_1594);
or U5933 (N_5933,N_2944,N_2294);
and U5934 (N_5934,N_906,N_2184);
nand U5935 (N_5935,N_2479,N_911);
or U5936 (N_5936,N_351,N_1172);
nor U5937 (N_5937,N_416,N_2325);
and U5938 (N_5938,N_1058,N_956);
and U5939 (N_5939,N_1950,N_341);
or U5940 (N_5940,N_1180,N_2593);
nand U5941 (N_5941,N_342,N_1052);
nor U5942 (N_5942,N_2274,N_1469);
and U5943 (N_5943,N_1215,N_2600);
or U5944 (N_5944,N_1401,N_2988);
or U5945 (N_5945,N_2573,N_905);
xnor U5946 (N_5946,N_1105,N_1065);
and U5947 (N_5947,N_1171,N_1750);
and U5948 (N_5948,N_2278,N_2478);
or U5949 (N_5949,N_2975,N_1248);
and U5950 (N_5950,N_1574,N_189);
nor U5951 (N_5951,N_1538,N_489);
nand U5952 (N_5952,N_1210,N_2115);
nand U5953 (N_5953,N_119,N_1293);
and U5954 (N_5954,N_157,N_387);
nor U5955 (N_5955,N_668,N_661);
or U5956 (N_5956,N_518,N_335);
nand U5957 (N_5957,N_2869,N_2973);
nand U5958 (N_5958,N_1983,N_2730);
nand U5959 (N_5959,N_380,N_2909);
nor U5960 (N_5960,N_2086,N_1599);
or U5961 (N_5961,N_649,N_464);
nand U5962 (N_5962,N_1096,N_731);
and U5963 (N_5963,N_770,N_1270);
nand U5964 (N_5964,N_2702,N_2628);
nor U5965 (N_5965,N_937,N_498);
or U5966 (N_5966,N_657,N_2264);
nor U5967 (N_5967,N_49,N_609);
nor U5968 (N_5968,N_2955,N_2185);
nor U5969 (N_5969,N_2634,N_444);
nand U5970 (N_5970,N_1659,N_1669);
nor U5971 (N_5971,N_2237,N_1463);
and U5972 (N_5972,N_2210,N_106);
nand U5973 (N_5973,N_240,N_1157);
nand U5974 (N_5974,N_2882,N_556);
nand U5975 (N_5975,N_1687,N_1700);
nor U5976 (N_5976,N_980,N_919);
or U5977 (N_5977,N_83,N_1349);
and U5978 (N_5978,N_686,N_320);
nor U5979 (N_5979,N_53,N_1700);
or U5980 (N_5980,N_1190,N_1516);
nor U5981 (N_5981,N_1052,N_337);
xnor U5982 (N_5982,N_1772,N_2624);
or U5983 (N_5983,N_2642,N_2029);
and U5984 (N_5984,N_2719,N_122);
nor U5985 (N_5985,N_2185,N_39);
or U5986 (N_5986,N_1395,N_2477);
nor U5987 (N_5987,N_1125,N_86);
nor U5988 (N_5988,N_2558,N_2323);
or U5989 (N_5989,N_2814,N_1288);
and U5990 (N_5990,N_59,N_1372);
xor U5991 (N_5991,N_2296,N_2538);
or U5992 (N_5992,N_366,N_2550);
and U5993 (N_5993,N_1036,N_1945);
or U5994 (N_5994,N_2535,N_127);
and U5995 (N_5995,N_2570,N_2803);
nand U5996 (N_5996,N_734,N_1869);
or U5997 (N_5997,N_1252,N_543);
and U5998 (N_5998,N_2621,N_472);
nor U5999 (N_5999,N_881,N_1683);
nor U6000 (N_6000,N_4135,N_5414);
and U6001 (N_6001,N_5326,N_3749);
nand U6002 (N_6002,N_4612,N_4207);
or U6003 (N_6003,N_3972,N_5155);
nor U6004 (N_6004,N_5954,N_4358);
nand U6005 (N_6005,N_5944,N_4393);
and U6006 (N_6006,N_5718,N_4403);
nand U6007 (N_6007,N_4430,N_5128);
nor U6008 (N_6008,N_5329,N_3504);
nand U6009 (N_6009,N_3337,N_5118);
nor U6010 (N_6010,N_4708,N_4072);
and U6011 (N_6011,N_3732,N_4411);
nand U6012 (N_6012,N_3718,N_5038);
or U6013 (N_6013,N_5767,N_4660);
or U6014 (N_6014,N_5911,N_5417);
or U6015 (N_6015,N_5806,N_4920);
nand U6016 (N_6016,N_5217,N_5487);
or U6017 (N_6017,N_3459,N_5597);
nand U6018 (N_6018,N_5776,N_4374);
and U6019 (N_6019,N_5212,N_5664);
xnor U6020 (N_6020,N_3555,N_5448);
and U6021 (N_6021,N_5822,N_5109);
or U6022 (N_6022,N_3675,N_5532);
nor U6023 (N_6023,N_4657,N_3082);
or U6024 (N_6024,N_4617,N_3456);
and U6025 (N_6025,N_5492,N_5385);
and U6026 (N_6026,N_5669,N_4241);
and U6027 (N_6027,N_4132,N_5022);
or U6028 (N_6028,N_5769,N_4850);
or U6029 (N_6029,N_4454,N_4165);
nand U6030 (N_6030,N_5552,N_4450);
and U6031 (N_6031,N_4714,N_4339);
nand U6032 (N_6032,N_3104,N_5710);
or U6033 (N_6033,N_3697,N_3430);
and U6034 (N_6034,N_4995,N_3823);
and U6035 (N_6035,N_3349,N_3310);
and U6036 (N_6036,N_3470,N_3515);
and U6037 (N_6037,N_4844,N_3371);
xnor U6038 (N_6038,N_3530,N_3256);
nand U6039 (N_6039,N_5379,N_4967);
or U6040 (N_6040,N_4020,N_5571);
and U6041 (N_6041,N_5538,N_4666);
xnor U6042 (N_6042,N_4401,N_5603);
and U6043 (N_6043,N_3519,N_5953);
or U6044 (N_6044,N_5051,N_5026);
nor U6045 (N_6045,N_5549,N_3672);
nand U6046 (N_6046,N_4774,N_4114);
or U6047 (N_6047,N_3626,N_3221);
or U6048 (N_6048,N_4410,N_3159);
and U6049 (N_6049,N_5488,N_4476);
nand U6050 (N_6050,N_5061,N_4895);
and U6051 (N_6051,N_4100,N_4286);
and U6052 (N_6052,N_4890,N_3360);
and U6053 (N_6053,N_3854,N_5279);
nand U6054 (N_6054,N_4434,N_3200);
and U6055 (N_6055,N_4574,N_5010);
or U6056 (N_6056,N_3034,N_5519);
or U6057 (N_6057,N_3063,N_4356);
or U6058 (N_6058,N_5435,N_4394);
and U6059 (N_6059,N_3368,N_3378);
or U6060 (N_6060,N_5274,N_4716);
nand U6061 (N_6061,N_4999,N_3801);
and U6062 (N_6062,N_4550,N_4070);
nor U6063 (N_6063,N_5447,N_5007);
or U6064 (N_6064,N_5221,N_5736);
and U6065 (N_6065,N_5638,N_3413);
or U6066 (N_6066,N_3653,N_5497);
and U6067 (N_6067,N_3988,N_3856);
xor U6068 (N_6068,N_5514,N_4876);
or U6069 (N_6069,N_3589,N_5608);
and U6070 (N_6070,N_5582,N_5804);
nand U6071 (N_6071,N_3648,N_4795);
and U6072 (N_6072,N_5885,N_4773);
nor U6073 (N_6073,N_5614,N_4889);
nor U6074 (N_6074,N_3240,N_3217);
or U6075 (N_6075,N_3879,N_5180);
nor U6076 (N_6076,N_4663,N_4470);
and U6077 (N_6077,N_4661,N_5122);
and U6078 (N_6078,N_4233,N_5153);
nand U6079 (N_6079,N_5306,N_5512);
nand U6080 (N_6080,N_4246,N_3620);
nor U6081 (N_6081,N_3521,N_4051);
nand U6082 (N_6082,N_3486,N_5275);
or U6083 (N_6083,N_4524,N_5255);
nand U6084 (N_6084,N_5339,N_4271);
nor U6085 (N_6085,N_3436,N_5420);
nor U6086 (N_6086,N_4564,N_5360);
or U6087 (N_6087,N_5357,N_5528);
or U6088 (N_6088,N_3405,N_3911);
nand U6089 (N_6089,N_5244,N_5292);
nor U6090 (N_6090,N_5475,N_3334);
and U6091 (N_6091,N_3354,N_5042);
or U6092 (N_6092,N_3272,N_5593);
and U6093 (N_6093,N_3674,N_5886);
and U6094 (N_6094,N_3095,N_5152);
nand U6095 (N_6095,N_5317,N_4636);
or U6096 (N_6096,N_5300,N_4749);
and U6097 (N_6097,N_5063,N_3579);
and U6098 (N_6098,N_5267,N_5580);
nand U6099 (N_6099,N_3422,N_4928);
and U6100 (N_6100,N_4047,N_3918);
nand U6101 (N_6101,N_5008,N_4518);
or U6102 (N_6102,N_4644,N_3618);
and U6103 (N_6103,N_3925,N_4382);
xor U6104 (N_6104,N_4802,N_3587);
or U6105 (N_6105,N_3943,N_5733);
nand U6106 (N_6106,N_5330,N_3287);
nor U6107 (N_6107,N_3543,N_3263);
nor U6108 (N_6108,N_4916,N_4863);
xnor U6109 (N_6109,N_3971,N_3940);
and U6110 (N_6110,N_4109,N_3963);
or U6111 (N_6111,N_4436,N_3094);
or U6112 (N_6112,N_4162,N_5559);
nor U6113 (N_6113,N_5199,N_5511);
nor U6114 (N_6114,N_4260,N_5649);
and U6115 (N_6115,N_4579,N_4231);
xnor U6116 (N_6116,N_3317,N_4329);
nand U6117 (N_6117,N_3609,N_4192);
nand U6118 (N_6118,N_3717,N_5974);
nor U6119 (N_6119,N_4061,N_3212);
nor U6120 (N_6120,N_3731,N_3125);
and U6121 (N_6121,N_5728,N_5505);
or U6122 (N_6122,N_3264,N_5772);
nor U6123 (N_6123,N_3214,N_4658);
nor U6124 (N_6124,N_5095,N_4723);
or U6125 (N_6125,N_5749,N_4623);
and U6126 (N_6126,N_4408,N_3556);
and U6127 (N_6127,N_3818,N_4487);
nand U6128 (N_6128,N_5369,N_4944);
and U6129 (N_6129,N_3130,N_3072);
and U6130 (N_6130,N_4614,N_3280);
nor U6131 (N_6131,N_3944,N_4053);
or U6132 (N_6132,N_4010,N_3733);
and U6133 (N_6133,N_3143,N_3399);
and U6134 (N_6134,N_3931,N_4908);
or U6135 (N_6135,N_4050,N_5590);
or U6136 (N_6136,N_3651,N_5864);
nand U6137 (N_6137,N_5151,N_4502);
and U6138 (N_6138,N_4370,N_5518);
nand U6139 (N_6139,N_4855,N_4040);
xor U6140 (N_6140,N_5302,N_3137);
or U6141 (N_6141,N_3656,N_5003);
and U6142 (N_6142,N_4551,N_5052);
nand U6143 (N_6143,N_3475,N_4979);
or U6144 (N_6144,N_4297,N_4957);
and U6145 (N_6145,N_3296,N_4811);
nor U6146 (N_6146,N_4156,N_4019);
nor U6147 (N_6147,N_5851,N_3951);
and U6148 (N_6148,N_5522,N_3313);
or U6149 (N_6149,N_4864,N_4990);
nand U6150 (N_6150,N_3324,N_3301);
or U6151 (N_6151,N_4289,N_4484);
nand U6152 (N_6152,N_5237,N_5539);
nor U6153 (N_6153,N_5135,N_3690);
or U6154 (N_6154,N_3339,N_4672);
nand U6155 (N_6155,N_5945,N_4390);
nand U6156 (N_6156,N_3336,N_5923);
nor U6157 (N_6157,N_3984,N_5148);
or U6158 (N_6158,N_5111,N_5101);
or U6159 (N_6159,N_5353,N_4664);
and U6160 (N_6160,N_5730,N_3631);
nand U6161 (N_6161,N_4234,N_3634);
or U6162 (N_6162,N_3919,N_3231);
or U6163 (N_6163,N_5999,N_4939);
or U6164 (N_6164,N_3204,N_5948);
and U6165 (N_6165,N_3734,N_4413);
or U6166 (N_6166,N_4177,N_4331);
or U6167 (N_6167,N_3945,N_4712);
or U6168 (N_6168,N_5783,N_5691);
nand U6169 (N_6169,N_3490,N_3489);
or U6170 (N_6170,N_4938,N_3719);
xor U6171 (N_6171,N_3291,N_4062);
nor U6172 (N_6172,N_4333,N_3821);
or U6173 (N_6173,N_5693,N_5560);
or U6174 (N_6174,N_4093,N_3670);
nor U6175 (N_6175,N_3380,N_5645);
nor U6176 (N_6176,N_3414,N_3182);
nand U6177 (N_6177,N_5651,N_3767);
and U6178 (N_6178,N_5181,N_4540);
or U6179 (N_6179,N_4589,N_4490);
nand U6180 (N_6180,N_4302,N_5219);
nand U6181 (N_6181,N_4075,N_5112);
nand U6182 (N_6182,N_5790,N_4818);
or U6183 (N_6183,N_5106,N_4198);
or U6184 (N_6184,N_5717,N_3786);
nor U6185 (N_6185,N_4480,N_3529);
nand U6186 (N_6186,N_5335,N_3882);
nand U6187 (N_6187,N_5070,N_4477);
nand U6188 (N_6188,N_3056,N_5110);
nor U6189 (N_6189,N_4178,N_5609);
nand U6190 (N_6190,N_5928,N_3228);
and U6191 (N_6191,N_5156,N_5228);
or U6192 (N_6192,N_4236,N_5652);
nor U6193 (N_6193,N_4710,N_4251);
nor U6194 (N_6194,N_4378,N_5982);
and U6195 (N_6195,N_5470,N_3260);
nand U6196 (N_6196,N_3139,N_3596);
nor U6197 (N_6197,N_5039,N_3561);
and U6198 (N_6198,N_5424,N_5879);
and U6199 (N_6199,N_4486,N_4686);
xor U6200 (N_6200,N_5281,N_5458);
nor U6201 (N_6201,N_4639,N_4254);
or U6202 (N_6202,N_4046,N_4185);
and U6203 (N_6203,N_5338,N_4910);
nor U6204 (N_6204,N_4744,N_5639);
nand U6205 (N_6205,N_3538,N_3491);
and U6206 (N_6206,N_5348,N_3169);
or U6207 (N_6207,N_4580,N_3744);
nor U6208 (N_6208,N_4201,N_4513);
or U6209 (N_6209,N_4959,N_4348);
or U6210 (N_6210,N_3271,N_5239);
or U6211 (N_6211,N_3016,N_4536);
or U6212 (N_6212,N_5214,N_4497);
and U6213 (N_6213,N_5410,N_4258);
or U6214 (N_6214,N_4735,N_3031);
nor U6215 (N_6215,N_3300,N_5293);
nor U6216 (N_6216,N_3533,N_5189);
nor U6217 (N_6217,N_3111,N_3659);
nand U6218 (N_6218,N_4154,N_3708);
and U6219 (N_6219,N_4845,N_3539);
and U6220 (N_6220,N_3472,N_3764);
nand U6221 (N_6221,N_3974,N_3434);
xnor U6222 (N_6222,N_4711,N_3702);
or U6223 (N_6223,N_3583,N_5149);
or U6224 (N_6224,N_3637,N_5397);
and U6225 (N_6225,N_5299,N_4142);
or U6226 (N_6226,N_3868,N_4960);
nand U6227 (N_6227,N_5079,N_3040);
and U6228 (N_6228,N_4553,N_3006);
or U6229 (N_6229,N_4103,N_3549);
nor U6230 (N_6230,N_3437,N_3950);
and U6231 (N_6231,N_5831,N_4973);
nor U6232 (N_6232,N_4618,N_4298);
or U6233 (N_6233,N_4772,N_4210);
and U6234 (N_6234,N_5671,N_3014);
nand U6235 (N_6235,N_3728,N_5235);
nand U6236 (N_6236,N_4029,N_3048);
or U6237 (N_6237,N_4698,N_3450);
and U6238 (N_6238,N_4321,N_5890);
and U6239 (N_6239,N_3921,N_3975);
or U6240 (N_6240,N_3989,N_5898);
or U6241 (N_6241,N_5754,N_3585);
nor U6242 (N_6242,N_3018,N_4404);
nor U6243 (N_6243,N_3180,N_3067);
and U6244 (N_6244,N_5677,N_5133);
nor U6245 (N_6245,N_3630,N_4343);
or U6246 (N_6246,N_3799,N_3148);
nand U6247 (N_6247,N_3790,N_5753);
nor U6248 (N_6248,N_5167,N_5014);
nand U6249 (N_6249,N_3232,N_4069);
nand U6250 (N_6250,N_3327,N_5025);
nand U6251 (N_6251,N_5252,N_3484);
nand U6252 (N_6252,N_4533,N_3815);
and U6253 (N_6253,N_5980,N_5527);
nand U6254 (N_6254,N_5506,N_3129);
nand U6255 (N_6255,N_4126,N_5197);
or U6256 (N_6256,N_4566,N_5610);
xor U6257 (N_6257,N_4906,N_3848);
or U6258 (N_6258,N_3900,N_3723);
or U6259 (N_6259,N_4738,N_5752);
or U6260 (N_6260,N_4351,N_5304);
or U6261 (N_6261,N_4164,N_4439);
and U6262 (N_6262,N_4734,N_3106);
nor U6263 (N_6263,N_5035,N_4037);
and U6264 (N_6264,N_3429,N_3443);
or U6265 (N_6265,N_5673,N_5144);
nand U6266 (N_6266,N_4598,N_4720);
and U6267 (N_6267,N_4904,N_5637);
and U6268 (N_6268,N_5810,N_4615);
nand U6269 (N_6269,N_3069,N_3101);
xnor U6270 (N_6270,N_5823,N_5942);
or U6271 (N_6271,N_3866,N_5108);
or U6272 (N_6272,N_5588,N_5005);
or U6273 (N_6273,N_3132,N_3622);
nand U6274 (N_6274,N_5927,N_4252);
and U6275 (N_6275,N_4030,N_4542);
or U6276 (N_6276,N_5602,N_3604);
nand U6277 (N_6277,N_4721,N_3927);
nand U6278 (N_6278,N_5346,N_4512);
xnor U6279 (N_6279,N_3865,N_3615);
or U6280 (N_6280,N_3320,N_3477);
or U6281 (N_6281,N_5596,N_3178);
nor U6282 (N_6282,N_3760,N_4226);
or U6283 (N_6283,N_5843,N_3568);
nor U6284 (N_6284,N_4974,N_5784);
nand U6285 (N_6285,N_3128,N_5740);
nand U6286 (N_6286,N_4823,N_3559);
or U6287 (N_6287,N_3558,N_5365);
nor U6288 (N_6288,N_5315,N_3294);
nor U6289 (N_6289,N_5502,N_3857);
nor U6290 (N_6290,N_4642,N_3557);
or U6291 (N_6291,N_4651,N_5091);
nand U6292 (N_6292,N_4785,N_5553);
nor U6293 (N_6293,N_4678,N_5382);
or U6294 (N_6294,N_3150,N_4459);
or U6295 (N_6295,N_5012,N_4364);
xor U6296 (N_6296,N_4911,N_4527);
or U6297 (N_6297,N_4360,N_3121);
or U6298 (N_6298,N_5263,N_3058);
nor U6299 (N_6299,N_5159,N_4143);
nand U6300 (N_6300,N_3782,N_4288);
nor U6301 (N_6301,N_5479,N_4872);
or U6302 (N_6302,N_5732,N_3729);
and U6303 (N_6303,N_3142,N_5918);
nor U6304 (N_6304,N_4846,N_4954);
or U6305 (N_6305,N_3374,N_4746);
and U6306 (N_6306,N_3677,N_3224);
nor U6307 (N_6307,N_3134,N_4966);
nor U6308 (N_6308,N_4753,N_5179);
nand U6309 (N_6309,N_5828,N_3164);
nand U6310 (N_6310,N_3157,N_4627);
nand U6311 (N_6311,N_4853,N_5543);
and U6312 (N_6312,N_4211,N_5647);
and U6313 (N_6313,N_3353,N_4577);
or U6314 (N_6314,N_5940,N_5257);
nand U6315 (N_6315,N_5320,N_5866);
and U6316 (N_6316,N_4758,N_5876);
and U6317 (N_6317,N_4670,N_3955);
or U6318 (N_6318,N_5620,N_3898);
nor U6319 (N_6319,N_3662,N_4932);
nor U6320 (N_6320,N_3131,N_3278);
and U6321 (N_6321,N_4743,N_5727);
and U6322 (N_6322,N_4862,N_4150);
and U6323 (N_6323,N_5625,N_4923);
nand U6324 (N_6324,N_5373,N_4385);
or U6325 (N_6325,N_4510,N_3474);
and U6326 (N_6326,N_5973,N_4389);
nand U6327 (N_6327,N_5950,N_4941);
nor U6328 (N_6328,N_4452,N_4015);
or U6329 (N_6329,N_3079,N_3175);
or U6330 (N_6330,N_3304,N_4197);
and U6331 (N_6331,N_4174,N_4665);
nor U6332 (N_6332,N_3766,N_4056);
and U6333 (N_6333,N_4812,N_4461);
nand U6334 (N_6334,N_4294,N_3994);
and U6335 (N_6335,N_4986,N_5642);
nor U6336 (N_6336,N_3810,N_4320);
nor U6337 (N_6337,N_4687,N_4697);
and U6338 (N_6338,N_3065,N_4695);
nand U6339 (N_6339,N_3481,N_5062);
and U6340 (N_6340,N_5814,N_4115);
nand U6341 (N_6341,N_5707,N_4208);
or U6342 (N_6342,N_3889,N_5644);
xnor U6343 (N_6343,N_4996,N_4309);
nand U6344 (N_6344,N_5738,N_3505);
nand U6345 (N_6345,N_4306,N_5551);
nand U6346 (N_6346,N_3545,N_5611);
and U6347 (N_6347,N_4544,N_5816);
xnor U6348 (N_6348,N_3683,N_5870);
nand U6349 (N_6349,N_4755,N_4763);
and U6350 (N_6350,N_3638,N_5943);
or U6351 (N_6351,N_3852,N_5524);
nor U6352 (N_6352,N_5194,N_3303);
nand U6353 (N_6353,N_3840,N_4031);
or U6354 (N_6354,N_4146,N_4530);
and U6355 (N_6355,N_4914,N_3597);
or U6356 (N_6356,N_4278,N_4138);
or U6357 (N_6357,N_3384,N_3306);
and U6358 (N_6358,N_4692,N_4464);
or U6359 (N_6359,N_4969,N_3356);
and U6360 (N_6360,N_3483,N_4011);
and U6361 (N_6361,N_4677,N_4303);
nor U6362 (N_6362,N_5993,N_5462);
and U6363 (N_6363,N_4407,N_4794);
and U6364 (N_6364,N_4905,N_3883);
or U6365 (N_6365,N_5697,N_4781);
or U6366 (N_6366,N_5599,N_5795);
or U6367 (N_6367,N_5905,N_3293);
and U6368 (N_6368,N_5557,N_4770);
nor U6369 (N_6369,N_3133,N_5157);
and U6370 (N_6370,N_5023,N_4901);
nor U6371 (N_6371,N_4313,N_5705);
and U6372 (N_6372,N_5834,N_3107);
and U6373 (N_6373,N_4330,N_3100);
nand U6374 (N_6374,N_5457,N_4406);
nand U6375 (N_6375,N_4593,N_5634);
nand U6376 (N_6376,N_4520,N_3447);
or U6377 (N_6377,N_3551,N_4222);
or U6378 (N_6378,N_3794,N_5238);
xor U6379 (N_6379,N_4237,N_4261);
nand U6380 (N_6380,N_5480,N_3938);
nor U6381 (N_6381,N_4843,N_5242);
and U6382 (N_6382,N_5248,N_4507);
nor U6383 (N_6383,N_3657,N_4526);
or U6384 (N_6384,N_4423,N_3248);
nand U6385 (N_6385,N_3935,N_4819);
or U6386 (N_6386,N_4806,N_4937);
nor U6387 (N_6387,N_4022,N_3661);
and U6388 (N_6388,N_4879,N_5979);
nand U6389 (N_6389,N_5461,N_4491);
nor U6390 (N_6390,N_3404,N_3331);
nand U6391 (N_6391,N_3689,N_4334);
and U6392 (N_6392,N_4683,N_4556);
nand U6393 (N_6393,N_4722,N_3563);
or U6394 (N_6394,N_4097,N_4894);
nor U6395 (N_6395,N_3052,N_5631);
or U6396 (N_6396,N_4568,N_5124);
nor U6397 (N_6397,N_5465,N_3881);
or U6398 (N_6398,N_4948,N_3508);
nand U6399 (N_6399,N_5399,N_3791);
nand U6400 (N_6400,N_4765,N_4805);
nor U6401 (N_6401,N_3276,N_5800);
nor U6402 (N_6402,N_3088,N_5037);
nor U6403 (N_6403,N_5321,N_3588);
nor U6404 (N_6404,N_4212,N_5722);
nand U6405 (N_6405,N_4545,N_4747);
and U6406 (N_6406,N_3873,N_4104);
and U6407 (N_6407,N_5449,N_5425);
nor U6408 (N_6408,N_4506,N_3814);
nor U6409 (N_6409,N_5706,N_4444);
nand U6410 (N_6410,N_3230,N_5380);
nand U6411 (N_6411,N_5550,N_3887);
nor U6412 (N_6412,N_5680,N_5836);
or U6413 (N_6413,N_4638,N_4004);
nor U6414 (N_6414,N_3893,N_5997);
and U6415 (N_6415,N_3019,N_3314);
nand U6416 (N_6416,N_4715,N_3438);
nor U6417 (N_6417,N_4124,N_3420);
nand U6418 (N_6418,N_3837,N_3614);
nand U6419 (N_6419,N_5604,N_4569);
and U6420 (N_6420,N_4293,N_5046);
or U6421 (N_6421,N_4012,N_5970);
nand U6422 (N_6422,N_4492,N_3516);
nand U6423 (N_6423,N_3466,N_4264);
and U6424 (N_6424,N_5992,N_4919);
and U6425 (N_6425,N_4368,N_5454);
nand U6426 (N_6426,N_5481,N_5598);
nand U6427 (N_6427,N_3344,N_4341);
nor U6428 (N_6428,N_3996,N_3109);
nand U6429 (N_6429,N_4592,N_4118);
nor U6430 (N_6430,N_4227,N_3784);
or U6431 (N_6431,N_5441,N_3956);
and U6432 (N_6432,N_4869,N_3196);
or U6433 (N_6433,N_3454,N_5139);
nand U6434 (N_6434,N_4860,N_4788);
nor U6435 (N_6435,N_5585,N_3346);
nor U6436 (N_6436,N_5071,N_4007);
nor U6437 (N_6437,N_3026,N_5307);
and U6438 (N_6438,N_3347,N_3363);
nand U6439 (N_6439,N_3383,N_5947);
and U6440 (N_6440,N_5711,N_5075);
or U6441 (N_6441,N_5907,N_3282);
nor U6442 (N_6442,N_3275,N_4183);
and U6443 (N_6443,N_4676,N_4961);
or U6444 (N_6444,N_5114,N_3904);
and U6445 (N_6445,N_3798,N_3813);
and U6446 (N_6446,N_4988,N_4412);
or U6447 (N_6447,N_5283,N_5234);
nor U6448 (N_6448,N_3412,N_3395);
nor U6449 (N_6449,N_4228,N_4312);
or U6450 (N_6450,N_4120,N_3890);
or U6451 (N_6451,N_5266,N_4601);
and U6452 (N_6452,N_5791,N_5374);
nor U6453 (N_6453,N_4367,N_4980);
and U6454 (N_6454,N_5618,N_4789);
nand U6455 (N_6455,N_5098,N_5378);
and U6456 (N_6456,N_3647,N_5251);
or U6457 (N_6457,N_3820,N_4455);
nand U6458 (N_6458,N_3241,N_4926);
and U6459 (N_6459,N_3833,N_4764);
or U6460 (N_6460,N_5452,N_4418);
or U6461 (N_6461,N_5759,N_3135);
xnor U6462 (N_6462,N_3195,N_3165);
nor U6463 (N_6463,N_3548,N_4603);
nand U6464 (N_6464,N_5616,N_5429);
nor U6465 (N_6465,N_5643,N_5858);
nor U6466 (N_6466,N_3845,N_3747);
and U6467 (N_6467,N_4259,N_5510);
and U6468 (N_6468,N_3788,N_5920);
nor U6469 (N_6469,N_3394,N_3599);
and U6470 (N_6470,N_4684,N_3902);
nand U6471 (N_6471,N_4122,N_5996);
xnor U6472 (N_6472,N_4694,N_5324);
or U6473 (N_6473,N_5725,N_4503);
or U6474 (N_6474,N_5704,N_3629);
or U6475 (N_6475,N_5142,N_3701);
or U6476 (N_6476,N_4884,N_4305);
nor U6477 (N_6477,N_3355,N_5842);
or U6478 (N_6478,N_3838,N_4859);
nand U6479 (N_6479,N_3997,N_3335);
nor U6480 (N_6480,N_5246,N_3119);
or U6481 (N_6481,N_4693,N_5720);
and U6482 (N_6482,N_4921,N_4335);
nor U6483 (N_6483,N_3460,N_5764);
or U6484 (N_6484,N_5305,N_5629);
nor U6485 (N_6485,N_3161,N_5896);
and U6486 (N_6486,N_4912,N_4955);
nor U6487 (N_6487,N_4445,N_5427);
or U6488 (N_6488,N_5029,N_5393);
nor U6489 (N_6489,N_3993,N_5744);
or U6490 (N_6490,N_5177,N_3036);
or U6491 (N_6491,N_5838,N_5100);
or U6492 (N_6492,N_3105,N_3736);
nor U6493 (N_6493,N_3608,N_5793);
or U6494 (N_6494,N_5987,N_4121);
or U6495 (N_6495,N_4607,N_4308);
nand U6496 (N_6496,N_3261,N_4169);
or U6497 (N_6497,N_5656,N_5984);
and U6498 (N_6498,N_5434,N_5983);
and U6499 (N_6499,N_4620,N_4605);
and U6500 (N_6500,N_3062,N_3365);
nor U6501 (N_6501,N_4379,N_4968);
nor U6502 (N_6502,N_4371,N_4915);
nand U6503 (N_6503,N_5807,N_5047);
and U6504 (N_6504,N_5847,N_5683);
nand U6505 (N_6505,N_3144,N_4473);
nor U6506 (N_6506,N_4189,N_3907);
nor U6507 (N_6507,N_5956,N_4994);
or U6508 (N_6508,N_5391,N_3093);
nand U6509 (N_6509,N_5341,N_4127);
and U6510 (N_6510,N_3511,N_5533);
nand U6511 (N_6511,N_3899,N_5595);
nor U6512 (N_6512,N_4778,N_3692);
nor U6513 (N_6513,N_4827,N_4239);
and U6514 (N_6514,N_3562,N_3496);
xor U6515 (N_6515,N_5965,N_3461);
nor U6516 (N_6516,N_4054,N_5349);
nand U6517 (N_6517,N_4052,N_4633);
xor U6518 (N_6518,N_4362,N_3464);
nand U6519 (N_6519,N_4391,N_5056);
nand U6520 (N_6520,N_5895,N_3375);
xor U6521 (N_6521,N_5674,N_3712);
or U6522 (N_6522,N_4943,N_4776);
nor U6523 (N_6523,N_4756,N_5981);
nand U6524 (N_6524,N_3612,N_3909);
nor U6525 (N_6525,N_4078,N_4984);
nand U6526 (N_6526,N_5601,N_3849);
and U6527 (N_6527,N_3087,N_4496);
and U6528 (N_6528,N_3085,N_3739);
or U6529 (N_6529,N_5739,N_3939);
or U6530 (N_6530,N_3435,N_3001);
and U6531 (N_6531,N_5205,N_5938);
nand U6532 (N_6532,N_4304,N_5438);
or U6533 (N_6533,N_3074,N_5286);
and U6534 (N_6534,N_3992,N_4907);
nand U6535 (N_6535,N_5405,N_4307);
or U6536 (N_6536,N_5259,N_5520);
and U6537 (N_6537,N_5829,N_3581);
nor U6538 (N_6538,N_4337,N_5282);
and U6539 (N_6539,N_3742,N_5929);
nand U6540 (N_6540,N_5129,N_4557);
nor U6541 (N_6541,N_5624,N_5174);
nand U6542 (N_6542,N_5227,N_5937);
nor U6543 (N_6543,N_4700,N_4397);
and U6544 (N_6544,N_3526,N_5442);
and U6545 (N_6545,N_5358,N_4216);
nand U6546 (N_6546,N_4088,N_3510);
or U6547 (N_6547,N_5613,N_4942);
or U6548 (N_6548,N_5568,N_5021);
and U6549 (N_6549,N_4993,N_5696);
nor U6550 (N_6550,N_4483,N_3572);
and U6551 (N_6551,N_3817,N_3808);
nor U6552 (N_6552,N_4847,N_3639);
nor U6553 (N_6553,N_5269,N_3283);
nor U6554 (N_6554,N_4108,N_5268);
nor U6555 (N_6555,N_4437,N_3610);
nand U6556 (N_6556,N_3402,N_4475);
nand U6557 (N_6557,N_5555,N_3655);
nand U6558 (N_6558,N_3400,N_5781);
nor U6559 (N_6559,N_5474,N_5432);
nand U6560 (N_6560,N_3348,N_3698);
nor U6561 (N_6561,N_5158,N_4885);
and U6562 (N_6562,N_3621,N_5779);
nor U6563 (N_6563,N_3758,N_4970);
xor U6564 (N_6564,N_3326,N_3658);
nor U6565 (N_6565,N_4982,N_5600);
or U6566 (N_6566,N_3554,N_4600);
xnor U6567 (N_6567,N_5473,N_3696);
and U6568 (N_6568,N_5932,N_5952);
nand U6569 (N_6569,N_5411,N_3401);
nand U6570 (N_6570,N_4582,N_3836);
nand U6571 (N_6571,N_5857,N_5160);
nand U6572 (N_6572,N_5925,N_5163);
nor U6573 (N_6573,N_5531,N_4091);
or U6574 (N_6574,N_5794,N_4933);
nand U6575 (N_6575,N_4137,N_4023);
nor U6576 (N_6576,N_4680,N_4028);
or U6577 (N_6577,N_4349,N_4956);
nor U6578 (N_6578,N_4365,N_4498);
or U6579 (N_6579,N_4558,N_5428);
nand U6580 (N_6580,N_3623,N_4696);
nor U6581 (N_6581,N_5771,N_5418);
and U6582 (N_6582,N_4733,N_5826);
or U6583 (N_6583,N_3565,N_5808);
nand U6584 (N_6584,N_3279,N_3020);
nor U6585 (N_6585,N_3783,N_4026);
nand U6586 (N_6586,N_5641,N_3770);
or U6587 (N_6587,N_3340,N_4645);
and U6588 (N_6588,N_5439,N_3913);
and U6589 (N_6589,N_5536,N_4560);
and U6590 (N_6590,N_4086,N_4373);
and U6591 (N_6591,N_4591,N_3908);
or U6592 (N_6592,N_4255,N_4099);
xnor U6593 (N_6593,N_5291,N_4472);
and U6594 (N_6594,N_5688,N_5240);
or U6595 (N_6595,N_4095,N_4581);
and U6596 (N_6596,N_3205,N_3000);
and U6597 (N_6597,N_3524,N_3153);
or U6598 (N_6598,N_5666,N_5729);
and U6599 (N_6599,N_5362,N_3537);
nor U6600 (N_6600,N_4338,N_4301);
or U6601 (N_6601,N_5731,N_3924);
or U6602 (N_6602,N_5265,N_5757);
nor U6603 (N_6603,N_4171,N_3929);
nor U6604 (N_6604,N_4123,N_5686);
nand U6605 (N_6605,N_3376,N_5853);
or U6606 (N_6606,N_5574,N_5355);
or U6607 (N_6607,N_4669,N_3222);
and U6608 (N_6608,N_3194,N_3691);
and U6609 (N_6609,N_5935,N_3177);
or U6610 (N_6610,N_4153,N_4427);
nor U6611 (N_6611,N_5384,N_3081);
nor U6612 (N_6612,N_5825,N_4173);
nor U6613 (N_6613,N_4702,N_5200);
nand U6614 (N_6614,N_5569,N_5490);
nor U6615 (N_6615,N_3167,N_5173);
or U6616 (N_6616,N_3762,N_5909);
or U6617 (N_6617,N_5587,N_4883);
or U6618 (N_6618,N_4748,N_5653);
and U6619 (N_6619,N_3928,N_4800);
and U6620 (N_6620,N_4626,N_4713);
and U6621 (N_6621,N_5060,N_3179);
or U6622 (N_6622,N_3390,N_3591);
nand U6623 (N_6623,N_3010,N_4148);
nor U6624 (N_6624,N_3410,N_3147);
nand U6625 (N_6625,N_5607,N_5366);
nor U6626 (N_6626,N_3149,N_5137);
and U6627 (N_6627,N_5001,N_3958);
and U6628 (N_6628,N_3960,N_5913);
nor U6629 (N_6629,N_3022,N_4991);
or U6630 (N_6630,N_4383,N_3892);
or U6631 (N_6631,N_5284,N_5670);
or U6632 (N_6632,N_5066,N_4160);
and U6633 (N_6633,N_4158,N_4425);
and U6634 (N_6634,N_5661,N_3755);
and U6635 (N_6635,N_3961,N_5494);
and U6636 (N_6636,N_5774,N_4760);
and U6637 (N_6637,N_3290,N_4066);
nor U6638 (N_6638,N_4344,N_5832);
and U6639 (N_6639,N_4021,N_3964);
xor U6640 (N_6640,N_3267,N_4032);
and U6641 (N_6641,N_4590,N_4036);
or U6642 (N_6642,N_5815,N_3835);
or U6643 (N_6643,N_3407,N_5786);
or U6644 (N_6644,N_3013,N_5724);
nor U6645 (N_6645,N_4369,N_4814);
nand U6646 (N_6646,N_5395,N_4049);
or U6647 (N_6647,N_4829,N_3227);
nor U6648 (N_6648,N_5930,N_4648);
nand U6649 (N_6649,N_5541,N_4548);
xor U6650 (N_6650,N_5883,N_3915);
or U6651 (N_6651,N_3665,N_5233);
and U6652 (N_6652,N_5176,N_5899);
and U6653 (N_6653,N_3166,N_3032);
nand U6654 (N_6654,N_3574,N_3954);
nand U6655 (N_6655,N_5663,N_4098);
or U6656 (N_6656,N_5322,N_4946);
and U6657 (N_6657,N_3015,N_3752);
and U6658 (N_6658,N_4424,N_3715);
nor U6659 (N_6659,N_3080,N_4936);
nand U6660 (N_6660,N_4217,N_3136);
nor U6661 (N_6661,N_4668,N_3068);
nor U6662 (N_6662,N_5204,N_4388);
nand U6663 (N_6663,N_3342,N_4728);
nor U6664 (N_6664,N_3640,N_3252);
and U6665 (N_6665,N_3979,N_4731);
or U6666 (N_6666,N_5209,N_4586);
nor U6667 (N_6667,N_4699,N_4583);
or U6668 (N_6668,N_5941,N_5295);
or U6669 (N_6669,N_3059,N_3903);
or U6670 (N_6670,N_5682,N_3841);
nor U6671 (N_6671,N_3498,N_5018);
or U6672 (N_6672,N_4754,N_5562);
nand U6673 (N_6673,N_5798,N_4602);
nor U6674 (N_6674,N_5978,N_3937);
and U6675 (N_6675,N_5926,N_5565);
or U6676 (N_6676,N_5865,N_4813);
or U6677 (N_6677,N_5699,N_5824);
nand U6678 (N_6678,N_4740,N_4039);
nor U6679 (N_6679,N_5030,N_5090);
and U6680 (N_6680,N_5313,N_4505);
nor U6681 (N_6681,N_5998,N_4327);
and U6682 (N_6682,N_5827,N_5626);
nand U6683 (N_6683,N_4446,N_4232);
nand U6684 (N_6684,N_4253,N_4930);
or U6685 (N_6685,N_3108,N_4958);
or U6686 (N_6686,N_3819,N_3053);
and U6687 (N_6687,N_4654,N_3600);
nor U6688 (N_6688,N_5623,N_5545);
nand U6689 (N_6689,N_5975,N_3999);
nand U6690 (N_6690,N_3341,N_5741);
and U6691 (N_6691,N_4613,N_3724);
or U6692 (N_6692,N_4628,N_3190);
and U6693 (N_6693,N_4539,N_3002);
or U6694 (N_6694,N_3880,N_4256);
or U6695 (N_6695,N_5903,N_4317);
nand U6696 (N_6696,N_3876,N_5521);
nor U6697 (N_6697,N_3738,N_4479);
nor U6698 (N_6698,N_3455,N_3171);
nor U6699 (N_6699,N_5924,N_5635);
nor U6700 (N_6700,N_5206,N_4284);
nand U6701 (N_6701,N_4347,N_5440);
and U6702 (N_6702,N_5354,N_5388);
or U6703 (N_6703,N_3544,N_4820);
nor U6704 (N_6704,N_4963,N_3864);
nand U6705 (N_6705,N_4918,N_3501);
nor U6706 (N_6706,N_4671,N_5650);
nor U6707 (N_6707,N_3448,N_5657);
or U6708 (N_6708,N_5777,N_3269);
or U6709 (N_6709,N_5278,N_5024);
nand U6710 (N_6710,N_4571,N_4622);
nor U6711 (N_6711,N_3488,N_3513);
nor U6712 (N_6712,N_3187,N_5398);
or U6713 (N_6713,N_3071,N_3926);
and U6714 (N_6714,N_4440,N_5534);
and U6715 (N_6715,N_5032,N_5121);
nand U6716 (N_6716,N_3787,N_3494);
and U6717 (N_6717,N_5554,N_3185);
nor U6718 (N_6718,N_5033,N_3547);
and U6719 (N_6719,N_4426,N_4608);
nand U6720 (N_6720,N_4060,N_5573);
or U6721 (N_6721,N_3302,N_5679);
nor U6722 (N_6722,N_4068,N_5383);
and U6723 (N_6723,N_5850,N_4398);
xor U6724 (N_6724,N_4230,N_5130);
nor U6725 (N_6725,N_5094,N_5716);
nand U6726 (N_6726,N_5034,N_5298);
or U6727 (N_6727,N_5168,N_5083);
nand U6728 (N_6728,N_3532,N_5994);
nand U6729 (N_6729,N_3449,N_5530);
nand U6730 (N_6730,N_3700,N_4875);
and U6731 (N_6731,N_4345,N_3382);
nand U6732 (N_6732,N_4751,N_4783);
and U6733 (N_6733,N_4596,N_4065);
nor U6734 (N_6734,N_3669,N_3254);
or U6735 (N_6735,N_4113,N_4191);
and U6736 (N_6736,N_4541,N_5000);
nor U6737 (N_6737,N_3440,N_4886);
or U6738 (N_6738,N_5210,N_4117);
and U6739 (N_6739,N_5561,N_3318);
or U6740 (N_6740,N_4927,N_4554);
nor U6741 (N_6741,N_4295,N_4131);
nor U6742 (N_6742,N_3590,N_4266);
and U6743 (N_6743,N_3469,N_4691);
and U6744 (N_6744,N_3916,N_5077);
nor U6745 (N_6745,N_5912,N_3030);
nor U6746 (N_6746,N_3411,N_3831);
nand U6747 (N_6747,N_3215,N_5072);
and U6748 (N_6748,N_5036,N_3253);
or U6749 (N_6749,N_4352,N_3602);
nand U6750 (N_6750,N_4585,N_4978);
nor U6751 (N_6751,N_5015,N_4900);
or U6752 (N_6752,N_5367,N_4247);
or U6753 (N_6753,N_4257,N_3704);
nand U6754 (N_6754,N_4471,N_3917);
nand U6755 (N_6755,N_4975,N_5443);
or U6756 (N_6756,N_3207,N_3684);
and U6757 (N_6757,N_5892,N_3246);
xnor U6758 (N_6758,N_5803,N_5855);
nand U6759 (N_6759,N_5544,N_4856);
nand U6760 (N_6760,N_3037,N_3576);
nand U6761 (N_6761,N_3042,N_3932);
nand U6762 (N_6762,N_4206,N_5147);
and U6763 (N_6763,N_3522,N_4460);
or U6764 (N_6764,N_3235,N_3021);
nand U6765 (N_6765,N_3566,N_3192);
or U6766 (N_6766,N_4106,N_3540);
nor U6767 (N_6767,N_4567,N_3352);
and U6768 (N_6768,N_5676,N_5044);
nor U6769 (N_6769,N_5583,N_5041);
and U6770 (N_6770,N_3332,N_4048);
nand U6771 (N_6771,N_5048,N_3518);
and U6772 (N_6772,N_4199,N_3942);
nand U6773 (N_6773,N_4801,N_5390);
xor U6774 (N_6774,N_4449,N_4316);
and U6775 (N_6775,N_3663,N_3258);
or U6776 (N_6776,N_3778,N_4609);
and U6777 (N_6777,N_4353,N_4935);
xnor U6778 (N_6778,N_5586,N_4270);
nor U6779 (N_6779,N_4523,N_5684);
nand U6780 (N_6780,N_4729,N_3245);
or U6781 (N_6781,N_3553,N_3673);
nor U6782 (N_6782,N_3811,N_3444);
nor U6783 (N_6783,N_4448,N_3870);
and U6784 (N_6784,N_3236,N_5309);
nor U6785 (N_6785,N_5389,N_4396);
nor U6786 (N_6786,N_3580,N_3403);
and U6787 (N_6787,N_5423,N_5316);
nor U6788 (N_6788,N_5922,N_4858);
or U6789 (N_6789,N_4166,N_5809);
and U6790 (N_6790,N_4815,N_4899);
nand U6791 (N_6791,N_3867,N_5419);
or U6792 (N_6792,N_3546,N_3906);
nor U6793 (N_6793,N_3298,N_3385);
or U6794 (N_6794,N_5220,N_3706);
nand U6795 (N_6795,N_4964,N_5936);
or U6796 (N_6796,N_5289,N_4417);
nor U6797 (N_6797,N_4981,N_3424);
or U6798 (N_6798,N_4202,N_3967);
or U6799 (N_6799,N_3028,N_5331);
and U6800 (N_6800,N_3707,N_4840);
nand U6801 (N_6801,N_3694,N_4094);
nor U6802 (N_6802,N_3268,N_4467);
or U6803 (N_6803,N_5086,N_3397);
nand U6804 (N_6804,N_5547,N_5190);
and U6805 (N_6805,N_4504,N_5271);
xor U6806 (N_6806,N_5049,N_4119);
nor U6807 (N_6807,N_4561,N_4690);
and U6808 (N_6808,N_3391,N_3995);
nand U6809 (N_6809,N_5849,N_4929);
nand U6810 (N_6810,N_4500,N_4213);
and U6811 (N_6811,N_5361,N_4870);
nor U6812 (N_6812,N_4925,N_3646);
and U6813 (N_6813,N_3219,N_3441);
and U6814 (N_6814,N_3754,N_3796);
and U6815 (N_6815,N_4777,N_5337);
nand U6816 (N_6816,N_4205,N_5088);
nor U6817 (N_6817,N_4102,N_5213);
or U6818 (N_6818,N_5819,N_5087);
nand U6819 (N_6819,N_5746,N_5523);
nor U6820 (N_6820,N_3055,N_5359);
and U6821 (N_6821,N_3047,N_4064);
and U6822 (N_6822,N_4273,N_4562);
nand U6823 (N_6823,N_5931,N_3078);
and U6824 (N_6824,N_5314,N_3807);
xnor U6825 (N_6825,N_5198,N_5660);
nand U6826 (N_6826,N_5364,N_3163);
and U6827 (N_6827,N_5356,N_4898);
or U6828 (N_6828,N_4000,N_4336);
nand U6829 (N_6829,N_4018,N_4080);
or U6830 (N_6830,N_5171,N_4013);
or U6831 (N_6831,N_3757,N_4441);
nand U6832 (N_6832,N_4107,N_5537);
nor U6833 (N_6833,N_5667,N_5564);
nand U6834 (N_6834,N_3726,N_3751);
and U6835 (N_6835,N_5408,N_5915);
or U6836 (N_6836,N_3247,N_3181);
nor U6837 (N_6837,N_3824,N_5887);
or U6838 (N_6838,N_3027,N_4868);
or U6839 (N_6839,N_4570,N_3969);
or U6840 (N_6840,N_3425,N_3570);
nor U6841 (N_6841,N_4149,N_5964);
nand U6842 (N_6842,N_5606,N_5165);
or U6843 (N_6843,N_4494,N_3611);
or U6844 (N_6844,N_3038,N_5906);
or U6845 (N_6845,N_5801,N_4144);
and U6846 (N_6846,N_5078,N_5763);
and U6847 (N_6847,N_5460,N_4277);
nor U6848 (N_6848,N_3209,N_3982);
and U6849 (N_6849,N_3502,N_3509);
nand U6850 (N_6850,N_3569,N_4837);
or U6851 (N_6851,N_3506,N_3652);
nand U6852 (N_6852,N_4867,N_4641);
or U6853 (N_6853,N_3057,N_3688);
nor U6854 (N_6854,N_5485,N_3644);
nand U6855 (N_6855,N_3632,N_5080);
nand U6856 (N_6856,N_3567,N_5622);
nor U6857 (N_6857,N_4717,N_3442);
and U6858 (N_6858,N_4193,N_3061);
or U6859 (N_6859,N_4058,N_4705);
and U6860 (N_6860,N_5280,N_5507);
and U6861 (N_6861,N_3364,N_5726);
or U6862 (N_6862,N_4204,N_3946);
nor U6863 (N_6863,N_3284,N_5131);
and U6864 (N_6864,N_5343,N_3682);
nand U6865 (N_6865,N_5894,N_3295);
or U6866 (N_6866,N_3480,N_4395);
or U6867 (N_6867,N_3064,N_5211);
nand U6868 (N_6868,N_5839,N_4214);
nor U6869 (N_6869,N_4782,N_4363);
nand U6870 (N_6870,N_4848,N_5869);
or U6871 (N_6871,N_3850,N_4399);
or U6872 (N_6872,N_3528,N_4809);
or U6873 (N_6873,N_4357,N_4485);
and U6874 (N_6874,N_4647,N_3809);
or U6875 (N_6875,N_3023,N_5345);
or U6876 (N_6876,N_5848,N_4897);
and U6877 (N_6877,N_4141,N_4831);
or U6878 (N_6878,N_3152,N_4830);
nor U6879 (N_6879,N_5186,N_3202);
and U6880 (N_6880,N_4101,N_3863);
and U6881 (N_6881,N_4750,N_5040);
nand U6882 (N_6882,N_3914,N_4167);
nor U6883 (N_6883,N_4752,N_3004);
or U6884 (N_6884,N_4400,N_3145);
or U6885 (N_6885,N_4134,N_4874);
and U6886 (N_6886,N_5579,N_5208);
or U6887 (N_6887,N_3603,N_5004);
nand U6888 (N_6888,N_3664,N_4457);
or U6889 (N_6889,N_5377,N_5662);
nor U6890 (N_6890,N_3859,N_5297);
and U6891 (N_6891,N_3124,N_4432);
nand U6892 (N_6892,N_3468,N_4025);
nand U6893 (N_6893,N_5789,N_4909);
nand U6894 (N_6894,N_3507,N_3922);
nor U6895 (N_6895,N_3322,N_5143);
nor U6896 (N_6896,N_3710,N_4775);
and U6897 (N_6897,N_4268,N_3118);
nand U6898 (N_6898,N_4768,N_4194);
nand U6899 (N_6899,N_4092,N_3650);
and U6900 (N_6900,N_5615,N_3605);
nor U6901 (N_6901,N_3573,N_4186);
or U6902 (N_6902,N_4611,N_4616);
or U6903 (N_6903,N_5796,N_4525);
or U6904 (N_6904,N_3858,N_5939);
nand U6905 (N_6905,N_5216,N_4276);
xnor U6906 (N_6906,N_5104,N_4219);
nor U6907 (N_6907,N_5333,N_5581);
and U6908 (N_6908,N_3281,N_4016);
nand U6909 (N_6909,N_3033,N_5476);
or U6910 (N_6910,N_3843,N_3896);
xnor U6911 (N_6911,N_4761,N_3463);
and U6912 (N_6912,N_4630,N_4634);
nand U6913 (N_6913,N_5910,N_3560);
nor U6914 (N_6914,N_4709,N_5690);
nor U6915 (N_6915,N_3842,N_5762);
and U6916 (N_6916,N_5301,N_3389);
nand U6917 (N_6917,N_3421,N_3832);
and U6918 (N_6918,N_5893,N_5862);
and U6919 (N_6919,N_4105,N_5169);
or U6920 (N_6920,N_5117,N_5126);
nand U6921 (N_6921,N_3527,N_5880);
xnor U6922 (N_6922,N_5059,N_4111);
and U6923 (N_6923,N_4799,N_5277);
nor U6924 (N_6924,N_4346,N_3457);
and U6925 (N_6925,N_3897,N_4534);
nor U6926 (N_6926,N_3977,N_4810);
nand U6927 (N_6927,N_5218,N_5873);
nor U6928 (N_6928,N_3753,N_3577);
nand U6929 (N_6929,N_3685,N_3270);
nand U6930 (N_6930,N_4350,N_4771);
nand U6931 (N_6931,N_5758,N_3183);
nor U6932 (N_6932,N_5576,N_4808);
and U6933 (N_6933,N_3381,N_5437);
nor U6934 (N_6934,N_5272,N_4063);
and U6935 (N_6935,N_4766,N_5681);
nand U6936 (N_6936,N_3482,N_3433);
or U6937 (N_6937,N_5963,N_3377);
or U6938 (N_6938,N_3936,N_4625);
nor U6939 (N_6939,N_5466,N_3846);
and U6940 (N_6940,N_4325,N_3359);
and U6941 (N_6941,N_3792,N_5276);
xnor U6942 (N_6942,N_4576,N_5185);
nor U6943 (N_6943,N_4200,N_4468);
nor U6944 (N_6944,N_3601,N_4983);
or U6945 (N_6945,N_4474,N_5068);
and U6946 (N_6946,N_5860,N_3713);
nand U6947 (N_6947,N_3351,N_5646);
nor U6948 (N_6948,N_5436,N_5955);
nand U6949 (N_6949,N_4832,N_4089);
nor U6950 (N_6950,N_3361,N_4244);
nor U6951 (N_6951,N_3110,N_4055);
or U6952 (N_6952,N_3523,N_4857);
nor U6953 (N_6953,N_5020,N_4387);
and U6954 (N_6954,N_5976,N_3251);
and U6955 (N_6955,N_5594,N_4575);
or U6956 (N_6956,N_4887,N_5636);
nor U6957 (N_6957,N_3308,N_5773);
nor U6958 (N_6958,N_5572,N_4034);
and U6959 (N_6959,N_5187,N_4182);
xnor U6960 (N_6960,N_3886,N_3720);
nor U6961 (N_6961,N_4632,N_5988);
or U6962 (N_6962,N_5589,N_5175);
and U6963 (N_6963,N_4300,N_4299);
and U6964 (N_6964,N_4917,N_3198);
or U6965 (N_6965,N_4465,N_4737);
and U6966 (N_6966,N_3830,N_4573);
or U6967 (N_6967,N_3328,N_5563);
nor U6968 (N_6968,N_3073,N_5630);
or U6969 (N_6969,N_5821,N_4081);
or U6970 (N_6970,N_3851,N_5407);
or U6971 (N_6971,N_3193,N_3981);
or U6972 (N_6972,N_3957,N_5172);
nand U6973 (N_6973,N_4865,N_3262);
nor U6974 (N_6974,N_3160,N_4517);
or U6975 (N_6975,N_5381,N_4688);
nor U6976 (N_6976,N_3743,N_5231);
and U6977 (N_6977,N_5065,N_4643);
nor U6978 (N_6978,N_5064,N_4265);
or U6979 (N_6979,N_4243,N_4552);
nor U6980 (N_6980,N_3011,N_4310);
and U6981 (N_6981,N_4949,N_3316);
and U6982 (N_6982,N_3012,N_3578);
or U6983 (N_6983,N_3070,N_3321);
or U6984 (N_6984,N_3968,N_4133);
and U6985 (N_6985,N_4762,N_3393);
xor U6986 (N_6986,N_3199,N_5404);
nor U6987 (N_6987,N_4287,N_3117);
and U6988 (N_6988,N_4002,N_3976);
and U6989 (N_6989,N_5556,N_5877);
and U6990 (N_6990,N_5203,N_5558);
nand U6991 (N_6991,N_4071,N_5069);
nand U6992 (N_6992,N_5971,N_5245);
xnor U6993 (N_6993,N_4724,N_5058);
nand U6994 (N_6994,N_4381,N_5312);
nor U6995 (N_6995,N_4597,N_4017);
nand U6996 (N_6996,N_3286,N_5396);
nand U6997 (N_6997,N_3878,N_5723);
and U6998 (N_6998,N_5508,N_5472);
or U6999 (N_6999,N_4290,N_4458);
nand U7000 (N_7000,N_3329,N_4488);
nor U7001 (N_7001,N_4913,N_5372);
or U7002 (N_7002,N_5516,N_5351);
and U7003 (N_7003,N_5768,N_4175);
or U7004 (N_7004,N_4224,N_5972);
nor U7005 (N_7005,N_3367,N_4985);
nor U7006 (N_7006,N_3007,N_4249);
nor U7007 (N_7007,N_3970,N_4861);
or U7008 (N_7008,N_4421,N_5426);
nand U7009 (N_7009,N_3191,N_3985);
nor U7010 (N_7010,N_5867,N_3826);
nand U7011 (N_7011,N_5446,N_5116);
nor U7012 (N_7012,N_3952,N_3086);
or U7013 (N_7013,N_4521,N_3667);
nor U7014 (N_7014,N_5258,N_5260);
nor U7015 (N_7015,N_3756,N_5578);
or U7016 (N_7016,N_3234,N_5191);
and U7017 (N_7017,N_3184,N_4392);
nand U7018 (N_7018,N_3005,N_5659);
nor U7019 (N_7019,N_3497,N_3409);
nor U7020 (N_7020,N_3920,N_3098);
nor U7021 (N_7021,N_3319,N_3607);
nand U7022 (N_7022,N_3947,N_5115);
xor U7023 (N_7023,N_5665,N_4807);
and U7024 (N_7024,N_4640,N_5009);
nor U7025 (N_7025,N_4319,N_3771);
or U7026 (N_7026,N_3138,N_5612);
nand U7027 (N_7027,N_4242,N_5105);
nand U7028 (N_7028,N_4793,N_5136);
nor U7029 (N_7029,N_5946,N_5525);
and U7030 (N_7030,N_3705,N_4209);
nor U7031 (N_7031,N_5835,N_5756);
and U7032 (N_7032,N_3099,N_3800);
nor U7033 (N_7033,N_4326,N_5323);
nand U7034 (N_7034,N_5344,N_5119);
nand U7035 (N_7035,N_5127,N_4361);
and U7036 (N_7036,N_5188,N_5743);
xnor U7037 (N_7037,N_4128,N_3333);
or U7038 (N_7038,N_5619,N_3812);
nand U7039 (N_7039,N_4817,N_5140);
and U7040 (N_7040,N_4610,N_4281);
or U7041 (N_7041,N_4821,N_5575);
nor U7042 (N_7042,N_4797,N_4535);
nor U7043 (N_7043,N_5350,N_5463);
xnor U7044 (N_7044,N_4951,N_4176);
nand U7045 (N_7045,N_5145,N_4587);
or U7046 (N_7046,N_3934,N_4549);
and U7047 (N_7047,N_4235,N_4402);
and U7048 (N_7048,N_3635,N_3686);
nor U7049 (N_7049,N_3445,N_4798);
xor U7050 (N_7050,N_4414,N_3220);
nor U7051 (N_7051,N_4652,N_4161);
nor U7052 (N_7052,N_5236,N_3197);
nor U7053 (N_7053,N_3680,N_4804);
nor U7054 (N_7054,N_5394,N_5694);
nand U7055 (N_7055,N_3895,N_4852);
xor U7056 (N_7056,N_5503,N_5714);
nand U7057 (N_7057,N_3987,N_3649);
nand U7058 (N_7058,N_4340,N_4478);
or U7059 (N_7059,N_5247,N_5483);
nor U7060 (N_7060,N_4791,N_5232);
nor U7061 (N_7061,N_5201,N_4682);
nand U7062 (N_7062,N_3711,N_5811);
and U7063 (N_7063,N_4922,N_3292);
and U7064 (N_7064,N_5495,N_5401);
nor U7065 (N_7065,N_4838,N_5617);
or U7066 (N_7066,N_4741,N_5017);
and U7067 (N_7067,N_3492,N_4129);
nor U7068 (N_7068,N_4003,N_4155);
or U7069 (N_7069,N_4538,N_3097);
and U7070 (N_7070,N_3627,N_4987);
and U7071 (N_7071,N_3083,N_4035);
nand U7072 (N_7072,N_5097,N_4419);
or U7073 (N_7073,N_4689,N_5761);
or U7074 (N_7074,N_4274,N_4429);
or U7075 (N_7075,N_3584,N_5249);
or U7076 (N_7076,N_5416,N_4836);
or U7077 (N_7077,N_5863,N_4619);
nor U7078 (N_7078,N_5431,N_3776);
or U7079 (N_7079,N_3871,N_5074);
nor U7080 (N_7080,N_3861,N_5856);
and U7081 (N_7081,N_5102,N_5202);
nor U7082 (N_7082,N_3714,N_3839);
nand U7083 (N_7083,N_5859,N_3309);
and U7084 (N_7084,N_4386,N_5833);
xor U7085 (N_7085,N_3041,N_4279);
or U7086 (N_7086,N_3552,N_5370);
nor U7087 (N_7087,N_4736,N_3415);
nor U7088 (N_7088,N_4096,N_5477);
or U7089 (N_7089,N_4151,N_5708);
and U7090 (N_7090,N_3024,N_3990);
nor U7091 (N_7091,N_4180,N_4787);
nor U7092 (N_7092,N_3617,N_4079);
and U7093 (N_7093,N_5150,N_3373);
or U7094 (N_7094,N_4780,N_4655);
nor U7095 (N_7095,N_5775,N_4172);
nand U7096 (N_7096,N_5493,N_5123);
or U7097 (N_7097,N_5628,N_3123);
nand U7098 (N_7098,N_4220,N_4006);
or U7099 (N_7099,N_3888,N_5712);
nor U7100 (N_7100,N_5016,N_5456);
nor U7101 (N_7101,N_5884,N_5229);
nand U7102 (N_7102,N_4311,N_4824);
nand U7103 (N_7103,N_3535,N_4631);
nor U7104 (N_7104,N_5904,N_5195);
nor U7105 (N_7105,N_5529,N_3514);
or U7106 (N_7106,N_3793,N_4896);
nor U7107 (N_7107,N_3829,N_3534);
or U7108 (N_7108,N_5261,N_3759);
nand U7109 (N_7109,N_5968,N_4447);
and U7110 (N_7110,N_3146,N_4184);
and U7111 (N_7111,N_5897,N_5745);
or U7112 (N_7112,N_4511,N_5222);
nor U7113 (N_7113,N_3330,N_3828);
nor U7114 (N_7114,N_5914,N_5415);
or U7115 (N_7115,N_3151,N_3439);
and U7116 (N_7116,N_4495,N_4759);
and U7117 (N_7117,N_3966,N_3017);
xnor U7118 (N_7118,N_4851,N_5054);
and U7119 (N_7119,N_5715,N_5854);
nand U7120 (N_7120,N_4674,N_4971);
or U7121 (N_7121,N_4673,N_5089);
and U7122 (N_7122,N_3297,N_3338);
and U7123 (N_7123,N_3678,N_4537);
nand U7124 (N_7124,N_5900,N_4803);
nor U7125 (N_7125,N_5368,N_4952);
nor U7126 (N_7126,N_3485,N_5287);
xor U7127 (N_7127,N_3910,N_4816);
nor U7128 (N_7128,N_5073,N_5957);
nor U7129 (N_7129,N_5755,N_5376);
nor U7130 (N_7130,N_4902,N_5780);
nor U7131 (N_7131,N_4225,N_5363);
nor U7132 (N_7132,N_5467,N_3874);
and U7133 (N_7133,N_3417,N_5878);
nor U7134 (N_7134,N_5099,N_3091);
or U7135 (N_7135,N_5120,N_4546);
nand U7136 (N_7136,N_5141,N_5486);
nor U7137 (N_7137,N_3189,N_3894);
nor U7138 (N_7138,N_5655,N_4163);
nor U7139 (N_7139,N_3884,N_4057);
or U7140 (N_7140,N_4248,N_4977);
nand U7141 (N_7141,N_5535,N_3387);
nand U7142 (N_7142,N_3242,N_3727);
or U7143 (N_7143,N_5294,N_5875);
and U7144 (N_7144,N_3785,N_4572);
nor U7145 (N_7145,N_4588,N_4354);
nor U7146 (N_7146,N_3312,N_5459);
or U7147 (N_7147,N_5250,N_5332);
nand U7148 (N_7148,N_4532,N_4790);
nor U7149 (N_7149,N_3168,N_5489);
nand U7150 (N_7150,N_4038,N_5499);
or U7151 (N_7151,N_5917,N_4090);
nor U7152 (N_7152,N_5334,N_3779);
or U7153 (N_7153,N_4085,N_5802);
nand U7154 (N_7154,N_4318,N_3531);
nor U7155 (N_7155,N_3141,N_3847);
nor U7156 (N_7156,N_4727,N_5695);
nor U7157 (N_7157,N_3325,N_4931);
and U7158 (N_7158,N_3465,N_3213);
and U7159 (N_7159,N_4377,N_5496);
nand U7160 (N_7160,N_3860,N_5818);
and U7161 (N_7161,N_4372,N_4681);
or U7162 (N_7162,N_3029,N_4033);
and U7163 (N_7163,N_5840,N_4223);
nor U7164 (N_7164,N_3103,N_5995);
nor U7165 (N_7165,N_3885,N_5813);
and U7166 (N_7166,N_5817,N_5096);
and U7167 (N_7167,N_5469,N_4528);
and U7168 (N_7168,N_4420,N_3703);
or U7169 (N_7169,N_3408,N_5966);
and U7170 (N_7170,N_3462,N_3471);
nand U7171 (N_7171,N_4547,N_5273);
and U7172 (N_7172,N_4604,N_3446);
nor U7173 (N_7173,N_3049,N_3288);
nor U7174 (N_7174,N_3060,N_4442);
and U7175 (N_7175,N_5750,N_3089);
xnor U7176 (N_7176,N_3008,N_3285);
or U7177 (N_7177,N_3419,N_3582);
nand U7178 (N_7178,N_4849,N_5687);
nand U7179 (N_7179,N_5076,N_5542);
or U7180 (N_7180,N_5805,N_3781);
nor U7181 (N_7181,N_5782,N_3423);
nor U7182 (N_7182,N_5747,N_3855);
and U7183 (N_7183,N_4283,N_4646);
or U7184 (N_7184,N_4508,N_3035);
nor U7185 (N_7185,N_4882,N_3816);
or U7186 (N_7186,N_5792,N_3406);
or U7187 (N_7187,N_4074,N_4481);
and U7188 (N_7188,N_3980,N_5765);
or U7189 (N_7189,N_4730,N_3458);
or U7190 (N_7190,N_5006,N_4168);
and U7191 (N_7191,N_3479,N_3780);
xor U7192 (N_7192,N_3962,N_4005);
nand U7193 (N_7193,N_3500,N_4834);
nor U7194 (N_7194,N_3345,N_4462);
nor U7195 (N_7195,N_3102,N_5031);
nand U7196 (N_7196,N_5760,N_4624);
nor U7197 (N_7197,N_3277,N_5325);
nor U7198 (N_7198,N_5183,N_4565);
nor U7199 (N_7199,N_3973,N_3077);
and U7200 (N_7200,N_3172,N_3499);
or U7201 (N_7201,N_3208,N_5422);
nand U7202 (N_7202,N_5567,N_5290);
or U7203 (N_7203,N_3633,N_5933);
and U7204 (N_7204,N_4950,N_5960);
xor U7205 (N_7205,N_4514,N_4992);
or U7206 (N_7206,N_4706,N_3173);
nand U7207 (N_7207,N_3775,N_4629);
nand U7208 (N_7208,N_3571,N_4043);
and U7209 (N_7209,N_3140,N_3542);
nand U7210 (N_7210,N_5392,N_3096);
or U7211 (N_7211,N_5478,N_4009);
and U7212 (N_7212,N_5409,N_3238);
and U7213 (N_7213,N_4221,N_3467);
and U7214 (N_7214,N_5698,N_3076);
and U7215 (N_7215,N_3211,N_3473);
nand U7216 (N_7216,N_3203,N_3045);
xnor U7217 (N_7217,N_5125,N_4888);
or U7218 (N_7218,N_5548,N_4433);
and U7219 (N_7219,N_4578,N_4833);
nand U7220 (N_7220,N_3299,N_4084);
and U7221 (N_7221,N_5225,N_4285);
or U7222 (N_7222,N_4784,N_4218);
xor U7223 (N_7223,N_3495,N_4116);
or U7224 (N_7224,N_4008,N_3636);
or U7225 (N_7225,N_4136,N_4769);
nor U7226 (N_7226,N_5468,N_3216);
nor U7227 (N_7227,N_3418,N_3265);
or U7228 (N_7228,N_3643,N_5934);
nor U7229 (N_7229,N_3905,N_3797);
xnor U7230 (N_7230,N_3763,N_5230);
nor U7231 (N_7231,N_5352,N_4275);
nor U7232 (N_7232,N_5868,N_5134);
and U7233 (N_7233,N_5027,N_4529);
and U7234 (N_7234,N_5166,N_5591);
nor U7235 (N_7235,N_4267,N_5675);
and U7236 (N_7236,N_3550,N_3687);
or U7237 (N_7237,N_3991,N_3307);
xnor U7238 (N_7238,N_4584,N_4726);
nor U7239 (N_7239,N_3478,N_4409);
and U7240 (N_7240,N_5444,N_4044);
or U7241 (N_7241,N_5977,N_4262);
or U7242 (N_7242,N_4181,N_4489);
nor U7243 (N_7243,N_4940,N_4675);
nand U7244 (N_7244,N_5778,N_5500);
nand U7245 (N_7245,N_5874,N_3229);
nand U7246 (N_7246,N_4828,N_4229);
and U7247 (N_7247,N_5672,N_5621);
and U7248 (N_7248,N_3113,N_3737);
or U7249 (N_7249,N_5308,N_3606);
nor U7250 (N_7250,N_4466,N_5951);
or U7251 (N_7251,N_5788,N_4826);
nand U7252 (N_7252,N_5288,N_3586);
or U7253 (N_7253,N_5837,N_3825);
or U7254 (N_7254,N_5570,N_3009);
nor U7255 (N_7255,N_4792,N_5082);
and U7256 (N_7256,N_4322,N_4718);
and U7257 (N_7257,N_3226,N_3452);
and U7258 (N_7258,N_3721,N_4893);
nor U7259 (N_7259,N_5400,N_3681);
nand U7260 (N_7260,N_5002,N_5797);
nand U7261 (N_7261,N_5402,N_3223);
nand U7262 (N_7262,N_5515,N_5371);
or U7263 (N_7263,N_4422,N_4110);
and U7264 (N_7264,N_4083,N_4324);
nand U7265 (N_7265,N_5043,N_4559);
nor U7266 (N_7266,N_3891,N_3949);
nand U7267 (N_7267,N_5019,N_4976);
and U7268 (N_7268,N_5844,N_3453);
or U7269 (N_7269,N_5889,N_3237);
and U7270 (N_7270,N_5421,N_4087);
nor U7271 (N_7271,N_4359,N_3427);
nor U7272 (N_7272,N_3043,N_5342);
nand U7273 (N_7273,N_5081,N_3370);
nand U7274 (N_7274,N_5011,N_4531);
or U7275 (N_7275,N_3730,N_4280);
nand U7276 (N_7276,N_3805,N_3266);
and U7277 (N_7277,N_3668,N_3709);
nand U7278 (N_7278,N_5050,N_4296);
nor U7279 (N_7279,N_3372,N_3386);
nand U7280 (N_7280,N_3126,N_5028);
and U7281 (N_7281,N_4203,N_3671);
nor U7282 (N_7282,N_3311,N_4891);
and U7283 (N_7283,N_5375,N_3619);
nand U7284 (N_7284,N_3772,N_3170);
nand U7285 (N_7285,N_4272,N_5471);
nor U7286 (N_7286,N_3116,N_5959);
or U7287 (N_7287,N_4112,N_3725);
and U7288 (N_7288,N_5336,N_3525);
or U7289 (N_7289,N_3517,N_4854);
nand U7290 (N_7290,N_4042,N_4650);
and U7291 (N_7291,N_3795,N_5841);
or U7292 (N_7292,N_5770,N_3255);
nor U7293 (N_7293,N_4140,N_3750);
nor U7294 (N_7294,N_4989,N_5067);
nand U7295 (N_7295,N_5403,N_5310);
nand U7296 (N_7296,N_3075,N_5296);
and U7297 (N_7297,N_4159,N_5742);
xor U7298 (N_7298,N_5881,N_4384);
or U7299 (N_7299,N_5701,N_5540);
and U7300 (N_7300,N_3396,N_4482);
xor U7301 (N_7301,N_5577,N_3156);
or U7302 (N_7302,N_5318,N_4594);
nor U7303 (N_7303,N_5328,N_4027);
and U7304 (N_7304,N_3693,N_4170);
or U7305 (N_7305,N_5713,N_5057);
nand U7306 (N_7306,N_5605,N_4880);
or U7307 (N_7307,N_5161,N_4873);
and U7308 (N_7308,N_4659,N_3206);
or U7309 (N_7309,N_4962,N_3777);
xor U7310 (N_7310,N_4947,N_4157);
nor U7311 (N_7311,N_5689,N_4621);
nor U7312 (N_7312,N_5455,N_4282);
nand U7313 (N_7313,N_3250,N_5846);
and U7314 (N_7314,N_5787,N_3827);
and U7315 (N_7315,N_3092,N_3025);
nand U7316 (N_7316,N_3520,N_4215);
and U7317 (N_7317,N_5700,N_4892);
or U7318 (N_7318,N_4190,N_5908);
nor U7319 (N_7319,N_5719,N_4679);
nor U7320 (N_7320,N_4822,N_4667);
nand U7321 (N_7321,N_5092,N_5450);
and U7322 (N_7322,N_5921,N_3930);
nor U7323 (N_7323,N_3941,N_3066);
or U7324 (N_7324,N_3357,N_5748);
and U7325 (N_7325,N_4238,N_5632);
and U7326 (N_7326,N_5709,N_5285);
nor U7327 (N_7327,N_4732,N_3592);
nor U7328 (N_7328,N_5498,N_3769);
nand U7329 (N_7329,N_5178,N_3188);
nand U7330 (N_7330,N_4463,N_3162);
or U7331 (N_7331,N_3054,N_4328);
and U7332 (N_7332,N_3761,N_3745);
and U7333 (N_7333,N_3642,N_3575);
and U7334 (N_7334,N_4082,N_4179);
or U7335 (N_7335,N_4519,N_5207);
or U7336 (N_7336,N_5164,N_4501);
nor U7337 (N_7337,N_3243,N_5053);
and U7338 (N_7338,N_5882,N_4077);
or U7339 (N_7339,N_5433,N_3046);
and U7340 (N_7340,N_3426,N_5226);
nor U7341 (N_7341,N_3259,N_3154);
nand U7342 (N_7342,N_3593,N_5224);
nand U7343 (N_7343,N_5045,N_5509);
and U7344 (N_7344,N_5891,N_5464);
nand U7345 (N_7345,N_5013,N_5340);
or U7346 (N_7346,N_3641,N_4323);
nand U7347 (N_7347,N_5215,N_5949);
nand U7348 (N_7348,N_3722,N_5658);
nand U7349 (N_7349,N_3044,N_3186);
nand U7350 (N_7350,N_4263,N_5347);
nor U7351 (N_7351,N_3654,N_3765);
and U7352 (N_7352,N_3392,N_3695);
and U7353 (N_7353,N_5484,N_4877);
nand U7354 (N_7354,N_3249,N_3366);
and U7355 (N_7355,N_4871,N_3625);
and U7356 (N_7356,N_3388,N_3716);
or U7357 (N_7357,N_3774,N_4599);
nor U7358 (N_7358,N_5916,N_3120);
nor U7359 (N_7359,N_4945,N_3986);
nor U7360 (N_7360,N_4924,N_5243);
or U7361 (N_7361,N_4188,N_5678);
nand U7362 (N_7362,N_5737,N_3158);
nand U7363 (N_7363,N_3901,N_3746);
or U7364 (N_7364,N_4656,N_3923);
or U7365 (N_7365,N_5654,N_4493);
nand U7366 (N_7366,N_5820,N_4376);
nor U7367 (N_7367,N_4779,N_4522);
nor U7368 (N_7368,N_5584,N_4366);
nor U7369 (N_7369,N_4147,N_5084);
or U7370 (N_7370,N_5182,N_4998);
and U7371 (N_7371,N_3912,N_4653);
nor U7372 (N_7372,N_4451,N_4745);
nand U7373 (N_7373,N_4555,N_4881);
and U7374 (N_7374,N_3416,N_5162);
nand U7375 (N_7375,N_3176,N_3844);
or U7376 (N_7376,N_5192,N_4332);
or U7377 (N_7377,N_4315,N_5958);
nand U7378 (N_7378,N_4145,N_4469);
nor U7379 (N_7379,N_3039,N_4059);
nand U7380 (N_7380,N_3323,N_3218);
or U7381 (N_7381,N_4903,N_4152);
and U7382 (N_7382,N_5967,N_4965);
and U7383 (N_7383,N_5989,N_5872);
nand U7384 (N_7384,N_5103,N_5113);
or U7385 (N_7385,N_4250,N_4606);
and U7386 (N_7386,N_5107,N_4796);
or U7387 (N_7387,N_4001,N_5303);
or U7388 (N_7388,N_4701,N_3789);
nand U7389 (N_7389,N_4453,N_5256);
nand U7390 (N_7390,N_3741,N_5413);
or U7391 (N_7391,N_3155,N_3998);
or U7392 (N_7392,N_3660,N_3432);
nand U7393 (N_7393,N_3233,N_3503);
nand U7394 (N_7394,N_4499,N_3379);
and U7395 (N_7395,N_3679,N_3676);
or U7396 (N_7396,N_4878,N_3210);
or U7397 (N_7397,N_5888,N_3875);
and U7398 (N_7398,N_3273,N_4125);
or U7399 (N_7399,N_4662,N_5196);
or U7400 (N_7400,N_4067,N_3933);
or U7401 (N_7401,N_5513,N_3431);
and U7402 (N_7402,N_4130,N_5055);
and U7403 (N_7403,N_5919,N_5592);
and U7404 (N_7404,N_3536,N_4767);
and U7405 (N_7405,N_4435,N_5406);
or U7406 (N_7406,N_5253,N_3090);
nor U7407 (N_7407,N_4431,N_3978);
and U7408 (N_7408,N_3803,N_3122);
nor U7409 (N_7409,N_4725,N_3289);
nor U7410 (N_7410,N_5546,N_3740);
or U7411 (N_7411,N_4839,N_4835);
and U7412 (N_7412,N_4516,N_5901);
and U7413 (N_7413,N_3869,N_5852);
nor U7414 (N_7414,N_5969,N_3616);
or U7415 (N_7415,N_3564,N_4972);
or U7416 (N_7416,N_5703,N_4786);
and U7417 (N_7417,N_3595,N_5735);
and U7418 (N_7418,N_3362,N_4509);
and U7419 (N_7419,N_3115,N_4595);
nor U7420 (N_7420,N_5702,N_5986);
or U7421 (N_7421,N_4456,N_4997);
nand U7422 (N_7422,N_5991,N_4076);
or U7423 (N_7423,N_3699,N_3853);
and U7424 (N_7424,N_4139,N_4245);
or U7425 (N_7425,N_5845,N_5223);
nor U7426 (N_7426,N_5430,N_4415);
or U7427 (N_7427,N_3822,N_3953);
nand U7428 (N_7428,N_3802,N_3768);
nor U7429 (N_7429,N_5648,N_4841);
nor U7430 (N_7430,N_5154,N_4014);
nand U7431 (N_7431,N_3666,N_5482);
nor U7432 (N_7432,N_3257,N_3628);
and U7433 (N_7433,N_3493,N_3350);
and U7434 (N_7434,N_3428,N_4703);
and U7435 (N_7435,N_3114,N_4292);
or U7436 (N_7436,N_4045,N_5193);
nand U7437 (N_7437,N_5871,N_3983);
or U7438 (N_7438,N_3959,N_3512);
or U7439 (N_7439,N_5085,N_5627);
nand U7440 (N_7440,N_4707,N_5962);
or U7441 (N_7441,N_5387,N_5985);
nor U7442 (N_7442,N_4416,N_4187);
or U7443 (N_7443,N_5640,N_3084);
nor U7444 (N_7444,N_3358,N_5093);
or U7445 (N_7445,N_3773,N_5721);
and U7446 (N_7446,N_5451,N_4375);
or U7447 (N_7447,N_4443,N_4240);
and U7448 (N_7448,N_3645,N_3748);
and U7449 (N_7449,N_5184,N_3476);
and U7450 (N_7450,N_3735,N_3804);
nor U7451 (N_7451,N_5262,N_5132);
nand U7452 (N_7452,N_4405,N_4739);
or U7453 (N_7453,N_3834,N_3050);
and U7454 (N_7454,N_5566,N_5327);
nand U7455 (N_7455,N_3541,N_5633);
and U7456 (N_7456,N_4685,N_4637);
nor U7457 (N_7457,N_4380,N_5785);
and U7458 (N_7458,N_3487,N_4515);
nor U7459 (N_7459,N_3051,N_5902);
nor U7460 (N_7460,N_3343,N_4269);
nor U7461 (N_7461,N_5138,N_5241);
nor U7462 (N_7462,N_5445,N_5453);
nor U7463 (N_7463,N_3201,N_3624);
nor U7464 (N_7464,N_5170,N_5734);
xnor U7465 (N_7465,N_4866,N_5491);
nor U7466 (N_7466,N_4314,N_3613);
and U7467 (N_7467,N_4842,N_4195);
and U7468 (N_7468,N_4041,N_4024);
or U7469 (N_7469,N_3806,N_5861);
or U7470 (N_7470,N_4742,N_5692);
nand U7471 (N_7471,N_4825,N_5685);
nor U7472 (N_7472,N_3244,N_4543);
or U7473 (N_7473,N_5504,N_3965);
or U7474 (N_7474,N_5751,N_5146);
nor U7475 (N_7475,N_3877,N_4355);
xnor U7476 (N_7476,N_5668,N_4428);
and U7477 (N_7477,N_3451,N_5270);
nor U7478 (N_7478,N_5812,N_3003);
nand U7479 (N_7479,N_5412,N_5799);
nor U7480 (N_7480,N_4196,N_3862);
or U7481 (N_7481,N_3305,N_5990);
nor U7482 (N_7482,N_3174,N_3315);
and U7483 (N_7483,N_3127,N_3225);
nand U7484 (N_7484,N_5501,N_4438);
nand U7485 (N_7485,N_4704,N_4719);
nor U7486 (N_7486,N_3594,N_4073);
nand U7487 (N_7487,N_5386,N_5264);
or U7488 (N_7488,N_5961,N_4953);
nand U7489 (N_7489,N_4342,N_5311);
nand U7490 (N_7490,N_3369,N_4934);
nor U7491 (N_7491,N_3112,N_4649);
and U7492 (N_7492,N_5517,N_5254);
or U7493 (N_7493,N_4563,N_5319);
nand U7494 (N_7494,N_4291,N_3239);
nor U7495 (N_7495,N_4635,N_3948);
and U7496 (N_7496,N_4757,N_3598);
nand U7497 (N_7497,N_3398,N_5830);
nor U7498 (N_7498,N_5766,N_5526);
nor U7499 (N_7499,N_3274,N_3872);
or U7500 (N_7500,N_4030,N_4988);
and U7501 (N_7501,N_5695,N_5544);
xnor U7502 (N_7502,N_3678,N_4200);
and U7503 (N_7503,N_4126,N_5648);
nor U7504 (N_7504,N_5938,N_3143);
nor U7505 (N_7505,N_5560,N_5869);
xor U7506 (N_7506,N_5437,N_4623);
or U7507 (N_7507,N_3124,N_5787);
xnor U7508 (N_7508,N_5763,N_4976);
and U7509 (N_7509,N_3390,N_5119);
and U7510 (N_7510,N_3137,N_4939);
or U7511 (N_7511,N_3646,N_5840);
nor U7512 (N_7512,N_5934,N_3244);
nor U7513 (N_7513,N_4184,N_5276);
nand U7514 (N_7514,N_5604,N_3291);
nor U7515 (N_7515,N_4871,N_5437);
nor U7516 (N_7516,N_5179,N_5841);
and U7517 (N_7517,N_5265,N_4350);
or U7518 (N_7518,N_4129,N_4767);
nor U7519 (N_7519,N_3585,N_5613);
and U7520 (N_7520,N_5979,N_5139);
or U7521 (N_7521,N_5281,N_3298);
nor U7522 (N_7522,N_4294,N_4148);
or U7523 (N_7523,N_4200,N_4981);
or U7524 (N_7524,N_5419,N_5501);
nand U7525 (N_7525,N_4384,N_5877);
nand U7526 (N_7526,N_5168,N_3047);
or U7527 (N_7527,N_4784,N_4714);
nor U7528 (N_7528,N_5517,N_3705);
nand U7529 (N_7529,N_3973,N_4037);
nand U7530 (N_7530,N_4144,N_4914);
or U7531 (N_7531,N_4061,N_5175);
and U7532 (N_7532,N_4464,N_5028);
nand U7533 (N_7533,N_5245,N_3085);
or U7534 (N_7534,N_5058,N_5568);
nor U7535 (N_7535,N_4821,N_3885);
and U7536 (N_7536,N_4072,N_3976);
and U7537 (N_7537,N_4000,N_3562);
nand U7538 (N_7538,N_5297,N_4826);
and U7539 (N_7539,N_3554,N_3158);
nor U7540 (N_7540,N_5324,N_5259);
nand U7541 (N_7541,N_5703,N_5962);
nand U7542 (N_7542,N_4523,N_3188);
nand U7543 (N_7543,N_4124,N_3606);
or U7544 (N_7544,N_4634,N_4399);
nor U7545 (N_7545,N_5247,N_4370);
nor U7546 (N_7546,N_3170,N_4440);
nor U7547 (N_7547,N_5023,N_4080);
or U7548 (N_7548,N_3148,N_3722);
nand U7549 (N_7549,N_3251,N_4799);
nor U7550 (N_7550,N_3873,N_3126);
nand U7551 (N_7551,N_4138,N_4351);
or U7552 (N_7552,N_4054,N_4095);
nor U7553 (N_7553,N_4435,N_4321);
and U7554 (N_7554,N_4219,N_4706);
or U7555 (N_7555,N_3239,N_5676);
nand U7556 (N_7556,N_3243,N_3137);
nor U7557 (N_7557,N_4883,N_4305);
or U7558 (N_7558,N_4060,N_5083);
nor U7559 (N_7559,N_5119,N_4905);
nand U7560 (N_7560,N_3770,N_4678);
nand U7561 (N_7561,N_5494,N_3234);
nand U7562 (N_7562,N_3698,N_4119);
nor U7563 (N_7563,N_5456,N_5403);
nor U7564 (N_7564,N_5027,N_5853);
and U7565 (N_7565,N_5981,N_5276);
and U7566 (N_7566,N_4903,N_5883);
nand U7567 (N_7567,N_4827,N_5801);
or U7568 (N_7568,N_3296,N_4833);
nand U7569 (N_7569,N_5544,N_3504);
nor U7570 (N_7570,N_4248,N_5945);
and U7571 (N_7571,N_3083,N_5492);
nor U7572 (N_7572,N_5364,N_4466);
and U7573 (N_7573,N_3412,N_5623);
nor U7574 (N_7574,N_3106,N_5051);
or U7575 (N_7575,N_3485,N_4453);
nor U7576 (N_7576,N_3301,N_4235);
nor U7577 (N_7577,N_5126,N_3032);
and U7578 (N_7578,N_4342,N_3953);
and U7579 (N_7579,N_3499,N_5917);
nand U7580 (N_7580,N_5047,N_3888);
nor U7581 (N_7581,N_5820,N_5839);
nand U7582 (N_7582,N_5539,N_5411);
nor U7583 (N_7583,N_5107,N_3689);
nor U7584 (N_7584,N_5341,N_5493);
nor U7585 (N_7585,N_4606,N_4915);
nor U7586 (N_7586,N_5564,N_5742);
and U7587 (N_7587,N_4960,N_4242);
nand U7588 (N_7588,N_4438,N_3945);
or U7589 (N_7589,N_3652,N_5406);
nand U7590 (N_7590,N_4964,N_5910);
nand U7591 (N_7591,N_3995,N_3259);
or U7592 (N_7592,N_5730,N_3827);
and U7593 (N_7593,N_4018,N_3928);
nor U7594 (N_7594,N_3831,N_5200);
nand U7595 (N_7595,N_3744,N_3738);
nand U7596 (N_7596,N_3360,N_4806);
and U7597 (N_7597,N_5775,N_5901);
and U7598 (N_7598,N_4400,N_3834);
nor U7599 (N_7599,N_5500,N_3505);
nand U7600 (N_7600,N_5403,N_3523);
or U7601 (N_7601,N_4959,N_3185);
nand U7602 (N_7602,N_4192,N_3565);
nand U7603 (N_7603,N_4817,N_4839);
or U7604 (N_7604,N_5113,N_4443);
nor U7605 (N_7605,N_4380,N_3451);
or U7606 (N_7606,N_5533,N_4077);
nor U7607 (N_7607,N_4813,N_5102);
and U7608 (N_7608,N_3727,N_3506);
nor U7609 (N_7609,N_5995,N_4471);
or U7610 (N_7610,N_4225,N_3648);
or U7611 (N_7611,N_4761,N_5012);
and U7612 (N_7612,N_5151,N_5185);
and U7613 (N_7613,N_4905,N_5631);
or U7614 (N_7614,N_4684,N_3514);
nand U7615 (N_7615,N_4422,N_5090);
nor U7616 (N_7616,N_3633,N_3193);
nand U7617 (N_7617,N_4619,N_4385);
nor U7618 (N_7618,N_3861,N_5865);
or U7619 (N_7619,N_5075,N_4019);
and U7620 (N_7620,N_4289,N_5608);
and U7621 (N_7621,N_3697,N_4267);
nor U7622 (N_7622,N_5337,N_3385);
and U7623 (N_7623,N_3518,N_4513);
nand U7624 (N_7624,N_3297,N_5224);
or U7625 (N_7625,N_4479,N_3714);
nor U7626 (N_7626,N_4306,N_3000);
nor U7627 (N_7627,N_3455,N_4130);
nor U7628 (N_7628,N_4277,N_5016);
nand U7629 (N_7629,N_4428,N_4120);
nand U7630 (N_7630,N_4693,N_5022);
nand U7631 (N_7631,N_3570,N_5580);
and U7632 (N_7632,N_3238,N_4341);
and U7633 (N_7633,N_3542,N_5545);
or U7634 (N_7634,N_4268,N_5461);
and U7635 (N_7635,N_4275,N_3462);
nor U7636 (N_7636,N_5746,N_5192);
nor U7637 (N_7637,N_5388,N_3582);
or U7638 (N_7638,N_3702,N_4288);
and U7639 (N_7639,N_3980,N_3998);
and U7640 (N_7640,N_5979,N_4362);
nor U7641 (N_7641,N_5211,N_3010);
and U7642 (N_7642,N_3642,N_3870);
and U7643 (N_7643,N_3716,N_3315);
or U7644 (N_7644,N_4877,N_4678);
nor U7645 (N_7645,N_4453,N_4781);
nor U7646 (N_7646,N_5600,N_4557);
or U7647 (N_7647,N_4266,N_4072);
nor U7648 (N_7648,N_5532,N_3517);
xnor U7649 (N_7649,N_3102,N_4944);
nand U7650 (N_7650,N_3332,N_3288);
nand U7651 (N_7651,N_3429,N_5287);
and U7652 (N_7652,N_4391,N_5571);
nand U7653 (N_7653,N_5892,N_4558);
and U7654 (N_7654,N_4889,N_3583);
nand U7655 (N_7655,N_3638,N_3531);
nor U7656 (N_7656,N_3758,N_5306);
and U7657 (N_7657,N_4921,N_5125);
nand U7658 (N_7658,N_3148,N_4023);
or U7659 (N_7659,N_5808,N_3141);
nand U7660 (N_7660,N_5995,N_5875);
and U7661 (N_7661,N_5241,N_5246);
or U7662 (N_7662,N_5174,N_3715);
nand U7663 (N_7663,N_5903,N_4888);
and U7664 (N_7664,N_5929,N_5631);
nand U7665 (N_7665,N_5815,N_3406);
nand U7666 (N_7666,N_5608,N_5349);
nand U7667 (N_7667,N_3980,N_4293);
and U7668 (N_7668,N_5697,N_3949);
and U7669 (N_7669,N_3079,N_3153);
or U7670 (N_7670,N_5652,N_5991);
and U7671 (N_7671,N_3361,N_5843);
nor U7672 (N_7672,N_5438,N_3710);
or U7673 (N_7673,N_5818,N_5467);
or U7674 (N_7674,N_3810,N_3279);
nand U7675 (N_7675,N_5570,N_3610);
or U7676 (N_7676,N_4471,N_5545);
nand U7677 (N_7677,N_3745,N_5813);
and U7678 (N_7678,N_4427,N_5518);
nor U7679 (N_7679,N_3407,N_3459);
and U7680 (N_7680,N_4652,N_4303);
nand U7681 (N_7681,N_4259,N_3152);
nand U7682 (N_7682,N_4147,N_4813);
nor U7683 (N_7683,N_3611,N_3453);
or U7684 (N_7684,N_5766,N_4459);
nand U7685 (N_7685,N_4678,N_3810);
or U7686 (N_7686,N_3483,N_4277);
nor U7687 (N_7687,N_4278,N_3689);
and U7688 (N_7688,N_3248,N_4401);
nor U7689 (N_7689,N_4897,N_5783);
nand U7690 (N_7690,N_5389,N_4570);
nand U7691 (N_7691,N_5443,N_4402);
or U7692 (N_7692,N_4193,N_5218);
and U7693 (N_7693,N_3557,N_5672);
and U7694 (N_7694,N_4799,N_3443);
nand U7695 (N_7695,N_4703,N_3507);
or U7696 (N_7696,N_4407,N_3180);
nand U7697 (N_7697,N_5515,N_5177);
nand U7698 (N_7698,N_3602,N_5528);
and U7699 (N_7699,N_4498,N_5468);
nor U7700 (N_7700,N_3802,N_4135);
and U7701 (N_7701,N_4972,N_5573);
nor U7702 (N_7702,N_3548,N_5532);
nor U7703 (N_7703,N_4082,N_5683);
and U7704 (N_7704,N_3983,N_5610);
and U7705 (N_7705,N_5901,N_5954);
and U7706 (N_7706,N_5320,N_4560);
nor U7707 (N_7707,N_5457,N_3300);
or U7708 (N_7708,N_5576,N_4425);
nor U7709 (N_7709,N_3957,N_5222);
and U7710 (N_7710,N_3926,N_3435);
nor U7711 (N_7711,N_5248,N_4536);
or U7712 (N_7712,N_4086,N_3203);
nor U7713 (N_7713,N_4545,N_3509);
nor U7714 (N_7714,N_3676,N_3258);
nor U7715 (N_7715,N_5359,N_4907);
nor U7716 (N_7716,N_5414,N_3531);
or U7717 (N_7717,N_5186,N_3279);
nor U7718 (N_7718,N_3587,N_5093);
nor U7719 (N_7719,N_5346,N_5530);
and U7720 (N_7720,N_3757,N_3821);
or U7721 (N_7721,N_5832,N_5513);
nand U7722 (N_7722,N_3182,N_5714);
and U7723 (N_7723,N_3908,N_5142);
or U7724 (N_7724,N_5720,N_3265);
nor U7725 (N_7725,N_3328,N_4761);
nor U7726 (N_7726,N_5741,N_4726);
and U7727 (N_7727,N_5048,N_3361);
and U7728 (N_7728,N_3991,N_5084);
or U7729 (N_7729,N_3509,N_4346);
nand U7730 (N_7730,N_4681,N_3022);
nand U7731 (N_7731,N_5529,N_3557);
nand U7732 (N_7732,N_4928,N_5359);
nor U7733 (N_7733,N_3294,N_4736);
nor U7734 (N_7734,N_4834,N_5785);
nand U7735 (N_7735,N_4373,N_3511);
nand U7736 (N_7736,N_5329,N_4632);
or U7737 (N_7737,N_4697,N_4392);
nor U7738 (N_7738,N_3430,N_5410);
nand U7739 (N_7739,N_5856,N_3097);
and U7740 (N_7740,N_5666,N_4133);
nand U7741 (N_7741,N_5590,N_5616);
nand U7742 (N_7742,N_5401,N_5421);
or U7743 (N_7743,N_3409,N_4004);
or U7744 (N_7744,N_5381,N_3046);
nor U7745 (N_7745,N_3400,N_3440);
xor U7746 (N_7746,N_3875,N_4746);
and U7747 (N_7747,N_5634,N_5994);
nor U7748 (N_7748,N_3916,N_5675);
and U7749 (N_7749,N_4836,N_3480);
xnor U7750 (N_7750,N_3925,N_4478);
nor U7751 (N_7751,N_3677,N_3976);
and U7752 (N_7752,N_3838,N_5824);
nor U7753 (N_7753,N_3829,N_3992);
xnor U7754 (N_7754,N_4852,N_4629);
or U7755 (N_7755,N_5987,N_3430);
and U7756 (N_7756,N_5738,N_3227);
nand U7757 (N_7757,N_3823,N_5895);
nor U7758 (N_7758,N_4716,N_3684);
or U7759 (N_7759,N_5521,N_5862);
nor U7760 (N_7760,N_3600,N_4060);
and U7761 (N_7761,N_3240,N_5969);
and U7762 (N_7762,N_3695,N_4053);
nand U7763 (N_7763,N_5575,N_3204);
xor U7764 (N_7764,N_4126,N_5337);
nor U7765 (N_7765,N_4486,N_5295);
nand U7766 (N_7766,N_5256,N_3873);
nor U7767 (N_7767,N_3223,N_3911);
nor U7768 (N_7768,N_3796,N_5486);
or U7769 (N_7769,N_3092,N_4708);
and U7770 (N_7770,N_5452,N_4669);
or U7771 (N_7771,N_4339,N_3416);
nand U7772 (N_7772,N_4056,N_5162);
nor U7773 (N_7773,N_3570,N_4736);
nand U7774 (N_7774,N_5242,N_3183);
nor U7775 (N_7775,N_3676,N_4336);
nand U7776 (N_7776,N_5564,N_3548);
or U7777 (N_7777,N_5466,N_3445);
and U7778 (N_7778,N_4668,N_3343);
nand U7779 (N_7779,N_3611,N_3512);
and U7780 (N_7780,N_5223,N_5171);
nand U7781 (N_7781,N_5328,N_4522);
nor U7782 (N_7782,N_4019,N_5402);
and U7783 (N_7783,N_4401,N_5743);
nor U7784 (N_7784,N_4445,N_5435);
and U7785 (N_7785,N_5280,N_3709);
nor U7786 (N_7786,N_4552,N_5130);
nand U7787 (N_7787,N_5674,N_4912);
and U7788 (N_7788,N_5078,N_4809);
nand U7789 (N_7789,N_3082,N_5964);
or U7790 (N_7790,N_5496,N_4514);
nor U7791 (N_7791,N_5448,N_5614);
nand U7792 (N_7792,N_3174,N_5810);
nand U7793 (N_7793,N_4075,N_4484);
nor U7794 (N_7794,N_5595,N_4867);
or U7795 (N_7795,N_4384,N_5111);
nor U7796 (N_7796,N_3798,N_3778);
or U7797 (N_7797,N_5923,N_3249);
nor U7798 (N_7798,N_3768,N_4574);
and U7799 (N_7799,N_3545,N_5234);
nor U7800 (N_7800,N_4989,N_5154);
nand U7801 (N_7801,N_5620,N_4220);
xnor U7802 (N_7802,N_5844,N_4032);
and U7803 (N_7803,N_4191,N_5235);
nor U7804 (N_7804,N_3100,N_4294);
nand U7805 (N_7805,N_4571,N_4070);
nor U7806 (N_7806,N_5394,N_3200);
nand U7807 (N_7807,N_3047,N_5561);
and U7808 (N_7808,N_4165,N_5019);
and U7809 (N_7809,N_4257,N_3492);
nand U7810 (N_7810,N_5841,N_5645);
or U7811 (N_7811,N_5400,N_5337);
nand U7812 (N_7812,N_3845,N_3148);
or U7813 (N_7813,N_5115,N_4593);
and U7814 (N_7814,N_3295,N_4408);
or U7815 (N_7815,N_4840,N_5482);
nand U7816 (N_7816,N_3504,N_5687);
nor U7817 (N_7817,N_3240,N_5628);
nor U7818 (N_7818,N_3997,N_5280);
nand U7819 (N_7819,N_4702,N_5466);
nand U7820 (N_7820,N_3989,N_4982);
nor U7821 (N_7821,N_4527,N_5465);
xnor U7822 (N_7822,N_4044,N_3147);
nand U7823 (N_7823,N_4988,N_3940);
nor U7824 (N_7824,N_4833,N_3431);
nor U7825 (N_7825,N_3860,N_5983);
nor U7826 (N_7826,N_4384,N_5602);
nand U7827 (N_7827,N_3773,N_3874);
nand U7828 (N_7828,N_5444,N_4208);
and U7829 (N_7829,N_3596,N_5498);
nand U7830 (N_7830,N_3152,N_5187);
nor U7831 (N_7831,N_3027,N_4461);
nand U7832 (N_7832,N_5110,N_4753);
or U7833 (N_7833,N_5457,N_4978);
or U7834 (N_7834,N_4185,N_3311);
nand U7835 (N_7835,N_4267,N_5748);
or U7836 (N_7836,N_5647,N_5047);
nand U7837 (N_7837,N_3676,N_4377);
or U7838 (N_7838,N_5132,N_3242);
or U7839 (N_7839,N_3487,N_5981);
nand U7840 (N_7840,N_3201,N_4685);
nor U7841 (N_7841,N_3763,N_4588);
nor U7842 (N_7842,N_5744,N_5674);
or U7843 (N_7843,N_5193,N_5617);
and U7844 (N_7844,N_5598,N_5372);
and U7845 (N_7845,N_5963,N_4329);
or U7846 (N_7846,N_3825,N_5079);
xnor U7847 (N_7847,N_3128,N_5999);
and U7848 (N_7848,N_5854,N_5013);
or U7849 (N_7849,N_3297,N_3607);
nand U7850 (N_7850,N_3855,N_3266);
or U7851 (N_7851,N_4558,N_4138);
nor U7852 (N_7852,N_5575,N_5143);
nand U7853 (N_7853,N_3096,N_4955);
or U7854 (N_7854,N_3242,N_4403);
nand U7855 (N_7855,N_3971,N_3918);
and U7856 (N_7856,N_5405,N_5256);
nand U7857 (N_7857,N_4529,N_3898);
or U7858 (N_7858,N_5951,N_5225);
nand U7859 (N_7859,N_4074,N_5518);
and U7860 (N_7860,N_4314,N_3397);
xnor U7861 (N_7861,N_3516,N_5609);
and U7862 (N_7862,N_5239,N_5885);
and U7863 (N_7863,N_4570,N_5048);
or U7864 (N_7864,N_5109,N_3203);
or U7865 (N_7865,N_3679,N_3883);
nand U7866 (N_7866,N_5259,N_4319);
and U7867 (N_7867,N_3134,N_4911);
nand U7868 (N_7868,N_4487,N_3749);
and U7869 (N_7869,N_4912,N_5428);
or U7870 (N_7870,N_5728,N_5225);
nor U7871 (N_7871,N_5666,N_5883);
nor U7872 (N_7872,N_3738,N_5368);
and U7873 (N_7873,N_4961,N_4609);
nand U7874 (N_7874,N_4111,N_3734);
and U7875 (N_7875,N_5512,N_5718);
or U7876 (N_7876,N_5701,N_5189);
nor U7877 (N_7877,N_3094,N_5257);
and U7878 (N_7878,N_3563,N_4595);
nand U7879 (N_7879,N_3384,N_4632);
and U7880 (N_7880,N_5065,N_3977);
and U7881 (N_7881,N_4118,N_5645);
nor U7882 (N_7882,N_4937,N_5848);
and U7883 (N_7883,N_4055,N_4012);
nand U7884 (N_7884,N_3372,N_5940);
and U7885 (N_7885,N_5722,N_3513);
nor U7886 (N_7886,N_5890,N_3225);
nor U7887 (N_7887,N_5972,N_5894);
or U7888 (N_7888,N_5255,N_3295);
and U7889 (N_7889,N_4551,N_4667);
or U7890 (N_7890,N_5555,N_3817);
nor U7891 (N_7891,N_3695,N_4954);
nor U7892 (N_7892,N_4497,N_4895);
and U7893 (N_7893,N_4100,N_4166);
nand U7894 (N_7894,N_3153,N_5074);
and U7895 (N_7895,N_4399,N_5338);
and U7896 (N_7896,N_4701,N_3420);
nor U7897 (N_7897,N_3235,N_3379);
nand U7898 (N_7898,N_3552,N_4232);
or U7899 (N_7899,N_4287,N_4544);
nand U7900 (N_7900,N_3992,N_5582);
nor U7901 (N_7901,N_3749,N_4558);
or U7902 (N_7902,N_3605,N_3976);
nand U7903 (N_7903,N_3839,N_4110);
nor U7904 (N_7904,N_4297,N_3900);
and U7905 (N_7905,N_3730,N_5978);
or U7906 (N_7906,N_3577,N_5779);
nand U7907 (N_7907,N_3861,N_4500);
and U7908 (N_7908,N_3674,N_3015);
nand U7909 (N_7909,N_5474,N_4566);
or U7910 (N_7910,N_5908,N_5934);
nand U7911 (N_7911,N_5384,N_3975);
nor U7912 (N_7912,N_4829,N_5504);
and U7913 (N_7913,N_4820,N_5218);
or U7914 (N_7914,N_3841,N_4288);
and U7915 (N_7915,N_3949,N_3076);
and U7916 (N_7916,N_5007,N_4025);
or U7917 (N_7917,N_3084,N_4983);
and U7918 (N_7918,N_3939,N_4594);
and U7919 (N_7919,N_5123,N_5932);
nor U7920 (N_7920,N_4569,N_4230);
nand U7921 (N_7921,N_4138,N_5489);
nand U7922 (N_7922,N_4975,N_5320);
and U7923 (N_7923,N_3792,N_4507);
or U7924 (N_7924,N_3226,N_4012);
nand U7925 (N_7925,N_3141,N_3300);
nand U7926 (N_7926,N_4583,N_4940);
xor U7927 (N_7927,N_5596,N_3241);
nand U7928 (N_7928,N_3873,N_3871);
and U7929 (N_7929,N_4987,N_4164);
or U7930 (N_7930,N_5878,N_4704);
and U7931 (N_7931,N_5513,N_3181);
and U7932 (N_7932,N_5994,N_4154);
and U7933 (N_7933,N_3835,N_4825);
nor U7934 (N_7934,N_3473,N_3928);
or U7935 (N_7935,N_5484,N_5926);
nor U7936 (N_7936,N_3127,N_4499);
or U7937 (N_7937,N_5249,N_3732);
nor U7938 (N_7938,N_5575,N_5812);
or U7939 (N_7939,N_3901,N_5884);
and U7940 (N_7940,N_3428,N_3345);
nor U7941 (N_7941,N_3783,N_5663);
nand U7942 (N_7942,N_3054,N_4377);
or U7943 (N_7943,N_4225,N_5096);
and U7944 (N_7944,N_3739,N_5127);
nor U7945 (N_7945,N_4275,N_4335);
nand U7946 (N_7946,N_4498,N_4535);
nor U7947 (N_7947,N_3028,N_3324);
nand U7948 (N_7948,N_3929,N_4898);
or U7949 (N_7949,N_5653,N_4088);
or U7950 (N_7950,N_3854,N_5536);
and U7951 (N_7951,N_3163,N_3959);
nor U7952 (N_7952,N_3998,N_5621);
nand U7953 (N_7953,N_5306,N_4446);
nor U7954 (N_7954,N_5556,N_5122);
nor U7955 (N_7955,N_3455,N_3342);
nor U7956 (N_7956,N_3764,N_5355);
and U7957 (N_7957,N_5625,N_5572);
or U7958 (N_7958,N_5223,N_4465);
and U7959 (N_7959,N_5423,N_4469);
nor U7960 (N_7960,N_5926,N_3094);
and U7961 (N_7961,N_3990,N_3065);
nand U7962 (N_7962,N_3880,N_5944);
or U7963 (N_7963,N_3304,N_4651);
and U7964 (N_7964,N_4638,N_5925);
nand U7965 (N_7965,N_4902,N_5010);
and U7966 (N_7966,N_4965,N_5299);
nor U7967 (N_7967,N_3969,N_4162);
xnor U7968 (N_7968,N_5876,N_5885);
nand U7969 (N_7969,N_4394,N_3457);
nor U7970 (N_7970,N_5526,N_3421);
or U7971 (N_7971,N_3704,N_4555);
or U7972 (N_7972,N_5162,N_4771);
nor U7973 (N_7973,N_4147,N_4750);
nand U7974 (N_7974,N_5289,N_5280);
nor U7975 (N_7975,N_5279,N_4878);
and U7976 (N_7976,N_5159,N_5460);
nor U7977 (N_7977,N_3582,N_5517);
or U7978 (N_7978,N_5468,N_3072);
nor U7979 (N_7979,N_4883,N_5526);
or U7980 (N_7980,N_3287,N_3293);
or U7981 (N_7981,N_5515,N_3832);
nand U7982 (N_7982,N_3526,N_3476);
nor U7983 (N_7983,N_3504,N_3734);
and U7984 (N_7984,N_4681,N_4761);
and U7985 (N_7985,N_5017,N_4610);
nor U7986 (N_7986,N_3520,N_5800);
or U7987 (N_7987,N_4860,N_5317);
xnor U7988 (N_7988,N_5486,N_3037);
or U7989 (N_7989,N_3181,N_5033);
and U7990 (N_7990,N_4298,N_4761);
and U7991 (N_7991,N_4321,N_5868);
or U7992 (N_7992,N_4676,N_3484);
or U7993 (N_7993,N_5292,N_4131);
and U7994 (N_7994,N_5190,N_4238);
or U7995 (N_7995,N_5313,N_5759);
or U7996 (N_7996,N_4859,N_5309);
or U7997 (N_7997,N_3409,N_3829);
xnor U7998 (N_7998,N_5040,N_4779);
nand U7999 (N_7999,N_5367,N_3776);
or U8000 (N_8000,N_4739,N_3710);
xor U8001 (N_8001,N_5390,N_5862);
and U8002 (N_8002,N_4552,N_5618);
and U8003 (N_8003,N_3138,N_5828);
nand U8004 (N_8004,N_3430,N_3034);
or U8005 (N_8005,N_3768,N_4685);
nor U8006 (N_8006,N_4580,N_4000);
nor U8007 (N_8007,N_5341,N_5638);
or U8008 (N_8008,N_3020,N_5226);
nand U8009 (N_8009,N_3529,N_3624);
nor U8010 (N_8010,N_5149,N_3126);
and U8011 (N_8011,N_4935,N_5741);
and U8012 (N_8012,N_5847,N_3136);
nand U8013 (N_8013,N_3873,N_4589);
or U8014 (N_8014,N_5910,N_5882);
or U8015 (N_8015,N_4726,N_3307);
or U8016 (N_8016,N_3240,N_3513);
and U8017 (N_8017,N_3146,N_3165);
nor U8018 (N_8018,N_5439,N_3531);
and U8019 (N_8019,N_3160,N_5743);
nand U8020 (N_8020,N_5993,N_3839);
and U8021 (N_8021,N_4926,N_3693);
nand U8022 (N_8022,N_3367,N_3495);
nor U8023 (N_8023,N_5454,N_4741);
nand U8024 (N_8024,N_5262,N_5406);
nor U8025 (N_8025,N_4609,N_5068);
xnor U8026 (N_8026,N_3924,N_3925);
or U8027 (N_8027,N_4399,N_5342);
xor U8028 (N_8028,N_5824,N_3314);
nand U8029 (N_8029,N_5393,N_3026);
nand U8030 (N_8030,N_3205,N_3517);
nor U8031 (N_8031,N_5297,N_3753);
nor U8032 (N_8032,N_5141,N_5973);
nand U8033 (N_8033,N_3448,N_5310);
nor U8034 (N_8034,N_4675,N_3537);
nand U8035 (N_8035,N_3903,N_5101);
nand U8036 (N_8036,N_5326,N_5895);
and U8037 (N_8037,N_4343,N_4800);
nand U8038 (N_8038,N_4460,N_5539);
nor U8039 (N_8039,N_3716,N_3406);
nand U8040 (N_8040,N_4709,N_5867);
and U8041 (N_8041,N_5336,N_5796);
or U8042 (N_8042,N_3554,N_5080);
and U8043 (N_8043,N_4174,N_4651);
or U8044 (N_8044,N_3613,N_4348);
nor U8045 (N_8045,N_4272,N_5323);
and U8046 (N_8046,N_3534,N_5516);
nor U8047 (N_8047,N_3657,N_3885);
nand U8048 (N_8048,N_4294,N_3364);
nand U8049 (N_8049,N_3065,N_3295);
or U8050 (N_8050,N_5984,N_4712);
or U8051 (N_8051,N_5277,N_4068);
nand U8052 (N_8052,N_5983,N_5429);
or U8053 (N_8053,N_4288,N_5687);
nor U8054 (N_8054,N_4968,N_4705);
and U8055 (N_8055,N_3042,N_4184);
nand U8056 (N_8056,N_5869,N_3344);
nand U8057 (N_8057,N_5819,N_4544);
and U8058 (N_8058,N_3014,N_5318);
or U8059 (N_8059,N_4714,N_4101);
nand U8060 (N_8060,N_4694,N_5092);
nand U8061 (N_8061,N_3735,N_3339);
or U8062 (N_8062,N_3790,N_5379);
nor U8063 (N_8063,N_3120,N_5007);
nand U8064 (N_8064,N_3132,N_3698);
nand U8065 (N_8065,N_3447,N_3317);
or U8066 (N_8066,N_5654,N_5222);
nor U8067 (N_8067,N_4373,N_4560);
xnor U8068 (N_8068,N_3332,N_3586);
or U8069 (N_8069,N_5409,N_5604);
or U8070 (N_8070,N_5427,N_5468);
nor U8071 (N_8071,N_4839,N_4335);
nor U8072 (N_8072,N_4300,N_5938);
xnor U8073 (N_8073,N_3890,N_3090);
or U8074 (N_8074,N_4427,N_3612);
and U8075 (N_8075,N_5166,N_3296);
and U8076 (N_8076,N_4917,N_5195);
nand U8077 (N_8077,N_3706,N_3971);
nor U8078 (N_8078,N_3959,N_3415);
and U8079 (N_8079,N_5781,N_3458);
nand U8080 (N_8080,N_4088,N_5075);
nor U8081 (N_8081,N_3053,N_3947);
or U8082 (N_8082,N_4122,N_5691);
or U8083 (N_8083,N_5036,N_5548);
or U8084 (N_8084,N_4206,N_5425);
nand U8085 (N_8085,N_3327,N_4723);
and U8086 (N_8086,N_4362,N_4692);
and U8087 (N_8087,N_5395,N_4405);
or U8088 (N_8088,N_4687,N_3339);
and U8089 (N_8089,N_3079,N_4734);
and U8090 (N_8090,N_4159,N_4956);
and U8091 (N_8091,N_4164,N_5934);
or U8092 (N_8092,N_4373,N_3913);
nor U8093 (N_8093,N_4050,N_5936);
and U8094 (N_8094,N_4700,N_3137);
nor U8095 (N_8095,N_4289,N_4547);
nor U8096 (N_8096,N_4398,N_5391);
and U8097 (N_8097,N_3207,N_5154);
nor U8098 (N_8098,N_4158,N_4782);
nand U8099 (N_8099,N_5407,N_4738);
or U8100 (N_8100,N_3557,N_4160);
or U8101 (N_8101,N_5437,N_3743);
or U8102 (N_8102,N_5326,N_3913);
nor U8103 (N_8103,N_4445,N_3710);
nor U8104 (N_8104,N_3226,N_5973);
nor U8105 (N_8105,N_4525,N_3993);
and U8106 (N_8106,N_3108,N_5579);
or U8107 (N_8107,N_3514,N_4812);
nand U8108 (N_8108,N_4874,N_4424);
or U8109 (N_8109,N_5664,N_3591);
nor U8110 (N_8110,N_3772,N_5790);
or U8111 (N_8111,N_5850,N_5790);
or U8112 (N_8112,N_5643,N_5806);
and U8113 (N_8113,N_5898,N_5932);
or U8114 (N_8114,N_4182,N_3126);
nor U8115 (N_8115,N_5087,N_3707);
nor U8116 (N_8116,N_5025,N_4112);
and U8117 (N_8117,N_5043,N_4598);
nand U8118 (N_8118,N_3704,N_5718);
nor U8119 (N_8119,N_4014,N_4200);
and U8120 (N_8120,N_5715,N_5621);
and U8121 (N_8121,N_3022,N_3415);
and U8122 (N_8122,N_4982,N_4870);
and U8123 (N_8123,N_5134,N_5848);
and U8124 (N_8124,N_4454,N_3042);
or U8125 (N_8125,N_5565,N_3886);
nor U8126 (N_8126,N_3830,N_4149);
nor U8127 (N_8127,N_5020,N_5337);
and U8128 (N_8128,N_3715,N_5917);
xor U8129 (N_8129,N_3401,N_5272);
xor U8130 (N_8130,N_4027,N_3030);
nor U8131 (N_8131,N_4855,N_5864);
nor U8132 (N_8132,N_4683,N_4440);
nor U8133 (N_8133,N_3551,N_5428);
nand U8134 (N_8134,N_4730,N_5499);
nand U8135 (N_8135,N_5441,N_4729);
nor U8136 (N_8136,N_5209,N_4260);
nor U8137 (N_8137,N_4374,N_3832);
or U8138 (N_8138,N_5818,N_4579);
nand U8139 (N_8139,N_3752,N_4128);
or U8140 (N_8140,N_5145,N_5569);
and U8141 (N_8141,N_4160,N_5186);
xnor U8142 (N_8142,N_3922,N_3769);
or U8143 (N_8143,N_4198,N_3252);
nand U8144 (N_8144,N_3002,N_5644);
nand U8145 (N_8145,N_3934,N_5401);
or U8146 (N_8146,N_4921,N_4550);
nor U8147 (N_8147,N_4727,N_3782);
or U8148 (N_8148,N_4331,N_5263);
or U8149 (N_8149,N_3803,N_5251);
or U8150 (N_8150,N_5397,N_4260);
nand U8151 (N_8151,N_5952,N_5740);
and U8152 (N_8152,N_4622,N_3091);
nand U8153 (N_8153,N_5707,N_3398);
nor U8154 (N_8154,N_5419,N_3034);
xnor U8155 (N_8155,N_3312,N_3225);
nor U8156 (N_8156,N_3941,N_4978);
or U8157 (N_8157,N_4301,N_5840);
and U8158 (N_8158,N_5338,N_5410);
nor U8159 (N_8159,N_3968,N_3128);
or U8160 (N_8160,N_4008,N_5762);
or U8161 (N_8161,N_5928,N_5861);
or U8162 (N_8162,N_4134,N_5843);
nor U8163 (N_8163,N_3826,N_3654);
nand U8164 (N_8164,N_3495,N_5066);
nand U8165 (N_8165,N_4905,N_5878);
nor U8166 (N_8166,N_4760,N_4355);
or U8167 (N_8167,N_5270,N_4217);
nand U8168 (N_8168,N_5294,N_5304);
nand U8169 (N_8169,N_4938,N_5357);
nor U8170 (N_8170,N_4361,N_5020);
nor U8171 (N_8171,N_5095,N_5391);
and U8172 (N_8172,N_4929,N_3963);
nor U8173 (N_8173,N_4913,N_3515);
or U8174 (N_8174,N_3711,N_5483);
nor U8175 (N_8175,N_3164,N_5750);
or U8176 (N_8176,N_3726,N_5226);
nor U8177 (N_8177,N_4062,N_3639);
nor U8178 (N_8178,N_5199,N_5886);
nor U8179 (N_8179,N_4607,N_5014);
nand U8180 (N_8180,N_5955,N_5536);
nand U8181 (N_8181,N_4260,N_3455);
and U8182 (N_8182,N_5048,N_4473);
nor U8183 (N_8183,N_5849,N_4162);
or U8184 (N_8184,N_5849,N_5785);
nor U8185 (N_8185,N_5757,N_4147);
nand U8186 (N_8186,N_5841,N_3050);
or U8187 (N_8187,N_5628,N_3526);
or U8188 (N_8188,N_5107,N_5469);
and U8189 (N_8189,N_3786,N_4852);
nand U8190 (N_8190,N_4528,N_5151);
nor U8191 (N_8191,N_3135,N_5464);
nand U8192 (N_8192,N_4444,N_3755);
nor U8193 (N_8193,N_4700,N_3017);
or U8194 (N_8194,N_4055,N_3822);
and U8195 (N_8195,N_3946,N_5936);
nor U8196 (N_8196,N_4852,N_5134);
nand U8197 (N_8197,N_3609,N_4498);
or U8198 (N_8198,N_5357,N_4467);
nor U8199 (N_8199,N_3657,N_4573);
and U8200 (N_8200,N_3319,N_3688);
or U8201 (N_8201,N_3928,N_4767);
and U8202 (N_8202,N_3314,N_3374);
nand U8203 (N_8203,N_5261,N_4431);
nand U8204 (N_8204,N_5835,N_5067);
and U8205 (N_8205,N_4901,N_5095);
and U8206 (N_8206,N_4979,N_4164);
or U8207 (N_8207,N_5168,N_4037);
nor U8208 (N_8208,N_3256,N_4026);
or U8209 (N_8209,N_5758,N_4208);
or U8210 (N_8210,N_5998,N_4736);
and U8211 (N_8211,N_5749,N_4337);
xor U8212 (N_8212,N_4528,N_4943);
nand U8213 (N_8213,N_5438,N_5115);
nor U8214 (N_8214,N_4537,N_4445);
and U8215 (N_8215,N_4967,N_3951);
nand U8216 (N_8216,N_5207,N_5862);
nor U8217 (N_8217,N_3059,N_3397);
or U8218 (N_8218,N_3165,N_5550);
nor U8219 (N_8219,N_4173,N_4418);
nor U8220 (N_8220,N_3019,N_3741);
nand U8221 (N_8221,N_5175,N_4851);
nand U8222 (N_8222,N_4673,N_3749);
nor U8223 (N_8223,N_4819,N_5998);
or U8224 (N_8224,N_4552,N_3303);
or U8225 (N_8225,N_5574,N_5361);
nand U8226 (N_8226,N_3386,N_5138);
nor U8227 (N_8227,N_3727,N_4642);
and U8228 (N_8228,N_5470,N_4724);
nand U8229 (N_8229,N_4536,N_4777);
and U8230 (N_8230,N_3722,N_4912);
nor U8231 (N_8231,N_5767,N_3868);
or U8232 (N_8232,N_3769,N_4759);
and U8233 (N_8233,N_3821,N_3341);
and U8234 (N_8234,N_4704,N_4766);
nand U8235 (N_8235,N_5655,N_4941);
nand U8236 (N_8236,N_3131,N_4018);
nand U8237 (N_8237,N_4934,N_3885);
nand U8238 (N_8238,N_4425,N_3635);
nor U8239 (N_8239,N_3301,N_5526);
or U8240 (N_8240,N_3348,N_5265);
and U8241 (N_8241,N_3135,N_3272);
and U8242 (N_8242,N_3943,N_5702);
nand U8243 (N_8243,N_4576,N_5519);
nor U8244 (N_8244,N_5009,N_4566);
and U8245 (N_8245,N_5258,N_4427);
nor U8246 (N_8246,N_5076,N_3956);
and U8247 (N_8247,N_3763,N_5568);
nor U8248 (N_8248,N_4139,N_3913);
or U8249 (N_8249,N_4848,N_3703);
or U8250 (N_8250,N_5291,N_4620);
or U8251 (N_8251,N_5834,N_3531);
nand U8252 (N_8252,N_3566,N_4574);
or U8253 (N_8253,N_3005,N_5169);
or U8254 (N_8254,N_4212,N_5873);
and U8255 (N_8255,N_3337,N_3807);
and U8256 (N_8256,N_4558,N_3518);
nor U8257 (N_8257,N_3086,N_4785);
nor U8258 (N_8258,N_4936,N_3768);
nor U8259 (N_8259,N_5922,N_4637);
or U8260 (N_8260,N_5614,N_5386);
nor U8261 (N_8261,N_5041,N_4614);
xnor U8262 (N_8262,N_4454,N_4270);
or U8263 (N_8263,N_4295,N_3368);
nand U8264 (N_8264,N_3260,N_4957);
and U8265 (N_8265,N_3673,N_3700);
and U8266 (N_8266,N_5708,N_4610);
nand U8267 (N_8267,N_3945,N_4323);
and U8268 (N_8268,N_3044,N_3847);
or U8269 (N_8269,N_4835,N_4325);
nand U8270 (N_8270,N_3859,N_3146);
xor U8271 (N_8271,N_3815,N_5124);
or U8272 (N_8272,N_3433,N_5521);
and U8273 (N_8273,N_3639,N_4988);
nor U8274 (N_8274,N_3019,N_4166);
or U8275 (N_8275,N_5673,N_3215);
and U8276 (N_8276,N_3766,N_5409);
nor U8277 (N_8277,N_3875,N_4217);
nor U8278 (N_8278,N_5506,N_3778);
and U8279 (N_8279,N_5329,N_5722);
and U8280 (N_8280,N_5546,N_3642);
and U8281 (N_8281,N_4610,N_4724);
nand U8282 (N_8282,N_3413,N_4639);
nor U8283 (N_8283,N_5610,N_3712);
nor U8284 (N_8284,N_5168,N_4542);
and U8285 (N_8285,N_4776,N_4285);
nand U8286 (N_8286,N_3583,N_4359);
or U8287 (N_8287,N_5932,N_3405);
or U8288 (N_8288,N_5133,N_5006);
and U8289 (N_8289,N_3010,N_4218);
nand U8290 (N_8290,N_3272,N_4627);
or U8291 (N_8291,N_4655,N_3765);
nand U8292 (N_8292,N_5505,N_5665);
nand U8293 (N_8293,N_3079,N_3893);
nand U8294 (N_8294,N_5251,N_4359);
nor U8295 (N_8295,N_3267,N_4454);
or U8296 (N_8296,N_4318,N_3570);
nor U8297 (N_8297,N_5059,N_4305);
or U8298 (N_8298,N_4395,N_4592);
or U8299 (N_8299,N_5588,N_5860);
nand U8300 (N_8300,N_3929,N_4255);
nand U8301 (N_8301,N_3764,N_3070);
and U8302 (N_8302,N_3985,N_3712);
or U8303 (N_8303,N_5207,N_3202);
and U8304 (N_8304,N_4038,N_5359);
nor U8305 (N_8305,N_3545,N_4454);
nor U8306 (N_8306,N_4021,N_3788);
nor U8307 (N_8307,N_4364,N_5214);
nor U8308 (N_8308,N_4587,N_4240);
or U8309 (N_8309,N_3424,N_4330);
nor U8310 (N_8310,N_4022,N_3170);
and U8311 (N_8311,N_3366,N_4449);
nor U8312 (N_8312,N_3213,N_3991);
and U8313 (N_8313,N_4112,N_5231);
nand U8314 (N_8314,N_3344,N_5437);
or U8315 (N_8315,N_4728,N_4680);
nor U8316 (N_8316,N_3664,N_4873);
and U8317 (N_8317,N_4515,N_5462);
xnor U8318 (N_8318,N_3531,N_5224);
nand U8319 (N_8319,N_4286,N_5010);
and U8320 (N_8320,N_4253,N_5075);
nor U8321 (N_8321,N_3495,N_4937);
nor U8322 (N_8322,N_3618,N_5464);
and U8323 (N_8323,N_4560,N_3850);
nor U8324 (N_8324,N_4320,N_4721);
or U8325 (N_8325,N_4528,N_3074);
or U8326 (N_8326,N_5028,N_3108);
nor U8327 (N_8327,N_4028,N_4388);
nor U8328 (N_8328,N_4840,N_4992);
nor U8329 (N_8329,N_5489,N_3888);
nand U8330 (N_8330,N_4215,N_4649);
xor U8331 (N_8331,N_5702,N_3296);
and U8332 (N_8332,N_3717,N_5971);
nor U8333 (N_8333,N_4558,N_4956);
or U8334 (N_8334,N_4198,N_5253);
nor U8335 (N_8335,N_5086,N_4227);
nor U8336 (N_8336,N_3130,N_3748);
nand U8337 (N_8337,N_4401,N_4242);
xor U8338 (N_8338,N_3601,N_4727);
and U8339 (N_8339,N_4283,N_5703);
and U8340 (N_8340,N_3180,N_5845);
nand U8341 (N_8341,N_4674,N_3891);
and U8342 (N_8342,N_4171,N_5061);
nor U8343 (N_8343,N_3042,N_3063);
nand U8344 (N_8344,N_3246,N_5400);
nand U8345 (N_8345,N_4234,N_4827);
nor U8346 (N_8346,N_5705,N_4671);
or U8347 (N_8347,N_3092,N_3266);
nor U8348 (N_8348,N_5968,N_5325);
nand U8349 (N_8349,N_3845,N_4093);
nand U8350 (N_8350,N_5360,N_3192);
and U8351 (N_8351,N_4918,N_5345);
or U8352 (N_8352,N_5070,N_5789);
and U8353 (N_8353,N_5059,N_3592);
nor U8354 (N_8354,N_4958,N_5088);
or U8355 (N_8355,N_4238,N_4811);
or U8356 (N_8356,N_4844,N_3011);
nor U8357 (N_8357,N_3325,N_5048);
nor U8358 (N_8358,N_3143,N_5248);
xnor U8359 (N_8359,N_4804,N_4979);
nor U8360 (N_8360,N_4084,N_4631);
nor U8361 (N_8361,N_4611,N_3479);
and U8362 (N_8362,N_3487,N_3158);
nor U8363 (N_8363,N_3749,N_3652);
nor U8364 (N_8364,N_5305,N_4996);
or U8365 (N_8365,N_5186,N_5255);
and U8366 (N_8366,N_3587,N_4719);
nor U8367 (N_8367,N_5495,N_5588);
and U8368 (N_8368,N_4528,N_4822);
nor U8369 (N_8369,N_3399,N_5454);
xnor U8370 (N_8370,N_5045,N_3850);
and U8371 (N_8371,N_4252,N_3862);
or U8372 (N_8372,N_4257,N_3473);
nor U8373 (N_8373,N_3564,N_3842);
or U8374 (N_8374,N_4692,N_5593);
or U8375 (N_8375,N_4626,N_5817);
nand U8376 (N_8376,N_4249,N_5452);
and U8377 (N_8377,N_4547,N_4379);
and U8378 (N_8378,N_3114,N_4079);
xnor U8379 (N_8379,N_5974,N_4267);
nand U8380 (N_8380,N_4609,N_3005);
and U8381 (N_8381,N_4702,N_5901);
xnor U8382 (N_8382,N_4904,N_4993);
nor U8383 (N_8383,N_5133,N_3432);
or U8384 (N_8384,N_3957,N_4726);
nand U8385 (N_8385,N_4317,N_5500);
nand U8386 (N_8386,N_3616,N_5008);
or U8387 (N_8387,N_5204,N_4224);
and U8388 (N_8388,N_4149,N_4202);
or U8389 (N_8389,N_3162,N_3007);
nand U8390 (N_8390,N_3232,N_4748);
or U8391 (N_8391,N_4260,N_4309);
nand U8392 (N_8392,N_5757,N_3683);
and U8393 (N_8393,N_5042,N_5998);
nand U8394 (N_8394,N_5190,N_4189);
nand U8395 (N_8395,N_5846,N_5571);
and U8396 (N_8396,N_5732,N_4047);
or U8397 (N_8397,N_4670,N_4040);
nand U8398 (N_8398,N_4665,N_4709);
or U8399 (N_8399,N_4094,N_3762);
nor U8400 (N_8400,N_3196,N_4684);
nor U8401 (N_8401,N_3966,N_4854);
and U8402 (N_8402,N_4584,N_3677);
xor U8403 (N_8403,N_5502,N_5902);
or U8404 (N_8404,N_3606,N_4354);
nand U8405 (N_8405,N_4728,N_3395);
and U8406 (N_8406,N_4757,N_5100);
nand U8407 (N_8407,N_5863,N_3467);
or U8408 (N_8408,N_4975,N_3966);
and U8409 (N_8409,N_5580,N_3478);
or U8410 (N_8410,N_4685,N_4393);
nor U8411 (N_8411,N_4598,N_4829);
nand U8412 (N_8412,N_4952,N_4077);
nand U8413 (N_8413,N_3397,N_5623);
or U8414 (N_8414,N_5793,N_5678);
and U8415 (N_8415,N_4098,N_3821);
and U8416 (N_8416,N_3745,N_4723);
or U8417 (N_8417,N_5222,N_4735);
nand U8418 (N_8418,N_4915,N_4242);
nand U8419 (N_8419,N_4941,N_4995);
nor U8420 (N_8420,N_5908,N_3858);
nand U8421 (N_8421,N_3647,N_4051);
and U8422 (N_8422,N_5728,N_4673);
nand U8423 (N_8423,N_4363,N_3791);
nand U8424 (N_8424,N_3566,N_3452);
nand U8425 (N_8425,N_3005,N_5890);
or U8426 (N_8426,N_3058,N_3175);
or U8427 (N_8427,N_3712,N_3232);
or U8428 (N_8428,N_5260,N_4487);
and U8429 (N_8429,N_5050,N_4648);
nand U8430 (N_8430,N_5428,N_3342);
and U8431 (N_8431,N_5794,N_4763);
or U8432 (N_8432,N_4744,N_4708);
or U8433 (N_8433,N_5972,N_5313);
nor U8434 (N_8434,N_5036,N_3403);
nor U8435 (N_8435,N_3341,N_5003);
nand U8436 (N_8436,N_3344,N_4316);
or U8437 (N_8437,N_3639,N_3575);
nor U8438 (N_8438,N_3087,N_5562);
xor U8439 (N_8439,N_3603,N_5859);
nand U8440 (N_8440,N_3574,N_5508);
and U8441 (N_8441,N_3784,N_5860);
nand U8442 (N_8442,N_5475,N_5938);
nand U8443 (N_8443,N_5178,N_3793);
nand U8444 (N_8444,N_4552,N_3273);
and U8445 (N_8445,N_5358,N_4110);
nor U8446 (N_8446,N_5546,N_5719);
and U8447 (N_8447,N_3907,N_3777);
or U8448 (N_8448,N_5070,N_5900);
or U8449 (N_8449,N_4736,N_4227);
nor U8450 (N_8450,N_3947,N_3393);
or U8451 (N_8451,N_3190,N_3579);
nor U8452 (N_8452,N_3331,N_3552);
nand U8453 (N_8453,N_3326,N_4053);
nand U8454 (N_8454,N_5607,N_4555);
nor U8455 (N_8455,N_3219,N_4047);
nand U8456 (N_8456,N_4539,N_4153);
or U8457 (N_8457,N_5787,N_4805);
nor U8458 (N_8458,N_3639,N_4952);
nor U8459 (N_8459,N_3929,N_3647);
nor U8460 (N_8460,N_5702,N_4594);
nor U8461 (N_8461,N_4045,N_5311);
or U8462 (N_8462,N_4455,N_3064);
nand U8463 (N_8463,N_5178,N_3553);
nor U8464 (N_8464,N_4929,N_3490);
and U8465 (N_8465,N_4914,N_3376);
or U8466 (N_8466,N_4558,N_4695);
nand U8467 (N_8467,N_5250,N_5339);
or U8468 (N_8468,N_3336,N_4472);
or U8469 (N_8469,N_4036,N_4676);
or U8470 (N_8470,N_5398,N_4310);
and U8471 (N_8471,N_5808,N_4356);
and U8472 (N_8472,N_3731,N_3517);
nand U8473 (N_8473,N_5356,N_3628);
nand U8474 (N_8474,N_5811,N_4884);
nor U8475 (N_8475,N_5056,N_5311);
nand U8476 (N_8476,N_3823,N_5700);
nand U8477 (N_8477,N_3300,N_5543);
nand U8478 (N_8478,N_3306,N_3022);
nand U8479 (N_8479,N_4874,N_3155);
nand U8480 (N_8480,N_5465,N_4398);
nand U8481 (N_8481,N_4124,N_5130);
xnor U8482 (N_8482,N_3490,N_5092);
nor U8483 (N_8483,N_3879,N_4202);
and U8484 (N_8484,N_4697,N_3208);
or U8485 (N_8485,N_4106,N_3068);
or U8486 (N_8486,N_4331,N_5638);
and U8487 (N_8487,N_5001,N_5933);
nand U8488 (N_8488,N_3727,N_4038);
and U8489 (N_8489,N_4091,N_3656);
nand U8490 (N_8490,N_4821,N_3257);
nand U8491 (N_8491,N_5665,N_5729);
and U8492 (N_8492,N_3829,N_3860);
and U8493 (N_8493,N_5731,N_5959);
or U8494 (N_8494,N_5158,N_5116);
nor U8495 (N_8495,N_4247,N_5811);
and U8496 (N_8496,N_3291,N_3594);
nor U8497 (N_8497,N_5383,N_5047);
and U8498 (N_8498,N_3000,N_5449);
or U8499 (N_8499,N_3852,N_4797);
or U8500 (N_8500,N_4429,N_5018);
or U8501 (N_8501,N_4625,N_5824);
xnor U8502 (N_8502,N_4852,N_3902);
nor U8503 (N_8503,N_4493,N_3441);
or U8504 (N_8504,N_5464,N_3032);
nor U8505 (N_8505,N_4893,N_5096);
or U8506 (N_8506,N_4763,N_4164);
nand U8507 (N_8507,N_3820,N_5143);
nor U8508 (N_8508,N_3858,N_4736);
and U8509 (N_8509,N_3176,N_4915);
or U8510 (N_8510,N_4945,N_5062);
nand U8511 (N_8511,N_5935,N_3423);
and U8512 (N_8512,N_4734,N_5112);
or U8513 (N_8513,N_4377,N_4522);
nor U8514 (N_8514,N_4052,N_5388);
or U8515 (N_8515,N_5607,N_4458);
nor U8516 (N_8516,N_5485,N_5995);
and U8517 (N_8517,N_3374,N_3251);
nand U8518 (N_8518,N_3001,N_3700);
nor U8519 (N_8519,N_3404,N_5103);
nand U8520 (N_8520,N_4376,N_5658);
nor U8521 (N_8521,N_3736,N_5722);
nor U8522 (N_8522,N_5859,N_3782);
nor U8523 (N_8523,N_3614,N_4972);
and U8524 (N_8524,N_3564,N_4157);
nor U8525 (N_8525,N_3786,N_5106);
and U8526 (N_8526,N_5132,N_4557);
nor U8527 (N_8527,N_4663,N_4745);
nand U8528 (N_8528,N_3489,N_3018);
or U8529 (N_8529,N_4605,N_3807);
or U8530 (N_8530,N_5658,N_3300);
nor U8531 (N_8531,N_5132,N_5397);
or U8532 (N_8532,N_5196,N_5915);
and U8533 (N_8533,N_4803,N_4540);
nand U8534 (N_8534,N_4249,N_3956);
nand U8535 (N_8535,N_5265,N_3280);
and U8536 (N_8536,N_4637,N_5375);
or U8537 (N_8537,N_3440,N_3828);
or U8538 (N_8538,N_3947,N_5699);
and U8539 (N_8539,N_4874,N_4083);
or U8540 (N_8540,N_5366,N_5753);
and U8541 (N_8541,N_4934,N_4417);
or U8542 (N_8542,N_3257,N_4485);
or U8543 (N_8543,N_4232,N_4510);
nand U8544 (N_8544,N_3641,N_5493);
and U8545 (N_8545,N_3911,N_5757);
and U8546 (N_8546,N_4948,N_5762);
nand U8547 (N_8547,N_3836,N_5529);
or U8548 (N_8548,N_3407,N_3947);
and U8549 (N_8549,N_3753,N_4430);
xnor U8550 (N_8550,N_5499,N_3830);
nor U8551 (N_8551,N_5180,N_5311);
nand U8552 (N_8552,N_4216,N_4913);
and U8553 (N_8553,N_4624,N_3364);
nor U8554 (N_8554,N_3261,N_5394);
or U8555 (N_8555,N_3499,N_4130);
nor U8556 (N_8556,N_3599,N_3836);
nand U8557 (N_8557,N_3232,N_3244);
or U8558 (N_8558,N_5371,N_3076);
or U8559 (N_8559,N_3008,N_3735);
or U8560 (N_8560,N_3923,N_4244);
nor U8561 (N_8561,N_3285,N_4649);
or U8562 (N_8562,N_3793,N_5013);
and U8563 (N_8563,N_5831,N_4855);
nor U8564 (N_8564,N_4463,N_3854);
nand U8565 (N_8565,N_4379,N_3279);
nor U8566 (N_8566,N_3227,N_3188);
or U8567 (N_8567,N_3559,N_3739);
nor U8568 (N_8568,N_4082,N_4530);
and U8569 (N_8569,N_5365,N_5033);
nand U8570 (N_8570,N_3723,N_4656);
nor U8571 (N_8571,N_3648,N_4320);
or U8572 (N_8572,N_3956,N_4581);
nor U8573 (N_8573,N_4939,N_5335);
nor U8574 (N_8574,N_5785,N_5204);
or U8575 (N_8575,N_3533,N_3216);
and U8576 (N_8576,N_4350,N_5622);
nor U8577 (N_8577,N_3306,N_3729);
and U8578 (N_8578,N_3225,N_5468);
or U8579 (N_8579,N_5138,N_3840);
and U8580 (N_8580,N_3469,N_3911);
or U8581 (N_8581,N_5719,N_4747);
or U8582 (N_8582,N_4632,N_4832);
nor U8583 (N_8583,N_3325,N_4501);
nor U8584 (N_8584,N_5297,N_5898);
and U8585 (N_8585,N_4584,N_5726);
and U8586 (N_8586,N_4265,N_4610);
xnor U8587 (N_8587,N_3151,N_4012);
nor U8588 (N_8588,N_3264,N_3744);
and U8589 (N_8589,N_3353,N_3261);
or U8590 (N_8590,N_3001,N_4302);
nor U8591 (N_8591,N_3493,N_3716);
and U8592 (N_8592,N_4939,N_3431);
nor U8593 (N_8593,N_3314,N_5677);
and U8594 (N_8594,N_5632,N_4601);
or U8595 (N_8595,N_5246,N_5796);
nand U8596 (N_8596,N_3728,N_5107);
and U8597 (N_8597,N_4980,N_4549);
and U8598 (N_8598,N_5721,N_4649);
nor U8599 (N_8599,N_4838,N_4014);
nor U8600 (N_8600,N_4670,N_4039);
nand U8601 (N_8601,N_5846,N_4174);
or U8602 (N_8602,N_5258,N_5389);
or U8603 (N_8603,N_3617,N_3282);
nor U8604 (N_8604,N_3144,N_5334);
nand U8605 (N_8605,N_4901,N_4902);
nand U8606 (N_8606,N_5739,N_5758);
nand U8607 (N_8607,N_4266,N_3308);
and U8608 (N_8608,N_4061,N_3322);
or U8609 (N_8609,N_4932,N_5603);
nand U8610 (N_8610,N_5013,N_5820);
nor U8611 (N_8611,N_3379,N_4619);
nor U8612 (N_8612,N_4578,N_3240);
nor U8613 (N_8613,N_3072,N_3826);
or U8614 (N_8614,N_5940,N_4965);
nor U8615 (N_8615,N_3454,N_4585);
or U8616 (N_8616,N_3089,N_5537);
nor U8617 (N_8617,N_4313,N_3904);
nor U8618 (N_8618,N_3816,N_4093);
and U8619 (N_8619,N_4664,N_3217);
nand U8620 (N_8620,N_3326,N_5424);
nor U8621 (N_8621,N_3033,N_4694);
and U8622 (N_8622,N_5912,N_3128);
or U8623 (N_8623,N_4330,N_3396);
or U8624 (N_8624,N_5695,N_3111);
nor U8625 (N_8625,N_4272,N_5535);
or U8626 (N_8626,N_3094,N_3903);
or U8627 (N_8627,N_5248,N_5989);
or U8628 (N_8628,N_5905,N_5355);
or U8629 (N_8629,N_3214,N_5156);
or U8630 (N_8630,N_5732,N_4389);
or U8631 (N_8631,N_5313,N_4648);
nand U8632 (N_8632,N_5995,N_5553);
or U8633 (N_8633,N_4427,N_4481);
nor U8634 (N_8634,N_4140,N_5391);
or U8635 (N_8635,N_3053,N_3546);
nor U8636 (N_8636,N_4862,N_5946);
and U8637 (N_8637,N_5939,N_3093);
and U8638 (N_8638,N_3252,N_5952);
and U8639 (N_8639,N_3383,N_5742);
nand U8640 (N_8640,N_5244,N_4125);
or U8641 (N_8641,N_5048,N_4945);
nand U8642 (N_8642,N_5153,N_3682);
nand U8643 (N_8643,N_5772,N_5458);
nor U8644 (N_8644,N_4191,N_5772);
or U8645 (N_8645,N_3854,N_3892);
and U8646 (N_8646,N_3415,N_5511);
nand U8647 (N_8647,N_3012,N_3310);
xor U8648 (N_8648,N_4183,N_5029);
or U8649 (N_8649,N_3630,N_5552);
and U8650 (N_8650,N_4296,N_4867);
or U8651 (N_8651,N_4270,N_5975);
nand U8652 (N_8652,N_3490,N_5127);
and U8653 (N_8653,N_3784,N_5767);
nor U8654 (N_8654,N_5184,N_3917);
and U8655 (N_8655,N_3110,N_3197);
and U8656 (N_8656,N_4474,N_5375);
nand U8657 (N_8657,N_4315,N_4844);
and U8658 (N_8658,N_5661,N_4650);
nand U8659 (N_8659,N_4233,N_4950);
nor U8660 (N_8660,N_5312,N_3515);
nand U8661 (N_8661,N_3634,N_3162);
or U8662 (N_8662,N_3713,N_4963);
and U8663 (N_8663,N_5700,N_3104);
nand U8664 (N_8664,N_4585,N_5886);
nand U8665 (N_8665,N_3943,N_4718);
and U8666 (N_8666,N_4495,N_5740);
or U8667 (N_8667,N_5722,N_5377);
nand U8668 (N_8668,N_3041,N_4804);
or U8669 (N_8669,N_4692,N_5012);
and U8670 (N_8670,N_4532,N_4129);
and U8671 (N_8671,N_5851,N_4278);
nor U8672 (N_8672,N_4877,N_3047);
nand U8673 (N_8673,N_5198,N_4712);
and U8674 (N_8674,N_3565,N_3353);
nor U8675 (N_8675,N_4667,N_3071);
nand U8676 (N_8676,N_5404,N_3348);
nand U8677 (N_8677,N_3640,N_3450);
or U8678 (N_8678,N_4667,N_4860);
nand U8679 (N_8679,N_3083,N_3420);
or U8680 (N_8680,N_4235,N_4682);
nand U8681 (N_8681,N_4716,N_3854);
nor U8682 (N_8682,N_5087,N_3048);
xnor U8683 (N_8683,N_5867,N_4136);
nand U8684 (N_8684,N_3402,N_4875);
or U8685 (N_8685,N_3575,N_3447);
and U8686 (N_8686,N_5285,N_3013);
and U8687 (N_8687,N_4707,N_3467);
nor U8688 (N_8688,N_4884,N_3942);
and U8689 (N_8689,N_3121,N_5713);
nand U8690 (N_8690,N_5323,N_5567);
and U8691 (N_8691,N_5899,N_3773);
nand U8692 (N_8692,N_5761,N_5393);
nand U8693 (N_8693,N_5824,N_5994);
or U8694 (N_8694,N_3100,N_5438);
nor U8695 (N_8695,N_4455,N_5364);
nor U8696 (N_8696,N_4857,N_4027);
nand U8697 (N_8697,N_5358,N_3027);
xor U8698 (N_8698,N_5211,N_5595);
nand U8699 (N_8699,N_5661,N_4536);
or U8700 (N_8700,N_5220,N_5756);
nand U8701 (N_8701,N_4675,N_5388);
nor U8702 (N_8702,N_5418,N_5987);
or U8703 (N_8703,N_5411,N_4712);
and U8704 (N_8704,N_5940,N_4834);
or U8705 (N_8705,N_4920,N_3810);
nor U8706 (N_8706,N_5854,N_3252);
and U8707 (N_8707,N_3459,N_5119);
and U8708 (N_8708,N_4074,N_3991);
nor U8709 (N_8709,N_5888,N_5585);
nor U8710 (N_8710,N_5368,N_5695);
or U8711 (N_8711,N_3930,N_4835);
and U8712 (N_8712,N_3417,N_5001);
or U8713 (N_8713,N_3587,N_4973);
nand U8714 (N_8714,N_3278,N_3654);
or U8715 (N_8715,N_3334,N_4425);
nand U8716 (N_8716,N_4631,N_4777);
nand U8717 (N_8717,N_3638,N_3052);
and U8718 (N_8718,N_5099,N_5070);
and U8719 (N_8719,N_5506,N_4468);
and U8720 (N_8720,N_4416,N_3763);
and U8721 (N_8721,N_5140,N_5275);
nand U8722 (N_8722,N_4589,N_4298);
or U8723 (N_8723,N_5518,N_5558);
nor U8724 (N_8724,N_3725,N_3364);
nor U8725 (N_8725,N_5545,N_5667);
or U8726 (N_8726,N_4811,N_3057);
or U8727 (N_8727,N_4621,N_4140);
or U8728 (N_8728,N_5599,N_4167);
or U8729 (N_8729,N_4852,N_5111);
and U8730 (N_8730,N_4013,N_3726);
nand U8731 (N_8731,N_5668,N_3389);
nor U8732 (N_8732,N_4098,N_5131);
or U8733 (N_8733,N_3467,N_3268);
nor U8734 (N_8734,N_5920,N_4082);
nand U8735 (N_8735,N_5124,N_3217);
nand U8736 (N_8736,N_4280,N_4393);
and U8737 (N_8737,N_5247,N_4365);
nand U8738 (N_8738,N_4402,N_4999);
nor U8739 (N_8739,N_3958,N_4768);
and U8740 (N_8740,N_5786,N_4480);
and U8741 (N_8741,N_4573,N_3104);
nand U8742 (N_8742,N_3528,N_5355);
nand U8743 (N_8743,N_5442,N_4961);
nor U8744 (N_8744,N_4548,N_3189);
nand U8745 (N_8745,N_4691,N_3392);
nor U8746 (N_8746,N_5375,N_5209);
nand U8747 (N_8747,N_3361,N_4747);
nor U8748 (N_8748,N_5013,N_4502);
nor U8749 (N_8749,N_5570,N_3881);
or U8750 (N_8750,N_4055,N_3508);
or U8751 (N_8751,N_5438,N_5276);
and U8752 (N_8752,N_3013,N_4361);
and U8753 (N_8753,N_3755,N_4501);
and U8754 (N_8754,N_3517,N_3884);
or U8755 (N_8755,N_5967,N_3293);
nand U8756 (N_8756,N_4582,N_4519);
and U8757 (N_8757,N_5818,N_5477);
nand U8758 (N_8758,N_5569,N_4955);
or U8759 (N_8759,N_4168,N_3060);
or U8760 (N_8760,N_3757,N_5518);
nand U8761 (N_8761,N_5000,N_3506);
nor U8762 (N_8762,N_5985,N_5028);
nor U8763 (N_8763,N_4898,N_3570);
or U8764 (N_8764,N_4738,N_3694);
nor U8765 (N_8765,N_4392,N_5161);
nand U8766 (N_8766,N_5844,N_4369);
and U8767 (N_8767,N_5677,N_3804);
nand U8768 (N_8768,N_3815,N_5618);
nand U8769 (N_8769,N_4145,N_4844);
xnor U8770 (N_8770,N_5889,N_3595);
nor U8771 (N_8771,N_5964,N_4706);
nor U8772 (N_8772,N_4134,N_3392);
nand U8773 (N_8773,N_5639,N_3069);
and U8774 (N_8774,N_5101,N_4957);
or U8775 (N_8775,N_3977,N_5855);
nor U8776 (N_8776,N_5693,N_4312);
nor U8777 (N_8777,N_3792,N_4988);
nand U8778 (N_8778,N_3810,N_4850);
nand U8779 (N_8779,N_5556,N_4054);
nor U8780 (N_8780,N_4639,N_5675);
and U8781 (N_8781,N_3436,N_3245);
nor U8782 (N_8782,N_4117,N_4087);
nor U8783 (N_8783,N_5370,N_5921);
nand U8784 (N_8784,N_4945,N_3786);
or U8785 (N_8785,N_5155,N_3475);
nor U8786 (N_8786,N_5509,N_5289);
and U8787 (N_8787,N_4376,N_3339);
or U8788 (N_8788,N_3608,N_3549);
nand U8789 (N_8789,N_5056,N_5638);
or U8790 (N_8790,N_4405,N_3646);
nand U8791 (N_8791,N_3974,N_5117);
and U8792 (N_8792,N_3500,N_5099);
nor U8793 (N_8793,N_4688,N_3562);
xnor U8794 (N_8794,N_3418,N_3174);
nor U8795 (N_8795,N_5261,N_5179);
nor U8796 (N_8796,N_3159,N_4729);
or U8797 (N_8797,N_3573,N_4690);
and U8798 (N_8798,N_3145,N_3874);
xor U8799 (N_8799,N_5395,N_3565);
and U8800 (N_8800,N_3444,N_4965);
nor U8801 (N_8801,N_5351,N_4996);
nand U8802 (N_8802,N_5782,N_4223);
nand U8803 (N_8803,N_5709,N_5504);
nor U8804 (N_8804,N_3579,N_5983);
xor U8805 (N_8805,N_3947,N_3472);
or U8806 (N_8806,N_5598,N_5960);
and U8807 (N_8807,N_5498,N_4555);
or U8808 (N_8808,N_3701,N_5200);
nor U8809 (N_8809,N_4981,N_3232);
or U8810 (N_8810,N_4828,N_4573);
nor U8811 (N_8811,N_4514,N_3333);
nand U8812 (N_8812,N_3837,N_5617);
nand U8813 (N_8813,N_3956,N_4287);
nor U8814 (N_8814,N_4525,N_5409);
or U8815 (N_8815,N_5501,N_4263);
or U8816 (N_8816,N_4178,N_4861);
or U8817 (N_8817,N_3543,N_5878);
and U8818 (N_8818,N_5019,N_5533);
or U8819 (N_8819,N_5635,N_4790);
nor U8820 (N_8820,N_5719,N_4136);
nor U8821 (N_8821,N_4696,N_5711);
nor U8822 (N_8822,N_3326,N_5445);
nand U8823 (N_8823,N_4492,N_3856);
nand U8824 (N_8824,N_3110,N_4235);
xnor U8825 (N_8825,N_3185,N_4266);
or U8826 (N_8826,N_4848,N_5098);
nand U8827 (N_8827,N_4960,N_4359);
or U8828 (N_8828,N_4469,N_4058);
or U8829 (N_8829,N_4761,N_4335);
and U8830 (N_8830,N_3060,N_3543);
and U8831 (N_8831,N_4269,N_5592);
and U8832 (N_8832,N_4061,N_5488);
nand U8833 (N_8833,N_4426,N_5396);
nor U8834 (N_8834,N_3249,N_3313);
nor U8835 (N_8835,N_4222,N_5680);
nand U8836 (N_8836,N_5160,N_3058);
and U8837 (N_8837,N_4339,N_4176);
nor U8838 (N_8838,N_4567,N_3944);
nor U8839 (N_8839,N_5825,N_5787);
xnor U8840 (N_8840,N_3760,N_4515);
and U8841 (N_8841,N_3640,N_3823);
nor U8842 (N_8842,N_3653,N_3549);
nor U8843 (N_8843,N_3225,N_5517);
nor U8844 (N_8844,N_3544,N_5888);
nand U8845 (N_8845,N_3293,N_3512);
or U8846 (N_8846,N_4032,N_3884);
xor U8847 (N_8847,N_4979,N_5228);
nand U8848 (N_8848,N_5730,N_5024);
nor U8849 (N_8849,N_4637,N_3924);
or U8850 (N_8850,N_4885,N_5162);
nor U8851 (N_8851,N_4845,N_5351);
nor U8852 (N_8852,N_3081,N_3185);
nand U8853 (N_8853,N_3268,N_4976);
or U8854 (N_8854,N_5234,N_5279);
and U8855 (N_8855,N_3753,N_3281);
or U8856 (N_8856,N_4432,N_3695);
or U8857 (N_8857,N_3240,N_5291);
and U8858 (N_8858,N_4591,N_3177);
nand U8859 (N_8859,N_3495,N_3579);
or U8860 (N_8860,N_4374,N_3378);
nor U8861 (N_8861,N_5686,N_4738);
or U8862 (N_8862,N_3269,N_3508);
nor U8863 (N_8863,N_4597,N_3935);
or U8864 (N_8864,N_5335,N_4473);
xor U8865 (N_8865,N_3042,N_4718);
nor U8866 (N_8866,N_4017,N_4282);
nand U8867 (N_8867,N_3895,N_5080);
nor U8868 (N_8868,N_5717,N_4399);
or U8869 (N_8869,N_3702,N_5421);
and U8870 (N_8870,N_3073,N_5248);
nand U8871 (N_8871,N_5187,N_5197);
and U8872 (N_8872,N_3342,N_5991);
nand U8873 (N_8873,N_3035,N_4824);
nor U8874 (N_8874,N_4429,N_4747);
nand U8875 (N_8875,N_5059,N_3766);
and U8876 (N_8876,N_4312,N_3446);
and U8877 (N_8877,N_3514,N_5292);
or U8878 (N_8878,N_3744,N_3875);
and U8879 (N_8879,N_3494,N_3422);
nand U8880 (N_8880,N_3206,N_4124);
nand U8881 (N_8881,N_4496,N_3168);
nand U8882 (N_8882,N_3179,N_5671);
xnor U8883 (N_8883,N_3379,N_4360);
or U8884 (N_8884,N_3890,N_4764);
or U8885 (N_8885,N_4505,N_5522);
nor U8886 (N_8886,N_4018,N_5506);
nor U8887 (N_8887,N_5250,N_5728);
nand U8888 (N_8888,N_5932,N_5503);
or U8889 (N_8889,N_4416,N_3445);
nor U8890 (N_8890,N_4820,N_3923);
xnor U8891 (N_8891,N_3986,N_5183);
and U8892 (N_8892,N_5515,N_5958);
or U8893 (N_8893,N_5624,N_3905);
nor U8894 (N_8894,N_5791,N_4470);
nand U8895 (N_8895,N_4186,N_3751);
nor U8896 (N_8896,N_3435,N_5485);
nand U8897 (N_8897,N_5582,N_5254);
or U8898 (N_8898,N_3629,N_4011);
nor U8899 (N_8899,N_3292,N_5308);
and U8900 (N_8900,N_3855,N_4080);
xnor U8901 (N_8901,N_5818,N_4683);
or U8902 (N_8902,N_4673,N_4722);
nand U8903 (N_8903,N_3415,N_4174);
xnor U8904 (N_8904,N_5946,N_3791);
or U8905 (N_8905,N_4148,N_4460);
nand U8906 (N_8906,N_3938,N_5970);
and U8907 (N_8907,N_4607,N_3627);
or U8908 (N_8908,N_3986,N_3748);
nand U8909 (N_8909,N_5328,N_3202);
or U8910 (N_8910,N_3821,N_3228);
or U8911 (N_8911,N_3778,N_3133);
nor U8912 (N_8912,N_5325,N_3285);
xor U8913 (N_8913,N_4137,N_4673);
xnor U8914 (N_8914,N_5376,N_5442);
or U8915 (N_8915,N_5491,N_5328);
nand U8916 (N_8916,N_4647,N_4690);
xnor U8917 (N_8917,N_4137,N_3470);
nand U8918 (N_8918,N_5311,N_4303);
nor U8919 (N_8919,N_4022,N_3448);
nor U8920 (N_8920,N_5624,N_3976);
nor U8921 (N_8921,N_3589,N_4302);
and U8922 (N_8922,N_5887,N_4742);
and U8923 (N_8923,N_4332,N_3910);
and U8924 (N_8924,N_5970,N_5389);
nand U8925 (N_8925,N_4290,N_4888);
nand U8926 (N_8926,N_4552,N_5854);
nand U8927 (N_8927,N_4403,N_4232);
and U8928 (N_8928,N_4644,N_3781);
and U8929 (N_8929,N_3219,N_3831);
or U8930 (N_8930,N_5971,N_5978);
nand U8931 (N_8931,N_3711,N_4429);
or U8932 (N_8932,N_5955,N_3710);
or U8933 (N_8933,N_4995,N_5065);
and U8934 (N_8934,N_5384,N_5986);
nand U8935 (N_8935,N_4460,N_5123);
or U8936 (N_8936,N_4032,N_4697);
or U8937 (N_8937,N_4459,N_3631);
xnor U8938 (N_8938,N_3359,N_3411);
nor U8939 (N_8939,N_5787,N_4209);
and U8940 (N_8940,N_3103,N_3301);
nor U8941 (N_8941,N_5011,N_5238);
nand U8942 (N_8942,N_4235,N_5422);
nor U8943 (N_8943,N_4863,N_3787);
or U8944 (N_8944,N_5618,N_3912);
and U8945 (N_8945,N_5511,N_4447);
and U8946 (N_8946,N_4778,N_3675);
nor U8947 (N_8947,N_4324,N_3952);
or U8948 (N_8948,N_4417,N_3564);
and U8949 (N_8949,N_3216,N_5549);
and U8950 (N_8950,N_3802,N_3872);
and U8951 (N_8951,N_5092,N_3296);
nor U8952 (N_8952,N_5413,N_3896);
nor U8953 (N_8953,N_4714,N_5202);
nand U8954 (N_8954,N_3312,N_4194);
and U8955 (N_8955,N_5024,N_3940);
or U8956 (N_8956,N_5746,N_3107);
and U8957 (N_8957,N_4597,N_3704);
or U8958 (N_8958,N_5453,N_4510);
nor U8959 (N_8959,N_4169,N_4512);
nand U8960 (N_8960,N_3857,N_5867);
or U8961 (N_8961,N_3195,N_4942);
nand U8962 (N_8962,N_4439,N_3306);
and U8963 (N_8963,N_5190,N_4281);
nor U8964 (N_8964,N_4291,N_3333);
and U8965 (N_8965,N_4289,N_3108);
and U8966 (N_8966,N_3852,N_4306);
nand U8967 (N_8967,N_3345,N_3944);
nor U8968 (N_8968,N_5345,N_5628);
or U8969 (N_8969,N_5298,N_5351);
or U8970 (N_8970,N_5627,N_5405);
nand U8971 (N_8971,N_5949,N_3509);
and U8972 (N_8972,N_4003,N_4802);
or U8973 (N_8973,N_5772,N_5824);
or U8974 (N_8974,N_4005,N_4529);
or U8975 (N_8975,N_4800,N_4911);
or U8976 (N_8976,N_5337,N_4378);
nor U8977 (N_8977,N_3004,N_4381);
or U8978 (N_8978,N_3537,N_5996);
nand U8979 (N_8979,N_5996,N_5311);
and U8980 (N_8980,N_3517,N_5490);
nand U8981 (N_8981,N_4386,N_3320);
and U8982 (N_8982,N_4812,N_3220);
nand U8983 (N_8983,N_5426,N_5564);
nand U8984 (N_8984,N_3835,N_5372);
nor U8985 (N_8985,N_4816,N_4332);
nor U8986 (N_8986,N_3624,N_3687);
nor U8987 (N_8987,N_3002,N_4661);
or U8988 (N_8988,N_5212,N_4889);
nand U8989 (N_8989,N_4683,N_5109);
nor U8990 (N_8990,N_4009,N_5770);
nor U8991 (N_8991,N_4588,N_3978);
and U8992 (N_8992,N_5331,N_5507);
or U8993 (N_8993,N_3016,N_4495);
nand U8994 (N_8994,N_5415,N_5843);
nor U8995 (N_8995,N_4207,N_5556);
or U8996 (N_8996,N_3274,N_5069);
xor U8997 (N_8997,N_5843,N_4350);
nor U8998 (N_8998,N_5268,N_5386);
and U8999 (N_8999,N_5931,N_5207);
and U9000 (N_9000,N_6677,N_7617);
xnor U9001 (N_9001,N_8654,N_6022);
or U9002 (N_9002,N_7542,N_7075);
nand U9003 (N_9003,N_8817,N_6526);
or U9004 (N_9004,N_6553,N_7262);
xnor U9005 (N_9005,N_6953,N_8498);
nor U9006 (N_9006,N_8433,N_7777);
nand U9007 (N_9007,N_8326,N_8823);
nor U9008 (N_9008,N_6619,N_7279);
nand U9009 (N_9009,N_8562,N_8656);
nand U9010 (N_9010,N_8800,N_8329);
or U9011 (N_9011,N_6997,N_7315);
nor U9012 (N_9012,N_8331,N_8455);
nand U9013 (N_9013,N_6719,N_8615);
nand U9014 (N_9014,N_8537,N_6468);
and U9015 (N_9015,N_8001,N_7120);
nor U9016 (N_9016,N_7354,N_7398);
nand U9017 (N_9017,N_6494,N_6636);
and U9018 (N_9018,N_7888,N_7083);
nand U9019 (N_9019,N_8905,N_7108);
and U9020 (N_9020,N_8200,N_8922);
or U9021 (N_9021,N_6752,N_8602);
nand U9022 (N_9022,N_7805,N_7025);
nor U9023 (N_9023,N_6747,N_6753);
nand U9024 (N_9024,N_6174,N_8875);
or U9025 (N_9025,N_6579,N_6888);
or U9026 (N_9026,N_7961,N_8270);
nor U9027 (N_9027,N_8332,N_6709);
and U9028 (N_9028,N_8842,N_8906);
and U9029 (N_9029,N_6640,N_8179);
and U9030 (N_9030,N_8940,N_8581);
or U9031 (N_9031,N_7107,N_7055);
xnor U9032 (N_9032,N_8890,N_6019);
and U9033 (N_9033,N_8567,N_8106);
or U9034 (N_9034,N_6339,N_8677);
or U9035 (N_9035,N_7143,N_6875);
nand U9036 (N_9036,N_6679,N_8802);
and U9037 (N_9037,N_7875,N_8555);
or U9038 (N_9038,N_7010,N_8864);
and U9039 (N_9039,N_6401,N_7548);
nor U9040 (N_9040,N_6728,N_8419);
and U9041 (N_9041,N_7205,N_8969);
nand U9042 (N_9042,N_7463,N_6958);
or U9043 (N_9043,N_7067,N_8724);
and U9044 (N_9044,N_7167,N_7795);
nor U9045 (N_9045,N_7399,N_8160);
and U9046 (N_9046,N_7586,N_8369);
or U9047 (N_9047,N_7868,N_6721);
nor U9048 (N_9048,N_7700,N_8208);
nand U9049 (N_9049,N_8595,N_8682);
and U9050 (N_9050,N_6484,N_7724);
or U9051 (N_9051,N_6147,N_8354);
and U9052 (N_9052,N_8314,N_8895);
nand U9053 (N_9053,N_7639,N_6871);
nor U9054 (N_9054,N_8673,N_6480);
nor U9055 (N_9055,N_7475,N_8281);
nor U9056 (N_9056,N_7421,N_8668);
and U9057 (N_9057,N_6540,N_6437);
nand U9058 (N_9058,N_8630,N_8702);
or U9059 (N_9059,N_8911,N_7782);
and U9060 (N_9060,N_7145,N_6055);
or U9061 (N_9061,N_8097,N_6667);
and U9062 (N_9062,N_8457,N_6221);
and U9063 (N_9063,N_8954,N_7390);
nand U9064 (N_9064,N_6985,N_7349);
nor U9065 (N_9065,N_7892,N_6078);
nor U9066 (N_9066,N_7134,N_7059);
nand U9067 (N_9067,N_6268,N_8356);
or U9068 (N_9068,N_7719,N_7987);
nor U9069 (N_9069,N_7230,N_6510);
nand U9070 (N_9070,N_6968,N_8662);
nand U9071 (N_9071,N_8564,N_7515);
or U9072 (N_9072,N_7984,N_6954);
nand U9073 (N_9073,N_8578,N_7268);
nor U9074 (N_9074,N_6706,N_6511);
or U9075 (N_9075,N_7213,N_6796);
nand U9076 (N_9076,N_6172,N_7871);
nor U9077 (N_9077,N_8177,N_6797);
nor U9078 (N_9078,N_6190,N_8453);
nor U9079 (N_9079,N_7710,N_6546);
and U9080 (N_9080,N_6199,N_7093);
and U9081 (N_9081,N_6737,N_8180);
and U9082 (N_9082,N_8610,N_6804);
nor U9083 (N_9083,N_6854,N_7171);
nand U9084 (N_9084,N_8308,N_6945);
nand U9085 (N_9085,N_6780,N_8254);
or U9086 (N_9086,N_7273,N_7793);
and U9087 (N_9087,N_6328,N_8941);
or U9088 (N_9088,N_6482,N_7540);
or U9089 (N_9089,N_8278,N_8717);
or U9090 (N_9090,N_7085,N_6101);
nor U9091 (N_9091,N_8410,N_7731);
nor U9092 (N_9092,N_7910,N_7543);
or U9093 (N_9093,N_7392,N_6836);
nor U9094 (N_9094,N_7712,N_8653);
and U9095 (N_9095,N_7549,N_7382);
and U9096 (N_9096,N_7507,N_7411);
nor U9097 (N_9097,N_6094,N_6334);
or U9098 (N_9098,N_7842,N_7624);
or U9099 (N_9099,N_8183,N_8402);
and U9100 (N_9100,N_7184,N_8822);
nor U9101 (N_9101,N_7900,N_6966);
or U9102 (N_9102,N_7594,N_6451);
nand U9103 (N_9103,N_8299,N_6273);
or U9104 (N_9104,N_7469,N_6472);
nand U9105 (N_9105,N_6456,N_7080);
nor U9106 (N_9106,N_7658,N_6637);
nand U9107 (N_9107,N_7631,N_8047);
nand U9108 (N_9108,N_8328,N_7448);
nor U9109 (N_9109,N_7996,N_8252);
and U9110 (N_9110,N_7118,N_8833);
and U9111 (N_9111,N_8919,N_7481);
or U9112 (N_9112,N_7921,N_7880);
nand U9113 (N_9113,N_8342,N_8313);
and U9114 (N_9114,N_6378,N_7284);
nand U9115 (N_9115,N_7529,N_6941);
or U9116 (N_9116,N_8704,N_7730);
nand U9117 (N_9117,N_8083,N_8579);
nor U9118 (N_9118,N_6974,N_8709);
or U9119 (N_9119,N_7394,N_7049);
nand U9120 (N_9120,N_8442,N_6869);
nor U9121 (N_9121,N_8789,N_6149);
and U9122 (N_9122,N_7478,N_7445);
or U9123 (N_9123,N_7992,N_6478);
nand U9124 (N_9124,N_6056,N_6322);
or U9125 (N_9125,N_8867,N_7454);
xor U9126 (N_9126,N_8745,N_6403);
nor U9127 (N_9127,N_8845,N_8014);
nand U9128 (N_9128,N_6371,N_6145);
nand U9129 (N_9129,N_7063,N_6369);
or U9130 (N_9130,N_6093,N_6414);
nor U9131 (N_9131,N_8675,N_8752);
nor U9132 (N_9132,N_6028,N_6891);
nand U9133 (N_9133,N_8269,N_7783);
and U9134 (N_9134,N_8257,N_7460);
nor U9135 (N_9135,N_6878,N_8306);
nand U9136 (N_9136,N_7938,N_6042);
or U9137 (N_9137,N_8207,N_6604);
and U9138 (N_9138,N_6315,N_7068);
nor U9139 (N_9139,N_7653,N_8046);
or U9140 (N_9140,N_6711,N_8736);
and U9141 (N_9141,N_6877,N_7416);
or U9142 (N_9142,N_6260,N_7372);
xor U9143 (N_9143,N_8396,N_7287);
nor U9144 (N_9144,N_6845,N_7129);
nand U9145 (N_9145,N_8035,N_8510);
nor U9146 (N_9146,N_8995,N_6560);
nand U9147 (N_9147,N_8855,N_7765);
nor U9148 (N_9148,N_6951,N_7060);
xnor U9149 (N_9149,N_8244,N_8321);
and U9150 (N_9150,N_7571,N_7916);
nor U9151 (N_9151,N_8840,N_7810);
or U9152 (N_9152,N_8617,N_6748);
or U9153 (N_9153,N_7231,N_7796);
nor U9154 (N_9154,N_6184,N_8202);
and U9155 (N_9155,N_7029,N_7749);
nand U9156 (N_9156,N_6206,N_7032);
and U9157 (N_9157,N_8366,N_7491);
or U9158 (N_9158,N_8527,N_7401);
nor U9159 (N_9159,N_6496,N_7590);
and U9160 (N_9160,N_7807,N_8848);
nor U9161 (N_9161,N_6072,N_8378);
or U9162 (N_9162,N_6876,N_7191);
or U9163 (N_9163,N_7747,N_8598);
and U9164 (N_9164,N_6285,N_6499);
and U9165 (N_9165,N_8156,N_7275);
nor U9166 (N_9166,N_7691,N_7189);
nand U9167 (N_9167,N_8074,N_7726);
and U9168 (N_9168,N_8377,N_6799);
nand U9169 (N_9169,N_6517,N_7744);
or U9170 (N_9170,N_8703,N_6960);
nand U9171 (N_9171,N_7260,N_6448);
and U9172 (N_9172,N_7896,N_7277);
or U9173 (N_9173,N_8769,N_7127);
and U9174 (N_9174,N_7226,N_8126);
and U9175 (N_9175,N_8151,N_7434);
or U9176 (N_9176,N_7019,N_8808);
and U9177 (N_9177,N_6251,N_7355);
and U9178 (N_9178,N_8081,N_7022);
or U9179 (N_9179,N_7014,N_6544);
or U9180 (N_9180,N_6734,N_8013);
nor U9181 (N_9181,N_7674,N_7076);
nand U9182 (N_9182,N_7945,N_7114);
or U9183 (N_9183,N_6815,N_7560);
and U9184 (N_9184,N_6107,N_6761);
nand U9185 (N_9185,N_6750,N_6057);
and U9186 (N_9186,N_8871,N_7435);
nor U9187 (N_9187,N_7610,N_7736);
and U9188 (N_9188,N_6427,N_8627);
or U9189 (N_9189,N_7286,N_6702);
xnor U9190 (N_9190,N_7577,N_7099);
and U9191 (N_9191,N_7570,N_6408);
or U9192 (N_9192,N_6185,N_6930);
nand U9193 (N_9193,N_8909,N_6025);
nor U9194 (N_9194,N_7005,N_7418);
nor U9195 (N_9195,N_8549,N_8176);
and U9196 (N_9196,N_7671,N_7288);
or U9197 (N_9197,N_8529,N_6880);
nor U9198 (N_9198,N_6584,N_6811);
nand U9199 (N_9199,N_7211,N_7247);
or U9200 (N_9200,N_6128,N_7637);
and U9201 (N_9201,N_8107,N_6950);
or U9202 (N_9202,N_8137,N_8622);
and U9203 (N_9203,N_6281,N_8633);
and U9204 (N_9204,N_6029,N_8665);
nand U9205 (N_9205,N_8155,N_8372);
or U9206 (N_9206,N_6908,N_7633);
and U9207 (N_9207,N_8394,N_8893);
nor U9208 (N_9208,N_8659,N_7697);
and U9209 (N_9209,N_7026,N_6065);
nor U9210 (N_9210,N_6806,N_6755);
nand U9211 (N_9211,N_7340,N_6017);
and U9212 (N_9212,N_7131,N_6062);
nor U9213 (N_9213,N_6572,N_7879);
nand U9214 (N_9214,N_8818,N_8411);
and U9215 (N_9215,N_8612,N_8978);
and U9216 (N_9216,N_8168,N_7538);
and U9217 (N_9217,N_7696,N_6381);
nor U9218 (N_9218,N_7950,N_7034);
and U9219 (N_9219,N_6547,N_7789);
nor U9220 (N_9220,N_6602,N_7834);
nand U9221 (N_9221,N_6488,N_6539);
nor U9222 (N_9222,N_8773,N_6650);
nor U9223 (N_9223,N_6193,N_8507);
or U9224 (N_9224,N_6698,N_8072);
xor U9225 (N_9225,N_8288,N_7997);
and U9226 (N_9226,N_6186,N_8199);
and U9227 (N_9227,N_8437,N_6862);
nand U9228 (N_9228,N_8084,N_6112);
or U9229 (N_9229,N_6872,N_6230);
and U9230 (N_9230,N_8258,N_8215);
nand U9231 (N_9231,N_7373,N_8028);
nor U9232 (N_9232,N_8184,N_6077);
nand U9233 (N_9233,N_6674,N_8436);
nor U9234 (N_9234,N_8981,N_6583);
nor U9235 (N_9235,N_7500,N_7556);
nand U9236 (N_9236,N_6148,N_8094);
or U9237 (N_9237,N_8222,N_8649);
or U9238 (N_9238,N_7035,N_8664);
nand U9239 (N_9239,N_6117,N_6994);
or U9240 (N_9240,N_6743,N_8040);
or U9241 (N_9241,N_8974,N_6764);
nor U9242 (N_9242,N_6326,N_7256);
nor U9243 (N_9243,N_7584,N_7044);
nor U9244 (N_9244,N_8261,N_6097);
and U9245 (N_9245,N_8486,N_8553);
nand U9246 (N_9246,N_7539,N_7461);
or U9247 (N_9247,N_6599,N_6794);
nand U9248 (N_9248,N_8629,N_8078);
or U9249 (N_9249,N_7821,N_7592);
nand U9250 (N_9250,N_6988,N_6914);
nand U9251 (N_9251,N_8899,N_7715);
nor U9252 (N_9252,N_6576,N_6449);
or U9253 (N_9253,N_7985,N_7863);
or U9254 (N_9254,N_6311,N_7196);
or U9255 (N_9255,N_8353,N_7212);
or U9256 (N_9256,N_8631,N_8341);
or U9257 (N_9257,N_7497,N_7186);
nor U9258 (N_9258,N_6129,N_7018);
or U9259 (N_9259,N_6307,N_6259);
or U9260 (N_9260,N_8472,N_7762);
and U9261 (N_9261,N_6061,N_8089);
and U9262 (N_9262,N_6790,N_7894);
nand U9263 (N_9263,N_8772,N_8054);
nand U9264 (N_9264,N_7562,N_7133);
nor U9265 (N_9265,N_7255,N_6342);
nor U9266 (N_9266,N_8849,N_7408);
and U9267 (N_9267,N_7439,N_7521);
nand U9268 (N_9268,N_6864,N_8286);
nand U9269 (N_9269,N_8965,N_8755);
nand U9270 (N_9270,N_7787,N_7927);
and U9271 (N_9271,N_8406,N_7425);
or U9272 (N_9272,N_6689,N_8706);
or U9273 (N_9273,N_8671,N_7754);
or U9274 (N_9274,N_7358,N_6242);
nor U9275 (N_9275,N_8193,N_7723);
or U9276 (N_9276,N_8016,N_6942);
and U9277 (N_9277,N_8707,N_8563);
or U9278 (N_9278,N_6421,N_7904);
nor U9279 (N_9279,N_7020,N_7876);
or U9280 (N_9280,N_7944,N_8582);
or U9281 (N_9281,N_6781,N_6161);
and U9282 (N_9282,N_7155,N_6883);
or U9283 (N_9283,N_8383,N_7977);
or U9284 (N_9284,N_7006,N_6944);
nor U9285 (N_9285,N_6388,N_6046);
nand U9286 (N_9286,N_6948,N_7257);
or U9287 (N_9287,N_7649,N_6926);
and U9288 (N_9288,N_7137,N_8195);
nor U9289 (N_9289,N_6582,N_7857);
nor U9290 (N_9290,N_7021,N_7300);
or U9291 (N_9291,N_8454,N_7199);
or U9292 (N_9292,N_6506,N_8782);
nand U9293 (N_9293,N_7442,N_6973);
and U9294 (N_9294,N_6075,N_7561);
nand U9295 (N_9295,N_8721,N_6071);
or U9296 (N_9296,N_7732,N_6932);
nand U9297 (N_9297,N_8647,N_7811);
or U9298 (N_9298,N_8470,N_8690);
xnor U9299 (N_9299,N_8648,N_6309);
or U9300 (N_9300,N_6049,N_6445);
or U9301 (N_9301,N_7149,N_7533);
or U9302 (N_9302,N_6085,N_6996);
nor U9303 (N_9303,N_6059,N_8018);
nor U9304 (N_9304,N_7283,N_6398);
or U9305 (N_9305,N_6137,N_8539);
and U9306 (N_9306,N_6138,N_8655);
xnor U9307 (N_9307,N_6696,N_8775);
and U9308 (N_9308,N_8946,N_6348);
and U9309 (N_9309,N_7430,N_7669);
and U9310 (N_9310,N_8999,N_8735);
or U9311 (N_9311,N_6171,N_6670);
nor U9312 (N_9312,N_8082,N_8841);
nand U9313 (N_9313,N_6157,N_7780);
or U9314 (N_9314,N_8642,N_6471);
or U9315 (N_9315,N_7753,N_7690);
xnor U9316 (N_9316,N_8431,N_6598);
and U9317 (N_9317,N_6947,N_8614);
nand U9318 (N_9318,N_7384,N_6007);
or U9319 (N_9319,N_8283,N_8449);
nor U9320 (N_9320,N_8776,N_7956);
nor U9321 (N_9321,N_7013,N_6500);
or U9322 (N_9322,N_7410,N_7417);
or U9323 (N_9323,N_7641,N_7499);
or U9324 (N_9324,N_8583,N_8282);
and U9325 (N_9325,N_6601,N_8915);
nand U9326 (N_9326,N_6635,N_7245);
and U9327 (N_9327,N_7935,N_6125);
or U9328 (N_9328,N_7221,N_8316);
and U9329 (N_9329,N_8294,N_8639);
or U9330 (N_9330,N_8189,N_6651);
and U9331 (N_9331,N_7852,N_7017);
or U9332 (N_9332,N_8778,N_8588);
or U9333 (N_9333,N_6243,N_7140);
or U9334 (N_9334,N_7490,N_7534);
and U9335 (N_9335,N_6937,N_7431);
nor U9336 (N_9336,N_7670,N_8474);
and U9337 (N_9337,N_8159,N_8570);
nor U9338 (N_9338,N_7725,N_7383);
or U9339 (N_9339,N_7816,N_6912);
nor U9340 (N_9340,N_6036,N_7917);
nand U9341 (N_9341,N_7089,N_6336);
nand U9342 (N_9342,N_8125,N_7193);
or U9343 (N_9343,N_8584,N_7240);
nand U9344 (N_9344,N_6585,N_7924);
nand U9345 (N_9345,N_6548,N_7328);
xnor U9346 (N_9346,N_6407,N_8497);
and U9347 (N_9347,N_7367,N_8214);
nor U9348 (N_9348,N_8153,N_6209);
nand U9349 (N_9349,N_6039,N_6113);
nand U9350 (N_9350,N_8145,N_8446);
or U9351 (N_9351,N_8743,N_6789);
nand U9352 (N_9352,N_7389,N_6319);
and U9353 (N_9353,N_8506,N_7508);
nand U9354 (N_9354,N_8504,N_7667);
or U9355 (N_9355,N_8146,N_8813);
nand U9356 (N_9356,N_6530,N_6383);
nand U9357 (N_9357,N_8070,N_6776);
nor U9358 (N_9358,N_8438,N_6158);
nor U9359 (N_9359,N_7960,N_8414);
nand U9360 (N_9360,N_6305,N_6267);
nor U9361 (N_9361,N_8050,N_8916);
or U9362 (N_9362,N_6358,N_6751);
and U9363 (N_9363,N_6578,N_8501);
nor U9364 (N_9364,N_7139,N_6939);
and U9365 (N_9365,N_6826,N_7166);
nand U9366 (N_9366,N_7037,N_7727);
or U9367 (N_9367,N_8407,N_6045);
and U9368 (N_9368,N_7902,N_7764);
and U9369 (N_9369,N_7648,N_6785);
nor U9370 (N_9370,N_8161,N_6524);
or U9371 (N_9371,N_8440,N_7299);
and U9372 (N_9372,N_8357,N_6214);
and U9373 (N_9373,N_6005,N_6132);
or U9374 (N_9374,N_7689,N_6135);
nand U9375 (N_9375,N_6018,N_6343);
and U9376 (N_9376,N_7832,N_8968);
nor U9377 (N_9377,N_8336,N_8024);
or U9378 (N_9378,N_7665,N_7920);
or U9379 (N_9379,N_6264,N_6424);
nor U9380 (N_9380,N_6928,N_6216);
nor U9381 (N_9381,N_6215,N_8427);
nand U9382 (N_9382,N_6416,N_6226);
or U9383 (N_9383,N_6282,N_8480);
and U9384 (N_9384,N_6187,N_6453);
or U9385 (N_9385,N_6618,N_6123);
nor U9386 (N_9386,N_6505,N_7619);
xnor U9387 (N_9387,N_8093,N_7074);
and U9388 (N_9388,N_7046,N_6295);
or U9389 (N_9389,N_8491,N_8192);
xnor U9390 (N_9390,N_8122,N_8903);
or U9391 (N_9391,N_7568,N_8317);
nand U9392 (N_9392,N_8646,N_7940);
or U9393 (N_9393,N_8929,N_7298);
nor U9394 (N_9394,N_8548,N_8170);
or U9395 (N_9395,N_7885,N_6773);
and U9396 (N_9396,N_8132,N_8080);
nor U9397 (N_9397,N_8619,N_6512);
or U9398 (N_9398,N_7263,N_6527);
nand U9399 (N_9399,N_7760,N_8991);
or U9400 (N_9400,N_8730,N_8275);
nor U9401 (N_9401,N_6066,N_7348);
nor U9402 (N_9402,N_6054,N_8099);
nand U9403 (N_9403,N_7951,N_8263);
and U9404 (N_9404,N_7342,N_6008);
nor U9405 (N_9405,N_6608,N_6182);
nor U9406 (N_9406,N_8699,N_6962);
or U9407 (N_9407,N_8908,N_8305);
nand U9408 (N_9408,N_6442,N_6000);
nand U9409 (N_9409,N_8220,N_8542);
and U9410 (N_9410,N_8815,N_8520);
xnor U9411 (N_9411,N_8450,N_8987);
nor U9412 (N_9412,N_6812,N_6096);
or U9413 (N_9413,N_7827,N_7370);
or U9414 (N_9414,N_7467,N_8345);
or U9415 (N_9415,N_7535,N_8262);
nand U9416 (N_9416,N_7906,N_8688);
nand U9417 (N_9417,N_6324,N_7176);
nand U9418 (N_9418,N_8951,N_6967);
and U9419 (N_9419,N_8605,N_7701);
or U9420 (N_9420,N_8277,N_6177);
nand U9421 (N_9421,N_7003,N_7147);
nor U9422 (N_9422,N_8043,N_7489);
nand U9423 (N_9423,N_6367,N_6009);
and U9424 (N_9424,N_8577,N_8700);
nor U9425 (N_9425,N_8375,N_8053);
and U9426 (N_9426,N_6197,N_6705);
or U9427 (N_9427,N_7102,N_7400);
nand U9428 (N_9428,N_7239,N_7415);
and U9429 (N_9429,N_8874,N_6657);
or U9430 (N_9430,N_7041,N_8826);
and U9431 (N_9431,N_8493,N_7936);
and U9432 (N_9432,N_6133,N_6217);
nand U9433 (N_9433,N_7476,N_7859);
nand U9434 (N_9434,N_8012,N_7301);
or U9435 (N_9435,N_7662,N_8144);
nand U9436 (N_9436,N_7803,N_7282);
and U9437 (N_9437,N_6194,N_8120);
or U9438 (N_9438,N_6498,N_8993);
nand U9439 (N_9439,N_8618,N_7357);
or U9440 (N_9440,N_7195,N_6518);
nor U9441 (N_9441,N_6580,N_8300);
nand U9442 (N_9442,N_7073,N_8166);
or U9443 (N_9443,N_7739,N_7159);
nand U9444 (N_9444,N_6536,N_6676);
or U9445 (N_9445,N_8695,N_7208);
nor U9446 (N_9446,N_8112,N_8967);
nand U9447 (N_9447,N_6115,N_8212);
nor U9448 (N_9448,N_7048,N_6909);
or U9449 (N_9449,N_7338,N_6116);
xor U9450 (N_9450,N_7962,N_7650);
nor U9451 (N_9451,N_8361,N_8680);
and U9452 (N_9452,N_6219,N_7520);
nand U9453 (N_9453,N_6374,N_7835);
or U9454 (N_9454,N_6245,N_6090);
nand U9455 (N_9455,N_6220,N_7874);
nor U9456 (N_9456,N_6616,N_7031);
nand U9457 (N_9457,N_8381,N_6362);
nor U9458 (N_9458,N_6644,N_8997);
xor U9459 (N_9459,N_7513,N_7387);
nand U9460 (N_9460,N_7038,N_8092);
and U9461 (N_9461,N_7368,N_6410);
or U9462 (N_9462,N_7845,N_7216);
nor U9463 (N_9463,N_7993,N_7982);
and U9464 (N_9464,N_8711,N_6853);
and U9465 (N_9465,N_7306,N_8141);
nand U9466 (N_9466,N_6550,N_7381);
or U9467 (N_9467,N_6058,N_6870);
or U9468 (N_9468,N_6641,N_7905);
nand U9469 (N_9469,N_7321,N_7546);
and U9470 (N_9470,N_7607,N_7661);
nand U9471 (N_9471,N_7095,N_8744);
nand U9472 (N_9472,N_8872,N_6122);
and U9473 (N_9473,N_7779,N_6188);
and U9474 (N_9474,N_8169,N_7999);
and U9475 (N_9475,N_8108,N_7000);
and U9476 (N_9476,N_7970,N_6418);
nor U9477 (N_9477,N_7363,N_6255);
and U9478 (N_9478,N_8526,N_6715);
or U9479 (N_9479,N_8061,N_8398);
nor U9480 (N_9480,N_6879,N_6068);
and U9481 (N_9481,N_6035,N_7353);
nor U9482 (N_9482,N_7578,N_6614);
and U9483 (N_9483,N_8000,N_7840);
nand U9484 (N_9484,N_6593,N_7580);
or U9485 (N_9485,N_6856,N_7583);
and U9486 (N_9486,N_6554,N_7356);
nand U9487 (N_9487,N_7822,N_8291);
nand U9488 (N_9488,N_8386,N_6377);
nand U9489 (N_9489,N_8681,N_8777);
nor U9490 (N_9490,N_7437,N_8931);
nor U9491 (N_9491,N_6159,N_6088);
nand U9492 (N_9492,N_8110,N_6433);
or U9493 (N_9493,N_6142,N_7419);
or U9494 (N_9494,N_6963,N_8927);
nand U9495 (N_9495,N_7750,N_7138);
and U9496 (N_9496,N_8531,N_6531);
and U9497 (N_9497,N_7153,N_8621);
nand U9498 (N_9498,N_6570,N_8670);
nand U9499 (N_9499,N_7350,N_6777);
or U9500 (N_9500,N_8888,N_7406);
nor U9501 (N_9501,N_8889,N_7331);
and U9502 (N_9502,N_6464,N_6998);
nand U9503 (N_9503,N_8364,N_6402);
nor U9504 (N_9504,N_7559,N_8458);
nor U9505 (N_9505,N_8373,N_8322);
nand U9506 (N_9506,N_7271,N_7391);
nand U9507 (N_9507,N_7065,N_6757);
nor U9508 (N_9508,N_7494,N_7907);
xnor U9509 (N_9509,N_7506,N_8284);
xnor U9510 (N_9510,N_7327,N_7495);
nor U9511 (N_9511,N_6353,N_6581);
nor U9512 (N_9512,N_6455,N_8421);
nand U9513 (N_9513,N_7264,N_6766);
xor U9514 (N_9514,N_6687,N_6995);
or U9515 (N_9515,N_7453,N_8413);
nor U9516 (N_9516,N_6386,N_6083);
nand U9517 (N_9517,N_7484,N_6392);
nand U9518 (N_9518,N_8733,N_8580);
nand U9519 (N_9519,N_6917,N_8479);
or U9520 (N_9520,N_8712,N_7774);
and U9521 (N_9521,N_7558,N_7440);
nor U9522 (N_9522,N_6541,N_8992);
and U9523 (N_9523,N_6787,N_7527);
nor U9524 (N_9524,N_6098,N_6033);
nor U9525 (N_9525,N_8754,N_6759);
xor U9526 (N_9526,N_6528,N_6020);
nand U9527 (N_9527,N_6935,N_8887);
nor U9528 (N_9528,N_7635,N_7613);
or U9529 (N_9529,N_7308,N_7359);
or U9530 (N_9530,N_8608,N_7595);
or U9531 (N_9531,N_8293,N_7265);
nor U9532 (N_9532,N_8188,N_8359);
and U9533 (N_9533,N_6979,N_8124);
nor U9534 (N_9534,N_7173,N_7930);
nor U9535 (N_9535,N_6770,N_7378);
nand U9536 (N_9536,N_8209,N_6529);
nand U9537 (N_9537,N_8661,N_7519);
nor U9538 (N_9538,N_6659,N_6800);
or U9539 (N_9539,N_8259,N_6725);
nand U9540 (N_9540,N_6905,N_7554);
and U9541 (N_9541,N_6292,N_7676);
xnor U9542 (N_9542,N_8063,N_6744);
nor U9543 (N_9543,N_7250,N_7849);
and U9544 (N_9544,N_8518,N_7998);
xor U9545 (N_9545,N_7232,N_6628);
and U9546 (N_9546,N_8439,N_8121);
and U9547 (N_9547,N_8725,N_8561);
or U9548 (N_9548,N_8766,N_8689);
nand U9549 (N_9549,N_8761,N_7165);
nor U9550 (N_9550,N_8623,N_7567);
nor U9551 (N_9551,N_7593,N_8774);
nor U9552 (N_9552,N_8515,N_7311);
nand U9553 (N_9553,N_8004,N_6851);
nand U9554 (N_9554,N_7456,N_8938);
and U9555 (N_9555,N_7867,N_8245);
or U9556 (N_9556,N_6809,N_7274);
nor U9557 (N_9557,N_8424,N_6425);
and U9558 (N_9558,N_7123,N_8425);
nor U9559 (N_9559,N_7575,N_6565);
and U9560 (N_9560,N_7062,N_8850);
and U9561 (N_9561,N_8380,N_8240);
and U9562 (N_9562,N_6070,N_8741);
nand U9563 (N_9563,N_8865,N_7101);
and U9564 (N_9564,N_8478,N_7488);
nand U9565 (N_9565,N_6952,N_6503);
and U9566 (N_9566,N_8311,N_8651);
nor U9567 (N_9567,N_8937,N_6890);
xnor U9568 (N_9568,N_7925,N_6830);
nand U9569 (N_9569,N_6210,N_6222);
xor U9570 (N_9570,N_7703,N_7707);
or U9571 (N_9571,N_8988,N_8934);
nor U9572 (N_9572,N_6986,N_6936);
nor U9573 (N_9573,N_6886,N_8544);
and U9574 (N_9574,N_6666,N_8750);
xnor U9575 (N_9575,N_6831,N_8123);
or U9576 (N_9576,N_6218,N_7225);
nand U9577 (N_9577,N_8022,N_8363);
or U9578 (N_9578,N_6459,N_6733);
xnor U9579 (N_9579,N_6249,N_7677);
nand U9580 (N_9580,N_7319,N_8298);
xor U9581 (N_9581,N_7786,N_6467);
nand U9582 (N_9582,N_8678,N_8205);
nand U9583 (N_9583,N_8190,N_8109);
and U9584 (N_9584,N_7652,N_7609);
nand U9585 (N_9585,N_8597,N_7883);
nor U9586 (N_9586,N_8370,N_7148);
nand U9587 (N_9587,N_8175,N_7626);
and U9588 (N_9588,N_6726,N_8576);
nand U9589 (N_9589,N_7812,N_8429);
and U9590 (N_9590,N_7293,N_6846);
and U9591 (N_9591,N_7252,N_8897);
or U9592 (N_9592,N_8181,N_7423);
nand U9593 (N_9593,N_6643,N_7973);
or U9594 (N_9594,N_6349,N_6724);
or U9595 (N_9595,N_6300,N_8901);
or U9596 (N_9596,N_6920,N_8592);
or U9597 (N_9597,N_8601,N_8869);
and U9598 (N_9598,N_8451,N_6284);
nand U9599 (N_9599,N_8447,N_6756);
or U9600 (N_9600,N_7828,N_6825);
and U9601 (N_9601,N_7097,N_8599);
and U9602 (N_9602,N_6861,N_6680);
and U9603 (N_9603,N_8918,N_6898);
or U9604 (N_9604,N_7544,N_6927);
nor U9605 (N_9605,N_7207,N_8545);
and U9606 (N_9606,N_7470,N_8977);
nand U9607 (N_9607,N_7873,N_6192);
and U9608 (N_9608,N_6525,N_6151);
and U9609 (N_9609,N_8471,N_8225);
nor U9610 (N_9610,N_6280,N_7053);
nor U9611 (N_9611,N_6064,N_8163);
and U9612 (N_9612,N_6286,N_7913);
nor U9613 (N_9613,N_7210,N_8473);
nor U9614 (N_9614,N_7722,N_7142);
and U9615 (N_9615,N_6720,N_6204);
nor U9616 (N_9616,N_6782,N_7092);
or U9617 (N_9617,N_8679,N_8960);
nor U9618 (N_9618,N_7181,N_8783);
or U9619 (N_9619,N_7040,N_7078);
or U9620 (N_9620,N_8950,N_6537);
nand U9621 (N_9621,N_8045,N_6538);
nor U9622 (N_9622,N_6462,N_7033);
nor U9623 (N_9623,N_7402,N_7487);
and U9624 (N_9624,N_6603,N_8031);
or U9625 (N_9625,N_7228,N_7644);
or U9626 (N_9626,N_7157,N_6638);
or U9627 (N_9627,N_6191,N_7188);
nand U9628 (N_9628,N_7030,N_8324);
and U9629 (N_9629,N_7931,N_7889);
nand U9630 (N_9630,N_6195,N_7455);
nor U9631 (N_9631,N_8719,N_6178);
and U9632 (N_9632,N_6841,N_7830);
nand U9633 (N_9633,N_6139,N_8138);
nand U9634 (N_9634,N_8831,N_6551);
nor U9635 (N_9635,N_7361,N_6993);
nand U9636 (N_9636,N_6975,N_7655);
and U9637 (N_9637,N_7711,N_6663);
or U9638 (N_9638,N_7128,N_8158);
nor U9639 (N_9639,N_8339,N_8793);
or U9640 (N_9640,N_6254,N_8056);
or U9641 (N_9641,N_7452,N_8218);
and U9642 (N_9642,N_8663,N_8734);
nand U9643 (N_9643,N_6360,N_8959);
and U9644 (N_9644,N_6850,N_6814);
nor U9645 (N_9645,N_6263,N_7995);
and U9646 (N_9646,N_7323,N_8803);
nor U9647 (N_9647,N_6807,N_7869);
nand U9648 (N_9648,N_8385,N_6034);
nand U9649 (N_9649,N_6736,N_6359);
or U9650 (N_9650,N_8384,N_6592);
nor U9651 (N_9651,N_8828,N_8945);
and U9652 (N_9652,N_6321,N_7024);
nor U9653 (N_9653,N_8315,N_8465);
or U9654 (N_9654,N_8795,N_6571);
and U9655 (N_9655,N_8185,N_8891);
nor U9656 (N_9656,N_8071,N_8591);
nor U9657 (N_9657,N_7066,N_8611);
nand U9658 (N_9658,N_6738,N_7596);
or U9659 (N_9659,N_6276,N_7451);
and U9660 (N_9660,N_8227,N_6984);
and U9661 (N_9661,N_7862,N_8676);
nand U9662 (N_9662,N_8697,N_7865);
and U9663 (N_9663,N_6559,N_6639);
and U9664 (N_9664,N_6232,N_7163);
nor U9665 (N_9665,N_7981,N_6169);
and U9666 (N_9666,N_6533,N_7178);
nor U9667 (N_9667,N_7124,N_6340);
nor U9668 (N_9668,N_8034,N_8508);
and U9669 (N_9669,N_8575,N_7929);
and U9670 (N_9670,N_6892,N_8186);
or U9671 (N_9671,N_6735,N_7685);
nor U9672 (N_9672,N_7895,N_7237);
nor U9673 (N_9673,N_8551,N_6523);
or U9674 (N_9674,N_6274,N_6352);
nand U9675 (N_9675,N_8973,N_8923);
and U9676 (N_9676,N_6802,N_6160);
nand U9677 (N_9677,N_6957,N_8150);
and U9678 (N_9678,N_8514,N_7706);
nand U9679 (N_9679,N_7932,N_6212);
xnor U9680 (N_9680,N_7002,N_8635);
and U9681 (N_9681,N_7587,N_8130);
and U9682 (N_9682,N_6843,N_8710);
and U9683 (N_9683,N_6417,N_6155);
nor U9684 (N_9684,N_8434,N_7809);
or U9685 (N_9685,N_8904,N_6457);
or U9686 (N_9686,N_7643,N_7611);
nand U9687 (N_9687,N_7926,N_7958);
and U9688 (N_9688,N_6513,N_6233);
nor U9689 (N_9689,N_6397,N_6982);
and U9690 (N_9690,N_8976,N_8779);
xor U9691 (N_9691,N_6605,N_7241);
nand U9692 (N_9692,N_7721,N_7433);
and U9693 (N_9693,N_7766,N_8522);
xnor U9694 (N_9694,N_7819,N_7187);
or U9695 (N_9695,N_7152,N_6109);
nand U9696 (N_9696,N_8296,N_6391);
nor U9697 (N_9697,N_7132,N_6649);
nand U9698 (N_9698,N_8644,N_6015);
nor U9699 (N_9699,N_6350,N_7937);
or U9700 (N_9700,N_7007,N_7269);
nand U9701 (N_9701,N_7861,N_6646);
nand U9702 (N_9702,N_8528,N_6250);
or U9703 (N_9703,N_6818,N_7347);
or U9704 (N_9704,N_7980,N_8516);
or U9705 (N_9705,N_8174,N_6771);
xor U9706 (N_9706,N_6832,N_6476);
or U9707 (N_9707,N_8740,N_7295);
and U9708 (N_9708,N_6949,N_8076);
nand U9709 (N_9709,N_6568,N_8693);
nand U9710 (N_9710,N_7716,N_6819);
or U9711 (N_9711,N_7088,N_7377);
nand U9712 (N_9712,N_6881,N_7657);
nand U9713 (N_9713,N_8786,N_6380);
nor U9714 (N_9714,N_6201,N_6144);
or U9715 (N_9715,N_8898,N_8015);
xor U9716 (N_9716,N_6612,N_6697);
or U9717 (N_9717,N_7605,N_6681);
nand U9718 (N_9718,N_8878,N_6627);
and U9719 (N_9719,N_8509,N_6712);
or U9720 (N_9720,N_7238,N_8371);
nor U9721 (N_9721,N_7682,N_7125);
and U9722 (N_9722,N_6857,N_6283);
nand U9723 (N_9723,N_8418,N_6312);
or U9724 (N_9724,N_7965,N_7141);
nand U9725 (N_9725,N_8468,N_7881);
and U9726 (N_9726,N_7343,N_7899);
and U9727 (N_9727,N_7839,N_7458);
nor U9728 (N_9728,N_6784,N_7280);
nand U9729 (N_9729,N_6980,N_7438);
or U9730 (N_9730,N_7224,N_8051);
nand U9731 (N_9731,N_6971,N_8705);
and U9732 (N_9732,N_7776,N_6897);
nor U9733 (N_9733,N_7393,N_6567);
or U9734 (N_9734,N_7976,N_6758);
and U9735 (N_9735,N_7249,N_8533);
nor U9736 (N_9736,N_8235,N_6906);
nor U9737 (N_9737,N_6345,N_8127);
nor U9738 (N_9738,N_8103,N_7854);
nand U9739 (N_9739,N_7504,N_6450);
nor U9740 (N_9740,N_7922,N_7975);
or U9741 (N_9741,N_7557,N_8821);
nor U9742 (N_9742,N_7890,N_8302);
and U9743 (N_9743,N_6099,N_8086);
or U9744 (N_9744,N_6454,N_8297);
or U9745 (N_9745,N_8173,N_6707);
nand U9746 (N_9746,N_8096,N_8672);
nor U9747 (N_9747,N_6717,N_6821);
nor U9748 (N_9748,N_8566,N_7693);
and U9749 (N_9749,N_6596,N_7798);
nand U9750 (N_9750,N_8892,N_8010);
nor U9751 (N_9751,N_6452,N_8738);
nand U9752 (N_9752,N_7773,N_7949);
or U9753 (N_9753,N_6431,N_6376);
or U9754 (N_9754,N_7115,N_6074);
nand U9755 (N_9755,N_8606,N_6817);
and U9756 (N_9756,N_7206,N_8422);
xor U9757 (N_9757,N_8834,N_6839);
nor U9758 (N_9758,N_6594,N_7517);
and U9759 (N_9759,N_8805,N_7329);
and U9760 (N_9760,N_7352,N_6396);
nor U9761 (N_9761,N_8312,N_8133);
and U9762 (N_9762,N_7934,N_7135);
nand U9763 (N_9763,N_8285,N_8607);
nor U9764 (N_9764,N_7266,N_8019);
nand U9765 (N_9765,N_6718,N_8814);
nand U9766 (N_9766,N_6589,N_6855);
or U9767 (N_9767,N_7229,N_7045);
and U9768 (N_9768,N_6346,N_6907);
and U9769 (N_9769,N_8983,N_8837);
nor U9770 (N_9770,N_7952,N_7536);
or U9771 (N_9771,N_8948,N_8233);
or U9772 (N_9772,N_8448,N_8844);
nor U9773 (N_9773,N_6786,N_8804);
nand U9774 (N_9774,N_7105,N_8289);
nand U9775 (N_9775,N_6170,N_7694);
and U9776 (N_9776,N_6976,N_7680);
and U9777 (N_9777,N_8280,N_8477);
or U9778 (N_9778,N_6704,N_7638);
and U9779 (N_9779,N_6772,N_7618);
or U9780 (N_9780,N_6532,N_8253);
or U9781 (N_9781,N_8131,N_6146);
nor U9782 (N_9782,N_6032,N_7528);
nand U9783 (N_9783,N_8287,N_6793);
or U9784 (N_9784,N_8279,N_8970);
or U9785 (N_9785,N_6126,N_8115);
nand U9786 (N_9786,N_7156,N_8863);
or U9787 (N_9787,N_6956,N_7698);
and U9788 (N_9788,N_7681,N_7692);
or U9789 (N_9789,N_7623,N_8652);
and U9790 (N_9790,N_8069,N_6882);
and U9791 (N_9791,N_6929,N_8781);
nand U9792 (N_9792,N_8066,N_6095);
or U9793 (N_9793,N_8464,N_8502);
and U9794 (N_9794,N_7509,N_8986);
nor U9795 (N_9795,N_6121,N_8246);
nand U9796 (N_9796,N_8512,N_7911);
nand U9797 (N_9797,N_8505,N_8264);
nand U9798 (N_9798,N_8460,N_7162);
xor U9799 (N_9799,N_8428,N_8023);
nand U9800 (N_9800,N_7505,N_7449);
nor U9801 (N_9801,N_8077,N_8241);
or U9802 (N_9802,N_8896,N_8223);
and U9803 (N_9803,N_7775,N_6634);
or U9804 (N_9804,N_7683,N_6901);
or U9805 (N_9805,N_6465,N_6867);
nor U9806 (N_9806,N_6683,N_7325);
or U9807 (N_9807,N_7646,N_7502);
nor U9808 (N_9808,N_7668,N_8039);
and U9809 (N_9809,N_8729,N_6556);
nand U9810 (N_9810,N_8393,N_7564);
nor U9811 (N_9811,N_6685,N_7818);
nand U9812 (N_9812,N_6535,N_6765);
or U9813 (N_9813,N_8204,N_8481);
nand U9814 (N_9814,N_8866,N_8452);
nand U9815 (N_9815,N_6461,N_8139);
nor U9816 (N_9816,N_8490,N_8221);
nand U9817 (N_9817,N_6919,N_7227);
or U9818 (N_9818,N_8667,N_7466);
nand U9819 (N_9819,N_6458,N_7887);
nor U9820 (N_9820,N_8105,N_7622);
nand U9821 (N_9821,N_8467,N_6289);
nor U9822 (N_9822,N_8732,N_7272);
and U9823 (N_9823,N_8532,N_6323);
or U9824 (N_9824,N_6729,N_6355);
and U9825 (N_9825,N_8052,N_6624);
nand U9826 (N_9826,N_6965,N_8310);
and U9827 (N_9827,N_8405,N_6501);
nor U9828 (N_9828,N_7177,N_6208);
or U9829 (N_9829,N_7532,N_8162);
nor U9830 (N_9830,N_6317,N_6269);
and U9831 (N_9831,N_6924,N_6330);
and U9832 (N_9832,N_8882,N_6196);
nand U9833 (N_9833,N_6406,N_7959);
and U9834 (N_9834,N_7720,N_6648);
nor U9835 (N_9835,N_7215,N_6516);
and U9836 (N_9836,N_6202,N_7675);
nor U9837 (N_9837,N_7154,N_8914);
nor U9838 (N_9838,N_7663,N_7785);
or U9839 (N_9839,N_8256,N_7695);
or U9840 (N_9840,N_7150,N_6858);
and U9841 (N_9841,N_8017,N_7313);
or U9842 (N_9842,N_8975,N_7042);
nor U9843 (N_9843,N_8171,N_8990);
nand U9844 (N_9844,N_8964,N_8747);
nand U9845 (N_9845,N_8900,N_8101);
nand U9846 (N_9846,N_6012,N_6167);
nor U9847 (N_9847,N_7791,N_6329);
or U9848 (N_9848,N_7254,N_8910);
or U9849 (N_9849,N_8036,N_7994);
nand U9850 (N_9850,N_6768,N_8098);
and U9851 (N_9851,N_6405,N_8824);
nor U9852 (N_9852,N_7824,N_6239);
and U9853 (N_9853,N_8198,N_8691);
xnor U9854 (N_9854,N_7968,N_7464);
and U9855 (N_9855,N_7914,N_7820);
nand U9856 (N_9856,N_7482,N_7728);
and U9857 (N_9857,N_8157,N_6444);
or U9858 (N_9858,N_6296,N_8790);
or U9859 (N_9859,N_6168,N_6915);
nand U9860 (N_9860,N_6240,N_8737);
and U9861 (N_9861,N_7422,N_8838);
nor U9862 (N_9862,N_8389,N_6610);
nand U9863 (N_9863,N_8870,N_8059);
or U9864 (N_9864,N_7214,N_8660);
and U9865 (N_9865,N_6692,N_7427);
and U9866 (N_9866,N_6470,N_6069);
nand U9867 (N_9867,N_7886,N_7784);
nand U9868 (N_9868,N_8041,N_8492);
or U9869 (N_9869,N_6660,N_8854);
nor U9870 (N_9870,N_8113,N_7823);
nand U9871 (N_9871,N_7537,N_8488);
or U9872 (N_9872,N_6272,N_8829);
and U9873 (N_9873,N_8634,N_6708);
nand U9874 (N_9874,N_6265,N_7420);
nor U9875 (N_9875,N_7983,N_6294);
nand U9876 (N_9876,N_8559,N_6668);
or U9877 (N_9877,N_6082,N_8351);
nor U9878 (N_9878,N_7770,N_8928);
nand U9879 (N_9879,N_8271,N_8309);
and U9880 (N_9880,N_8213,N_6590);
nand U9881 (N_9881,N_7640,N_7376);
and U9882 (N_9882,N_6140,N_8694);
and U9883 (N_9883,N_6373,N_6852);
nand U9884 (N_9884,N_8962,N_7404);
nor U9885 (N_9885,N_6918,N_8812);
and U9886 (N_9886,N_7011,N_8065);
or U9887 (N_9887,N_7569,N_7702);
nand U9888 (N_9888,N_6645,N_6002);
and U9889 (N_9889,N_6303,N_6562);
and U9890 (N_9890,N_6834,N_6102);
nor U9891 (N_9891,N_8435,N_6314);
nand U9892 (N_9892,N_8825,N_6549);
and U9893 (N_9893,N_8002,N_8716);
nor U9894 (N_9894,N_7366,N_6563);
and U9895 (N_9895,N_8787,N_8503);
nand U9896 (N_9896,N_7733,N_7183);
nor U9897 (N_9897,N_7942,N_7525);
and U9898 (N_9898,N_6180,N_8753);
or U9899 (N_9899,N_8304,N_7572);
or U9900 (N_9900,N_8685,N_8519);
or U9901 (N_9901,N_8996,N_8947);
or U9902 (N_9902,N_7413,N_8636);
or U9903 (N_9903,N_8683,N_6502);
nand U9904 (N_9904,N_6351,N_8152);
and U9905 (N_9905,N_8167,N_7117);
and U9906 (N_9906,N_8191,N_6100);
nor U9907 (N_9907,N_7236,N_7388);
nand U9908 (N_9908,N_7741,N_6591);
nor U9909 (N_9909,N_8536,N_8613);
nor U9910 (N_9910,N_6763,N_7203);
or U9911 (N_9911,N_7735,N_8883);
and U9912 (N_9912,N_8550,N_7086);
and U9913 (N_9913,N_6181,N_8861);
nand U9914 (N_9914,N_6298,N_8994);
and U9915 (N_9915,N_6361,N_6310);
and U9916 (N_9916,N_8088,N_8547);
nand U9917 (N_9917,N_7332,N_6474);
nor U9918 (N_9918,N_8217,N_7918);
nor U9919 (N_9919,N_6014,N_7672);
nand U9920 (N_9920,N_6978,N_8925);
nand U9921 (N_9921,N_6320,N_7316);
nand U9922 (N_9922,N_7219,N_6091);
nor U9923 (N_9923,N_7379,N_6435);
nand U9924 (N_9924,N_7310,N_7180);
and U9925 (N_9925,N_7457,N_8907);
or U9926 (N_9926,N_6896,N_6060);
or U9927 (N_9927,N_7737,N_8172);
xor U9928 (N_9928,N_7802,N_6087);
nor U9929 (N_9929,N_7553,N_8456);
nand U9930 (N_9930,N_6769,N_6393);
nand U9931 (N_9931,N_7113,N_8469);
nor U9932 (N_9932,N_7351,N_6597);
and U9933 (N_9933,N_6943,N_7027);
and U9934 (N_9934,N_8420,N_8236);
nand U9935 (N_9935,N_7853,N_8347);
nand U9936 (N_9936,N_8589,N_8718);
and U9937 (N_9937,N_7825,N_7659);
nor U9938 (N_9938,N_6290,N_7201);
and U9939 (N_9939,N_8443,N_7485);
or U9940 (N_9940,N_8956,N_7004);
or U9941 (N_9941,N_7901,N_8114);
or U9942 (N_9942,N_8620,N_8290);
or U9943 (N_9943,N_7815,N_6244);
nor U9944 (N_9944,N_8224,N_6288);
and U9945 (N_9945,N_8165,N_7336);
or U9946 (N_9946,N_8009,N_6466);
nor U9947 (N_9947,N_7686,N_7322);
nand U9948 (N_9948,N_6653,N_7043);
xor U9949 (N_9949,N_7111,N_7218);
nor U9950 (N_9950,N_7057,N_6792);
and U9951 (N_9951,N_6647,N_6654);
nand U9952 (N_9952,N_6004,N_6308);
or U9953 (N_9953,N_8201,N_6150);
nor U9954 (N_9954,N_8989,N_8641);
nand U9955 (N_9955,N_8090,N_8846);
or U9956 (N_9956,N_7632,N_7602);
nor U9957 (N_9957,N_7664,N_6569);
and U9958 (N_9958,N_8349,N_7344);
or U9959 (N_9959,N_6399,N_6363);
nand U9960 (N_9960,N_6625,N_6803);
nand U9961 (N_9961,N_7738,N_6731);
nor U9962 (N_9962,N_8247,N_6910);
or U9963 (N_9963,N_7185,N_8816);
or U9964 (N_9964,N_6278,N_8585);
nand U9965 (N_9965,N_8810,N_6428);
and U9966 (N_9966,N_7050,N_6412);
nor U9967 (N_9967,N_7826,N_7547);
and U9968 (N_9968,N_7459,N_7380);
or U9969 (N_9969,N_6318,N_8572);
nand U9970 (N_9970,N_7052,N_8376);
and U9971 (N_9971,N_6762,N_7576);
and U9972 (N_9972,N_8273,N_8027);
or U9973 (N_9973,N_6205,N_8650);
or U9974 (N_9974,N_6332,N_7168);
or U9975 (N_9975,N_6561,N_7989);
and U9976 (N_9976,N_8219,N_7028);
or U9977 (N_9977,N_7291,N_6114);
and U9978 (N_9978,N_8511,N_8196);
nand U9979 (N_9979,N_6933,N_8111);
nor U9980 (N_9980,N_6023,N_8276);
or U9981 (N_9981,N_8475,N_7778);
or U9982 (N_9982,N_8415,N_7745);
and U9983 (N_9983,N_6778,N_7281);
nand U9984 (N_9984,N_6740,N_6900);
and U9985 (N_9985,N_7621,N_8573);
nand U9986 (N_9986,N_6631,N_7465);
nand U9987 (N_9987,N_6483,N_8228);
or U9988 (N_9988,N_8554,N_7001);
nor U9989 (N_9989,N_7740,N_7278);
or U9990 (N_9990,N_8379,N_7915);
nand U9991 (N_9991,N_7443,N_6024);
and U9992 (N_9992,N_8292,N_7708);
and U9993 (N_9993,N_7579,N_8770);
and U9994 (N_9994,N_8958,N_6873);
and U9995 (N_9995,N_6682,N_8587);
nand U9996 (N_9996,N_8523,N_8365);
nor U9997 (N_9997,N_6489,N_8858);
nor U9998 (N_9998,N_8229,N_6485);
nand U9999 (N_9999,N_6969,N_7297);
or U10000 (N_10000,N_7943,N_6543);
nor U10001 (N_10001,N_8768,N_6555);
and U10002 (N_10002,N_7759,N_7794);
or U10003 (N_10003,N_6492,N_6675);
and U10004 (N_10004,N_7531,N_7908);
nand U10005 (N_10005,N_6163,N_7294);
or U10006 (N_10006,N_8320,N_7261);
or U10007 (N_10007,N_8924,N_8568);
nor U10008 (N_10008,N_7190,N_6938);
or U10009 (N_10009,N_7551,N_7036);
xor U10010 (N_10010,N_7116,N_8541);
or U10011 (N_10011,N_7444,N_8806);
or U10012 (N_10012,N_6106,N_6623);
and U10013 (N_10013,N_7223,N_6262);
or U10014 (N_10014,N_8557,N_6235);
nand U10015 (N_10015,N_6534,N_6490);
nand U10016 (N_10016,N_7182,N_6946);
and U10017 (N_10017,N_8792,N_7912);
nand U10018 (N_10018,N_6394,N_7337);
or U10019 (N_10019,N_6211,N_6179);
and U10020 (N_10020,N_6991,N_6691);
or U10021 (N_10021,N_7751,N_8408);
or U10022 (N_10022,N_6213,N_7630);
or U10023 (N_10023,N_8020,N_6652);
nor U10024 (N_10024,N_6105,N_6899);
nor U10025 (N_10025,N_8530,N_8535);
nor U10026 (N_10026,N_6699,N_8495);
and U10027 (N_10027,N_6143,N_7518);
nand U10028 (N_10028,N_8091,N_6134);
and U10029 (N_10029,N_6063,N_6426);
nor U10030 (N_10030,N_6621,N_7979);
xnor U10031 (N_10031,N_8135,N_7047);
or U10032 (N_10032,N_6413,N_8935);
nor U10033 (N_10033,N_7429,N_8060);
nor U10034 (N_10034,N_7523,N_7878);
nor U10035 (N_10035,N_6824,N_6779);
nand U10036 (N_10036,N_8338,N_7909);
and U10037 (N_10037,N_6297,N_7591);
nand U10038 (N_10038,N_8827,N_8596);
nand U10039 (N_10039,N_8726,N_6600);
or U10040 (N_10040,N_6382,N_8785);
nor U10041 (N_10041,N_7079,N_7654);
or U10042 (N_10042,N_6154,N_6152);
nand U10043 (N_10043,N_7317,N_7829);
nor U10044 (N_10044,N_6783,N_7345);
or U10045 (N_10045,N_7860,N_6419);
xnor U10046 (N_10046,N_8687,N_7971);
and U10047 (N_10047,N_6990,N_6895);
nand U10048 (N_10048,N_8552,N_7395);
or U10049 (N_10049,N_6916,N_8525);
nor U10050 (N_10050,N_6774,N_6629);
nor U10051 (N_10051,N_8148,N_7645);
nor U10052 (N_10052,N_7170,N_7808);
or U10053 (N_10053,N_8851,N_6798);
nand U10054 (N_10054,N_7069,N_6338);
nor U10055 (N_10055,N_6688,N_6835);
and U10056 (N_10056,N_8367,N_7941);
or U10057 (N_10057,N_6104,N_6234);
xnor U10058 (N_10058,N_7312,N_6423);
nor U10059 (N_10059,N_6354,N_8971);
and U10060 (N_10060,N_6566,N_8197);
and U10061 (N_10061,N_8794,N_6722);
and U10062 (N_10062,N_7988,N_7893);
and U10063 (N_10063,N_8698,N_8476);
nand U10064 (N_10064,N_8025,N_8210);
or U10065 (N_10065,N_6742,N_7891);
nand U10066 (N_10066,N_8343,N_7369);
nor U10067 (N_10067,N_6111,N_6333);
nand U10068 (N_10068,N_6261,N_8586);
and U10069 (N_10069,N_6823,N_6238);
nand U10070 (N_10070,N_6124,N_7172);
or U10071 (N_10071,N_7781,N_7403);
or U10072 (N_10072,N_7158,N_8758);
nor U10073 (N_10073,N_8272,N_7285);
nand U10074 (N_10074,N_8295,N_6840);
or U10075 (N_10075,N_6231,N_7884);
nor U10076 (N_10076,N_8463,N_8543);
and U10077 (N_10077,N_6130,N_8917);
xor U10078 (N_10078,N_8226,N_8149);
or U10079 (N_10079,N_7628,N_8445);
nand U10080 (N_10080,N_8048,N_7972);
or U10081 (N_10081,N_8301,N_6237);
and U10082 (N_10082,N_7364,N_6655);
or U10083 (N_10083,N_6795,N_6754);
nor U10084 (N_10084,N_7096,N_6327);
or U10085 (N_10085,N_8731,N_8843);
nand U10086 (N_10086,N_6987,N_6656);
nor U10087 (N_10087,N_6922,N_7882);
or U10088 (N_10088,N_7790,N_7194);
or U10089 (N_10089,N_8714,N_6131);
nor U10090 (N_10090,N_8334,N_6732);
nand U10091 (N_10091,N_8885,N_7589);
or U10092 (N_10092,N_8560,N_8360);
nor U10093 (N_10093,N_8392,N_6256);
or U10094 (N_10094,N_8998,N_8032);
nor U10095 (N_10095,N_7169,N_8604);
nand U10096 (N_10096,N_7743,N_7705);
nand U10097 (N_10097,N_8085,N_7015);
nand U10098 (N_10098,N_8759,N_8645);
nor U10099 (N_10099,N_6477,N_8058);
or U10100 (N_10100,N_8943,N_8260);
nand U10101 (N_10101,N_8494,N_6671);
and U10102 (N_10102,N_6520,N_6507);
and U10103 (N_10103,N_7526,N_8764);
xor U10104 (N_10104,N_8274,N_6258);
or U10105 (N_10105,N_6609,N_6011);
nand U10106 (N_10106,N_7954,N_6844);
or U10107 (N_10107,N_6356,N_8044);
and U10108 (N_10108,N_8942,N_8142);
nor U10109 (N_10109,N_6859,N_6316);
nor U10110 (N_10110,N_7371,N_7039);
nand U10111 (N_10111,N_7939,N_6165);
xnor U10112 (N_10112,N_8021,N_7772);
nand U10113 (N_10113,N_6439,N_8944);
nor U10114 (N_10114,N_6573,N_8708);
or U10115 (N_10115,N_7106,N_8243);
nor U10116 (N_10116,N_7752,N_8762);
and U10117 (N_10117,N_6509,N_6642);
and U10118 (N_10118,N_8232,N_6545);
nor U10119 (N_10119,N_8348,N_7235);
or U10120 (N_10120,N_7841,N_8902);
nand U10121 (N_10121,N_8307,N_8666);
nor U10122 (N_10122,N_8616,N_6223);
or U10123 (N_10123,N_8067,N_6052);
nor U10124 (N_10124,N_8955,N_7164);
nand U10125 (N_10125,N_6617,N_6030);
and U10126 (N_10126,N_7991,N_6801);
or U10127 (N_10127,N_7386,N_6048);
nor U10128 (N_10128,N_8713,N_6013);
nor U10129 (N_10129,N_6073,N_7756);
nand U10130 (N_10130,N_6120,N_7217);
and U10131 (N_10131,N_8104,N_8860);
and U10132 (N_10132,N_8517,N_6849);
xnor U10133 (N_10133,N_8546,N_8876);
nand U10134 (N_10134,N_8936,N_6775);
or U10135 (N_10135,N_7446,N_7846);
or U10136 (N_10136,N_8426,N_6746);
or U10137 (N_10137,N_6542,N_7009);
or U10138 (N_10138,N_6357,N_7799);
nand U10139 (N_10139,N_7601,N_8852);
nand U10140 (N_10140,N_6404,N_6473);
and U10141 (N_10141,N_6086,N_7850);
or U10142 (N_10142,N_8643,N_6370);
nand U10143 (N_10143,N_6118,N_8862);
or U10144 (N_10144,N_7964,N_8839);
and U10145 (N_10145,N_8811,N_7614);
and U10146 (N_10146,N_8417,N_8231);
nor U10147 (N_10147,N_6041,N_6865);
nand U10148 (N_10148,N_8857,N_8416);
nand U10149 (N_10149,N_8820,N_8590);
and U10150 (N_10150,N_7688,N_6611);
nor U10151 (N_10151,N_8638,N_8686);
and U10152 (N_10152,N_7758,N_7246);
or U10153 (N_10153,N_7330,N_8739);
or U10154 (N_10154,N_7679,N_6384);
nand U10155 (N_10155,N_6277,N_6690);
nand U10156 (N_10156,N_7472,N_7814);
nand U10157 (N_10157,N_6266,N_7248);
nand U10158 (N_10158,N_7493,N_8784);
xnor U10159 (N_10159,N_7574,N_6925);
nand U10160 (N_10160,N_6760,N_6080);
nor U10161 (N_10161,N_7870,N_7858);
and U10162 (N_10162,N_8068,N_7290);
or U10163 (N_10163,N_8095,N_7292);
xor U10164 (N_10164,N_7522,N_8556);
nand U10165 (N_10165,N_7603,N_8268);
and U10166 (N_10166,N_8984,N_6366);
or U10167 (N_10167,N_6820,N_8178);
nor U10168 (N_10168,N_7606,N_7986);
or U10169 (N_10169,N_8496,N_6430);
and U10170 (N_10170,N_8234,N_7084);
xnor U10171 (N_10171,N_6684,N_8625);
nand U10172 (N_10172,N_7362,N_6923);
nand U10173 (N_10173,N_7436,N_8856);
nor U10174 (N_10174,N_8807,N_8797);
nor U10175 (N_10175,N_8346,N_6229);
and U10176 (N_10176,N_8333,N_6479);
nand U10177 (N_10177,N_7598,N_6127);
and U10178 (N_10178,N_7151,N_6434);
nor U10179 (N_10179,N_7963,N_7501);
or U10180 (N_10180,N_8674,N_6198);
nor U10181 (N_10181,N_7304,N_7817);
or U10182 (N_10182,N_8011,N_6887);
nor U10183 (N_10183,N_7836,N_6810);
and U10184 (N_10184,N_8242,N_8265);
nand U10185 (N_10185,N_8780,N_6860);
and U10186 (N_10186,N_6813,N_6620);
nand U10187 (N_10187,N_6693,N_6521);
nor U10188 (N_10188,N_7978,N_6972);
nor U10189 (N_10189,N_7699,N_6436);
or U10190 (N_10190,N_7634,N_8203);
or U10191 (N_10191,N_8594,N_8409);
or U10192 (N_10192,N_8216,N_6868);
nand U10193 (N_10193,N_6714,N_8500);
nor U10194 (N_10194,N_6203,N_6153);
nor U10195 (N_10195,N_7061,N_6270);
or U10196 (N_10196,N_7175,N_6344);
nor U10197 (N_10197,N_8720,N_6959);
and U10198 (N_10198,N_7081,N_8003);
nor U10199 (N_10199,N_8763,N_6626);
and U10200 (N_10200,N_7479,N_7324);
nor U10201 (N_10201,N_8521,N_6141);
nand U10202 (N_10202,N_7365,N_7259);
or U10203 (N_10203,N_7582,N_7072);
or U10204 (N_10204,N_6275,N_6469);
nand U10205 (N_10205,N_6304,N_7748);
or U10206 (N_10206,N_7447,N_6495);
and U10207 (N_10207,N_7608,N_8116);
nand U10208 (N_10208,N_7642,N_6497);
and U10209 (N_10209,N_8182,N_6390);
and U10210 (N_10210,N_7746,N_6828);
nand U10211 (N_10211,N_6767,N_8513);
nor U10212 (N_10212,N_6847,N_7684);
nor U10213 (N_10213,N_6741,N_6347);
nor U10214 (N_10214,N_8485,N_6252);
nand U10215 (N_10215,N_8100,N_6228);
and U10216 (N_10216,N_7872,N_8727);
nand U10217 (N_10217,N_6885,N_8558);
and U10218 (N_10218,N_7174,N_7146);
nand U10219 (N_10219,N_7955,N_6108);
and U10220 (N_10220,N_7687,N_6664);
nand U10221 (N_10221,N_8323,N_7222);
or U10222 (N_10222,N_6700,N_6299);
and U10223 (N_10223,N_8953,N_6341);
nor U10224 (N_10224,N_8194,N_8939);
or U10225 (N_10225,N_8624,N_6040);
and U10226 (N_10226,N_6837,N_8248);
or U10227 (N_10227,N_8932,N_8684);
and U10228 (N_10228,N_6287,N_7432);
nand U10229 (N_10229,N_8791,N_6089);
and U10230 (N_10230,N_6552,N_8387);
or U10231 (N_10231,N_8836,N_8239);
and U10232 (N_10232,N_7581,N_8757);
nor U10233 (N_10233,N_6415,N_8658);
or U10234 (N_10234,N_7087,N_6658);
nand U10235 (N_10235,N_7769,N_7729);
nand U10236 (N_10236,N_7209,N_6337);
and U10237 (N_10237,N_8388,N_6429);
nand U10238 (N_10238,N_8250,N_6701);
nand U10239 (N_10239,N_8756,N_6519);
and U10240 (N_10240,N_6460,N_6911);
xor U10241 (N_10241,N_8524,N_7233);
nand U10242 (N_10242,N_6225,N_6110);
and U10243 (N_10243,N_7251,N_6730);
nand U10244 (N_10244,N_8466,N_7409);
nor U10245 (N_10245,N_6162,N_7717);
nand U10246 (N_10246,N_7474,N_8038);
nor U10247 (N_10247,N_7341,N_7616);
nand U10248 (N_10248,N_7709,N_8788);
nand U10249 (N_10249,N_6999,N_8853);
and U10250 (N_10250,N_8482,N_6447);
nand U10251 (N_10251,N_8669,N_8006);
nand U10252 (N_10252,N_8330,N_7597);
nand U10253 (N_10253,N_6486,N_7673);
nor U10254 (N_10254,N_7604,N_7801);
and U10255 (N_10255,N_7585,N_6236);
nand U10256 (N_10256,N_8412,N_6508);
nor U10257 (N_10257,N_8963,N_7309);
or U10258 (N_10258,N_8395,N_6387);
nor U10259 (N_10259,N_8267,N_8574);
nor U10260 (N_10260,N_8881,N_8352);
nor U10261 (N_10261,N_8859,N_6595);
or U10262 (N_10262,N_8118,N_8237);
nand U10263 (N_10263,N_6893,N_6977);
or U10264 (N_10264,N_7660,N_6364);
or U10265 (N_10265,N_8164,N_7755);
or U10266 (N_10266,N_7552,N_7851);
or U10267 (N_10267,N_7864,N_7058);
nand U10268 (N_10268,N_8483,N_7339);
nor U10269 (N_10269,N_6749,N_7843);
nor U10270 (N_10270,N_7831,N_7550);
nand U10271 (N_10271,N_7946,N_7335);
and U10272 (N_10272,N_8799,N_8632);
or U10273 (N_10273,N_7767,N_7126);
nand U10274 (N_10274,N_7612,N_6084);
or U10275 (N_10275,N_6136,N_7600);
nand U10276 (N_10276,N_7761,N_6463);
and U10277 (N_10277,N_8055,N_7197);
nand U10278 (N_10278,N_6031,N_7714);
nor U10279 (N_10279,N_6400,N_6713);
and U10280 (N_10280,N_8340,N_8982);
nand U10281 (N_10281,N_6440,N_7837);
nand U10282 (N_10282,N_7450,N_8140);
nor U10283 (N_10283,N_7757,N_8049);
xor U10284 (N_10284,N_7012,N_7813);
nand U10285 (N_10285,N_7947,N_7742);
and U10286 (N_10286,N_6119,N_6175);
xor U10287 (N_10287,N_8266,N_7071);
nand U10288 (N_10288,N_8569,N_8005);
nand U10289 (N_10289,N_7407,N_7243);
nand U10290 (N_10290,N_6672,N_7656);
xnor U10291 (N_10291,N_8728,N_6838);
or U10292 (N_10292,N_8696,N_8499);
xnor U10293 (N_10293,N_8462,N_7098);
or U10294 (N_10294,N_6379,N_7396);
xor U10295 (N_10295,N_6863,N_8399);
nand U10296 (N_10296,N_6695,N_6558);
nor U10297 (N_10297,N_7647,N_8877);
and U10298 (N_10298,N_8350,N_7666);
or U10299 (N_10299,N_8251,N_8147);
or U10300 (N_10300,N_7990,N_6279);
and U10301 (N_10301,N_7405,N_6805);
nor U10302 (N_10302,N_7477,N_6678);
nand U10303 (N_10303,N_6016,N_7091);
xnor U10304 (N_10304,N_6992,N_6694);
nor U10305 (N_10305,N_8835,N_7462);
or U10306 (N_10306,N_7346,N_8154);
nor U10307 (N_10307,N_7923,N_8007);
and U10308 (N_10308,N_7797,N_7838);
nand U10309 (N_10309,N_6564,N_6808);
nor U10310 (N_10310,N_6200,N_6889);
or U10311 (N_10311,N_8957,N_8715);
nand U10312 (N_10312,N_7800,N_6001);
nand U10313 (N_10313,N_7771,N_7678);
or U10314 (N_10314,N_8886,N_7094);
or U10315 (N_10315,N_7198,N_6302);
nand U10316 (N_10316,N_6894,N_8143);
and U10317 (N_10317,N_6913,N_6156);
nor U10318 (N_10318,N_8571,N_6487);
nor U10319 (N_10319,N_8626,N_6301);
nand U10320 (N_10320,N_7788,N_8444);
nand U10321 (N_10321,N_7267,N_7496);
or U10322 (N_10322,N_8760,N_8042);
xnor U10323 (N_10323,N_7948,N_7898);
nand U10324 (N_10324,N_8879,N_7426);
nor U10325 (N_10325,N_8484,N_8609);
and U10326 (N_10326,N_8628,N_8751);
or U10327 (N_10327,N_8489,N_8933);
nand U10328 (N_10328,N_7933,N_7204);
and U10329 (N_10329,N_6257,N_6325);
nor U10330 (N_10330,N_7768,N_8033);
or U10331 (N_10331,N_7806,N_6522);
xnor U10332 (N_10332,N_7627,N_6662);
and U10333 (N_10333,N_7503,N_8238);
nand U10334 (N_10334,N_7064,N_8355);
or U10335 (N_10335,N_6866,N_8980);
and U10336 (N_10336,N_8979,N_6833);
or U10337 (N_10337,N_8128,N_7121);
or U10338 (N_10338,N_7100,N_7512);
nor U10339 (N_10339,N_7588,N_7524);
nand U10340 (N_10340,N_6921,N_7957);
and U10341 (N_10341,N_7563,N_6574);
nand U10342 (N_10342,N_8926,N_8920);
or U10343 (N_10343,N_8368,N_8830);
and U10344 (N_10344,N_7833,N_8742);
nand U10345 (N_10345,N_7397,N_7855);
and U10346 (N_10346,N_7077,N_8075);
and U10347 (N_10347,N_8390,N_6842);
nor U10348 (N_10348,N_6884,N_8441);
and U10349 (N_10349,N_6931,N_7792);
nor U10350 (N_10350,N_7112,N_7471);
nor U10351 (N_10351,N_6003,N_8303);
nor U10352 (N_10352,N_6027,N_6365);
xnor U10353 (N_10353,N_6389,N_6432);
nand U10354 (N_10354,N_7130,N_6613);
and U10355 (N_10355,N_6271,N_6446);
nor U10356 (N_10356,N_7202,N_8397);
nand U10357 (N_10357,N_6241,N_8723);
nor U10358 (N_10358,N_6633,N_6981);
or U10359 (N_10359,N_8325,N_7599);
nand U10360 (N_10360,N_7326,N_7545);
and U10361 (N_10361,N_7385,N_6673);
or U10362 (N_10362,N_8461,N_6176);
and U10363 (N_10363,N_7473,N_6902);
and U10364 (N_10364,N_7498,N_7510);
xnor U10365 (N_10365,N_8335,N_8894);
and U10366 (N_10366,N_8062,N_6606);
or U10367 (N_10367,N_8749,N_6475);
nand U10368 (N_10368,N_7334,N_8819);
and U10369 (N_10369,N_6079,N_7651);
nand U10370 (N_10370,N_7051,N_6043);
and U10371 (N_10371,N_8230,N_7966);
nor U10372 (N_10372,N_8079,N_8966);
or U10373 (N_10373,N_6103,N_7161);
nor U10374 (N_10374,N_8318,N_8404);
nand U10375 (N_10375,N_6248,N_7974);
xor U10376 (N_10376,N_8487,N_7104);
and U10377 (N_10377,N_7428,N_7848);
nor U10378 (N_10378,N_6441,N_6038);
or U10379 (N_10379,N_8637,N_6438);
nand U10380 (N_10380,N_7530,N_6409);
nand U10381 (N_10381,N_8538,N_8136);
nor U10382 (N_10382,N_6716,N_7718);
nor U10383 (N_10383,N_6822,N_6044);
or U10384 (N_10384,N_6934,N_6422);
or U10385 (N_10385,N_8912,N_7734);
nand U10386 (N_10386,N_6306,N_7054);
or U10387 (N_10387,N_7919,N_8206);
nand U10388 (N_10388,N_7070,N_6514);
nor U10389 (N_10389,N_6491,N_8030);
and U10390 (N_10390,N_7483,N_7258);
nand U10391 (N_10391,N_8603,N_8640);
nor U10392 (N_10392,N_8211,N_6964);
or U10393 (N_10393,N_8771,N_6788);
or U10394 (N_10394,N_8798,N_8722);
nand U10395 (N_10395,N_6375,N_6076);
and U10396 (N_10396,N_6293,N_8029);
or U10397 (N_10397,N_7270,N_6622);
or U10398 (N_10398,N_7110,N_6067);
or U10399 (N_10399,N_8801,N_6577);
or U10400 (N_10400,N_8868,N_7511);
nand U10401 (N_10401,N_8057,N_6586);
nor U10402 (N_10402,N_7967,N_7565);
nor U10403 (N_10403,N_6247,N_7320);
and U10404 (N_10404,N_8847,N_6739);
or U10405 (N_10405,N_8026,N_8913);
nand U10406 (N_10406,N_8657,N_6006);
nor U10407 (N_10407,N_7414,N_7234);
or U10408 (N_10408,N_6420,N_7541);
nor U10409 (N_10409,N_8593,N_6395);
or U10410 (N_10410,N_7296,N_6745);
or U10411 (N_10411,N_6848,N_7023);
or U10412 (N_10412,N_6727,N_7844);
nand U10413 (N_10413,N_6368,N_6686);
nand U10414 (N_10414,N_7220,N_7136);
nand U10415 (N_10415,N_7244,N_6335);
or U10416 (N_10416,N_8134,N_7374);
or U10417 (N_10417,N_7514,N_8952);
or U10418 (N_10418,N_7625,N_6227);
nand U10419 (N_10419,N_8701,N_6411);
nor U10420 (N_10420,N_7847,N_8985);
nand U10421 (N_10421,N_6207,N_6443);
nor U10422 (N_10422,N_6669,N_7486);
or U10423 (N_10423,N_8961,N_6313);
and U10424 (N_10424,N_7314,N_7008);
nand U10425 (N_10425,N_8930,N_6224);
or U10426 (N_10426,N_8949,N_6493);
nor U10427 (N_10427,N_8767,N_6515);
nand U10428 (N_10428,N_8374,N_8064);
or U10429 (N_10429,N_7969,N_6983);
nor U10430 (N_10430,N_7056,N_6026);
or U10431 (N_10431,N_8746,N_8401);
and U10432 (N_10432,N_7333,N_6050);
xnor U10433 (N_10433,N_8873,N_6874);
or U10434 (N_10434,N_6903,N_7897);
or U10435 (N_10435,N_7179,N_7566);
nor U10436 (N_10436,N_8117,N_8129);
nand U10437 (N_10437,N_6630,N_6904);
and U10438 (N_10438,N_7303,N_6081);
or U10439 (N_10439,N_6385,N_8382);
and U10440 (N_10440,N_7160,N_6189);
nand U10441 (N_10441,N_8362,N_8540);
nand U10442 (N_10442,N_8102,N_6372);
nor U10443 (N_10443,N_7953,N_8403);
nand U10444 (N_10444,N_7016,N_6575);
and U10445 (N_10445,N_7856,N_7573);
nand U10446 (N_10446,N_7082,N_6173);
or U10447 (N_10447,N_6557,N_8692);
nor U10448 (N_10448,N_6940,N_7615);
and U10449 (N_10449,N_8037,N_7441);
nor U10450 (N_10450,N_6021,N_7144);
nand U10451 (N_10451,N_7276,N_6588);
nand U10452 (N_10452,N_7289,N_6183);
and U10453 (N_10453,N_8087,N_6791);
nor U10454 (N_10454,N_8073,N_8119);
or U10455 (N_10455,N_8337,N_8534);
and U10456 (N_10456,N_6827,N_6047);
nor U10457 (N_10457,N_7424,N_7620);
nand U10458 (N_10458,N_7480,N_6710);
nand U10459 (N_10459,N_8344,N_6164);
nand U10460 (N_10460,N_8972,N_6504);
or U10461 (N_10461,N_7375,N_6615);
nand U10462 (N_10462,N_8327,N_6661);
nand U10463 (N_10463,N_6246,N_8832);
nand U10464 (N_10464,N_7192,N_7468);
or U10465 (N_10465,N_8884,N_8809);
nor U10466 (N_10466,N_6970,N_6816);
nor U10467 (N_10467,N_6587,N_6010);
and U10468 (N_10468,N_7713,N_6955);
nor U10469 (N_10469,N_8187,N_6607);
or U10470 (N_10470,N_6703,N_8423);
and U10471 (N_10471,N_8400,N_7804);
and U10472 (N_10472,N_7305,N_7318);
nor U10473 (N_10473,N_7877,N_8249);
and U10474 (N_10474,N_7492,N_7629);
and U10475 (N_10475,N_7119,N_7109);
nor U10476 (N_10476,N_6989,N_7704);
nand U10477 (N_10477,N_6961,N_8008);
nand U10478 (N_10478,N_6051,N_7903);
or U10479 (N_10479,N_8255,N_6291);
or U10480 (N_10480,N_7307,N_6166);
and U10481 (N_10481,N_7090,N_6829);
or U10482 (N_10482,N_7103,N_7763);
or U10483 (N_10483,N_7302,N_8430);
nand U10484 (N_10484,N_7516,N_8459);
nand U10485 (N_10485,N_7360,N_8880);
or U10486 (N_10486,N_8565,N_7866);
or U10487 (N_10487,N_6092,N_7412);
nand U10488 (N_10488,N_7200,N_6632);
or U10489 (N_10489,N_8765,N_7555);
or U10490 (N_10490,N_6253,N_7122);
and U10491 (N_10491,N_6053,N_8432);
nor U10492 (N_10492,N_6037,N_7928);
and U10493 (N_10493,N_7242,N_8796);
nand U10494 (N_10494,N_7636,N_8600);
nand U10495 (N_10495,N_7253,N_6331);
and U10496 (N_10496,N_8921,N_8391);
nand U10497 (N_10497,N_6665,N_8748);
or U10498 (N_10498,N_8358,N_6481);
nand U10499 (N_10499,N_8319,N_6723);
or U10500 (N_10500,N_8405,N_8878);
nor U10501 (N_10501,N_8062,N_6535);
or U10502 (N_10502,N_6706,N_7565);
and U10503 (N_10503,N_7690,N_7446);
and U10504 (N_10504,N_6775,N_8416);
or U10505 (N_10505,N_6184,N_7973);
or U10506 (N_10506,N_6116,N_8007);
and U10507 (N_10507,N_7060,N_7896);
or U10508 (N_10508,N_8827,N_7243);
nand U10509 (N_10509,N_7051,N_6141);
and U10510 (N_10510,N_7446,N_7764);
xnor U10511 (N_10511,N_7878,N_8614);
or U10512 (N_10512,N_6096,N_8227);
nor U10513 (N_10513,N_6753,N_6262);
and U10514 (N_10514,N_8698,N_8882);
nor U10515 (N_10515,N_8198,N_7197);
and U10516 (N_10516,N_6986,N_6359);
and U10517 (N_10517,N_6667,N_6367);
and U10518 (N_10518,N_8104,N_7359);
nor U10519 (N_10519,N_7374,N_7781);
or U10520 (N_10520,N_7292,N_7195);
and U10521 (N_10521,N_6539,N_7066);
nand U10522 (N_10522,N_7589,N_7134);
nor U10523 (N_10523,N_8788,N_6424);
and U10524 (N_10524,N_8696,N_8629);
nand U10525 (N_10525,N_8156,N_7787);
and U10526 (N_10526,N_8732,N_8073);
nor U10527 (N_10527,N_7863,N_6622);
and U10528 (N_10528,N_8840,N_8904);
and U10529 (N_10529,N_6282,N_8239);
and U10530 (N_10530,N_7024,N_6135);
and U10531 (N_10531,N_8186,N_7836);
nor U10532 (N_10532,N_8654,N_7381);
and U10533 (N_10533,N_7229,N_7994);
and U10534 (N_10534,N_6602,N_6296);
and U10535 (N_10535,N_7488,N_6693);
or U10536 (N_10536,N_8452,N_6584);
nand U10537 (N_10537,N_8908,N_6979);
nand U10538 (N_10538,N_6917,N_8523);
and U10539 (N_10539,N_7359,N_6360);
nor U10540 (N_10540,N_7891,N_8558);
and U10541 (N_10541,N_6028,N_7669);
xnor U10542 (N_10542,N_8343,N_6416);
or U10543 (N_10543,N_6436,N_8314);
nand U10544 (N_10544,N_6180,N_8898);
and U10545 (N_10545,N_7002,N_8160);
nor U10546 (N_10546,N_8563,N_8971);
and U10547 (N_10547,N_7193,N_7961);
nand U10548 (N_10548,N_7071,N_8368);
or U10549 (N_10549,N_7497,N_8322);
or U10550 (N_10550,N_7930,N_8335);
nand U10551 (N_10551,N_7779,N_6298);
or U10552 (N_10552,N_8663,N_7392);
or U10553 (N_10553,N_8129,N_6983);
or U10554 (N_10554,N_7723,N_7773);
nor U10555 (N_10555,N_7242,N_8501);
and U10556 (N_10556,N_7000,N_6502);
nand U10557 (N_10557,N_6277,N_8407);
and U10558 (N_10558,N_6240,N_8768);
nand U10559 (N_10559,N_6478,N_8989);
nand U10560 (N_10560,N_7941,N_7820);
or U10561 (N_10561,N_8806,N_8973);
or U10562 (N_10562,N_8019,N_7123);
or U10563 (N_10563,N_7511,N_8427);
or U10564 (N_10564,N_6373,N_7006);
nor U10565 (N_10565,N_6078,N_7698);
nor U10566 (N_10566,N_6188,N_6727);
xnor U10567 (N_10567,N_7432,N_6588);
or U10568 (N_10568,N_8917,N_8704);
and U10569 (N_10569,N_8749,N_6733);
nor U10570 (N_10570,N_6610,N_6339);
or U10571 (N_10571,N_8224,N_8666);
and U10572 (N_10572,N_7871,N_7196);
and U10573 (N_10573,N_7881,N_6734);
nand U10574 (N_10574,N_6448,N_8733);
or U10575 (N_10575,N_8104,N_6102);
and U10576 (N_10576,N_6993,N_7192);
or U10577 (N_10577,N_8253,N_8769);
nand U10578 (N_10578,N_6619,N_8705);
nand U10579 (N_10579,N_7371,N_6137);
nand U10580 (N_10580,N_7026,N_8768);
or U10581 (N_10581,N_7581,N_6718);
nand U10582 (N_10582,N_6372,N_6263);
and U10583 (N_10583,N_7777,N_6910);
nand U10584 (N_10584,N_7749,N_7998);
and U10585 (N_10585,N_6157,N_8612);
nor U10586 (N_10586,N_6938,N_6572);
and U10587 (N_10587,N_6404,N_6436);
or U10588 (N_10588,N_7640,N_7162);
nor U10589 (N_10589,N_7915,N_7664);
and U10590 (N_10590,N_7237,N_7920);
or U10591 (N_10591,N_7729,N_8588);
or U10592 (N_10592,N_7866,N_7256);
and U10593 (N_10593,N_6253,N_7527);
or U10594 (N_10594,N_6536,N_7622);
and U10595 (N_10595,N_7394,N_6335);
nand U10596 (N_10596,N_7086,N_8655);
or U10597 (N_10597,N_8369,N_7631);
nor U10598 (N_10598,N_6852,N_7564);
or U10599 (N_10599,N_6537,N_6674);
and U10600 (N_10600,N_8573,N_6712);
nor U10601 (N_10601,N_6884,N_6531);
or U10602 (N_10602,N_6117,N_8140);
or U10603 (N_10603,N_8031,N_6679);
nor U10604 (N_10604,N_7714,N_7935);
and U10605 (N_10605,N_6575,N_6505);
and U10606 (N_10606,N_6530,N_7312);
and U10607 (N_10607,N_6797,N_6981);
or U10608 (N_10608,N_8289,N_8923);
or U10609 (N_10609,N_7530,N_8877);
or U10610 (N_10610,N_8108,N_8156);
nand U10611 (N_10611,N_8836,N_6285);
nand U10612 (N_10612,N_8061,N_7613);
or U10613 (N_10613,N_8349,N_6078);
and U10614 (N_10614,N_7185,N_8015);
nand U10615 (N_10615,N_6666,N_7713);
nor U10616 (N_10616,N_7350,N_7258);
xor U10617 (N_10617,N_7072,N_6273);
nand U10618 (N_10618,N_7311,N_6425);
or U10619 (N_10619,N_8407,N_6635);
nor U10620 (N_10620,N_8214,N_6951);
or U10621 (N_10621,N_6119,N_8016);
and U10622 (N_10622,N_6440,N_7885);
nor U10623 (N_10623,N_6255,N_8262);
or U10624 (N_10624,N_8608,N_8282);
nand U10625 (N_10625,N_8126,N_6796);
nor U10626 (N_10626,N_8862,N_6653);
nor U10627 (N_10627,N_6285,N_8918);
nand U10628 (N_10628,N_6970,N_7006);
xor U10629 (N_10629,N_8811,N_6085);
and U10630 (N_10630,N_6674,N_6494);
and U10631 (N_10631,N_7836,N_6862);
nand U10632 (N_10632,N_6692,N_6562);
nand U10633 (N_10633,N_7223,N_8438);
or U10634 (N_10634,N_8939,N_7756);
or U10635 (N_10635,N_7228,N_7879);
or U10636 (N_10636,N_6825,N_6822);
nor U10637 (N_10637,N_7752,N_8055);
and U10638 (N_10638,N_7709,N_8185);
nand U10639 (N_10639,N_6498,N_7758);
and U10640 (N_10640,N_6251,N_6246);
and U10641 (N_10641,N_8264,N_7097);
nor U10642 (N_10642,N_8291,N_7802);
and U10643 (N_10643,N_6166,N_8680);
nand U10644 (N_10644,N_8769,N_8109);
nand U10645 (N_10645,N_7730,N_8214);
or U10646 (N_10646,N_6753,N_8667);
or U10647 (N_10647,N_8335,N_8434);
or U10648 (N_10648,N_6641,N_6006);
and U10649 (N_10649,N_6716,N_7129);
nor U10650 (N_10650,N_7694,N_7796);
or U10651 (N_10651,N_6726,N_6847);
and U10652 (N_10652,N_7997,N_6054);
and U10653 (N_10653,N_6107,N_8880);
nor U10654 (N_10654,N_6288,N_6978);
xor U10655 (N_10655,N_8579,N_8096);
or U10656 (N_10656,N_7566,N_7156);
and U10657 (N_10657,N_8657,N_7947);
or U10658 (N_10658,N_7888,N_8069);
and U10659 (N_10659,N_6849,N_7123);
nand U10660 (N_10660,N_7368,N_6085);
and U10661 (N_10661,N_6071,N_8235);
nor U10662 (N_10662,N_8160,N_8395);
nand U10663 (N_10663,N_6734,N_6232);
or U10664 (N_10664,N_7282,N_7773);
nand U10665 (N_10665,N_7167,N_8759);
nand U10666 (N_10666,N_6655,N_6450);
nor U10667 (N_10667,N_6453,N_8109);
nand U10668 (N_10668,N_8605,N_6461);
or U10669 (N_10669,N_8005,N_7084);
nor U10670 (N_10670,N_6465,N_7903);
nor U10671 (N_10671,N_6331,N_8918);
nor U10672 (N_10672,N_8136,N_7473);
or U10673 (N_10673,N_8192,N_8163);
nor U10674 (N_10674,N_6186,N_8808);
and U10675 (N_10675,N_6857,N_7593);
or U10676 (N_10676,N_6149,N_6213);
nand U10677 (N_10677,N_7389,N_6662);
and U10678 (N_10678,N_7948,N_6220);
or U10679 (N_10679,N_6772,N_8557);
nand U10680 (N_10680,N_6472,N_6389);
or U10681 (N_10681,N_8918,N_6609);
and U10682 (N_10682,N_6350,N_6064);
nand U10683 (N_10683,N_6778,N_8444);
nand U10684 (N_10684,N_7937,N_6022);
nand U10685 (N_10685,N_8276,N_8996);
nor U10686 (N_10686,N_6634,N_7705);
and U10687 (N_10687,N_8891,N_6625);
nor U10688 (N_10688,N_8028,N_6664);
and U10689 (N_10689,N_7612,N_7811);
and U10690 (N_10690,N_6554,N_8210);
and U10691 (N_10691,N_7094,N_7913);
or U10692 (N_10692,N_6702,N_8616);
nor U10693 (N_10693,N_6595,N_6530);
nand U10694 (N_10694,N_6287,N_6039);
and U10695 (N_10695,N_6937,N_7828);
or U10696 (N_10696,N_7894,N_6001);
and U10697 (N_10697,N_7663,N_6592);
nor U10698 (N_10698,N_7226,N_6178);
nand U10699 (N_10699,N_6602,N_7414);
nand U10700 (N_10700,N_7659,N_7938);
and U10701 (N_10701,N_8554,N_7737);
xnor U10702 (N_10702,N_7986,N_6723);
and U10703 (N_10703,N_6857,N_8623);
or U10704 (N_10704,N_7490,N_7123);
nor U10705 (N_10705,N_8464,N_7351);
nor U10706 (N_10706,N_7377,N_7016);
or U10707 (N_10707,N_8923,N_6899);
nand U10708 (N_10708,N_8095,N_8096);
and U10709 (N_10709,N_7253,N_7452);
or U10710 (N_10710,N_6692,N_6667);
and U10711 (N_10711,N_7478,N_7484);
nor U10712 (N_10712,N_8865,N_7876);
or U10713 (N_10713,N_8547,N_7513);
nand U10714 (N_10714,N_8342,N_6828);
and U10715 (N_10715,N_6022,N_6168);
nor U10716 (N_10716,N_6263,N_6046);
xor U10717 (N_10717,N_7846,N_7553);
nor U10718 (N_10718,N_8998,N_8004);
nor U10719 (N_10719,N_6204,N_7723);
and U10720 (N_10720,N_7691,N_7660);
nor U10721 (N_10721,N_6886,N_7628);
nor U10722 (N_10722,N_6778,N_6668);
nor U10723 (N_10723,N_7981,N_7821);
nor U10724 (N_10724,N_6403,N_6147);
and U10725 (N_10725,N_6706,N_7620);
or U10726 (N_10726,N_7723,N_7328);
nand U10727 (N_10727,N_7482,N_6692);
nand U10728 (N_10728,N_7761,N_6400);
nor U10729 (N_10729,N_7632,N_6959);
nand U10730 (N_10730,N_8921,N_6262);
xor U10731 (N_10731,N_6799,N_7487);
and U10732 (N_10732,N_7774,N_6003);
and U10733 (N_10733,N_7437,N_8861);
xnor U10734 (N_10734,N_7881,N_7589);
nand U10735 (N_10735,N_7756,N_8045);
or U10736 (N_10736,N_8039,N_8730);
nand U10737 (N_10737,N_6551,N_7248);
or U10738 (N_10738,N_6014,N_8156);
and U10739 (N_10739,N_6808,N_6191);
nand U10740 (N_10740,N_6949,N_8628);
and U10741 (N_10741,N_6649,N_7061);
nor U10742 (N_10742,N_6209,N_8771);
and U10743 (N_10743,N_6637,N_7118);
and U10744 (N_10744,N_6730,N_6764);
nand U10745 (N_10745,N_8760,N_7437);
nor U10746 (N_10746,N_7665,N_8289);
and U10747 (N_10747,N_8280,N_6692);
or U10748 (N_10748,N_6103,N_6732);
and U10749 (N_10749,N_6166,N_8707);
and U10750 (N_10750,N_6621,N_8754);
nand U10751 (N_10751,N_8986,N_7925);
nand U10752 (N_10752,N_7580,N_8381);
and U10753 (N_10753,N_6066,N_6899);
xnor U10754 (N_10754,N_7346,N_7359);
and U10755 (N_10755,N_8947,N_8495);
xor U10756 (N_10756,N_7714,N_7827);
and U10757 (N_10757,N_6986,N_6422);
nor U10758 (N_10758,N_7210,N_7236);
nor U10759 (N_10759,N_6677,N_6242);
and U10760 (N_10760,N_7542,N_6964);
or U10761 (N_10761,N_7116,N_8168);
nor U10762 (N_10762,N_6269,N_6301);
xnor U10763 (N_10763,N_8481,N_8229);
and U10764 (N_10764,N_6602,N_7437);
nor U10765 (N_10765,N_7948,N_8302);
nand U10766 (N_10766,N_7630,N_8022);
nor U10767 (N_10767,N_7393,N_8702);
or U10768 (N_10768,N_7798,N_8131);
nand U10769 (N_10769,N_7121,N_8287);
and U10770 (N_10770,N_8870,N_7691);
or U10771 (N_10771,N_8732,N_8640);
and U10772 (N_10772,N_7333,N_6965);
nor U10773 (N_10773,N_6255,N_6742);
and U10774 (N_10774,N_6514,N_6238);
or U10775 (N_10775,N_6659,N_8911);
nand U10776 (N_10776,N_6626,N_7806);
nand U10777 (N_10777,N_6172,N_8902);
or U10778 (N_10778,N_6084,N_7908);
or U10779 (N_10779,N_6891,N_6781);
nand U10780 (N_10780,N_6022,N_6950);
nand U10781 (N_10781,N_7715,N_8196);
nor U10782 (N_10782,N_6594,N_7444);
and U10783 (N_10783,N_8255,N_6459);
nand U10784 (N_10784,N_8333,N_6383);
and U10785 (N_10785,N_8762,N_6923);
or U10786 (N_10786,N_7840,N_6772);
and U10787 (N_10787,N_6499,N_8097);
and U10788 (N_10788,N_6228,N_6803);
nand U10789 (N_10789,N_6998,N_8774);
nand U10790 (N_10790,N_6253,N_8037);
nand U10791 (N_10791,N_7151,N_8342);
or U10792 (N_10792,N_7529,N_7971);
and U10793 (N_10793,N_8019,N_6766);
and U10794 (N_10794,N_8504,N_8124);
nor U10795 (N_10795,N_8995,N_8748);
or U10796 (N_10796,N_8299,N_6159);
and U10797 (N_10797,N_6064,N_8719);
and U10798 (N_10798,N_7487,N_7538);
nand U10799 (N_10799,N_6012,N_8968);
and U10800 (N_10800,N_6393,N_7568);
nor U10801 (N_10801,N_6253,N_6861);
or U10802 (N_10802,N_6284,N_8689);
nand U10803 (N_10803,N_6589,N_8474);
nand U10804 (N_10804,N_7583,N_6041);
or U10805 (N_10805,N_7679,N_6044);
and U10806 (N_10806,N_7637,N_7078);
nor U10807 (N_10807,N_7239,N_8431);
or U10808 (N_10808,N_7923,N_8321);
nand U10809 (N_10809,N_6243,N_6246);
and U10810 (N_10810,N_6787,N_7674);
or U10811 (N_10811,N_6498,N_6885);
nand U10812 (N_10812,N_6621,N_8807);
nand U10813 (N_10813,N_8886,N_8623);
nor U10814 (N_10814,N_8654,N_7910);
nor U10815 (N_10815,N_6739,N_8677);
or U10816 (N_10816,N_8177,N_7565);
nor U10817 (N_10817,N_7142,N_6298);
nand U10818 (N_10818,N_7154,N_7968);
or U10819 (N_10819,N_6577,N_8400);
nor U10820 (N_10820,N_7366,N_7709);
nand U10821 (N_10821,N_8610,N_8737);
and U10822 (N_10822,N_8040,N_8517);
or U10823 (N_10823,N_7686,N_7040);
nand U10824 (N_10824,N_7359,N_8085);
nor U10825 (N_10825,N_7788,N_8803);
or U10826 (N_10826,N_8474,N_6068);
nand U10827 (N_10827,N_8874,N_8986);
nor U10828 (N_10828,N_8706,N_8927);
or U10829 (N_10829,N_7250,N_7888);
and U10830 (N_10830,N_8872,N_6990);
nand U10831 (N_10831,N_7083,N_6922);
or U10832 (N_10832,N_8497,N_8486);
and U10833 (N_10833,N_7223,N_8197);
and U10834 (N_10834,N_6291,N_7561);
nand U10835 (N_10835,N_7308,N_8873);
nand U10836 (N_10836,N_7595,N_8258);
nor U10837 (N_10837,N_6675,N_6917);
and U10838 (N_10838,N_8796,N_7892);
or U10839 (N_10839,N_8252,N_7291);
nand U10840 (N_10840,N_6045,N_6600);
and U10841 (N_10841,N_8705,N_8516);
and U10842 (N_10842,N_7597,N_7329);
nor U10843 (N_10843,N_7408,N_6841);
or U10844 (N_10844,N_8706,N_8318);
or U10845 (N_10845,N_6018,N_6086);
and U10846 (N_10846,N_8607,N_8799);
nand U10847 (N_10847,N_7088,N_8759);
and U10848 (N_10848,N_6041,N_7724);
or U10849 (N_10849,N_6433,N_6556);
or U10850 (N_10850,N_8094,N_6644);
and U10851 (N_10851,N_7776,N_8954);
and U10852 (N_10852,N_6013,N_6465);
nor U10853 (N_10853,N_6561,N_6866);
and U10854 (N_10854,N_8935,N_6135);
nor U10855 (N_10855,N_7894,N_8257);
nand U10856 (N_10856,N_8635,N_6297);
and U10857 (N_10857,N_6641,N_7700);
nor U10858 (N_10858,N_8468,N_6365);
nand U10859 (N_10859,N_6016,N_6106);
and U10860 (N_10860,N_8936,N_6442);
or U10861 (N_10861,N_8125,N_6933);
nor U10862 (N_10862,N_6462,N_6268);
or U10863 (N_10863,N_8397,N_6706);
and U10864 (N_10864,N_6782,N_6056);
and U10865 (N_10865,N_8972,N_8577);
or U10866 (N_10866,N_8839,N_6481);
or U10867 (N_10867,N_8408,N_6174);
nor U10868 (N_10868,N_8994,N_8877);
and U10869 (N_10869,N_6517,N_7135);
nand U10870 (N_10870,N_8344,N_7957);
and U10871 (N_10871,N_8673,N_6763);
or U10872 (N_10872,N_8749,N_8807);
and U10873 (N_10873,N_6797,N_6952);
and U10874 (N_10874,N_6971,N_7329);
and U10875 (N_10875,N_6684,N_8438);
or U10876 (N_10876,N_7729,N_8524);
nand U10877 (N_10877,N_8557,N_7789);
or U10878 (N_10878,N_8979,N_7371);
or U10879 (N_10879,N_8833,N_6487);
and U10880 (N_10880,N_7434,N_8223);
or U10881 (N_10881,N_8681,N_7962);
nand U10882 (N_10882,N_6268,N_6200);
nand U10883 (N_10883,N_6064,N_7236);
nor U10884 (N_10884,N_7132,N_6090);
nand U10885 (N_10885,N_7030,N_8258);
nand U10886 (N_10886,N_6455,N_8593);
and U10887 (N_10887,N_8223,N_7656);
or U10888 (N_10888,N_8432,N_6671);
or U10889 (N_10889,N_8584,N_6926);
nor U10890 (N_10890,N_8545,N_8540);
or U10891 (N_10891,N_7484,N_6479);
or U10892 (N_10892,N_8619,N_7746);
xor U10893 (N_10893,N_8707,N_6926);
or U10894 (N_10894,N_6453,N_8313);
nor U10895 (N_10895,N_8595,N_6725);
or U10896 (N_10896,N_6239,N_7181);
nor U10897 (N_10897,N_8575,N_8619);
or U10898 (N_10898,N_8899,N_8988);
or U10899 (N_10899,N_6463,N_8077);
nor U10900 (N_10900,N_8861,N_6817);
nor U10901 (N_10901,N_8035,N_7991);
or U10902 (N_10902,N_8717,N_8025);
nor U10903 (N_10903,N_6058,N_6628);
nor U10904 (N_10904,N_7244,N_7653);
xor U10905 (N_10905,N_6347,N_6535);
and U10906 (N_10906,N_6421,N_8717);
or U10907 (N_10907,N_8491,N_8677);
or U10908 (N_10908,N_7239,N_7656);
nand U10909 (N_10909,N_8002,N_6659);
nor U10910 (N_10910,N_6643,N_7693);
nor U10911 (N_10911,N_6335,N_8384);
and U10912 (N_10912,N_8400,N_7678);
nor U10913 (N_10913,N_6052,N_8215);
and U10914 (N_10914,N_8452,N_8480);
and U10915 (N_10915,N_7656,N_7807);
and U10916 (N_10916,N_6200,N_6202);
and U10917 (N_10917,N_7084,N_7301);
and U10918 (N_10918,N_6957,N_6792);
and U10919 (N_10919,N_6429,N_6701);
and U10920 (N_10920,N_8519,N_8114);
and U10921 (N_10921,N_7721,N_8353);
nor U10922 (N_10922,N_7930,N_7895);
xnor U10923 (N_10923,N_7797,N_6091);
or U10924 (N_10924,N_8956,N_7371);
or U10925 (N_10925,N_8691,N_7684);
or U10926 (N_10926,N_6134,N_7451);
nor U10927 (N_10927,N_7354,N_7112);
nand U10928 (N_10928,N_6353,N_6296);
nor U10929 (N_10929,N_7793,N_7459);
and U10930 (N_10930,N_6861,N_8737);
nand U10931 (N_10931,N_7519,N_7251);
or U10932 (N_10932,N_7819,N_7011);
or U10933 (N_10933,N_7465,N_6999);
or U10934 (N_10934,N_6220,N_8406);
and U10935 (N_10935,N_8246,N_8231);
or U10936 (N_10936,N_6512,N_6708);
nand U10937 (N_10937,N_7393,N_8108);
nand U10938 (N_10938,N_6911,N_6260);
or U10939 (N_10939,N_7996,N_8391);
nor U10940 (N_10940,N_6836,N_8893);
or U10941 (N_10941,N_8797,N_7176);
nor U10942 (N_10942,N_7767,N_7534);
and U10943 (N_10943,N_8948,N_8768);
nand U10944 (N_10944,N_6871,N_7258);
nand U10945 (N_10945,N_6201,N_8515);
or U10946 (N_10946,N_6192,N_8257);
and U10947 (N_10947,N_6378,N_7220);
nand U10948 (N_10948,N_6846,N_7804);
nor U10949 (N_10949,N_6079,N_7695);
or U10950 (N_10950,N_7789,N_7156);
and U10951 (N_10951,N_7572,N_7133);
or U10952 (N_10952,N_7313,N_6954);
or U10953 (N_10953,N_8307,N_6323);
nor U10954 (N_10954,N_6283,N_7586);
and U10955 (N_10955,N_6875,N_6490);
nand U10956 (N_10956,N_7806,N_8993);
or U10957 (N_10957,N_7093,N_7239);
nand U10958 (N_10958,N_6427,N_8556);
and U10959 (N_10959,N_7091,N_8522);
nor U10960 (N_10960,N_6164,N_7343);
and U10961 (N_10961,N_6260,N_7414);
and U10962 (N_10962,N_8585,N_8074);
nand U10963 (N_10963,N_6697,N_7242);
nor U10964 (N_10964,N_7679,N_7136);
and U10965 (N_10965,N_6793,N_6888);
or U10966 (N_10966,N_8747,N_7865);
xnor U10967 (N_10967,N_8739,N_7725);
and U10968 (N_10968,N_6862,N_8661);
or U10969 (N_10969,N_6318,N_6029);
nor U10970 (N_10970,N_7951,N_8749);
nor U10971 (N_10971,N_8729,N_8992);
nor U10972 (N_10972,N_8595,N_8288);
or U10973 (N_10973,N_8723,N_6464);
or U10974 (N_10974,N_6041,N_6908);
nor U10975 (N_10975,N_6307,N_6246);
and U10976 (N_10976,N_7929,N_7611);
nor U10977 (N_10977,N_6899,N_7860);
nor U10978 (N_10978,N_8250,N_8563);
nor U10979 (N_10979,N_7232,N_8502);
xor U10980 (N_10980,N_6361,N_8985);
nor U10981 (N_10981,N_8081,N_6189);
nor U10982 (N_10982,N_8496,N_7432);
nand U10983 (N_10983,N_6716,N_6633);
nor U10984 (N_10984,N_7561,N_8679);
nand U10985 (N_10985,N_6866,N_7140);
nor U10986 (N_10986,N_6326,N_8264);
nor U10987 (N_10987,N_8938,N_6285);
nor U10988 (N_10988,N_7539,N_8530);
nand U10989 (N_10989,N_8931,N_8684);
nand U10990 (N_10990,N_7080,N_6308);
or U10991 (N_10991,N_7010,N_6879);
nor U10992 (N_10992,N_6436,N_7943);
and U10993 (N_10993,N_6396,N_6854);
nand U10994 (N_10994,N_6261,N_8340);
nor U10995 (N_10995,N_7354,N_6610);
nor U10996 (N_10996,N_7206,N_6538);
xnor U10997 (N_10997,N_6399,N_7815);
or U10998 (N_10998,N_7821,N_8895);
or U10999 (N_10999,N_8862,N_7595);
and U11000 (N_11000,N_7787,N_6682);
or U11001 (N_11001,N_7530,N_6398);
or U11002 (N_11002,N_8215,N_8121);
nor U11003 (N_11003,N_8715,N_7606);
nor U11004 (N_11004,N_8722,N_8746);
nor U11005 (N_11005,N_8691,N_7247);
nor U11006 (N_11006,N_6382,N_8749);
nor U11007 (N_11007,N_8142,N_8288);
nor U11008 (N_11008,N_6205,N_8656);
or U11009 (N_11009,N_7810,N_8272);
or U11010 (N_11010,N_8410,N_8884);
nand U11011 (N_11011,N_6273,N_7207);
nor U11012 (N_11012,N_7510,N_6965);
nor U11013 (N_11013,N_7250,N_7006);
and U11014 (N_11014,N_8411,N_6844);
and U11015 (N_11015,N_8841,N_8599);
and U11016 (N_11016,N_7509,N_6716);
nand U11017 (N_11017,N_6459,N_8162);
and U11018 (N_11018,N_6264,N_8939);
nand U11019 (N_11019,N_8754,N_7029);
or U11020 (N_11020,N_7009,N_6513);
or U11021 (N_11021,N_7567,N_6359);
and U11022 (N_11022,N_8705,N_7455);
and U11023 (N_11023,N_7749,N_7796);
or U11024 (N_11024,N_7761,N_8296);
or U11025 (N_11025,N_6552,N_8626);
and U11026 (N_11026,N_6898,N_6272);
nor U11027 (N_11027,N_7579,N_8217);
nand U11028 (N_11028,N_6784,N_8258);
nand U11029 (N_11029,N_8336,N_8942);
nand U11030 (N_11030,N_6945,N_7328);
and U11031 (N_11031,N_7512,N_6814);
nand U11032 (N_11032,N_8229,N_7882);
and U11033 (N_11033,N_7889,N_8980);
and U11034 (N_11034,N_8249,N_8266);
and U11035 (N_11035,N_6154,N_8441);
and U11036 (N_11036,N_7932,N_6445);
or U11037 (N_11037,N_7256,N_7307);
or U11038 (N_11038,N_7625,N_7936);
and U11039 (N_11039,N_8375,N_8437);
or U11040 (N_11040,N_8707,N_7828);
and U11041 (N_11041,N_6210,N_7911);
and U11042 (N_11042,N_6432,N_7812);
or U11043 (N_11043,N_8483,N_7634);
nor U11044 (N_11044,N_7472,N_8170);
or U11045 (N_11045,N_6748,N_6866);
and U11046 (N_11046,N_6092,N_7211);
nand U11047 (N_11047,N_7298,N_7178);
and U11048 (N_11048,N_7730,N_6396);
xnor U11049 (N_11049,N_7342,N_8227);
nor U11050 (N_11050,N_7101,N_7640);
and U11051 (N_11051,N_7016,N_8898);
nand U11052 (N_11052,N_8316,N_8126);
and U11053 (N_11053,N_8664,N_6896);
or U11054 (N_11054,N_8331,N_7884);
and U11055 (N_11055,N_8536,N_6669);
and U11056 (N_11056,N_6873,N_6697);
and U11057 (N_11057,N_7351,N_7655);
nand U11058 (N_11058,N_8479,N_7772);
or U11059 (N_11059,N_8289,N_6316);
nand U11060 (N_11060,N_8979,N_8768);
nand U11061 (N_11061,N_7532,N_6067);
xor U11062 (N_11062,N_8882,N_7788);
xor U11063 (N_11063,N_7159,N_8742);
or U11064 (N_11064,N_6169,N_8780);
nand U11065 (N_11065,N_7977,N_7513);
nand U11066 (N_11066,N_7283,N_8697);
nor U11067 (N_11067,N_6608,N_8954);
and U11068 (N_11068,N_7605,N_6200);
and U11069 (N_11069,N_7277,N_7605);
or U11070 (N_11070,N_7048,N_6635);
nor U11071 (N_11071,N_7598,N_7362);
nor U11072 (N_11072,N_7011,N_8769);
nor U11073 (N_11073,N_7761,N_8004);
nand U11074 (N_11074,N_8933,N_8542);
or U11075 (N_11075,N_8363,N_7628);
and U11076 (N_11076,N_6013,N_6903);
nor U11077 (N_11077,N_7830,N_7639);
nand U11078 (N_11078,N_7250,N_6907);
or U11079 (N_11079,N_8630,N_6080);
nand U11080 (N_11080,N_6964,N_8100);
or U11081 (N_11081,N_6220,N_7469);
nor U11082 (N_11082,N_7302,N_8941);
and U11083 (N_11083,N_7683,N_6061);
nor U11084 (N_11084,N_6063,N_6341);
and U11085 (N_11085,N_7259,N_7821);
and U11086 (N_11086,N_6517,N_7440);
or U11087 (N_11087,N_7098,N_7218);
and U11088 (N_11088,N_6383,N_8151);
or U11089 (N_11089,N_8543,N_7801);
and U11090 (N_11090,N_8986,N_8993);
and U11091 (N_11091,N_8131,N_8326);
and U11092 (N_11092,N_6927,N_8005);
nand U11093 (N_11093,N_7868,N_8655);
and U11094 (N_11094,N_8235,N_7492);
and U11095 (N_11095,N_8416,N_7728);
nor U11096 (N_11096,N_8728,N_8148);
or U11097 (N_11097,N_8876,N_8586);
nand U11098 (N_11098,N_6394,N_6814);
nand U11099 (N_11099,N_8981,N_6244);
and U11100 (N_11100,N_8305,N_6279);
and U11101 (N_11101,N_8050,N_7389);
nor U11102 (N_11102,N_8962,N_6019);
or U11103 (N_11103,N_7860,N_8892);
nor U11104 (N_11104,N_7744,N_6792);
and U11105 (N_11105,N_8178,N_7336);
or U11106 (N_11106,N_8145,N_7650);
and U11107 (N_11107,N_7837,N_6235);
and U11108 (N_11108,N_8524,N_7822);
or U11109 (N_11109,N_6580,N_6512);
and U11110 (N_11110,N_6211,N_8604);
or U11111 (N_11111,N_7868,N_8949);
nand U11112 (N_11112,N_7984,N_7160);
nand U11113 (N_11113,N_8332,N_7002);
nand U11114 (N_11114,N_6681,N_7377);
nor U11115 (N_11115,N_7501,N_7677);
nor U11116 (N_11116,N_6532,N_7409);
nand U11117 (N_11117,N_6422,N_6622);
nor U11118 (N_11118,N_7463,N_6166);
or U11119 (N_11119,N_6161,N_6644);
or U11120 (N_11120,N_7625,N_6440);
nor U11121 (N_11121,N_8346,N_8840);
nor U11122 (N_11122,N_6112,N_8762);
nand U11123 (N_11123,N_8969,N_6297);
or U11124 (N_11124,N_7649,N_7111);
and U11125 (N_11125,N_6691,N_7705);
nor U11126 (N_11126,N_6313,N_8959);
or U11127 (N_11127,N_6132,N_6145);
nand U11128 (N_11128,N_6147,N_8834);
or U11129 (N_11129,N_7274,N_8199);
or U11130 (N_11130,N_7498,N_7536);
nor U11131 (N_11131,N_8301,N_6098);
or U11132 (N_11132,N_6440,N_7394);
or U11133 (N_11133,N_8641,N_6355);
nand U11134 (N_11134,N_6807,N_8395);
nand U11135 (N_11135,N_8734,N_7886);
nor U11136 (N_11136,N_7613,N_7690);
or U11137 (N_11137,N_6365,N_7110);
nor U11138 (N_11138,N_8286,N_7117);
nand U11139 (N_11139,N_7915,N_8040);
nor U11140 (N_11140,N_7278,N_6548);
nor U11141 (N_11141,N_8554,N_7702);
or U11142 (N_11142,N_6852,N_6970);
xor U11143 (N_11143,N_7606,N_7983);
and U11144 (N_11144,N_8088,N_6704);
nand U11145 (N_11145,N_7261,N_6128);
and U11146 (N_11146,N_6903,N_8115);
and U11147 (N_11147,N_7008,N_6815);
nor U11148 (N_11148,N_6336,N_6322);
or U11149 (N_11149,N_8343,N_6370);
nor U11150 (N_11150,N_7243,N_6580);
nor U11151 (N_11151,N_7023,N_8788);
and U11152 (N_11152,N_6639,N_7001);
nand U11153 (N_11153,N_8006,N_7936);
or U11154 (N_11154,N_6608,N_6052);
nand U11155 (N_11155,N_8946,N_7344);
and U11156 (N_11156,N_7101,N_6874);
and U11157 (N_11157,N_8076,N_7870);
nand U11158 (N_11158,N_7502,N_7255);
or U11159 (N_11159,N_8866,N_7349);
nand U11160 (N_11160,N_6359,N_6965);
nand U11161 (N_11161,N_7345,N_6576);
or U11162 (N_11162,N_6764,N_8611);
and U11163 (N_11163,N_7002,N_7204);
or U11164 (N_11164,N_7596,N_8674);
and U11165 (N_11165,N_6197,N_8720);
nor U11166 (N_11166,N_8459,N_8533);
nand U11167 (N_11167,N_6170,N_8509);
nor U11168 (N_11168,N_8076,N_6796);
or U11169 (N_11169,N_6404,N_8982);
nand U11170 (N_11170,N_6917,N_6219);
or U11171 (N_11171,N_7758,N_6279);
nor U11172 (N_11172,N_7450,N_7844);
nand U11173 (N_11173,N_6060,N_6340);
nand U11174 (N_11174,N_7400,N_6530);
nor U11175 (N_11175,N_7626,N_7250);
and U11176 (N_11176,N_8637,N_7436);
or U11177 (N_11177,N_8942,N_8514);
nor U11178 (N_11178,N_7412,N_8504);
or U11179 (N_11179,N_7145,N_8582);
nand U11180 (N_11180,N_8639,N_7690);
or U11181 (N_11181,N_7131,N_7895);
or U11182 (N_11182,N_6770,N_7949);
or U11183 (N_11183,N_6229,N_7488);
nand U11184 (N_11184,N_8240,N_8644);
or U11185 (N_11185,N_8036,N_8225);
nor U11186 (N_11186,N_8941,N_6232);
nor U11187 (N_11187,N_6703,N_7706);
and U11188 (N_11188,N_6014,N_8383);
xor U11189 (N_11189,N_6414,N_7010);
and U11190 (N_11190,N_7470,N_8766);
nor U11191 (N_11191,N_8217,N_8438);
or U11192 (N_11192,N_8014,N_7236);
and U11193 (N_11193,N_7656,N_6354);
nand U11194 (N_11194,N_8537,N_8797);
or U11195 (N_11195,N_6205,N_7623);
and U11196 (N_11196,N_6420,N_8350);
nand U11197 (N_11197,N_7793,N_6408);
nor U11198 (N_11198,N_6600,N_6532);
or U11199 (N_11199,N_6777,N_8398);
or U11200 (N_11200,N_7045,N_6025);
or U11201 (N_11201,N_6969,N_6901);
or U11202 (N_11202,N_7990,N_6332);
or U11203 (N_11203,N_7000,N_8452);
or U11204 (N_11204,N_6728,N_7883);
nand U11205 (N_11205,N_8641,N_7516);
nand U11206 (N_11206,N_7465,N_8445);
or U11207 (N_11207,N_8371,N_8186);
nor U11208 (N_11208,N_8918,N_6889);
and U11209 (N_11209,N_8967,N_8327);
nand U11210 (N_11210,N_7965,N_8284);
nand U11211 (N_11211,N_6187,N_6177);
nor U11212 (N_11212,N_7044,N_8396);
nor U11213 (N_11213,N_6522,N_8827);
nand U11214 (N_11214,N_7920,N_6100);
nor U11215 (N_11215,N_6794,N_7749);
nor U11216 (N_11216,N_7083,N_6989);
nand U11217 (N_11217,N_8360,N_6236);
xnor U11218 (N_11218,N_7146,N_8658);
nand U11219 (N_11219,N_6384,N_8425);
nor U11220 (N_11220,N_8415,N_6049);
and U11221 (N_11221,N_7324,N_6810);
nor U11222 (N_11222,N_6994,N_7731);
and U11223 (N_11223,N_7853,N_8342);
or U11224 (N_11224,N_7936,N_6726);
or U11225 (N_11225,N_7882,N_7030);
nand U11226 (N_11226,N_8143,N_7930);
nand U11227 (N_11227,N_7275,N_7246);
nor U11228 (N_11228,N_7021,N_8091);
nor U11229 (N_11229,N_8197,N_8256);
nand U11230 (N_11230,N_6278,N_8803);
nor U11231 (N_11231,N_8680,N_8409);
nand U11232 (N_11232,N_8464,N_6920);
and U11233 (N_11233,N_6098,N_8851);
and U11234 (N_11234,N_7718,N_6824);
nand U11235 (N_11235,N_8545,N_8549);
nor U11236 (N_11236,N_7730,N_7818);
or U11237 (N_11237,N_7767,N_7580);
or U11238 (N_11238,N_6997,N_7855);
nor U11239 (N_11239,N_6159,N_8473);
and U11240 (N_11240,N_7893,N_8098);
and U11241 (N_11241,N_7166,N_6228);
or U11242 (N_11242,N_6873,N_7376);
or U11243 (N_11243,N_8429,N_6319);
and U11244 (N_11244,N_8072,N_6816);
and U11245 (N_11245,N_6398,N_6487);
or U11246 (N_11246,N_7321,N_6871);
nor U11247 (N_11247,N_8944,N_7623);
xor U11248 (N_11248,N_8396,N_6312);
nand U11249 (N_11249,N_6371,N_8796);
and U11250 (N_11250,N_7592,N_8321);
nand U11251 (N_11251,N_7155,N_6782);
nand U11252 (N_11252,N_8033,N_6351);
or U11253 (N_11253,N_6555,N_8040);
nand U11254 (N_11254,N_7872,N_6347);
nand U11255 (N_11255,N_6355,N_7988);
or U11256 (N_11256,N_7080,N_6240);
and U11257 (N_11257,N_8161,N_6636);
nand U11258 (N_11258,N_8245,N_8060);
and U11259 (N_11259,N_7792,N_6242);
and U11260 (N_11260,N_6492,N_8269);
and U11261 (N_11261,N_8240,N_6660);
nor U11262 (N_11262,N_7907,N_6551);
nor U11263 (N_11263,N_8347,N_8911);
nand U11264 (N_11264,N_6094,N_8860);
and U11265 (N_11265,N_8752,N_8939);
and U11266 (N_11266,N_6802,N_8697);
nor U11267 (N_11267,N_6035,N_7023);
and U11268 (N_11268,N_6071,N_7009);
or U11269 (N_11269,N_7198,N_7015);
nand U11270 (N_11270,N_6509,N_8015);
nor U11271 (N_11271,N_8657,N_8376);
nor U11272 (N_11272,N_8549,N_6433);
nor U11273 (N_11273,N_6521,N_6737);
and U11274 (N_11274,N_8689,N_6676);
nor U11275 (N_11275,N_7801,N_7464);
and U11276 (N_11276,N_8751,N_8740);
nor U11277 (N_11277,N_7816,N_8368);
nor U11278 (N_11278,N_7905,N_8118);
nor U11279 (N_11279,N_7587,N_7781);
or U11280 (N_11280,N_7233,N_7373);
xnor U11281 (N_11281,N_7262,N_6432);
xor U11282 (N_11282,N_7343,N_6966);
or U11283 (N_11283,N_7429,N_7590);
nor U11284 (N_11284,N_7185,N_8858);
and U11285 (N_11285,N_6072,N_7200);
nand U11286 (N_11286,N_8830,N_7974);
nor U11287 (N_11287,N_7902,N_7709);
and U11288 (N_11288,N_7665,N_7875);
nand U11289 (N_11289,N_8608,N_8369);
nand U11290 (N_11290,N_8964,N_8015);
and U11291 (N_11291,N_8760,N_7617);
and U11292 (N_11292,N_7080,N_6891);
nand U11293 (N_11293,N_8323,N_7247);
nor U11294 (N_11294,N_6854,N_8173);
nor U11295 (N_11295,N_7668,N_7439);
nor U11296 (N_11296,N_8682,N_8284);
and U11297 (N_11297,N_7417,N_8399);
nor U11298 (N_11298,N_6557,N_8394);
nand U11299 (N_11299,N_7209,N_8971);
nor U11300 (N_11300,N_7961,N_6913);
and U11301 (N_11301,N_6354,N_8898);
xor U11302 (N_11302,N_8186,N_7546);
or U11303 (N_11303,N_7314,N_6225);
and U11304 (N_11304,N_8157,N_6281);
or U11305 (N_11305,N_7004,N_8152);
nand U11306 (N_11306,N_8056,N_8500);
and U11307 (N_11307,N_6811,N_7583);
and U11308 (N_11308,N_6135,N_6536);
nor U11309 (N_11309,N_7114,N_6778);
and U11310 (N_11310,N_6857,N_6634);
nand U11311 (N_11311,N_6748,N_7406);
xor U11312 (N_11312,N_7855,N_6688);
nor U11313 (N_11313,N_7360,N_7211);
nor U11314 (N_11314,N_6427,N_7253);
or U11315 (N_11315,N_6386,N_8613);
or U11316 (N_11316,N_6380,N_7557);
and U11317 (N_11317,N_8589,N_7729);
or U11318 (N_11318,N_8602,N_6860);
and U11319 (N_11319,N_6404,N_7564);
nand U11320 (N_11320,N_8498,N_7801);
nor U11321 (N_11321,N_6178,N_7431);
nor U11322 (N_11322,N_7240,N_6040);
or U11323 (N_11323,N_7471,N_8145);
xnor U11324 (N_11324,N_7898,N_6288);
or U11325 (N_11325,N_6916,N_8915);
or U11326 (N_11326,N_7069,N_6701);
nand U11327 (N_11327,N_8506,N_6582);
and U11328 (N_11328,N_6558,N_7001);
and U11329 (N_11329,N_8711,N_7561);
and U11330 (N_11330,N_7950,N_7788);
xor U11331 (N_11331,N_7426,N_8066);
nor U11332 (N_11332,N_7515,N_8414);
and U11333 (N_11333,N_7780,N_8268);
nor U11334 (N_11334,N_8966,N_7379);
or U11335 (N_11335,N_6977,N_7977);
or U11336 (N_11336,N_8561,N_8187);
or U11337 (N_11337,N_7493,N_8311);
or U11338 (N_11338,N_7868,N_8222);
nand U11339 (N_11339,N_8995,N_6706);
or U11340 (N_11340,N_6240,N_7496);
nor U11341 (N_11341,N_6069,N_8086);
or U11342 (N_11342,N_8707,N_7150);
and U11343 (N_11343,N_8419,N_6580);
and U11344 (N_11344,N_6796,N_7260);
and U11345 (N_11345,N_7134,N_8488);
and U11346 (N_11346,N_7684,N_8478);
nand U11347 (N_11347,N_7283,N_7929);
nor U11348 (N_11348,N_6960,N_8123);
or U11349 (N_11349,N_8711,N_8147);
nand U11350 (N_11350,N_6506,N_7781);
nand U11351 (N_11351,N_8075,N_8379);
or U11352 (N_11352,N_8414,N_6400);
nor U11353 (N_11353,N_6266,N_6377);
nand U11354 (N_11354,N_6582,N_7740);
or U11355 (N_11355,N_6318,N_7977);
nor U11356 (N_11356,N_8834,N_7171);
nand U11357 (N_11357,N_7840,N_7446);
nor U11358 (N_11358,N_6507,N_7463);
and U11359 (N_11359,N_7873,N_7658);
nor U11360 (N_11360,N_6566,N_8156);
or U11361 (N_11361,N_7145,N_6519);
or U11362 (N_11362,N_7439,N_8810);
or U11363 (N_11363,N_8890,N_8375);
nand U11364 (N_11364,N_6348,N_6343);
or U11365 (N_11365,N_8097,N_6205);
nor U11366 (N_11366,N_8464,N_7507);
and U11367 (N_11367,N_7562,N_8529);
and U11368 (N_11368,N_7554,N_8744);
nand U11369 (N_11369,N_7588,N_6616);
and U11370 (N_11370,N_6085,N_7396);
nor U11371 (N_11371,N_6828,N_7411);
and U11372 (N_11372,N_7762,N_6802);
and U11373 (N_11373,N_7717,N_7688);
and U11374 (N_11374,N_8006,N_6729);
or U11375 (N_11375,N_7710,N_8740);
nor U11376 (N_11376,N_6633,N_8350);
and U11377 (N_11377,N_7801,N_7633);
or U11378 (N_11378,N_8748,N_6941);
nor U11379 (N_11379,N_7741,N_6005);
and U11380 (N_11380,N_6255,N_8255);
or U11381 (N_11381,N_6717,N_6600);
or U11382 (N_11382,N_8338,N_6373);
or U11383 (N_11383,N_6966,N_6516);
and U11384 (N_11384,N_6648,N_6723);
or U11385 (N_11385,N_7983,N_6438);
nor U11386 (N_11386,N_7100,N_8048);
nand U11387 (N_11387,N_6223,N_7931);
nor U11388 (N_11388,N_8933,N_7716);
nand U11389 (N_11389,N_6623,N_8334);
and U11390 (N_11390,N_6087,N_6094);
nor U11391 (N_11391,N_7087,N_7757);
and U11392 (N_11392,N_7493,N_8513);
xnor U11393 (N_11393,N_8792,N_6162);
xnor U11394 (N_11394,N_6300,N_8898);
and U11395 (N_11395,N_7979,N_8474);
nor U11396 (N_11396,N_8776,N_6877);
nand U11397 (N_11397,N_6898,N_7113);
or U11398 (N_11398,N_6150,N_7327);
nor U11399 (N_11399,N_7926,N_8504);
nor U11400 (N_11400,N_6803,N_8908);
xor U11401 (N_11401,N_6011,N_6052);
and U11402 (N_11402,N_6626,N_7168);
nor U11403 (N_11403,N_7107,N_7066);
nor U11404 (N_11404,N_7735,N_6126);
nor U11405 (N_11405,N_6441,N_6622);
and U11406 (N_11406,N_8829,N_7211);
nor U11407 (N_11407,N_7496,N_6129);
and U11408 (N_11408,N_8767,N_6306);
and U11409 (N_11409,N_7716,N_8577);
and U11410 (N_11410,N_7014,N_7845);
nor U11411 (N_11411,N_8833,N_7913);
and U11412 (N_11412,N_6225,N_7185);
nand U11413 (N_11413,N_8829,N_7751);
nor U11414 (N_11414,N_7693,N_7654);
or U11415 (N_11415,N_8286,N_6051);
or U11416 (N_11416,N_7469,N_7988);
or U11417 (N_11417,N_8671,N_7719);
and U11418 (N_11418,N_7806,N_7347);
nand U11419 (N_11419,N_7844,N_8231);
nor U11420 (N_11420,N_7085,N_6036);
nor U11421 (N_11421,N_8054,N_7004);
nor U11422 (N_11422,N_6366,N_7286);
or U11423 (N_11423,N_7648,N_8279);
and U11424 (N_11424,N_7571,N_7495);
and U11425 (N_11425,N_8620,N_7299);
and U11426 (N_11426,N_6332,N_7690);
and U11427 (N_11427,N_7376,N_7794);
nor U11428 (N_11428,N_6160,N_6458);
and U11429 (N_11429,N_7779,N_8342);
nand U11430 (N_11430,N_6637,N_7257);
nand U11431 (N_11431,N_7045,N_6165);
or U11432 (N_11432,N_6862,N_8904);
and U11433 (N_11433,N_7349,N_7929);
xor U11434 (N_11434,N_8084,N_8055);
nand U11435 (N_11435,N_8107,N_6100);
or U11436 (N_11436,N_8490,N_7375);
nor U11437 (N_11437,N_6980,N_8634);
nor U11438 (N_11438,N_7230,N_6743);
and U11439 (N_11439,N_7834,N_6565);
or U11440 (N_11440,N_7078,N_6868);
nand U11441 (N_11441,N_6441,N_6914);
nand U11442 (N_11442,N_7492,N_8485);
and U11443 (N_11443,N_8365,N_8675);
nor U11444 (N_11444,N_8519,N_8962);
nor U11445 (N_11445,N_6589,N_8415);
or U11446 (N_11446,N_6072,N_6086);
or U11447 (N_11447,N_6487,N_6374);
or U11448 (N_11448,N_6259,N_8758);
or U11449 (N_11449,N_8012,N_7461);
nor U11450 (N_11450,N_7965,N_7841);
or U11451 (N_11451,N_6873,N_6834);
xor U11452 (N_11452,N_8397,N_6286);
or U11453 (N_11453,N_8145,N_6647);
nand U11454 (N_11454,N_6742,N_6020);
or U11455 (N_11455,N_7470,N_6061);
and U11456 (N_11456,N_8689,N_8926);
nor U11457 (N_11457,N_8710,N_6309);
nor U11458 (N_11458,N_6929,N_8200);
and U11459 (N_11459,N_8183,N_6223);
nand U11460 (N_11460,N_8733,N_8568);
nand U11461 (N_11461,N_8713,N_7400);
xnor U11462 (N_11462,N_6899,N_8779);
and U11463 (N_11463,N_8423,N_6460);
or U11464 (N_11464,N_8246,N_6987);
or U11465 (N_11465,N_7012,N_8740);
and U11466 (N_11466,N_7995,N_7611);
nor U11467 (N_11467,N_6926,N_7635);
nand U11468 (N_11468,N_7964,N_6309);
nor U11469 (N_11469,N_6685,N_8165);
nor U11470 (N_11470,N_6285,N_6903);
and U11471 (N_11471,N_7675,N_6142);
or U11472 (N_11472,N_6366,N_7464);
nor U11473 (N_11473,N_8101,N_8937);
and U11474 (N_11474,N_6206,N_7492);
and U11475 (N_11475,N_6958,N_6857);
and U11476 (N_11476,N_6793,N_6134);
or U11477 (N_11477,N_7081,N_6601);
or U11478 (N_11478,N_7892,N_7554);
nor U11479 (N_11479,N_8216,N_6046);
and U11480 (N_11480,N_8154,N_7835);
and U11481 (N_11481,N_6893,N_6496);
or U11482 (N_11482,N_6401,N_8612);
or U11483 (N_11483,N_7765,N_6617);
nor U11484 (N_11484,N_7837,N_8718);
nor U11485 (N_11485,N_7305,N_8266);
nand U11486 (N_11486,N_8104,N_8051);
nand U11487 (N_11487,N_6297,N_6556);
nor U11488 (N_11488,N_8864,N_6088);
or U11489 (N_11489,N_7598,N_6160);
or U11490 (N_11490,N_6088,N_8133);
or U11491 (N_11491,N_6195,N_6501);
and U11492 (N_11492,N_6430,N_6860);
or U11493 (N_11493,N_6014,N_8155);
nor U11494 (N_11494,N_8461,N_7407);
nand U11495 (N_11495,N_8924,N_7536);
or U11496 (N_11496,N_7813,N_6386);
or U11497 (N_11497,N_6223,N_7793);
nand U11498 (N_11498,N_7063,N_6684);
and U11499 (N_11499,N_6729,N_6775);
and U11500 (N_11500,N_8308,N_6333);
nand U11501 (N_11501,N_6913,N_7883);
xnor U11502 (N_11502,N_7165,N_6325);
and U11503 (N_11503,N_8230,N_7622);
and U11504 (N_11504,N_8629,N_7804);
nand U11505 (N_11505,N_8901,N_7033);
nor U11506 (N_11506,N_8629,N_6227);
or U11507 (N_11507,N_6999,N_6438);
nor U11508 (N_11508,N_7173,N_6549);
or U11509 (N_11509,N_8273,N_7503);
and U11510 (N_11510,N_8241,N_7375);
xor U11511 (N_11511,N_7209,N_6924);
and U11512 (N_11512,N_8907,N_6480);
xor U11513 (N_11513,N_7640,N_8644);
nand U11514 (N_11514,N_7504,N_7611);
nor U11515 (N_11515,N_7177,N_8195);
or U11516 (N_11516,N_6994,N_8969);
nand U11517 (N_11517,N_6664,N_6326);
xnor U11518 (N_11518,N_6034,N_6395);
nand U11519 (N_11519,N_8164,N_7502);
or U11520 (N_11520,N_8618,N_6780);
or U11521 (N_11521,N_7732,N_8021);
nor U11522 (N_11522,N_8341,N_7782);
nand U11523 (N_11523,N_7852,N_7527);
and U11524 (N_11524,N_8971,N_6901);
or U11525 (N_11525,N_6943,N_6643);
xor U11526 (N_11526,N_8085,N_6785);
and U11527 (N_11527,N_6563,N_7317);
xnor U11528 (N_11528,N_8267,N_8423);
and U11529 (N_11529,N_8727,N_6818);
nand U11530 (N_11530,N_6003,N_6140);
nor U11531 (N_11531,N_8396,N_6754);
xnor U11532 (N_11532,N_8804,N_7284);
and U11533 (N_11533,N_8501,N_6061);
and U11534 (N_11534,N_6860,N_8736);
and U11535 (N_11535,N_8708,N_8774);
and U11536 (N_11536,N_6278,N_8811);
nand U11537 (N_11537,N_8812,N_6771);
or U11538 (N_11538,N_8264,N_7890);
and U11539 (N_11539,N_7449,N_8884);
or U11540 (N_11540,N_6646,N_7709);
and U11541 (N_11541,N_7734,N_6408);
and U11542 (N_11542,N_6488,N_8076);
and U11543 (N_11543,N_8416,N_7077);
and U11544 (N_11544,N_6078,N_6630);
and U11545 (N_11545,N_8949,N_7722);
nor U11546 (N_11546,N_8380,N_8570);
nand U11547 (N_11547,N_6732,N_7882);
and U11548 (N_11548,N_7178,N_8558);
or U11549 (N_11549,N_7997,N_7169);
nand U11550 (N_11550,N_6910,N_8998);
nand U11551 (N_11551,N_7637,N_6175);
nor U11552 (N_11552,N_8060,N_7407);
nand U11553 (N_11553,N_7616,N_6531);
nand U11554 (N_11554,N_7537,N_8970);
nor U11555 (N_11555,N_6871,N_8945);
or U11556 (N_11556,N_7767,N_8023);
or U11557 (N_11557,N_7661,N_8521);
nor U11558 (N_11558,N_8331,N_7262);
xnor U11559 (N_11559,N_7332,N_7700);
nor U11560 (N_11560,N_7973,N_6311);
or U11561 (N_11561,N_8359,N_7176);
nor U11562 (N_11562,N_8796,N_8136);
nand U11563 (N_11563,N_7469,N_8295);
xnor U11564 (N_11564,N_6159,N_6784);
and U11565 (N_11565,N_6589,N_6817);
nand U11566 (N_11566,N_8175,N_8882);
nand U11567 (N_11567,N_8331,N_8663);
or U11568 (N_11568,N_6295,N_7018);
nand U11569 (N_11569,N_7015,N_6659);
nand U11570 (N_11570,N_8483,N_7480);
nor U11571 (N_11571,N_8063,N_6641);
or U11572 (N_11572,N_7248,N_6324);
xnor U11573 (N_11573,N_6948,N_6367);
and U11574 (N_11574,N_7342,N_6717);
nor U11575 (N_11575,N_7335,N_6292);
nand U11576 (N_11576,N_6456,N_8644);
nand U11577 (N_11577,N_8135,N_8985);
and U11578 (N_11578,N_7444,N_6974);
nor U11579 (N_11579,N_8897,N_8064);
and U11580 (N_11580,N_7171,N_7785);
and U11581 (N_11581,N_7176,N_6598);
nand U11582 (N_11582,N_7427,N_7560);
xor U11583 (N_11583,N_7727,N_7715);
nor U11584 (N_11584,N_7804,N_7693);
nand U11585 (N_11585,N_8054,N_7717);
or U11586 (N_11586,N_6325,N_6103);
nor U11587 (N_11587,N_6650,N_8144);
nor U11588 (N_11588,N_6273,N_6857);
nor U11589 (N_11589,N_7338,N_6192);
or U11590 (N_11590,N_8425,N_8104);
nand U11591 (N_11591,N_8066,N_7457);
and U11592 (N_11592,N_6346,N_6452);
nand U11593 (N_11593,N_6887,N_8543);
nand U11594 (N_11594,N_6763,N_7362);
or U11595 (N_11595,N_7037,N_8193);
and U11596 (N_11596,N_7451,N_6791);
and U11597 (N_11597,N_6906,N_8314);
nand U11598 (N_11598,N_7482,N_7749);
nand U11599 (N_11599,N_8168,N_8316);
or U11600 (N_11600,N_7341,N_7400);
and U11601 (N_11601,N_7986,N_6406);
and U11602 (N_11602,N_8218,N_8340);
nor U11603 (N_11603,N_7127,N_6466);
or U11604 (N_11604,N_7199,N_7180);
or U11605 (N_11605,N_7566,N_8145);
nand U11606 (N_11606,N_6677,N_7414);
nand U11607 (N_11607,N_7388,N_7251);
nor U11608 (N_11608,N_7426,N_7756);
and U11609 (N_11609,N_6050,N_6746);
or U11610 (N_11610,N_7456,N_8383);
or U11611 (N_11611,N_6215,N_6543);
nor U11612 (N_11612,N_6585,N_8359);
nand U11613 (N_11613,N_8930,N_7807);
and U11614 (N_11614,N_6141,N_7417);
nand U11615 (N_11615,N_8811,N_8348);
nand U11616 (N_11616,N_8946,N_8455);
or U11617 (N_11617,N_7534,N_7132);
xnor U11618 (N_11618,N_6596,N_8491);
nand U11619 (N_11619,N_8336,N_7360);
nand U11620 (N_11620,N_6322,N_7381);
nor U11621 (N_11621,N_8677,N_6035);
or U11622 (N_11622,N_8703,N_6826);
nand U11623 (N_11623,N_8177,N_6038);
or U11624 (N_11624,N_8160,N_6351);
and U11625 (N_11625,N_7700,N_7432);
and U11626 (N_11626,N_6044,N_7343);
nand U11627 (N_11627,N_6980,N_7641);
or U11628 (N_11628,N_8190,N_6863);
and U11629 (N_11629,N_6962,N_8313);
nand U11630 (N_11630,N_7692,N_8482);
or U11631 (N_11631,N_6116,N_8489);
nand U11632 (N_11632,N_6862,N_6413);
or U11633 (N_11633,N_8074,N_6797);
or U11634 (N_11634,N_7305,N_7499);
nand U11635 (N_11635,N_8994,N_6268);
or U11636 (N_11636,N_6423,N_8571);
nand U11637 (N_11637,N_7873,N_8950);
or U11638 (N_11638,N_6755,N_8328);
or U11639 (N_11639,N_6023,N_8303);
xnor U11640 (N_11640,N_6229,N_8880);
and U11641 (N_11641,N_6550,N_8029);
nand U11642 (N_11642,N_8311,N_7248);
or U11643 (N_11643,N_7616,N_6266);
or U11644 (N_11644,N_7038,N_6077);
or U11645 (N_11645,N_6706,N_7000);
or U11646 (N_11646,N_6329,N_7404);
nor U11647 (N_11647,N_8002,N_7563);
and U11648 (N_11648,N_6801,N_6844);
or U11649 (N_11649,N_8878,N_6395);
nor U11650 (N_11650,N_8505,N_7706);
or U11651 (N_11651,N_7331,N_6290);
nand U11652 (N_11652,N_8634,N_6863);
and U11653 (N_11653,N_8596,N_8091);
nor U11654 (N_11654,N_6899,N_8031);
nand U11655 (N_11655,N_7473,N_8141);
and U11656 (N_11656,N_6370,N_7505);
nand U11657 (N_11657,N_8088,N_7202);
nand U11658 (N_11658,N_8551,N_7966);
nand U11659 (N_11659,N_8649,N_8299);
and U11660 (N_11660,N_8960,N_8447);
or U11661 (N_11661,N_6199,N_6853);
nor U11662 (N_11662,N_6820,N_8039);
or U11663 (N_11663,N_6294,N_8135);
nand U11664 (N_11664,N_7917,N_6872);
nor U11665 (N_11665,N_7984,N_8967);
nor U11666 (N_11666,N_6302,N_7225);
and U11667 (N_11667,N_8746,N_6876);
nor U11668 (N_11668,N_6889,N_6159);
and U11669 (N_11669,N_6449,N_6090);
nor U11670 (N_11670,N_8794,N_8176);
and U11671 (N_11671,N_8600,N_8186);
nand U11672 (N_11672,N_6271,N_7904);
xnor U11673 (N_11673,N_7213,N_6717);
nand U11674 (N_11674,N_8637,N_7696);
nand U11675 (N_11675,N_8605,N_6669);
nor U11676 (N_11676,N_7077,N_6700);
and U11677 (N_11677,N_6205,N_7811);
and U11678 (N_11678,N_8710,N_8004);
nor U11679 (N_11679,N_7137,N_7967);
nand U11680 (N_11680,N_8216,N_8386);
nand U11681 (N_11681,N_7938,N_8206);
or U11682 (N_11682,N_7788,N_6416);
nor U11683 (N_11683,N_7457,N_7389);
nand U11684 (N_11684,N_7443,N_7619);
nor U11685 (N_11685,N_6671,N_6400);
nor U11686 (N_11686,N_7111,N_7345);
nand U11687 (N_11687,N_8074,N_8055);
nor U11688 (N_11688,N_8734,N_7740);
nor U11689 (N_11689,N_8260,N_7809);
or U11690 (N_11690,N_7573,N_8516);
nor U11691 (N_11691,N_7809,N_7576);
nor U11692 (N_11692,N_6753,N_8991);
and U11693 (N_11693,N_8602,N_7791);
nor U11694 (N_11694,N_8884,N_8870);
or U11695 (N_11695,N_7013,N_7057);
nor U11696 (N_11696,N_8807,N_8839);
nor U11697 (N_11697,N_7729,N_8947);
or U11698 (N_11698,N_6514,N_6160);
or U11699 (N_11699,N_8637,N_7798);
nor U11700 (N_11700,N_6363,N_7873);
and U11701 (N_11701,N_6515,N_7357);
nor U11702 (N_11702,N_8015,N_8552);
nand U11703 (N_11703,N_7386,N_7702);
or U11704 (N_11704,N_8221,N_7697);
nand U11705 (N_11705,N_6697,N_6389);
nor U11706 (N_11706,N_7395,N_7907);
and U11707 (N_11707,N_8142,N_6890);
or U11708 (N_11708,N_7462,N_7488);
or U11709 (N_11709,N_7593,N_7584);
or U11710 (N_11710,N_8549,N_7948);
nor U11711 (N_11711,N_7355,N_6002);
or U11712 (N_11712,N_8970,N_8504);
nor U11713 (N_11713,N_7932,N_8549);
nand U11714 (N_11714,N_6229,N_8647);
nand U11715 (N_11715,N_6216,N_8136);
nor U11716 (N_11716,N_8894,N_7734);
nor U11717 (N_11717,N_6114,N_6335);
and U11718 (N_11718,N_8276,N_8942);
xnor U11719 (N_11719,N_7739,N_6573);
or U11720 (N_11720,N_8826,N_7450);
nand U11721 (N_11721,N_6299,N_7725);
xor U11722 (N_11722,N_8270,N_8851);
or U11723 (N_11723,N_6691,N_6956);
nor U11724 (N_11724,N_6396,N_7423);
nor U11725 (N_11725,N_8850,N_7388);
nor U11726 (N_11726,N_6185,N_7313);
nor U11727 (N_11727,N_8939,N_7558);
nand U11728 (N_11728,N_6684,N_7730);
or U11729 (N_11729,N_7965,N_7633);
nor U11730 (N_11730,N_8635,N_6782);
and U11731 (N_11731,N_8887,N_7564);
or U11732 (N_11732,N_8658,N_6243);
nand U11733 (N_11733,N_6557,N_7786);
nand U11734 (N_11734,N_6055,N_6250);
or U11735 (N_11735,N_8381,N_7618);
and U11736 (N_11736,N_6555,N_6276);
nand U11737 (N_11737,N_8142,N_8675);
nand U11738 (N_11738,N_6084,N_8718);
nor U11739 (N_11739,N_6676,N_8462);
nor U11740 (N_11740,N_7824,N_6086);
xor U11741 (N_11741,N_6771,N_6410);
nor U11742 (N_11742,N_6165,N_6699);
nor U11743 (N_11743,N_7635,N_8131);
nand U11744 (N_11744,N_6028,N_7584);
or U11745 (N_11745,N_8073,N_7550);
or U11746 (N_11746,N_7238,N_8181);
or U11747 (N_11747,N_6802,N_6619);
nand U11748 (N_11748,N_7915,N_6809);
and U11749 (N_11749,N_6013,N_8735);
nand U11750 (N_11750,N_7141,N_7508);
nor U11751 (N_11751,N_8142,N_8298);
and U11752 (N_11752,N_6602,N_6346);
and U11753 (N_11753,N_8578,N_6100);
nor U11754 (N_11754,N_7540,N_6348);
nor U11755 (N_11755,N_7993,N_6462);
and U11756 (N_11756,N_7675,N_7029);
nand U11757 (N_11757,N_8052,N_6821);
nor U11758 (N_11758,N_7033,N_7882);
or U11759 (N_11759,N_7637,N_7930);
nor U11760 (N_11760,N_6185,N_8344);
and U11761 (N_11761,N_6977,N_6152);
nand U11762 (N_11762,N_6766,N_8732);
nor U11763 (N_11763,N_7150,N_6257);
nand U11764 (N_11764,N_8810,N_7803);
or U11765 (N_11765,N_6192,N_8969);
and U11766 (N_11766,N_7753,N_8582);
nor U11767 (N_11767,N_8382,N_8836);
xor U11768 (N_11768,N_7821,N_6907);
or U11769 (N_11769,N_6552,N_7195);
or U11770 (N_11770,N_6444,N_6883);
nor U11771 (N_11771,N_7357,N_6971);
and U11772 (N_11772,N_7547,N_8263);
and U11773 (N_11773,N_8349,N_8862);
or U11774 (N_11774,N_7187,N_7650);
or U11775 (N_11775,N_6851,N_7975);
nor U11776 (N_11776,N_8757,N_8746);
and U11777 (N_11777,N_7935,N_7747);
nor U11778 (N_11778,N_8938,N_7157);
nor U11779 (N_11779,N_8529,N_6550);
and U11780 (N_11780,N_7104,N_8456);
and U11781 (N_11781,N_8675,N_7275);
nor U11782 (N_11782,N_7840,N_6524);
nand U11783 (N_11783,N_8487,N_8332);
nor U11784 (N_11784,N_8510,N_8831);
or U11785 (N_11785,N_7800,N_6211);
and U11786 (N_11786,N_6320,N_8347);
and U11787 (N_11787,N_6952,N_8471);
nor U11788 (N_11788,N_8348,N_8084);
nor U11789 (N_11789,N_6282,N_7605);
and U11790 (N_11790,N_7485,N_6647);
nor U11791 (N_11791,N_6486,N_8462);
and U11792 (N_11792,N_8864,N_7542);
and U11793 (N_11793,N_7448,N_6591);
nor U11794 (N_11794,N_6135,N_6597);
nor U11795 (N_11795,N_8569,N_8381);
nor U11796 (N_11796,N_6299,N_8963);
or U11797 (N_11797,N_8589,N_6200);
or U11798 (N_11798,N_7743,N_7462);
nand U11799 (N_11799,N_7268,N_7500);
and U11800 (N_11800,N_8557,N_7787);
or U11801 (N_11801,N_7302,N_8632);
or U11802 (N_11802,N_8281,N_6485);
or U11803 (N_11803,N_8646,N_6336);
and U11804 (N_11804,N_7863,N_7458);
nand U11805 (N_11805,N_8593,N_6400);
nand U11806 (N_11806,N_6067,N_6520);
nor U11807 (N_11807,N_8082,N_8815);
and U11808 (N_11808,N_7458,N_8657);
or U11809 (N_11809,N_7654,N_8026);
or U11810 (N_11810,N_7954,N_8294);
nand U11811 (N_11811,N_8270,N_8315);
or U11812 (N_11812,N_6850,N_6216);
and U11813 (N_11813,N_6709,N_7021);
or U11814 (N_11814,N_8540,N_8166);
nor U11815 (N_11815,N_7110,N_7727);
or U11816 (N_11816,N_7892,N_7450);
and U11817 (N_11817,N_7640,N_8800);
and U11818 (N_11818,N_7909,N_8327);
and U11819 (N_11819,N_7986,N_6241);
nand U11820 (N_11820,N_6464,N_7985);
or U11821 (N_11821,N_7257,N_7721);
or U11822 (N_11822,N_6907,N_8266);
nor U11823 (N_11823,N_7415,N_7682);
and U11824 (N_11824,N_7746,N_7117);
or U11825 (N_11825,N_6181,N_7217);
nor U11826 (N_11826,N_7406,N_7984);
and U11827 (N_11827,N_7146,N_7630);
nand U11828 (N_11828,N_6277,N_7957);
or U11829 (N_11829,N_6393,N_6581);
or U11830 (N_11830,N_6049,N_6549);
and U11831 (N_11831,N_6059,N_6600);
nand U11832 (N_11832,N_8448,N_6421);
or U11833 (N_11833,N_6895,N_6197);
nand U11834 (N_11834,N_7684,N_8896);
nor U11835 (N_11835,N_6378,N_7455);
and U11836 (N_11836,N_7037,N_7748);
nor U11837 (N_11837,N_8854,N_7025);
nand U11838 (N_11838,N_7487,N_7423);
nand U11839 (N_11839,N_6752,N_6797);
or U11840 (N_11840,N_8428,N_8736);
nor U11841 (N_11841,N_8293,N_6276);
or U11842 (N_11842,N_6082,N_8480);
or U11843 (N_11843,N_6003,N_6137);
nand U11844 (N_11844,N_8496,N_7344);
and U11845 (N_11845,N_8155,N_6347);
nand U11846 (N_11846,N_6473,N_8005);
and U11847 (N_11847,N_6255,N_6007);
or U11848 (N_11848,N_7382,N_7553);
and U11849 (N_11849,N_6203,N_7872);
nand U11850 (N_11850,N_8356,N_7301);
nand U11851 (N_11851,N_8854,N_7821);
nor U11852 (N_11852,N_6820,N_6533);
nor U11853 (N_11853,N_7894,N_8289);
nand U11854 (N_11854,N_6989,N_6144);
or U11855 (N_11855,N_8221,N_8765);
nor U11856 (N_11856,N_6489,N_7494);
nand U11857 (N_11857,N_7046,N_6144);
nand U11858 (N_11858,N_7776,N_6987);
nand U11859 (N_11859,N_6649,N_8590);
and U11860 (N_11860,N_6534,N_8769);
or U11861 (N_11861,N_7885,N_6310);
and U11862 (N_11862,N_7727,N_8215);
or U11863 (N_11863,N_7852,N_7200);
and U11864 (N_11864,N_8564,N_6989);
and U11865 (N_11865,N_6341,N_6205);
nand U11866 (N_11866,N_6773,N_7363);
and U11867 (N_11867,N_8867,N_8172);
and U11868 (N_11868,N_8281,N_7381);
nor U11869 (N_11869,N_8422,N_7788);
xor U11870 (N_11870,N_8805,N_7953);
or U11871 (N_11871,N_8262,N_7961);
nor U11872 (N_11872,N_8557,N_6887);
nand U11873 (N_11873,N_8940,N_7016);
or U11874 (N_11874,N_8750,N_8744);
and U11875 (N_11875,N_7863,N_6227);
or U11876 (N_11876,N_7829,N_7771);
and U11877 (N_11877,N_6648,N_6102);
nand U11878 (N_11878,N_6101,N_8532);
and U11879 (N_11879,N_6242,N_8040);
nor U11880 (N_11880,N_7083,N_8562);
nand U11881 (N_11881,N_7953,N_7039);
nand U11882 (N_11882,N_8419,N_7625);
or U11883 (N_11883,N_8386,N_8534);
nor U11884 (N_11884,N_7478,N_7081);
xor U11885 (N_11885,N_7611,N_7853);
and U11886 (N_11886,N_7456,N_7862);
and U11887 (N_11887,N_7397,N_7450);
and U11888 (N_11888,N_6181,N_8064);
nand U11889 (N_11889,N_7210,N_7186);
xnor U11890 (N_11890,N_8304,N_8308);
nor U11891 (N_11891,N_7400,N_6471);
nor U11892 (N_11892,N_7408,N_8462);
or U11893 (N_11893,N_8850,N_8077);
nor U11894 (N_11894,N_6966,N_8039);
nor U11895 (N_11895,N_7164,N_8618);
and U11896 (N_11896,N_6850,N_7543);
and U11897 (N_11897,N_8911,N_6861);
nand U11898 (N_11898,N_7551,N_7614);
nor U11899 (N_11899,N_7179,N_6204);
nand U11900 (N_11900,N_8050,N_6443);
or U11901 (N_11901,N_7537,N_8273);
and U11902 (N_11902,N_8873,N_7312);
nand U11903 (N_11903,N_8697,N_7511);
nand U11904 (N_11904,N_8796,N_6022);
nor U11905 (N_11905,N_7514,N_7930);
or U11906 (N_11906,N_7548,N_7520);
or U11907 (N_11907,N_8327,N_6162);
or U11908 (N_11908,N_7403,N_8041);
xor U11909 (N_11909,N_7034,N_7197);
and U11910 (N_11910,N_8668,N_7514);
and U11911 (N_11911,N_7142,N_7159);
nor U11912 (N_11912,N_8041,N_6873);
xnor U11913 (N_11913,N_6662,N_6748);
nor U11914 (N_11914,N_7295,N_8905);
xor U11915 (N_11915,N_6419,N_6935);
nand U11916 (N_11916,N_8536,N_6847);
or U11917 (N_11917,N_7486,N_7575);
and U11918 (N_11918,N_7531,N_8831);
xnor U11919 (N_11919,N_7415,N_7626);
nor U11920 (N_11920,N_8491,N_7456);
nand U11921 (N_11921,N_8597,N_6902);
nand U11922 (N_11922,N_8967,N_7804);
xor U11923 (N_11923,N_6074,N_6544);
nor U11924 (N_11924,N_7964,N_7260);
nor U11925 (N_11925,N_6430,N_6486);
or U11926 (N_11926,N_8144,N_6185);
nand U11927 (N_11927,N_8105,N_8167);
nor U11928 (N_11928,N_6715,N_7701);
nand U11929 (N_11929,N_6029,N_7531);
and U11930 (N_11930,N_8572,N_7985);
and U11931 (N_11931,N_8726,N_8398);
nor U11932 (N_11932,N_6844,N_8321);
and U11933 (N_11933,N_8662,N_7137);
and U11934 (N_11934,N_8042,N_7163);
nor U11935 (N_11935,N_6663,N_8565);
nand U11936 (N_11936,N_6747,N_7300);
or U11937 (N_11937,N_8475,N_6868);
and U11938 (N_11938,N_8793,N_6839);
and U11939 (N_11939,N_8921,N_6925);
nor U11940 (N_11940,N_6871,N_7812);
and U11941 (N_11941,N_8087,N_6959);
nor U11942 (N_11942,N_7160,N_6947);
nand U11943 (N_11943,N_7322,N_8363);
or U11944 (N_11944,N_6274,N_7720);
or U11945 (N_11945,N_6479,N_6454);
nor U11946 (N_11946,N_8057,N_6197);
nand U11947 (N_11947,N_8483,N_6024);
and U11948 (N_11948,N_7870,N_6865);
or U11949 (N_11949,N_7727,N_8927);
nor U11950 (N_11950,N_6212,N_6911);
or U11951 (N_11951,N_6199,N_6234);
nand U11952 (N_11952,N_6270,N_8142);
nor U11953 (N_11953,N_7226,N_7364);
nand U11954 (N_11954,N_6706,N_8683);
xor U11955 (N_11955,N_6401,N_8812);
nand U11956 (N_11956,N_7964,N_8122);
nor U11957 (N_11957,N_8316,N_8898);
nand U11958 (N_11958,N_7472,N_8613);
and U11959 (N_11959,N_6748,N_8961);
or U11960 (N_11960,N_6315,N_6894);
nor U11961 (N_11961,N_6518,N_8462);
or U11962 (N_11962,N_8607,N_6397);
and U11963 (N_11963,N_6803,N_7392);
or U11964 (N_11964,N_8871,N_6459);
or U11965 (N_11965,N_8461,N_7899);
and U11966 (N_11966,N_6001,N_6593);
xor U11967 (N_11967,N_7401,N_8578);
nand U11968 (N_11968,N_6772,N_6509);
or U11969 (N_11969,N_7886,N_8498);
nand U11970 (N_11970,N_8771,N_8559);
nor U11971 (N_11971,N_7699,N_6585);
nand U11972 (N_11972,N_8132,N_7257);
and U11973 (N_11973,N_7789,N_8261);
and U11974 (N_11974,N_8175,N_8000);
or U11975 (N_11975,N_7548,N_7211);
nand U11976 (N_11976,N_8594,N_6059);
and U11977 (N_11977,N_6111,N_7933);
and U11978 (N_11978,N_7155,N_6493);
and U11979 (N_11979,N_7169,N_6717);
nand U11980 (N_11980,N_7508,N_7246);
and U11981 (N_11981,N_8159,N_7718);
or U11982 (N_11982,N_7037,N_7264);
nand U11983 (N_11983,N_7209,N_6034);
nand U11984 (N_11984,N_6396,N_7561);
nor U11985 (N_11985,N_7597,N_8420);
nor U11986 (N_11986,N_8000,N_7230);
or U11987 (N_11987,N_6666,N_7181);
and U11988 (N_11988,N_7912,N_7408);
nand U11989 (N_11989,N_7634,N_6415);
nor U11990 (N_11990,N_8746,N_8544);
xnor U11991 (N_11991,N_7019,N_6025);
or U11992 (N_11992,N_6105,N_6233);
nor U11993 (N_11993,N_8478,N_8601);
nor U11994 (N_11994,N_8461,N_7512);
nor U11995 (N_11995,N_6303,N_6912);
or U11996 (N_11996,N_7008,N_6054);
or U11997 (N_11997,N_8674,N_7962);
or U11998 (N_11998,N_6851,N_6444);
and U11999 (N_11999,N_7838,N_8001);
and U12000 (N_12000,N_11015,N_9203);
and U12001 (N_12001,N_9906,N_10058);
nand U12002 (N_12002,N_9517,N_10668);
or U12003 (N_12003,N_11264,N_11886);
nand U12004 (N_12004,N_10967,N_10009);
and U12005 (N_12005,N_9980,N_11004);
or U12006 (N_12006,N_10021,N_9212);
or U12007 (N_12007,N_10913,N_11801);
nor U12008 (N_12008,N_11349,N_10951);
nand U12009 (N_12009,N_9849,N_9874);
or U12010 (N_12010,N_9033,N_11928);
or U12011 (N_12011,N_10977,N_10347);
nor U12012 (N_12012,N_11609,N_11002);
nor U12013 (N_12013,N_11777,N_11547);
and U12014 (N_12014,N_9218,N_11205);
or U12015 (N_12015,N_10811,N_10640);
nand U12016 (N_12016,N_11499,N_9286);
or U12017 (N_12017,N_10428,N_10275);
xor U12018 (N_12018,N_9144,N_10548);
or U12019 (N_12019,N_10720,N_9423);
nor U12020 (N_12020,N_11936,N_10316);
and U12021 (N_12021,N_9532,N_10943);
or U12022 (N_12022,N_10629,N_11644);
or U12023 (N_12023,N_9529,N_10429);
and U12024 (N_12024,N_10826,N_9773);
and U12025 (N_12025,N_10795,N_11857);
and U12026 (N_12026,N_9097,N_10910);
nand U12027 (N_12027,N_9186,N_9544);
nand U12028 (N_12028,N_10060,N_11301);
xor U12029 (N_12029,N_9657,N_11027);
nor U12030 (N_12030,N_10872,N_9655);
and U12031 (N_12031,N_10160,N_10049);
or U12032 (N_12032,N_11241,N_11270);
nand U12033 (N_12033,N_11025,N_9077);
nand U12034 (N_12034,N_11808,N_11505);
nand U12035 (N_12035,N_9567,N_9010);
nand U12036 (N_12036,N_11810,N_11398);
xor U12037 (N_12037,N_10961,N_10442);
and U12038 (N_12038,N_11195,N_10769);
or U12039 (N_12039,N_9954,N_9891);
nand U12040 (N_12040,N_11838,N_11493);
and U12041 (N_12041,N_9949,N_9416);
and U12042 (N_12042,N_9042,N_10713);
or U12043 (N_12043,N_9045,N_9519);
or U12044 (N_12044,N_10878,N_9070);
nor U12045 (N_12045,N_9306,N_9153);
and U12046 (N_12046,N_10023,N_9249);
and U12047 (N_12047,N_9852,N_11321);
nor U12048 (N_12048,N_11334,N_9453);
or U12049 (N_12049,N_9391,N_10241);
nor U12050 (N_12050,N_10088,N_10729);
and U12051 (N_12051,N_9412,N_10156);
nand U12052 (N_12052,N_10935,N_11249);
and U12053 (N_12053,N_11864,N_10902);
and U12054 (N_12054,N_10922,N_11145);
and U12055 (N_12055,N_10243,N_11157);
and U12056 (N_12056,N_10227,N_9679);
nor U12057 (N_12057,N_10999,N_9482);
and U12058 (N_12058,N_9802,N_11440);
nor U12059 (N_12059,N_10360,N_11546);
nand U12060 (N_12060,N_10784,N_11737);
nand U12061 (N_12061,N_11716,N_11039);
and U12062 (N_12062,N_10451,N_10365);
nor U12063 (N_12063,N_9104,N_9041);
or U12064 (N_12064,N_11675,N_10046);
nand U12065 (N_12065,N_11283,N_11688);
and U12066 (N_12066,N_10828,N_9078);
or U12067 (N_12067,N_11481,N_9654);
nand U12068 (N_12068,N_10586,N_10940);
or U12069 (N_12069,N_9316,N_11436);
and U12070 (N_12070,N_9639,N_9673);
or U12071 (N_12071,N_10947,N_10962);
nor U12072 (N_12072,N_11828,N_10276);
and U12073 (N_12073,N_10973,N_9014);
nand U12074 (N_12074,N_9715,N_10186);
or U12075 (N_12075,N_11381,N_11146);
and U12076 (N_12076,N_11405,N_11459);
or U12077 (N_12077,N_9653,N_9812);
and U12078 (N_12078,N_9081,N_10771);
or U12079 (N_12079,N_10105,N_10263);
nand U12080 (N_12080,N_10136,N_11946);
nand U12081 (N_12081,N_11295,N_10081);
and U12082 (N_12082,N_10928,N_10906);
and U12083 (N_12083,N_9707,N_11686);
nor U12084 (N_12084,N_11367,N_10344);
nand U12085 (N_12085,N_11587,N_9119);
nor U12086 (N_12086,N_9926,N_10749);
and U12087 (N_12087,N_10636,N_11066);
or U12088 (N_12088,N_9462,N_9205);
nand U12089 (N_12089,N_11791,N_9513);
nor U12090 (N_12090,N_9016,N_11739);
and U12091 (N_12091,N_9420,N_11939);
or U12092 (N_12092,N_9247,N_9349);
or U12093 (N_12093,N_11319,N_10370);
nor U12094 (N_12094,N_10897,N_11050);
nor U12095 (N_12095,N_9074,N_11412);
nor U12096 (N_12096,N_11140,N_10296);
nor U12097 (N_12097,N_9694,N_11265);
nand U12098 (N_12098,N_11339,N_10268);
and U12099 (N_12099,N_9989,N_10318);
nand U12100 (N_12100,N_11306,N_9115);
or U12101 (N_12101,N_10780,N_10546);
and U12102 (N_12102,N_11384,N_9388);
and U12103 (N_12103,N_11389,N_10917);
nand U12104 (N_12104,N_11707,N_9684);
or U12105 (N_12105,N_11313,N_9151);
nor U12106 (N_12106,N_9063,N_10398);
xnor U12107 (N_12107,N_11409,N_9121);
xnor U12108 (N_12108,N_9711,N_10498);
nand U12109 (N_12109,N_11057,N_11985);
and U12110 (N_12110,N_11151,N_9032);
and U12111 (N_12111,N_11600,N_9035);
and U12112 (N_12112,N_10484,N_11179);
and U12113 (N_12113,N_9739,N_11136);
and U12114 (N_12114,N_9860,N_11294);
nand U12115 (N_12115,N_11997,N_11377);
nand U12116 (N_12116,N_10992,N_10624);
nor U12117 (N_12117,N_10824,N_9375);
and U12118 (N_12118,N_10016,N_9541);
and U12119 (N_12119,N_10787,N_11959);
and U12120 (N_12120,N_9333,N_10882);
nand U12121 (N_12121,N_9187,N_11812);
or U12122 (N_12122,N_11898,N_10687);
nand U12123 (N_12123,N_10474,N_11927);
nand U12124 (N_12124,N_9405,N_11013);
nor U12125 (N_12125,N_9809,N_11322);
and U12126 (N_12126,N_10252,N_10452);
nor U12127 (N_12127,N_10020,N_9551);
or U12128 (N_12128,N_9626,N_9629);
nor U12129 (N_12129,N_10323,N_9433);
nor U12130 (N_12130,N_9856,N_10108);
and U12131 (N_12131,N_10834,N_11636);
and U12132 (N_12132,N_11361,N_9603);
nand U12133 (N_12133,N_11121,N_10114);
nand U12134 (N_12134,N_9426,N_11512);
nor U12135 (N_12135,N_11980,N_11388);
and U12136 (N_12136,N_9220,N_9830);
nand U12137 (N_12137,N_11112,N_9861);
nand U12138 (N_12138,N_11530,N_9263);
and U12139 (N_12139,N_11622,N_11837);
nand U12140 (N_12140,N_9443,N_11841);
and U12141 (N_12141,N_10265,N_10554);
or U12142 (N_12142,N_9120,N_11433);
and U12143 (N_12143,N_11401,N_9368);
nor U12144 (N_12144,N_9646,N_11943);
or U12145 (N_12145,N_11764,N_11047);
and U12146 (N_12146,N_9634,N_9566);
nor U12147 (N_12147,N_11593,N_11703);
xnor U12148 (N_12148,N_9092,N_9067);
or U12149 (N_12149,N_11890,N_10682);
or U12150 (N_12150,N_11494,N_11536);
or U12151 (N_12151,N_10357,N_10424);
nor U12152 (N_12152,N_10532,N_11503);
or U12153 (N_12153,N_9219,N_11244);
and U12154 (N_12154,N_11176,N_11310);
nor U12155 (N_12155,N_9130,N_10255);
or U12156 (N_12156,N_11395,N_10577);
xor U12157 (N_12157,N_11007,N_11803);
nand U12158 (N_12158,N_9757,N_11442);
or U12159 (N_12159,N_9281,N_9387);
nand U12160 (N_12160,N_11059,N_9805);
or U12161 (N_12161,N_9586,N_10773);
or U12162 (N_12162,N_10007,N_10195);
nor U12163 (N_12163,N_10655,N_9876);
nand U12164 (N_12164,N_9733,N_11983);
nand U12165 (N_12165,N_10519,N_10793);
nor U12166 (N_12166,N_11202,N_10813);
nor U12167 (N_12167,N_11895,N_9918);
and U12168 (N_12168,N_9914,N_9300);
xor U12169 (N_12169,N_9013,N_9478);
nand U12170 (N_12170,N_10403,N_11345);
or U12171 (N_12171,N_10753,N_11920);
or U12172 (N_12172,N_9688,N_11460);
and U12173 (N_12173,N_9133,N_10991);
or U12174 (N_12174,N_9952,N_11141);
nor U12175 (N_12175,N_11156,N_11095);
and U12176 (N_12176,N_9438,N_9278);
xor U12177 (N_12177,N_9029,N_9997);
nand U12178 (N_12178,N_10619,N_9641);
and U12179 (N_12179,N_9870,N_9554);
or U12180 (N_12180,N_10697,N_9331);
nor U12181 (N_12181,N_10670,N_11323);
nand U12182 (N_12182,N_11477,N_11563);
and U12183 (N_12183,N_11403,N_10379);
nor U12184 (N_12184,N_11570,N_10236);
or U12185 (N_12185,N_9284,N_10884);
nand U12186 (N_12186,N_11839,N_9038);
or U12187 (N_12187,N_10100,N_10129);
nor U12188 (N_12188,N_9088,N_11844);
or U12189 (N_12189,N_10896,N_11934);
and U12190 (N_12190,N_10775,N_9259);
and U12191 (N_12191,N_11374,N_11250);
xor U12192 (N_12192,N_9742,N_9666);
nand U12193 (N_12193,N_10311,N_9756);
nor U12194 (N_12194,N_11291,N_11019);
nor U12195 (N_12195,N_9789,N_9037);
nand U12196 (N_12196,N_11240,N_9533);
or U12197 (N_12197,N_11260,N_10385);
nand U12198 (N_12198,N_9209,N_9938);
nand U12199 (N_12199,N_10675,N_9040);
nor U12200 (N_12200,N_9486,N_11743);
or U12201 (N_12201,N_11944,N_9882);
xor U12202 (N_12202,N_10639,N_9525);
or U12203 (N_12203,N_11124,N_9524);
nor U12204 (N_12204,N_9647,N_10680);
nand U12205 (N_12205,N_10240,N_9935);
nor U12206 (N_12206,N_9108,N_9008);
or U12207 (N_12207,N_9518,N_10008);
and U12208 (N_12208,N_11128,N_10116);
nor U12209 (N_12209,N_9394,N_9516);
and U12210 (N_12210,N_11282,N_10409);
nor U12211 (N_12211,N_9880,N_11525);
nor U12212 (N_12212,N_11571,N_10730);
or U12213 (N_12213,N_11557,N_10259);
nand U12214 (N_12214,N_9061,N_9815);
nand U12215 (N_12215,N_11598,N_10517);
or U12216 (N_12216,N_10731,N_11788);
nor U12217 (N_12217,N_9776,N_9210);
or U12218 (N_12218,N_10469,N_9528);
and U12219 (N_12219,N_9591,N_10916);
and U12220 (N_12220,N_9840,N_11298);
xnor U12221 (N_12221,N_10281,N_10701);
and U12222 (N_12222,N_10959,N_11624);
or U12223 (N_12223,N_9183,N_10703);
nand U12224 (N_12224,N_9966,N_10950);
nor U12225 (N_12225,N_10396,N_10445);
nor U12226 (N_12226,N_11233,N_11269);
or U12227 (N_12227,N_10974,N_10755);
nor U12228 (N_12228,N_9977,N_10399);
and U12229 (N_12229,N_11211,N_11439);
nand U12230 (N_12230,N_10301,N_11451);
nand U12231 (N_12231,N_10644,N_9582);
nor U12232 (N_12232,N_11560,N_10455);
nor U12233 (N_12233,N_10096,N_9396);
and U12234 (N_12234,N_9879,N_11206);
nand U12235 (N_12235,N_9595,N_10039);
and U12236 (N_12236,N_9777,N_9126);
nor U12237 (N_12237,N_11420,N_11018);
or U12238 (N_12238,N_9139,N_10177);
or U12239 (N_12239,N_10602,N_11474);
nor U12240 (N_12240,N_11664,N_9923);
or U12241 (N_12241,N_10812,N_10918);
or U12242 (N_12242,N_11304,N_11376);
nor U12243 (N_12243,N_11663,N_10339);
nor U12244 (N_12244,N_11346,N_10170);
or U12245 (N_12245,N_11642,N_9577);
nor U12246 (N_12246,N_9251,N_9473);
nand U12247 (N_12247,N_10306,N_11667);
or U12248 (N_12248,N_10605,N_11639);
or U12249 (N_12249,N_10119,N_11520);
nand U12250 (N_12250,N_9283,N_9746);
nand U12251 (N_12251,N_10065,N_11231);
or U12252 (N_12252,N_9147,N_9310);
nand U12253 (N_12253,N_11650,N_9969);
and U12254 (N_12254,N_9837,N_11134);
or U12255 (N_12255,N_11713,N_9542);
and U12256 (N_12256,N_11062,N_9982);
nand U12257 (N_12257,N_9571,N_9208);
nor U12258 (N_12258,N_11511,N_11786);
nand U12259 (N_12259,N_9071,N_9034);
nand U12260 (N_12260,N_11976,N_10791);
nand U12261 (N_12261,N_9995,N_10647);
nor U12262 (N_12262,N_11278,N_9295);
xnor U12263 (N_12263,N_10457,N_9028);
or U12264 (N_12264,N_9617,N_9652);
xnor U12265 (N_12265,N_10262,N_9157);
nand U12266 (N_12266,N_11868,N_10909);
nand U12267 (N_12267,N_10535,N_11252);
or U12268 (N_12268,N_9325,N_10745);
nand U12269 (N_12269,N_10831,N_10657);
nor U12270 (N_12270,N_9811,N_10835);
or U12271 (N_12271,N_9452,N_11613);
and U12272 (N_12272,N_10052,N_10584);
nor U12273 (N_12273,N_9797,N_10401);
nand U12274 (N_12274,N_11101,N_9987);
nor U12275 (N_12275,N_11757,N_9568);
and U12276 (N_12276,N_9668,N_9361);
or U12277 (N_12277,N_9553,N_11931);
or U12278 (N_12278,N_9373,N_11445);
and U12279 (N_12279,N_9143,N_10972);
and U12280 (N_12280,N_10860,N_11251);
or U12281 (N_12281,N_11907,N_9523);
nor U12282 (N_12282,N_9392,N_11776);
and U12283 (N_12283,N_10249,N_10743);
nor U12284 (N_12284,N_9583,N_10271);
and U12285 (N_12285,N_11924,N_9853);
nand U12286 (N_12286,N_10799,N_11834);
or U12287 (N_12287,N_10069,N_11578);
nor U12288 (N_12288,N_9999,N_11726);
or U12289 (N_12289,N_11165,N_10239);
nand U12290 (N_12290,N_9352,N_9522);
nand U12291 (N_12291,N_9890,N_9863);
or U12292 (N_12292,N_10673,N_10971);
or U12293 (N_12293,N_10635,N_11496);
or U12294 (N_12294,N_11872,N_11649);
or U12295 (N_12295,N_9446,N_11399);
or U12296 (N_12296,N_10561,N_9448);
nor U12297 (N_12297,N_11422,N_11161);
nor U12298 (N_12298,N_9044,N_9507);
and U12299 (N_12299,N_10145,N_10213);
nand U12300 (N_12300,N_10198,N_9743);
xnor U12301 (N_12301,N_10381,N_11091);
nand U12302 (N_12302,N_11859,N_11665);
nand U12303 (N_12303,N_9735,N_10801);
nor U12304 (N_12304,N_11977,N_11216);
and U12305 (N_12305,N_10404,N_11333);
xor U12306 (N_12306,N_11080,N_9344);
and U12307 (N_12307,N_11592,N_9217);
or U12308 (N_12308,N_10120,N_11783);
nor U12309 (N_12309,N_11831,N_9998);
or U12310 (N_12310,N_9953,N_11689);
xor U12311 (N_12311,N_10297,N_11109);
or U12312 (N_12312,N_9136,N_10142);
nor U12313 (N_12313,N_11227,N_10707);
nand U12314 (N_12314,N_9576,N_11006);
and U12315 (N_12315,N_11933,N_10865);
nand U12316 (N_12316,N_10643,N_10989);
xor U12317 (N_12317,N_9764,N_11654);
or U12318 (N_12318,N_9332,N_9318);
and U12319 (N_12319,N_10201,N_11540);
xnor U12320 (N_12320,N_10901,N_10110);
nand U12321 (N_12321,N_10969,N_9941);
and U12322 (N_12322,N_9798,N_9992);
or U12323 (N_12323,N_11288,N_11795);
nand U12324 (N_12324,N_10157,N_11880);
nand U12325 (N_12325,N_11212,N_11628);
nand U12326 (N_12326,N_11850,N_10762);
nand U12327 (N_12327,N_10855,N_11660);
or U12328 (N_12328,N_11379,N_10964);
nand U12329 (N_12329,N_11854,N_11698);
or U12330 (N_12330,N_10211,N_11896);
nor U12331 (N_12331,N_10165,N_10842);
and U12332 (N_12332,N_9340,N_9729);
nor U12333 (N_12333,N_10449,N_9500);
nand U12334 (N_12334,N_11465,N_10738);
nand U12335 (N_12335,N_11584,N_11210);
and U12336 (N_12336,N_10509,N_11279);
nor U12337 (N_12337,N_9095,N_9674);
or U12338 (N_12338,N_9640,N_11517);
nor U12339 (N_12339,N_9622,N_10036);
nor U12340 (N_12340,N_11873,N_11461);
and U12341 (N_12341,N_9085,N_10045);
nor U12342 (N_12342,N_9824,N_9925);
and U12343 (N_12343,N_11894,N_10471);
or U12344 (N_12344,N_11117,N_11064);
nand U12345 (N_12345,N_10180,N_11397);
and U12346 (N_12346,N_9197,N_11608);
nand U12347 (N_12347,N_10557,N_11138);
nand U12348 (N_12348,N_10463,N_10514);
or U12349 (N_12349,N_9514,N_9030);
nand U12350 (N_12350,N_9866,N_11352);
xnor U12351 (N_12351,N_9971,N_10139);
or U12352 (N_12352,N_10290,N_10153);
nor U12353 (N_12353,N_9298,N_9003);
nand U12354 (N_12354,N_10540,N_10274);
and U12355 (N_12355,N_10032,N_11965);
or U12356 (N_12356,N_9105,N_9697);
and U12357 (N_12357,N_10544,N_9223);
nor U12358 (N_12358,N_9575,N_10287);
and U12359 (N_12359,N_9842,N_10526);
xor U12360 (N_12360,N_11676,N_10957);
nor U12361 (N_12361,N_10194,N_9341);
nor U12362 (N_12362,N_11234,N_11763);
nand U12363 (N_12363,N_11090,N_10161);
or U12364 (N_12364,N_10233,N_10212);
nand U12365 (N_12365,N_9555,N_10015);
nor U12366 (N_12366,N_10374,N_9459);
xor U12367 (N_12367,N_10770,N_11324);
nor U12368 (N_12368,N_9226,N_11428);
or U12369 (N_12369,N_11070,N_11094);
nand U12370 (N_12370,N_10847,N_10123);
nand U12371 (N_12371,N_11558,N_11438);
and U12372 (N_12372,N_11341,N_10664);
nand U12373 (N_12373,N_9921,N_9176);
nand U12374 (N_12374,N_11790,N_11149);
or U12375 (N_12375,N_10234,N_10353);
nand U12376 (N_12376,N_9169,N_9950);
nand U12377 (N_12377,N_9896,N_11652);
nor U12378 (N_12378,N_10545,N_9023);
and U12379 (N_12379,N_9312,N_11378);
nor U12380 (N_12380,N_11537,N_10927);
or U12381 (N_12381,N_11552,N_10543);
and U12382 (N_12382,N_10313,N_10141);
nor U12383 (N_12383,N_11522,N_10012);
or U12384 (N_12384,N_10516,N_11147);
nor U12385 (N_12385,N_11605,N_9470);
and U12386 (N_12386,N_9948,N_10871);
nand U12387 (N_12387,N_10574,N_9821);
nor U12388 (N_12388,N_11975,N_10754);
nand U12389 (N_12389,N_11132,N_10616);
and U12390 (N_12390,N_11960,N_10846);
and U12391 (N_12391,N_10696,N_10070);
or U12392 (N_12392,N_10623,N_10302);
nand U12393 (N_12393,N_10090,N_11286);
nor U12394 (N_12394,N_11340,N_11887);
nor U12395 (N_12395,N_9053,N_9690);
nor U12396 (N_12396,N_11498,N_9850);
nor U12397 (N_12397,N_11023,N_11296);
nor U12398 (N_12398,N_10143,N_11350);
nand U12399 (N_12399,N_9436,N_11708);
xor U12400 (N_12400,N_11060,N_11866);
nand U12401 (N_12401,N_10852,N_9774);
nand U12402 (N_12402,N_9763,N_9540);
nand U12403 (N_12403,N_11507,N_11317);
nor U12404 (N_12404,N_10102,N_9745);
nand U12405 (N_12405,N_9080,N_11072);
nor U12406 (N_12406,N_9844,N_9868);
nand U12407 (N_12407,N_11549,N_9857);
nand U12408 (N_12408,N_9785,N_11787);
nor U12409 (N_12409,N_10218,N_9211);
and U12410 (N_12410,N_9499,N_11266);
nand U12411 (N_12411,N_10440,N_11368);
and U12412 (N_12412,N_11115,N_9432);
nand U12413 (N_12413,N_11579,N_9350);
nor U12414 (N_12414,N_9000,N_10541);
nor U12415 (N_12415,N_11355,N_9910);
nand U12416 (N_12416,N_9963,N_9796);
or U12417 (N_12417,N_9727,N_10341);
nor U12418 (N_12418,N_11103,N_11012);
or U12419 (N_12419,N_11423,N_10465);
nand U12420 (N_12420,N_10948,N_10373);
and U12421 (N_12421,N_11394,N_10216);
nand U12422 (N_12422,N_9930,N_10209);
and U12423 (N_12423,N_11483,N_9501);
nand U12424 (N_12424,N_10406,N_10372);
nor U12425 (N_12425,N_11926,N_9710);
nor U12426 (N_12426,N_9002,N_11921);
nand U12427 (N_12427,N_10470,N_10077);
nor U12428 (N_12428,N_10003,N_11524);
nand U12429 (N_12429,N_11691,N_11848);
and U12430 (N_12430,N_9348,N_10072);
nor U12431 (N_12431,N_11447,N_11443);
and U12432 (N_12432,N_10646,N_9703);
nand U12433 (N_12433,N_10258,N_10614);
nor U12434 (N_12434,N_9813,N_10053);
or U12435 (N_12435,N_10400,N_10024);
nor U12436 (N_12436,N_10589,N_11198);
nand U12437 (N_12437,N_11556,N_11169);
nor U12438 (N_12438,N_10037,N_10576);
nor U12439 (N_12439,N_10472,N_10923);
nand U12440 (N_12440,N_9267,N_11318);
and U12441 (N_12441,N_11135,N_9939);
nand U12442 (N_12442,N_11534,N_11327);
nor U12443 (N_12443,N_9826,N_11935);
or U12444 (N_12444,N_10609,N_11220);
nand U12445 (N_12445,N_10479,N_9322);
nor U12446 (N_12446,N_10818,N_10611);
nor U12447 (N_12447,N_11596,N_9454);
nor U12448 (N_12448,N_11017,N_9810);
nand U12449 (N_12449,N_11336,N_9965);
and U12450 (N_12450,N_9353,N_11771);
nand U12451 (N_12451,N_9804,N_10591);
or U12452 (N_12452,N_11998,N_11792);
and U12453 (N_12453,N_9200,N_11919);
nand U12454 (N_12454,N_11245,N_11464);
and U12455 (N_12455,N_10529,N_10308);
and U12456 (N_12456,N_10987,N_10908);
xnor U12457 (N_12457,N_10757,N_9851);
nand U12458 (N_12458,N_9122,N_10531);
nand U12459 (N_12459,N_9932,N_9427);
or U12460 (N_12460,N_10245,N_11102);
nand U12461 (N_12461,N_11554,N_9545);
nor U12462 (N_12462,N_9422,N_10111);
and U12463 (N_12463,N_10778,N_11818);
and U12464 (N_12464,N_10420,N_11865);
and U12465 (N_12465,N_10331,N_11166);
nor U12466 (N_12466,N_9605,N_10988);
or U12467 (N_12467,N_11670,N_9548);
xor U12468 (N_12468,N_9994,N_10002);
or U12469 (N_12469,N_10953,N_11200);
or U12470 (N_12470,N_9457,N_10558);
xnor U12471 (N_12471,N_11375,N_9667);
nor U12472 (N_12472,N_10966,N_10315);
and U12473 (N_12473,N_9580,N_10392);
and U12474 (N_12474,N_11967,N_9321);
nor U12475 (N_12475,N_9645,N_11001);
and U12476 (N_12476,N_9201,N_9164);
and U12477 (N_12477,N_10975,N_11480);
xnor U12478 (N_12478,N_10314,N_9556);
nor U12479 (N_12479,N_9409,N_9117);
nand U12480 (N_12480,N_11833,N_10718);
or U12481 (N_12481,N_9794,N_9708);
and U12482 (N_12482,N_11988,N_11116);
and U12483 (N_12483,N_10340,N_10995);
nor U12484 (N_12484,N_11038,N_11823);
nand U12485 (N_12485,N_10683,N_11470);
and U12486 (N_12486,N_11621,N_11954);
or U12487 (N_12487,N_9942,N_11566);
and U12488 (N_12488,N_11261,N_9159);
nor U12489 (N_12489,N_11213,N_9466);
nand U12490 (N_12490,N_11574,N_10464);
nor U12491 (N_12491,N_10772,N_11947);
nor U12492 (N_12492,N_11760,N_9455);
or U12493 (N_12493,N_10562,N_11427);
and U12494 (N_12494,N_10175,N_10924);
or U12495 (N_12495,N_9335,N_9717);
nor U12496 (N_12496,N_10330,N_11819);
nor U12497 (N_12497,N_9007,N_9277);
and U12498 (N_12498,N_9246,N_9364);
and U12499 (N_12499,N_9195,N_11604);
or U12500 (N_12500,N_11674,N_9878);
or U12501 (N_12501,N_11658,N_9698);
and U12502 (N_12502,N_9451,N_10494);
or U12503 (N_12503,N_9598,N_9425);
nor U12504 (N_12504,N_9728,N_11131);
or U12505 (N_12505,N_11731,N_10740);
or U12506 (N_12506,N_11254,N_9628);
nand U12507 (N_12507,N_9682,N_10886);
nor U12508 (N_12508,N_9407,N_10080);
nor U12509 (N_12509,N_11230,N_9428);
nor U12510 (N_12510,N_10349,N_9530);
nor U12511 (N_12511,N_9893,N_10607);
or U12512 (N_12512,N_10719,N_10618);
nand U12513 (N_12513,N_11187,N_10615);
xor U12514 (N_12514,N_11178,N_11893);
and U12515 (N_12515,N_10407,N_10527);
nor U12516 (N_12516,N_11292,N_11449);
or U12517 (N_12517,N_11561,N_11223);
and U12518 (N_12518,N_11785,N_9398);
or U12519 (N_12519,N_10383,N_9858);
or U12520 (N_12520,N_9846,N_10027);
or U12521 (N_12521,N_9146,N_10371);
and U12522 (N_12522,N_9975,N_10497);
or U12523 (N_12523,N_10863,N_10106);
or U12524 (N_12524,N_10760,N_10642);
or U12525 (N_12525,N_11901,N_11431);
nand U12526 (N_12526,N_11130,N_11542);
or U12527 (N_12527,N_9477,N_10931);
nor U12528 (N_12528,N_9661,N_10728);
nand U12529 (N_12529,N_10246,N_10343);
nor U12530 (N_12530,N_9520,N_11454);
or U12531 (N_12531,N_10706,N_9389);
and U12532 (N_12532,N_9747,N_11402);
xor U12533 (N_12533,N_9957,N_9260);
or U12534 (N_12534,N_9493,N_11577);
nand U12535 (N_12535,N_11247,N_10149);
nor U12536 (N_12536,N_9149,N_10571);
nand U12537 (N_12537,N_10700,N_9606);
nor U12538 (N_12538,N_9103,N_10648);
and U12539 (N_12539,N_9922,N_9314);
nand U12540 (N_12540,N_11906,N_10487);
xor U12541 (N_12541,N_11168,N_11661);
or U12542 (N_12542,N_9637,N_10205);
nand U12543 (N_12543,N_11243,N_10152);
or U12544 (N_12544,N_10125,N_9463);
or U12545 (N_12545,N_11816,N_11041);
nand U12546 (N_12546,N_9456,N_9700);
or U12547 (N_12547,N_9589,N_11827);
nand U12548 (N_12548,N_9892,N_9806);
or U12549 (N_12549,N_11366,N_10176);
nand U12550 (N_12550,N_10768,N_11863);
or U12551 (N_12551,N_10051,N_10892);
and U12552 (N_12552,N_10217,N_10395);
and U12553 (N_12553,N_11780,N_11074);
and U12554 (N_12554,N_11773,N_11633);
nand U12555 (N_12555,N_9073,N_9549);
or U12556 (N_12556,N_9687,N_10355);
and U12557 (N_12557,N_9231,N_9358);
xor U12558 (N_12558,N_11765,N_10521);
and U12559 (N_12559,N_10253,N_10984);
and U12560 (N_12560,N_11905,N_10716);
or U12561 (N_12561,N_10098,N_10503);
or U12562 (N_12562,N_11748,N_10665);
nand U12563 (N_12563,N_10364,N_10836);
nand U12564 (N_12564,N_9370,N_11990);
nor U12565 (N_12565,N_9736,N_11516);
and U12566 (N_12566,N_10441,N_11910);
nor U12567 (N_12567,N_11413,N_9511);
nor U12568 (N_12568,N_9170,N_9887);
and U12569 (N_12569,N_10759,N_10530);
nand U12570 (N_12570,N_9955,N_10490);
or U12571 (N_12571,N_9495,N_11750);
or U12572 (N_12572,N_11616,N_11365);
or U12573 (N_12573,N_10534,N_10288);
nor U12574 (N_12574,N_11815,N_10324);
nor U12575 (N_12575,N_10278,N_11048);
nand U12576 (N_12576,N_9280,N_11991);
nor U12577 (N_12577,N_9109,N_10229);
and U12578 (N_12578,N_9384,N_11159);
and U12579 (N_12579,N_10030,N_10256);
nand U12580 (N_12580,N_9920,N_11559);
or U12581 (N_12581,N_9258,N_10013);
nand U12582 (N_12582,N_9397,N_10468);
nor U12583 (N_12583,N_11183,N_9497);
or U12584 (N_12584,N_9761,N_11606);
and U12585 (N_12585,N_9188,N_11089);
nand U12586 (N_12586,N_10466,N_10210);
and U12587 (N_12587,N_10504,N_9440);
nand U12588 (N_12588,N_11016,N_10815);
nand U12589 (N_12589,N_11271,N_11918);
and U12590 (N_12590,N_11419,N_9967);
and U12591 (N_12591,N_10934,N_11607);
nor U12592 (N_12592,N_9399,N_10669);
nand U12593 (N_12593,N_11680,N_11802);
nand U12594 (N_12594,N_9945,N_11805);
and U12595 (N_12595,N_11582,N_11637);
nand U12596 (N_12596,N_9276,N_9616);
or U12597 (N_12597,N_10654,N_10875);
and U12598 (N_12598,N_9415,N_9928);
or U12599 (N_12599,N_11741,N_9828);
and U12600 (N_12600,N_11036,N_11862);
nand U12601 (N_12601,N_9791,N_11031);
and U12602 (N_12602,N_9885,N_9574);
or U12603 (N_12603,N_10300,N_11035);
nor U12604 (N_12604,N_10478,N_10499);
nand U12605 (N_12605,N_11881,N_9515);
nor U12606 (N_12606,N_10378,N_9235);
nand U12607 (N_12607,N_9302,N_9770);
nor U12608 (N_12608,N_11441,N_11701);
nand U12609 (N_12609,N_11902,N_9600);
or U12610 (N_12610,N_10617,N_10715);
or U12611 (N_12611,N_9778,N_11372);
nand U12612 (N_12612,N_11185,N_11751);
or U12613 (N_12613,N_11953,N_11297);
nand U12614 (N_12614,N_11585,N_10781);
xor U12615 (N_12615,N_9241,N_9148);
nand U12616 (N_12616,N_11127,N_11753);
nor U12617 (N_12617,N_11065,N_10949);
nor U12618 (N_12618,N_11793,N_10518);
nor U12619 (N_12619,N_10461,N_10097);
or U12620 (N_12620,N_11719,N_9052);
and U12621 (N_12621,N_11672,N_10926);
or U12622 (N_12622,N_10079,N_11514);
nand U12623 (N_12623,N_10849,N_9199);
nor U12624 (N_12624,N_9716,N_10031);
and U12625 (N_12625,N_9469,N_10725);
and U12626 (N_12626,N_10402,N_11014);
or U12627 (N_12627,N_11312,N_11029);
nand U12628 (N_12628,N_10193,N_11817);
and U12629 (N_12629,N_10393,N_11343);
nand U12630 (N_12630,N_10853,N_10423);
and U12631 (N_12631,N_11067,N_9083);
and U12632 (N_12632,N_9604,N_11821);
nand U12633 (N_12633,N_11214,N_11899);
nor U12634 (N_12634,N_11369,N_9198);
nand U12635 (N_12635,N_9867,N_10197);
nor U12636 (N_12636,N_10155,N_11876);
nand U12637 (N_12637,N_9632,N_9021);
and U12638 (N_12638,N_10181,N_11603);
or U12639 (N_12639,N_11623,N_9380);
or U12640 (N_12640,N_9292,N_9274);
nor U12641 (N_12641,N_10628,N_9897);
and U12642 (N_12642,N_9725,N_10397);
nand U12643 (N_12643,N_9547,N_11945);
and U12644 (N_12644,N_9369,N_9383);
nor U12645 (N_12645,N_9173,N_9196);
or U12646 (N_12646,N_11256,N_9327);
nand U12647 (N_12647,N_9584,N_10590);
nor U12648 (N_12648,N_11677,N_11425);
or U12649 (N_12649,N_9245,N_9124);
nand U12650 (N_12650,N_9419,N_11342);
and U12651 (N_12651,N_11885,N_9505);
nand U12652 (N_12652,N_11575,N_11527);
nand U12653 (N_12653,N_10270,N_10981);
or U12654 (N_12654,N_11075,N_11738);
or U12655 (N_12655,N_10238,N_10620);
and U12656 (N_12656,N_9678,N_9702);
nor U12657 (N_12657,N_11925,N_11434);
nand U12658 (N_12658,N_10893,N_10085);
nor U12659 (N_12659,N_10130,N_9787);
or U12660 (N_12660,N_11594,N_11192);
nand U12661 (N_12661,N_10220,N_9114);
and U12662 (N_12662,N_10645,N_11174);
or U12663 (N_12663,N_10547,N_9229);
nor U12664 (N_12664,N_11989,N_11982);
nand U12665 (N_12665,N_11647,N_11962);
and U12666 (N_12666,N_11188,N_9672);
nor U12667 (N_12667,N_10333,N_11937);
nand U12668 (N_12668,N_11614,N_10492);
or U12669 (N_12669,N_9434,N_10633);
nor U12670 (N_12670,N_10507,N_10358);
or U12671 (N_12671,N_11706,N_10879);
nand U12672 (N_12672,N_11853,N_11122);
xnor U12673 (N_12673,N_9834,N_11509);
nor U12674 (N_12674,N_11456,N_10336);
nor U12675 (N_12675,N_10312,N_9253);
or U12676 (N_12676,N_9376,N_10764);
nand U12677 (N_12677,N_10208,N_10215);
nor U12678 (N_12678,N_11635,N_11835);
and U12679 (N_12679,N_9346,N_10954);
nor U12680 (N_12680,N_10226,N_10641);
nand U12681 (N_12681,N_10418,N_9270);
nand U12682 (N_12682,N_9190,N_11900);
and U12683 (N_12683,N_9110,N_9573);
and U12684 (N_12684,N_9755,N_10733);
nand U12685 (N_12685,N_11662,N_9512);
nor U12686 (N_12686,N_10785,N_10056);
nor U12687 (N_12687,N_11497,N_10783);
and U12688 (N_12688,N_10979,N_10539);
or U12689 (N_12689,N_11555,N_9731);
or U12690 (N_12690,N_10608,N_10280);
nand U12691 (N_12691,N_9102,N_10870);
nor U12692 (N_12692,N_10978,N_11468);
or U12693 (N_12693,N_11970,N_9001);
and U12694 (N_12694,N_11330,N_10866);
nand U12695 (N_12695,N_11797,N_11385);
or U12696 (N_12696,N_10598,N_11867);
or U12697 (N_12697,N_9521,N_11186);
or U12698 (N_12698,N_10659,N_10171);
nor U12699 (N_12699,N_11589,N_9509);
and U12700 (N_12700,N_9011,N_11508);
and U12701 (N_12701,N_10076,N_10985);
and U12702 (N_12702,N_11519,N_9101);
or U12703 (N_12703,N_11472,N_11583);
and U12704 (N_12704,N_9202,N_11693);
and U12705 (N_12705,N_10078,N_10025);
and U12706 (N_12706,N_9820,N_9162);
nor U12707 (N_12707,N_10382,N_9768);
nor U12708 (N_12708,N_9360,N_10174);
and U12709 (N_12709,N_11302,N_9712);
and U12710 (N_12710,N_9754,N_10495);
and U12711 (N_12711,N_10612,N_9172);
nand U12712 (N_12712,N_10501,N_11999);
nor U12713 (N_12713,N_10004,N_10101);
or U12714 (N_12714,N_10094,N_9597);
and U12715 (N_12715,N_10282,N_9326);
and U12716 (N_12716,N_10711,N_10091);
nand U12717 (N_12717,N_11932,N_10083);
nor U12718 (N_12718,N_10695,N_9911);
or U12719 (N_12719,N_9753,N_9875);
or U12720 (N_12720,N_9658,N_11028);
nand U12721 (N_12721,N_9683,N_9429);
and U12722 (N_12722,N_11126,N_11526);
or U12723 (N_12723,N_11581,N_10942);
nor U12724 (N_12724,N_11300,N_9961);
or U12725 (N_12725,N_11332,N_11718);
and U12726 (N_12726,N_9086,N_9585);
xnor U12727 (N_12727,N_9907,N_9113);
nor U12728 (N_12728,N_10794,N_11337);
or U12729 (N_12729,N_11201,N_10792);
nand U12730 (N_12730,N_9884,N_11155);
or U12731 (N_12731,N_10377,N_9401);
nand U12732 (N_12732,N_11085,N_11215);
nor U12733 (N_12733,N_11889,N_9612);
nor U12734 (N_12734,N_11150,N_10858);
nor U12735 (N_12735,N_10103,N_11453);
or U12736 (N_12736,N_9006,N_9165);
nand U12737 (N_12737,N_9330,N_11908);
nor U12738 (N_12738,N_11160,N_10427);
and U12739 (N_12739,N_11408,N_10059);
nor U12740 (N_12740,N_10167,N_11551);
or U12741 (N_12741,N_9602,N_9472);
nor U12742 (N_12742,N_11285,N_10196);
and U12743 (N_12743,N_9623,N_11204);
nor U12744 (N_12744,N_10437,N_11504);
nand U12745 (N_12745,N_10414,N_9758);
or U12746 (N_12746,N_9618,N_9250);
and U12747 (N_12747,N_10997,N_10915);
or U12748 (N_12748,N_9100,N_11118);
and U12749 (N_12749,N_9015,N_10260);
and U12750 (N_12750,N_11891,N_11034);
nand U12751 (N_12751,N_11010,N_10285);
or U12752 (N_12752,N_10325,N_11715);
and U12753 (N_12753,N_9624,N_10159);
and U12754 (N_12754,N_9154,N_11040);
nand U12755 (N_12755,N_11011,N_9301);
and U12756 (N_12756,N_11320,N_10447);
and U12757 (N_12757,N_10084,N_11772);
nor U12758 (N_12758,N_9243,N_9379);
nand U12759 (N_12759,N_9257,N_11189);
or U12760 (N_12760,N_11197,N_10638);
or U12761 (N_12761,N_9898,N_9854);
nand U12762 (N_12762,N_10816,N_10837);
and U12763 (N_12763,N_9651,N_9779);
or U12764 (N_12764,N_10237,N_10435);
nand U12765 (N_12765,N_10073,N_11964);
nand U12766 (N_12766,N_11380,N_10678);
and U12767 (N_12767,N_9413,N_10421);
or U12768 (N_12768,N_10786,N_10726);
nand U12769 (N_12769,N_9468,N_10968);
or U12770 (N_12770,N_10485,N_11851);
or U12771 (N_12771,N_9160,N_9089);
and U12772 (N_12772,N_10874,N_9307);
nand U12773 (N_12773,N_9442,N_10880);
or U12774 (N_12774,N_9663,N_10187);
and U12775 (N_12775,N_9638,N_9385);
and U12776 (N_12776,N_11699,N_10721);
nand U12777 (N_12777,N_10476,N_10830);
nand U12778 (N_12778,N_9627,N_9762);
or U12779 (N_12779,N_10304,N_11915);
and U12780 (N_12780,N_9271,N_10838);
nor U12781 (N_12781,N_10568,N_11284);
or U12782 (N_12782,N_10767,N_10790);
nand U12783 (N_12783,N_9940,N_9025);
nand U12784 (N_12784,N_11564,N_10299);
or U12785 (N_12785,N_11452,N_10335);
nand U12786 (N_12786,N_9546,N_11709);
and U12787 (N_12787,N_10462,N_11569);
and U12788 (N_12788,N_9182,N_11722);
and U12789 (N_12789,N_9783,N_10192);
nor U12790 (N_12790,N_10182,N_9024);
and U12791 (N_12791,N_9978,N_11255);
and U12792 (N_12792,N_9901,N_10074);
xor U12793 (N_12793,N_9252,N_10899);
and U12794 (N_12794,N_9099,N_10634);
or U12795 (N_12795,N_10907,N_9780);
nand U12796 (N_12796,N_10829,N_9781);
or U12797 (N_12797,N_11721,N_9976);
or U12798 (N_12798,N_11228,N_11775);
nor U12799 (N_12799,N_9215,N_11154);
nor U12800 (N_12800,N_9635,N_9607);
and U12801 (N_12801,N_10844,N_11049);
nor U12802 (N_12802,N_11779,N_11725);
nor U12803 (N_12803,N_10266,N_10348);
nor U12804 (N_12804,N_9899,N_11287);
nor U12805 (N_12805,N_11360,N_10553);
or U12806 (N_12806,N_9204,N_11110);
nor U12807 (N_12807,N_9750,N_11125);
and U12808 (N_12808,N_10267,N_10134);
nand U12809 (N_12809,N_10298,N_9069);
nor U12810 (N_12810,N_11455,N_11759);
and U12811 (N_12811,N_10888,N_11640);
and U12812 (N_12812,N_9734,N_11359);
nand U12813 (N_12813,N_10825,N_11590);
and U12814 (N_12814,N_9990,N_10164);
nor U12815 (N_12815,N_11673,N_10861);
and U12816 (N_12816,N_11922,N_11770);
and U12817 (N_12817,N_9290,N_10709);
nor U12818 (N_12818,N_9272,N_11364);
or U12819 (N_12819,N_9004,N_11129);
or U12820 (N_12820,N_9587,N_11437);
nor U12821 (N_12821,N_9931,N_9788);
nor U12822 (N_12822,N_10986,N_10214);
and U12823 (N_12823,N_10413,N_10202);
and U12824 (N_12824,N_11177,N_9959);
nor U12825 (N_12825,N_11754,N_10087);
and U12826 (N_12826,N_11407,N_10505);
and U12827 (N_12827,N_10765,N_9418);
or U12828 (N_12828,N_9564,N_9299);
and U12829 (N_12829,N_9670,N_11463);
and U12830 (N_12830,N_9740,N_11711);
nand U12831 (N_12831,N_10674,N_10699);
and U12832 (N_12832,N_10146,N_11798);
or U12833 (N_12833,N_11217,N_9150);
or U12834 (N_12834,N_11978,N_11576);
and U12835 (N_12835,N_9166,N_10154);
nor U12836 (N_12836,N_10150,N_9018);
nor U12837 (N_12837,N_11500,N_9904);
and U12838 (N_12838,N_10168,N_11601);
and U12839 (N_12839,N_9973,N_9508);
and U12840 (N_12840,N_11383,N_11356);
or U12841 (N_12841,N_10843,N_11353);
nand U12842 (N_12842,N_9951,N_9458);
or U12843 (N_12843,N_9288,N_10320);
nand U12844 (N_12844,N_9686,N_9347);
and U12845 (N_12845,N_10579,N_9917);
nand U12846 (N_12846,N_11695,N_9382);
or U12847 (N_12847,N_10677,N_9615);
or U12848 (N_12848,N_9693,N_10895);
nand U12849 (N_12849,N_9179,N_11714);
nand U12850 (N_12850,N_9471,N_10556);
nand U12851 (N_12851,N_9527,N_11104);
and U12852 (N_12852,N_10511,N_10019);
nor U12853 (N_12853,N_11942,N_10774);
nand U12854 (N_12854,N_10712,N_9881);
and U12855 (N_12855,N_9072,N_9264);
and U12856 (N_12856,N_10185,N_11591);
and U12857 (N_12857,N_11535,N_9135);
nand U12858 (N_12858,N_11171,N_11479);
and U12859 (N_12859,N_9793,N_10292);
or U12860 (N_12860,N_11024,N_9234);
nand U12861 (N_12861,N_9817,N_10805);
nand U12862 (N_12862,N_9662,N_11646);
and U12863 (N_12863,N_11084,N_11148);
and U12864 (N_12864,N_10944,N_10273);
or U12865 (N_12865,N_10563,N_11730);
nor U12866 (N_12866,N_11051,N_10005);
xnor U12867 (N_12867,N_11539,N_11488);
nor U12868 (N_12868,N_9760,N_11411);
and U12869 (N_12869,N_9833,N_9506);
or U12870 (N_12870,N_9191,N_10722);
nand U12871 (N_12871,N_9060,N_9094);
nor U12872 (N_12872,N_9558,N_10506);
nor U12873 (N_12873,N_9228,N_10067);
and U12874 (N_12874,N_11973,N_9066);
and U12875 (N_12875,N_9504,N_10089);
nand U12876 (N_12876,N_11232,N_11248);
nand U12877 (N_12877,N_10600,N_11467);
and U12878 (N_12878,N_9137,N_10434);
and U12879 (N_12879,N_9648,N_9282);
and U12880 (N_12880,N_11246,N_9562);
or U12881 (N_12881,N_10391,N_10894);
nor U12882 (N_12882,N_9181,N_11163);
or U12883 (N_12883,N_9578,N_11870);
or U12884 (N_12884,N_11184,N_9561);
nand U12885 (N_12885,N_9979,N_11705);
nor U12886 (N_12886,N_11756,N_11523);
nand U12887 (N_12887,N_9404,N_10279);
and U12888 (N_12888,N_10533,N_9378);
nor U12889 (N_12889,N_9972,N_11518);
nand U12890 (N_12890,N_9633,N_11329);
nor U12891 (N_12891,N_11774,N_11392);
or U12892 (N_12892,N_10459,N_11972);
and U12893 (N_12893,N_10436,N_11700);
and U12894 (N_12894,N_10779,N_9116);
nor U12895 (N_12895,N_9536,N_9650);
nor U12896 (N_12896,N_11842,N_10068);
nor U12897 (N_12897,N_9795,N_10334);
and U12898 (N_12898,N_10172,N_10235);
and U12899 (N_12899,N_10809,N_9611);
nand U12900 (N_12900,N_11796,N_11694);
or U12901 (N_12901,N_10685,N_11631);
and U12902 (N_12902,N_11133,N_11955);
and U12903 (N_12903,N_9129,N_9649);
nor U12904 (N_12904,N_11897,N_10033);
and U12905 (N_12905,N_11299,N_10735);
nand U12906 (N_12906,N_10660,N_9588);
or U12907 (N_12907,N_10822,N_11435);
nor U12908 (N_12908,N_11450,N_11096);
nor U12909 (N_12909,N_11846,N_10204);
or U12910 (N_12910,N_9929,N_9185);
nor U12911 (N_12911,N_11446,N_11820);
or U12912 (N_12912,N_9784,N_9665);
or U12913 (N_12913,N_11855,N_10876);
nor U12914 (N_12914,N_10921,N_10512);
or U12915 (N_12915,N_10929,N_11417);
and U12916 (N_12916,N_11565,N_11669);
nand U12917 (N_12917,N_11325,N_9214);
and U12918 (N_12918,N_11533,N_10310);
and U12919 (N_12919,N_9475,N_9134);
nor U12920 (N_12920,N_11903,N_10454);
nor U12921 (N_12921,N_10135,N_10859);
nor U12922 (N_12922,N_11697,N_10121);
and U12923 (N_12923,N_11789,N_10883);
nor U12924 (N_12924,N_10970,N_9381);
nor U12925 (N_12925,N_10158,N_9479);
and U12926 (N_12926,N_11348,N_11257);
and U12927 (N_12927,N_10789,N_11046);
nor U12928 (N_12928,N_11263,N_10128);
or U12929 (N_12929,N_10133,N_9090);
or U12930 (N_12930,N_9933,N_9909);
or U12931 (N_12931,N_9417,N_11755);
or U12932 (N_12932,N_10840,N_11548);
nand U12933 (N_12933,N_10993,N_9393);
nand U12934 (N_12934,N_9800,N_11487);
or U12935 (N_12935,N_10093,N_9769);
and U12936 (N_12936,N_10063,N_10580);
and U12937 (N_12937,N_10649,N_11458);
nand U12938 (N_12938,N_9184,N_9142);
and U12939 (N_12939,N_9131,N_10329);
or U12940 (N_12940,N_10148,N_11949);
and U12941 (N_12941,N_11811,N_10751);
nand U12942 (N_12942,N_10651,N_10604);
and U12943 (N_12943,N_11729,N_10368);
or U12944 (N_12944,N_9819,N_9465);
or U12945 (N_12945,N_9993,N_10332);
xnor U12946 (N_12946,N_9079,N_11836);
or U12947 (N_12947,N_11822,N_9356);
nor U12948 (N_12948,N_9807,N_11651);
and U12949 (N_12949,N_11105,N_10676);
nor U12950 (N_12950,N_11088,N_11077);
and U12951 (N_12951,N_11501,N_9675);
nand U12952 (N_12952,N_11275,N_11612);
or U12953 (N_12953,N_10958,N_11963);
or U12954 (N_12954,N_10572,N_10467);
or U12955 (N_12955,N_9503,N_11021);
or U12956 (N_12956,N_10508,N_10748);
nand U12957 (N_12957,N_9403,N_11869);
and U12958 (N_12958,N_10862,N_11767);
nand U12959 (N_12959,N_10588,N_10803);
nand U12960 (N_12960,N_9236,N_11416);
or U12961 (N_12961,N_11830,N_9118);
and U12962 (N_12962,N_10307,N_11825);
nand U12963 (N_12963,N_9752,N_11641);
or U12964 (N_12964,N_11181,N_10188);
nand U12965 (N_12965,N_10147,N_11806);
nor U12966 (N_12966,N_10937,N_10387);
nor U12967 (N_12967,N_10050,N_10939);
nand U12968 (N_12968,N_9339,N_10679);
and U12969 (N_12969,N_9319,N_11638);
or U12970 (N_12970,N_9996,N_11111);
nand U12971 (N_12971,N_11098,N_10113);
and U12972 (N_12972,N_9464,N_9790);
or U12973 (N_12973,N_10848,N_10477);
or U12974 (N_12974,N_9986,N_11475);
nor U12975 (N_12975,N_10489,N_9526);
nor U12976 (N_12976,N_9937,N_9488);
or U12977 (N_12977,N_9991,N_9213);
and U12978 (N_12978,N_10802,N_9916);
nor U12979 (N_12979,N_10596,N_11054);
nand U12980 (N_12980,N_11164,N_9098);
and U12981 (N_12981,N_9227,N_11506);
nand U12982 (N_12982,N_11766,N_9424);
and U12983 (N_12983,N_9230,N_11347);
and U12984 (N_12984,N_10369,N_10248);
nand U12985 (N_12985,N_9981,N_11370);
or U12986 (N_12986,N_11562,N_11550);
nand U12987 (N_12987,N_10362,N_10191);
nand U12988 (N_12988,N_10173,N_9046);
nor U12989 (N_12989,N_9767,N_11882);
nand U12990 (N_12990,N_9766,N_10806);
nand U12991 (N_12991,N_11746,N_11107);
nor U12992 (N_12992,N_10996,N_9273);
nor U12993 (N_12993,N_10582,N_9822);
nor U12994 (N_12994,N_9569,N_10925);
nand U12995 (N_12995,N_9355,N_10746);
or U12996 (N_12996,N_9279,N_10475);
nand U12997 (N_12997,N_9342,N_10631);
nor U12998 (N_12998,N_11032,N_10496);
or U12999 (N_12999,N_11914,N_11666);
nor U13000 (N_13000,N_10734,N_11826);
or U13001 (N_13001,N_10137,N_10322);
nor U13002 (N_13002,N_11242,N_11814);
and U13003 (N_13003,N_10744,N_10417);
nand U13004 (N_13004,N_10277,N_9491);
or U13005 (N_13005,N_11153,N_10938);
nand U13006 (N_13006,N_10426,N_11078);
nor U13007 (N_13007,N_11532,N_9194);
nor U13008 (N_13008,N_9161,N_10006);
nand U13009 (N_13009,N_9946,N_10776);
nand U13010 (N_13010,N_9689,N_11293);
and U13011 (N_13011,N_11196,N_9390);
nand U13012 (N_13012,N_10144,N_11410);
nand U13013 (N_13013,N_10515,N_11113);
xnor U13014 (N_13014,N_10798,N_11229);
and U13015 (N_13015,N_9865,N_10658);
nand U13016 (N_13016,N_10903,N_11734);
nand U13017 (N_13017,N_11005,N_9631);
nor U13018 (N_13018,N_10389,N_9354);
nor U13019 (N_13019,N_10169,N_11358);
and U13020 (N_13020,N_10854,N_9192);
and U13021 (N_13021,N_10284,N_11106);
nand U13022 (N_13022,N_9039,N_11020);
and U13023 (N_13023,N_11940,N_9193);
or U13024 (N_13024,N_9027,N_11992);
and U13025 (N_13025,N_9304,N_9803);
and U13026 (N_13026,N_10637,N_11432);
nor U13027 (N_13027,N_11305,N_10444);
nand U13028 (N_13028,N_10412,N_10663);
or U13029 (N_13029,N_10000,N_9848);
nand U13030 (N_13030,N_11203,N_10286);
nand U13031 (N_13031,N_9696,N_9847);
nor U13032 (N_13032,N_11749,N_9439);
and U13033 (N_13033,N_9845,N_10055);
nor U13034 (N_13034,N_11426,N_9449);
nor U13035 (N_13035,N_10552,N_10062);
nor U13036 (N_13036,N_10082,N_9411);
and U13037 (N_13037,N_10573,N_11878);
and U13038 (N_13038,N_9489,N_11682);
and U13039 (N_13039,N_10867,N_10887);
nor U13040 (N_13040,N_11045,N_10338);
and U13041 (N_13041,N_10621,N_9772);
or U13042 (N_13042,N_11491,N_10850);
xor U13043 (N_13043,N_9579,N_9444);
or U13044 (N_13044,N_11762,N_10481);
nor U13045 (N_13045,N_11087,N_11079);
or U13046 (N_13046,N_11338,N_9476);
nand U13047 (N_13047,N_10207,N_9864);
or U13048 (N_13048,N_10528,N_10043);
nor U13049 (N_13049,N_10936,N_10242);
nand U13050 (N_13050,N_9374,N_9216);
nand U13051 (N_13051,N_9320,N_10118);
nand U13052 (N_13052,N_9207,N_11404);
and U13053 (N_13053,N_10693,N_9168);
nor U13054 (N_13054,N_10885,N_9905);
or U13055 (N_13055,N_11086,N_10450);
and U13056 (N_13056,N_9123,N_9233);
nand U13057 (N_13057,N_11545,N_10820);
or U13058 (N_13058,N_9726,N_9676);
nand U13059 (N_13059,N_11076,N_10328);
nand U13060 (N_13060,N_11671,N_10295);
and U13061 (N_13061,N_11071,N_10422);
nand U13062 (N_13062,N_9093,N_10565);
or U13063 (N_13063,N_10224,N_10732);
nor U13064 (N_13064,N_10011,N_9296);
nand U13065 (N_13065,N_11602,N_11199);
nand U13066 (N_13066,N_9009,N_10017);
and U13067 (N_13067,N_11736,N_9225);
or U13068 (N_13068,N_11813,N_9983);
and U13069 (N_13069,N_10321,N_11387);
or U13070 (N_13070,N_10914,N_10223);
or U13071 (N_13071,N_11627,N_10761);
nor U13072 (N_13072,N_9539,N_9560);
and U13073 (N_13073,N_10522,N_10814);
nor U13074 (N_13074,N_9156,N_9543);
nor U13075 (N_13075,N_10599,N_9895);
nand U13076 (N_13076,N_10071,N_10109);
nor U13077 (N_13077,N_9888,N_9919);
and U13078 (N_13078,N_9889,N_11315);
or U13079 (N_13079,N_10839,N_11892);
or U13080 (N_13080,N_10500,N_11710);
nand U13081 (N_13081,N_11717,N_10587);
or U13082 (N_13082,N_10250,N_9724);
nand U13083 (N_13083,N_11769,N_10692);
nor U13084 (N_13084,N_10955,N_10671);
nor U13085 (N_13085,N_11744,N_9677);
nand U13086 (N_13086,N_11619,N_11429);
or U13087 (N_13087,N_9943,N_9613);
or U13088 (N_13088,N_10911,N_9447);
nand U13089 (N_13089,N_9550,N_10667);
xnor U13090 (N_13090,N_11143,N_9367);
or U13091 (N_13091,N_10303,N_9958);
and U13092 (N_13092,N_9054,N_11222);
nor U13093 (N_13093,N_10384,N_9309);
and U13094 (N_13094,N_10705,N_11391);
nor U13095 (N_13095,N_10807,N_9685);
or U13096 (N_13096,N_10661,N_9357);
xor U13097 (N_13097,N_9450,N_11055);
nor U13098 (N_13098,N_11768,N_10980);
nand U13099 (N_13099,N_10291,N_9487);
nor U13100 (N_13100,N_9621,N_11704);
nand U13101 (N_13101,N_10035,N_10856);
and U13102 (N_13102,N_9057,N_9268);
or U13103 (N_13103,N_11236,N_11218);
and U13104 (N_13104,N_9474,N_10206);
or U13105 (N_13105,N_9704,N_11877);
nor U13106 (N_13106,N_11344,N_10827);
nand U13107 (N_13107,N_10857,N_10603);
or U13108 (N_13108,N_11611,N_10873);
nor U13109 (N_13109,N_10625,N_10714);
nor U13110 (N_13110,N_9601,N_9155);
nor U13111 (N_13111,N_10054,N_11800);
xnor U13112 (N_13112,N_11849,N_9862);
and U13113 (N_13113,N_10652,N_9087);
or U13114 (N_13114,N_11484,N_10998);
nand U13115 (N_13115,N_10581,N_11884);
nand U13116 (N_13116,N_11495,N_11044);
or U13117 (N_13117,N_10990,N_11486);
nand U13118 (N_13118,N_9402,N_10578);
or U13119 (N_13119,N_11471,N_11277);
and U13120 (N_13120,N_9799,N_10622);
or U13121 (N_13121,N_11995,N_10804);
or U13122 (N_13122,N_9883,N_9681);
or U13123 (N_13123,N_9956,N_10376);
nor U13124 (N_13124,N_10626,N_9664);
or U13125 (N_13125,N_11108,N_11784);
nand U13126 (N_13126,N_9964,N_11513);
and U13127 (N_13127,N_11311,N_11362);
and U13128 (N_13128,N_11490,N_10653);
or U13129 (N_13129,N_10456,N_10132);
nand U13130 (N_13130,N_11952,N_11538);
nand U13131 (N_13131,N_10758,N_9351);
xor U13132 (N_13132,N_10189,N_9068);
and U13133 (N_13133,N_11219,N_9720);
and U13134 (N_13134,N_10486,N_11740);
or U13135 (N_13135,N_10513,N_10057);
nor U13136 (N_13136,N_9498,N_9328);
or U13137 (N_13137,N_11309,N_10566);
or U13138 (N_13138,N_9043,N_10419);
xor U13139 (N_13139,N_9749,N_11712);
nor U13140 (N_13140,N_11845,N_10666);
and U13141 (N_13141,N_9502,N_9051);
and U13142 (N_13142,N_11476,N_11373);
or U13143 (N_13143,N_11382,N_9022);
nand U13144 (N_13144,N_10868,N_9408);
nor U13145 (N_13145,N_10151,N_9317);
nor U13146 (N_13146,N_11056,N_10394);
and U13147 (N_13147,N_10305,N_10851);
or U13148 (N_13148,N_11875,N_11904);
nand U13149 (N_13149,N_10630,N_9839);
and U13150 (N_13150,N_9315,N_10289);
nand U13151 (N_13151,N_9371,N_9744);
or U13152 (N_13152,N_10845,N_9985);
nand U13153 (N_13153,N_9293,N_9338);
or U13154 (N_13154,N_11492,N_11371);
or U13155 (N_13155,N_10458,N_10346);
or U13156 (N_13156,N_11861,N_11618);
or U13157 (N_13157,N_11617,N_10737);
and U13158 (N_13158,N_10976,N_11328);
nor U13159 (N_13159,N_10864,N_10254);
nor U13160 (N_13160,N_10904,N_11489);
nor U13161 (N_13161,N_9636,N_10570);
or U13162 (N_13162,N_11938,N_9660);
nor U13163 (N_13163,N_11595,N_10001);
nand U13164 (N_13164,N_11415,N_9125);
nor U13165 (N_13165,N_11687,N_11852);
nor U13166 (N_13166,N_10264,N_9275);
and U13167 (N_13167,N_10261,N_10411);
or U13168 (N_13168,N_10473,N_11957);
nand U13169 (N_13169,N_11681,N_10502);
nand U13170 (N_13170,N_11259,N_10945);
nor U13171 (N_13171,N_11728,N_9659);
nor U13172 (N_13172,N_9871,N_10595);
nor U13173 (N_13173,N_9255,N_11473);
nand U13174 (N_13174,N_9873,N_11599);
or U13175 (N_13175,N_9297,N_11847);
xor U13176 (N_13176,N_10689,N_10583);
nor U13177 (N_13177,N_9537,N_11588);
and U13178 (N_13178,N_10510,N_11840);
and U13179 (N_13179,N_11061,N_11690);
nor U13180 (N_13180,N_9222,N_11424);
nand U13181 (N_13181,N_11732,N_9174);
nor U13182 (N_13182,N_9902,N_9461);
nor U13183 (N_13183,N_11761,N_11073);
and U13184 (N_13184,N_11052,N_11735);
and U13185 (N_13185,N_11386,N_11273);
or U13186 (N_13186,N_10823,N_9816);
and U13187 (N_13187,N_10788,N_11657);
or U13188 (N_13188,N_9107,N_9823);
or U13189 (N_13189,N_11824,N_9570);
or U13190 (N_13190,N_9494,N_11478);
nor U13191 (N_13191,N_10756,N_9323);
nand U13192 (N_13192,N_9838,N_11531);
nand U13193 (N_13193,N_9531,N_11303);
and U13194 (N_13194,N_9128,N_9254);
nand U13195 (N_13195,N_9377,N_9145);
nand U13196 (N_13196,N_11238,N_9096);
and U13197 (N_13197,N_10956,N_10782);
or U13198 (N_13198,N_11724,N_10405);
and U13199 (N_13199,N_10832,N_11331);
nand U13200 (N_13200,N_9261,N_11685);
nor U13201 (N_13201,N_9206,N_11274);
or U13202 (N_13202,N_11629,N_11193);
nand U13203 (N_13203,N_11871,N_11580);
or U13204 (N_13204,N_11979,N_11929);
nand U13205 (N_13205,N_9262,N_10691);
xor U13206 (N_13206,N_10283,N_9701);
nor U13207 (N_13207,N_11948,N_9467);
and U13208 (N_13208,N_11042,N_10034);
nor U13209 (N_13209,N_9718,N_11615);
or U13210 (N_13210,N_10416,N_10225);
or U13211 (N_13211,N_10112,N_9005);
or U13212 (N_13212,N_11544,N_10018);
and U13213 (N_13213,N_10061,N_10575);
nor U13214 (N_13214,N_11253,N_11632);
and U13215 (N_13215,N_11860,N_10041);
or U13216 (N_13216,N_10536,N_10890);
xnor U13217 (N_13217,N_10965,N_11390);
or U13218 (N_13218,N_9189,N_11485);
and U13219 (N_13219,N_11009,N_10742);
nor U13220 (N_13220,N_9552,N_11172);
or U13221 (N_13221,N_10946,N_10800);
nand U13222 (N_13222,N_9557,N_10390);
or U13223 (N_13223,N_11119,N_9431);
and U13224 (N_13224,N_10549,N_10117);
nand U13225 (N_13225,N_10038,N_10433);
nor U13226 (N_13226,N_10350,N_10430);
nand U13227 (N_13227,N_11396,N_10066);
and U13228 (N_13228,N_10388,N_11053);
nor U13229 (N_13229,N_11752,N_11653);
and U13230 (N_13230,N_10542,N_9435);
and U13231 (N_13231,N_9289,N_11421);
nand U13232 (N_13232,N_10585,N_9801);
or U13233 (N_13233,N_11684,N_11916);
or U13234 (N_13234,N_11093,N_11807);
or U13235 (N_13235,N_9224,N_10337);
and U13236 (N_13236,N_11745,N_10231);
nand U13237 (N_13237,N_11209,N_9538);
nor U13238 (N_13238,N_9908,N_11123);
nand U13239 (N_13239,N_11033,N_9372);
nand U13240 (N_13240,N_9695,N_9759);
and U13241 (N_13241,N_11182,N_11008);
and U13242 (N_13242,N_9395,N_10048);
nor U13243 (N_13243,N_10184,N_9699);
nand U13244 (N_13244,N_10930,N_11099);
nand U13245 (N_13245,N_9565,N_9265);
and U13246 (N_13246,N_11225,N_10425);
nand U13247 (N_13247,N_10819,N_10203);
nand U13248 (N_13248,N_11781,N_11224);
nand U13249 (N_13249,N_11586,N_10127);
and U13250 (N_13250,N_10960,N_11026);
nor U13251 (N_13251,N_9912,N_9020);
nor U13252 (N_13252,N_9775,N_11568);
or U13253 (N_13253,N_9814,N_10766);
or U13254 (N_13254,N_9483,N_11162);
or U13255 (N_13255,N_10010,N_10796);
and U13256 (N_13256,N_11521,N_9366);
nor U13257 (N_13257,N_9480,N_9140);
and U13258 (N_13258,N_11272,N_11742);
nor U13259 (N_13259,N_11226,N_9324);
nand U13260 (N_13260,N_10952,N_9329);
and U13261 (N_13261,N_10736,N_11620);
nor U13262 (N_13262,N_11363,N_9669);
nor U13263 (N_13263,N_10380,N_11567);
nand U13264 (N_13264,N_10162,N_11466);
nor U13265 (N_13265,N_9620,N_10727);
and U13266 (N_13266,N_9730,N_11858);
and U13267 (N_13267,N_9808,N_10095);
nor U13268 (N_13268,N_11208,N_10448);
or U13269 (N_13269,N_10228,N_9960);
nand U13270 (N_13270,N_10889,N_9827);
nor U13271 (N_13271,N_9180,N_9709);
nand U13272 (N_13272,N_11994,N_10190);
nand U13273 (N_13273,N_11986,N_10408);
and U13274 (N_13274,N_9308,N_9031);
or U13275 (N_13275,N_11114,N_10272);
or U13276 (N_13276,N_9609,N_9614);
nor U13277 (N_13277,N_9291,N_9765);
nand U13278 (N_13278,N_11081,N_9714);
and U13279 (N_13279,N_11400,N_10559);
or U13280 (N_13280,N_9610,N_10681);
nand U13281 (N_13281,N_11354,N_9877);
or U13282 (N_13282,N_9737,N_10222);
nor U13283 (N_13283,N_10739,N_9859);
nand U13284 (N_13284,N_11268,N_11335);
xnor U13285 (N_13285,N_10410,N_9058);
and U13286 (N_13286,N_9240,N_10366);
nand U13287 (N_13287,N_11482,N_9294);
or U13288 (N_13288,N_9825,N_11414);
or U13289 (N_13289,N_11794,N_9141);
and U13290 (N_13290,N_11573,N_9266);
nor U13291 (N_13291,N_9535,N_9026);
or U13292 (N_13292,N_10345,N_9843);
nor U13293 (N_13293,N_11969,N_11276);
or U13294 (N_13294,N_9841,N_11951);
and U13295 (N_13295,N_10538,N_9630);
nor U13296 (N_13296,N_11648,N_10199);
and U13297 (N_13297,N_10124,N_9106);
and U13298 (N_13298,N_10483,N_10047);
nand U13299 (N_13299,N_10221,N_10040);
or U13300 (N_13300,N_11974,N_11175);
and U13301 (N_13301,N_9691,N_10594);
or U13302 (N_13302,N_10750,N_9285);
or U13303 (N_13303,N_10523,N_11941);
or U13304 (N_13304,N_9343,N_10431);
nand U13305 (N_13305,N_10443,N_11307);
or U13306 (N_13306,N_11083,N_9049);
nor U13307 (N_13307,N_11923,N_10075);
xor U13308 (N_13308,N_9886,N_10747);
nand U13309 (N_13309,N_9619,N_9311);
and U13310 (N_13310,N_9581,N_9437);
nor U13311 (N_13311,N_9386,N_11541);
and U13312 (N_13312,N_9111,N_9178);
nor U13313 (N_13313,N_11643,N_11655);
or U13314 (N_13314,N_10092,N_11832);
xnor U13315 (N_13315,N_9947,N_11958);
nand U13316 (N_13316,N_10099,N_9572);
nor U13317 (N_13317,N_9362,N_11879);
and U13318 (N_13318,N_9915,N_11267);
or U13319 (N_13319,N_10593,N_11144);
nand U13320 (N_13320,N_9047,N_11634);
and U13321 (N_13321,N_9594,N_9855);
nand U13322 (N_13322,N_9934,N_11804);
nor U13323 (N_13323,N_10537,N_10163);
or U13324 (N_13324,N_10257,N_10841);
or U13325 (N_13325,N_10131,N_10741);
or U13326 (N_13326,N_10317,N_9244);
or U13327 (N_13327,N_11778,N_9248);
xor U13328 (N_13328,N_11829,N_11630);
and U13329 (N_13329,N_11758,N_9741);
or U13330 (N_13330,N_11237,N_9831);
and U13331 (N_13331,N_10480,N_9706);
and U13332 (N_13332,N_9163,N_11152);
or U13333 (N_13333,N_10251,N_10994);
and U13334 (N_13334,N_10363,N_11418);
nand U13335 (N_13335,N_10717,N_9056);
and U13336 (N_13336,N_10166,N_11120);
nor U13337 (N_13337,N_11809,N_9625);
nor U13338 (N_13338,N_11326,N_9590);
or U13339 (N_13339,N_11502,N_11956);
nand U13340 (N_13340,N_10898,N_9599);
or U13341 (N_13341,N_9869,N_9988);
or U13342 (N_13342,N_10763,N_9492);
or U13343 (N_13343,N_9643,N_9642);
nor U13344 (N_13344,N_9924,N_9936);
nand U13345 (N_13345,N_9829,N_10869);
or U13346 (N_13346,N_10183,N_11626);
nor U13347 (N_13347,N_9894,N_10933);
nand U13348 (N_13348,N_10122,N_10460);
nor U13349 (N_13349,N_9748,N_10613);
nor U13350 (N_13350,N_10309,N_9237);
xor U13351 (N_13351,N_9713,N_9242);
and U13352 (N_13352,N_9771,N_10386);
nor U13353 (N_13353,N_10912,N_10817);
nor U13354 (N_13354,N_9596,N_11971);
and U13355 (N_13355,N_10900,N_10698);
or U13356 (N_13356,N_10104,N_10627);
or U13357 (N_13357,N_11281,N_11679);
xnor U13358 (N_13358,N_10982,N_9287);
and U13359 (N_13359,N_9221,N_11022);
and U13360 (N_13360,N_9239,N_10891);
nand U13361 (N_13361,N_11912,N_10672);
and U13362 (N_13362,N_9303,N_11221);
nor U13363 (N_13363,N_10294,N_9336);
and U13364 (N_13364,N_11190,N_11069);
or U13365 (N_13365,N_11659,N_9012);
or U13366 (N_13366,N_11843,N_11515);
or U13367 (N_13367,N_10232,N_11158);
or U13368 (N_13368,N_10606,N_10247);
or U13369 (N_13369,N_11968,N_9721);
nand U13370 (N_13370,N_10567,N_11173);
and U13371 (N_13371,N_10710,N_10482);
nor U13372 (N_13372,N_10140,N_11258);
or U13373 (N_13373,N_9719,N_11610);
nand U13374 (N_13374,N_9019,N_11030);
nor U13375 (N_13375,N_9345,N_11262);
nor U13376 (N_13376,N_10269,N_9365);
and U13377 (N_13377,N_10126,N_9974);
nor U13378 (N_13378,N_10808,N_10446);
or U13379 (N_13379,N_10493,N_10014);
nand U13380 (N_13380,N_11316,N_9084);
nor U13381 (N_13381,N_9334,N_9510);
nand U13382 (N_13382,N_11180,N_10920);
xor U13383 (N_13383,N_10488,N_11092);
nand U13384 (N_13384,N_10026,N_9481);
and U13385 (N_13385,N_11678,N_11911);
nor U13386 (N_13386,N_11191,N_10432);
and U13387 (N_13387,N_9363,N_10723);
nand U13388 (N_13388,N_10491,N_10833);
or U13389 (N_13389,N_11290,N_10724);
nor U13390 (N_13390,N_11097,N_10107);
and U13391 (N_13391,N_10551,N_10797);
nor U13392 (N_13392,N_10684,N_11142);
nor U13393 (N_13393,N_9593,N_9075);
or U13394 (N_13394,N_11457,N_11529);
nand U13395 (N_13395,N_9608,N_11510);
or U13396 (N_13396,N_10230,N_11727);
xor U13397 (N_13397,N_10932,N_10555);
nand U13398 (N_13398,N_11723,N_9112);
xor U13399 (N_13399,N_9970,N_9900);
nor U13400 (N_13400,N_11528,N_10351);
or U13401 (N_13401,N_9962,N_9738);
nor U13402 (N_13402,N_9082,N_11207);
nand U13403 (N_13403,N_11462,N_11917);
nand U13404 (N_13404,N_11597,N_11625);
or U13405 (N_13405,N_11137,N_10569);
nand U13406 (N_13406,N_9017,N_9127);
and U13407 (N_13407,N_11913,N_9036);
xnor U13408 (N_13408,N_9835,N_11289);
or U13409 (N_13409,N_11393,N_10520);
nor U13410 (N_13410,N_9337,N_10777);
nor U13411 (N_13411,N_11553,N_11448);
nor U13412 (N_13412,N_11961,N_11981);
nand U13413 (N_13413,N_9872,N_10597);
nor U13414 (N_13414,N_10821,N_9732);
and U13415 (N_13415,N_11444,N_10138);
nand U13416 (N_13416,N_10359,N_10178);
nand U13417 (N_13417,N_9238,N_9723);
and U13418 (N_13418,N_10415,N_10524);
nor U13419 (N_13419,N_9076,N_11043);
xor U13420 (N_13420,N_9421,N_11782);
or U13421 (N_13421,N_11909,N_11987);
xor U13422 (N_13422,N_9786,N_9792);
nand U13423 (N_13423,N_9496,N_9256);
nand U13424 (N_13424,N_11950,N_10905);
or U13425 (N_13425,N_9671,N_11799);
nand U13426 (N_13426,N_10702,N_10560);
or U13427 (N_13427,N_10601,N_10361);
and U13428 (N_13428,N_10881,N_9406);
and U13429 (N_13429,N_10708,N_10356);
or U13430 (N_13430,N_9313,N_10327);
and U13431 (N_13431,N_10064,N_10326);
nand U13432 (N_13432,N_10550,N_11308);
or U13433 (N_13433,N_10919,N_9430);
and U13434 (N_13434,N_10941,N_9050);
nand U13435 (N_13435,N_10044,N_9927);
and U13436 (N_13436,N_11702,N_11058);
and U13437 (N_13437,N_10439,N_9490);
or U13438 (N_13438,N_9065,N_9091);
or U13439 (N_13439,N_11984,N_9158);
or U13440 (N_13440,N_9441,N_9152);
or U13441 (N_13441,N_11351,N_9680);
nor U13442 (N_13442,N_11082,N_10983);
and U13443 (N_13443,N_9055,N_11314);
and U13444 (N_13444,N_10342,N_11469);
nand U13445 (N_13445,N_9414,N_9485);
xor U13446 (N_13446,N_11068,N_9832);
nor U13447 (N_13447,N_10704,N_9059);
nand U13448 (N_13448,N_10688,N_9359);
or U13449 (N_13449,N_10752,N_9782);
nor U13450 (N_13450,N_9644,N_10686);
nand U13451 (N_13451,N_9692,N_11100);
nor U13452 (N_13452,N_10564,N_9305);
nand U13453 (N_13453,N_9656,N_9410);
and U13454 (N_13454,N_9177,N_11235);
or U13455 (N_13455,N_10022,N_9722);
and U13456 (N_13456,N_11645,N_11930);
xor U13457 (N_13457,N_10694,N_9484);
nor U13458 (N_13458,N_11543,N_11239);
or U13459 (N_13459,N_10367,N_11696);
or U13460 (N_13460,N_9836,N_9232);
nor U13461 (N_13461,N_10963,N_9062);
or U13462 (N_13462,N_10592,N_9064);
nor U13463 (N_13463,N_11280,N_11037);
nand U13464 (N_13464,N_10632,N_9175);
nand U13465 (N_13465,N_10610,N_9269);
or U13466 (N_13466,N_11063,N_10354);
xor U13467 (N_13467,N_10438,N_9705);
or U13468 (N_13468,N_9944,N_10690);
nor U13469 (N_13469,N_10028,N_10453);
or U13470 (N_13470,N_11406,N_10650);
nor U13471 (N_13471,N_10115,N_9534);
or U13472 (N_13472,N_10375,N_11733);
or U13473 (N_13473,N_11996,N_9913);
nand U13474 (N_13474,N_11668,N_10877);
nand U13475 (N_13475,N_11656,N_9563);
and U13476 (N_13476,N_9818,N_10200);
and U13477 (N_13477,N_10293,N_9984);
nor U13478 (N_13478,N_9400,N_10042);
nor U13479 (N_13479,N_9445,N_10810);
and U13480 (N_13480,N_11003,N_9559);
xor U13481 (N_13481,N_9167,N_10662);
nand U13482 (N_13482,N_9592,N_11720);
nand U13483 (N_13483,N_9751,N_11993);
nor U13484 (N_13484,N_10086,N_9968);
and U13485 (N_13485,N_10244,N_11572);
and U13486 (N_13486,N_10219,N_9138);
and U13487 (N_13487,N_9132,N_10319);
and U13488 (N_13488,N_11139,N_10525);
nor U13489 (N_13489,N_11874,N_11430);
or U13490 (N_13490,N_11747,N_11000);
nand U13491 (N_13491,N_9048,N_11966);
or U13492 (N_13492,N_11170,N_11683);
nand U13493 (N_13493,N_11194,N_9460);
nor U13494 (N_13494,N_10352,N_10179);
and U13495 (N_13495,N_11167,N_9903);
nand U13496 (N_13496,N_11692,N_10656);
nor U13497 (N_13497,N_11856,N_10029);
nor U13498 (N_13498,N_11357,N_11888);
nand U13499 (N_13499,N_11883,N_9171);
nor U13500 (N_13500,N_11490,N_11602);
and U13501 (N_13501,N_10498,N_11060);
nand U13502 (N_13502,N_11090,N_11463);
or U13503 (N_13503,N_10233,N_10051);
and U13504 (N_13504,N_10023,N_10141);
and U13505 (N_13505,N_10225,N_11642);
or U13506 (N_13506,N_11840,N_9327);
nand U13507 (N_13507,N_9397,N_9288);
nor U13508 (N_13508,N_11030,N_10669);
or U13509 (N_13509,N_10201,N_11661);
nand U13510 (N_13510,N_11497,N_9273);
nor U13511 (N_13511,N_11131,N_9986);
or U13512 (N_13512,N_10271,N_9995);
or U13513 (N_13513,N_9935,N_10687);
or U13514 (N_13514,N_10115,N_10694);
or U13515 (N_13515,N_10511,N_11301);
and U13516 (N_13516,N_9050,N_10388);
and U13517 (N_13517,N_11837,N_10510);
nand U13518 (N_13518,N_10912,N_9020);
and U13519 (N_13519,N_9102,N_11132);
and U13520 (N_13520,N_10683,N_10756);
and U13521 (N_13521,N_9666,N_11206);
nor U13522 (N_13522,N_10998,N_10331);
nor U13523 (N_13523,N_9642,N_9593);
or U13524 (N_13524,N_11724,N_9603);
nand U13525 (N_13525,N_11326,N_9456);
and U13526 (N_13526,N_11919,N_11303);
xor U13527 (N_13527,N_10915,N_11471);
nor U13528 (N_13528,N_10831,N_9737);
nor U13529 (N_13529,N_11719,N_11380);
nand U13530 (N_13530,N_10210,N_10266);
and U13531 (N_13531,N_11868,N_9547);
nor U13532 (N_13532,N_11007,N_9334);
or U13533 (N_13533,N_10049,N_10919);
and U13534 (N_13534,N_9884,N_10736);
and U13535 (N_13535,N_10595,N_9270);
or U13536 (N_13536,N_10613,N_10916);
nand U13537 (N_13537,N_9469,N_10786);
nand U13538 (N_13538,N_10764,N_10039);
nor U13539 (N_13539,N_10735,N_11951);
nor U13540 (N_13540,N_11516,N_10310);
nor U13541 (N_13541,N_10214,N_10208);
nand U13542 (N_13542,N_11402,N_11937);
nand U13543 (N_13543,N_11304,N_9217);
and U13544 (N_13544,N_11974,N_11148);
nand U13545 (N_13545,N_11010,N_10293);
nor U13546 (N_13546,N_10792,N_10395);
or U13547 (N_13547,N_10062,N_9267);
and U13548 (N_13548,N_11729,N_9644);
or U13549 (N_13549,N_9613,N_11142);
nor U13550 (N_13550,N_11311,N_11579);
nor U13551 (N_13551,N_11566,N_9708);
nand U13552 (N_13552,N_11507,N_11862);
and U13553 (N_13553,N_9028,N_9713);
or U13554 (N_13554,N_9828,N_10642);
nand U13555 (N_13555,N_9908,N_10531);
and U13556 (N_13556,N_9679,N_10336);
nor U13557 (N_13557,N_10338,N_9031);
nand U13558 (N_13558,N_11310,N_9425);
or U13559 (N_13559,N_10029,N_11153);
nor U13560 (N_13560,N_9138,N_10201);
nand U13561 (N_13561,N_10843,N_9823);
nand U13562 (N_13562,N_11547,N_10258);
and U13563 (N_13563,N_10539,N_9201);
or U13564 (N_13564,N_10942,N_10227);
xnor U13565 (N_13565,N_9406,N_9054);
or U13566 (N_13566,N_10107,N_11943);
and U13567 (N_13567,N_10900,N_11679);
or U13568 (N_13568,N_10820,N_11685);
or U13569 (N_13569,N_10222,N_11243);
nand U13570 (N_13570,N_9558,N_10680);
or U13571 (N_13571,N_11924,N_9936);
nand U13572 (N_13572,N_10314,N_9704);
and U13573 (N_13573,N_10647,N_11214);
nor U13574 (N_13574,N_10046,N_9391);
or U13575 (N_13575,N_10918,N_11917);
nand U13576 (N_13576,N_9899,N_10216);
nor U13577 (N_13577,N_11839,N_10725);
xnor U13578 (N_13578,N_10782,N_9092);
nor U13579 (N_13579,N_11421,N_9065);
or U13580 (N_13580,N_10374,N_11259);
and U13581 (N_13581,N_11483,N_11450);
and U13582 (N_13582,N_11460,N_10250);
or U13583 (N_13583,N_9998,N_10398);
and U13584 (N_13584,N_11893,N_10289);
and U13585 (N_13585,N_10359,N_11468);
nor U13586 (N_13586,N_9374,N_9251);
nor U13587 (N_13587,N_10811,N_10128);
or U13588 (N_13588,N_10791,N_10064);
nor U13589 (N_13589,N_11205,N_11487);
or U13590 (N_13590,N_11911,N_11317);
nor U13591 (N_13591,N_10400,N_10568);
nor U13592 (N_13592,N_11674,N_9200);
nor U13593 (N_13593,N_9087,N_10599);
and U13594 (N_13594,N_10083,N_10351);
or U13595 (N_13595,N_9860,N_11988);
nor U13596 (N_13596,N_11473,N_11650);
and U13597 (N_13597,N_10948,N_9895);
nand U13598 (N_13598,N_10662,N_9776);
nand U13599 (N_13599,N_9539,N_11196);
nand U13600 (N_13600,N_11080,N_9591);
or U13601 (N_13601,N_9856,N_9397);
xor U13602 (N_13602,N_10698,N_10603);
and U13603 (N_13603,N_9407,N_9390);
and U13604 (N_13604,N_11688,N_9828);
nand U13605 (N_13605,N_11775,N_10471);
or U13606 (N_13606,N_11207,N_11552);
or U13607 (N_13607,N_10757,N_11706);
nand U13608 (N_13608,N_9390,N_11204);
or U13609 (N_13609,N_11426,N_11630);
nor U13610 (N_13610,N_9368,N_10970);
nor U13611 (N_13611,N_9754,N_10764);
or U13612 (N_13612,N_9788,N_9822);
nor U13613 (N_13613,N_9784,N_10213);
nand U13614 (N_13614,N_10281,N_9864);
or U13615 (N_13615,N_11842,N_10840);
or U13616 (N_13616,N_11794,N_11349);
nand U13617 (N_13617,N_10619,N_9781);
and U13618 (N_13618,N_11435,N_10617);
and U13619 (N_13619,N_9818,N_10603);
nor U13620 (N_13620,N_10155,N_11478);
and U13621 (N_13621,N_10510,N_11651);
and U13622 (N_13622,N_9526,N_10598);
or U13623 (N_13623,N_10916,N_9466);
and U13624 (N_13624,N_10950,N_11082);
and U13625 (N_13625,N_11101,N_10509);
or U13626 (N_13626,N_10625,N_10544);
nand U13627 (N_13627,N_11281,N_11480);
nor U13628 (N_13628,N_10128,N_9735);
and U13629 (N_13629,N_10262,N_10897);
or U13630 (N_13630,N_9046,N_9638);
or U13631 (N_13631,N_10994,N_9168);
or U13632 (N_13632,N_10139,N_10670);
nand U13633 (N_13633,N_11212,N_10573);
nand U13634 (N_13634,N_9339,N_9988);
nand U13635 (N_13635,N_11724,N_9153);
and U13636 (N_13636,N_9814,N_10576);
or U13637 (N_13637,N_11785,N_9949);
and U13638 (N_13638,N_10725,N_10311);
and U13639 (N_13639,N_9056,N_9670);
or U13640 (N_13640,N_9988,N_11818);
xnor U13641 (N_13641,N_10497,N_11510);
nand U13642 (N_13642,N_9586,N_9784);
nor U13643 (N_13643,N_10493,N_10207);
nor U13644 (N_13644,N_9674,N_9855);
or U13645 (N_13645,N_11291,N_11769);
nand U13646 (N_13646,N_9835,N_9609);
nor U13647 (N_13647,N_9278,N_10233);
and U13648 (N_13648,N_10412,N_9440);
and U13649 (N_13649,N_10997,N_11570);
nand U13650 (N_13650,N_10319,N_10334);
nand U13651 (N_13651,N_9364,N_11616);
nand U13652 (N_13652,N_11773,N_10142);
nand U13653 (N_13653,N_9961,N_11612);
or U13654 (N_13654,N_11407,N_11655);
and U13655 (N_13655,N_10688,N_11010);
nand U13656 (N_13656,N_10719,N_11705);
or U13657 (N_13657,N_10363,N_10632);
or U13658 (N_13658,N_9364,N_10652);
or U13659 (N_13659,N_10068,N_9255);
nand U13660 (N_13660,N_11816,N_9388);
nor U13661 (N_13661,N_9189,N_9086);
nand U13662 (N_13662,N_10543,N_9015);
nand U13663 (N_13663,N_10851,N_10380);
and U13664 (N_13664,N_11873,N_10964);
or U13665 (N_13665,N_11510,N_9958);
and U13666 (N_13666,N_11634,N_11580);
or U13667 (N_13667,N_9005,N_11585);
and U13668 (N_13668,N_9740,N_9201);
nor U13669 (N_13669,N_10662,N_9739);
or U13670 (N_13670,N_9306,N_11406);
and U13671 (N_13671,N_9579,N_10113);
and U13672 (N_13672,N_10231,N_10895);
or U13673 (N_13673,N_10811,N_10025);
nor U13674 (N_13674,N_11265,N_10560);
or U13675 (N_13675,N_10991,N_9274);
or U13676 (N_13676,N_10284,N_9732);
nand U13677 (N_13677,N_9111,N_10232);
or U13678 (N_13678,N_10805,N_10066);
xnor U13679 (N_13679,N_9231,N_10720);
nor U13680 (N_13680,N_9847,N_10456);
nor U13681 (N_13681,N_9054,N_10869);
nand U13682 (N_13682,N_10019,N_10543);
and U13683 (N_13683,N_11126,N_11960);
or U13684 (N_13684,N_10516,N_11052);
nand U13685 (N_13685,N_11196,N_11929);
or U13686 (N_13686,N_11950,N_11525);
nor U13687 (N_13687,N_9982,N_11215);
or U13688 (N_13688,N_11381,N_9571);
nand U13689 (N_13689,N_10179,N_11821);
nor U13690 (N_13690,N_9050,N_9464);
and U13691 (N_13691,N_9909,N_10646);
and U13692 (N_13692,N_9273,N_9922);
nand U13693 (N_13693,N_10866,N_10064);
and U13694 (N_13694,N_11880,N_11631);
and U13695 (N_13695,N_10162,N_10389);
nand U13696 (N_13696,N_10402,N_9970);
or U13697 (N_13697,N_9431,N_9938);
nand U13698 (N_13698,N_10768,N_11149);
nor U13699 (N_13699,N_10175,N_11325);
nand U13700 (N_13700,N_11707,N_9679);
or U13701 (N_13701,N_9758,N_10125);
nand U13702 (N_13702,N_11398,N_10617);
and U13703 (N_13703,N_9906,N_10754);
and U13704 (N_13704,N_10373,N_9043);
or U13705 (N_13705,N_9044,N_10362);
nand U13706 (N_13706,N_10686,N_9914);
nor U13707 (N_13707,N_10725,N_9992);
and U13708 (N_13708,N_9721,N_11429);
nand U13709 (N_13709,N_9120,N_10987);
or U13710 (N_13710,N_10098,N_9697);
and U13711 (N_13711,N_9661,N_9212);
nor U13712 (N_13712,N_10493,N_11494);
xnor U13713 (N_13713,N_9386,N_10535);
and U13714 (N_13714,N_9371,N_9938);
or U13715 (N_13715,N_10939,N_11388);
and U13716 (N_13716,N_11511,N_11235);
and U13717 (N_13717,N_11768,N_11088);
and U13718 (N_13718,N_9955,N_10928);
and U13719 (N_13719,N_9723,N_10233);
nand U13720 (N_13720,N_11036,N_10211);
nand U13721 (N_13721,N_10492,N_9323);
or U13722 (N_13722,N_10478,N_9068);
nand U13723 (N_13723,N_11854,N_9798);
and U13724 (N_13724,N_10397,N_11826);
nor U13725 (N_13725,N_9032,N_9718);
nor U13726 (N_13726,N_10254,N_9682);
or U13727 (N_13727,N_9777,N_10618);
and U13728 (N_13728,N_9262,N_9076);
and U13729 (N_13729,N_10392,N_10248);
and U13730 (N_13730,N_11122,N_9110);
nand U13731 (N_13731,N_9195,N_10014);
nand U13732 (N_13732,N_9919,N_10420);
nand U13733 (N_13733,N_11528,N_10711);
nand U13734 (N_13734,N_9860,N_11709);
and U13735 (N_13735,N_11276,N_11501);
nand U13736 (N_13736,N_10769,N_11464);
or U13737 (N_13737,N_10148,N_9332);
and U13738 (N_13738,N_10320,N_9094);
nand U13739 (N_13739,N_11264,N_11491);
and U13740 (N_13740,N_11808,N_10638);
and U13741 (N_13741,N_11965,N_11901);
nor U13742 (N_13742,N_10460,N_10945);
or U13743 (N_13743,N_9992,N_9097);
or U13744 (N_13744,N_10378,N_9911);
and U13745 (N_13745,N_11693,N_11569);
or U13746 (N_13746,N_10847,N_11474);
or U13747 (N_13747,N_9293,N_10965);
or U13748 (N_13748,N_9352,N_11294);
and U13749 (N_13749,N_11529,N_9882);
nand U13750 (N_13750,N_10924,N_9796);
or U13751 (N_13751,N_10191,N_11349);
nand U13752 (N_13752,N_10869,N_9935);
nand U13753 (N_13753,N_9839,N_10405);
nor U13754 (N_13754,N_10617,N_11447);
nand U13755 (N_13755,N_11206,N_11296);
nand U13756 (N_13756,N_10144,N_10183);
nand U13757 (N_13757,N_9083,N_11450);
nor U13758 (N_13758,N_11052,N_11910);
nor U13759 (N_13759,N_10405,N_9323);
nand U13760 (N_13760,N_11736,N_10771);
nor U13761 (N_13761,N_11116,N_9269);
nand U13762 (N_13762,N_10451,N_10741);
nor U13763 (N_13763,N_9874,N_10450);
nand U13764 (N_13764,N_9189,N_11646);
nor U13765 (N_13765,N_9175,N_11747);
nor U13766 (N_13766,N_11891,N_9307);
or U13767 (N_13767,N_10356,N_11910);
or U13768 (N_13768,N_11251,N_11819);
nor U13769 (N_13769,N_10531,N_9416);
nor U13770 (N_13770,N_10140,N_9966);
or U13771 (N_13771,N_9367,N_11641);
or U13772 (N_13772,N_10347,N_9888);
nor U13773 (N_13773,N_11971,N_9708);
nand U13774 (N_13774,N_11539,N_11182);
or U13775 (N_13775,N_11078,N_10469);
nor U13776 (N_13776,N_9204,N_9147);
nor U13777 (N_13777,N_9663,N_9119);
nand U13778 (N_13778,N_10003,N_11937);
or U13779 (N_13779,N_11589,N_11849);
nand U13780 (N_13780,N_9389,N_10566);
nor U13781 (N_13781,N_9861,N_10329);
nand U13782 (N_13782,N_10743,N_11628);
nor U13783 (N_13783,N_11218,N_10205);
or U13784 (N_13784,N_11460,N_11082);
nor U13785 (N_13785,N_9283,N_11807);
nor U13786 (N_13786,N_9364,N_11611);
or U13787 (N_13787,N_10092,N_9335);
nor U13788 (N_13788,N_9581,N_11094);
nand U13789 (N_13789,N_10178,N_10508);
or U13790 (N_13790,N_11226,N_10378);
nand U13791 (N_13791,N_9369,N_10833);
or U13792 (N_13792,N_11815,N_11877);
nor U13793 (N_13793,N_11331,N_9742);
and U13794 (N_13794,N_10054,N_11510);
and U13795 (N_13795,N_11217,N_9030);
nor U13796 (N_13796,N_10608,N_10941);
nor U13797 (N_13797,N_9093,N_11397);
xnor U13798 (N_13798,N_11209,N_11574);
and U13799 (N_13799,N_9024,N_11793);
nor U13800 (N_13800,N_10288,N_11313);
nor U13801 (N_13801,N_11560,N_10968);
nand U13802 (N_13802,N_10632,N_10164);
nor U13803 (N_13803,N_9090,N_11797);
nor U13804 (N_13804,N_10552,N_9475);
nand U13805 (N_13805,N_10921,N_9150);
or U13806 (N_13806,N_10750,N_11787);
and U13807 (N_13807,N_11773,N_9291);
or U13808 (N_13808,N_11126,N_11558);
and U13809 (N_13809,N_10417,N_9241);
nor U13810 (N_13810,N_11884,N_11351);
and U13811 (N_13811,N_9195,N_10431);
nand U13812 (N_13812,N_9218,N_10657);
nor U13813 (N_13813,N_11636,N_9099);
nor U13814 (N_13814,N_11778,N_10267);
nor U13815 (N_13815,N_9430,N_9436);
and U13816 (N_13816,N_11727,N_10555);
nor U13817 (N_13817,N_10124,N_10249);
nor U13818 (N_13818,N_9701,N_9959);
or U13819 (N_13819,N_10884,N_10150);
or U13820 (N_13820,N_11351,N_11955);
and U13821 (N_13821,N_9054,N_10086);
and U13822 (N_13822,N_10852,N_10857);
nand U13823 (N_13823,N_10424,N_10584);
nand U13824 (N_13824,N_10429,N_10789);
nand U13825 (N_13825,N_10020,N_11824);
nor U13826 (N_13826,N_9880,N_9360);
nand U13827 (N_13827,N_10796,N_11894);
nand U13828 (N_13828,N_9767,N_10413);
nand U13829 (N_13829,N_9518,N_10257);
or U13830 (N_13830,N_9572,N_10090);
or U13831 (N_13831,N_11056,N_10760);
and U13832 (N_13832,N_10409,N_11017);
nand U13833 (N_13833,N_9937,N_11757);
nand U13834 (N_13834,N_10793,N_11787);
nor U13835 (N_13835,N_11764,N_10166);
nand U13836 (N_13836,N_10581,N_10277);
nor U13837 (N_13837,N_11558,N_10000);
nor U13838 (N_13838,N_10766,N_10866);
and U13839 (N_13839,N_11239,N_9974);
or U13840 (N_13840,N_9030,N_10857);
or U13841 (N_13841,N_9103,N_9420);
and U13842 (N_13842,N_10745,N_9767);
or U13843 (N_13843,N_9561,N_10074);
nand U13844 (N_13844,N_10509,N_11517);
and U13845 (N_13845,N_9502,N_11890);
nand U13846 (N_13846,N_10650,N_9384);
or U13847 (N_13847,N_11646,N_10521);
and U13848 (N_13848,N_11286,N_10587);
or U13849 (N_13849,N_10966,N_10110);
nor U13850 (N_13850,N_9405,N_9714);
xnor U13851 (N_13851,N_11405,N_10378);
or U13852 (N_13852,N_10334,N_9301);
and U13853 (N_13853,N_11020,N_10301);
or U13854 (N_13854,N_10517,N_9319);
nand U13855 (N_13855,N_10660,N_9990);
xnor U13856 (N_13856,N_10643,N_9391);
and U13857 (N_13857,N_11898,N_9712);
nand U13858 (N_13858,N_10741,N_10649);
nor U13859 (N_13859,N_10908,N_11881);
or U13860 (N_13860,N_9918,N_11085);
and U13861 (N_13861,N_11660,N_11004);
or U13862 (N_13862,N_11183,N_11084);
nor U13863 (N_13863,N_10580,N_11695);
and U13864 (N_13864,N_9380,N_11904);
or U13865 (N_13865,N_11974,N_10735);
or U13866 (N_13866,N_11110,N_11864);
nor U13867 (N_13867,N_10161,N_11593);
nand U13868 (N_13868,N_9873,N_9626);
or U13869 (N_13869,N_9854,N_9858);
and U13870 (N_13870,N_9214,N_9849);
or U13871 (N_13871,N_9553,N_10909);
nor U13872 (N_13872,N_10902,N_9257);
nand U13873 (N_13873,N_10445,N_11305);
nand U13874 (N_13874,N_11335,N_9136);
or U13875 (N_13875,N_9474,N_11335);
and U13876 (N_13876,N_9951,N_11004);
nand U13877 (N_13877,N_10668,N_10735);
nor U13878 (N_13878,N_10368,N_10322);
and U13879 (N_13879,N_9400,N_9850);
nand U13880 (N_13880,N_9441,N_11464);
or U13881 (N_13881,N_10471,N_10387);
xor U13882 (N_13882,N_9460,N_9105);
nand U13883 (N_13883,N_9390,N_10834);
nand U13884 (N_13884,N_9422,N_11006);
nor U13885 (N_13885,N_10799,N_11848);
nor U13886 (N_13886,N_11105,N_10260);
nand U13887 (N_13887,N_9948,N_10970);
or U13888 (N_13888,N_9482,N_9288);
or U13889 (N_13889,N_9379,N_11216);
or U13890 (N_13890,N_11955,N_11620);
nor U13891 (N_13891,N_11380,N_11073);
or U13892 (N_13892,N_9451,N_10662);
nand U13893 (N_13893,N_9476,N_10299);
nor U13894 (N_13894,N_10601,N_10295);
and U13895 (N_13895,N_9483,N_10882);
and U13896 (N_13896,N_11853,N_11913);
nor U13897 (N_13897,N_10010,N_10453);
nand U13898 (N_13898,N_9169,N_10708);
nor U13899 (N_13899,N_11929,N_10895);
or U13900 (N_13900,N_9800,N_10836);
nor U13901 (N_13901,N_9159,N_9553);
or U13902 (N_13902,N_9783,N_9377);
nor U13903 (N_13903,N_9262,N_11441);
or U13904 (N_13904,N_9472,N_9021);
nand U13905 (N_13905,N_9102,N_11268);
or U13906 (N_13906,N_10918,N_11782);
nor U13907 (N_13907,N_10458,N_10357);
and U13908 (N_13908,N_10645,N_9517);
and U13909 (N_13909,N_9589,N_10027);
and U13910 (N_13910,N_11826,N_11183);
nor U13911 (N_13911,N_9376,N_10399);
or U13912 (N_13912,N_11479,N_9265);
nor U13913 (N_13913,N_10689,N_10075);
nor U13914 (N_13914,N_10314,N_11044);
or U13915 (N_13915,N_11219,N_10653);
nor U13916 (N_13916,N_10258,N_11142);
nor U13917 (N_13917,N_9590,N_11631);
and U13918 (N_13918,N_9047,N_11545);
or U13919 (N_13919,N_9723,N_11349);
nand U13920 (N_13920,N_11783,N_11476);
and U13921 (N_13921,N_11971,N_9278);
nand U13922 (N_13922,N_10582,N_10359);
xor U13923 (N_13923,N_11556,N_9365);
or U13924 (N_13924,N_11523,N_9222);
nor U13925 (N_13925,N_11138,N_11017);
or U13926 (N_13926,N_10894,N_10352);
and U13927 (N_13927,N_10847,N_11154);
nand U13928 (N_13928,N_11806,N_9440);
and U13929 (N_13929,N_9722,N_11756);
or U13930 (N_13930,N_9013,N_10048);
or U13931 (N_13931,N_11007,N_10618);
nand U13932 (N_13932,N_11481,N_9177);
nor U13933 (N_13933,N_9479,N_11536);
nand U13934 (N_13934,N_9395,N_10308);
nor U13935 (N_13935,N_11456,N_10314);
and U13936 (N_13936,N_10067,N_9543);
or U13937 (N_13937,N_10981,N_10046);
or U13938 (N_13938,N_11631,N_11688);
nand U13939 (N_13939,N_9393,N_11667);
and U13940 (N_13940,N_11197,N_10179);
xnor U13941 (N_13941,N_10820,N_10169);
or U13942 (N_13942,N_9090,N_9065);
and U13943 (N_13943,N_11300,N_9820);
nand U13944 (N_13944,N_10498,N_11380);
and U13945 (N_13945,N_11447,N_10889);
nand U13946 (N_13946,N_10194,N_11922);
nand U13947 (N_13947,N_10164,N_11324);
or U13948 (N_13948,N_10707,N_11533);
nand U13949 (N_13949,N_10451,N_11907);
or U13950 (N_13950,N_11368,N_9463);
nor U13951 (N_13951,N_10285,N_11280);
or U13952 (N_13952,N_10506,N_10306);
nor U13953 (N_13953,N_9822,N_11585);
and U13954 (N_13954,N_10606,N_9412);
or U13955 (N_13955,N_10911,N_10400);
or U13956 (N_13956,N_11349,N_11985);
or U13957 (N_13957,N_10014,N_9555);
or U13958 (N_13958,N_11910,N_10953);
nand U13959 (N_13959,N_9405,N_11064);
or U13960 (N_13960,N_10921,N_9887);
nor U13961 (N_13961,N_11566,N_11594);
or U13962 (N_13962,N_11607,N_11076);
nor U13963 (N_13963,N_10609,N_10302);
nand U13964 (N_13964,N_11806,N_10041);
or U13965 (N_13965,N_11951,N_9663);
and U13966 (N_13966,N_11799,N_10497);
nor U13967 (N_13967,N_10482,N_9614);
nand U13968 (N_13968,N_9506,N_9228);
and U13969 (N_13969,N_11749,N_9513);
nand U13970 (N_13970,N_9846,N_9067);
nor U13971 (N_13971,N_9743,N_9695);
or U13972 (N_13972,N_11820,N_11423);
nand U13973 (N_13973,N_11110,N_11077);
nor U13974 (N_13974,N_11702,N_11039);
nand U13975 (N_13975,N_11006,N_9345);
nand U13976 (N_13976,N_9281,N_9794);
or U13977 (N_13977,N_10556,N_9551);
nand U13978 (N_13978,N_11318,N_10866);
xnor U13979 (N_13979,N_11229,N_9160);
and U13980 (N_13980,N_11667,N_10148);
nand U13981 (N_13981,N_9567,N_11691);
or U13982 (N_13982,N_11332,N_11314);
nor U13983 (N_13983,N_10864,N_10515);
nor U13984 (N_13984,N_11264,N_9673);
or U13985 (N_13985,N_11648,N_10759);
nor U13986 (N_13986,N_10870,N_10469);
and U13987 (N_13987,N_10240,N_11317);
nor U13988 (N_13988,N_9130,N_10650);
nor U13989 (N_13989,N_9772,N_9619);
and U13990 (N_13990,N_9213,N_11190);
nor U13991 (N_13991,N_9233,N_9537);
nand U13992 (N_13992,N_11399,N_9839);
nor U13993 (N_13993,N_11069,N_11315);
nor U13994 (N_13994,N_9955,N_9381);
or U13995 (N_13995,N_9818,N_11873);
and U13996 (N_13996,N_10328,N_9695);
nand U13997 (N_13997,N_9929,N_9983);
nand U13998 (N_13998,N_11033,N_9117);
nand U13999 (N_13999,N_10698,N_11605);
nand U14000 (N_14000,N_11154,N_10074);
nand U14001 (N_14001,N_11146,N_9317);
nand U14002 (N_14002,N_11919,N_11669);
or U14003 (N_14003,N_9837,N_10732);
nor U14004 (N_14004,N_11977,N_11652);
nor U14005 (N_14005,N_11585,N_10624);
and U14006 (N_14006,N_11232,N_9660);
or U14007 (N_14007,N_10257,N_10948);
and U14008 (N_14008,N_11417,N_11759);
nand U14009 (N_14009,N_9506,N_9347);
nor U14010 (N_14010,N_10824,N_9803);
nand U14011 (N_14011,N_9762,N_10817);
nand U14012 (N_14012,N_9656,N_9485);
nor U14013 (N_14013,N_10757,N_10914);
nor U14014 (N_14014,N_9436,N_11556);
nor U14015 (N_14015,N_11553,N_10919);
nand U14016 (N_14016,N_9687,N_11603);
and U14017 (N_14017,N_11841,N_11162);
and U14018 (N_14018,N_10635,N_11200);
or U14019 (N_14019,N_10667,N_11624);
and U14020 (N_14020,N_11140,N_11690);
nand U14021 (N_14021,N_9710,N_10122);
or U14022 (N_14022,N_9856,N_9847);
or U14023 (N_14023,N_10339,N_10930);
nor U14024 (N_14024,N_10358,N_11092);
or U14025 (N_14025,N_9177,N_10196);
or U14026 (N_14026,N_11948,N_10838);
nand U14027 (N_14027,N_11746,N_11429);
and U14028 (N_14028,N_9575,N_11469);
nor U14029 (N_14029,N_9702,N_9545);
and U14030 (N_14030,N_9250,N_9728);
nand U14031 (N_14031,N_11566,N_11006);
or U14032 (N_14032,N_11214,N_11863);
xnor U14033 (N_14033,N_10508,N_11319);
nor U14034 (N_14034,N_9431,N_10276);
or U14035 (N_14035,N_10393,N_10812);
or U14036 (N_14036,N_11291,N_11444);
nor U14037 (N_14037,N_9335,N_9614);
nor U14038 (N_14038,N_9859,N_9250);
or U14039 (N_14039,N_10927,N_10069);
and U14040 (N_14040,N_10662,N_9597);
or U14041 (N_14041,N_10070,N_11285);
nand U14042 (N_14042,N_10466,N_9573);
and U14043 (N_14043,N_9360,N_11436);
nand U14044 (N_14044,N_9127,N_9240);
nand U14045 (N_14045,N_11180,N_10524);
or U14046 (N_14046,N_9768,N_10888);
and U14047 (N_14047,N_9253,N_10764);
or U14048 (N_14048,N_9567,N_9183);
nand U14049 (N_14049,N_11705,N_10572);
and U14050 (N_14050,N_10277,N_9627);
nor U14051 (N_14051,N_11264,N_9780);
nand U14052 (N_14052,N_11271,N_10469);
nand U14053 (N_14053,N_11993,N_9584);
or U14054 (N_14054,N_9463,N_10139);
nor U14055 (N_14055,N_9218,N_11695);
or U14056 (N_14056,N_9853,N_9696);
nand U14057 (N_14057,N_11352,N_10042);
and U14058 (N_14058,N_9384,N_11830);
nor U14059 (N_14059,N_11512,N_10233);
and U14060 (N_14060,N_10446,N_11310);
nand U14061 (N_14061,N_9962,N_9121);
nand U14062 (N_14062,N_10025,N_9155);
and U14063 (N_14063,N_9379,N_10284);
or U14064 (N_14064,N_10683,N_10672);
or U14065 (N_14065,N_10871,N_11138);
nand U14066 (N_14066,N_11697,N_11483);
nand U14067 (N_14067,N_10041,N_9447);
nor U14068 (N_14068,N_10252,N_9668);
nand U14069 (N_14069,N_10359,N_11381);
and U14070 (N_14070,N_9492,N_9673);
or U14071 (N_14071,N_9137,N_11788);
or U14072 (N_14072,N_11236,N_11927);
or U14073 (N_14073,N_10414,N_9625);
and U14074 (N_14074,N_9697,N_10435);
xnor U14075 (N_14075,N_10468,N_10710);
or U14076 (N_14076,N_10243,N_10344);
nor U14077 (N_14077,N_11555,N_10017);
and U14078 (N_14078,N_10391,N_9719);
and U14079 (N_14079,N_11410,N_9145);
or U14080 (N_14080,N_9921,N_9704);
xnor U14081 (N_14081,N_11626,N_10597);
and U14082 (N_14082,N_10780,N_9714);
or U14083 (N_14083,N_10619,N_11627);
nand U14084 (N_14084,N_11489,N_10243);
and U14085 (N_14085,N_9736,N_11591);
nand U14086 (N_14086,N_11462,N_9198);
nand U14087 (N_14087,N_10956,N_10259);
and U14088 (N_14088,N_9371,N_11706);
nor U14089 (N_14089,N_10523,N_9726);
and U14090 (N_14090,N_10405,N_10595);
and U14091 (N_14091,N_11462,N_10119);
or U14092 (N_14092,N_11250,N_11474);
nand U14093 (N_14093,N_9907,N_11880);
and U14094 (N_14094,N_10956,N_9116);
and U14095 (N_14095,N_9021,N_10818);
or U14096 (N_14096,N_11143,N_10401);
nor U14097 (N_14097,N_10717,N_10384);
nand U14098 (N_14098,N_10607,N_10154);
and U14099 (N_14099,N_10668,N_10958);
or U14100 (N_14100,N_9930,N_10432);
or U14101 (N_14101,N_10927,N_10239);
or U14102 (N_14102,N_10952,N_10640);
nand U14103 (N_14103,N_9109,N_9881);
xnor U14104 (N_14104,N_9938,N_10025);
nand U14105 (N_14105,N_10919,N_10797);
nand U14106 (N_14106,N_10309,N_11636);
nor U14107 (N_14107,N_11790,N_10833);
nand U14108 (N_14108,N_9549,N_10934);
or U14109 (N_14109,N_10600,N_11469);
or U14110 (N_14110,N_10147,N_11320);
nor U14111 (N_14111,N_10811,N_10660);
xnor U14112 (N_14112,N_11030,N_9373);
or U14113 (N_14113,N_11013,N_11948);
and U14114 (N_14114,N_11018,N_9008);
or U14115 (N_14115,N_10111,N_9629);
nor U14116 (N_14116,N_11582,N_9696);
nand U14117 (N_14117,N_10861,N_10636);
or U14118 (N_14118,N_10404,N_11693);
or U14119 (N_14119,N_11385,N_10708);
and U14120 (N_14120,N_9829,N_10291);
nor U14121 (N_14121,N_9333,N_11251);
nor U14122 (N_14122,N_9221,N_11259);
or U14123 (N_14123,N_9455,N_11218);
nand U14124 (N_14124,N_9195,N_11976);
nor U14125 (N_14125,N_9648,N_11030);
or U14126 (N_14126,N_9940,N_9633);
nor U14127 (N_14127,N_10752,N_10334);
xnor U14128 (N_14128,N_11058,N_9678);
nand U14129 (N_14129,N_11256,N_9953);
nand U14130 (N_14130,N_9235,N_10208);
and U14131 (N_14131,N_10315,N_11736);
or U14132 (N_14132,N_9927,N_10956);
nor U14133 (N_14133,N_9124,N_9242);
and U14134 (N_14134,N_11630,N_11596);
nand U14135 (N_14135,N_11983,N_10519);
and U14136 (N_14136,N_9986,N_10127);
or U14137 (N_14137,N_10195,N_11237);
nor U14138 (N_14138,N_11072,N_9507);
and U14139 (N_14139,N_10132,N_10133);
xnor U14140 (N_14140,N_9093,N_11725);
xor U14141 (N_14141,N_10030,N_11390);
nor U14142 (N_14142,N_9217,N_10157);
nor U14143 (N_14143,N_10421,N_10683);
or U14144 (N_14144,N_9461,N_10159);
nand U14145 (N_14145,N_11402,N_10433);
or U14146 (N_14146,N_11768,N_9084);
nor U14147 (N_14147,N_11691,N_9409);
nand U14148 (N_14148,N_9287,N_10489);
and U14149 (N_14149,N_9253,N_10811);
nand U14150 (N_14150,N_9727,N_11556);
or U14151 (N_14151,N_9720,N_9308);
nand U14152 (N_14152,N_9526,N_9488);
and U14153 (N_14153,N_9506,N_9461);
nor U14154 (N_14154,N_10963,N_9482);
or U14155 (N_14155,N_9900,N_10199);
nand U14156 (N_14156,N_11419,N_11366);
or U14157 (N_14157,N_10274,N_10200);
nand U14158 (N_14158,N_9725,N_10382);
nand U14159 (N_14159,N_10442,N_10330);
and U14160 (N_14160,N_9613,N_10417);
and U14161 (N_14161,N_10619,N_9610);
nor U14162 (N_14162,N_11359,N_9758);
or U14163 (N_14163,N_9837,N_9596);
xnor U14164 (N_14164,N_10360,N_10084);
xor U14165 (N_14165,N_9895,N_11251);
nand U14166 (N_14166,N_9139,N_11151);
nand U14167 (N_14167,N_9218,N_10107);
and U14168 (N_14168,N_10728,N_9498);
or U14169 (N_14169,N_10442,N_11410);
nand U14170 (N_14170,N_11408,N_9752);
or U14171 (N_14171,N_9994,N_9019);
nor U14172 (N_14172,N_9760,N_11236);
nor U14173 (N_14173,N_10101,N_11561);
xor U14174 (N_14174,N_11289,N_9297);
nand U14175 (N_14175,N_9005,N_11150);
or U14176 (N_14176,N_9003,N_11818);
nor U14177 (N_14177,N_9834,N_11907);
or U14178 (N_14178,N_9005,N_10522);
nor U14179 (N_14179,N_10544,N_11768);
nand U14180 (N_14180,N_9180,N_11942);
nor U14181 (N_14181,N_10113,N_11250);
nor U14182 (N_14182,N_11545,N_10754);
or U14183 (N_14183,N_11041,N_9288);
or U14184 (N_14184,N_11783,N_10276);
xor U14185 (N_14185,N_10382,N_11720);
nand U14186 (N_14186,N_11763,N_9920);
nor U14187 (N_14187,N_11531,N_11019);
nor U14188 (N_14188,N_11085,N_10422);
or U14189 (N_14189,N_11574,N_11558);
nor U14190 (N_14190,N_9241,N_11947);
or U14191 (N_14191,N_11471,N_9451);
nand U14192 (N_14192,N_10584,N_10716);
nand U14193 (N_14193,N_11656,N_10685);
xnor U14194 (N_14194,N_11564,N_11756);
or U14195 (N_14195,N_9988,N_10724);
and U14196 (N_14196,N_11663,N_11466);
nand U14197 (N_14197,N_9370,N_11170);
and U14198 (N_14198,N_9469,N_9368);
and U14199 (N_14199,N_9515,N_9775);
and U14200 (N_14200,N_11777,N_11201);
nand U14201 (N_14201,N_9568,N_11016);
nand U14202 (N_14202,N_11867,N_10848);
nand U14203 (N_14203,N_10200,N_9926);
and U14204 (N_14204,N_10359,N_11644);
and U14205 (N_14205,N_9157,N_10658);
or U14206 (N_14206,N_9772,N_9747);
nor U14207 (N_14207,N_9664,N_11451);
or U14208 (N_14208,N_11036,N_9067);
or U14209 (N_14209,N_9235,N_11106);
nor U14210 (N_14210,N_10296,N_9214);
and U14211 (N_14211,N_10100,N_10389);
and U14212 (N_14212,N_9645,N_9608);
and U14213 (N_14213,N_10597,N_9780);
and U14214 (N_14214,N_9288,N_10113);
nor U14215 (N_14215,N_9953,N_11586);
or U14216 (N_14216,N_10963,N_9887);
and U14217 (N_14217,N_9476,N_10535);
and U14218 (N_14218,N_9446,N_10490);
nand U14219 (N_14219,N_10092,N_10260);
nand U14220 (N_14220,N_11246,N_10298);
and U14221 (N_14221,N_10204,N_9592);
or U14222 (N_14222,N_10680,N_11645);
and U14223 (N_14223,N_10041,N_9880);
and U14224 (N_14224,N_9428,N_11280);
nand U14225 (N_14225,N_11893,N_11170);
or U14226 (N_14226,N_10026,N_10111);
nor U14227 (N_14227,N_11082,N_9678);
nand U14228 (N_14228,N_10182,N_9820);
xor U14229 (N_14229,N_10581,N_11588);
nand U14230 (N_14230,N_11135,N_9713);
or U14231 (N_14231,N_11262,N_11917);
nor U14232 (N_14232,N_11601,N_9194);
nand U14233 (N_14233,N_10169,N_10320);
or U14234 (N_14234,N_11685,N_10268);
or U14235 (N_14235,N_9193,N_9929);
nand U14236 (N_14236,N_9397,N_9705);
nor U14237 (N_14237,N_10481,N_11794);
nand U14238 (N_14238,N_10694,N_11386);
nand U14239 (N_14239,N_10008,N_11687);
nand U14240 (N_14240,N_10505,N_10667);
or U14241 (N_14241,N_10605,N_9800);
nand U14242 (N_14242,N_10264,N_11862);
nor U14243 (N_14243,N_10036,N_9097);
or U14244 (N_14244,N_11028,N_9462);
nor U14245 (N_14245,N_11693,N_11621);
nand U14246 (N_14246,N_10341,N_10206);
nand U14247 (N_14247,N_10147,N_10194);
or U14248 (N_14248,N_10261,N_10437);
nor U14249 (N_14249,N_9320,N_10568);
nor U14250 (N_14250,N_11514,N_10214);
nor U14251 (N_14251,N_11243,N_9643);
or U14252 (N_14252,N_9783,N_9073);
nand U14253 (N_14253,N_9448,N_10054);
nor U14254 (N_14254,N_10046,N_10389);
nand U14255 (N_14255,N_9571,N_9732);
and U14256 (N_14256,N_10579,N_11088);
or U14257 (N_14257,N_9785,N_10800);
nand U14258 (N_14258,N_9660,N_11474);
nor U14259 (N_14259,N_9170,N_11830);
and U14260 (N_14260,N_11223,N_9931);
xnor U14261 (N_14261,N_9843,N_9455);
nor U14262 (N_14262,N_11139,N_11092);
nand U14263 (N_14263,N_11757,N_9216);
or U14264 (N_14264,N_11902,N_11127);
nor U14265 (N_14265,N_11764,N_9589);
nand U14266 (N_14266,N_11495,N_9887);
or U14267 (N_14267,N_10971,N_10848);
xnor U14268 (N_14268,N_11043,N_11678);
nand U14269 (N_14269,N_10050,N_9624);
nand U14270 (N_14270,N_9062,N_10419);
and U14271 (N_14271,N_10198,N_10242);
nor U14272 (N_14272,N_9929,N_9598);
and U14273 (N_14273,N_10580,N_9762);
and U14274 (N_14274,N_10572,N_10800);
xnor U14275 (N_14275,N_9056,N_9708);
or U14276 (N_14276,N_10861,N_11968);
or U14277 (N_14277,N_11602,N_10661);
nor U14278 (N_14278,N_9264,N_10314);
and U14279 (N_14279,N_11923,N_9256);
and U14280 (N_14280,N_10013,N_10903);
or U14281 (N_14281,N_10967,N_10946);
or U14282 (N_14282,N_11072,N_9560);
nor U14283 (N_14283,N_9541,N_9835);
and U14284 (N_14284,N_11870,N_10296);
nand U14285 (N_14285,N_11208,N_9341);
nand U14286 (N_14286,N_9273,N_9999);
and U14287 (N_14287,N_10762,N_11054);
and U14288 (N_14288,N_11591,N_10317);
or U14289 (N_14289,N_10109,N_9483);
nand U14290 (N_14290,N_10979,N_9221);
or U14291 (N_14291,N_11622,N_9264);
and U14292 (N_14292,N_10027,N_9759);
or U14293 (N_14293,N_10526,N_10761);
and U14294 (N_14294,N_10479,N_11816);
or U14295 (N_14295,N_9097,N_10681);
nand U14296 (N_14296,N_9607,N_9095);
or U14297 (N_14297,N_9036,N_9359);
nand U14298 (N_14298,N_9017,N_10498);
and U14299 (N_14299,N_10241,N_10159);
nor U14300 (N_14300,N_10393,N_9513);
and U14301 (N_14301,N_11187,N_11766);
nand U14302 (N_14302,N_9335,N_11983);
or U14303 (N_14303,N_10546,N_9115);
or U14304 (N_14304,N_11232,N_11953);
nand U14305 (N_14305,N_10165,N_11749);
and U14306 (N_14306,N_11987,N_9583);
or U14307 (N_14307,N_10139,N_11979);
nand U14308 (N_14308,N_9559,N_11950);
nor U14309 (N_14309,N_11610,N_9979);
and U14310 (N_14310,N_10523,N_11761);
and U14311 (N_14311,N_11453,N_10131);
nor U14312 (N_14312,N_11108,N_9351);
and U14313 (N_14313,N_9507,N_10469);
and U14314 (N_14314,N_9595,N_9122);
nor U14315 (N_14315,N_9809,N_10362);
and U14316 (N_14316,N_10214,N_10885);
and U14317 (N_14317,N_10302,N_11112);
nand U14318 (N_14318,N_10337,N_9466);
and U14319 (N_14319,N_11937,N_10733);
nor U14320 (N_14320,N_10252,N_9233);
nor U14321 (N_14321,N_10404,N_10892);
nor U14322 (N_14322,N_9230,N_10905);
and U14323 (N_14323,N_11675,N_10538);
nand U14324 (N_14324,N_9715,N_9545);
or U14325 (N_14325,N_9357,N_10274);
or U14326 (N_14326,N_11123,N_10853);
nor U14327 (N_14327,N_11788,N_9532);
or U14328 (N_14328,N_9409,N_9340);
nand U14329 (N_14329,N_10045,N_9873);
or U14330 (N_14330,N_9314,N_11396);
and U14331 (N_14331,N_11453,N_10269);
and U14332 (N_14332,N_9010,N_9198);
or U14333 (N_14333,N_11772,N_10830);
xnor U14334 (N_14334,N_9845,N_11602);
or U14335 (N_14335,N_11024,N_10963);
nor U14336 (N_14336,N_11976,N_9315);
nor U14337 (N_14337,N_9142,N_10010);
and U14338 (N_14338,N_10752,N_11336);
nor U14339 (N_14339,N_11211,N_10249);
or U14340 (N_14340,N_10729,N_11579);
and U14341 (N_14341,N_10333,N_11569);
nor U14342 (N_14342,N_10616,N_10136);
or U14343 (N_14343,N_9371,N_11311);
or U14344 (N_14344,N_10675,N_11188);
nor U14345 (N_14345,N_9972,N_9404);
nand U14346 (N_14346,N_10048,N_9912);
nor U14347 (N_14347,N_10434,N_9043);
and U14348 (N_14348,N_10741,N_9756);
or U14349 (N_14349,N_9838,N_10813);
nand U14350 (N_14350,N_9704,N_9380);
nor U14351 (N_14351,N_9226,N_9718);
or U14352 (N_14352,N_9986,N_11211);
and U14353 (N_14353,N_11264,N_9964);
nor U14354 (N_14354,N_9650,N_10485);
nand U14355 (N_14355,N_10959,N_10703);
nor U14356 (N_14356,N_11402,N_9312);
nand U14357 (N_14357,N_10791,N_11697);
xnor U14358 (N_14358,N_9969,N_9149);
nand U14359 (N_14359,N_10519,N_10730);
nor U14360 (N_14360,N_10108,N_11313);
nand U14361 (N_14361,N_10005,N_10319);
nor U14362 (N_14362,N_9808,N_11533);
xnor U14363 (N_14363,N_10080,N_10849);
and U14364 (N_14364,N_11020,N_10855);
and U14365 (N_14365,N_9269,N_10664);
nand U14366 (N_14366,N_9061,N_10285);
nand U14367 (N_14367,N_11972,N_10843);
nand U14368 (N_14368,N_9707,N_9599);
or U14369 (N_14369,N_10975,N_11453);
nor U14370 (N_14370,N_9392,N_10726);
nor U14371 (N_14371,N_9444,N_9270);
or U14372 (N_14372,N_11340,N_9401);
or U14373 (N_14373,N_9634,N_9480);
nand U14374 (N_14374,N_9536,N_9818);
nand U14375 (N_14375,N_10777,N_9699);
nand U14376 (N_14376,N_9477,N_9483);
nor U14377 (N_14377,N_10618,N_10829);
xor U14378 (N_14378,N_11129,N_10256);
nor U14379 (N_14379,N_11664,N_10173);
nor U14380 (N_14380,N_9124,N_10283);
and U14381 (N_14381,N_9913,N_10181);
nor U14382 (N_14382,N_11338,N_9577);
nand U14383 (N_14383,N_11950,N_9237);
nor U14384 (N_14384,N_9827,N_9057);
or U14385 (N_14385,N_10678,N_10242);
nand U14386 (N_14386,N_11855,N_11201);
xnor U14387 (N_14387,N_9218,N_11705);
or U14388 (N_14388,N_9111,N_11707);
nand U14389 (N_14389,N_11029,N_10035);
nor U14390 (N_14390,N_10919,N_9639);
and U14391 (N_14391,N_11546,N_10400);
nand U14392 (N_14392,N_10764,N_9380);
nor U14393 (N_14393,N_11658,N_9824);
or U14394 (N_14394,N_9671,N_11656);
or U14395 (N_14395,N_10135,N_10020);
and U14396 (N_14396,N_9519,N_11735);
nand U14397 (N_14397,N_10091,N_11183);
nand U14398 (N_14398,N_9857,N_9282);
or U14399 (N_14399,N_9922,N_10942);
or U14400 (N_14400,N_9306,N_9379);
nor U14401 (N_14401,N_10955,N_10968);
and U14402 (N_14402,N_10448,N_9580);
and U14403 (N_14403,N_9661,N_11572);
nand U14404 (N_14404,N_10440,N_11152);
xnor U14405 (N_14405,N_11776,N_10467);
nand U14406 (N_14406,N_9012,N_9502);
or U14407 (N_14407,N_9439,N_9910);
nand U14408 (N_14408,N_10187,N_10350);
or U14409 (N_14409,N_11226,N_11119);
nand U14410 (N_14410,N_11576,N_9160);
and U14411 (N_14411,N_10053,N_9152);
and U14412 (N_14412,N_9230,N_11874);
nor U14413 (N_14413,N_11606,N_10205);
and U14414 (N_14414,N_11300,N_9940);
nor U14415 (N_14415,N_9079,N_10636);
or U14416 (N_14416,N_11231,N_11755);
nand U14417 (N_14417,N_9684,N_11168);
or U14418 (N_14418,N_9967,N_11754);
nor U14419 (N_14419,N_10455,N_10462);
nor U14420 (N_14420,N_11752,N_10375);
nor U14421 (N_14421,N_9667,N_9254);
nor U14422 (N_14422,N_10252,N_10778);
and U14423 (N_14423,N_10230,N_10280);
nand U14424 (N_14424,N_11755,N_11654);
nor U14425 (N_14425,N_10940,N_9876);
nand U14426 (N_14426,N_10252,N_9330);
nand U14427 (N_14427,N_11311,N_9646);
nand U14428 (N_14428,N_9159,N_11429);
and U14429 (N_14429,N_11835,N_10680);
and U14430 (N_14430,N_11714,N_10893);
or U14431 (N_14431,N_11315,N_11220);
and U14432 (N_14432,N_9866,N_9842);
and U14433 (N_14433,N_9934,N_9218);
and U14434 (N_14434,N_11801,N_10265);
and U14435 (N_14435,N_9789,N_10924);
and U14436 (N_14436,N_10573,N_9393);
or U14437 (N_14437,N_10309,N_10430);
or U14438 (N_14438,N_10102,N_11588);
and U14439 (N_14439,N_9019,N_11899);
nand U14440 (N_14440,N_10842,N_10003);
and U14441 (N_14441,N_10056,N_10214);
xor U14442 (N_14442,N_9493,N_9877);
and U14443 (N_14443,N_9976,N_9770);
nand U14444 (N_14444,N_10308,N_11989);
and U14445 (N_14445,N_9592,N_10234);
or U14446 (N_14446,N_9995,N_11697);
nor U14447 (N_14447,N_9651,N_10085);
and U14448 (N_14448,N_9988,N_11755);
nand U14449 (N_14449,N_9993,N_10446);
or U14450 (N_14450,N_11952,N_10843);
or U14451 (N_14451,N_10499,N_10167);
and U14452 (N_14452,N_10728,N_9962);
nor U14453 (N_14453,N_9443,N_11128);
nor U14454 (N_14454,N_11307,N_11353);
nand U14455 (N_14455,N_9398,N_11000);
and U14456 (N_14456,N_10995,N_9326);
or U14457 (N_14457,N_11468,N_9624);
nor U14458 (N_14458,N_11307,N_9639);
nand U14459 (N_14459,N_9291,N_10060);
nand U14460 (N_14460,N_10312,N_10677);
nand U14461 (N_14461,N_11690,N_10360);
nand U14462 (N_14462,N_10733,N_10541);
or U14463 (N_14463,N_11390,N_10193);
xor U14464 (N_14464,N_10198,N_11265);
nor U14465 (N_14465,N_11179,N_11385);
and U14466 (N_14466,N_11425,N_10977);
nand U14467 (N_14467,N_9197,N_10034);
or U14468 (N_14468,N_9275,N_9827);
and U14469 (N_14469,N_9844,N_10364);
nand U14470 (N_14470,N_11284,N_11588);
or U14471 (N_14471,N_11979,N_9220);
nand U14472 (N_14472,N_9030,N_9046);
nand U14473 (N_14473,N_9691,N_10442);
and U14474 (N_14474,N_10905,N_10423);
and U14475 (N_14475,N_9902,N_11110);
nand U14476 (N_14476,N_10539,N_11201);
and U14477 (N_14477,N_11526,N_11278);
nand U14478 (N_14478,N_10174,N_9690);
or U14479 (N_14479,N_10036,N_11126);
and U14480 (N_14480,N_10879,N_11607);
nor U14481 (N_14481,N_9079,N_9297);
or U14482 (N_14482,N_10105,N_9109);
nor U14483 (N_14483,N_9166,N_9054);
and U14484 (N_14484,N_9346,N_10627);
nand U14485 (N_14485,N_9301,N_9605);
or U14486 (N_14486,N_10615,N_9911);
nor U14487 (N_14487,N_10006,N_11414);
nand U14488 (N_14488,N_11001,N_10492);
and U14489 (N_14489,N_9313,N_10990);
nor U14490 (N_14490,N_9077,N_11422);
nor U14491 (N_14491,N_9670,N_11668);
and U14492 (N_14492,N_9264,N_10074);
nand U14493 (N_14493,N_11892,N_9847);
nor U14494 (N_14494,N_9021,N_9243);
nand U14495 (N_14495,N_10781,N_11502);
and U14496 (N_14496,N_9693,N_9786);
nor U14497 (N_14497,N_11557,N_11309);
or U14498 (N_14498,N_11642,N_9618);
or U14499 (N_14499,N_10209,N_9079);
nor U14500 (N_14500,N_9779,N_11960);
nor U14501 (N_14501,N_11934,N_11052);
nand U14502 (N_14502,N_10819,N_11578);
nand U14503 (N_14503,N_9627,N_9706);
nand U14504 (N_14504,N_10966,N_11308);
nand U14505 (N_14505,N_10283,N_10598);
and U14506 (N_14506,N_10453,N_10261);
or U14507 (N_14507,N_10712,N_9802);
nor U14508 (N_14508,N_10491,N_10246);
nor U14509 (N_14509,N_10123,N_10217);
nand U14510 (N_14510,N_10960,N_10299);
nor U14511 (N_14511,N_10517,N_10101);
and U14512 (N_14512,N_10166,N_11069);
nand U14513 (N_14513,N_10229,N_11770);
and U14514 (N_14514,N_10014,N_10275);
or U14515 (N_14515,N_11706,N_10018);
or U14516 (N_14516,N_11183,N_9425);
and U14517 (N_14517,N_11873,N_10722);
or U14518 (N_14518,N_11848,N_10831);
and U14519 (N_14519,N_11919,N_11496);
and U14520 (N_14520,N_10870,N_10040);
nor U14521 (N_14521,N_11234,N_11717);
or U14522 (N_14522,N_9450,N_10172);
and U14523 (N_14523,N_11467,N_9492);
nor U14524 (N_14524,N_9569,N_11653);
xnor U14525 (N_14525,N_10778,N_11168);
nor U14526 (N_14526,N_9311,N_11829);
nor U14527 (N_14527,N_11489,N_9765);
and U14528 (N_14528,N_9929,N_11052);
nand U14529 (N_14529,N_9439,N_9769);
and U14530 (N_14530,N_11907,N_11084);
and U14531 (N_14531,N_11073,N_9137);
or U14532 (N_14532,N_10601,N_9284);
or U14533 (N_14533,N_9901,N_11678);
nand U14534 (N_14534,N_9345,N_9905);
or U14535 (N_14535,N_9285,N_9911);
or U14536 (N_14536,N_11258,N_10900);
and U14537 (N_14537,N_11643,N_11750);
nand U14538 (N_14538,N_11284,N_11881);
nand U14539 (N_14539,N_9522,N_9997);
nor U14540 (N_14540,N_9261,N_11430);
or U14541 (N_14541,N_11565,N_11437);
nand U14542 (N_14542,N_11999,N_9022);
or U14543 (N_14543,N_10063,N_9500);
or U14544 (N_14544,N_9682,N_9378);
and U14545 (N_14545,N_11202,N_9027);
nand U14546 (N_14546,N_11822,N_11186);
and U14547 (N_14547,N_11998,N_10790);
and U14548 (N_14548,N_11092,N_9214);
nor U14549 (N_14549,N_11168,N_9368);
nand U14550 (N_14550,N_9005,N_10529);
and U14551 (N_14551,N_9384,N_10796);
or U14552 (N_14552,N_11772,N_10146);
and U14553 (N_14553,N_10576,N_9769);
and U14554 (N_14554,N_10858,N_9738);
and U14555 (N_14555,N_11642,N_11417);
and U14556 (N_14556,N_9905,N_11947);
or U14557 (N_14557,N_9160,N_10151);
and U14558 (N_14558,N_11039,N_10638);
nand U14559 (N_14559,N_10479,N_10008);
nand U14560 (N_14560,N_10540,N_11400);
and U14561 (N_14561,N_10061,N_11187);
nand U14562 (N_14562,N_10977,N_11916);
and U14563 (N_14563,N_11498,N_11122);
or U14564 (N_14564,N_11929,N_10802);
nor U14565 (N_14565,N_10560,N_10730);
and U14566 (N_14566,N_10783,N_9758);
or U14567 (N_14567,N_9922,N_11576);
and U14568 (N_14568,N_9393,N_10746);
or U14569 (N_14569,N_10957,N_11563);
nor U14570 (N_14570,N_10802,N_11423);
or U14571 (N_14571,N_10410,N_10908);
and U14572 (N_14572,N_11619,N_9893);
and U14573 (N_14573,N_9865,N_11380);
xnor U14574 (N_14574,N_11407,N_9409);
or U14575 (N_14575,N_9482,N_9674);
or U14576 (N_14576,N_9310,N_9518);
nor U14577 (N_14577,N_10379,N_9125);
nand U14578 (N_14578,N_11884,N_10632);
nor U14579 (N_14579,N_9136,N_9827);
and U14580 (N_14580,N_9929,N_9379);
nor U14581 (N_14581,N_9493,N_10798);
nand U14582 (N_14582,N_9188,N_9445);
xnor U14583 (N_14583,N_10782,N_11619);
nand U14584 (N_14584,N_10355,N_11806);
nor U14585 (N_14585,N_9552,N_9180);
nand U14586 (N_14586,N_10287,N_9790);
or U14587 (N_14587,N_10863,N_9818);
or U14588 (N_14588,N_11593,N_10020);
nand U14589 (N_14589,N_11840,N_11220);
nand U14590 (N_14590,N_10208,N_11006);
and U14591 (N_14591,N_11758,N_10189);
nand U14592 (N_14592,N_10115,N_11280);
nor U14593 (N_14593,N_11465,N_9811);
and U14594 (N_14594,N_11536,N_11940);
and U14595 (N_14595,N_11691,N_11155);
nand U14596 (N_14596,N_9114,N_10782);
nand U14597 (N_14597,N_9193,N_10341);
or U14598 (N_14598,N_9675,N_9231);
and U14599 (N_14599,N_10112,N_10485);
nand U14600 (N_14600,N_11677,N_11791);
or U14601 (N_14601,N_9649,N_9252);
nor U14602 (N_14602,N_9995,N_9485);
nor U14603 (N_14603,N_10112,N_11453);
and U14604 (N_14604,N_10478,N_11612);
and U14605 (N_14605,N_10304,N_11328);
and U14606 (N_14606,N_10972,N_9905);
or U14607 (N_14607,N_10246,N_11923);
nor U14608 (N_14608,N_11758,N_11169);
or U14609 (N_14609,N_9566,N_11786);
nor U14610 (N_14610,N_9635,N_11552);
nand U14611 (N_14611,N_11381,N_10536);
or U14612 (N_14612,N_11436,N_11957);
nand U14613 (N_14613,N_9486,N_11153);
or U14614 (N_14614,N_10435,N_9638);
and U14615 (N_14615,N_11460,N_9430);
and U14616 (N_14616,N_10159,N_10790);
or U14617 (N_14617,N_11566,N_10244);
or U14618 (N_14618,N_11896,N_10352);
or U14619 (N_14619,N_11729,N_10549);
nor U14620 (N_14620,N_9129,N_10762);
xor U14621 (N_14621,N_11777,N_9597);
nand U14622 (N_14622,N_10943,N_11378);
and U14623 (N_14623,N_10470,N_9083);
or U14624 (N_14624,N_10166,N_9737);
and U14625 (N_14625,N_11674,N_9323);
or U14626 (N_14626,N_9895,N_11315);
xor U14627 (N_14627,N_11543,N_11939);
nand U14628 (N_14628,N_10512,N_9086);
nand U14629 (N_14629,N_9352,N_10956);
or U14630 (N_14630,N_11570,N_9687);
and U14631 (N_14631,N_10070,N_9719);
or U14632 (N_14632,N_11423,N_10016);
or U14633 (N_14633,N_10950,N_9505);
nor U14634 (N_14634,N_9676,N_9860);
or U14635 (N_14635,N_11650,N_11059);
and U14636 (N_14636,N_9466,N_9007);
nor U14637 (N_14637,N_10013,N_11306);
nor U14638 (N_14638,N_11978,N_11473);
nor U14639 (N_14639,N_11505,N_10814);
or U14640 (N_14640,N_9565,N_10086);
and U14641 (N_14641,N_10927,N_11476);
or U14642 (N_14642,N_11043,N_11695);
or U14643 (N_14643,N_9725,N_11371);
or U14644 (N_14644,N_9877,N_10278);
nor U14645 (N_14645,N_10034,N_10792);
and U14646 (N_14646,N_10830,N_10395);
and U14647 (N_14647,N_9616,N_9711);
nand U14648 (N_14648,N_9781,N_10599);
or U14649 (N_14649,N_9414,N_11444);
nor U14650 (N_14650,N_11120,N_10913);
nand U14651 (N_14651,N_10116,N_9031);
xnor U14652 (N_14652,N_10114,N_10908);
or U14653 (N_14653,N_11281,N_9727);
nand U14654 (N_14654,N_11765,N_11137);
nor U14655 (N_14655,N_11894,N_9034);
and U14656 (N_14656,N_9375,N_9470);
or U14657 (N_14657,N_11267,N_10068);
and U14658 (N_14658,N_9224,N_11489);
and U14659 (N_14659,N_11454,N_10016);
nand U14660 (N_14660,N_9079,N_10390);
and U14661 (N_14661,N_9153,N_10238);
nand U14662 (N_14662,N_11618,N_11828);
and U14663 (N_14663,N_10953,N_11575);
nand U14664 (N_14664,N_11592,N_9794);
nand U14665 (N_14665,N_11786,N_10447);
nor U14666 (N_14666,N_10079,N_10998);
or U14667 (N_14667,N_11822,N_11576);
or U14668 (N_14668,N_11476,N_10535);
or U14669 (N_14669,N_10207,N_11424);
nor U14670 (N_14670,N_10825,N_11085);
and U14671 (N_14671,N_9136,N_9297);
and U14672 (N_14672,N_11316,N_11146);
nand U14673 (N_14673,N_11396,N_11865);
nor U14674 (N_14674,N_11247,N_11920);
nor U14675 (N_14675,N_11367,N_10929);
and U14676 (N_14676,N_10935,N_11712);
and U14677 (N_14677,N_10074,N_11413);
and U14678 (N_14678,N_9860,N_9059);
nand U14679 (N_14679,N_9958,N_11969);
nor U14680 (N_14680,N_9956,N_11497);
and U14681 (N_14681,N_9768,N_11648);
and U14682 (N_14682,N_11710,N_10326);
nand U14683 (N_14683,N_10907,N_10507);
nor U14684 (N_14684,N_10738,N_10706);
and U14685 (N_14685,N_9531,N_9821);
nor U14686 (N_14686,N_10220,N_11894);
nor U14687 (N_14687,N_11363,N_9699);
or U14688 (N_14688,N_9078,N_11420);
or U14689 (N_14689,N_11033,N_11540);
or U14690 (N_14690,N_9679,N_11398);
xor U14691 (N_14691,N_11718,N_10490);
nor U14692 (N_14692,N_9208,N_10863);
and U14693 (N_14693,N_9263,N_10869);
and U14694 (N_14694,N_11865,N_10590);
nor U14695 (N_14695,N_9890,N_11587);
nor U14696 (N_14696,N_10314,N_9028);
and U14697 (N_14697,N_9899,N_10976);
nand U14698 (N_14698,N_9232,N_10223);
nor U14699 (N_14699,N_11222,N_10571);
nor U14700 (N_14700,N_10906,N_11422);
and U14701 (N_14701,N_9478,N_10912);
nand U14702 (N_14702,N_9505,N_9135);
nand U14703 (N_14703,N_10207,N_11137);
or U14704 (N_14704,N_11683,N_11137);
and U14705 (N_14705,N_10038,N_9938);
xor U14706 (N_14706,N_10098,N_9687);
nor U14707 (N_14707,N_11603,N_11938);
nor U14708 (N_14708,N_11018,N_10321);
or U14709 (N_14709,N_10884,N_9654);
nor U14710 (N_14710,N_9544,N_11004);
nor U14711 (N_14711,N_10535,N_9002);
or U14712 (N_14712,N_10178,N_9105);
nand U14713 (N_14713,N_9377,N_11311);
and U14714 (N_14714,N_11665,N_10209);
nor U14715 (N_14715,N_9338,N_11782);
or U14716 (N_14716,N_10509,N_11571);
nand U14717 (N_14717,N_11309,N_11766);
and U14718 (N_14718,N_11351,N_9970);
nand U14719 (N_14719,N_11292,N_10447);
and U14720 (N_14720,N_11286,N_11033);
nand U14721 (N_14721,N_10298,N_9093);
nand U14722 (N_14722,N_11953,N_11235);
and U14723 (N_14723,N_9895,N_10533);
nor U14724 (N_14724,N_10531,N_10583);
or U14725 (N_14725,N_9892,N_11543);
nand U14726 (N_14726,N_9917,N_10711);
xor U14727 (N_14727,N_11654,N_9946);
or U14728 (N_14728,N_11227,N_9804);
and U14729 (N_14729,N_9681,N_9744);
and U14730 (N_14730,N_11463,N_11650);
or U14731 (N_14731,N_9816,N_10976);
nor U14732 (N_14732,N_10395,N_9292);
nor U14733 (N_14733,N_9172,N_10420);
and U14734 (N_14734,N_11521,N_9137);
nand U14735 (N_14735,N_11402,N_10238);
and U14736 (N_14736,N_10038,N_9380);
nor U14737 (N_14737,N_10063,N_9667);
nor U14738 (N_14738,N_9850,N_9545);
or U14739 (N_14739,N_9874,N_9444);
nor U14740 (N_14740,N_9945,N_11900);
nand U14741 (N_14741,N_11941,N_9287);
nand U14742 (N_14742,N_11332,N_9867);
or U14743 (N_14743,N_10681,N_10078);
nor U14744 (N_14744,N_9845,N_9887);
or U14745 (N_14745,N_11085,N_11378);
and U14746 (N_14746,N_10983,N_10181);
or U14747 (N_14747,N_11785,N_9419);
or U14748 (N_14748,N_11069,N_9309);
nand U14749 (N_14749,N_9086,N_11825);
or U14750 (N_14750,N_9723,N_11968);
xnor U14751 (N_14751,N_10250,N_10887);
nor U14752 (N_14752,N_9497,N_9357);
nand U14753 (N_14753,N_9290,N_10351);
or U14754 (N_14754,N_9036,N_9710);
and U14755 (N_14755,N_10075,N_11890);
nor U14756 (N_14756,N_9871,N_9614);
nor U14757 (N_14757,N_9519,N_10125);
or U14758 (N_14758,N_11269,N_11833);
or U14759 (N_14759,N_10144,N_9176);
nor U14760 (N_14760,N_10576,N_11306);
nor U14761 (N_14761,N_9933,N_10086);
nand U14762 (N_14762,N_11762,N_9965);
and U14763 (N_14763,N_10765,N_9212);
nor U14764 (N_14764,N_11089,N_10640);
and U14765 (N_14765,N_10346,N_11310);
and U14766 (N_14766,N_10841,N_9685);
nor U14767 (N_14767,N_9622,N_10164);
nand U14768 (N_14768,N_11277,N_11743);
and U14769 (N_14769,N_11276,N_10989);
nand U14770 (N_14770,N_9660,N_10893);
nand U14771 (N_14771,N_10676,N_9349);
or U14772 (N_14772,N_10141,N_10020);
nand U14773 (N_14773,N_10336,N_10188);
and U14774 (N_14774,N_11099,N_11048);
nand U14775 (N_14775,N_10342,N_11617);
nand U14776 (N_14776,N_11248,N_9913);
nand U14777 (N_14777,N_10893,N_10692);
nand U14778 (N_14778,N_11025,N_9790);
or U14779 (N_14779,N_9436,N_9477);
nor U14780 (N_14780,N_10571,N_9375);
nor U14781 (N_14781,N_9998,N_10540);
and U14782 (N_14782,N_9882,N_11838);
and U14783 (N_14783,N_11584,N_9680);
or U14784 (N_14784,N_11101,N_10447);
nand U14785 (N_14785,N_9271,N_9903);
or U14786 (N_14786,N_9608,N_10341);
or U14787 (N_14787,N_10296,N_10767);
nand U14788 (N_14788,N_11489,N_9674);
nor U14789 (N_14789,N_11380,N_9894);
or U14790 (N_14790,N_11688,N_10680);
nor U14791 (N_14791,N_10156,N_11691);
nor U14792 (N_14792,N_9188,N_11642);
nand U14793 (N_14793,N_9583,N_9513);
nor U14794 (N_14794,N_11526,N_9000);
and U14795 (N_14795,N_11976,N_11141);
and U14796 (N_14796,N_10496,N_11754);
nand U14797 (N_14797,N_10879,N_11436);
or U14798 (N_14798,N_11259,N_11679);
nor U14799 (N_14799,N_10107,N_9200);
and U14800 (N_14800,N_9528,N_11871);
nand U14801 (N_14801,N_11579,N_10918);
or U14802 (N_14802,N_10994,N_11439);
or U14803 (N_14803,N_9674,N_9312);
and U14804 (N_14804,N_10595,N_9609);
nor U14805 (N_14805,N_10250,N_11767);
nor U14806 (N_14806,N_9498,N_11522);
or U14807 (N_14807,N_10090,N_9155);
and U14808 (N_14808,N_10970,N_9490);
or U14809 (N_14809,N_9597,N_11672);
and U14810 (N_14810,N_9240,N_9163);
xnor U14811 (N_14811,N_11828,N_11887);
xnor U14812 (N_14812,N_9355,N_10515);
or U14813 (N_14813,N_11213,N_11963);
nor U14814 (N_14814,N_10888,N_9988);
or U14815 (N_14815,N_11054,N_11137);
and U14816 (N_14816,N_11934,N_11806);
xor U14817 (N_14817,N_11468,N_11429);
or U14818 (N_14818,N_10375,N_10260);
nor U14819 (N_14819,N_11680,N_10236);
nor U14820 (N_14820,N_11118,N_11482);
or U14821 (N_14821,N_9982,N_10530);
nor U14822 (N_14822,N_9032,N_11293);
nor U14823 (N_14823,N_10127,N_11674);
nand U14824 (N_14824,N_9604,N_11153);
and U14825 (N_14825,N_10131,N_11699);
and U14826 (N_14826,N_10453,N_10839);
or U14827 (N_14827,N_10167,N_10902);
or U14828 (N_14828,N_10852,N_9175);
or U14829 (N_14829,N_10809,N_10053);
or U14830 (N_14830,N_10158,N_9927);
nand U14831 (N_14831,N_10220,N_10175);
nor U14832 (N_14832,N_9107,N_10747);
and U14833 (N_14833,N_9004,N_10082);
or U14834 (N_14834,N_10322,N_11018);
nor U14835 (N_14835,N_9089,N_9166);
and U14836 (N_14836,N_10228,N_10781);
or U14837 (N_14837,N_9414,N_11562);
nor U14838 (N_14838,N_11671,N_11236);
and U14839 (N_14839,N_11684,N_11958);
and U14840 (N_14840,N_10000,N_11254);
nor U14841 (N_14841,N_9945,N_9992);
nand U14842 (N_14842,N_10814,N_9331);
and U14843 (N_14843,N_10928,N_9159);
and U14844 (N_14844,N_9805,N_11860);
or U14845 (N_14845,N_11625,N_11127);
nand U14846 (N_14846,N_10237,N_10566);
nand U14847 (N_14847,N_10803,N_11065);
nand U14848 (N_14848,N_10263,N_9251);
or U14849 (N_14849,N_9755,N_9019);
and U14850 (N_14850,N_9709,N_9339);
nand U14851 (N_14851,N_10014,N_9688);
nand U14852 (N_14852,N_10714,N_9490);
or U14853 (N_14853,N_10821,N_9711);
and U14854 (N_14854,N_10100,N_10223);
nand U14855 (N_14855,N_9841,N_10137);
nor U14856 (N_14856,N_11868,N_9336);
or U14857 (N_14857,N_10864,N_11698);
and U14858 (N_14858,N_11992,N_10713);
nor U14859 (N_14859,N_9550,N_9934);
and U14860 (N_14860,N_9283,N_11275);
and U14861 (N_14861,N_9489,N_10153);
nor U14862 (N_14862,N_11314,N_9176);
nor U14863 (N_14863,N_10432,N_11050);
nand U14864 (N_14864,N_10617,N_9747);
and U14865 (N_14865,N_9658,N_11604);
or U14866 (N_14866,N_11456,N_10499);
or U14867 (N_14867,N_9157,N_10408);
and U14868 (N_14868,N_10454,N_11387);
and U14869 (N_14869,N_9701,N_11262);
nand U14870 (N_14870,N_11031,N_10270);
or U14871 (N_14871,N_11379,N_9225);
nor U14872 (N_14872,N_9860,N_9033);
nor U14873 (N_14873,N_11750,N_10944);
nand U14874 (N_14874,N_9108,N_9082);
nor U14875 (N_14875,N_10714,N_11032);
nor U14876 (N_14876,N_11762,N_11143);
nand U14877 (N_14877,N_9134,N_11246);
nand U14878 (N_14878,N_11358,N_10740);
and U14879 (N_14879,N_11137,N_10370);
or U14880 (N_14880,N_10800,N_10280);
nand U14881 (N_14881,N_10418,N_10302);
or U14882 (N_14882,N_10983,N_11083);
and U14883 (N_14883,N_9476,N_10111);
and U14884 (N_14884,N_9892,N_9454);
nand U14885 (N_14885,N_9261,N_11278);
or U14886 (N_14886,N_11513,N_9009);
xor U14887 (N_14887,N_11834,N_11288);
or U14888 (N_14888,N_11373,N_9966);
nand U14889 (N_14889,N_9640,N_11273);
or U14890 (N_14890,N_10237,N_11039);
and U14891 (N_14891,N_10207,N_10336);
nor U14892 (N_14892,N_10048,N_10590);
or U14893 (N_14893,N_9533,N_10501);
nor U14894 (N_14894,N_10478,N_11444);
nor U14895 (N_14895,N_10772,N_9411);
and U14896 (N_14896,N_11550,N_9757);
xnor U14897 (N_14897,N_11348,N_10426);
nor U14898 (N_14898,N_9637,N_10400);
and U14899 (N_14899,N_10869,N_11147);
nand U14900 (N_14900,N_9321,N_10494);
nor U14901 (N_14901,N_9729,N_10899);
or U14902 (N_14902,N_11756,N_10563);
nor U14903 (N_14903,N_11743,N_9151);
and U14904 (N_14904,N_9545,N_11518);
nand U14905 (N_14905,N_11118,N_9424);
nand U14906 (N_14906,N_11714,N_10723);
and U14907 (N_14907,N_9245,N_10698);
or U14908 (N_14908,N_9332,N_11828);
nand U14909 (N_14909,N_9118,N_11698);
and U14910 (N_14910,N_9812,N_10394);
nor U14911 (N_14911,N_10224,N_11999);
and U14912 (N_14912,N_10153,N_10662);
and U14913 (N_14913,N_9762,N_10287);
and U14914 (N_14914,N_10757,N_10832);
nand U14915 (N_14915,N_10548,N_11852);
and U14916 (N_14916,N_11642,N_10193);
and U14917 (N_14917,N_11010,N_11522);
and U14918 (N_14918,N_9059,N_11863);
nand U14919 (N_14919,N_11819,N_9208);
and U14920 (N_14920,N_9060,N_10603);
nand U14921 (N_14921,N_11861,N_10174);
nor U14922 (N_14922,N_10754,N_11096);
or U14923 (N_14923,N_11416,N_9874);
or U14924 (N_14924,N_9814,N_9967);
nand U14925 (N_14925,N_10416,N_10136);
or U14926 (N_14926,N_9287,N_11203);
xor U14927 (N_14927,N_9934,N_11019);
or U14928 (N_14928,N_11040,N_10711);
or U14929 (N_14929,N_10438,N_10346);
nand U14930 (N_14930,N_11534,N_9431);
nand U14931 (N_14931,N_9383,N_10207);
nor U14932 (N_14932,N_10504,N_9770);
nor U14933 (N_14933,N_9747,N_9643);
and U14934 (N_14934,N_11651,N_9792);
nor U14935 (N_14935,N_10889,N_11604);
nor U14936 (N_14936,N_10447,N_10845);
nand U14937 (N_14937,N_10693,N_11935);
nor U14938 (N_14938,N_10516,N_11584);
nor U14939 (N_14939,N_9718,N_10904);
and U14940 (N_14940,N_9658,N_10287);
and U14941 (N_14941,N_10082,N_9222);
nand U14942 (N_14942,N_10547,N_10674);
nor U14943 (N_14943,N_11234,N_11425);
and U14944 (N_14944,N_10674,N_10670);
nor U14945 (N_14945,N_10066,N_11265);
nand U14946 (N_14946,N_10743,N_9427);
or U14947 (N_14947,N_11709,N_11888);
nand U14948 (N_14948,N_10222,N_10679);
and U14949 (N_14949,N_9293,N_11552);
or U14950 (N_14950,N_11428,N_11817);
or U14951 (N_14951,N_9157,N_11664);
nor U14952 (N_14952,N_11093,N_9533);
nand U14953 (N_14953,N_9083,N_11444);
nor U14954 (N_14954,N_10715,N_9527);
or U14955 (N_14955,N_11811,N_11437);
nor U14956 (N_14956,N_11624,N_10158);
and U14957 (N_14957,N_11457,N_11881);
nand U14958 (N_14958,N_11249,N_10411);
and U14959 (N_14959,N_10789,N_9334);
and U14960 (N_14960,N_10029,N_10374);
and U14961 (N_14961,N_10636,N_9794);
nor U14962 (N_14962,N_9407,N_9432);
and U14963 (N_14963,N_11170,N_10597);
nor U14964 (N_14964,N_11043,N_9692);
nor U14965 (N_14965,N_10255,N_10123);
nor U14966 (N_14966,N_10391,N_10472);
and U14967 (N_14967,N_9782,N_10380);
and U14968 (N_14968,N_11703,N_10495);
or U14969 (N_14969,N_10803,N_11023);
and U14970 (N_14970,N_9700,N_9213);
xor U14971 (N_14971,N_11134,N_10722);
nor U14972 (N_14972,N_11637,N_11395);
nor U14973 (N_14973,N_10620,N_11798);
and U14974 (N_14974,N_9305,N_10648);
nand U14975 (N_14975,N_10739,N_11366);
or U14976 (N_14976,N_10621,N_11535);
nand U14977 (N_14977,N_10084,N_11483);
nor U14978 (N_14978,N_9049,N_10528);
and U14979 (N_14979,N_9129,N_11802);
and U14980 (N_14980,N_11155,N_10367);
nor U14981 (N_14981,N_11504,N_10129);
or U14982 (N_14982,N_10528,N_9397);
nand U14983 (N_14983,N_10655,N_11812);
and U14984 (N_14984,N_11295,N_10076);
nand U14985 (N_14985,N_9141,N_10762);
or U14986 (N_14986,N_9058,N_10518);
nand U14987 (N_14987,N_9678,N_9631);
nor U14988 (N_14988,N_11460,N_11465);
or U14989 (N_14989,N_10893,N_9743);
nand U14990 (N_14990,N_10850,N_10327);
and U14991 (N_14991,N_9780,N_10837);
and U14992 (N_14992,N_10298,N_9577);
and U14993 (N_14993,N_9657,N_11103);
nor U14994 (N_14994,N_9620,N_10467);
or U14995 (N_14995,N_10395,N_11686);
nand U14996 (N_14996,N_9585,N_9827);
and U14997 (N_14997,N_10835,N_11240);
or U14998 (N_14998,N_10190,N_11469);
nor U14999 (N_14999,N_9417,N_11808);
nand UO_0 (O_0,N_12447,N_14826);
nand UO_1 (O_1,N_14741,N_13156);
nand UO_2 (O_2,N_14437,N_14816);
or UO_3 (O_3,N_13966,N_14180);
and UO_4 (O_4,N_12199,N_13237);
or UO_5 (O_5,N_12403,N_12802);
nand UO_6 (O_6,N_13525,N_12218);
or UO_7 (O_7,N_14687,N_14022);
and UO_8 (O_8,N_12937,N_13694);
nor UO_9 (O_9,N_12239,N_14218);
nor UO_10 (O_10,N_14173,N_14755);
or UO_11 (O_11,N_14266,N_12381);
nor UO_12 (O_12,N_12864,N_12269);
and UO_13 (O_13,N_13843,N_14272);
or UO_14 (O_14,N_14518,N_12254);
and UO_15 (O_15,N_14041,N_13984);
and UO_16 (O_16,N_13306,N_13889);
and UO_17 (O_17,N_13832,N_13482);
or UO_18 (O_18,N_14896,N_12703);
or UO_19 (O_19,N_12493,N_12357);
nor UO_20 (O_20,N_13125,N_12607);
and UO_21 (O_21,N_12674,N_12328);
or UO_22 (O_22,N_12073,N_13249);
nor UO_23 (O_23,N_12972,N_13548);
nor UO_24 (O_24,N_14210,N_12927);
nor UO_25 (O_25,N_13019,N_12477);
or UO_26 (O_26,N_12234,N_14724);
nand UO_27 (O_27,N_13483,N_14413);
nand UO_28 (O_28,N_13211,N_13786);
nand UO_29 (O_29,N_12185,N_13908);
nor UO_30 (O_30,N_13437,N_12696);
or UO_31 (O_31,N_12536,N_13754);
or UO_32 (O_32,N_12048,N_14564);
or UO_33 (O_33,N_14791,N_13205);
and UO_34 (O_34,N_12065,N_14350);
nor UO_35 (O_35,N_12443,N_14613);
and UO_36 (O_36,N_12208,N_14371);
or UO_37 (O_37,N_12260,N_12110);
nand UO_38 (O_38,N_14348,N_14986);
nand UO_39 (O_39,N_13982,N_13932);
nand UO_40 (O_40,N_14061,N_13104);
and UO_41 (O_41,N_13815,N_12890);
and UO_42 (O_42,N_14148,N_13480);
or UO_43 (O_43,N_12648,N_13383);
and UO_44 (O_44,N_13481,N_12631);
nand UO_45 (O_45,N_12911,N_13813);
or UO_46 (O_46,N_12406,N_12288);
nand UO_47 (O_47,N_14628,N_12999);
nor UO_48 (O_48,N_12960,N_14404);
and UO_49 (O_49,N_12202,N_12723);
nand UO_50 (O_50,N_14122,N_12826);
nor UO_51 (O_51,N_13496,N_13329);
nor UO_52 (O_52,N_13326,N_12318);
and UO_53 (O_53,N_12622,N_13254);
xor UO_54 (O_54,N_12635,N_14839);
nor UO_55 (O_55,N_13448,N_13102);
and UO_56 (O_56,N_14159,N_13723);
or UO_57 (O_57,N_13484,N_13007);
xor UO_58 (O_58,N_14191,N_12616);
and UO_59 (O_59,N_12554,N_14807);
or UO_60 (O_60,N_12700,N_12259);
and UO_61 (O_61,N_14860,N_12051);
or UO_62 (O_62,N_13705,N_14196);
or UO_63 (O_63,N_12873,N_12418);
nor UO_64 (O_64,N_14994,N_13041);
and UO_65 (O_65,N_14474,N_14060);
and UO_66 (O_66,N_13914,N_12896);
nand UO_67 (O_67,N_12498,N_14871);
nor UO_68 (O_68,N_12919,N_13364);
or UO_69 (O_69,N_13945,N_13658);
or UO_70 (O_70,N_12987,N_14231);
or UO_71 (O_71,N_14009,N_13228);
nor UO_72 (O_72,N_14273,N_14537);
and UO_73 (O_73,N_12738,N_12449);
nor UO_74 (O_74,N_12766,N_13569);
nand UO_75 (O_75,N_14144,N_12128);
and UO_76 (O_76,N_13256,N_14514);
and UO_77 (O_77,N_14566,N_12285);
nand UO_78 (O_78,N_12138,N_13162);
nor UO_79 (O_79,N_14547,N_14677);
nor UO_80 (O_80,N_14252,N_12358);
nor UO_81 (O_81,N_13416,N_12681);
nor UO_82 (O_82,N_13076,N_12124);
and UO_83 (O_83,N_14961,N_12568);
and UO_84 (O_84,N_14658,N_13352);
nor UO_85 (O_85,N_12430,N_14449);
xor UO_86 (O_86,N_14975,N_13467);
nor UO_87 (O_87,N_13030,N_12533);
or UO_88 (O_88,N_12074,N_12215);
and UO_89 (O_89,N_12029,N_14453);
nand UO_90 (O_90,N_14088,N_13736);
nor UO_91 (O_91,N_13108,N_13086);
and UO_92 (O_92,N_12977,N_14419);
nor UO_93 (O_93,N_14854,N_12435);
nor UO_94 (O_94,N_13940,N_14500);
and UO_95 (O_95,N_13682,N_14104);
nor UO_96 (O_96,N_12899,N_14605);
nand UO_97 (O_97,N_12998,N_14722);
or UO_98 (O_98,N_14501,N_12323);
nand UO_99 (O_99,N_13486,N_13857);
or UO_100 (O_100,N_14209,N_13181);
or UO_101 (O_101,N_13021,N_12510);
or UO_102 (O_102,N_12350,N_13426);
nand UO_103 (O_103,N_14825,N_12344);
and UO_104 (O_104,N_12278,N_13113);
nor UO_105 (O_105,N_14053,N_12816);
or UO_106 (O_106,N_14249,N_13592);
or UO_107 (O_107,N_14242,N_12274);
nor UO_108 (O_108,N_14369,N_12803);
and UO_109 (O_109,N_13056,N_12572);
nor UO_110 (O_110,N_14264,N_14351);
nor UO_111 (O_111,N_14539,N_14884);
nor UO_112 (O_112,N_12518,N_13906);
nor UO_113 (O_113,N_14923,N_12419);
or UO_114 (O_114,N_14582,N_12308);
nand UO_115 (O_115,N_13570,N_14590);
nor UO_116 (O_116,N_14407,N_13839);
or UO_117 (O_117,N_13109,N_13728);
nor UO_118 (O_118,N_14044,N_14202);
nand UO_119 (O_119,N_14892,N_12827);
nor UO_120 (O_120,N_12421,N_14377);
nor UO_121 (O_121,N_14666,N_14378);
or UO_122 (O_122,N_13542,N_14522);
nor UO_123 (O_123,N_13866,N_12395);
nand UO_124 (O_124,N_12502,N_14805);
nor UO_125 (O_125,N_14997,N_14320);
or UO_126 (O_126,N_14757,N_12535);
or UO_127 (O_127,N_12428,N_13063);
nand UO_128 (O_128,N_14129,N_13385);
and UO_129 (O_129,N_12321,N_12543);
and UO_130 (O_130,N_14108,N_12106);
or UO_131 (O_131,N_12530,N_14995);
or UO_132 (O_132,N_14817,N_14346);
nand UO_133 (O_133,N_12052,N_13530);
xor UO_134 (O_134,N_12783,N_13847);
or UO_135 (O_135,N_12851,N_12066);
or UO_136 (O_136,N_12653,N_12480);
and UO_137 (O_137,N_14505,N_14705);
nor UO_138 (O_138,N_14296,N_14462);
and UO_139 (O_139,N_13436,N_12086);
nor UO_140 (O_140,N_12769,N_14802);
nand UO_141 (O_141,N_14003,N_12503);
or UO_142 (O_142,N_13663,N_12295);
or UO_143 (O_143,N_13708,N_13586);
and UO_144 (O_144,N_12767,N_14559);
nand UO_145 (O_145,N_13065,N_14420);
nor UO_146 (O_146,N_13495,N_14852);
or UO_147 (O_147,N_12024,N_13639);
xor UO_148 (O_148,N_13500,N_12594);
nand UO_149 (O_149,N_13430,N_13576);
nand UO_150 (O_150,N_13809,N_14103);
nor UO_151 (O_151,N_12817,N_14552);
nor UO_152 (O_152,N_13686,N_14524);
nor UO_153 (O_153,N_13036,N_12404);
nor UO_154 (O_154,N_13291,N_12087);
nor UO_155 (O_155,N_12348,N_14841);
nor UO_156 (O_156,N_13928,N_13829);
nor UO_157 (O_157,N_14806,N_12885);
nand UO_158 (O_158,N_13697,N_12524);
nor UO_159 (O_159,N_12854,N_13774);
or UO_160 (O_160,N_12354,N_13250);
or UO_161 (O_161,N_12279,N_13709);
nand UO_162 (O_162,N_14598,N_12157);
and UO_163 (O_163,N_12845,N_14054);
nand UO_164 (O_164,N_13025,N_12057);
nand UO_165 (O_165,N_14151,N_14592);
nand UO_166 (O_166,N_14957,N_14573);
and UO_167 (O_167,N_12326,N_13078);
nor UO_168 (O_168,N_14908,N_14709);
nor UO_169 (O_169,N_12744,N_13240);
and UO_170 (O_170,N_13931,N_14527);
and UO_171 (O_171,N_14314,N_12242);
nor UO_172 (O_172,N_12601,N_12256);
and UO_173 (O_173,N_14738,N_12169);
nand UO_174 (O_174,N_14714,N_12667);
and UO_175 (O_175,N_13511,N_14255);
and UO_176 (O_176,N_12553,N_13729);
and UO_177 (O_177,N_13018,N_14344);
and UO_178 (O_178,N_12929,N_14930);
or UO_179 (O_179,N_14546,N_12223);
nand UO_180 (O_180,N_13028,N_14747);
nand UO_181 (O_181,N_13376,N_13695);
nor UO_182 (O_182,N_14683,N_12091);
nor UO_183 (O_183,N_14192,N_13775);
nand UO_184 (O_184,N_12356,N_13475);
or UO_185 (O_185,N_13010,N_13219);
and UO_186 (O_186,N_14007,N_13583);
or UO_187 (O_187,N_14693,N_14834);
nand UO_188 (O_188,N_13182,N_13652);
and UO_189 (O_189,N_12808,N_13547);
or UO_190 (O_190,N_13257,N_12232);
or UO_191 (O_191,N_14604,N_12782);
nor UO_192 (O_192,N_13133,N_13630);
and UO_193 (O_193,N_12955,N_12132);
nand UO_194 (O_194,N_13455,N_13360);
nand UO_195 (O_195,N_14058,N_14772);
nor UO_196 (O_196,N_12991,N_14265);
and UO_197 (O_197,N_14890,N_12585);
nand UO_198 (O_198,N_14645,N_12710);
and UO_199 (O_199,N_14018,N_14558);
nor UO_200 (O_200,N_12969,N_12322);
or UO_201 (O_201,N_12345,N_13821);
or UO_202 (O_202,N_14381,N_12470);
nor UO_203 (O_203,N_14118,N_13699);
nor UO_204 (O_204,N_13788,N_14996);
nand UO_205 (O_205,N_14691,N_14864);
and UO_206 (O_206,N_14535,N_14868);
or UO_207 (O_207,N_12108,N_13068);
xor UO_208 (O_208,N_13354,N_14876);
or UO_209 (O_209,N_12819,N_13094);
nand UO_210 (O_210,N_13097,N_14284);
nor UO_211 (O_211,N_14447,N_12033);
nor UO_212 (O_212,N_14328,N_14660);
or UO_213 (O_213,N_13606,N_13804);
nand UO_214 (O_214,N_14780,N_12399);
nand UO_215 (O_215,N_14782,N_12677);
or UO_216 (O_216,N_12486,N_13992);
or UO_217 (O_217,N_13668,N_14595);
nor UO_218 (O_218,N_12003,N_13447);
and UO_219 (O_219,N_13653,N_14245);
or UO_220 (O_220,N_12732,N_13346);
nor UO_221 (O_221,N_12499,N_14033);
nand UO_222 (O_222,N_12591,N_13185);
xor UO_223 (O_223,N_13989,N_12574);
and UO_224 (O_224,N_14149,N_13994);
and UO_225 (O_225,N_14833,N_14174);
nor UO_226 (O_226,N_13335,N_14811);
or UO_227 (O_227,N_12760,N_12483);
or UO_228 (O_228,N_13636,N_12820);
or UO_229 (O_229,N_12016,N_12730);
and UO_230 (O_230,N_12402,N_14386);
nor UO_231 (O_231,N_13521,N_13340);
nor UO_232 (O_232,N_14313,N_12140);
and UO_233 (O_233,N_13252,N_13757);
nand UO_234 (O_234,N_13072,N_13502);
and UO_235 (O_235,N_12335,N_13504);
or UO_236 (O_236,N_12712,N_13136);
or UO_237 (O_237,N_13339,N_13137);
and UO_238 (O_238,N_12595,N_13266);
nand UO_239 (O_239,N_14080,N_14365);
and UO_240 (O_240,N_12832,N_12941);
nand UO_241 (O_241,N_13017,N_12107);
and UO_242 (O_242,N_12975,N_12966);
or UO_243 (O_243,N_12475,N_12456);
nand UO_244 (O_244,N_12867,N_12928);
or UO_245 (O_245,N_14119,N_14197);
xnor UO_246 (O_246,N_13207,N_12726);
and UO_247 (O_247,N_14203,N_12604);
nor UO_248 (O_248,N_13602,N_12784);
nand UO_249 (O_249,N_13357,N_13979);
or UO_250 (O_250,N_14525,N_13292);
and UO_251 (O_251,N_14471,N_12670);
nor UO_252 (O_252,N_12014,N_13465);
nor UO_253 (O_253,N_12233,N_13913);
and UO_254 (O_254,N_13750,N_13564);
nor UO_255 (O_255,N_14797,N_13273);
or UO_256 (O_256,N_14679,N_12482);
and UO_257 (O_257,N_13002,N_12913);
xnor UO_258 (O_258,N_12367,N_12045);
nor UO_259 (O_259,N_13693,N_12944);
xnor UO_260 (O_260,N_14713,N_13559);
or UO_261 (O_261,N_12142,N_13283);
nand UO_262 (O_262,N_13883,N_12935);
or UO_263 (O_263,N_13048,N_12090);
and UO_264 (O_264,N_13118,N_14297);
nand UO_265 (O_265,N_13865,N_14241);
nand UO_266 (O_266,N_14486,N_13196);
and UO_267 (O_267,N_13479,N_12365);
nand UO_268 (O_268,N_14803,N_13373);
and UO_269 (O_269,N_12342,N_12985);
nor UO_270 (O_270,N_14484,N_12838);
nand UO_271 (O_271,N_14176,N_12191);
or UO_272 (O_272,N_12876,N_12139);
and UO_273 (O_273,N_12440,N_13477);
nand UO_274 (O_274,N_13626,N_13791);
and UO_275 (O_275,N_14861,N_14831);
nor UO_276 (O_276,N_14697,N_12325);
and UO_277 (O_277,N_12619,N_14214);
or UO_278 (O_278,N_12165,N_13445);
xnor UO_279 (O_279,N_14682,N_14819);
nor UO_280 (O_280,N_13272,N_14944);
and UO_281 (O_281,N_13314,N_14257);
nand UO_282 (O_282,N_14850,N_13609);
nor UO_283 (O_283,N_13905,N_12303);
xor UO_284 (O_284,N_13515,N_13616);
and UO_285 (O_285,N_14376,N_12789);
and UO_286 (O_286,N_13935,N_14251);
and UO_287 (O_287,N_13080,N_13618);
nor UO_288 (O_288,N_14097,N_14671);
nor UO_289 (O_289,N_13659,N_13006);
nor UO_290 (O_290,N_13440,N_14312);
or UO_291 (O_291,N_13087,N_12579);
or UO_292 (O_292,N_12474,N_14082);
nand UO_293 (O_293,N_14665,N_14828);
and UO_294 (O_294,N_14565,N_13270);
or UO_295 (O_295,N_14795,N_12171);
and UO_296 (O_296,N_14125,N_13566);
nor UO_297 (O_297,N_13154,N_12265);
nand UO_298 (O_298,N_12000,N_12450);
or UO_299 (O_299,N_12801,N_14787);
nor UO_300 (O_300,N_13869,N_14792);
nor UO_301 (O_301,N_14620,N_14062);
and UO_302 (O_302,N_14416,N_13581);
nand UO_303 (O_303,N_13469,N_13789);
and UO_304 (O_304,N_13026,N_13478);
and UO_305 (O_305,N_12753,N_12061);
nand UO_306 (O_306,N_14327,N_12241);
and UO_307 (O_307,N_12981,N_12756);
nor UO_308 (O_308,N_12547,N_12079);
or UO_309 (O_309,N_13785,N_14425);
or UO_310 (O_310,N_13224,N_14382);
and UO_311 (O_311,N_12940,N_14881);
or UO_312 (O_312,N_13735,N_12751);
nor UO_313 (O_313,N_12060,N_12485);
nand UO_314 (O_314,N_13062,N_12668);
or UO_315 (O_315,N_13546,N_12264);
xor UO_316 (O_316,N_13202,N_13749);
and UO_317 (O_317,N_13431,N_13064);
and UO_318 (O_318,N_13886,N_13132);
or UO_319 (O_319,N_12740,N_13999);
and UO_320 (O_320,N_14659,N_14725);
nor UO_321 (O_321,N_12041,N_13929);
nor UO_322 (O_322,N_14409,N_12366);
or UO_323 (O_323,N_12145,N_13424);
nand UO_324 (O_324,N_14719,N_12961);
nand UO_325 (O_325,N_13607,N_13603);
nand UO_326 (O_326,N_14905,N_13055);
nor UO_327 (O_327,N_14135,N_13432);
nor UO_328 (O_328,N_12031,N_12207);
xnor UO_329 (O_329,N_13105,N_13212);
and UO_330 (O_330,N_12620,N_13214);
or UO_331 (O_331,N_12497,N_13040);
and UO_332 (O_332,N_12878,N_13328);
nand UO_333 (O_333,N_12912,N_13834);
and UO_334 (O_334,N_14676,N_13873);
or UO_335 (O_335,N_13733,N_12638);
and UO_336 (O_336,N_14161,N_12022);
nor UO_337 (O_337,N_14601,N_13816);
and UO_338 (O_338,N_13327,N_14672);
or UO_339 (O_339,N_12811,N_14389);
or UO_340 (O_340,N_14095,N_12408);
or UO_341 (O_341,N_13678,N_13554);
nand UO_342 (O_342,N_13150,N_12597);
and UO_343 (O_343,N_14767,N_12204);
and UO_344 (O_344,N_14275,N_12608);
or UO_345 (O_345,N_13389,N_14579);
nand UO_346 (O_346,N_13814,N_14749);
nand UO_347 (O_347,N_12229,N_12646);
and UO_348 (O_348,N_13271,N_12283);
and UO_349 (O_349,N_12695,N_12665);
nand UO_350 (O_350,N_13011,N_12689);
or UO_351 (O_351,N_12180,N_13321);
nor UO_352 (O_352,N_12775,N_13684);
or UO_353 (O_353,N_13580,N_12945);
xnor UO_354 (O_354,N_13926,N_12174);
xnor UO_355 (O_355,N_13493,N_13656);
nor UO_356 (O_356,N_12821,N_12901);
or UO_357 (O_357,N_12167,N_12293);
nor UO_358 (O_358,N_13001,N_13732);
nor UO_359 (O_359,N_13751,N_14387);
nand UO_360 (O_360,N_12385,N_12289);
and UO_361 (O_361,N_14329,N_12096);
nand UO_362 (O_362,N_12075,N_13412);
and UO_363 (O_363,N_12313,N_13704);
nand UO_364 (O_364,N_13806,N_13597);
xnor UO_365 (O_365,N_14158,N_14942);
and UO_366 (O_366,N_14971,N_13474);
or UO_367 (O_367,N_12059,N_13057);
nand UO_368 (O_368,N_13771,N_14434);
or UO_369 (O_369,N_12198,N_14778);
nor UO_370 (O_370,N_13503,N_12752);
nand UO_371 (O_371,N_13146,N_13919);
nor UO_372 (O_372,N_12353,N_14362);
nor UO_373 (O_373,N_14692,N_14271);
xor UO_374 (O_374,N_12586,N_14038);
or UO_375 (O_375,N_12836,N_12237);
nand UO_376 (O_376,N_14359,N_14674);
and UO_377 (O_377,N_12522,N_12950);
nand UO_378 (O_378,N_12649,N_13689);
nand UO_379 (O_379,N_14510,N_13641);
nor UO_380 (O_380,N_13201,N_12825);
or UO_381 (O_381,N_14184,N_14065);
nand UO_382 (O_382,N_13160,N_13836);
nand UO_383 (O_383,N_12210,N_13655);
nand UO_384 (O_384,N_12206,N_13895);
nand UO_385 (O_385,N_13319,N_13574);
or UO_386 (O_386,N_14756,N_13882);
or UO_387 (O_387,N_14017,N_14475);
nor UO_388 (O_388,N_12959,N_14454);
nor UO_389 (O_389,N_14551,N_13022);
or UO_390 (O_390,N_12971,N_14446);
and UO_391 (O_391,N_12800,N_13297);
and UO_392 (O_392,N_14403,N_14305);
xor UO_393 (O_393,N_14987,N_12850);
nor UO_394 (O_394,N_14600,N_14550);
nand UO_395 (O_395,N_13888,N_14642);
nor UO_396 (O_396,N_14761,N_13463);
nor UO_397 (O_397,N_14766,N_12663);
nor UO_398 (O_398,N_14468,N_14762);
nand UO_399 (O_399,N_13174,N_14528);
and UO_400 (O_400,N_12580,N_13631);
and UO_401 (O_401,N_14057,N_12917);
and UO_402 (O_402,N_13520,N_13584);
or UO_403 (O_403,N_12228,N_12815);
and UO_404 (O_404,N_13755,N_13203);
nand UO_405 (O_405,N_13730,N_13288);
nand UO_406 (O_406,N_12077,N_14814);
and UO_407 (O_407,N_14147,N_12220);
nor UO_408 (O_408,N_14696,N_14294);
and UO_409 (O_409,N_14748,N_12954);
nor UO_410 (O_410,N_12887,N_14189);
or UO_411 (O_411,N_12039,N_13911);
nand UO_412 (O_412,N_13544,N_14545);
nor UO_413 (O_413,N_14163,N_14112);
nand UO_414 (O_414,N_14967,N_13965);
and UO_415 (O_415,N_12095,N_14972);
nor UO_416 (O_416,N_14343,N_13260);
nand UO_417 (O_417,N_13739,N_13851);
and UO_418 (O_418,N_13613,N_12355);
or UO_419 (O_419,N_13085,N_12363);
nand UO_420 (O_420,N_13608,N_14623);
nor UO_421 (O_421,N_13023,N_12170);
nand UO_422 (O_422,N_13286,N_14681);
and UO_423 (O_423,N_13782,N_12661);
nand UO_424 (O_424,N_12351,N_14589);
and UO_425 (O_425,N_13512,N_14920);
or UO_426 (O_426,N_14548,N_13582);
and UO_427 (O_427,N_14531,N_13177);
or UO_428 (O_428,N_13949,N_14445);
and UO_429 (O_429,N_14366,N_13805);
nand UO_430 (O_430,N_12694,N_13761);
or UO_431 (O_431,N_12201,N_12478);
nor UO_432 (O_432,N_14504,N_12794);
nor UO_433 (O_433,N_13420,N_14502);
xor UO_434 (O_434,N_13691,N_14012);
xor UO_435 (O_435,N_12371,N_12855);
and UO_436 (O_436,N_13439,N_13334);
nor UO_437 (O_437,N_14542,N_13961);
or UO_438 (O_438,N_13151,N_14624);
or UO_439 (O_439,N_14422,N_12629);
nand UO_440 (O_440,N_12921,N_13187);
or UO_441 (O_441,N_12286,N_12611);
nor UO_442 (O_442,N_14190,N_13054);
nand UO_443 (O_443,N_12405,N_13140);
nand UO_444 (O_444,N_13111,N_14295);
nand UO_445 (O_445,N_13082,N_14100);
or UO_446 (O_446,N_14170,N_13423);
and UO_447 (O_447,N_14578,N_12755);
and UO_448 (O_448,N_13550,N_13714);
nand UO_449 (O_449,N_12225,N_12882);
or UO_450 (O_450,N_14730,N_13959);
nor UO_451 (O_451,N_12588,N_12725);
and UO_452 (O_452,N_12292,N_13290);
or UO_453 (O_453,N_14509,N_13863);
or UO_454 (O_454,N_14110,N_12652);
and UO_455 (O_455,N_12846,N_13666);
or UO_456 (O_456,N_14866,N_13179);
and UO_457 (O_457,N_12644,N_14084);
nand UO_458 (O_458,N_13665,N_13849);
nand UO_459 (O_459,N_13706,N_14048);
and UO_460 (O_460,N_12666,N_12392);
nor UO_461 (O_461,N_13244,N_13685);
or UO_462 (O_462,N_14145,N_13819);
or UO_463 (O_463,N_14947,N_13073);
and UO_464 (O_464,N_12872,N_14974);
or UO_465 (O_465,N_14611,N_12660);
and UO_466 (O_466,N_12227,N_13670);
and UO_467 (O_467,N_14028,N_14261);
and UO_468 (O_468,N_12672,N_12764);
and UO_469 (O_469,N_13858,N_14036);
or UO_470 (O_470,N_14345,N_12250);
and UO_471 (O_471,N_12916,N_14622);
nor UO_472 (O_472,N_13121,N_13936);
and UO_473 (O_473,N_14668,N_13840);
or UO_474 (O_474,N_12496,N_13210);
or UO_475 (O_475,N_14657,N_13059);
nand UO_476 (O_476,N_12545,N_13565);
nor UO_477 (O_477,N_14223,N_14776);
nor UO_478 (O_478,N_12777,N_13139);
and UO_479 (O_479,N_13920,N_13664);
or UO_480 (O_480,N_12517,N_12125);
nand UO_481 (O_481,N_12177,N_14532);
and UO_482 (O_482,N_12531,N_12092);
nor UO_483 (O_483,N_12281,N_13038);
nor UO_484 (O_484,N_12722,N_14759);
nand UO_485 (O_485,N_12748,N_12268);
or UO_486 (O_486,N_14931,N_13822);
nor UO_487 (O_487,N_12182,N_12391);
nor UO_488 (O_488,N_14325,N_12909);
nor UO_489 (O_489,N_14480,N_14310);
or UO_490 (O_490,N_13715,N_12506);
and UO_491 (O_491,N_13841,N_14243);
nand UO_492 (O_492,N_14185,N_14042);
nand UO_493 (O_493,N_13860,N_13088);
or UO_494 (O_494,N_14469,N_14689);
or UO_495 (O_495,N_14254,N_13418);
or UO_496 (O_496,N_14282,N_13830);
and UO_497 (O_497,N_14127,N_13594);
nor UO_498 (O_498,N_14179,N_14740);
or UO_499 (O_499,N_13452,N_12834);
and UO_500 (O_500,N_14763,N_12436);
nor UO_501 (O_501,N_12731,N_14225);
nand UO_502 (O_502,N_12790,N_13912);
xor UO_503 (O_503,N_12297,N_12143);
and UO_504 (O_504,N_13600,N_13368);
and UO_505 (O_505,N_12445,N_12918);
and UO_506 (O_506,N_12032,N_13222);
or UO_507 (O_507,N_12895,N_13589);
and UO_508 (O_508,N_12822,N_13531);
nor UO_509 (O_509,N_14607,N_14347);
nand UO_510 (O_510,N_13300,N_12637);
nor UO_511 (O_511,N_12063,N_13899);
or UO_512 (O_512,N_13324,N_13345);
or UO_513 (O_513,N_12609,N_12527);
nand UO_514 (O_514,N_13248,N_14114);
and UO_515 (O_515,N_13274,N_14970);
or UO_516 (O_516,N_13348,N_13127);
and UO_517 (O_517,N_13000,N_12951);
and UO_518 (O_518,N_12735,N_14609);
or UO_519 (O_519,N_12544,N_12623);
or UO_520 (O_520,N_12979,N_13066);
nor UO_521 (O_521,N_12739,N_12778);
nor UO_522 (O_522,N_12750,N_13438);
or UO_523 (O_523,N_13800,N_13534);
nor UO_524 (O_524,N_14315,N_14300);
nor UO_525 (O_525,N_12127,N_13585);
or UO_526 (O_526,N_12420,N_12394);
and UO_527 (O_527,N_14139,N_12809);
or UO_528 (O_528,N_12411,N_13762);
nor UO_529 (O_529,N_12294,N_12688);
xnor UO_530 (O_530,N_13285,N_13215);
nor UO_531 (O_531,N_12282,N_13386);
or UO_532 (O_532,N_14771,N_13110);
or UO_533 (O_533,N_14796,N_12307);
nand UO_534 (O_534,N_12062,N_12213);
or UO_535 (O_535,N_13753,N_12956);
nor UO_536 (O_536,N_13333,N_13625);
nor UO_537 (O_537,N_13667,N_14555);
or UO_538 (O_538,N_14616,N_12640);
or UO_539 (O_539,N_12072,N_12930);
nand UO_540 (O_540,N_12980,N_12549);
and UO_541 (O_541,N_13529,N_14383);
nor UO_542 (O_542,N_12673,N_12729);
nand UO_543 (O_543,N_13946,N_14517);
or UO_544 (O_544,N_13172,N_14669);
and UO_545 (O_545,N_14652,N_14123);
nand UO_546 (O_546,N_13159,N_12214);
nand UO_547 (O_547,N_13033,N_13363);
nand UO_548 (O_548,N_14259,N_13801);
nand UO_549 (O_549,N_13897,N_14783);
and UO_550 (O_550,N_13462,N_13535);
or UO_551 (O_551,N_14968,N_14293);
nand UO_552 (O_552,N_13269,N_12160);
nand UO_553 (O_553,N_12746,N_14291);
nor UO_554 (O_554,N_14699,N_13131);
or UO_555 (O_555,N_13640,N_14842);
or UO_556 (O_556,N_13081,N_14456);
or UO_557 (O_557,N_12575,N_12617);
or UO_558 (O_558,N_12742,N_13322);
xor UO_559 (O_559,N_14444,N_12134);
and UO_560 (O_560,N_14898,N_14143);
nor UO_561 (O_561,N_13168,N_12627);
nor UO_562 (O_562,N_13862,N_13450);
or UO_563 (O_563,N_14467,N_14770);
nor UO_564 (O_564,N_13323,N_14380);
or UO_565 (O_565,N_12556,N_12634);
and UO_566 (O_566,N_12787,N_14976);
or UO_567 (O_567,N_12953,N_12515);
nor UO_568 (O_568,N_13879,N_14168);
or UO_569 (O_569,N_14508,N_13282);
nor UO_570 (O_570,N_12902,N_13134);
nor UO_571 (O_571,N_12686,N_13122);
nor UO_572 (O_572,N_13939,N_14804);
nor UO_573 (O_573,N_12187,N_12511);
or UO_574 (O_574,N_12231,N_13366);
and UO_575 (O_575,N_14198,N_13461);
or UO_576 (O_576,N_12592,N_14650);
and UO_577 (O_577,N_12409,N_14081);
nand UO_578 (O_578,N_14718,N_13259);
nor UO_579 (O_579,N_13166,N_13925);
nor UO_580 (O_580,N_12571,N_14032);
and UO_581 (O_581,N_12874,N_12333);
nor UO_582 (O_582,N_13696,N_12044);
nand UO_583 (O_583,N_12166,N_13180);
and UO_584 (O_584,N_14673,N_13284);
nor UO_585 (O_585,N_13880,N_14808);
nor UO_586 (O_586,N_12104,N_13231);
nor UO_587 (O_587,N_13232,N_13293);
or UO_588 (O_588,N_14138,N_12757);
nand UO_589 (O_589,N_12563,N_14432);
or UO_590 (O_590,N_14618,N_14907);
nand UO_591 (O_591,N_13004,N_12034);
xor UO_592 (O_592,N_13008,N_13794);
and UO_593 (O_593,N_14980,N_12988);
or UO_594 (O_594,N_12973,N_12119);
nand UO_595 (O_595,N_13765,N_12984);
nor UO_596 (O_596,N_14339,N_14025);
or UO_597 (O_597,N_14865,N_13067);
or UO_598 (O_598,N_12133,N_13119);
nand UO_599 (O_599,N_13361,N_14331);
nand UO_600 (O_600,N_13902,N_12875);
nor UO_601 (O_601,N_14843,N_12932);
xor UO_602 (O_602,N_12249,N_13683);
or UO_603 (O_603,N_14832,N_13831);
and UO_604 (O_604,N_14227,N_13092);
nor UO_605 (O_605,N_13766,N_13473);
or UO_606 (O_606,N_13114,N_12488);
or UO_607 (O_607,N_14670,N_14649);
and UO_608 (O_608,N_14694,N_12512);
or UO_609 (O_609,N_12155,N_12192);
nor UO_610 (O_610,N_14936,N_14979);
or UO_611 (O_611,N_14047,N_12028);
nand UO_612 (O_612,N_14415,N_13674);
nand UO_613 (O_613,N_14274,N_14092);
or UO_614 (O_614,N_12791,N_13220);
and UO_615 (O_615,N_14617,N_14373);
nor UO_616 (O_616,N_14289,N_12219);
and UO_617 (O_617,N_14519,N_12209);
and UO_618 (O_618,N_13165,N_14324);
nor UO_619 (O_619,N_12765,N_12770);
and UO_620 (O_620,N_13987,N_14171);
nand UO_621 (O_621,N_13975,N_12144);
or UO_622 (O_622,N_13112,N_14512);
and UO_623 (O_623,N_13075,N_14793);
or UO_624 (O_624,N_14571,N_14002);
nor UO_625 (O_625,N_14130,N_13826);
or UO_626 (O_626,N_14529,N_13382);
nand UO_627 (O_627,N_13779,N_12632);
or UO_628 (O_628,N_13874,N_12844);
or UO_629 (O_629,N_12338,N_12625);
nor UO_630 (O_630,N_12541,N_13050);
or UO_631 (O_631,N_13891,N_13952);
and UO_632 (O_632,N_13149,N_14914);
and UO_633 (O_633,N_13797,N_12561);
nor UO_634 (O_634,N_13183,N_13144);
and UO_635 (O_635,N_12007,N_14384);
and UO_636 (O_636,N_13690,N_13850);
and UO_637 (O_637,N_14182,N_14809);
nand UO_638 (O_638,N_14030,N_12414);
nor UO_639 (O_639,N_14460,N_13610);
nand UO_640 (O_640,N_13748,N_13317);
nor UO_641 (O_641,N_12718,N_13218);
nand UO_642 (O_642,N_12175,N_14654);
nand UO_643 (O_643,N_14758,N_14101);
and UO_644 (O_644,N_14330,N_13457);
and UO_645 (O_645,N_14094,N_12481);
or UO_646 (O_646,N_14234,N_12939);
and UO_647 (O_647,N_14661,N_14520);
and UO_648 (O_648,N_13304,N_12576);
nor UO_649 (O_649,N_14553,N_14750);
and UO_650 (O_650,N_12070,N_14953);
nand UO_651 (O_651,N_12243,N_13648);
nor UO_652 (O_652,N_12389,N_14363);
or UO_653 (O_653,N_12866,N_14777);
or UO_654 (O_654,N_12733,N_13190);
nor UO_655 (O_655,N_13238,N_13116);
nor UO_656 (O_656,N_14603,N_12763);
nor UO_657 (O_657,N_14268,N_13229);
nand UO_658 (O_658,N_14248,N_13126);
or UO_659 (O_659,N_13350,N_13267);
nor UO_660 (O_660,N_14024,N_12013);
nor UO_661 (O_661,N_14894,N_14924);
nor UO_662 (O_662,N_12793,N_13184);
nand UO_663 (O_663,N_13161,N_14534);
or UO_664 (O_664,N_14169,N_13817);
nor UO_665 (O_665,N_13930,N_12257);
nor UO_666 (O_666,N_14071,N_14016);
nor UO_667 (O_667,N_14880,N_14442);
and UO_668 (O_668,N_14538,N_14496);
nand UO_669 (O_669,N_12799,N_13601);
nor UO_670 (O_670,N_13265,N_12555);
nor UO_671 (O_671,N_14039,N_14423);
and UO_672 (O_672,N_14536,N_14515);
and UO_673 (O_673,N_14862,N_14800);
nor UO_674 (O_674,N_12173,N_14729);
and UO_675 (O_675,N_12396,N_13356);
and UO_676 (O_676,N_12903,N_14647);
and UO_677 (O_677,N_12859,N_14250);
and UO_678 (O_678,N_12675,N_12252);
nor UO_679 (O_679,N_13910,N_14769);
and UO_680 (O_680,N_12329,N_14134);
nor UO_681 (O_681,N_12883,N_12301);
and UO_682 (O_682,N_13178,N_13167);
nand UO_683 (O_683,N_13957,N_12410);
xor UO_684 (O_684,N_13390,N_14483);
or UO_685 (O_685,N_12679,N_14247);
or UO_686 (O_686,N_13338,N_13264);
or UO_687 (O_687,N_14932,N_12830);
and UO_688 (O_688,N_14488,N_14981);
or UO_689 (O_689,N_13342,N_14064);
and UO_690 (O_690,N_14893,N_13428);
nand UO_691 (O_691,N_12603,N_13336);
or UO_692 (O_692,N_14006,N_13391);
nand UO_693 (O_693,N_13741,N_14226);
nand UO_694 (O_694,N_14421,N_14288);
or UO_695 (O_695,N_12501,N_12015);
xor UO_696 (O_696,N_12276,N_12010);
and UO_697 (O_697,N_14013,N_14530);
and UO_698 (O_698,N_13101,N_12030);
xnor UO_699 (O_699,N_14429,N_14165);
nor UO_700 (O_700,N_14606,N_12240);
or UO_701 (O_701,N_12442,N_13612);
nand UO_702 (O_702,N_14956,N_13349);
nand UO_703 (O_703,N_14557,N_12650);
xnor UO_704 (O_704,N_12970,N_12610);
xnor UO_705 (O_705,N_12310,N_14640);
and UO_706 (O_706,N_12476,N_12925);
nor UO_707 (O_707,N_12319,N_13556);
nor UO_708 (O_708,N_14311,N_12390);
and UO_709 (O_709,N_13053,N_12628);
or UO_710 (O_710,N_13387,N_13454);
nor UO_711 (O_711,N_13848,N_12304);
and UO_712 (O_712,N_12255,N_14935);
and UO_713 (O_713,N_12287,N_13216);
and UO_714 (O_714,N_13074,N_14374);
nor UO_715 (O_715,N_12457,N_12818);
or UO_716 (O_716,N_12468,N_13393);
nand UO_717 (O_717,N_14499,N_14260);
nand UO_718 (O_718,N_14457,N_13369);
nor UO_719 (O_719,N_13405,N_13921);
or UO_720 (O_720,N_12871,N_14785);
and UO_721 (O_721,N_14810,N_14233);
and UO_722 (O_722,N_13632,N_14070);
nor UO_723 (O_723,N_14745,N_13494);
nand UO_724 (O_724,N_13106,N_12415);
nand UO_725 (O_725,N_14838,N_12728);
nand UO_726 (O_726,N_14301,N_13927);
or UO_727 (O_727,N_12495,N_13093);
or UO_728 (O_728,N_14258,N_12302);
and UO_729 (O_729,N_12516,N_13646);
nor UO_730 (O_730,N_14736,N_14801);
nor UO_731 (O_731,N_14569,N_13492);
nand UO_732 (O_732,N_14102,N_14925);
nand UO_733 (O_733,N_12835,N_14178);
nor UO_734 (O_734,N_14688,N_13189);
or UO_735 (O_735,N_12100,N_14511);
nor UO_736 (O_736,N_14431,N_12749);
and UO_737 (O_737,N_13835,N_13532);
nor UO_738 (O_738,N_12275,N_12933);
or UO_739 (O_739,N_14615,N_13947);
and UO_740 (O_740,N_14614,N_14723);
and UO_741 (O_741,N_14703,N_13976);
nor UO_742 (O_742,N_14818,N_14391);
or UO_743 (O_743,N_13688,N_14799);
and UO_744 (O_744,N_14298,N_14922);
and UO_745 (O_745,N_12523,N_14938);
or UO_746 (O_746,N_12009,N_14638);
nor UO_747 (O_747,N_12747,N_13415);
nor UO_748 (O_748,N_14193,N_12768);
nor UO_749 (O_749,N_14988,N_12036);
nand UO_750 (O_750,N_12657,N_14340);
xor UO_751 (O_751,N_14636,N_14540);
nor UO_752 (O_752,N_13425,N_13472);
or UO_753 (O_753,N_12936,N_13505);
nand UO_754 (O_754,N_14490,N_14962);
nor UO_755 (O_755,N_12715,N_13411);
or UO_756 (O_756,N_12384,N_12983);
nor UO_757 (O_757,N_12886,N_13384);
nor UO_758 (O_758,N_12828,N_14086);
nand UO_759 (O_759,N_13540,N_14401);
and UO_760 (O_760,N_14280,N_12687);
nor UO_761 (O_761,N_14964,N_13402);
or UO_762 (O_762,N_12567,N_13123);
or UO_763 (O_763,N_14230,N_12655);
and UO_764 (O_764,N_12965,N_12774);
nor UO_765 (O_765,N_13325,N_14717);
or UO_766 (O_766,N_13042,N_14452);
or UO_767 (O_767,N_14302,N_13147);
nand UO_768 (O_768,N_14117,N_14238);
nand UO_769 (O_769,N_14116,N_12606);
or UO_770 (O_770,N_13192,N_13978);
or UO_771 (O_771,N_14989,N_12046);
or UO_772 (O_772,N_13488,N_14367);
or UO_773 (O_773,N_13983,N_13464);
or UO_774 (O_774,N_14211,N_12514);
xnor UO_775 (O_775,N_12131,N_14857);
nor UO_776 (O_776,N_13943,N_13115);
xnor UO_777 (O_777,N_12745,N_12088);
and UO_778 (O_778,N_12339,N_14851);
nand UO_779 (O_779,N_13555,N_13084);
or UO_780 (O_780,N_12184,N_12137);
or UO_781 (O_781,N_14427,N_12692);
nor UO_782 (O_782,N_12716,N_14883);
nor UO_783 (O_783,N_14632,N_14370);
or UO_784 (O_784,N_12413,N_13799);
and UO_785 (O_785,N_12097,N_14106);
nand UO_786 (O_786,N_13365,N_13698);
nor UO_787 (O_787,N_13239,N_12962);
and UO_788 (O_788,N_12719,N_13997);
nand UO_789 (O_789,N_12526,N_12785);
and UO_790 (O_790,N_13032,N_14411);
nor UO_791 (O_791,N_14948,N_12105);
or UO_792 (O_792,N_13128,N_13491);
nor UO_793 (O_793,N_14089,N_14237);
and UO_794 (O_794,N_12761,N_12314);
nand UO_795 (O_795,N_12277,N_12019);
or UO_796 (O_796,N_14891,N_14208);
and UO_797 (O_797,N_13117,N_12978);
and UO_798 (O_798,N_13024,N_13466);
nor UO_799 (O_799,N_14207,N_13990);
nand UO_800 (O_800,N_13209,N_12188);
or UO_801 (O_801,N_13768,N_14728);
nor UO_802 (O_802,N_14882,N_12190);
and UO_803 (O_803,N_13731,N_14352);
nand UO_804 (O_804,N_12025,N_12401);
nor UO_805 (O_805,N_12989,N_13312);
nand UO_806 (O_806,N_14612,N_13676);
or UO_807 (O_807,N_12795,N_13058);
xor UO_808 (O_808,N_12494,N_12893);
or UO_809 (O_809,N_14045,N_12957);
or UO_810 (O_810,N_13120,N_14844);
nor UO_811 (O_811,N_12002,N_14439);
or UO_812 (O_812,N_14879,N_14276);
nand UO_813 (O_813,N_12949,N_13344);
or UO_814 (O_814,N_13513,N_14115);
xnor UO_815 (O_815,N_13864,N_13644);
nand UO_816 (O_816,N_13560,N_14646);
nor UO_817 (O_817,N_14085,N_14859);
nor UO_818 (O_818,N_12071,N_14570);
or UO_819 (O_819,N_13468,N_13811);
or UO_820 (O_820,N_13876,N_14966);
nand UO_821 (O_821,N_13725,N_12263);
and UO_822 (O_822,N_13517,N_12361);
or UO_823 (O_823,N_14043,N_13577);
nor UO_824 (O_824,N_12709,N_14031);
or UO_825 (O_825,N_12425,N_12397);
and UO_826 (O_826,N_14653,N_13379);
or UO_827 (O_827,N_14175,N_14835);
nor UO_828 (O_828,N_13015,N_13974);
nor UO_829 (O_829,N_13784,N_14909);
nand UO_830 (O_830,N_14317,N_12315);
nor UO_831 (O_831,N_12186,N_12439);
nor UO_832 (O_832,N_12519,N_14754);
nor UO_833 (O_833,N_13654,N_13718);
nor UO_834 (O_834,N_12656,N_12720);
nand UO_835 (O_835,N_13635,N_14361);
or UO_836 (O_836,N_13924,N_14464);
nand UO_837 (O_837,N_14629,N_12235);
nor UO_838 (O_838,N_13510,N_13200);
nor UO_839 (O_839,N_12842,N_13650);
nand UO_840 (O_840,N_13394,N_12807);
nor UO_841 (O_841,N_14385,N_13221);
and UO_842 (O_842,N_14132,N_13153);
nor UO_843 (O_843,N_14829,N_12779);
and UO_844 (O_844,N_12441,N_13318);
nand UO_845 (O_845,N_13770,N_13489);
nor UO_846 (O_846,N_12711,N_13868);
or UO_847 (O_847,N_14212,N_14440);
and UO_848 (O_848,N_14959,N_13294);
nor UO_849 (O_849,N_12372,N_12343);
nor UO_850 (O_850,N_13487,N_13295);
and UO_851 (O_851,N_12189,N_14120);
and UO_852 (O_852,N_12327,N_13892);
nand UO_853 (O_853,N_13687,N_14109);
nor UO_854 (O_854,N_12161,N_12267);
nor UO_855 (O_855,N_12159,N_14008);
and UO_856 (O_856,N_13634,N_12316);
and UO_857 (O_857,N_14393,N_13241);
or UO_858 (O_858,N_14586,N_12550);
or UO_859 (O_859,N_14588,N_12566);
or UO_860 (O_860,N_14217,N_12993);
nor UO_861 (O_861,N_13545,N_13643);
and UO_862 (O_862,N_14029,N_14753);
xnor UO_863 (O_863,N_12528,N_12490);
nand UO_864 (O_864,N_13152,N_14798);
nand UO_865 (O_865,N_13406,N_12639);
nand UO_866 (O_866,N_13173,N_13679);
xnor UO_867 (O_867,N_12837,N_13549);
and UO_868 (O_868,N_13713,N_13760);
nand UO_869 (O_869,N_12111,N_12008);
nand UO_870 (O_870,N_13281,N_12798);
and UO_871 (O_871,N_14583,N_13158);
nand UO_872 (O_872,N_12004,N_14662);
and UO_873 (O_873,N_14399,N_13710);
and UO_874 (O_874,N_12922,N_12814);
or UO_875 (O_875,N_12261,N_14985);
or UO_876 (O_876,N_14973,N_12172);
and UO_877 (O_877,N_12271,N_12658);
or UO_878 (O_878,N_12432,N_14414);
xor UO_879 (O_879,N_12152,N_13476);
and UO_880 (O_880,N_13717,N_13591);
nand UO_881 (O_881,N_13395,N_12362);
nor UO_882 (O_882,N_12236,N_14395);
and UO_883 (O_883,N_12069,N_13009);
nand UO_884 (O_884,N_13701,N_14358);
or UO_885 (O_885,N_12312,N_14568);
nor UO_886 (O_886,N_12853,N_13341);
and UO_887 (O_887,N_13079,N_14544);
nor UO_888 (O_888,N_12135,N_12596);
nor UO_889 (O_889,N_12680,N_13901);
or UO_890 (O_890,N_14476,N_12245);
nor UO_891 (O_891,N_14641,N_12573);
nand UO_892 (O_892,N_13875,N_12986);
nand UO_893 (O_893,N_13337,N_14656);
or UO_894 (O_894,N_14812,N_13037);
nand UO_895 (O_895,N_14267,N_12934);
nand UO_896 (O_896,N_12915,N_14052);
or UO_897 (O_897,N_12452,N_13098);
or UO_898 (O_898,N_13796,N_14136);
or UO_899 (O_899,N_12453,N_13523);
and UO_900 (O_900,N_14774,N_12460);
nand UO_901 (O_901,N_14091,N_13619);
or UO_902 (O_902,N_13499,N_14887);
nor UO_903 (O_903,N_12534,N_14010);
nor UO_904 (O_904,N_12099,N_13343);
or UO_905 (O_905,N_14308,N_12713);
nor UO_906 (O_906,N_13590,N_14702);
nor UO_907 (O_907,N_13579,N_13621);
or UO_908 (O_908,N_13253,N_12708);
or UO_909 (O_909,N_14379,N_14737);
nor UO_910 (O_910,N_12183,N_12920);
or UO_911 (O_911,N_14911,N_14215);
or UO_912 (O_912,N_12221,N_14716);
or UO_913 (O_913,N_12772,N_13628);
nor UO_914 (O_914,N_12103,N_13245);
or UO_915 (O_915,N_12026,N_13567);
and UO_916 (O_916,N_12889,N_14364);
and UO_917 (O_917,N_12331,N_12997);
or UO_918 (O_918,N_12539,N_14937);
xor UO_919 (O_919,N_14172,N_14394);
or UO_920 (O_920,N_14067,N_13671);
nand UO_921 (O_921,N_12334,N_14072);
nor UO_922 (O_922,N_14141,N_12148);
xor UO_923 (O_923,N_12868,N_14066);
nand UO_924 (O_924,N_14577,N_14263);
or UO_925 (O_925,N_12847,N_14392);
or UO_926 (O_926,N_13627,N_14406);
and UO_927 (O_927,N_14200,N_12162);
or UO_928 (O_928,N_12848,N_13922);
nor UO_929 (O_929,N_13596,N_12806);
nand UO_930 (O_930,N_13091,N_13193);
and UO_931 (O_931,N_12863,N_13027);
nand UO_932 (O_932,N_14549,N_14927);
nand UO_933 (O_933,N_14201,N_12317);
nor UO_934 (O_934,N_13163,N_13853);
and UO_935 (O_935,N_13971,N_13915);
and UO_936 (O_936,N_12179,N_14873);
and UO_937 (O_937,N_14786,N_12704);
xor UO_938 (O_938,N_14478,N_14461);
and UO_939 (O_939,N_14035,N_13890);
nand UO_940 (O_940,N_14820,N_13528);
nand UO_941 (O_941,N_12011,N_12964);
nor UO_942 (O_942,N_14098,N_13649);
nand UO_943 (O_943,N_12862,N_13331);
nand UO_944 (O_944,N_12701,N_12147);
nor UO_945 (O_945,N_13962,N_14481);
nand UO_946 (O_946,N_13918,N_12224);
nand UO_947 (O_947,N_14644,N_14593);
and UO_948 (O_948,N_13988,N_14999);
xor UO_949 (O_949,N_12727,N_13509);
and UO_950 (O_950,N_13164,N_14885);
nor UO_951 (O_951,N_12852,N_12565);
or UO_952 (O_952,N_13916,N_13661);
nor UO_953 (O_953,N_12958,N_14704);
and UO_954 (O_954,N_13355,N_12849);
or UO_955 (O_955,N_12685,N_14051);
nor UO_956 (O_956,N_14602,N_14794);
nand UO_957 (O_957,N_14633,N_14224);
nor UO_958 (O_958,N_12266,N_13719);
nor UO_959 (O_959,N_12337,N_12116);
and UO_960 (O_960,N_12678,N_14355);
nor UO_961 (O_961,N_12058,N_13881);
nand UO_962 (O_962,N_12296,N_13722);
nor UO_963 (O_963,N_13005,N_12370);
or UO_964 (O_964,N_14027,N_13870);
or UO_965 (O_965,N_13599,N_13727);
and UO_966 (O_966,N_13884,N_13854);
nand UO_967 (O_967,N_13737,N_14680);
or UO_968 (O_968,N_13934,N_14913);
nor UO_969 (O_969,N_14026,N_12636);
nand UO_970 (O_970,N_12898,N_13280);
or UO_971 (O_971,N_14847,N_13370);
or UO_972 (O_972,N_14727,N_14575);
nor UO_973 (O_973,N_14710,N_12758);
or UO_974 (O_974,N_13604,N_12558);
and UO_975 (O_975,N_14715,N_14059);
nand UO_976 (O_976,N_14846,N_13740);
or UO_977 (O_977,N_13519,N_13060);
and UO_978 (O_978,N_13996,N_13490);
and UO_979 (O_979,N_12352,N_13401);
and UO_980 (O_980,N_12569,N_13933);
nand UO_981 (O_981,N_12856,N_14398);
nand UO_982 (O_982,N_13107,N_14195);
nand UO_983 (O_983,N_13793,N_14240);
or UO_984 (O_984,N_14836,N_13501);
nor UO_985 (O_985,N_14845,N_12926);
and UO_986 (O_986,N_14899,N_14943);
and UO_987 (O_987,N_12910,N_12943);
and UO_988 (O_988,N_12469,N_14368);
or UO_989 (O_989,N_13396,N_12247);
or UO_990 (O_990,N_12491,N_14167);
or UO_991 (O_991,N_14146,N_14643);
nand UO_992 (O_992,N_14576,N_12195);
nor UO_993 (O_993,N_13968,N_14760);
or UO_994 (O_994,N_12130,N_12464);
nor UO_995 (O_995,N_13077,N_13307);
or UO_996 (O_996,N_14430,N_14342);
nor UO_997 (O_997,N_12299,N_14412);
and UO_998 (O_998,N_14152,N_12341);
nor UO_999 (O_999,N_13278,N_12076);
and UO_1000 (O_1000,N_12599,N_12114);
and UO_1001 (O_1001,N_13377,N_14895);
nor UO_1002 (O_1002,N_14983,N_14246);
nand UO_1003 (O_1003,N_12582,N_14400);
nand UO_1004 (O_1004,N_13651,N_14270);
nand UO_1005 (O_1005,N_14277,N_14111);
xor UO_1006 (O_1006,N_14941,N_14177);
or UO_1007 (O_1007,N_14034,N_13867);
xnor UO_1008 (O_1008,N_12992,N_14698);
and UO_1009 (O_1009,N_14939,N_12248);
and UO_1010 (O_1010,N_14773,N_12164);
nand UO_1011 (O_1011,N_13362,N_12551);
nor UO_1012 (O_1012,N_12613,N_13980);
nand UO_1013 (O_1013,N_13378,N_13453);
xor UO_1014 (O_1014,N_14443,N_14194);
nor UO_1015 (O_1015,N_12176,N_14853);
and UO_1016 (O_1016,N_13204,N_13673);
nor UO_1017 (O_1017,N_14784,N_14487);
and UO_1018 (O_1018,N_14822,N_13313);
or UO_1019 (O_1019,N_14965,N_12976);
and UO_1020 (O_1020,N_13985,N_14133);
and UO_1021 (O_1021,N_13157,N_12129);
and UO_1022 (O_1022,N_13287,N_14919);
nor UO_1023 (O_1023,N_12444,N_13507);
nor UO_1024 (O_1024,N_12829,N_14685);
and UO_1025 (O_1025,N_12387,N_12451);
or UO_1026 (O_1026,N_12373,N_14397);
or UO_1027 (O_1027,N_13404,N_14077);
nand UO_1028 (O_1028,N_14993,N_12654);
or UO_1029 (O_1029,N_13958,N_13807);
and UO_1030 (O_1030,N_13443,N_12270);
or UO_1031 (O_1031,N_14513,N_14562);
and UO_1032 (O_1032,N_13170,N_13427);
or UO_1033 (O_1033,N_14594,N_14858);
or UO_1034 (O_1034,N_13142,N_13944);
nand UO_1035 (O_1035,N_14228,N_13186);
or UO_1036 (O_1036,N_14655,N_14912);
nand UO_1037 (O_1037,N_13742,N_13444);
nor UO_1038 (O_1038,N_14353,N_13572);
and UO_1039 (O_1039,N_13941,N_12805);
nand UO_1040 (O_1040,N_13029,N_12300);
or UO_1041 (O_1041,N_12860,N_13417);
nor UO_1042 (O_1042,N_12948,N_14867);
nand UO_1043 (O_1043,N_12120,N_12178);
and UO_1044 (O_1044,N_14764,N_14162);
or UO_1045 (O_1045,N_12446,N_12484);
nor UO_1046 (O_1046,N_12717,N_12141);
nand UO_1047 (O_1047,N_12118,N_14470);
and UO_1048 (O_1048,N_12967,N_13846);
and UO_1049 (O_1049,N_14503,N_13562);
nor UO_1050 (O_1050,N_12841,N_13838);
or UO_1051 (O_1051,N_13738,N_12386);
nand UO_1052 (O_1052,N_12364,N_12346);
or UO_1053 (O_1053,N_14954,N_13514);
nand UO_1054 (O_1054,N_13279,N_12870);
nor UO_1055 (O_1055,N_13518,N_12455);
or UO_1056 (O_1056,N_12067,N_13135);
nand UO_1057 (O_1057,N_14587,N_14150);
nand UO_1058 (O_1058,N_12924,N_12982);
or UO_1059 (O_1059,N_12309,N_13726);
nand UO_1060 (O_1060,N_14824,N_13798);
or UO_1061 (O_1061,N_12043,N_12047);
or UO_1062 (O_1062,N_12946,N_12005);
and UO_1063 (O_1063,N_13070,N_12633);
nand UO_1064 (O_1064,N_13090,N_13963);
or UO_1065 (O_1065,N_13330,N_13043);
or UO_1066 (O_1066,N_12126,N_14417);
or UO_1067 (O_1067,N_12466,N_13571);
nor UO_1068 (O_1068,N_13148,N_13459);
nor UO_1069 (O_1069,N_14621,N_14627);
nand UO_1070 (O_1070,N_14285,N_14648);
and UO_1071 (O_1071,N_12080,N_12858);
nand UO_1072 (O_1072,N_12542,N_14049);
or UO_1073 (O_1073,N_13764,N_13275);
nor UO_1074 (O_1074,N_12564,N_14619);
or UO_1075 (O_1075,N_13553,N_14900);
and UO_1076 (O_1076,N_13442,N_14338);
or UO_1077 (O_1077,N_12473,N_12330);
and UO_1078 (O_1078,N_12881,N_12509);
or UO_1079 (O_1079,N_12538,N_13552);
and UO_1080 (O_1080,N_14743,N_13230);
or UO_1081 (O_1081,N_12557,N_12900);
or UO_1082 (O_1082,N_12904,N_13894);
xnor UO_1083 (O_1083,N_13543,N_14073);
and UO_1084 (O_1084,N_13171,N_13497);
and UO_1085 (O_1085,N_13243,N_13624);
nor UO_1086 (O_1086,N_14541,N_14585);
nand UO_1087 (O_1087,N_13711,N_14482);
or UO_1088 (O_1088,N_14307,N_12379);
or UO_1089 (O_1089,N_12796,N_14186);
or UO_1090 (O_1090,N_14262,N_12194);
or UO_1091 (O_1091,N_13069,N_13937);
nor UO_1092 (O_1092,N_14695,N_13460);
nand UO_1093 (O_1093,N_14521,N_12626);
and UO_1094 (O_1094,N_14000,N_13226);
nand UO_1095 (O_1095,N_12947,N_14341);
nor UO_1096 (O_1096,N_12089,N_12865);
or UO_1097 (O_1097,N_13539,N_13233);
nand UO_1098 (O_1098,N_13449,N_12651);
or UO_1099 (O_1099,N_14303,N_14886);
or UO_1100 (O_1100,N_12884,N_14744);
nor UO_1101 (O_1101,N_12068,N_12552);
xnor UO_1102 (O_1102,N_12181,N_12492);
nor UO_1103 (O_1103,N_13044,N_13103);
nand UO_1104 (O_1104,N_13358,N_12578);
or UO_1105 (O_1105,N_12122,N_12149);
and UO_1106 (O_1106,N_12690,N_14978);
xor UO_1107 (O_1107,N_12532,N_13967);
and UO_1108 (O_1108,N_13506,N_12306);
and UO_1109 (O_1109,N_12336,N_14405);
nand UO_1110 (O_1110,N_12388,N_13955);
and UO_1111 (O_1111,N_13593,N_12605);
nor UO_1112 (O_1112,N_14963,N_12479);
and UO_1113 (O_1113,N_13538,N_14933);
nor UO_1114 (O_1114,N_13485,N_13446);
nor UO_1115 (O_1115,N_14731,N_14639);
xor UO_1116 (O_1116,N_13398,N_14849);
or UO_1117 (O_1117,N_13611,N_12205);
and UO_1118 (O_1118,N_14137,N_12598);
xor UO_1119 (O_1119,N_13422,N_12050);
nor UO_1120 (O_1120,N_13712,N_12743);
xnor UO_1121 (O_1121,N_13720,N_12272);
and UO_1122 (O_1122,N_14121,N_12431);
nand UO_1123 (O_1123,N_14156,N_14283);
nor UO_1124 (O_1124,N_14751,N_12618);
nand UO_1125 (O_1125,N_14625,N_14219);
nand UO_1126 (O_1126,N_12593,N_14458);
nand UO_1127 (O_1127,N_12458,N_14635);
nor UO_1128 (O_1128,N_13223,N_13953);
nand UO_1129 (O_1129,N_14984,N_13262);
nand UO_1130 (O_1130,N_14788,N_13498);
or UO_1131 (O_1131,N_13622,N_13777);
or UO_1132 (O_1132,N_12724,N_14436);
nor UO_1133 (O_1133,N_12702,N_14004);
nand UO_1134 (O_1134,N_12839,N_12200);
and UO_1135 (O_1135,N_13012,N_12952);
xor UO_1136 (O_1136,N_13268,N_12647);
nand UO_1137 (O_1137,N_14472,N_13311);
nand UO_1138 (O_1138,N_14929,N_13247);
and UO_1139 (O_1139,N_14848,N_13578);
xor UO_1140 (O_1140,N_13917,N_12513);
or UO_1141 (O_1141,N_14450,N_13700);
nor UO_1142 (O_1142,N_12426,N_13844);
nor UO_1143 (O_1143,N_13995,N_14584);
or UO_1144 (O_1144,N_14337,N_14005);
and UO_1145 (O_1145,N_13991,N_14244);
nand UO_1146 (O_1146,N_13938,N_14388);
nand UO_1147 (O_1147,N_13964,N_13434);
or UO_1148 (O_1148,N_12877,N_13175);
or UO_1149 (O_1149,N_13537,N_14187);
xnor UO_1150 (O_1150,N_14402,N_13758);
and UO_1151 (O_1151,N_12320,N_13408);
nor UO_1152 (O_1152,N_13802,N_13470);
and UO_1153 (O_1153,N_14078,N_12676);
and UO_1154 (O_1154,N_13145,N_13969);
and UO_1155 (O_1155,N_12520,N_13020);
nand UO_1156 (O_1156,N_13772,N_14543);
or UO_1157 (O_1157,N_12762,N_13660);
and UO_1158 (O_1158,N_12581,N_12376);
nand UO_1159 (O_1159,N_13143,N_13587);
nor UO_1160 (O_1160,N_14982,N_14459);
nor UO_1161 (O_1161,N_14815,N_12448);
or UO_1162 (O_1162,N_12888,N_13034);
nor UO_1163 (O_1163,N_14675,N_13217);
nand UO_1164 (O_1164,N_14732,N_14827);
and UO_1165 (O_1165,N_12662,N_14128);
or UO_1166 (O_1166,N_13255,N_13195);
and UO_1167 (O_1167,N_13429,N_13138);
nand UO_1168 (O_1168,N_13769,N_14426);
or UO_1169 (O_1169,N_14372,N_14046);
nand UO_1170 (O_1170,N_13605,N_14926);
or UO_1171 (O_1171,N_14229,N_14563);
or UO_1172 (O_1172,N_14733,N_12707);
or UO_1173 (O_1173,N_13970,N_14055);
and UO_1174 (O_1174,N_14142,N_14591);
and UO_1175 (O_1175,N_14477,N_12153);
and UO_1176 (O_1176,N_12006,N_12151);
and UO_1177 (O_1177,N_13551,N_14916);
nor UO_1178 (O_1178,N_14952,N_12471);
nand UO_1179 (O_1179,N_12504,N_13598);
or UO_1180 (O_1180,N_14286,N_13234);
nand UO_1181 (O_1181,N_12963,N_12880);
or UO_1182 (O_1182,N_13263,N_13208);
and UO_1183 (O_1183,N_14126,N_14019);
or UO_1184 (O_1184,N_14667,N_12253);
and UO_1185 (O_1185,N_12056,N_14256);
nand UO_1186 (O_1186,N_14023,N_12102);
and UO_1187 (O_1187,N_12905,N_14915);
nor UO_1188 (O_1188,N_14183,N_12546);
and UO_1189 (O_1189,N_13441,N_12021);
nand UO_1190 (O_1190,N_13993,N_12771);
and UO_1191 (O_1191,N_13855,N_12369);
or UO_1192 (O_1192,N_13923,N_13763);
or UO_1193 (O_1193,N_13129,N_13071);
nand UO_1194 (O_1194,N_13095,N_14079);
and UO_1195 (O_1195,N_13051,N_13898);
or UO_1196 (O_1196,N_14533,N_14056);
or UO_1197 (O_1197,N_12094,N_13818);
or UO_1198 (O_1198,N_12222,N_13013);
nor UO_1199 (O_1199,N_14507,N_13845);
or UO_1200 (O_1200,N_13031,N_14489);
and UO_1201 (O_1201,N_12291,N_12570);
or UO_1202 (O_1202,N_13657,N_13629);
and UO_1203 (O_1203,N_14199,N_14014);
nor UO_1204 (O_1204,N_12781,N_12508);
nand UO_1205 (O_1205,N_14768,N_14707);
or UO_1206 (O_1206,N_13315,N_13795);
nand UO_1207 (O_1207,N_14205,N_13227);
nand UO_1208 (O_1208,N_14360,N_12869);
and UO_1209 (O_1209,N_13878,N_13909);
nand UO_1210 (O_1210,N_12562,N_14498);
nor UO_1211 (O_1211,N_13856,N_14040);
nand UO_1212 (O_1212,N_12461,N_14424);
and UO_1213 (O_1213,N_12642,N_14626);
and UO_1214 (O_1214,N_13124,N_13332);
nand UO_1215 (O_1215,N_14479,N_13199);
nand UO_1216 (O_1216,N_14099,N_12136);
or UO_1217 (O_1217,N_13046,N_12230);
or UO_1218 (O_1218,N_12083,N_12085);
nor UO_1219 (O_1219,N_13298,N_14869);
nor UO_1220 (O_1220,N_14506,N_12600);
nor UO_1221 (O_1221,N_12671,N_14068);
and UO_1222 (O_1222,N_12923,N_12968);
nor UO_1223 (O_1223,N_14290,N_13558);
nor UO_1224 (O_1224,N_14991,N_12683);
or UO_1225 (O_1225,N_14323,N_12525);
nor UO_1226 (O_1226,N_12892,N_12560);
or UO_1227 (O_1227,N_14155,N_13563);
nand UO_1228 (O_1228,N_14789,N_14318);
or UO_1229 (O_1229,N_12810,N_13824);
or UO_1230 (O_1230,N_13588,N_12559);
or UO_1231 (O_1231,N_12459,N_12630);
nor UO_1232 (O_1232,N_12156,N_13303);
or UO_1233 (O_1233,N_13302,N_13956);
and UO_1234 (O_1234,N_14154,N_13451);
nor UO_1235 (O_1235,N_12374,N_12383);
nor UO_1236 (O_1236,N_13397,N_13724);
nor UO_1237 (O_1237,N_12251,N_13526);
nand UO_1238 (O_1238,N_14433,N_14428);
nand UO_1239 (O_1239,N_14074,N_13756);
nor UO_1240 (O_1240,N_12012,N_14928);
xnor UO_1241 (O_1241,N_12462,N_13374);
nand UO_1242 (O_1242,N_14711,N_14204);
nor UO_1243 (O_1243,N_12427,N_14813);
nand UO_1244 (O_1244,N_13827,N_14181);
nor UO_1245 (O_1245,N_13852,N_12375);
nor UO_1246 (O_1246,N_14775,N_13261);
nand UO_1247 (O_1247,N_12759,N_12023);
nand UO_1248 (O_1248,N_12037,N_12537);
and UO_1249 (O_1249,N_14221,N_13251);
or UO_1250 (O_1250,N_13637,N_13301);
and UO_1251 (O_1251,N_13310,N_13568);
nand UO_1252 (O_1252,N_13213,N_13872);
or UO_1253 (O_1253,N_14950,N_12691);
and UO_1254 (O_1254,N_13308,N_13900);
nand UO_1255 (O_1255,N_12017,N_13808);
nor UO_1256 (O_1256,N_14686,N_12664);
nand UO_1257 (O_1257,N_14904,N_14441);
nor UO_1258 (O_1258,N_12737,N_14096);
or UO_1259 (O_1259,N_14917,N_14701);
nor UO_1260 (O_1260,N_13825,N_13014);
nor UO_1261 (O_1261,N_14945,N_12054);
and UO_1262 (O_1262,N_14269,N_12831);
and UO_1263 (O_1263,N_14610,N_13960);
nor UO_1264 (O_1264,N_13877,N_14526);
xnor UO_1265 (O_1265,N_12990,N_13954);
or UO_1266 (O_1266,N_14299,N_13052);
nand UO_1267 (O_1267,N_12705,N_12773);
nor UO_1268 (O_1268,N_13372,N_14581);
and UO_1269 (O_1269,N_14561,N_14069);
and UO_1270 (O_1270,N_12463,N_12942);
nor UO_1271 (O_1271,N_12714,N_14306);
or UO_1272 (O_1272,N_14556,N_13703);
nor UO_1273 (O_1273,N_13100,N_12669);
nand UO_1274 (O_1274,N_13977,N_12380);
and UO_1275 (O_1275,N_14874,N_12212);
or UO_1276 (O_1276,N_12055,N_12018);
nand UO_1277 (O_1277,N_12398,N_14678);
or UO_1278 (O_1278,N_13096,N_13887);
or UO_1279 (O_1279,N_14332,N_12529);
xnor UO_1280 (O_1280,N_12340,N_12879);
xor UO_1281 (O_1281,N_12641,N_12377);
nand UO_1282 (O_1282,N_13623,N_12049);
xnor UO_1283 (O_1283,N_14608,N_14349);
nor UO_1284 (O_1284,N_14213,N_14903);
or UO_1285 (O_1285,N_13400,N_12123);
and UO_1286 (O_1286,N_14951,N_13188);
and UO_1287 (O_1287,N_12038,N_12472);
or UO_1288 (O_1288,N_12040,N_13859);
and UO_1289 (O_1289,N_14877,N_14572);
nand UO_1290 (O_1290,N_12280,N_12273);
nand UO_1291 (O_1291,N_14083,N_12053);
or UO_1292 (O_1292,N_13638,N_12093);
nor UO_1293 (O_1293,N_12698,N_13536);
or UO_1294 (O_1294,N_14336,N_14700);
or UO_1295 (O_1295,N_12994,N_14708);
nor UO_1296 (O_1296,N_12693,N_13615);
and UO_1297 (O_1297,N_14220,N_14969);
or UO_1298 (O_1298,N_14408,N_13861);
nand UO_1299 (O_1299,N_13236,N_12500);
nand UO_1300 (O_1300,N_12163,N_14721);
nor UO_1301 (O_1301,N_13045,N_13003);
and UO_1302 (O_1302,N_13516,N_13647);
nor UO_1303 (O_1303,N_14902,N_13998);
or UO_1304 (O_1304,N_13235,N_14015);
or UO_1305 (O_1305,N_12382,N_13780);
nor UO_1306 (O_1306,N_12001,N_12489);
and UO_1307 (O_1307,N_12507,N_12840);
nand UO_1308 (O_1308,N_13409,N_12305);
or UO_1309 (O_1309,N_13633,N_12699);
or UO_1310 (O_1310,N_14304,N_13541);
and UO_1311 (O_1311,N_14823,N_13614);
nand UO_1312 (O_1312,N_12645,N_14222);
or UO_1313 (O_1313,N_13299,N_14235);
nor UO_1314 (O_1314,N_14921,N_13783);
and UO_1315 (O_1315,N_14087,N_13981);
nand UO_1316 (O_1316,N_12454,N_14206);
or UO_1317 (O_1317,N_13620,N_14076);
nand UO_1318 (O_1318,N_12368,N_14494);
nor UO_1319 (O_1319,N_13745,N_14466);
and UO_1320 (O_1320,N_13399,N_13743);
nand UO_1321 (O_1321,N_13595,N_13803);
or UO_1322 (O_1322,N_13508,N_14232);
nand UO_1323 (O_1323,N_12590,N_13225);
and UO_1324 (O_1324,N_12906,N_12891);
and UO_1325 (O_1325,N_14567,N_12521);
and UO_1326 (O_1326,N_14870,N_14790);
or UO_1327 (O_1327,N_12246,N_13367);
or UO_1328 (O_1328,N_12721,N_14491);
nor UO_1329 (O_1329,N_12078,N_14837);
nand UO_1330 (O_1330,N_12938,N_13375);
nand UO_1331 (O_1331,N_14493,N_14020);
or UO_1332 (O_1332,N_14279,N_14316);
or UO_1333 (O_1333,N_13242,N_13787);
nand UO_1334 (O_1334,N_12158,N_12824);
nor UO_1335 (O_1335,N_12914,N_14375);
and UO_1336 (O_1336,N_13258,N_14292);
or UO_1337 (O_1337,N_14906,N_12833);
nand UO_1338 (O_1338,N_13309,N_14830);
nor UO_1339 (O_1339,N_12027,N_12823);
or UO_1340 (O_1340,N_14897,N_13810);
and UO_1341 (O_1341,N_13130,N_12196);
and UO_1342 (O_1342,N_13885,N_12262);
nor UO_1343 (O_1343,N_13823,N_13904);
or UO_1344 (O_1344,N_14554,N_14321);
nand UO_1345 (O_1345,N_14960,N_13561);
nor UO_1346 (O_1346,N_12324,N_12203);
and UO_1347 (O_1347,N_14495,N_13388);
or UO_1348 (O_1348,N_13677,N_14664);
nand UO_1349 (O_1349,N_13681,N_14560);
and UO_1350 (O_1350,N_12684,N_12035);
nor UO_1351 (O_1351,N_12417,N_13435);
xnor UO_1352 (O_1352,N_13276,N_13410);
and UO_1353 (O_1353,N_12897,N_14418);
or UO_1354 (O_1354,N_14574,N_13575);
or UO_1355 (O_1355,N_13792,N_13524);
or UO_1356 (O_1356,N_14901,N_12754);
or UO_1357 (O_1357,N_14597,N_13744);
nand UO_1358 (O_1358,N_14990,N_14021);
nor UO_1359 (O_1359,N_13296,N_13197);
nand UO_1360 (O_1360,N_14746,N_12115);
nor UO_1361 (O_1361,N_13702,N_12084);
and UO_1362 (O_1362,N_13747,N_13573);
or UO_1363 (O_1363,N_14734,N_12101);
nand UO_1364 (O_1364,N_13016,N_14356);
or UO_1365 (O_1365,N_14451,N_12615);
or UO_1366 (O_1366,N_12736,N_13986);
nor UO_1367 (O_1367,N_14742,N_12995);
or UO_1368 (O_1368,N_12706,N_12780);
and UO_1369 (O_1369,N_14166,N_12117);
nor UO_1370 (O_1370,N_14630,N_14958);
nand UO_1371 (O_1371,N_12424,N_12393);
or UO_1372 (O_1372,N_14319,N_14281);
or UO_1373 (O_1373,N_13456,N_14821);
nor UO_1374 (O_1374,N_14435,N_14438);
nand UO_1375 (O_1375,N_14878,N_12861);
and UO_1376 (O_1376,N_12416,N_14140);
xnor UO_1377 (O_1377,N_13061,N_12487);
and UO_1378 (O_1378,N_14463,N_14236);
or UO_1379 (O_1379,N_14309,N_12797);
nor UO_1380 (O_1380,N_13471,N_12857);
or UO_1381 (O_1381,N_14781,N_12433);
or UO_1382 (O_1382,N_14335,N_14497);
or UO_1383 (O_1383,N_13669,N_14523);
or UO_1384 (O_1384,N_12020,N_12907);
nand UO_1385 (O_1385,N_14977,N_14596);
nand UO_1386 (O_1386,N_13392,N_13662);
or UO_1387 (O_1387,N_12741,N_12682);
nor UO_1388 (O_1388,N_13721,N_13790);
and UO_1389 (O_1389,N_13951,N_14354);
xor UO_1390 (O_1390,N_12621,N_13305);
nor UO_1391 (O_1391,N_12776,N_14287);
nand UO_1392 (O_1392,N_12788,N_12587);
nand UO_1393 (O_1393,N_13320,N_13039);
nand UO_1394 (O_1394,N_12359,N_14157);
nor UO_1395 (O_1395,N_13907,N_14910);
nor UO_1396 (O_1396,N_12412,N_14863);
nand UO_1397 (O_1397,N_14334,N_12284);
xnor UO_1398 (O_1398,N_13371,N_12423);
and UO_1399 (O_1399,N_13421,N_14113);
or UO_1400 (O_1400,N_13533,N_13734);
nand UO_1401 (O_1401,N_13089,N_13833);
nor UO_1402 (O_1402,N_14690,N_12548);
nor UO_1403 (O_1403,N_12589,N_14516);
nand UO_1404 (O_1404,N_14465,N_13380);
nor UO_1405 (O_1405,N_14333,N_12974);
nand UO_1406 (O_1406,N_14188,N_13527);
and UO_1407 (O_1407,N_12238,N_14946);
nor UO_1408 (O_1408,N_12813,N_13141);
nand UO_1409 (O_1409,N_14107,N_14779);
or UO_1410 (O_1410,N_13557,N_12812);
or UO_1411 (O_1411,N_14949,N_14726);
nor UO_1412 (O_1412,N_13812,N_14160);
nor UO_1413 (O_1413,N_12211,N_13716);
and UO_1414 (O_1414,N_13680,N_14357);
nand UO_1415 (O_1415,N_13896,N_14706);
or UO_1416 (O_1416,N_14888,N_13973);
nor UO_1417 (O_1417,N_13419,N_12349);
and UO_1418 (O_1418,N_14410,N_14131);
and UO_1419 (O_1419,N_14239,N_13194);
nor UO_1420 (O_1420,N_12146,N_12290);
and UO_1421 (O_1421,N_13828,N_13169);
nand UO_1422 (O_1422,N_13359,N_14631);
nand UO_1423 (O_1423,N_14875,N_14955);
xnor UO_1424 (O_1424,N_12583,N_14992);
and UO_1425 (O_1425,N_12154,N_14684);
nand UO_1426 (O_1426,N_12311,N_12429);
nor UO_1427 (O_1427,N_13767,N_14855);
nand UO_1428 (O_1428,N_13820,N_12217);
nor UO_1429 (O_1429,N_12197,N_13871);
and UO_1430 (O_1430,N_14001,N_14216);
nor UO_1431 (O_1431,N_12804,N_14037);
nor UO_1432 (O_1432,N_14396,N_13642);
nor UO_1433 (O_1433,N_12614,N_13414);
or UO_1434 (O_1434,N_12438,N_12407);
nor UO_1435 (O_1435,N_13155,N_14663);
nand UO_1436 (O_1436,N_13707,N_12109);
and UO_1437 (O_1437,N_14253,N_13692);
and UO_1438 (O_1438,N_13759,N_13781);
nor UO_1439 (O_1439,N_13351,N_13645);
nor UO_1440 (O_1440,N_14063,N_12540);
or UO_1441 (O_1441,N_13837,N_14326);
or UO_1442 (O_1442,N_13893,N_12467);
nor UO_1443 (O_1443,N_13972,N_13776);
nor UO_1444 (O_1444,N_13316,N_12422);
and UO_1445 (O_1445,N_12400,N_14164);
nand UO_1446 (O_1446,N_14153,N_12244);
xor UO_1447 (O_1447,N_13403,N_14390);
nand UO_1448 (O_1448,N_13950,N_14840);
nand UO_1449 (O_1449,N_13099,N_13522);
or UO_1450 (O_1450,N_12996,N_14322);
and UO_1451 (O_1451,N_13752,N_12226);
nand UO_1452 (O_1452,N_13381,N_13347);
nor UO_1453 (O_1453,N_12360,N_14448);
or UO_1454 (O_1454,N_13353,N_12193);
or UO_1455 (O_1455,N_13206,N_12612);
nand UO_1456 (O_1456,N_14934,N_12113);
nor UO_1457 (O_1457,N_12931,N_12216);
nor UO_1458 (O_1458,N_12792,N_14278);
xnor UO_1459 (O_1459,N_14599,N_13176);
nand UO_1460 (O_1460,N_14739,N_13413);
nor UO_1461 (O_1461,N_13903,N_13458);
and UO_1462 (O_1462,N_13198,N_13083);
or UO_1463 (O_1463,N_12894,N_12843);
and UO_1464 (O_1464,N_13035,N_13746);
nand UO_1465 (O_1465,N_12734,N_12786);
or UO_1466 (O_1466,N_14637,N_12437);
and UO_1467 (O_1467,N_12602,N_12908);
and UO_1468 (O_1468,N_12258,N_13773);
nand UO_1469 (O_1469,N_13842,N_14090);
nor UO_1470 (O_1470,N_14918,N_13433);
and UO_1471 (O_1471,N_14889,N_14752);
or UO_1472 (O_1472,N_12378,N_14720);
nand UO_1473 (O_1473,N_14998,N_12150);
nor UO_1474 (O_1474,N_12121,N_12064);
or UO_1475 (O_1475,N_14940,N_14093);
nand UO_1476 (O_1476,N_14050,N_14455);
nand UO_1477 (O_1477,N_12465,N_12505);
nor UO_1478 (O_1478,N_13191,N_13942);
nand UO_1479 (O_1479,N_12112,N_12697);
nand UO_1480 (O_1480,N_12643,N_12577);
or UO_1481 (O_1481,N_12659,N_13675);
nor UO_1482 (O_1482,N_13778,N_12081);
and UO_1483 (O_1483,N_12042,N_14075);
nand UO_1484 (O_1484,N_13246,N_13289);
and UO_1485 (O_1485,N_12347,N_13407);
and UO_1486 (O_1486,N_13277,N_14124);
and UO_1487 (O_1487,N_14856,N_14492);
nand UO_1488 (O_1488,N_12624,N_14580);
xnor UO_1489 (O_1489,N_12082,N_14011);
nor UO_1490 (O_1490,N_14712,N_13948);
and UO_1491 (O_1491,N_14872,N_13617);
and UO_1492 (O_1492,N_12332,N_14634);
nor UO_1493 (O_1493,N_14105,N_14735);
or UO_1494 (O_1494,N_14651,N_13672);
and UO_1495 (O_1495,N_14765,N_13047);
nor UO_1496 (O_1496,N_12584,N_12434);
nor UO_1497 (O_1497,N_14485,N_12298);
or UO_1498 (O_1498,N_12168,N_14473);
nand UO_1499 (O_1499,N_12098,N_13049);
or UO_1500 (O_1500,N_13510,N_12875);
and UO_1501 (O_1501,N_13573,N_13917);
or UO_1502 (O_1502,N_13338,N_13630);
and UO_1503 (O_1503,N_13132,N_13713);
or UO_1504 (O_1504,N_13342,N_12851);
or UO_1505 (O_1505,N_12896,N_13740);
nor UO_1506 (O_1506,N_12648,N_13767);
and UO_1507 (O_1507,N_13906,N_14856);
and UO_1508 (O_1508,N_13476,N_13871);
nand UO_1509 (O_1509,N_13958,N_12425);
nor UO_1510 (O_1510,N_14380,N_13592);
nor UO_1511 (O_1511,N_12966,N_13316);
nor UO_1512 (O_1512,N_13363,N_12385);
nand UO_1513 (O_1513,N_12942,N_13154);
nand UO_1514 (O_1514,N_14958,N_12824);
or UO_1515 (O_1515,N_12243,N_13490);
and UO_1516 (O_1516,N_13316,N_14506);
nand UO_1517 (O_1517,N_13203,N_13440);
or UO_1518 (O_1518,N_12339,N_12617);
nor UO_1519 (O_1519,N_14716,N_14465);
nand UO_1520 (O_1520,N_14325,N_13117);
and UO_1521 (O_1521,N_13918,N_12972);
and UO_1522 (O_1522,N_14130,N_14687);
or UO_1523 (O_1523,N_13898,N_13213);
nor UO_1524 (O_1524,N_13392,N_14965);
nor UO_1525 (O_1525,N_14476,N_12677);
or UO_1526 (O_1526,N_13609,N_13328);
nor UO_1527 (O_1527,N_14619,N_12445);
and UO_1528 (O_1528,N_14498,N_12813);
or UO_1529 (O_1529,N_13431,N_12017);
nor UO_1530 (O_1530,N_12927,N_14865);
nand UO_1531 (O_1531,N_13428,N_12491);
nand UO_1532 (O_1532,N_12491,N_14526);
nor UO_1533 (O_1533,N_13481,N_12251);
nor UO_1534 (O_1534,N_14212,N_14607);
nand UO_1535 (O_1535,N_13848,N_14961);
and UO_1536 (O_1536,N_13655,N_13430);
nor UO_1537 (O_1537,N_12437,N_12285);
and UO_1538 (O_1538,N_12944,N_12374);
or UO_1539 (O_1539,N_13333,N_14220);
and UO_1540 (O_1540,N_12008,N_14119);
nor UO_1541 (O_1541,N_14061,N_14766);
or UO_1542 (O_1542,N_13219,N_14309);
or UO_1543 (O_1543,N_12616,N_12319);
nand UO_1544 (O_1544,N_12327,N_14401);
nand UO_1545 (O_1545,N_12069,N_13334);
and UO_1546 (O_1546,N_13223,N_12033);
or UO_1547 (O_1547,N_12382,N_14639);
nand UO_1548 (O_1548,N_12489,N_12633);
nand UO_1549 (O_1549,N_13543,N_12049);
or UO_1550 (O_1550,N_12127,N_14313);
or UO_1551 (O_1551,N_12575,N_14372);
and UO_1552 (O_1552,N_14934,N_13610);
or UO_1553 (O_1553,N_14129,N_12094);
nand UO_1554 (O_1554,N_14645,N_13969);
or UO_1555 (O_1555,N_13352,N_13278);
nor UO_1556 (O_1556,N_12422,N_12003);
nor UO_1557 (O_1557,N_14499,N_14854);
or UO_1558 (O_1558,N_14094,N_13763);
nand UO_1559 (O_1559,N_13494,N_13535);
and UO_1560 (O_1560,N_14350,N_12967);
nand UO_1561 (O_1561,N_13747,N_13168);
and UO_1562 (O_1562,N_12972,N_14672);
nor UO_1563 (O_1563,N_12089,N_12054);
nor UO_1564 (O_1564,N_12569,N_13027);
nand UO_1565 (O_1565,N_14402,N_12579);
or UO_1566 (O_1566,N_12926,N_12657);
nor UO_1567 (O_1567,N_14275,N_13336);
nand UO_1568 (O_1568,N_13834,N_12180);
nor UO_1569 (O_1569,N_12871,N_14746);
and UO_1570 (O_1570,N_13760,N_14264);
and UO_1571 (O_1571,N_14161,N_13553);
and UO_1572 (O_1572,N_12835,N_14353);
and UO_1573 (O_1573,N_12774,N_13473);
or UO_1574 (O_1574,N_14827,N_14370);
nand UO_1575 (O_1575,N_13963,N_14187);
nand UO_1576 (O_1576,N_13743,N_14295);
or UO_1577 (O_1577,N_14818,N_14591);
nor UO_1578 (O_1578,N_14231,N_12894);
or UO_1579 (O_1579,N_13363,N_13885);
or UO_1580 (O_1580,N_12260,N_14414);
and UO_1581 (O_1581,N_14045,N_14092);
nand UO_1582 (O_1582,N_13952,N_13775);
nand UO_1583 (O_1583,N_12282,N_12586);
nor UO_1584 (O_1584,N_14053,N_14283);
and UO_1585 (O_1585,N_14122,N_14897);
nand UO_1586 (O_1586,N_12875,N_12429);
nor UO_1587 (O_1587,N_14772,N_14152);
nand UO_1588 (O_1588,N_13109,N_12332);
or UO_1589 (O_1589,N_12301,N_12976);
and UO_1590 (O_1590,N_13706,N_12709);
nand UO_1591 (O_1591,N_14484,N_12720);
and UO_1592 (O_1592,N_14776,N_14972);
nor UO_1593 (O_1593,N_14613,N_14588);
and UO_1594 (O_1594,N_14414,N_12293);
and UO_1595 (O_1595,N_12426,N_13757);
nor UO_1596 (O_1596,N_12527,N_13302);
or UO_1597 (O_1597,N_12403,N_12837);
nor UO_1598 (O_1598,N_14416,N_12695);
nand UO_1599 (O_1599,N_14289,N_13595);
xor UO_1600 (O_1600,N_14883,N_13629);
nand UO_1601 (O_1601,N_14689,N_13175);
xor UO_1602 (O_1602,N_12242,N_13898);
nor UO_1603 (O_1603,N_12450,N_14711);
or UO_1604 (O_1604,N_12605,N_13785);
and UO_1605 (O_1605,N_14465,N_12101);
nor UO_1606 (O_1606,N_13903,N_13457);
and UO_1607 (O_1607,N_12322,N_14671);
nor UO_1608 (O_1608,N_13206,N_12479);
nor UO_1609 (O_1609,N_13436,N_13550);
and UO_1610 (O_1610,N_13184,N_13480);
nand UO_1611 (O_1611,N_13693,N_12383);
or UO_1612 (O_1612,N_14994,N_14172);
nor UO_1613 (O_1613,N_12336,N_13276);
xnor UO_1614 (O_1614,N_14655,N_12279);
or UO_1615 (O_1615,N_13794,N_13221);
and UO_1616 (O_1616,N_13908,N_13870);
nor UO_1617 (O_1617,N_13816,N_13745);
nor UO_1618 (O_1618,N_13357,N_13293);
nand UO_1619 (O_1619,N_12853,N_12266);
or UO_1620 (O_1620,N_12978,N_12615);
or UO_1621 (O_1621,N_13807,N_12710);
nand UO_1622 (O_1622,N_13833,N_13042);
and UO_1623 (O_1623,N_12570,N_12568);
nor UO_1624 (O_1624,N_12063,N_14154);
or UO_1625 (O_1625,N_12505,N_14291);
or UO_1626 (O_1626,N_13198,N_12401);
nor UO_1627 (O_1627,N_14683,N_14376);
xor UO_1628 (O_1628,N_12926,N_14044);
nand UO_1629 (O_1629,N_14096,N_12324);
nand UO_1630 (O_1630,N_14025,N_13655);
nor UO_1631 (O_1631,N_13641,N_12395);
and UO_1632 (O_1632,N_13416,N_13767);
nor UO_1633 (O_1633,N_12744,N_12956);
or UO_1634 (O_1634,N_14423,N_13324);
or UO_1635 (O_1635,N_13504,N_14366);
and UO_1636 (O_1636,N_13615,N_13855);
or UO_1637 (O_1637,N_12571,N_12628);
nand UO_1638 (O_1638,N_12321,N_14457);
or UO_1639 (O_1639,N_13510,N_13576);
nand UO_1640 (O_1640,N_13334,N_13090);
and UO_1641 (O_1641,N_14290,N_14213);
nand UO_1642 (O_1642,N_12522,N_12567);
or UO_1643 (O_1643,N_12500,N_13008);
nor UO_1644 (O_1644,N_12586,N_12286);
nand UO_1645 (O_1645,N_13122,N_14774);
and UO_1646 (O_1646,N_14523,N_14854);
nand UO_1647 (O_1647,N_14327,N_14348);
nor UO_1648 (O_1648,N_14655,N_14102);
nor UO_1649 (O_1649,N_14077,N_12653);
and UO_1650 (O_1650,N_13580,N_12717);
and UO_1651 (O_1651,N_12731,N_14945);
nor UO_1652 (O_1652,N_13269,N_13762);
and UO_1653 (O_1653,N_12926,N_14771);
xnor UO_1654 (O_1654,N_14316,N_13470);
and UO_1655 (O_1655,N_13143,N_12220);
nand UO_1656 (O_1656,N_13481,N_12629);
nor UO_1657 (O_1657,N_13863,N_13992);
nor UO_1658 (O_1658,N_13478,N_12804);
or UO_1659 (O_1659,N_14979,N_12617);
nor UO_1660 (O_1660,N_12334,N_12142);
nor UO_1661 (O_1661,N_13478,N_12960);
or UO_1662 (O_1662,N_13050,N_13622);
nor UO_1663 (O_1663,N_13031,N_12848);
nand UO_1664 (O_1664,N_12236,N_12831);
and UO_1665 (O_1665,N_14370,N_12108);
nor UO_1666 (O_1666,N_14339,N_13279);
nor UO_1667 (O_1667,N_14453,N_12671);
xor UO_1668 (O_1668,N_13846,N_13932);
nor UO_1669 (O_1669,N_14735,N_13225);
nor UO_1670 (O_1670,N_14726,N_13404);
or UO_1671 (O_1671,N_13701,N_13618);
nand UO_1672 (O_1672,N_14613,N_14985);
or UO_1673 (O_1673,N_12407,N_13110);
and UO_1674 (O_1674,N_13552,N_13852);
and UO_1675 (O_1675,N_12838,N_14292);
or UO_1676 (O_1676,N_12708,N_12244);
and UO_1677 (O_1677,N_13431,N_13736);
nor UO_1678 (O_1678,N_13784,N_14834);
nand UO_1679 (O_1679,N_14724,N_14340);
nand UO_1680 (O_1680,N_14780,N_14448);
and UO_1681 (O_1681,N_14859,N_12591);
and UO_1682 (O_1682,N_14698,N_14795);
or UO_1683 (O_1683,N_12163,N_14047);
and UO_1684 (O_1684,N_13181,N_12225);
or UO_1685 (O_1685,N_12334,N_12416);
and UO_1686 (O_1686,N_12855,N_13415);
and UO_1687 (O_1687,N_12268,N_12299);
nor UO_1688 (O_1688,N_12180,N_14081);
xor UO_1689 (O_1689,N_12178,N_12654);
and UO_1690 (O_1690,N_13169,N_12990);
and UO_1691 (O_1691,N_13447,N_12276);
nand UO_1692 (O_1692,N_14975,N_13732);
and UO_1693 (O_1693,N_14925,N_12609);
and UO_1694 (O_1694,N_12892,N_14714);
nand UO_1695 (O_1695,N_12104,N_14308);
nand UO_1696 (O_1696,N_13008,N_14709);
or UO_1697 (O_1697,N_12994,N_14742);
nor UO_1698 (O_1698,N_13362,N_14972);
nand UO_1699 (O_1699,N_12615,N_12968);
or UO_1700 (O_1700,N_14502,N_13484);
and UO_1701 (O_1701,N_13851,N_12813);
and UO_1702 (O_1702,N_13729,N_12087);
or UO_1703 (O_1703,N_13435,N_14956);
xor UO_1704 (O_1704,N_13156,N_12730);
and UO_1705 (O_1705,N_13288,N_14931);
nor UO_1706 (O_1706,N_14928,N_12248);
nor UO_1707 (O_1707,N_14482,N_12698);
and UO_1708 (O_1708,N_12206,N_14330);
or UO_1709 (O_1709,N_14739,N_13851);
nand UO_1710 (O_1710,N_13506,N_14349);
or UO_1711 (O_1711,N_12049,N_13337);
nand UO_1712 (O_1712,N_13886,N_12129);
and UO_1713 (O_1713,N_12466,N_14128);
or UO_1714 (O_1714,N_13115,N_13228);
or UO_1715 (O_1715,N_12553,N_14513);
nor UO_1716 (O_1716,N_14355,N_14993);
nand UO_1717 (O_1717,N_14147,N_14933);
nand UO_1718 (O_1718,N_12789,N_14797);
or UO_1719 (O_1719,N_14475,N_14831);
or UO_1720 (O_1720,N_12741,N_12067);
or UO_1721 (O_1721,N_14225,N_12922);
and UO_1722 (O_1722,N_14099,N_12343);
nor UO_1723 (O_1723,N_14871,N_13196);
and UO_1724 (O_1724,N_12229,N_14333);
nand UO_1725 (O_1725,N_13947,N_14977);
or UO_1726 (O_1726,N_12490,N_13720);
or UO_1727 (O_1727,N_14522,N_12055);
nor UO_1728 (O_1728,N_12986,N_13311);
nand UO_1729 (O_1729,N_13283,N_12961);
nor UO_1730 (O_1730,N_13099,N_14462);
nor UO_1731 (O_1731,N_13466,N_14145);
nor UO_1732 (O_1732,N_12591,N_13269);
nor UO_1733 (O_1733,N_12671,N_12921);
nand UO_1734 (O_1734,N_12292,N_12789);
and UO_1735 (O_1735,N_13480,N_13044);
nor UO_1736 (O_1736,N_12798,N_12485);
nand UO_1737 (O_1737,N_14334,N_12467);
and UO_1738 (O_1738,N_12524,N_13137);
nand UO_1739 (O_1739,N_12324,N_13037);
nand UO_1740 (O_1740,N_14127,N_12821);
or UO_1741 (O_1741,N_13591,N_12167);
or UO_1742 (O_1742,N_12143,N_13419);
nand UO_1743 (O_1743,N_14814,N_13460);
nor UO_1744 (O_1744,N_14139,N_13978);
and UO_1745 (O_1745,N_14031,N_12569);
nand UO_1746 (O_1746,N_14557,N_12580);
or UO_1747 (O_1747,N_14213,N_14168);
or UO_1748 (O_1748,N_14667,N_14792);
and UO_1749 (O_1749,N_14358,N_14906);
and UO_1750 (O_1750,N_14645,N_12547);
nor UO_1751 (O_1751,N_14011,N_14453);
nand UO_1752 (O_1752,N_12856,N_14782);
or UO_1753 (O_1753,N_13552,N_14039);
nor UO_1754 (O_1754,N_13041,N_12551);
nor UO_1755 (O_1755,N_14894,N_13060);
and UO_1756 (O_1756,N_12370,N_12857);
and UO_1757 (O_1757,N_13304,N_13957);
nand UO_1758 (O_1758,N_12080,N_14624);
and UO_1759 (O_1759,N_13569,N_12216);
and UO_1760 (O_1760,N_13473,N_13262);
nor UO_1761 (O_1761,N_14161,N_13578);
or UO_1762 (O_1762,N_14973,N_14490);
nand UO_1763 (O_1763,N_12827,N_12230);
or UO_1764 (O_1764,N_12080,N_13652);
nand UO_1765 (O_1765,N_13274,N_14704);
or UO_1766 (O_1766,N_14215,N_12156);
nand UO_1767 (O_1767,N_12534,N_14168);
and UO_1768 (O_1768,N_13181,N_12775);
and UO_1769 (O_1769,N_12450,N_14269);
nand UO_1770 (O_1770,N_12644,N_13754);
nand UO_1771 (O_1771,N_14997,N_14487);
nand UO_1772 (O_1772,N_12057,N_13690);
and UO_1773 (O_1773,N_14930,N_13582);
nor UO_1774 (O_1774,N_14951,N_13829);
nand UO_1775 (O_1775,N_13682,N_12287);
nand UO_1776 (O_1776,N_14867,N_12386);
nor UO_1777 (O_1777,N_13237,N_12541);
and UO_1778 (O_1778,N_13961,N_12529);
nor UO_1779 (O_1779,N_14711,N_12582);
nor UO_1780 (O_1780,N_12504,N_14246);
nor UO_1781 (O_1781,N_12085,N_14202);
and UO_1782 (O_1782,N_12287,N_14692);
and UO_1783 (O_1783,N_12629,N_12309);
nor UO_1784 (O_1784,N_14177,N_12739);
and UO_1785 (O_1785,N_12705,N_13030);
nand UO_1786 (O_1786,N_14277,N_13670);
nor UO_1787 (O_1787,N_12403,N_14214);
nand UO_1788 (O_1788,N_13326,N_14264);
and UO_1789 (O_1789,N_13043,N_13024);
and UO_1790 (O_1790,N_14570,N_14394);
nand UO_1791 (O_1791,N_14980,N_12193);
nand UO_1792 (O_1792,N_14162,N_12501);
and UO_1793 (O_1793,N_14468,N_12525);
and UO_1794 (O_1794,N_13971,N_14888);
nand UO_1795 (O_1795,N_13748,N_13117);
nor UO_1796 (O_1796,N_13306,N_13618);
and UO_1797 (O_1797,N_12163,N_13919);
and UO_1798 (O_1798,N_13013,N_13719);
nor UO_1799 (O_1799,N_14881,N_12910);
xnor UO_1800 (O_1800,N_13291,N_14092);
or UO_1801 (O_1801,N_13106,N_12153);
or UO_1802 (O_1802,N_13701,N_14986);
and UO_1803 (O_1803,N_13733,N_12773);
nor UO_1804 (O_1804,N_12995,N_13623);
or UO_1805 (O_1805,N_12754,N_13929);
nor UO_1806 (O_1806,N_14355,N_13178);
or UO_1807 (O_1807,N_14586,N_12370);
and UO_1808 (O_1808,N_14276,N_12391);
nor UO_1809 (O_1809,N_14854,N_13550);
and UO_1810 (O_1810,N_13509,N_14775);
and UO_1811 (O_1811,N_13031,N_14076);
and UO_1812 (O_1812,N_12058,N_13499);
and UO_1813 (O_1813,N_14555,N_14449);
nor UO_1814 (O_1814,N_12576,N_14739);
nand UO_1815 (O_1815,N_13049,N_14805);
or UO_1816 (O_1816,N_14010,N_14809);
nand UO_1817 (O_1817,N_14945,N_12275);
and UO_1818 (O_1818,N_13076,N_12459);
and UO_1819 (O_1819,N_14380,N_14804);
nand UO_1820 (O_1820,N_14070,N_12165);
or UO_1821 (O_1821,N_14346,N_14903);
nor UO_1822 (O_1822,N_12137,N_13746);
and UO_1823 (O_1823,N_14888,N_13481);
nor UO_1824 (O_1824,N_13568,N_14433);
or UO_1825 (O_1825,N_13998,N_12120);
nor UO_1826 (O_1826,N_14946,N_13944);
nor UO_1827 (O_1827,N_14849,N_12914);
nor UO_1828 (O_1828,N_12824,N_12755);
and UO_1829 (O_1829,N_14096,N_14047);
nor UO_1830 (O_1830,N_13442,N_12402);
nor UO_1831 (O_1831,N_14729,N_12114);
nand UO_1832 (O_1832,N_14685,N_13732);
or UO_1833 (O_1833,N_12508,N_14648);
and UO_1834 (O_1834,N_12821,N_13079);
nand UO_1835 (O_1835,N_12999,N_14169);
xnor UO_1836 (O_1836,N_12273,N_12461);
nor UO_1837 (O_1837,N_12644,N_12865);
or UO_1838 (O_1838,N_14587,N_12844);
nor UO_1839 (O_1839,N_14810,N_12363);
nor UO_1840 (O_1840,N_13202,N_12452);
or UO_1841 (O_1841,N_14573,N_14224);
nor UO_1842 (O_1842,N_13779,N_14548);
or UO_1843 (O_1843,N_13728,N_14982);
and UO_1844 (O_1844,N_12600,N_12795);
xor UO_1845 (O_1845,N_12171,N_13797);
nor UO_1846 (O_1846,N_13544,N_14992);
nor UO_1847 (O_1847,N_12082,N_12494);
and UO_1848 (O_1848,N_14798,N_12144);
xor UO_1849 (O_1849,N_12435,N_13785);
nor UO_1850 (O_1850,N_14832,N_13652);
or UO_1851 (O_1851,N_14190,N_12087);
nor UO_1852 (O_1852,N_13340,N_12116);
nand UO_1853 (O_1853,N_13190,N_12470);
nor UO_1854 (O_1854,N_12951,N_12616);
and UO_1855 (O_1855,N_12869,N_12459);
nor UO_1856 (O_1856,N_13326,N_14280);
and UO_1857 (O_1857,N_14374,N_13885);
nand UO_1858 (O_1858,N_14616,N_14395);
and UO_1859 (O_1859,N_14937,N_12018);
nand UO_1860 (O_1860,N_13999,N_14708);
and UO_1861 (O_1861,N_12103,N_13654);
and UO_1862 (O_1862,N_12955,N_12423);
nand UO_1863 (O_1863,N_12200,N_12941);
nand UO_1864 (O_1864,N_13930,N_13201);
nand UO_1865 (O_1865,N_12418,N_14086);
nor UO_1866 (O_1866,N_14338,N_12826);
nor UO_1867 (O_1867,N_14854,N_14789);
or UO_1868 (O_1868,N_14098,N_13361);
nor UO_1869 (O_1869,N_14097,N_13637);
nand UO_1870 (O_1870,N_13114,N_12660);
or UO_1871 (O_1871,N_14804,N_14539);
nor UO_1872 (O_1872,N_13560,N_12873);
or UO_1873 (O_1873,N_13307,N_14446);
or UO_1874 (O_1874,N_13598,N_14445);
or UO_1875 (O_1875,N_12930,N_13349);
or UO_1876 (O_1876,N_12284,N_13070);
nand UO_1877 (O_1877,N_13049,N_13627);
and UO_1878 (O_1878,N_13566,N_13546);
and UO_1879 (O_1879,N_12138,N_13014);
and UO_1880 (O_1880,N_13179,N_13037);
and UO_1881 (O_1881,N_14686,N_13176);
or UO_1882 (O_1882,N_13669,N_13684);
and UO_1883 (O_1883,N_13794,N_12115);
nor UO_1884 (O_1884,N_13652,N_14476);
xor UO_1885 (O_1885,N_13337,N_13385);
or UO_1886 (O_1886,N_12468,N_13708);
nor UO_1887 (O_1887,N_14719,N_14859);
or UO_1888 (O_1888,N_12106,N_12983);
and UO_1889 (O_1889,N_14503,N_13791);
nor UO_1890 (O_1890,N_14622,N_13196);
nor UO_1891 (O_1891,N_13383,N_14116);
nor UO_1892 (O_1892,N_13868,N_13841);
and UO_1893 (O_1893,N_12522,N_14200);
xor UO_1894 (O_1894,N_13924,N_13329);
and UO_1895 (O_1895,N_12770,N_13631);
nand UO_1896 (O_1896,N_12705,N_13757);
or UO_1897 (O_1897,N_14932,N_12287);
nor UO_1898 (O_1898,N_13149,N_12853);
and UO_1899 (O_1899,N_12353,N_14666);
nor UO_1900 (O_1900,N_14874,N_12570);
nor UO_1901 (O_1901,N_14037,N_13480);
and UO_1902 (O_1902,N_12615,N_14096);
nand UO_1903 (O_1903,N_14428,N_13019);
xnor UO_1904 (O_1904,N_14731,N_12523);
nor UO_1905 (O_1905,N_14433,N_13280);
nand UO_1906 (O_1906,N_14070,N_14454);
nand UO_1907 (O_1907,N_12686,N_14985);
nor UO_1908 (O_1908,N_12577,N_12366);
and UO_1909 (O_1909,N_12784,N_14672);
and UO_1910 (O_1910,N_13184,N_14942);
xor UO_1911 (O_1911,N_13815,N_14956);
and UO_1912 (O_1912,N_12439,N_12260);
and UO_1913 (O_1913,N_14957,N_12138);
nand UO_1914 (O_1914,N_12251,N_13261);
or UO_1915 (O_1915,N_12161,N_14471);
nand UO_1916 (O_1916,N_14024,N_13366);
or UO_1917 (O_1917,N_13467,N_14933);
nand UO_1918 (O_1918,N_12871,N_12060);
and UO_1919 (O_1919,N_12981,N_12473);
and UO_1920 (O_1920,N_14714,N_12163);
or UO_1921 (O_1921,N_13120,N_12590);
nor UO_1922 (O_1922,N_13511,N_14210);
nand UO_1923 (O_1923,N_12162,N_14071);
or UO_1924 (O_1924,N_12438,N_14164);
or UO_1925 (O_1925,N_14044,N_14181);
nand UO_1926 (O_1926,N_14262,N_14566);
and UO_1927 (O_1927,N_13868,N_14792);
and UO_1928 (O_1928,N_13763,N_12433);
nand UO_1929 (O_1929,N_14780,N_12627);
nor UO_1930 (O_1930,N_12062,N_14614);
nor UO_1931 (O_1931,N_14978,N_14701);
nor UO_1932 (O_1932,N_14360,N_13374);
xnor UO_1933 (O_1933,N_13787,N_12163);
nor UO_1934 (O_1934,N_14837,N_12213);
xor UO_1935 (O_1935,N_12543,N_12022);
or UO_1936 (O_1936,N_12502,N_13438);
or UO_1937 (O_1937,N_13923,N_13876);
nor UO_1938 (O_1938,N_12971,N_14937);
nand UO_1939 (O_1939,N_14943,N_12985);
and UO_1940 (O_1940,N_12840,N_14916);
or UO_1941 (O_1941,N_14069,N_14838);
or UO_1942 (O_1942,N_12866,N_13987);
or UO_1943 (O_1943,N_14020,N_14831);
nand UO_1944 (O_1944,N_14738,N_12110);
nand UO_1945 (O_1945,N_13991,N_13842);
nor UO_1946 (O_1946,N_14455,N_14901);
and UO_1947 (O_1947,N_13757,N_12159);
and UO_1948 (O_1948,N_13397,N_12847);
and UO_1949 (O_1949,N_13251,N_14582);
nand UO_1950 (O_1950,N_12780,N_14446);
nand UO_1951 (O_1951,N_14712,N_14554);
nand UO_1952 (O_1952,N_12240,N_14549);
or UO_1953 (O_1953,N_12805,N_14019);
nand UO_1954 (O_1954,N_14241,N_14984);
nor UO_1955 (O_1955,N_14463,N_13901);
xnor UO_1956 (O_1956,N_14560,N_13014);
or UO_1957 (O_1957,N_14962,N_14840);
and UO_1958 (O_1958,N_12576,N_13640);
nor UO_1959 (O_1959,N_14592,N_12866);
nor UO_1960 (O_1960,N_12846,N_12001);
nand UO_1961 (O_1961,N_14529,N_13445);
nor UO_1962 (O_1962,N_12372,N_12054);
or UO_1963 (O_1963,N_12022,N_13987);
nand UO_1964 (O_1964,N_12397,N_13494);
nor UO_1965 (O_1965,N_12821,N_14865);
and UO_1966 (O_1966,N_14894,N_12647);
and UO_1967 (O_1967,N_12149,N_14725);
nand UO_1968 (O_1968,N_12296,N_12892);
and UO_1969 (O_1969,N_14899,N_13231);
nor UO_1970 (O_1970,N_14922,N_12083);
xnor UO_1971 (O_1971,N_12708,N_14266);
or UO_1972 (O_1972,N_14221,N_14745);
or UO_1973 (O_1973,N_14450,N_14527);
and UO_1974 (O_1974,N_14051,N_12207);
or UO_1975 (O_1975,N_12214,N_13894);
nand UO_1976 (O_1976,N_12044,N_13690);
nor UO_1977 (O_1977,N_12799,N_14805);
or UO_1978 (O_1978,N_13554,N_13421);
and UO_1979 (O_1979,N_12995,N_13499);
nor UO_1980 (O_1980,N_14637,N_14377);
nor UO_1981 (O_1981,N_12454,N_14311);
and UO_1982 (O_1982,N_12147,N_12046);
or UO_1983 (O_1983,N_14548,N_13700);
nand UO_1984 (O_1984,N_14446,N_12743);
or UO_1985 (O_1985,N_12643,N_13676);
and UO_1986 (O_1986,N_12370,N_13449);
and UO_1987 (O_1987,N_12196,N_12989);
and UO_1988 (O_1988,N_14215,N_12286);
and UO_1989 (O_1989,N_12983,N_14270);
and UO_1990 (O_1990,N_12305,N_12295);
xnor UO_1991 (O_1991,N_14073,N_13711);
nor UO_1992 (O_1992,N_14183,N_12243);
nor UO_1993 (O_1993,N_13484,N_14367);
nand UO_1994 (O_1994,N_12884,N_13382);
xnor UO_1995 (O_1995,N_13709,N_13318);
and UO_1996 (O_1996,N_14038,N_12874);
xor UO_1997 (O_1997,N_14394,N_12888);
nand UO_1998 (O_1998,N_13198,N_12259);
and UO_1999 (O_1999,N_14256,N_14877);
endmodule