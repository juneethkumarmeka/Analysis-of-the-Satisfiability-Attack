module basic_750_5000_1000_5_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_85,In_488);
nor U1 (N_1,In_570,In_13);
nor U2 (N_2,In_90,In_377);
nor U3 (N_3,In_422,In_428);
or U4 (N_4,In_356,In_418);
and U5 (N_5,In_330,In_693);
and U6 (N_6,In_541,In_650);
nand U7 (N_7,In_140,In_740);
or U8 (N_8,In_273,In_358);
nand U9 (N_9,In_331,In_383);
and U10 (N_10,In_146,In_456);
nand U11 (N_11,In_133,In_127);
or U12 (N_12,In_74,In_348);
and U13 (N_13,In_228,In_439);
and U14 (N_14,In_26,In_593);
and U15 (N_15,In_100,In_103);
or U16 (N_16,In_705,In_297);
nand U17 (N_17,In_296,In_659);
nand U18 (N_18,In_32,In_65);
nand U19 (N_19,In_204,In_282);
and U20 (N_20,In_8,In_138);
and U21 (N_21,In_697,In_568);
or U22 (N_22,In_76,In_279);
nor U23 (N_23,In_575,In_9);
nor U24 (N_24,In_84,In_641);
nand U25 (N_25,In_125,In_467);
nand U26 (N_26,In_443,In_231);
nand U27 (N_27,In_426,In_445);
nand U28 (N_28,In_70,In_58);
and U29 (N_29,In_724,In_63);
and U30 (N_30,In_116,In_4);
nor U31 (N_31,In_291,In_598);
and U32 (N_32,In_537,In_741);
or U33 (N_33,In_684,In_548);
nand U34 (N_34,In_366,In_216);
or U35 (N_35,In_118,In_491);
or U36 (N_36,In_674,In_66);
and U37 (N_37,In_159,In_478);
or U38 (N_38,In_551,In_723);
and U39 (N_39,In_458,In_122);
and U40 (N_40,In_645,In_80);
or U41 (N_41,In_86,In_303);
nor U42 (N_42,In_171,In_544);
nand U43 (N_43,In_218,In_529);
xnor U44 (N_44,In_599,In_276);
nand U45 (N_45,In_226,In_75);
or U46 (N_46,In_397,In_446);
or U47 (N_47,In_308,In_534);
or U48 (N_48,In_485,In_481);
or U49 (N_49,In_324,In_689);
or U50 (N_50,In_523,In_703);
xor U51 (N_51,In_555,In_380);
nand U52 (N_52,In_245,In_421);
and U53 (N_53,In_442,In_346);
and U54 (N_54,In_253,In_81);
nor U55 (N_55,In_50,In_314);
nor U56 (N_56,In_37,In_293);
and U57 (N_57,In_730,In_547);
or U58 (N_58,In_666,In_620);
or U59 (N_59,In_704,In_25);
nand U60 (N_60,In_427,In_170);
nand U61 (N_61,In_419,In_295);
nand U62 (N_62,In_440,In_721);
nand U63 (N_63,In_482,In_142);
and U64 (N_64,In_135,In_67);
and U65 (N_65,In_670,In_248);
nand U66 (N_66,In_344,In_338);
and U67 (N_67,In_38,In_686);
and U68 (N_68,In_737,In_267);
and U69 (N_69,In_350,In_112);
and U70 (N_70,In_72,In_389);
or U71 (N_71,In_649,In_225);
and U72 (N_72,In_286,In_287);
nor U73 (N_73,In_40,In_718);
and U74 (N_74,In_34,In_474);
and U75 (N_75,In_414,In_706);
and U76 (N_76,In_315,In_434);
nor U77 (N_77,In_243,In_516);
and U78 (N_78,In_317,In_359);
nand U79 (N_79,In_610,In_515);
and U80 (N_80,In_708,In_265);
and U81 (N_81,In_97,In_585);
and U82 (N_82,In_318,In_169);
nor U83 (N_83,In_734,In_640);
nor U84 (N_84,In_99,In_545);
nor U85 (N_85,In_405,In_128);
nand U86 (N_86,In_518,In_29);
nand U87 (N_87,In_46,In_190);
nand U88 (N_88,In_540,In_676);
nand U89 (N_89,In_465,In_633);
nor U90 (N_90,In_347,In_381);
or U91 (N_91,In_357,In_141);
and U92 (N_92,In_20,In_137);
xnor U93 (N_93,In_55,In_672);
or U94 (N_94,In_449,In_96);
or U95 (N_95,In_432,In_305);
nor U96 (N_96,In_307,In_259);
nor U97 (N_97,In_2,In_238);
nor U98 (N_98,In_749,In_725);
nor U99 (N_99,In_56,In_514);
and U100 (N_100,In_617,In_433);
or U101 (N_101,In_503,In_31);
nand U102 (N_102,In_747,In_250);
and U103 (N_103,In_251,In_661);
nor U104 (N_104,In_208,In_664);
or U105 (N_105,In_384,In_24);
or U106 (N_106,In_455,In_326);
or U107 (N_107,In_214,In_742);
nand U108 (N_108,In_584,In_452);
or U109 (N_109,In_416,In_490);
or U110 (N_110,In_471,In_412);
nand U111 (N_111,In_546,In_313);
or U112 (N_112,In_473,In_187);
or U113 (N_113,In_163,In_513);
xnor U114 (N_114,In_487,In_576);
nand U115 (N_115,In_271,In_385);
and U116 (N_116,In_508,In_425);
nor U117 (N_117,In_586,In_589);
or U118 (N_118,In_205,In_158);
and U119 (N_119,In_219,In_378);
and U120 (N_120,In_130,In_626);
nor U121 (N_121,In_373,In_164);
or U122 (N_122,In_506,In_454);
or U123 (N_123,In_212,In_521);
or U124 (N_124,In_281,In_634);
and U125 (N_125,In_677,In_323);
and U126 (N_126,In_531,In_600);
nor U127 (N_127,In_582,In_539);
xnor U128 (N_128,In_681,In_210);
or U129 (N_129,In_517,In_200);
nor U130 (N_130,In_622,In_211);
nand U131 (N_131,In_108,In_566);
nand U132 (N_132,In_727,In_327);
nor U133 (N_133,In_499,In_345);
or U134 (N_134,In_404,In_209);
xnor U135 (N_135,In_731,In_429);
nor U136 (N_136,In_42,In_448);
nor U137 (N_137,In_451,In_290);
nand U138 (N_138,In_193,In_647);
or U139 (N_139,In_289,In_424);
nand U140 (N_140,In_95,In_16);
or U141 (N_141,In_501,In_564);
or U142 (N_142,In_89,In_302);
nand U143 (N_143,In_147,In_520);
nor U144 (N_144,In_646,In_355);
nand U145 (N_145,In_410,In_553);
or U146 (N_146,In_696,In_408);
nand U147 (N_147,In_54,In_614);
and U148 (N_148,In_607,In_68);
and U149 (N_149,In_104,In_463);
nand U150 (N_150,In_561,In_370);
nand U151 (N_151,In_574,In_709);
nand U152 (N_152,In_504,In_682);
nor U153 (N_153,In_401,In_192);
nor U154 (N_154,In_143,In_395);
and U155 (N_155,In_688,In_136);
xnor U156 (N_156,In_538,In_157);
nor U157 (N_157,In_93,In_354);
nand U158 (N_158,In_549,In_325);
xnor U159 (N_159,In_707,In_519);
xnor U160 (N_160,In_241,In_382);
or U161 (N_161,In_583,In_733);
nand U162 (N_162,In_294,In_628);
nand U163 (N_163,In_461,In_167);
xnor U164 (N_164,In_420,In_280);
nor U165 (N_165,In_145,In_713);
or U166 (N_166,In_64,In_699);
or U167 (N_167,In_423,In_675);
nand U168 (N_168,In_19,In_719);
or U169 (N_169,In_18,In_196);
and U170 (N_170,In_83,In_222);
or U171 (N_171,In_444,In_624);
or U172 (N_172,In_14,In_235);
and U173 (N_173,In_562,In_73);
xor U174 (N_174,In_114,In_154);
and U175 (N_175,In_11,In_71);
nand U176 (N_176,In_375,In_581);
nor U177 (N_177,In_217,In_476);
or U178 (N_178,In_363,In_556);
nand U179 (N_179,In_316,In_602);
or U180 (N_180,In_186,In_695);
and U181 (N_181,In_284,In_726);
nand U182 (N_182,In_21,In_340);
and U183 (N_183,In_694,In_413);
nor U184 (N_184,In_691,In_229);
or U185 (N_185,In_144,In_621);
nand U186 (N_186,In_257,In_542);
nand U187 (N_187,In_657,In_181);
nor U188 (N_188,In_198,In_464);
nor U189 (N_189,In_559,In_715);
or U190 (N_190,In_470,In_386);
nand U191 (N_191,In_59,In_61);
and U192 (N_192,In_106,In_391);
or U193 (N_193,In_392,In_179);
or U194 (N_194,In_603,In_60);
and U195 (N_195,In_269,In_616);
nand U196 (N_196,In_285,In_132);
or U197 (N_197,In_342,In_472);
or U198 (N_198,In_105,In_654);
nand U199 (N_199,In_1,In_590);
nor U200 (N_200,In_255,In_215);
and U201 (N_201,In_717,In_189);
nor U202 (N_202,In_417,In_435);
or U203 (N_203,In_258,In_44);
nor U204 (N_204,In_17,In_438);
and U205 (N_205,In_367,In_552);
nor U206 (N_206,In_150,In_644);
or U207 (N_207,In_92,In_609);
and U208 (N_208,In_399,In_195);
or U209 (N_209,In_690,In_403);
nor U210 (N_210,In_606,In_700);
and U211 (N_211,In_129,In_224);
nand U212 (N_212,In_246,In_283);
and U213 (N_213,In_685,In_663);
or U214 (N_214,In_662,In_353);
nand U215 (N_215,In_535,In_123);
and U216 (N_216,In_415,In_45);
nor U217 (N_217,In_374,In_494);
or U218 (N_218,In_394,In_304);
nand U219 (N_219,In_227,In_489);
or U220 (N_220,In_550,In_716);
or U221 (N_221,In_746,In_149);
or U222 (N_222,In_328,In_139);
nand U223 (N_223,In_35,In_220);
nand U224 (N_224,In_495,In_201);
nand U225 (N_225,In_202,In_630);
and U226 (N_226,In_232,In_631);
nor U227 (N_227,In_10,In_580);
and U228 (N_228,In_165,In_447);
and U229 (N_229,In_197,In_743);
nand U230 (N_230,In_369,In_162);
nor U231 (N_231,In_310,In_62);
xnor U232 (N_232,In_173,In_23);
nor U233 (N_233,In_450,In_230);
nand U234 (N_234,In_311,In_236);
and U235 (N_235,In_82,In_642);
nor U236 (N_236,In_720,In_636);
and U237 (N_237,In_364,In_275);
and U238 (N_238,In_680,In_254);
and U239 (N_239,In_333,In_745);
nor U240 (N_240,In_702,In_110);
or U241 (N_241,In_469,In_526);
nor U242 (N_242,In_79,In_505);
nand U243 (N_243,In_563,In_185);
nand U244 (N_244,In_402,In_183);
and U245 (N_245,In_270,In_47);
nand U246 (N_246,In_319,In_388);
and U247 (N_247,In_627,In_161);
or U248 (N_248,In_22,In_48);
nor U249 (N_249,In_595,In_671);
and U250 (N_250,In_572,In_278);
or U251 (N_251,In_479,In_460);
and U252 (N_252,In_252,In_372);
nor U253 (N_253,In_166,In_390);
nor U254 (N_254,In_396,In_368);
or U255 (N_255,In_571,In_365);
nand U256 (N_256,In_36,In_309);
nand U257 (N_257,In_191,In_57);
nor U258 (N_258,In_41,In_507);
nor U259 (N_259,In_288,In_532);
nand U260 (N_260,In_27,In_653);
nand U261 (N_261,In_522,In_618);
and U262 (N_262,In_667,In_605);
or U263 (N_263,In_613,In_502);
nor U264 (N_264,In_554,In_441);
or U265 (N_265,In_665,In_692);
and U266 (N_266,In_52,In_69);
nand U267 (N_267,In_411,In_406);
and U268 (N_268,In_437,In_635);
nor U269 (N_269,In_431,In_329);
nor U270 (N_270,In_119,In_277);
or U271 (N_271,In_632,In_321);
and U272 (N_272,In_459,In_7);
and U273 (N_273,In_673,In_376);
nand U274 (N_274,In_336,In_729);
or U275 (N_275,In_178,In_530);
and U276 (N_276,In_242,In_320);
and U277 (N_277,In_172,In_160);
nor U278 (N_278,In_184,In_739);
nand U279 (N_279,In_379,In_188);
nand U280 (N_280,In_30,In_577);
and U281 (N_281,In_528,In_339);
nand U282 (N_282,In_261,In_651);
and U283 (N_283,In_234,In_560);
nor U284 (N_284,In_203,In_120);
nand U285 (N_285,In_527,In_728);
nor U286 (N_286,In_371,In_223);
or U287 (N_287,In_484,In_77);
nor U288 (N_288,In_639,In_262);
nand U289 (N_289,In_687,In_175);
nor U290 (N_290,In_194,In_496);
nand U291 (N_291,In_714,In_510);
or U292 (N_292,In_237,In_512);
nand U293 (N_293,In_615,In_486);
or U294 (N_294,In_596,In_409);
nand U295 (N_295,In_565,In_592);
nor U296 (N_296,In_156,In_407);
and U297 (N_297,In_131,In_679);
and U298 (N_298,In_398,In_78);
nor U299 (N_299,In_206,In_360);
nand U300 (N_300,In_722,In_115);
xnor U301 (N_301,In_710,In_155);
or U302 (N_302,In_623,In_268);
nor U303 (N_303,In_525,In_352);
nor U304 (N_304,In_591,In_98);
and U305 (N_305,In_263,In_301);
and U306 (N_306,In_588,In_109);
nor U307 (N_307,In_669,In_604);
nor U308 (N_308,In_180,In_87);
and U309 (N_309,In_678,In_711);
or U310 (N_310,In_611,In_477);
and U311 (N_311,In_306,In_264);
and U312 (N_312,In_637,In_299);
or U313 (N_313,In_53,In_608);
nand U314 (N_314,In_334,In_466);
nand U315 (N_315,In_655,In_698);
xnor U316 (N_316,In_49,In_569);
nand U317 (N_317,In_660,In_643);
nand U318 (N_318,In_343,In_249);
nand U319 (N_319,In_744,In_579);
nor U320 (N_320,In_6,In_738);
or U321 (N_321,In_601,In_735);
xor U322 (N_322,In_0,In_199);
nand U323 (N_323,In_28,In_430);
nand U324 (N_324,In_612,In_475);
nand U325 (N_325,In_341,In_524);
nor U326 (N_326,In_619,In_94);
nand U327 (N_327,In_573,In_648);
and U328 (N_328,In_5,In_736);
and U329 (N_329,In_256,In_292);
or U330 (N_330,In_240,In_51);
and U331 (N_331,In_124,In_177);
nand U332 (N_332,In_3,In_168);
nor U333 (N_333,In_126,In_652);
nand U334 (N_334,In_247,In_121);
nor U335 (N_335,In_102,In_543);
nor U336 (N_336,In_625,In_151);
nand U337 (N_337,In_33,In_536);
and U338 (N_338,In_492,In_312);
or U339 (N_339,In_337,In_400);
nor U340 (N_340,In_597,In_393);
and U341 (N_341,In_468,In_683);
nor U342 (N_342,In_39,In_533);
or U343 (N_343,In_213,In_176);
nor U344 (N_344,In_436,In_335);
nor U345 (N_345,In_15,In_349);
or U346 (N_346,In_656,In_594);
or U347 (N_347,In_557,In_658);
or U348 (N_348,In_362,In_509);
nand U349 (N_349,In_701,In_668);
and U350 (N_350,In_567,In_480);
and U351 (N_351,In_260,In_117);
nand U352 (N_352,In_12,In_511);
nor U353 (N_353,In_221,In_483);
nor U354 (N_354,In_587,In_298);
or U355 (N_355,In_712,In_88);
nor U356 (N_356,In_153,In_493);
nand U357 (N_357,In_272,In_732);
xor U358 (N_358,In_101,In_91);
or U359 (N_359,In_361,In_387);
nand U360 (N_360,In_152,In_322);
nor U361 (N_361,In_462,In_274);
and U362 (N_362,In_351,In_638);
and U363 (N_363,In_266,In_300);
or U364 (N_364,In_148,In_239);
nor U365 (N_365,In_453,In_244);
nand U366 (N_366,In_748,In_500);
or U367 (N_367,In_207,In_182);
nor U368 (N_368,In_43,In_498);
or U369 (N_369,In_233,In_332);
and U370 (N_370,In_457,In_497);
nand U371 (N_371,In_134,In_174);
nor U372 (N_372,In_558,In_629);
nand U373 (N_373,In_113,In_578);
or U374 (N_374,In_111,In_107);
and U375 (N_375,In_405,In_330);
xor U376 (N_376,In_264,In_332);
or U377 (N_377,In_280,In_36);
nor U378 (N_378,In_626,In_275);
nor U379 (N_379,In_734,In_369);
and U380 (N_380,In_37,In_396);
nand U381 (N_381,In_533,In_188);
nor U382 (N_382,In_28,In_551);
nor U383 (N_383,In_683,In_688);
and U384 (N_384,In_47,In_284);
nor U385 (N_385,In_749,In_591);
or U386 (N_386,In_498,In_162);
nor U387 (N_387,In_640,In_716);
or U388 (N_388,In_522,In_64);
or U389 (N_389,In_531,In_453);
or U390 (N_390,In_301,In_511);
and U391 (N_391,In_574,In_438);
nor U392 (N_392,In_163,In_429);
or U393 (N_393,In_33,In_302);
and U394 (N_394,In_616,In_163);
nor U395 (N_395,In_489,In_355);
nand U396 (N_396,In_623,In_332);
or U397 (N_397,In_276,In_383);
nor U398 (N_398,In_413,In_741);
or U399 (N_399,In_542,In_85);
nor U400 (N_400,In_377,In_598);
or U401 (N_401,In_152,In_161);
nand U402 (N_402,In_479,In_419);
and U403 (N_403,In_436,In_374);
or U404 (N_404,In_101,In_717);
nand U405 (N_405,In_87,In_553);
and U406 (N_406,In_475,In_217);
and U407 (N_407,In_597,In_598);
or U408 (N_408,In_272,In_506);
nor U409 (N_409,In_210,In_44);
nand U410 (N_410,In_313,In_258);
nor U411 (N_411,In_3,In_82);
or U412 (N_412,In_133,In_72);
or U413 (N_413,In_168,In_497);
and U414 (N_414,In_245,In_690);
or U415 (N_415,In_558,In_309);
or U416 (N_416,In_621,In_691);
and U417 (N_417,In_680,In_718);
or U418 (N_418,In_14,In_639);
nor U419 (N_419,In_497,In_229);
and U420 (N_420,In_329,In_224);
nand U421 (N_421,In_464,In_542);
and U422 (N_422,In_545,In_748);
and U423 (N_423,In_260,In_164);
and U424 (N_424,In_149,In_441);
and U425 (N_425,In_100,In_437);
nand U426 (N_426,In_689,In_42);
nor U427 (N_427,In_320,In_538);
or U428 (N_428,In_442,In_713);
nand U429 (N_429,In_305,In_365);
nor U430 (N_430,In_481,In_459);
or U431 (N_431,In_95,In_51);
and U432 (N_432,In_501,In_555);
or U433 (N_433,In_523,In_444);
nand U434 (N_434,In_301,In_735);
and U435 (N_435,In_364,In_458);
or U436 (N_436,In_92,In_252);
nor U437 (N_437,In_628,In_9);
and U438 (N_438,In_132,In_687);
nor U439 (N_439,In_713,In_628);
or U440 (N_440,In_653,In_626);
nor U441 (N_441,In_383,In_152);
nor U442 (N_442,In_709,In_90);
nor U443 (N_443,In_727,In_150);
or U444 (N_444,In_210,In_554);
and U445 (N_445,In_42,In_85);
or U446 (N_446,In_265,In_665);
nor U447 (N_447,In_526,In_41);
and U448 (N_448,In_50,In_583);
nand U449 (N_449,In_25,In_705);
and U450 (N_450,In_222,In_517);
nand U451 (N_451,In_493,In_615);
nand U452 (N_452,In_600,In_264);
nand U453 (N_453,In_471,In_672);
nand U454 (N_454,In_660,In_11);
nand U455 (N_455,In_182,In_492);
nand U456 (N_456,In_271,In_282);
or U457 (N_457,In_192,In_61);
xor U458 (N_458,In_279,In_552);
nand U459 (N_459,In_625,In_623);
xor U460 (N_460,In_153,In_460);
nand U461 (N_461,In_748,In_145);
and U462 (N_462,In_675,In_124);
or U463 (N_463,In_72,In_670);
nor U464 (N_464,In_537,In_185);
or U465 (N_465,In_627,In_257);
nor U466 (N_466,In_19,In_486);
nor U467 (N_467,In_596,In_408);
nor U468 (N_468,In_331,In_17);
and U469 (N_469,In_584,In_286);
nor U470 (N_470,In_499,In_222);
nand U471 (N_471,In_567,In_315);
and U472 (N_472,In_192,In_107);
or U473 (N_473,In_481,In_720);
or U474 (N_474,In_374,In_702);
and U475 (N_475,In_557,In_257);
nor U476 (N_476,In_568,In_168);
nor U477 (N_477,In_216,In_670);
and U478 (N_478,In_269,In_67);
nand U479 (N_479,In_52,In_582);
nor U480 (N_480,In_222,In_426);
nor U481 (N_481,In_576,In_489);
nand U482 (N_482,In_657,In_221);
and U483 (N_483,In_568,In_709);
or U484 (N_484,In_173,In_436);
and U485 (N_485,In_536,In_399);
nand U486 (N_486,In_14,In_314);
nor U487 (N_487,In_716,In_115);
nor U488 (N_488,In_748,In_429);
nor U489 (N_489,In_555,In_300);
nor U490 (N_490,In_157,In_638);
or U491 (N_491,In_552,In_317);
xnor U492 (N_492,In_549,In_418);
and U493 (N_493,In_330,In_169);
and U494 (N_494,In_562,In_406);
nand U495 (N_495,In_621,In_722);
and U496 (N_496,In_415,In_498);
nor U497 (N_497,In_502,In_339);
and U498 (N_498,In_237,In_39);
nor U499 (N_499,In_534,In_107);
or U500 (N_500,In_712,In_159);
or U501 (N_501,In_601,In_508);
nor U502 (N_502,In_558,In_725);
nor U503 (N_503,In_712,In_222);
nand U504 (N_504,In_222,In_22);
nor U505 (N_505,In_313,In_182);
and U506 (N_506,In_199,In_192);
nor U507 (N_507,In_535,In_371);
nand U508 (N_508,In_472,In_195);
nor U509 (N_509,In_719,In_282);
or U510 (N_510,In_302,In_344);
and U511 (N_511,In_703,In_456);
or U512 (N_512,In_592,In_616);
nor U513 (N_513,In_262,In_313);
nor U514 (N_514,In_548,In_101);
or U515 (N_515,In_551,In_453);
nor U516 (N_516,In_615,In_23);
nand U517 (N_517,In_258,In_185);
nor U518 (N_518,In_442,In_477);
or U519 (N_519,In_469,In_326);
nor U520 (N_520,In_629,In_447);
or U521 (N_521,In_425,In_387);
nor U522 (N_522,In_134,In_649);
nor U523 (N_523,In_515,In_93);
and U524 (N_524,In_328,In_240);
nor U525 (N_525,In_243,In_17);
or U526 (N_526,In_123,In_148);
and U527 (N_527,In_217,In_80);
and U528 (N_528,In_126,In_50);
nor U529 (N_529,In_235,In_491);
or U530 (N_530,In_187,In_29);
or U531 (N_531,In_631,In_177);
nor U532 (N_532,In_338,In_630);
nand U533 (N_533,In_265,In_433);
or U534 (N_534,In_391,In_524);
or U535 (N_535,In_362,In_127);
or U536 (N_536,In_133,In_262);
nor U537 (N_537,In_159,In_83);
or U538 (N_538,In_629,In_444);
nor U539 (N_539,In_253,In_577);
nand U540 (N_540,In_712,In_527);
nor U541 (N_541,In_438,In_80);
or U542 (N_542,In_56,In_467);
nor U543 (N_543,In_215,In_40);
or U544 (N_544,In_422,In_73);
and U545 (N_545,In_351,In_231);
nand U546 (N_546,In_334,In_181);
or U547 (N_547,In_729,In_548);
nor U548 (N_548,In_397,In_743);
or U549 (N_549,In_236,In_443);
or U550 (N_550,In_141,In_315);
nand U551 (N_551,In_236,In_344);
nor U552 (N_552,In_628,In_390);
nor U553 (N_553,In_691,In_653);
or U554 (N_554,In_378,In_682);
or U555 (N_555,In_31,In_125);
nor U556 (N_556,In_590,In_739);
nor U557 (N_557,In_130,In_49);
nand U558 (N_558,In_244,In_509);
nand U559 (N_559,In_398,In_651);
or U560 (N_560,In_430,In_182);
nor U561 (N_561,In_6,In_511);
and U562 (N_562,In_388,In_396);
nor U563 (N_563,In_722,In_733);
nor U564 (N_564,In_195,In_689);
and U565 (N_565,In_572,In_157);
nand U566 (N_566,In_404,In_40);
or U567 (N_567,In_46,In_731);
or U568 (N_568,In_468,In_318);
and U569 (N_569,In_542,In_657);
and U570 (N_570,In_154,In_457);
nand U571 (N_571,In_698,In_706);
and U572 (N_572,In_724,In_287);
and U573 (N_573,In_272,In_187);
nor U574 (N_574,In_264,In_254);
or U575 (N_575,In_556,In_652);
nor U576 (N_576,In_654,In_195);
or U577 (N_577,In_314,In_595);
xnor U578 (N_578,In_548,In_627);
nor U579 (N_579,In_323,In_110);
or U580 (N_580,In_101,In_547);
or U581 (N_581,In_520,In_438);
and U582 (N_582,In_408,In_191);
and U583 (N_583,In_55,In_422);
and U584 (N_584,In_738,In_401);
and U585 (N_585,In_332,In_608);
nand U586 (N_586,In_561,In_85);
nand U587 (N_587,In_313,In_456);
and U588 (N_588,In_583,In_62);
and U589 (N_589,In_412,In_705);
nor U590 (N_590,In_606,In_159);
nand U591 (N_591,In_320,In_544);
and U592 (N_592,In_321,In_729);
nand U593 (N_593,In_592,In_658);
and U594 (N_594,In_634,In_559);
and U595 (N_595,In_208,In_476);
nand U596 (N_596,In_201,In_542);
nand U597 (N_597,In_335,In_164);
nand U598 (N_598,In_697,In_162);
and U599 (N_599,In_484,In_667);
and U600 (N_600,In_556,In_616);
nor U601 (N_601,In_96,In_711);
and U602 (N_602,In_387,In_510);
nor U603 (N_603,In_502,In_266);
or U604 (N_604,In_453,In_485);
nor U605 (N_605,In_411,In_343);
nor U606 (N_606,In_67,In_501);
and U607 (N_607,In_49,In_154);
nor U608 (N_608,In_99,In_45);
nand U609 (N_609,In_275,In_77);
and U610 (N_610,In_728,In_451);
or U611 (N_611,In_168,In_146);
or U612 (N_612,In_208,In_94);
xor U613 (N_613,In_324,In_577);
nor U614 (N_614,In_34,In_173);
and U615 (N_615,In_271,In_338);
or U616 (N_616,In_594,In_302);
or U617 (N_617,In_110,In_119);
xor U618 (N_618,In_540,In_351);
nand U619 (N_619,In_188,In_273);
or U620 (N_620,In_414,In_348);
and U621 (N_621,In_674,In_373);
or U622 (N_622,In_144,In_633);
and U623 (N_623,In_499,In_60);
and U624 (N_624,In_312,In_25);
nand U625 (N_625,In_730,In_647);
or U626 (N_626,In_662,In_491);
nor U627 (N_627,In_617,In_553);
nand U628 (N_628,In_600,In_308);
nand U629 (N_629,In_182,In_464);
or U630 (N_630,In_380,In_626);
or U631 (N_631,In_171,In_504);
or U632 (N_632,In_78,In_42);
nand U633 (N_633,In_61,In_297);
nor U634 (N_634,In_343,In_182);
nand U635 (N_635,In_316,In_341);
nor U636 (N_636,In_346,In_589);
xor U637 (N_637,In_482,In_343);
or U638 (N_638,In_484,In_12);
or U639 (N_639,In_702,In_386);
nor U640 (N_640,In_261,In_116);
nand U641 (N_641,In_463,In_239);
nand U642 (N_642,In_629,In_355);
and U643 (N_643,In_519,In_739);
nand U644 (N_644,In_320,In_299);
nand U645 (N_645,In_600,In_76);
or U646 (N_646,In_32,In_383);
or U647 (N_647,In_507,In_187);
nand U648 (N_648,In_302,In_54);
nand U649 (N_649,In_418,In_210);
nand U650 (N_650,In_619,In_394);
or U651 (N_651,In_356,In_485);
and U652 (N_652,In_503,In_708);
and U653 (N_653,In_144,In_690);
and U654 (N_654,In_49,In_153);
nor U655 (N_655,In_209,In_712);
nand U656 (N_656,In_570,In_323);
nand U657 (N_657,In_303,In_355);
nand U658 (N_658,In_69,In_551);
and U659 (N_659,In_576,In_329);
and U660 (N_660,In_552,In_477);
and U661 (N_661,In_53,In_553);
or U662 (N_662,In_101,In_736);
or U663 (N_663,In_232,In_677);
nor U664 (N_664,In_202,In_85);
nand U665 (N_665,In_410,In_396);
nor U666 (N_666,In_126,In_108);
nor U667 (N_667,In_612,In_545);
nand U668 (N_668,In_199,In_731);
or U669 (N_669,In_253,In_182);
or U670 (N_670,In_66,In_714);
nor U671 (N_671,In_460,In_409);
nor U672 (N_672,In_598,In_32);
or U673 (N_673,In_524,In_352);
and U674 (N_674,In_108,In_731);
and U675 (N_675,In_95,In_536);
nor U676 (N_676,In_585,In_711);
nand U677 (N_677,In_68,In_480);
or U678 (N_678,In_731,In_556);
nor U679 (N_679,In_380,In_514);
nand U680 (N_680,In_217,In_146);
nand U681 (N_681,In_246,In_371);
or U682 (N_682,In_282,In_299);
or U683 (N_683,In_460,In_639);
or U684 (N_684,In_222,In_367);
or U685 (N_685,In_550,In_522);
nand U686 (N_686,In_272,In_247);
nand U687 (N_687,In_282,In_89);
or U688 (N_688,In_652,In_120);
or U689 (N_689,In_570,In_144);
nor U690 (N_690,In_146,In_705);
and U691 (N_691,In_473,In_304);
nand U692 (N_692,In_85,In_466);
and U693 (N_693,In_529,In_227);
nor U694 (N_694,In_388,In_5);
nor U695 (N_695,In_124,In_592);
and U696 (N_696,In_448,In_566);
and U697 (N_697,In_548,In_613);
or U698 (N_698,In_253,In_269);
nand U699 (N_699,In_243,In_51);
or U700 (N_700,In_646,In_587);
or U701 (N_701,In_297,In_680);
nand U702 (N_702,In_489,In_566);
nor U703 (N_703,In_477,In_643);
nor U704 (N_704,In_67,In_66);
nor U705 (N_705,In_670,In_492);
or U706 (N_706,In_459,In_340);
and U707 (N_707,In_163,In_358);
xnor U708 (N_708,In_321,In_430);
and U709 (N_709,In_716,In_693);
nor U710 (N_710,In_351,In_639);
or U711 (N_711,In_416,In_578);
xor U712 (N_712,In_681,In_172);
nor U713 (N_713,In_718,In_440);
and U714 (N_714,In_565,In_384);
nand U715 (N_715,In_15,In_426);
nor U716 (N_716,In_233,In_278);
nand U717 (N_717,In_481,In_465);
nand U718 (N_718,In_661,In_2);
nand U719 (N_719,In_178,In_559);
and U720 (N_720,In_13,In_14);
nand U721 (N_721,In_340,In_623);
xnor U722 (N_722,In_146,In_679);
or U723 (N_723,In_367,In_532);
or U724 (N_724,In_429,In_208);
nand U725 (N_725,In_402,In_718);
or U726 (N_726,In_53,In_87);
nand U727 (N_727,In_681,In_272);
nor U728 (N_728,In_528,In_72);
nor U729 (N_729,In_458,In_103);
or U730 (N_730,In_381,In_201);
and U731 (N_731,In_527,In_379);
nor U732 (N_732,In_204,In_177);
nor U733 (N_733,In_108,In_441);
nand U734 (N_734,In_337,In_167);
nand U735 (N_735,In_202,In_282);
nor U736 (N_736,In_642,In_90);
and U737 (N_737,In_742,In_267);
or U738 (N_738,In_519,In_173);
nand U739 (N_739,In_270,In_80);
nand U740 (N_740,In_467,In_584);
and U741 (N_741,In_465,In_244);
nand U742 (N_742,In_319,In_645);
and U743 (N_743,In_255,In_661);
and U744 (N_744,In_459,In_506);
nand U745 (N_745,In_237,In_387);
nor U746 (N_746,In_499,In_71);
or U747 (N_747,In_503,In_572);
and U748 (N_748,In_318,In_240);
nor U749 (N_749,In_414,In_260);
or U750 (N_750,In_471,In_705);
nor U751 (N_751,In_449,In_465);
xnor U752 (N_752,In_475,In_719);
or U753 (N_753,In_663,In_530);
or U754 (N_754,In_314,In_671);
nand U755 (N_755,In_253,In_129);
and U756 (N_756,In_661,In_492);
nor U757 (N_757,In_105,In_35);
nor U758 (N_758,In_10,In_655);
nand U759 (N_759,In_90,In_111);
and U760 (N_760,In_521,In_285);
or U761 (N_761,In_640,In_695);
nor U762 (N_762,In_440,In_427);
and U763 (N_763,In_145,In_604);
or U764 (N_764,In_416,In_320);
nand U765 (N_765,In_507,In_511);
and U766 (N_766,In_206,In_413);
or U767 (N_767,In_402,In_526);
nor U768 (N_768,In_268,In_519);
nand U769 (N_769,In_435,In_185);
and U770 (N_770,In_338,In_387);
or U771 (N_771,In_521,In_41);
and U772 (N_772,In_39,In_75);
nor U773 (N_773,In_17,In_355);
nand U774 (N_774,In_105,In_325);
nand U775 (N_775,In_230,In_560);
nor U776 (N_776,In_598,In_237);
nand U777 (N_777,In_383,In_471);
xor U778 (N_778,In_674,In_739);
or U779 (N_779,In_545,In_57);
or U780 (N_780,In_274,In_548);
nand U781 (N_781,In_461,In_5);
nor U782 (N_782,In_484,In_567);
nor U783 (N_783,In_372,In_669);
nor U784 (N_784,In_489,In_123);
nor U785 (N_785,In_645,In_513);
and U786 (N_786,In_678,In_716);
nand U787 (N_787,In_658,In_139);
or U788 (N_788,In_283,In_145);
nor U789 (N_789,In_74,In_355);
nor U790 (N_790,In_747,In_110);
and U791 (N_791,In_573,In_40);
nor U792 (N_792,In_703,In_378);
or U793 (N_793,In_264,In_79);
and U794 (N_794,In_232,In_185);
and U795 (N_795,In_202,In_639);
nand U796 (N_796,In_477,In_65);
and U797 (N_797,In_613,In_402);
nor U798 (N_798,In_293,In_7);
and U799 (N_799,In_74,In_688);
nand U800 (N_800,In_602,In_276);
and U801 (N_801,In_84,In_461);
nand U802 (N_802,In_401,In_548);
or U803 (N_803,In_293,In_343);
and U804 (N_804,In_513,In_514);
nor U805 (N_805,In_743,In_567);
and U806 (N_806,In_669,In_552);
and U807 (N_807,In_642,In_154);
nor U808 (N_808,In_166,In_418);
nand U809 (N_809,In_373,In_439);
or U810 (N_810,In_652,In_434);
nand U811 (N_811,In_677,In_282);
nand U812 (N_812,In_709,In_619);
nand U813 (N_813,In_337,In_713);
xor U814 (N_814,In_162,In_582);
nor U815 (N_815,In_338,In_86);
nand U816 (N_816,In_365,In_434);
nand U817 (N_817,In_157,In_176);
and U818 (N_818,In_67,In_22);
and U819 (N_819,In_26,In_631);
and U820 (N_820,In_693,In_295);
or U821 (N_821,In_327,In_600);
nand U822 (N_822,In_702,In_531);
nor U823 (N_823,In_300,In_90);
and U824 (N_824,In_728,In_208);
nand U825 (N_825,In_322,In_364);
nor U826 (N_826,In_24,In_106);
nor U827 (N_827,In_648,In_234);
nor U828 (N_828,In_481,In_280);
nand U829 (N_829,In_317,In_114);
nor U830 (N_830,In_15,In_485);
or U831 (N_831,In_496,In_173);
nand U832 (N_832,In_732,In_746);
nor U833 (N_833,In_33,In_3);
nand U834 (N_834,In_415,In_473);
xor U835 (N_835,In_354,In_542);
and U836 (N_836,In_273,In_619);
or U837 (N_837,In_40,In_156);
nand U838 (N_838,In_695,In_545);
and U839 (N_839,In_682,In_150);
and U840 (N_840,In_295,In_522);
nand U841 (N_841,In_303,In_643);
and U842 (N_842,In_705,In_477);
nor U843 (N_843,In_15,In_601);
or U844 (N_844,In_28,In_528);
nor U845 (N_845,In_296,In_15);
nand U846 (N_846,In_588,In_270);
and U847 (N_847,In_384,In_664);
nand U848 (N_848,In_735,In_706);
nor U849 (N_849,In_138,In_85);
nor U850 (N_850,In_153,In_550);
nand U851 (N_851,In_483,In_17);
nor U852 (N_852,In_77,In_7);
and U853 (N_853,In_465,In_716);
and U854 (N_854,In_600,In_172);
and U855 (N_855,In_662,In_719);
nor U856 (N_856,In_599,In_383);
and U857 (N_857,In_65,In_629);
and U858 (N_858,In_513,In_637);
nand U859 (N_859,In_432,In_730);
nand U860 (N_860,In_60,In_577);
or U861 (N_861,In_357,In_86);
nor U862 (N_862,In_303,In_604);
nand U863 (N_863,In_564,In_33);
and U864 (N_864,In_562,In_605);
and U865 (N_865,In_290,In_262);
nand U866 (N_866,In_36,In_270);
and U867 (N_867,In_406,In_12);
or U868 (N_868,In_418,In_635);
nor U869 (N_869,In_670,In_109);
and U870 (N_870,In_538,In_153);
nor U871 (N_871,In_343,In_723);
and U872 (N_872,In_578,In_591);
and U873 (N_873,In_547,In_597);
or U874 (N_874,In_67,In_589);
and U875 (N_875,In_312,In_695);
or U876 (N_876,In_621,In_557);
or U877 (N_877,In_15,In_119);
nor U878 (N_878,In_357,In_189);
and U879 (N_879,In_528,In_120);
xnor U880 (N_880,In_158,In_624);
or U881 (N_881,In_242,In_315);
and U882 (N_882,In_49,In_219);
nand U883 (N_883,In_743,In_735);
and U884 (N_884,In_152,In_354);
nor U885 (N_885,In_560,In_433);
and U886 (N_886,In_254,In_666);
nor U887 (N_887,In_93,In_673);
or U888 (N_888,In_94,In_75);
or U889 (N_889,In_341,In_211);
nor U890 (N_890,In_434,In_217);
or U891 (N_891,In_738,In_318);
and U892 (N_892,In_690,In_414);
or U893 (N_893,In_71,In_280);
nor U894 (N_894,In_44,In_193);
and U895 (N_895,In_537,In_611);
nor U896 (N_896,In_295,In_633);
and U897 (N_897,In_69,In_134);
or U898 (N_898,In_659,In_91);
or U899 (N_899,In_187,In_600);
nor U900 (N_900,In_129,In_346);
nor U901 (N_901,In_480,In_298);
or U902 (N_902,In_235,In_498);
nand U903 (N_903,In_441,In_519);
nand U904 (N_904,In_219,In_614);
nor U905 (N_905,In_258,In_60);
nor U906 (N_906,In_235,In_199);
or U907 (N_907,In_648,In_24);
nor U908 (N_908,In_649,In_27);
nand U909 (N_909,In_706,In_10);
nor U910 (N_910,In_466,In_457);
or U911 (N_911,In_149,In_595);
nor U912 (N_912,In_164,In_610);
nor U913 (N_913,In_176,In_246);
and U914 (N_914,In_74,In_424);
xnor U915 (N_915,In_356,In_303);
nand U916 (N_916,In_744,In_243);
nand U917 (N_917,In_160,In_198);
nor U918 (N_918,In_637,In_574);
nand U919 (N_919,In_402,In_703);
and U920 (N_920,In_476,In_154);
nand U921 (N_921,In_469,In_61);
nand U922 (N_922,In_165,In_456);
or U923 (N_923,In_722,In_268);
nor U924 (N_924,In_353,In_59);
nor U925 (N_925,In_629,In_246);
nand U926 (N_926,In_730,In_402);
nor U927 (N_927,In_727,In_749);
nor U928 (N_928,In_15,In_301);
nor U929 (N_929,In_462,In_409);
xor U930 (N_930,In_279,In_180);
or U931 (N_931,In_619,In_266);
or U932 (N_932,In_496,In_39);
nor U933 (N_933,In_530,In_608);
nor U934 (N_934,In_95,In_199);
nand U935 (N_935,In_738,In_252);
and U936 (N_936,In_228,In_576);
nand U937 (N_937,In_589,In_336);
or U938 (N_938,In_499,In_502);
nand U939 (N_939,In_466,In_19);
nor U940 (N_940,In_242,In_644);
or U941 (N_941,In_721,In_2);
or U942 (N_942,In_627,In_188);
and U943 (N_943,In_707,In_15);
and U944 (N_944,In_238,In_628);
and U945 (N_945,In_19,In_178);
nor U946 (N_946,In_413,In_13);
or U947 (N_947,In_85,In_17);
nand U948 (N_948,In_62,In_160);
and U949 (N_949,In_557,In_695);
nand U950 (N_950,In_1,In_558);
and U951 (N_951,In_51,In_504);
nor U952 (N_952,In_748,In_352);
nor U953 (N_953,In_228,In_736);
nor U954 (N_954,In_55,In_33);
nor U955 (N_955,In_546,In_94);
and U956 (N_956,In_259,In_323);
nand U957 (N_957,In_340,In_97);
nor U958 (N_958,In_328,In_634);
nor U959 (N_959,In_631,In_738);
nand U960 (N_960,In_487,In_129);
or U961 (N_961,In_689,In_183);
nor U962 (N_962,In_683,In_351);
nand U963 (N_963,In_362,In_262);
nand U964 (N_964,In_488,In_453);
or U965 (N_965,In_88,In_428);
nand U966 (N_966,In_47,In_327);
nand U967 (N_967,In_409,In_6);
nor U968 (N_968,In_77,In_510);
nor U969 (N_969,In_336,In_228);
nor U970 (N_970,In_617,In_88);
or U971 (N_971,In_302,In_616);
xnor U972 (N_972,In_369,In_643);
nand U973 (N_973,In_31,In_719);
or U974 (N_974,In_192,In_361);
nor U975 (N_975,In_695,In_143);
nand U976 (N_976,In_284,In_572);
nor U977 (N_977,In_268,In_300);
nand U978 (N_978,In_86,In_246);
nand U979 (N_979,In_443,In_584);
nor U980 (N_980,In_381,In_68);
nand U981 (N_981,In_653,In_426);
and U982 (N_982,In_85,In_25);
or U983 (N_983,In_47,In_335);
nand U984 (N_984,In_304,In_299);
and U985 (N_985,In_648,In_345);
and U986 (N_986,In_272,In_465);
or U987 (N_987,In_613,In_618);
xnor U988 (N_988,In_636,In_531);
and U989 (N_989,In_425,In_279);
nor U990 (N_990,In_58,In_42);
nand U991 (N_991,In_293,In_632);
and U992 (N_992,In_698,In_741);
or U993 (N_993,In_186,In_128);
or U994 (N_994,In_399,In_355);
and U995 (N_995,In_282,In_154);
and U996 (N_996,In_493,In_429);
or U997 (N_997,In_578,In_7);
and U998 (N_998,In_318,In_235);
nor U999 (N_999,In_470,In_253);
xnor U1000 (N_1000,N_950,N_843);
nor U1001 (N_1001,N_873,N_204);
or U1002 (N_1002,N_452,N_327);
nor U1003 (N_1003,N_37,N_460);
or U1004 (N_1004,N_122,N_223);
and U1005 (N_1005,N_287,N_389);
and U1006 (N_1006,N_170,N_675);
or U1007 (N_1007,N_709,N_713);
nand U1008 (N_1008,N_761,N_681);
or U1009 (N_1009,N_150,N_784);
nor U1010 (N_1010,N_616,N_774);
and U1011 (N_1011,N_356,N_371);
or U1012 (N_1012,N_173,N_752);
and U1013 (N_1013,N_956,N_145);
and U1014 (N_1014,N_509,N_545);
and U1015 (N_1015,N_680,N_78);
or U1016 (N_1016,N_350,N_504);
nand U1017 (N_1017,N_864,N_470);
xnor U1018 (N_1018,N_455,N_800);
xnor U1019 (N_1019,N_662,N_857);
nor U1020 (N_1020,N_505,N_706);
nor U1021 (N_1021,N_912,N_778);
nand U1022 (N_1022,N_921,N_406);
and U1023 (N_1023,N_941,N_157);
nand U1024 (N_1024,N_478,N_746);
nand U1025 (N_1025,N_253,N_334);
nand U1026 (N_1026,N_533,N_717);
nand U1027 (N_1027,N_887,N_523);
or U1028 (N_1028,N_386,N_298);
and U1029 (N_1029,N_314,N_937);
or U1030 (N_1030,N_485,N_898);
and U1031 (N_1031,N_495,N_359);
nor U1032 (N_1032,N_27,N_559);
nand U1033 (N_1033,N_127,N_890);
nand U1034 (N_1034,N_189,N_560);
nor U1035 (N_1035,N_648,N_538);
nor U1036 (N_1036,N_530,N_918);
nor U1037 (N_1037,N_259,N_349);
or U1038 (N_1038,N_823,N_914);
nand U1039 (N_1039,N_95,N_420);
nor U1040 (N_1040,N_771,N_610);
and U1041 (N_1041,N_454,N_922);
nand U1042 (N_1042,N_38,N_80);
nand U1043 (N_1043,N_656,N_753);
xnor U1044 (N_1044,N_839,N_989);
nand U1045 (N_1045,N_623,N_834);
or U1046 (N_1046,N_97,N_198);
or U1047 (N_1047,N_479,N_114);
or U1048 (N_1048,N_197,N_469);
or U1049 (N_1049,N_501,N_368);
nand U1050 (N_1050,N_388,N_531);
or U1051 (N_1051,N_930,N_614);
or U1052 (N_1052,N_468,N_280);
or U1053 (N_1053,N_190,N_273);
nand U1054 (N_1054,N_982,N_626);
nand U1055 (N_1055,N_385,N_894);
nor U1056 (N_1056,N_674,N_810);
nor U1057 (N_1057,N_540,N_836);
nor U1058 (N_1058,N_855,N_311);
nand U1059 (N_1059,N_442,N_975);
and U1060 (N_1060,N_397,N_377);
or U1061 (N_1061,N_443,N_965);
and U1062 (N_1062,N_715,N_831);
or U1063 (N_1063,N_510,N_536);
nand U1064 (N_1064,N_735,N_724);
nor U1065 (N_1065,N_883,N_867);
and U1066 (N_1066,N_727,N_801);
or U1067 (N_1067,N_720,N_983);
or U1068 (N_1068,N_151,N_811);
nor U1069 (N_1069,N_436,N_765);
nor U1070 (N_1070,N_427,N_116);
and U1071 (N_1071,N_878,N_144);
nand U1072 (N_1072,N_544,N_872);
and U1073 (N_1073,N_971,N_14);
nand U1074 (N_1074,N_790,N_696);
and U1075 (N_1075,N_26,N_324);
or U1076 (N_1076,N_275,N_938);
or U1077 (N_1077,N_863,N_591);
and U1078 (N_1078,N_686,N_734);
and U1079 (N_1079,N_16,N_340);
nand U1080 (N_1080,N_940,N_722);
nor U1081 (N_1081,N_848,N_94);
and U1082 (N_1082,N_98,N_453);
or U1083 (N_1083,N_457,N_174);
nor U1084 (N_1084,N_669,N_488);
nand U1085 (N_1085,N_998,N_758);
nand U1086 (N_1086,N_780,N_683);
nor U1087 (N_1087,N_240,N_243);
nand U1088 (N_1088,N_827,N_318);
nor U1089 (N_1089,N_900,N_805);
nand U1090 (N_1090,N_550,N_247);
xor U1091 (N_1091,N_302,N_3);
nand U1092 (N_1092,N_134,N_797);
nor U1093 (N_1093,N_136,N_730);
or U1094 (N_1094,N_104,N_56);
nand U1095 (N_1095,N_685,N_682);
and U1096 (N_1096,N_117,N_807);
or U1097 (N_1097,N_928,N_375);
and U1098 (N_1098,N_2,N_245);
nor U1099 (N_1099,N_160,N_407);
nand U1100 (N_1100,N_897,N_202);
and U1101 (N_1101,N_339,N_343);
and U1102 (N_1102,N_83,N_789);
and U1103 (N_1103,N_307,N_363);
nor U1104 (N_1104,N_361,N_796);
or U1105 (N_1105,N_188,N_191);
nor U1106 (N_1106,N_747,N_946);
or U1107 (N_1107,N_721,N_901);
and U1108 (N_1108,N_896,N_668);
nand U1109 (N_1109,N_647,N_216);
and U1110 (N_1110,N_714,N_885);
nand U1111 (N_1111,N_152,N_574);
and U1112 (N_1112,N_988,N_963);
and U1113 (N_1113,N_667,N_945);
or U1114 (N_1114,N_760,N_292);
and U1115 (N_1115,N_596,N_640);
and U1116 (N_1116,N_233,N_698);
nand U1117 (N_1117,N_519,N_953);
or U1118 (N_1118,N_512,N_132);
nor U1119 (N_1119,N_776,N_165);
nor U1120 (N_1120,N_281,N_909);
nor U1121 (N_1121,N_399,N_392);
and U1122 (N_1122,N_781,N_603);
nand U1123 (N_1123,N_858,N_105);
nand U1124 (N_1124,N_611,N_820);
and U1125 (N_1125,N_597,N_579);
or U1126 (N_1126,N_300,N_594);
nand U1127 (N_1127,N_237,N_756);
or U1128 (N_1128,N_75,N_426);
and U1129 (N_1129,N_659,N_907);
nand U1130 (N_1130,N_21,N_718);
and U1131 (N_1131,N_33,N_379);
nor U1132 (N_1132,N_120,N_353);
nor U1133 (N_1133,N_217,N_955);
or U1134 (N_1134,N_411,N_321);
and U1135 (N_1135,N_783,N_565);
and U1136 (N_1136,N_653,N_415);
or U1137 (N_1137,N_396,N_703);
and U1138 (N_1138,N_974,N_68);
nand U1139 (N_1139,N_218,N_64);
nand U1140 (N_1140,N_847,N_121);
nand U1141 (N_1141,N_258,N_459);
and U1142 (N_1142,N_507,N_642);
or U1143 (N_1143,N_743,N_13);
and U1144 (N_1144,N_141,N_499);
and U1145 (N_1145,N_187,N_936);
nand U1146 (N_1146,N_705,N_566);
nand U1147 (N_1147,N_486,N_36);
xnor U1148 (N_1148,N_200,N_414);
or U1149 (N_1149,N_658,N_993);
nor U1150 (N_1150,N_893,N_369);
or U1151 (N_1151,N_913,N_702);
and U1152 (N_1152,N_607,N_618);
and U1153 (N_1153,N_148,N_40);
and U1154 (N_1154,N_837,N_562);
nor U1155 (N_1155,N_39,N_90);
or U1156 (N_1156,N_335,N_973);
nor U1157 (N_1157,N_865,N_466);
nor U1158 (N_1158,N_193,N_215);
and U1159 (N_1159,N_8,N_808);
and U1160 (N_1160,N_976,N_582);
and U1161 (N_1161,N_299,N_429);
or U1162 (N_1162,N_627,N_31);
and U1163 (N_1163,N_358,N_35);
or U1164 (N_1164,N_333,N_91);
nor U1165 (N_1165,N_860,N_815);
nand U1166 (N_1166,N_589,N_646);
nand U1167 (N_1167,N_265,N_413);
nor U1168 (N_1168,N_73,N_986);
and U1169 (N_1169,N_410,N_214);
nand U1170 (N_1170,N_842,N_851);
nor U1171 (N_1171,N_347,N_85);
nand U1172 (N_1172,N_841,N_471);
xnor U1173 (N_1173,N_553,N_360);
nor U1174 (N_1174,N_556,N_641);
nand U1175 (N_1175,N_547,N_517);
or U1176 (N_1176,N_34,N_849);
and U1177 (N_1177,N_739,N_42);
and U1178 (N_1178,N_467,N_929);
and U1179 (N_1179,N_395,N_862);
and U1180 (N_1180,N_874,N_664);
nor U1181 (N_1181,N_111,N_309);
and U1182 (N_1182,N_393,N_248);
nand U1183 (N_1183,N_795,N_301);
and U1184 (N_1184,N_18,N_777);
nor U1185 (N_1185,N_767,N_629);
xor U1186 (N_1186,N_135,N_451);
nor U1187 (N_1187,N_403,N_764);
or U1188 (N_1188,N_516,N_101);
and U1189 (N_1189,N_923,N_72);
or U1190 (N_1190,N_346,N_390);
nor U1191 (N_1191,N_79,N_483);
nand U1192 (N_1192,N_665,N_163);
nand U1193 (N_1193,N_179,N_182);
and U1194 (N_1194,N_711,N_306);
and U1195 (N_1195,N_231,N_374);
nor U1196 (N_1196,N_645,N_252);
and U1197 (N_1197,N_100,N_364);
nand U1198 (N_1198,N_690,N_147);
nand U1199 (N_1199,N_112,N_477);
nand U1200 (N_1200,N_551,N_167);
nor U1201 (N_1201,N_438,N_159);
nor U1202 (N_1202,N_969,N_759);
nand U1203 (N_1203,N_813,N_944);
and U1204 (N_1204,N_405,N_661);
nor U1205 (N_1205,N_155,N_854);
xnor U1206 (N_1206,N_593,N_818);
nand U1207 (N_1207,N_274,N_329);
or U1208 (N_1208,N_323,N_769);
nand U1209 (N_1209,N_828,N_20);
and U1210 (N_1210,N_313,N_511);
xor U1211 (N_1211,N_272,N_497);
nand U1212 (N_1212,N_107,N_67);
and U1213 (N_1213,N_908,N_639);
nor U1214 (N_1214,N_180,N_979);
and U1215 (N_1215,N_564,N_161);
or U1216 (N_1216,N_183,N_524);
nand U1217 (N_1217,N_961,N_241);
nor U1218 (N_1218,N_490,N_87);
or U1219 (N_1219,N_916,N_201);
nor U1220 (N_1220,N_701,N_555);
and U1221 (N_1221,N_525,N_844);
or U1222 (N_1222,N_581,N_316);
and U1223 (N_1223,N_49,N_82);
xor U1224 (N_1224,N_732,N_425);
or U1225 (N_1225,N_745,N_169);
nor U1226 (N_1226,N_447,N_268);
or U1227 (N_1227,N_254,N_81);
nand U1228 (N_1228,N_17,N_370);
and U1229 (N_1229,N_554,N_348);
nor U1230 (N_1230,N_513,N_373);
or U1231 (N_1231,N_242,N_943);
or U1232 (N_1232,N_417,N_766);
nor U1233 (N_1233,N_870,N_617);
or U1234 (N_1234,N_644,N_376);
xor U1235 (N_1235,N_768,N_999);
nor U1236 (N_1236,N_598,N_716);
nand U1237 (N_1237,N_331,N_239);
or U1238 (N_1238,N_51,N_521);
nor U1239 (N_1239,N_880,N_773);
or U1240 (N_1240,N_297,N_32);
or U1241 (N_1241,N_322,N_0);
nand U1242 (N_1242,N_382,N_22);
and U1243 (N_1243,N_192,N_137);
nand U1244 (N_1244,N_125,N_877);
nor U1245 (N_1245,N_852,N_723);
and U1246 (N_1246,N_991,N_261);
and U1247 (N_1247,N_948,N_6);
nor U1248 (N_1248,N_557,N_431);
xor U1249 (N_1249,N_255,N_688);
nor U1250 (N_1250,N_599,N_508);
and U1251 (N_1251,N_178,N_177);
or U1252 (N_1252,N_448,N_12);
or U1253 (N_1253,N_61,N_932);
or U1254 (N_1254,N_54,N_402);
nand U1255 (N_1255,N_592,N_770);
and U1256 (N_1256,N_113,N_628);
nand U1257 (N_1257,N_619,N_899);
or U1258 (N_1258,N_139,N_622);
or U1259 (N_1259,N_354,N_528);
nor U1260 (N_1260,N_391,N_50);
and U1261 (N_1261,N_954,N_305);
nor U1262 (N_1262,N_604,N_595);
nor U1263 (N_1263,N_24,N_539);
or U1264 (N_1264,N_398,N_726);
or U1265 (N_1265,N_792,N_25);
nand U1266 (N_1266,N_225,N_271);
nor U1267 (N_1267,N_830,N_814);
nor U1268 (N_1268,N_997,N_269);
or U1269 (N_1269,N_224,N_381);
nor U1270 (N_1270,N_260,N_563);
nor U1271 (N_1271,N_11,N_130);
or U1272 (N_1272,N_220,N_279);
and U1273 (N_1273,N_636,N_845);
nand U1274 (N_1274,N_206,N_428);
nor U1275 (N_1275,N_196,N_164);
and U1276 (N_1276,N_60,N_691);
and U1277 (N_1277,N_568,N_939);
nand U1278 (N_1278,N_256,N_694);
and U1279 (N_1279,N_439,N_503);
and U1280 (N_1280,N_740,N_317);
nand U1281 (N_1281,N_352,N_630);
or U1282 (N_1282,N_213,N_338);
nand U1283 (N_1283,N_184,N_935);
nand U1284 (N_1284,N_951,N_583);
nor U1285 (N_1285,N_534,N_229);
nor U1286 (N_1286,N_19,N_672);
and U1287 (N_1287,N_473,N_621);
nor U1288 (N_1288,N_809,N_609);
nand U1289 (N_1289,N_942,N_58);
and U1290 (N_1290,N_494,N_409);
nand U1291 (N_1291,N_755,N_649);
and U1292 (N_1292,N_699,N_678);
or U1293 (N_1293,N_210,N_88);
nand U1294 (N_1294,N_126,N_433);
xnor U1295 (N_1295,N_791,N_124);
nor U1296 (N_1296,N_612,N_995);
and U1297 (N_1297,N_695,N_710);
or U1298 (N_1298,N_288,N_430);
nand U1299 (N_1299,N_804,N_283);
and U1300 (N_1300,N_689,N_310);
nor U1301 (N_1301,N_905,N_267);
nor U1302 (N_1302,N_859,N_960);
nor U1303 (N_1303,N_838,N_575);
or U1304 (N_1304,N_631,N_45);
and U1305 (N_1305,N_634,N_257);
and U1306 (N_1306,N_401,N_613);
nor U1307 (N_1307,N_146,N_156);
nand U1308 (N_1308,N_458,N_650);
nand U1309 (N_1309,N_154,N_70);
nor U1310 (N_1310,N_303,N_748);
or U1311 (N_1311,N_990,N_277);
nand U1312 (N_1312,N_138,N_493);
nand U1313 (N_1313,N_738,N_236);
nand U1314 (N_1314,N_652,N_981);
or U1315 (N_1315,N_480,N_886);
nor U1316 (N_1316,N_958,N_266);
and U1317 (N_1317,N_484,N_529);
nor U1318 (N_1318,N_131,N_569);
or U1319 (N_1319,N_829,N_378);
and U1320 (N_1320,N_558,N_449);
nand U1321 (N_1321,N_606,N_700);
and U1322 (N_1322,N_464,N_803);
xor U1323 (N_1323,N_185,N_199);
nand U1324 (N_1324,N_980,N_788);
or U1325 (N_1325,N_63,N_917);
or U1326 (N_1326,N_625,N_891);
nor U1327 (N_1327,N_671,N_978);
nor U1328 (N_1328,N_286,N_250);
nor U1329 (N_1329,N_546,N_881);
and U1330 (N_1330,N_638,N_294);
nor U1331 (N_1331,N_481,N_153);
or U1332 (N_1332,N_86,N_172);
nor U1333 (N_1333,N_380,N_866);
and U1334 (N_1334,N_707,N_5);
nor U1335 (N_1335,N_876,N_238);
nand U1336 (N_1336,N_437,N_320);
or U1337 (N_1337,N_624,N_344);
xor U1338 (N_1338,N_326,N_461);
nor U1339 (N_1339,N_234,N_643);
nor U1340 (N_1340,N_987,N_476);
nand U1341 (N_1341,N_456,N_296);
or U1342 (N_1342,N_549,N_889);
or U1343 (N_1343,N_902,N_142);
nand U1344 (N_1344,N_330,N_869);
nor U1345 (N_1345,N_351,N_149);
nand U1346 (N_1346,N_832,N_365);
and U1347 (N_1347,N_312,N_527);
nand U1348 (N_1348,N_434,N_925);
and U1349 (N_1349,N_543,N_475);
and U1350 (N_1350,N_487,N_416);
nand U1351 (N_1351,N_474,N_123);
nand U1352 (N_1352,N_328,N_176);
and U1353 (N_1353,N_319,N_423);
and U1354 (N_1354,N_76,N_221);
or U1355 (N_1355,N_66,N_875);
or U1356 (N_1356,N_1,N_514);
and U1357 (N_1357,N_219,N_526);
and U1358 (N_1358,N_226,N_518);
and U1359 (N_1359,N_687,N_840);
and U1360 (N_1360,N_884,N_552);
nand U1361 (N_1361,N_440,N_615);
and U1362 (N_1362,N_910,N_232);
and U1363 (N_1363,N_861,N_435);
and U1364 (N_1364,N_115,N_244);
and U1365 (N_1365,N_208,N_293);
and U1366 (N_1366,N_463,N_666);
nor U1367 (N_1367,N_833,N_588);
nand U1368 (N_1368,N_868,N_289);
xnor U1369 (N_1369,N_871,N_482);
or U1370 (N_1370,N_262,N_835);
and U1371 (N_1371,N_441,N_450);
nor U1372 (N_1372,N_491,N_285);
nand U1373 (N_1373,N_882,N_228);
or U1374 (N_1374,N_412,N_28);
and U1375 (N_1375,N_500,N_919);
and U1376 (N_1376,N_888,N_227);
nand U1377 (N_1377,N_602,N_315);
nand U1378 (N_1378,N_633,N_655);
nor U1379 (N_1379,N_207,N_119);
and U1380 (N_1380,N_444,N_972);
nor U1381 (N_1381,N_383,N_906);
and U1382 (N_1382,N_404,N_920);
nand U1383 (N_1383,N_48,N_222);
nor U1384 (N_1384,N_535,N_421);
nand U1385 (N_1385,N_733,N_52);
nand U1386 (N_1386,N_856,N_947);
or U1387 (N_1387,N_264,N_498);
nor U1388 (N_1388,N_572,N_570);
or U1389 (N_1389,N_637,N_775);
nand U1390 (N_1390,N_697,N_462);
and U1391 (N_1391,N_532,N_23);
nand U1392 (N_1392,N_194,N_506);
or U1393 (N_1393,N_915,N_171);
or U1394 (N_1394,N_561,N_43);
nor U1395 (N_1395,N_580,N_663);
and U1396 (N_1396,N_846,N_181);
nand U1397 (N_1397,N_654,N_586);
nor U1398 (N_1398,N_55,N_515);
and U1399 (N_1399,N_782,N_99);
nor U1400 (N_1400,N_600,N_492);
and U1401 (N_1401,N_737,N_341);
nor U1402 (N_1402,N_158,N_911);
or U1403 (N_1403,N_548,N_994);
nor U1404 (N_1404,N_71,N_342);
nand U1405 (N_1405,N_357,N_708);
nor U1406 (N_1406,N_542,N_741);
nor U1407 (N_1407,N_962,N_195);
nand U1408 (N_1408,N_282,N_608);
nand U1409 (N_1409,N_806,N_587);
nand U1410 (N_1410,N_605,N_657);
nor U1411 (N_1411,N_108,N_424);
or U1412 (N_1412,N_74,N_118);
or U1413 (N_1413,N_418,N_779);
or U1414 (N_1414,N_719,N_263);
and U1415 (N_1415,N_577,N_670);
nand U1416 (N_1416,N_620,N_822);
or U1417 (N_1417,N_445,N_143);
nor U1418 (N_1418,N_362,N_821);
nor U1419 (N_1419,N_931,N_4);
nand U1420 (N_1420,N_10,N_812);
and U1421 (N_1421,N_992,N_754);
xnor U1422 (N_1422,N_496,N_432);
nand U1423 (N_1423,N_996,N_53);
or U1424 (N_1424,N_601,N_46);
and U1425 (N_1425,N_794,N_904);
and U1426 (N_1426,N_337,N_793);
nor U1427 (N_1427,N_799,N_472);
or U1428 (N_1428,N_584,N_751);
or U1429 (N_1429,N_30,N_93);
or U1430 (N_1430,N_802,N_355);
and U1431 (N_1431,N_129,N_62);
nor U1432 (N_1432,N_29,N_952);
and U1433 (N_1433,N_203,N_270);
nand U1434 (N_1434,N_704,N_728);
or U1435 (N_1435,N_175,N_742);
nand U1436 (N_1436,N_762,N_372);
nand U1437 (N_1437,N_230,N_332);
or U1438 (N_1438,N_903,N_850);
and U1439 (N_1439,N_520,N_772);
and U1440 (N_1440,N_128,N_729);
or U1441 (N_1441,N_394,N_235);
and U1442 (N_1442,N_676,N_489);
nand U1443 (N_1443,N_957,N_970);
or U1444 (N_1444,N_926,N_166);
or U1445 (N_1445,N_47,N_573);
nand U1446 (N_1446,N_537,N_7);
and U1447 (N_1447,N_205,N_336);
or U1448 (N_1448,N_291,N_446);
nand U1449 (N_1449,N_276,N_384);
and U1450 (N_1450,N_968,N_879);
nand U1451 (N_1451,N_853,N_522);
nor U1452 (N_1452,N_679,N_736);
and U1453 (N_1453,N_966,N_308);
nor U1454 (N_1454,N_749,N_251);
or U1455 (N_1455,N_366,N_816);
or U1456 (N_1456,N_400,N_133);
nand U1457 (N_1457,N_725,N_96);
or U1458 (N_1458,N_387,N_465);
nor U1459 (N_1459,N_576,N_824);
or U1460 (N_1460,N_787,N_693);
and U1461 (N_1461,N_89,N_541);
nor U1462 (N_1462,N_977,N_106);
nand U1463 (N_1463,N_367,N_408);
or U1464 (N_1464,N_892,N_567);
and U1465 (N_1465,N_826,N_102);
nor U1466 (N_1466,N_712,N_786);
nand U1467 (N_1467,N_422,N_924);
or U1468 (N_1468,N_819,N_817);
or U1469 (N_1469,N_934,N_212);
and U1470 (N_1470,N_959,N_209);
nor U1471 (N_1471,N_927,N_211);
and U1472 (N_1472,N_798,N_84);
and U1473 (N_1473,N_660,N_949);
and U1474 (N_1474,N_284,N_325);
nand U1475 (N_1475,N_246,N_168);
nand U1476 (N_1476,N_41,N_278);
nor U1477 (N_1477,N_140,N_635);
and U1478 (N_1478,N_162,N_967);
nor U1479 (N_1479,N_419,N_673);
nor U1480 (N_1480,N_345,N_502);
nand U1481 (N_1481,N_785,N_57);
and U1482 (N_1482,N_677,N_110);
and U1483 (N_1483,N_590,N_757);
and U1484 (N_1484,N_585,N_578);
nand U1485 (N_1485,N_984,N_186);
and U1486 (N_1486,N_651,N_249);
nand U1487 (N_1487,N_731,N_692);
nor U1488 (N_1488,N_65,N_69);
nand U1489 (N_1489,N_15,N_985);
nand U1490 (N_1490,N_109,N_933);
nor U1491 (N_1491,N_750,N_77);
nor U1492 (N_1492,N_763,N_103);
or U1493 (N_1493,N_684,N_964);
and U1494 (N_1494,N_44,N_92);
xnor U1495 (N_1495,N_744,N_895);
xor U1496 (N_1496,N_290,N_9);
nand U1497 (N_1497,N_295,N_571);
or U1498 (N_1498,N_825,N_632);
nand U1499 (N_1499,N_59,N_304);
or U1500 (N_1500,N_0,N_742);
or U1501 (N_1501,N_577,N_159);
or U1502 (N_1502,N_863,N_368);
nand U1503 (N_1503,N_663,N_192);
or U1504 (N_1504,N_553,N_286);
xor U1505 (N_1505,N_828,N_532);
or U1506 (N_1506,N_691,N_358);
and U1507 (N_1507,N_882,N_566);
or U1508 (N_1508,N_56,N_795);
and U1509 (N_1509,N_695,N_918);
or U1510 (N_1510,N_907,N_192);
and U1511 (N_1511,N_698,N_445);
or U1512 (N_1512,N_146,N_912);
or U1513 (N_1513,N_869,N_883);
or U1514 (N_1514,N_768,N_154);
or U1515 (N_1515,N_811,N_688);
nand U1516 (N_1516,N_731,N_736);
nor U1517 (N_1517,N_200,N_992);
nand U1518 (N_1518,N_664,N_667);
nand U1519 (N_1519,N_110,N_980);
or U1520 (N_1520,N_853,N_237);
nand U1521 (N_1521,N_103,N_618);
nor U1522 (N_1522,N_109,N_216);
or U1523 (N_1523,N_508,N_291);
and U1524 (N_1524,N_562,N_233);
nor U1525 (N_1525,N_221,N_878);
nor U1526 (N_1526,N_81,N_754);
or U1527 (N_1527,N_291,N_303);
xor U1528 (N_1528,N_162,N_140);
and U1529 (N_1529,N_153,N_999);
and U1530 (N_1530,N_50,N_153);
and U1531 (N_1531,N_362,N_418);
nor U1532 (N_1532,N_40,N_938);
nor U1533 (N_1533,N_365,N_56);
and U1534 (N_1534,N_421,N_332);
nor U1535 (N_1535,N_353,N_958);
or U1536 (N_1536,N_288,N_735);
and U1537 (N_1537,N_471,N_828);
or U1538 (N_1538,N_908,N_421);
and U1539 (N_1539,N_454,N_458);
and U1540 (N_1540,N_663,N_882);
or U1541 (N_1541,N_475,N_101);
nor U1542 (N_1542,N_798,N_406);
nand U1543 (N_1543,N_292,N_623);
nand U1544 (N_1544,N_878,N_219);
nor U1545 (N_1545,N_777,N_891);
nand U1546 (N_1546,N_702,N_41);
and U1547 (N_1547,N_395,N_721);
and U1548 (N_1548,N_449,N_798);
or U1549 (N_1549,N_269,N_232);
and U1550 (N_1550,N_536,N_611);
or U1551 (N_1551,N_499,N_736);
nand U1552 (N_1552,N_443,N_331);
and U1553 (N_1553,N_921,N_679);
and U1554 (N_1554,N_752,N_776);
nand U1555 (N_1555,N_354,N_747);
nand U1556 (N_1556,N_505,N_155);
nor U1557 (N_1557,N_469,N_51);
nor U1558 (N_1558,N_706,N_329);
or U1559 (N_1559,N_650,N_834);
nor U1560 (N_1560,N_929,N_962);
nor U1561 (N_1561,N_572,N_630);
or U1562 (N_1562,N_915,N_970);
nand U1563 (N_1563,N_677,N_439);
and U1564 (N_1564,N_634,N_349);
and U1565 (N_1565,N_172,N_954);
or U1566 (N_1566,N_839,N_730);
and U1567 (N_1567,N_78,N_330);
or U1568 (N_1568,N_995,N_172);
xor U1569 (N_1569,N_440,N_920);
nor U1570 (N_1570,N_756,N_832);
nand U1571 (N_1571,N_346,N_338);
nor U1572 (N_1572,N_166,N_947);
or U1573 (N_1573,N_409,N_935);
and U1574 (N_1574,N_89,N_606);
nand U1575 (N_1575,N_598,N_138);
xnor U1576 (N_1576,N_165,N_282);
nand U1577 (N_1577,N_629,N_345);
or U1578 (N_1578,N_866,N_186);
or U1579 (N_1579,N_987,N_337);
or U1580 (N_1580,N_807,N_840);
nand U1581 (N_1581,N_465,N_270);
or U1582 (N_1582,N_581,N_141);
nand U1583 (N_1583,N_520,N_32);
and U1584 (N_1584,N_911,N_738);
or U1585 (N_1585,N_736,N_220);
or U1586 (N_1586,N_973,N_415);
xor U1587 (N_1587,N_652,N_360);
or U1588 (N_1588,N_718,N_723);
nand U1589 (N_1589,N_427,N_273);
nand U1590 (N_1590,N_186,N_870);
nand U1591 (N_1591,N_325,N_75);
nand U1592 (N_1592,N_357,N_33);
nand U1593 (N_1593,N_405,N_347);
nand U1594 (N_1594,N_841,N_566);
nor U1595 (N_1595,N_801,N_847);
or U1596 (N_1596,N_18,N_164);
nand U1597 (N_1597,N_674,N_292);
nor U1598 (N_1598,N_997,N_84);
and U1599 (N_1599,N_870,N_201);
or U1600 (N_1600,N_220,N_408);
nand U1601 (N_1601,N_916,N_332);
nor U1602 (N_1602,N_847,N_515);
or U1603 (N_1603,N_695,N_172);
nor U1604 (N_1604,N_287,N_258);
and U1605 (N_1605,N_454,N_938);
and U1606 (N_1606,N_734,N_288);
nor U1607 (N_1607,N_766,N_483);
and U1608 (N_1608,N_714,N_324);
and U1609 (N_1609,N_744,N_243);
xnor U1610 (N_1610,N_724,N_728);
xnor U1611 (N_1611,N_39,N_682);
or U1612 (N_1612,N_855,N_454);
nor U1613 (N_1613,N_678,N_123);
or U1614 (N_1614,N_998,N_851);
nand U1615 (N_1615,N_473,N_876);
nor U1616 (N_1616,N_209,N_4);
and U1617 (N_1617,N_568,N_323);
xnor U1618 (N_1618,N_50,N_394);
or U1619 (N_1619,N_342,N_355);
nor U1620 (N_1620,N_28,N_244);
or U1621 (N_1621,N_856,N_961);
nor U1622 (N_1622,N_440,N_888);
nor U1623 (N_1623,N_909,N_487);
and U1624 (N_1624,N_675,N_621);
nor U1625 (N_1625,N_260,N_919);
and U1626 (N_1626,N_844,N_691);
nor U1627 (N_1627,N_501,N_363);
nor U1628 (N_1628,N_891,N_138);
and U1629 (N_1629,N_677,N_873);
nand U1630 (N_1630,N_852,N_633);
nor U1631 (N_1631,N_119,N_213);
or U1632 (N_1632,N_876,N_524);
or U1633 (N_1633,N_670,N_253);
nor U1634 (N_1634,N_75,N_63);
nor U1635 (N_1635,N_780,N_361);
or U1636 (N_1636,N_113,N_306);
nor U1637 (N_1637,N_815,N_24);
nand U1638 (N_1638,N_233,N_136);
nor U1639 (N_1639,N_362,N_135);
nor U1640 (N_1640,N_826,N_939);
nor U1641 (N_1641,N_904,N_546);
or U1642 (N_1642,N_486,N_95);
nand U1643 (N_1643,N_876,N_89);
and U1644 (N_1644,N_185,N_807);
nor U1645 (N_1645,N_35,N_381);
and U1646 (N_1646,N_120,N_938);
nor U1647 (N_1647,N_502,N_934);
and U1648 (N_1648,N_419,N_472);
nor U1649 (N_1649,N_41,N_151);
nor U1650 (N_1650,N_460,N_21);
or U1651 (N_1651,N_618,N_951);
or U1652 (N_1652,N_385,N_221);
nand U1653 (N_1653,N_467,N_938);
nor U1654 (N_1654,N_723,N_191);
nand U1655 (N_1655,N_187,N_401);
nand U1656 (N_1656,N_786,N_919);
or U1657 (N_1657,N_984,N_996);
nor U1658 (N_1658,N_51,N_905);
nand U1659 (N_1659,N_86,N_650);
nor U1660 (N_1660,N_343,N_824);
nor U1661 (N_1661,N_280,N_902);
and U1662 (N_1662,N_193,N_391);
nor U1663 (N_1663,N_545,N_613);
nor U1664 (N_1664,N_495,N_876);
and U1665 (N_1665,N_98,N_457);
nor U1666 (N_1666,N_699,N_22);
nor U1667 (N_1667,N_415,N_876);
nor U1668 (N_1668,N_664,N_366);
nor U1669 (N_1669,N_120,N_140);
or U1670 (N_1670,N_966,N_366);
nor U1671 (N_1671,N_387,N_675);
nor U1672 (N_1672,N_944,N_977);
or U1673 (N_1673,N_78,N_766);
and U1674 (N_1674,N_433,N_257);
nand U1675 (N_1675,N_837,N_672);
and U1676 (N_1676,N_966,N_755);
xnor U1677 (N_1677,N_691,N_184);
and U1678 (N_1678,N_228,N_436);
or U1679 (N_1679,N_273,N_895);
nand U1680 (N_1680,N_47,N_605);
and U1681 (N_1681,N_875,N_622);
nand U1682 (N_1682,N_502,N_627);
or U1683 (N_1683,N_135,N_67);
and U1684 (N_1684,N_793,N_596);
or U1685 (N_1685,N_507,N_428);
and U1686 (N_1686,N_680,N_317);
nor U1687 (N_1687,N_942,N_315);
and U1688 (N_1688,N_279,N_396);
nand U1689 (N_1689,N_155,N_674);
nand U1690 (N_1690,N_300,N_458);
and U1691 (N_1691,N_422,N_160);
or U1692 (N_1692,N_129,N_323);
nand U1693 (N_1693,N_970,N_481);
and U1694 (N_1694,N_82,N_30);
nor U1695 (N_1695,N_402,N_666);
nand U1696 (N_1696,N_194,N_525);
or U1697 (N_1697,N_938,N_512);
or U1698 (N_1698,N_580,N_290);
and U1699 (N_1699,N_94,N_186);
and U1700 (N_1700,N_302,N_980);
or U1701 (N_1701,N_621,N_645);
nand U1702 (N_1702,N_382,N_529);
and U1703 (N_1703,N_634,N_110);
or U1704 (N_1704,N_741,N_209);
and U1705 (N_1705,N_607,N_414);
or U1706 (N_1706,N_695,N_859);
or U1707 (N_1707,N_16,N_825);
nor U1708 (N_1708,N_24,N_148);
nand U1709 (N_1709,N_512,N_694);
or U1710 (N_1710,N_35,N_585);
nand U1711 (N_1711,N_166,N_869);
and U1712 (N_1712,N_126,N_848);
nor U1713 (N_1713,N_933,N_728);
or U1714 (N_1714,N_309,N_913);
nor U1715 (N_1715,N_380,N_443);
and U1716 (N_1716,N_363,N_916);
and U1717 (N_1717,N_197,N_574);
and U1718 (N_1718,N_902,N_806);
and U1719 (N_1719,N_108,N_214);
nor U1720 (N_1720,N_538,N_255);
or U1721 (N_1721,N_165,N_686);
nand U1722 (N_1722,N_68,N_90);
and U1723 (N_1723,N_738,N_862);
and U1724 (N_1724,N_700,N_665);
nand U1725 (N_1725,N_415,N_733);
nor U1726 (N_1726,N_922,N_401);
nand U1727 (N_1727,N_100,N_221);
and U1728 (N_1728,N_559,N_953);
nor U1729 (N_1729,N_561,N_714);
nand U1730 (N_1730,N_496,N_973);
nor U1731 (N_1731,N_940,N_3);
or U1732 (N_1732,N_993,N_883);
nor U1733 (N_1733,N_879,N_142);
and U1734 (N_1734,N_482,N_546);
nor U1735 (N_1735,N_288,N_870);
or U1736 (N_1736,N_121,N_379);
xnor U1737 (N_1737,N_52,N_289);
nor U1738 (N_1738,N_775,N_79);
nor U1739 (N_1739,N_259,N_526);
and U1740 (N_1740,N_630,N_714);
nand U1741 (N_1741,N_784,N_94);
and U1742 (N_1742,N_531,N_551);
or U1743 (N_1743,N_7,N_742);
and U1744 (N_1744,N_303,N_23);
or U1745 (N_1745,N_530,N_756);
xnor U1746 (N_1746,N_669,N_843);
nand U1747 (N_1747,N_386,N_815);
or U1748 (N_1748,N_250,N_46);
or U1749 (N_1749,N_523,N_186);
nor U1750 (N_1750,N_809,N_371);
nand U1751 (N_1751,N_382,N_690);
nor U1752 (N_1752,N_322,N_854);
and U1753 (N_1753,N_154,N_949);
nand U1754 (N_1754,N_358,N_318);
nand U1755 (N_1755,N_988,N_547);
and U1756 (N_1756,N_792,N_762);
or U1757 (N_1757,N_351,N_260);
or U1758 (N_1758,N_960,N_920);
nor U1759 (N_1759,N_720,N_647);
nand U1760 (N_1760,N_43,N_113);
or U1761 (N_1761,N_670,N_800);
nor U1762 (N_1762,N_91,N_352);
nand U1763 (N_1763,N_157,N_286);
or U1764 (N_1764,N_321,N_746);
nand U1765 (N_1765,N_611,N_399);
or U1766 (N_1766,N_351,N_837);
nor U1767 (N_1767,N_486,N_363);
or U1768 (N_1768,N_580,N_164);
nand U1769 (N_1769,N_189,N_844);
and U1770 (N_1770,N_849,N_62);
and U1771 (N_1771,N_167,N_544);
xor U1772 (N_1772,N_783,N_329);
nor U1773 (N_1773,N_504,N_681);
nor U1774 (N_1774,N_730,N_903);
and U1775 (N_1775,N_711,N_13);
nand U1776 (N_1776,N_319,N_246);
nand U1777 (N_1777,N_312,N_400);
nor U1778 (N_1778,N_457,N_422);
nand U1779 (N_1779,N_51,N_610);
nor U1780 (N_1780,N_709,N_503);
nand U1781 (N_1781,N_555,N_508);
or U1782 (N_1782,N_649,N_367);
xnor U1783 (N_1783,N_287,N_71);
or U1784 (N_1784,N_629,N_321);
nand U1785 (N_1785,N_25,N_135);
nor U1786 (N_1786,N_531,N_102);
nor U1787 (N_1787,N_974,N_388);
nand U1788 (N_1788,N_120,N_825);
and U1789 (N_1789,N_647,N_223);
nand U1790 (N_1790,N_706,N_551);
nand U1791 (N_1791,N_770,N_900);
nand U1792 (N_1792,N_932,N_562);
or U1793 (N_1793,N_341,N_587);
and U1794 (N_1794,N_273,N_488);
and U1795 (N_1795,N_457,N_211);
or U1796 (N_1796,N_793,N_171);
and U1797 (N_1797,N_990,N_339);
xor U1798 (N_1798,N_748,N_424);
or U1799 (N_1799,N_835,N_995);
and U1800 (N_1800,N_486,N_992);
and U1801 (N_1801,N_801,N_468);
nor U1802 (N_1802,N_209,N_700);
and U1803 (N_1803,N_791,N_723);
or U1804 (N_1804,N_197,N_140);
xnor U1805 (N_1805,N_814,N_589);
nand U1806 (N_1806,N_508,N_78);
and U1807 (N_1807,N_704,N_463);
nor U1808 (N_1808,N_752,N_575);
nand U1809 (N_1809,N_431,N_724);
nand U1810 (N_1810,N_956,N_38);
nor U1811 (N_1811,N_279,N_836);
nor U1812 (N_1812,N_937,N_483);
xnor U1813 (N_1813,N_968,N_728);
xor U1814 (N_1814,N_469,N_509);
and U1815 (N_1815,N_402,N_56);
or U1816 (N_1816,N_713,N_220);
and U1817 (N_1817,N_852,N_39);
nor U1818 (N_1818,N_577,N_573);
nor U1819 (N_1819,N_794,N_742);
nand U1820 (N_1820,N_490,N_932);
and U1821 (N_1821,N_80,N_592);
and U1822 (N_1822,N_951,N_35);
nor U1823 (N_1823,N_469,N_802);
or U1824 (N_1824,N_359,N_110);
and U1825 (N_1825,N_782,N_916);
xnor U1826 (N_1826,N_918,N_6);
nor U1827 (N_1827,N_931,N_124);
or U1828 (N_1828,N_236,N_647);
and U1829 (N_1829,N_728,N_921);
nand U1830 (N_1830,N_513,N_568);
and U1831 (N_1831,N_77,N_956);
and U1832 (N_1832,N_555,N_133);
nor U1833 (N_1833,N_444,N_726);
nor U1834 (N_1834,N_499,N_448);
nand U1835 (N_1835,N_502,N_556);
or U1836 (N_1836,N_443,N_344);
and U1837 (N_1837,N_103,N_65);
and U1838 (N_1838,N_611,N_722);
or U1839 (N_1839,N_260,N_75);
nor U1840 (N_1840,N_151,N_536);
or U1841 (N_1841,N_638,N_921);
nor U1842 (N_1842,N_67,N_315);
nor U1843 (N_1843,N_67,N_473);
nand U1844 (N_1844,N_404,N_467);
nor U1845 (N_1845,N_676,N_213);
and U1846 (N_1846,N_668,N_979);
nand U1847 (N_1847,N_43,N_592);
and U1848 (N_1848,N_717,N_636);
nor U1849 (N_1849,N_589,N_712);
xnor U1850 (N_1850,N_499,N_733);
or U1851 (N_1851,N_802,N_12);
or U1852 (N_1852,N_942,N_625);
xnor U1853 (N_1853,N_996,N_861);
and U1854 (N_1854,N_676,N_186);
nand U1855 (N_1855,N_707,N_407);
nor U1856 (N_1856,N_744,N_757);
or U1857 (N_1857,N_255,N_9);
and U1858 (N_1858,N_288,N_356);
and U1859 (N_1859,N_529,N_784);
nand U1860 (N_1860,N_446,N_470);
nor U1861 (N_1861,N_490,N_94);
nor U1862 (N_1862,N_827,N_536);
nand U1863 (N_1863,N_41,N_54);
nand U1864 (N_1864,N_899,N_340);
and U1865 (N_1865,N_376,N_13);
or U1866 (N_1866,N_918,N_131);
nor U1867 (N_1867,N_115,N_868);
nor U1868 (N_1868,N_500,N_287);
or U1869 (N_1869,N_276,N_620);
nor U1870 (N_1870,N_168,N_92);
nand U1871 (N_1871,N_866,N_953);
nand U1872 (N_1872,N_537,N_856);
nor U1873 (N_1873,N_890,N_472);
nor U1874 (N_1874,N_380,N_35);
nor U1875 (N_1875,N_963,N_339);
nor U1876 (N_1876,N_83,N_954);
or U1877 (N_1877,N_186,N_906);
nor U1878 (N_1878,N_738,N_756);
and U1879 (N_1879,N_989,N_558);
and U1880 (N_1880,N_705,N_508);
nand U1881 (N_1881,N_155,N_223);
nor U1882 (N_1882,N_405,N_462);
nor U1883 (N_1883,N_679,N_419);
and U1884 (N_1884,N_845,N_152);
xnor U1885 (N_1885,N_741,N_472);
or U1886 (N_1886,N_135,N_578);
or U1887 (N_1887,N_91,N_156);
and U1888 (N_1888,N_247,N_552);
or U1889 (N_1889,N_251,N_996);
or U1890 (N_1890,N_923,N_259);
and U1891 (N_1891,N_731,N_241);
nor U1892 (N_1892,N_131,N_445);
nand U1893 (N_1893,N_461,N_186);
and U1894 (N_1894,N_868,N_300);
or U1895 (N_1895,N_951,N_8);
nand U1896 (N_1896,N_340,N_327);
xnor U1897 (N_1897,N_603,N_868);
nand U1898 (N_1898,N_251,N_519);
or U1899 (N_1899,N_858,N_871);
nor U1900 (N_1900,N_268,N_470);
nor U1901 (N_1901,N_833,N_318);
nand U1902 (N_1902,N_681,N_238);
nor U1903 (N_1903,N_468,N_235);
nand U1904 (N_1904,N_260,N_47);
and U1905 (N_1905,N_396,N_294);
or U1906 (N_1906,N_618,N_701);
or U1907 (N_1907,N_479,N_574);
xor U1908 (N_1908,N_19,N_663);
nand U1909 (N_1909,N_671,N_145);
or U1910 (N_1910,N_113,N_86);
nor U1911 (N_1911,N_128,N_59);
nor U1912 (N_1912,N_816,N_775);
and U1913 (N_1913,N_204,N_976);
or U1914 (N_1914,N_593,N_332);
or U1915 (N_1915,N_337,N_878);
nand U1916 (N_1916,N_525,N_928);
or U1917 (N_1917,N_68,N_784);
and U1918 (N_1918,N_597,N_692);
nor U1919 (N_1919,N_598,N_761);
or U1920 (N_1920,N_477,N_287);
nand U1921 (N_1921,N_115,N_999);
and U1922 (N_1922,N_885,N_494);
nand U1923 (N_1923,N_958,N_114);
or U1924 (N_1924,N_209,N_494);
nor U1925 (N_1925,N_25,N_84);
or U1926 (N_1926,N_511,N_887);
nand U1927 (N_1927,N_465,N_5);
and U1928 (N_1928,N_955,N_488);
and U1929 (N_1929,N_863,N_553);
nor U1930 (N_1930,N_520,N_41);
nand U1931 (N_1931,N_48,N_950);
nor U1932 (N_1932,N_77,N_766);
or U1933 (N_1933,N_759,N_290);
or U1934 (N_1934,N_49,N_399);
or U1935 (N_1935,N_476,N_602);
and U1936 (N_1936,N_829,N_960);
nand U1937 (N_1937,N_418,N_367);
nor U1938 (N_1938,N_990,N_994);
nand U1939 (N_1939,N_917,N_918);
nand U1940 (N_1940,N_458,N_849);
or U1941 (N_1941,N_905,N_716);
nand U1942 (N_1942,N_205,N_462);
or U1943 (N_1943,N_846,N_561);
nand U1944 (N_1944,N_741,N_312);
and U1945 (N_1945,N_803,N_53);
nand U1946 (N_1946,N_209,N_311);
nor U1947 (N_1947,N_526,N_346);
or U1948 (N_1948,N_958,N_145);
nand U1949 (N_1949,N_871,N_468);
and U1950 (N_1950,N_512,N_666);
or U1951 (N_1951,N_731,N_935);
and U1952 (N_1952,N_82,N_845);
and U1953 (N_1953,N_475,N_637);
and U1954 (N_1954,N_248,N_26);
or U1955 (N_1955,N_445,N_201);
xnor U1956 (N_1956,N_458,N_671);
and U1957 (N_1957,N_481,N_244);
or U1958 (N_1958,N_559,N_263);
and U1959 (N_1959,N_538,N_751);
or U1960 (N_1960,N_358,N_807);
nand U1961 (N_1961,N_337,N_629);
nand U1962 (N_1962,N_916,N_794);
xnor U1963 (N_1963,N_77,N_858);
or U1964 (N_1964,N_445,N_58);
nor U1965 (N_1965,N_72,N_118);
or U1966 (N_1966,N_559,N_751);
and U1967 (N_1967,N_587,N_477);
nor U1968 (N_1968,N_799,N_757);
nand U1969 (N_1969,N_270,N_67);
and U1970 (N_1970,N_328,N_930);
nand U1971 (N_1971,N_739,N_669);
nor U1972 (N_1972,N_650,N_773);
nor U1973 (N_1973,N_166,N_547);
nor U1974 (N_1974,N_586,N_436);
xnor U1975 (N_1975,N_139,N_226);
nor U1976 (N_1976,N_484,N_599);
or U1977 (N_1977,N_194,N_554);
and U1978 (N_1978,N_71,N_384);
or U1979 (N_1979,N_609,N_489);
nand U1980 (N_1980,N_382,N_662);
and U1981 (N_1981,N_656,N_25);
nor U1982 (N_1982,N_445,N_125);
and U1983 (N_1983,N_875,N_578);
and U1984 (N_1984,N_58,N_945);
or U1985 (N_1985,N_103,N_479);
nor U1986 (N_1986,N_601,N_436);
and U1987 (N_1987,N_124,N_223);
nor U1988 (N_1988,N_139,N_447);
and U1989 (N_1989,N_499,N_741);
nand U1990 (N_1990,N_744,N_636);
nor U1991 (N_1991,N_897,N_581);
nand U1992 (N_1992,N_297,N_137);
and U1993 (N_1993,N_983,N_687);
and U1994 (N_1994,N_839,N_809);
nand U1995 (N_1995,N_436,N_939);
or U1996 (N_1996,N_710,N_793);
nand U1997 (N_1997,N_989,N_571);
nand U1998 (N_1998,N_350,N_248);
or U1999 (N_1999,N_823,N_557);
nor U2000 (N_2000,N_1116,N_1813);
nor U2001 (N_2001,N_1866,N_1869);
or U2002 (N_2002,N_1946,N_1243);
nand U2003 (N_2003,N_1912,N_1321);
nand U2004 (N_2004,N_1009,N_1921);
nand U2005 (N_2005,N_1038,N_1470);
and U2006 (N_2006,N_1051,N_1205);
nand U2007 (N_2007,N_1824,N_1212);
nor U2008 (N_2008,N_1443,N_1827);
nand U2009 (N_2009,N_1119,N_1731);
nand U2010 (N_2010,N_1893,N_1623);
and U2011 (N_2011,N_1419,N_1666);
nand U2012 (N_2012,N_1357,N_1907);
and U2013 (N_2013,N_1180,N_1778);
nand U2014 (N_2014,N_1883,N_1988);
nor U2015 (N_2015,N_1717,N_1860);
and U2016 (N_2016,N_1398,N_1642);
and U2017 (N_2017,N_1908,N_1553);
and U2018 (N_2018,N_1071,N_1797);
and U2019 (N_2019,N_1564,N_1895);
nand U2020 (N_2020,N_1575,N_1150);
nor U2021 (N_2021,N_1736,N_1789);
nand U2022 (N_2022,N_1030,N_1591);
or U2023 (N_2023,N_1355,N_1184);
nor U2024 (N_2024,N_1663,N_1632);
and U2025 (N_2025,N_1492,N_1432);
and U2026 (N_2026,N_1236,N_1399);
nand U2027 (N_2027,N_1322,N_1719);
nor U2028 (N_2028,N_1111,N_1724);
and U2029 (N_2029,N_1950,N_1668);
or U2030 (N_2030,N_1889,N_1337);
or U2031 (N_2031,N_1699,N_1783);
nor U2032 (N_2032,N_1753,N_1124);
nor U2033 (N_2033,N_1216,N_1973);
nand U2034 (N_2034,N_1258,N_1605);
and U2035 (N_2035,N_1561,N_1906);
and U2036 (N_2036,N_1147,N_1734);
nor U2037 (N_2037,N_1195,N_1000);
nor U2038 (N_2038,N_1630,N_1655);
nand U2039 (N_2039,N_1132,N_1956);
nor U2040 (N_2040,N_1016,N_1414);
nor U2041 (N_2041,N_1214,N_1841);
and U2042 (N_2042,N_1742,N_1594);
and U2043 (N_2043,N_1615,N_1157);
and U2044 (N_2044,N_1552,N_1968);
or U2045 (N_2045,N_1376,N_1238);
nand U2046 (N_2046,N_1363,N_1217);
nor U2047 (N_2047,N_1385,N_1574);
and U2048 (N_2048,N_1659,N_1382);
nand U2049 (N_2049,N_1146,N_1381);
nand U2050 (N_2050,N_1453,N_1042);
and U2051 (N_2051,N_1580,N_1800);
or U2052 (N_2052,N_1513,N_1681);
nor U2053 (N_2053,N_1602,N_1823);
and U2054 (N_2054,N_1587,N_1577);
nor U2055 (N_2055,N_1662,N_1065);
nor U2056 (N_2056,N_1394,N_1529);
nor U2057 (N_2057,N_1518,N_1137);
or U2058 (N_2058,N_1899,N_1611);
and U2059 (N_2059,N_1250,N_1943);
or U2060 (N_2060,N_1253,N_1418);
nand U2061 (N_2061,N_1035,N_1330);
nor U2062 (N_2062,N_1786,N_1177);
and U2063 (N_2063,N_1245,N_1235);
and U2064 (N_2064,N_1807,N_1215);
nor U2065 (N_2065,N_1557,N_1885);
nor U2066 (N_2066,N_1306,N_1391);
nand U2067 (N_2067,N_1942,N_1339);
nor U2068 (N_2068,N_1311,N_1528);
or U2069 (N_2069,N_1372,N_1417);
nand U2070 (N_2070,N_1340,N_1098);
or U2071 (N_2071,N_1331,N_1095);
nor U2072 (N_2072,N_1343,N_1707);
xor U2073 (N_2073,N_1070,N_1684);
and U2074 (N_2074,N_1074,N_1679);
nand U2075 (N_2075,N_1107,N_1282);
or U2076 (N_2076,N_1750,N_1178);
nor U2077 (N_2077,N_1240,N_1023);
nor U2078 (N_2078,N_1440,N_1791);
nor U2079 (N_2079,N_1650,N_1556);
or U2080 (N_2080,N_1323,N_1901);
and U2081 (N_2081,N_1127,N_1708);
and U2082 (N_2082,N_1859,N_1692);
nor U2083 (N_2083,N_1104,N_1952);
or U2084 (N_2084,N_1006,N_1249);
and U2085 (N_2085,N_1936,N_1752);
nand U2086 (N_2086,N_1677,N_1350);
and U2087 (N_2087,N_1197,N_1795);
nor U2088 (N_2088,N_1631,N_1844);
nor U2089 (N_2089,N_1371,N_1229);
nand U2090 (N_2090,N_1903,N_1945);
or U2091 (N_2091,N_1255,N_1764);
nor U2092 (N_2092,N_1210,N_1272);
nand U2093 (N_2093,N_1838,N_1353);
and U2094 (N_2094,N_1491,N_1486);
nor U2095 (N_2095,N_1846,N_1011);
nand U2096 (N_2096,N_1588,N_1910);
and U2097 (N_2097,N_1967,N_1619);
nor U2098 (N_2098,N_1412,N_1316);
or U2099 (N_2099,N_1980,N_1687);
and U2100 (N_2100,N_1857,N_1896);
and U2101 (N_2101,N_1460,N_1920);
and U2102 (N_2102,N_1268,N_1975);
xor U2103 (N_2103,N_1590,N_1057);
and U2104 (N_2104,N_1077,N_1046);
and U2105 (N_2105,N_1850,N_1209);
xor U2106 (N_2106,N_1652,N_1308);
or U2107 (N_2107,N_1523,N_1179);
or U2108 (N_2108,N_1100,N_1025);
nand U2109 (N_2109,N_1407,N_1505);
nor U2110 (N_2110,N_1054,N_1779);
or U2111 (N_2111,N_1225,N_1913);
and U2112 (N_2112,N_1193,N_1081);
or U2113 (N_2113,N_1291,N_1780);
nor U2114 (N_2114,N_1754,N_1364);
nand U2115 (N_2115,N_1434,N_1113);
nand U2116 (N_2116,N_1140,N_1582);
nand U2117 (N_2117,N_1902,N_1856);
nor U2118 (N_2118,N_1464,N_1482);
nor U2119 (N_2119,N_1325,N_1676);
and U2120 (N_2120,N_1818,N_1252);
nand U2121 (N_2121,N_1320,N_1387);
nor U2122 (N_2122,N_1929,N_1263);
nand U2123 (N_2123,N_1073,N_1360);
and U2124 (N_2124,N_1836,N_1352);
and U2125 (N_2125,N_1114,N_1198);
or U2126 (N_2126,N_1176,N_1947);
or U2127 (N_2127,N_1251,N_1436);
nor U2128 (N_2128,N_1480,N_1785);
nand U2129 (N_2129,N_1925,N_1422);
nor U2130 (N_2130,N_1402,N_1037);
and U2131 (N_2131,N_1772,N_1415);
and U2132 (N_2132,N_1324,N_1390);
or U2133 (N_2133,N_1932,N_1256);
or U2134 (N_2134,N_1775,N_1586);
and U2135 (N_2135,N_1133,N_1917);
nor U2136 (N_2136,N_1284,N_1086);
nand U2137 (N_2137,N_1012,N_1052);
nand U2138 (N_2138,N_1288,N_1115);
or U2139 (N_2139,N_1169,N_1231);
nor U2140 (N_2140,N_1861,N_1622);
nor U2141 (N_2141,N_1832,N_1465);
xnor U2142 (N_2142,N_1093,N_1957);
and U2143 (N_2143,N_1690,N_1682);
nand U2144 (N_2144,N_1366,N_1110);
nand U2145 (N_2145,N_1303,N_1227);
and U2146 (N_2146,N_1468,N_1804);
or U2147 (N_2147,N_1633,N_1516);
and U2148 (N_2148,N_1597,N_1617);
nor U2149 (N_2149,N_1361,N_1842);
and U2150 (N_2150,N_1259,N_1875);
or U2151 (N_2151,N_1021,N_1266);
or U2152 (N_2152,N_1026,N_1641);
nand U2153 (N_2153,N_1928,N_1218);
and U2154 (N_2154,N_1508,N_1232);
or U2155 (N_2155,N_1446,N_1948);
nand U2156 (N_2156,N_1233,N_1884);
nand U2157 (N_2157,N_1442,N_1369);
xnor U2158 (N_2158,N_1413,N_1043);
nand U2159 (N_2159,N_1156,N_1853);
or U2160 (N_2160,N_1301,N_1854);
nand U2161 (N_2161,N_1539,N_1128);
nand U2162 (N_2162,N_1534,N_1858);
and U2163 (N_2163,N_1722,N_1566);
and U2164 (N_2164,N_1526,N_1743);
and U2165 (N_2165,N_1172,N_1739);
and U2166 (N_2166,N_1963,N_1969);
or U2167 (N_2167,N_1520,N_1168);
or U2168 (N_2168,N_1386,N_1976);
nand U2169 (N_2169,N_1773,N_1036);
nor U2170 (N_2170,N_1447,N_1636);
nor U2171 (N_2171,N_1525,N_1423);
or U2172 (N_2172,N_1994,N_1420);
or U2173 (N_2173,N_1267,N_1223);
nand U2174 (N_2174,N_1951,N_1013);
nor U2175 (N_2175,N_1456,N_1608);
and U2176 (N_2176,N_1166,N_1700);
xor U2177 (N_2177,N_1173,N_1709);
or U2178 (N_2178,N_1959,N_1135);
or U2179 (N_2179,N_1297,N_1509);
nor U2180 (N_2180,N_1159,N_1408);
nor U2181 (N_2181,N_1454,N_1714);
nor U2182 (N_2182,N_1444,N_1931);
and U2183 (N_2183,N_1524,N_1735);
or U2184 (N_2184,N_1222,N_1274);
nor U2185 (N_2185,N_1441,N_1938);
nor U2186 (N_2186,N_1723,N_1664);
or U2187 (N_2187,N_1145,N_1658);
and U2188 (N_2188,N_1558,N_1672);
nor U2189 (N_2189,N_1471,N_1033);
nand U2190 (N_2190,N_1892,N_1535);
nand U2191 (N_2191,N_1203,N_1768);
or U2192 (N_2192,N_1260,N_1990);
or U2193 (N_2193,N_1194,N_1985);
nor U2194 (N_2194,N_1759,N_1809);
and U2195 (N_2195,N_1230,N_1003);
or U2196 (N_2196,N_1143,N_1796);
and U2197 (N_2197,N_1733,N_1701);
and U2198 (N_2198,N_1629,N_1091);
or U2199 (N_2199,N_1880,N_1820);
nand U2200 (N_2200,N_1187,N_1351);
nor U2201 (N_2201,N_1439,N_1475);
xnor U2202 (N_2202,N_1315,N_1384);
nand U2203 (N_2203,N_1204,N_1527);
nor U2204 (N_2204,N_1695,N_1897);
or U2205 (N_2205,N_1915,N_1437);
or U2206 (N_2206,N_1181,N_1130);
nor U2207 (N_2207,N_1821,N_1716);
nand U2208 (N_2208,N_1694,N_1751);
or U2209 (N_2209,N_1326,N_1606);
or U2210 (N_2210,N_1469,N_1314);
xor U2211 (N_2211,N_1401,N_1776);
nor U2212 (N_2212,N_1058,N_1817);
and U2213 (N_2213,N_1871,N_1610);
nand U2214 (N_2214,N_1467,N_1448);
nand U2215 (N_2215,N_1109,N_1774);
nand U2216 (N_2216,N_1530,N_1424);
nor U2217 (N_2217,N_1257,N_1822);
nand U2218 (N_2218,N_1691,N_1544);
nor U2219 (N_2219,N_1830,N_1490);
and U2220 (N_2220,N_1649,N_1438);
nand U2221 (N_2221,N_1273,N_1031);
nand U2222 (N_2222,N_1550,N_1312);
or U2223 (N_2223,N_1609,N_1887);
nand U2224 (N_2224,N_1514,N_1923);
and U2225 (N_2225,N_1139,N_1503);
and U2226 (N_2226,N_1992,N_1603);
nor U2227 (N_2227,N_1264,N_1459);
nor U2228 (N_2228,N_1637,N_1092);
nand U2229 (N_2229,N_1890,N_1863);
nand U2230 (N_2230,N_1200,N_1870);
and U2231 (N_2231,N_1955,N_1275);
nand U2232 (N_2232,N_1653,N_1067);
nand U2233 (N_2233,N_1234,N_1262);
nor U2234 (N_2234,N_1290,N_1755);
or U2235 (N_2235,N_1334,N_1082);
nand U2236 (N_2236,N_1494,N_1152);
nor U2237 (N_2237,N_1450,N_1829);
nand U2238 (N_2238,N_1741,N_1329);
nor U2239 (N_2239,N_1981,N_1777);
or U2240 (N_2240,N_1919,N_1122);
and U2241 (N_2241,N_1487,N_1378);
nand U2242 (N_2242,N_1472,N_1872);
or U2243 (N_2243,N_1914,N_1451);
and U2244 (N_2244,N_1247,N_1909);
or U2245 (N_2245,N_1389,N_1004);
nand U2246 (N_2246,N_1474,N_1693);
or U2247 (N_2247,N_1511,N_1626);
nor U2248 (N_2248,N_1346,N_1196);
and U2249 (N_2249,N_1944,N_1961);
nor U2250 (N_2250,N_1121,N_1579);
or U2251 (N_2251,N_1497,N_1295);
and U2252 (N_2252,N_1686,N_1411);
or U2253 (N_2253,N_1965,N_1125);
nor U2254 (N_2254,N_1348,N_1292);
nor U2255 (N_2255,N_1999,N_1485);
nand U2256 (N_2256,N_1349,N_1192);
xor U2257 (N_2257,N_1254,N_1224);
and U2258 (N_2258,N_1241,N_1802);
nor U2259 (N_2259,N_1549,N_1112);
nor U2260 (N_2260,N_1983,N_1085);
nor U2261 (N_2261,N_1601,N_1103);
nor U2262 (N_2262,N_1918,N_1294);
xnor U2263 (N_2263,N_1228,N_1573);
nand U2264 (N_2264,N_1596,N_1495);
nand U2265 (N_2265,N_1812,N_1845);
nand U2266 (N_2266,N_1765,N_1747);
nand U2267 (N_2267,N_1201,N_1015);
and U2268 (N_2268,N_1296,N_1102);
nor U2269 (N_2269,N_1449,N_1770);
nand U2270 (N_2270,N_1834,N_1149);
and U2271 (N_2271,N_1019,N_1718);
and U2272 (N_2272,N_1839,N_1426);
nor U2273 (N_2273,N_1873,N_1744);
and U2274 (N_2274,N_1634,N_1583);
and U2275 (N_2275,N_1604,N_1359);
nor U2276 (N_2276,N_1713,N_1665);
nand U2277 (N_2277,N_1094,N_1138);
or U2278 (N_2278,N_1142,N_1506);
and U2279 (N_2279,N_1763,N_1900);
nand U2280 (N_2280,N_1568,N_1463);
and U2281 (N_2281,N_1239,N_1989);
or U2282 (N_2282,N_1270,N_1542);
nor U2283 (N_2283,N_1704,N_1749);
or U2284 (N_2284,N_1728,N_1816);
xor U2285 (N_2285,N_1377,N_1790);
nor U2286 (N_2286,N_1007,N_1310);
nand U2287 (N_2287,N_1851,N_1737);
and U2288 (N_2288,N_1721,N_1762);
and U2289 (N_2289,N_1811,N_1978);
nor U2290 (N_2290,N_1433,N_1281);
nor U2291 (N_2291,N_1600,N_1997);
and U2292 (N_2292,N_1072,N_1246);
nand U2293 (N_2293,N_1572,N_1429);
nor U2294 (N_2294,N_1926,N_1894);
nand U2295 (N_2295,N_1158,N_1045);
nand U2296 (N_2296,N_1064,N_1059);
and U2297 (N_2297,N_1476,N_1061);
nand U2298 (N_2298,N_1499,N_1174);
and U2299 (N_2299,N_1380,N_1696);
or U2300 (N_2300,N_1338,N_1280);
nand U2301 (N_2301,N_1101,N_1392);
and U2302 (N_2302,N_1996,N_1206);
nor U2303 (N_2303,N_1053,N_1569);
nand U2304 (N_2304,N_1027,N_1313);
and U2305 (N_2305,N_1271,N_1304);
nand U2306 (N_2306,N_1062,N_1548);
nor U2307 (N_2307,N_1202,N_1008);
or U2308 (N_2308,N_1484,N_1559);
nor U2309 (N_2309,N_1078,N_1589);
nand U2310 (N_2310,N_1409,N_1781);
or U2311 (N_2311,N_1657,N_1089);
xnor U2312 (N_2312,N_1720,N_1040);
nor U2313 (N_2313,N_1624,N_1090);
nor U2314 (N_2314,N_1675,N_1560);
nor U2315 (N_2315,N_1170,N_1567);
nand U2316 (N_2316,N_1876,N_1769);
nand U2317 (N_2317,N_1477,N_1712);
or U2318 (N_2318,N_1638,N_1164);
or U2319 (N_2319,N_1703,N_1317);
or U2320 (N_2320,N_1047,N_1729);
and U2321 (N_2321,N_1646,N_1727);
or U2322 (N_2322,N_1536,N_1801);
or U2323 (N_2323,N_1705,N_1358);
or U2324 (N_2324,N_1421,N_1680);
nand U2325 (N_2325,N_1396,N_1738);
nor U2326 (N_2326,N_1805,N_1862);
or U2327 (N_2327,N_1507,N_1592);
and U2328 (N_2328,N_1794,N_1671);
nand U2329 (N_2329,N_1105,N_1041);
nand U2330 (N_2330,N_1151,N_1784);
or U2331 (N_2331,N_1598,N_1625);
nor U2332 (N_2332,N_1798,N_1644);
or U2333 (N_2333,N_1761,N_1293);
and U2334 (N_2334,N_1466,N_1927);
nand U2335 (N_2335,N_1746,N_1984);
nand U2336 (N_2336,N_1847,N_1627);
nand U2337 (N_2337,N_1435,N_1397);
nor U2338 (N_2338,N_1706,N_1248);
nand U2339 (N_2339,N_1108,N_1024);
and U2340 (N_2340,N_1584,N_1670);
nor U2341 (N_2341,N_1510,N_1685);
nand U2342 (N_2342,N_1865,N_1154);
and U2343 (N_2343,N_1305,N_1898);
or U2344 (N_2344,N_1767,N_1533);
and U2345 (N_2345,N_1087,N_1581);
or U2346 (N_2346,N_1620,N_1877);
and U2347 (N_2347,N_1711,N_1017);
or U2348 (N_2348,N_1571,N_1966);
or U2349 (N_2349,N_1498,N_1083);
nand U2350 (N_2350,N_1962,N_1309);
nand U2351 (N_2351,N_1287,N_1079);
or U2352 (N_2352,N_1211,N_1522);
and U2353 (N_2353,N_1916,N_1055);
nand U2354 (N_2354,N_1585,N_1545);
nand U2355 (N_2355,N_1837,N_1080);
nor U2356 (N_2356,N_1123,N_1688);
nor U2357 (N_2357,N_1618,N_1874);
xor U2358 (N_2358,N_1050,N_1911);
or U2359 (N_2359,N_1342,N_1843);
and U2360 (N_2360,N_1954,N_1175);
nand U2361 (N_2361,N_1949,N_1300);
or U2362 (N_2362,N_1244,N_1425);
nor U2363 (N_2363,N_1792,N_1022);
nor U2364 (N_2364,N_1327,N_1757);
xnor U2365 (N_2365,N_1621,N_1828);
nor U2366 (N_2366,N_1673,N_1362);
nor U2367 (N_2367,N_1698,N_1998);
nand U2368 (N_2368,N_1825,N_1367);
and U2369 (N_2369,N_1787,N_1069);
nor U2370 (N_2370,N_1517,N_1635);
nor U2371 (N_2371,N_1835,N_1269);
nor U2372 (N_2372,N_1056,N_1279);
or U2373 (N_2373,N_1960,N_1144);
nor U2374 (N_2374,N_1010,N_1651);
and U2375 (N_2375,N_1368,N_1756);
nand U2376 (N_2376,N_1134,N_1674);
nand U2377 (N_2377,N_1760,N_1018);
nor U2378 (N_2378,N_1848,N_1163);
and U2379 (N_2379,N_1826,N_1924);
nor U2380 (N_2380,N_1972,N_1974);
and U2381 (N_2381,N_1613,N_1882);
nor U2382 (N_2382,N_1640,N_1136);
nand U2383 (N_2383,N_1683,N_1496);
nand U2384 (N_2384,N_1815,N_1808);
or U2385 (N_2385,N_1393,N_1643);
or U2386 (N_2386,N_1881,N_1958);
nor U2387 (N_2387,N_1547,N_1365);
nand U2388 (N_2388,N_1066,N_1002);
or U2389 (N_2389,N_1599,N_1732);
or U2390 (N_2390,N_1500,N_1068);
nor U2391 (N_2391,N_1261,N_1519);
nor U2392 (N_2392,N_1276,N_1878);
nor U2393 (N_2393,N_1199,N_1512);
and U2394 (N_2394,N_1639,N_1565);
or U2395 (N_2395,N_1431,N_1970);
nand U2396 (N_2396,N_1097,N_1515);
nand U2397 (N_2397,N_1648,N_1986);
or U2398 (N_2398,N_1277,N_1562);
nor U2399 (N_2399,N_1049,N_1531);
nor U2400 (N_2400,N_1479,N_1473);
or U2401 (N_2401,N_1730,N_1689);
nor U2402 (N_2402,N_1867,N_1160);
or U2403 (N_2403,N_1461,N_1532);
and U2404 (N_2404,N_1819,N_1864);
and U2405 (N_2405,N_1501,N_1289);
xor U2406 (N_2406,N_1715,N_1654);
nor U2407 (N_2407,N_1375,N_1120);
nor U2408 (N_2408,N_1406,N_1029);
and U2409 (N_2409,N_1934,N_1726);
or U2410 (N_2410,N_1126,N_1661);
and U2411 (N_2411,N_1803,N_1328);
nor U2412 (N_2412,N_1318,N_1647);
and U2413 (N_2413,N_1283,N_1940);
and U2414 (N_2414,N_1788,N_1725);
or U2415 (N_2415,N_1964,N_1278);
nor U2416 (N_2416,N_1096,N_1886);
nand U2417 (N_2417,N_1667,N_1403);
and U2418 (N_2418,N_1141,N_1678);
nand U2419 (N_2419,N_1578,N_1171);
or U2420 (N_2420,N_1374,N_1005);
or U2421 (N_2421,N_1554,N_1373);
or U2422 (N_2422,N_1307,N_1745);
or U2423 (N_2423,N_1182,N_1521);
and U2424 (N_2424,N_1131,N_1593);
and U2425 (N_2425,N_1766,N_1048);
nor U2426 (N_2426,N_1555,N_1855);
nand U2427 (N_2427,N_1265,N_1347);
and U2428 (N_2428,N_1319,N_1660);
or U2429 (N_2429,N_1607,N_1489);
nor U2430 (N_2430,N_1904,N_1207);
or U2431 (N_2431,N_1457,N_1930);
nand U2432 (N_2432,N_1993,N_1106);
nand U2433 (N_2433,N_1935,N_1118);
or U2434 (N_2434,N_1410,N_1335);
nand U2435 (N_2435,N_1849,N_1852);
nand U2436 (N_2436,N_1504,N_1060);
and U2437 (N_2437,N_1285,N_1888);
and U2438 (N_2438,N_1383,N_1833);
nand U2439 (N_2439,N_1483,N_1478);
nand U2440 (N_2440,N_1001,N_1044);
and U2441 (N_2441,N_1183,N_1810);
nand U2442 (N_2442,N_1576,N_1614);
nor U2443 (N_2443,N_1458,N_1987);
nor U2444 (N_2444,N_1831,N_1941);
nor U2445 (N_2445,N_1405,N_1190);
or U2446 (N_2446,N_1977,N_1299);
or U2447 (N_2447,N_1740,N_1748);
and U2448 (N_2448,N_1039,N_1537);
nand U2449 (N_2449,N_1185,N_1612);
xnor U2450 (N_2450,N_1286,N_1063);
or U2451 (N_2451,N_1645,N_1034);
xnor U2452 (N_2452,N_1416,N_1771);
nand U2453 (N_2453,N_1543,N_1117);
or U2454 (N_2454,N_1075,N_1979);
nor U2455 (N_2455,N_1481,N_1922);
and U2456 (N_2456,N_1445,N_1710);
and U2457 (N_2457,N_1991,N_1341);
and U2458 (N_2458,N_1616,N_1333);
or U2459 (N_2459,N_1937,N_1208);
nor U2460 (N_2460,N_1302,N_1840);
or U2461 (N_2461,N_1995,N_1799);
and U2462 (N_2462,N_1220,N_1226);
and U2463 (N_2463,N_1148,N_1905);
and U2464 (N_2464,N_1356,N_1379);
or U2465 (N_2465,N_1546,N_1400);
nand U2466 (N_2466,N_1971,N_1868);
and U2467 (N_2467,N_1563,N_1702);
nand U2468 (N_2468,N_1428,N_1345);
or U2469 (N_2469,N_1502,N_1462);
or U2470 (N_2470,N_1982,N_1488);
or U2471 (N_2471,N_1165,N_1155);
nand U2472 (N_2472,N_1332,N_1161);
or U2473 (N_2473,N_1879,N_1191);
nor U2474 (N_2474,N_1237,N_1088);
xnor U2475 (N_2475,N_1298,N_1162);
nor U2476 (N_2476,N_1219,N_1697);
or U2477 (N_2477,N_1427,N_1099);
nor U2478 (N_2478,N_1167,N_1032);
nand U2479 (N_2479,N_1939,N_1028);
nand U2480 (N_2480,N_1814,N_1953);
or U2481 (N_2481,N_1188,N_1344);
nand U2482 (N_2482,N_1541,N_1782);
nand U2483 (N_2483,N_1595,N_1493);
nor U2484 (N_2484,N_1153,N_1242);
xor U2485 (N_2485,N_1570,N_1669);
nand U2486 (N_2486,N_1806,N_1388);
or U2487 (N_2487,N_1430,N_1336);
and U2488 (N_2488,N_1221,N_1404);
or U2489 (N_2489,N_1014,N_1551);
or U2490 (N_2490,N_1020,N_1129);
nand U2491 (N_2491,N_1455,N_1758);
nor U2492 (N_2492,N_1540,N_1656);
and U2493 (N_2493,N_1793,N_1354);
and U2494 (N_2494,N_1186,N_1891);
nand U2495 (N_2495,N_1213,N_1538);
or U2496 (N_2496,N_1076,N_1628);
or U2497 (N_2497,N_1189,N_1933);
nand U2498 (N_2498,N_1370,N_1084);
or U2499 (N_2499,N_1395,N_1452);
and U2500 (N_2500,N_1217,N_1306);
and U2501 (N_2501,N_1127,N_1391);
and U2502 (N_2502,N_1192,N_1096);
or U2503 (N_2503,N_1952,N_1376);
nand U2504 (N_2504,N_1564,N_1060);
and U2505 (N_2505,N_1275,N_1649);
nor U2506 (N_2506,N_1507,N_1273);
nor U2507 (N_2507,N_1487,N_1950);
nor U2508 (N_2508,N_1617,N_1869);
or U2509 (N_2509,N_1263,N_1650);
nand U2510 (N_2510,N_1828,N_1006);
and U2511 (N_2511,N_1159,N_1742);
or U2512 (N_2512,N_1327,N_1122);
nand U2513 (N_2513,N_1847,N_1804);
nand U2514 (N_2514,N_1291,N_1776);
and U2515 (N_2515,N_1041,N_1540);
nor U2516 (N_2516,N_1122,N_1441);
and U2517 (N_2517,N_1380,N_1564);
nand U2518 (N_2518,N_1193,N_1471);
nand U2519 (N_2519,N_1131,N_1767);
and U2520 (N_2520,N_1186,N_1659);
and U2521 (N_2521,N_1205,N_1270);
or U2522 (N_2522,N_1228,N_1650);
or U2523 (N_2523,N_1945,N_1069);
or U2524 (N_2524,N_1384,N_1922);
and U2525 (N_2525,N_1814,N_1896);
or U2526 (N_2526,N_1788,N_1770);
or U2527 (N_2527,N_1642,N_1994);
or U2528 (N_2528,N_1678,N_1536);
and U2529 (N_2529,N_1171,N_1617);
nand U2530 (N_2530,N_1786,N_1845);
and U2531 (N_2531,N_1145,N_1263);
nand U2532 (N_2532,N_1171,N_1841);
xor U2533 (N_2533,N_1399,N_1705);
nand U2534 (N_2534,N_1466,N_1340);
and U2535 (N_2535,N_1812,N_1825);
nand U2536 (N_2536,N_1610,N_1802);
nor U2537 (N_2537,N_1245,N_1472);
or U2538 (N_2538,N_1774,N_1773);
nand U2539 (N_2539,N_1204,N_1432);
and U2540 (N_2540,N_1058,N_1325);
or U2541 (N_2541,N_1973,N_1236);
and U2542 (N_2542,N_1154,N_1341);
or U2543 (N_2543,N_1634,N_1094);
or U2544 (N_2544,N_1853,N_1696);
and U2545 (N_2545,N_1579,N_1337);
nor U2546 (N_2546,N_1592,N_1527);
and U2547 (N_2547,N_1077,N_1095);
nor U2548 (N_2548,N_1145,N_1862);
or U2549 (N_2549,N_1046,N_1110);
or U2550 (N_2550,N_1119,N_1557);
or U2551 (N_2551,N_1297,N_1206);
and U2552 (N_2552,N_1302,N_1353);
nand U2553 (N_2553,N_1891,N_1876);
and U2554 (N_2554,N_1532,N_1913);
nor U2555 (N_2555,N_1556,N_1938);
nand U2556 (N_2556,N_1889,N_1675);
and U2557 (N_2557,N_1779,N_1963);
and U2558 (N_2558,N_1513,N_1130);
and U2559 (N_2559,N_1593,N_1018);
and U2560 (N_2560,N_1585,N_1022);
nor U2561 (N_2561,N_1651,N_1283);
or U2562 (N_2562,N_1920,N_1336);
or U2563 (N_2563,N_1949,N_1652);
nor U2564 (N_2564,N_1105,N_1606);
and U2565 (N_2565,N_1498,N_1810);
and U2566 (N_2566,N_1630,N_1013);
nand U2567 (N_2567,N_1284,N_1251);
xor U2568 (N_2568,N_1904,N_1321);
nor U2569 (N_2569,N_1811,N_1835);
nand U2570 (N_2570,N_1181,N_1364);
and U2571 (N_2571,N_1245,N_1075);
nor U2572 (N_2572,N_1980,N_1301);
and U2573 (N_2573,N_1241,N_1334);
or U2574 (N_2574,N_1799,N_1235);
and U2575 (N_2575,N_1093,N_1064);
nand U2576 (N_2576,N_1267,N_1473);
or U2577 (N_2577,N_1258,N_1432);
or U2578 (N_2578,N_1345,N_1812);
nand U2579 (N_2579,N_1303,N_1853);
or U2580 (N_2580,N_1279,N_1059);
or U2581 (N_2581,N_1327,N_1940);
or U2582 (N_2582,N_1170,N_1730);
and U2583 (N_2583,N_1873,N_1106);
nand U2584 (N_2584,N_1831,N_1226);
nand U2585 (N_2585,N_1942,N_1252);
and U2586 (N_2586,N_1052,N_1873);
nand U2587 (N_2587,N_1549,N_1000);
nor U2588 (N_2588,N_1265,N_1877);
nor U2589 (N_2589,N_1749,N_1151);
and U2590 (N_2590,N_1366,N_1599);
nor U2591 (N_2591,N_1775,N_1152);
nor U2592 (N_2592,N_1578,N_1562);
and U2593 (N_2593,N_1208,N_1465);
nand U2594 (N_2594,N_1276,N_1950);
nor U2595 (N_2595,N_1119,N_1226);
nand U2596 (N_2596,N_1170,N_1150);
and U2597 (N_2597,N_1016,N_1187);
or U2598 (N_2598,N_1268,N_1942);
nand U2599 (N_2599,N_1595,N_1839);
or U2600 (N_2600,N_1366,N_1037);
nand U2601 (N_2601,N_1301,N_1548);
and U2602 (N_2602,N_1537,N_1331);
nor U2603 (N_2603,N_1062,N_1166);
nor U2604 (N_2604,N_1766,N_1544);
and U2605 (N_2605,N_1614,N_1476);
nor U2606 (N_2606,N_1686,N_1803);
and U2607 (N_2607,N_1140,N_1153);
nor U2608 (N_2608,N_1114,N_1852);
nor U2609 (N_2609,N_1262,N_1751);
or U2610 (N_2610,N_1871,N_1591);
or U2611 (N_2611,N_1844,N_1967);
nand U2612 (N_2612,N_1259,N_1197);
nor U2613 (N_2613,N_1640,N_1798);
or U2614 (N_2614,N_1353,N_1366);
nor U2615 (N_2615,N_1853,N_1951);
nand U2616 (N_2616,N_1737,N_1705);
and U2617 (N_2617,N_1058,N_1857);
xor U2618 (N_2618,N_1919,N_1688);
nor U2619 (N_2619,N_1198,N_1761);
nand U2620 (N_2620,N_1501,N_1158);
nor U2621 (N_2621,N_1603,N_1986);
nand U2622 (N_2622,N_1667,N_1878);
nor U2623 (N_2623,N_1613,N_1955);
and U2624 (N_2624,N_1139,N_1341);
or U2625 (N_2625,N_1876,N_1041);
or U2626 (N_2626,N_1192,N_1807);
or U2627 (N_2627,N_1466,N_1116);
and U2628 (N_2628,N_1684,N_1101);
and U2629 (N_2629,N_1808,N_1901);
nor U2630 (N_2630,N_1595,N_1781);
nand U2631 (N_2631,N_1898,N_1531);
nand U2632 (N_2632,N_1041,N_1811);
and U2633 (N_2633,N_1672,N_1825);
nor U2634 (N_2634,N_1980,N_1265);
or U2635 (N_2635,N_1573,N_1963);
nand U2636 (N_2636,N_1618,N_1036);
nor U2637 (N_2637,N_1315,N_1492);
or U2638 (N_2638,N_1999,N_1188);
nor U2639 (N_2639,N_1029,N_1919);
nor U2640 (N_2640,N_1380,N_1751);
nand U2641 (N_2641,N_1006,N_1822);
nor U2642 (N_2642,N_1362,N_1758);
and U2643 (N_2643,N_1925,N_1788);
nand U2644 (N_2644,N_1677,N_1076);
and U2645 (N_2645,N_1097,N_1434);
nor U2646 (N_2646,N_1993,N_1464);
or U2647 (N_2647,N_1992,N_1890);
nand U2648 (N_2648,N_1088,N_1764);
or U2649 (N_2649,N_1971,N_1876);
nor U2650 (N_2650,N_1653,N_1346);
nand U2651 (N_2651,N_1663,N_1656);
or U2652 (N_2652,N_1232,N_1423);
and U2653 (N_2653,N_1290,N_1451);
nor U2654 (N_2654,N_1163,N_1827);
xnor U2655 (N_2655,N_1814,N_1755);
and U2656 (N_2656,N_1614,N_1028);
nor U2657 (N_2657,N_1450,N_1884);
and U2658 (N_2658,N_1375,N_1774);
nor U2659 (N_2659,N_1296,N_1485);
nand U2660 (N_2660,N_1027,N_1102);
nor U2661 (N_2661,N_1428,N_1131);
nor U2662 (N_2662,N_1630,N_1996);
and U2663 (N_2663,N_1832,N_1016);
nor U2664 (N_2664,N_1128,N_1899);
and U2665 (N_2665,N_1787,N_1840);
or U2666 (N_2666,N_1350,N_1263);
nor U2667 (N_2667,N_1872,N_1244);
or U2668 (N_2668,N_1869,N_1088);
and U2669 (N_2669,N_1292,N_1097);
and U2670 (N_2670,N_1887,N_1365);
nor U2671 (N_2671,N_1420,N_1694);
or U2672 (N_2672,N_1220,N_1333);
nand U2673 (N_2673,N_1482,N_1988);
and U2674 (N_2674,N_1517,N_1945);
nand U2675 (N_2675,N_1481,N_1760);
nor U2676 (N_2676,N_1462,N_1752);
and U2677 (N_2677,N_1832,N_1299);
and U2678 (N_2678,N_1183,N_1900);
or U2679 (N_2679,N_1541,N_1990);
or U2680 (N_2680,N_1113,N_1995);
and U2681 (N_2681,N_1308,N_1875);
nor U2682 (N_2682,N_1920,N_1033);
nor U2683 (N_2683,N_1322,N_1481);
and U2684 (N_2684,N_1874,N_1420);
or U2685 (N_2685,N_1716,N_1418);
or U2686 (N_2686,N_1955,N_1173);
or U2687 (N_2687,N_1285,N_1154);
nor U2688 (N_2688,N_1289,N_1767);
nand U2689 (N_2689,N_1218,N_1182);
nand U2690 (N_2690,N_1370,N_1745);
or U2691 (N_2691,N_1689,N_1110);
nor U2692 (N_2692,N_1219,N_1886);
or U2693 (N_2693,N_1601,N_1811);
and U2694 (N_2694,N_1812,N_1847);
and U2695 (N_2695,N_1085,N_1957);
nor U2696 (N_2696,N_1930,N_1734);
or U2697 (N_2697,N_1993,N_1666);
nand U2698 (N_2698,N_1941,N_1290);
and U2699 (N_2699,N_1559,N_1754);
nor U2700 (N_2700,N_1607,N_1169);
or U2701 (N_2701,N_1453,N_1341);
or U2702 (N_2702,N_1483,N_1822);
nor U2703 (N_2703,N_1738,N_1536);
nand U2704 (N_2704,N_1642,N_1444);
nor U2705 (N_2705,N_1587,N_1959);
or U2706 (N_2706,N_1376,N_1747);
or U2707 (N_2707,N_1034,N_1073);
and U2708 (N_2708,N_1897,N_1258);
and U2709 (N_2709,N_1892,N_1743);
or U2710 (N_2710,N_1240,N_1080);
nor U2711 (N_2711,N_1863,N_1610);
nor U2712 (N_2712,N_1447,N_1290);
and U2713 (N_2713,N_1471,N_1272);
nand U2714 (N_2714,N_1752,N_1843);
and U2715 (N_2715,N_1500,N_1901);
nand U2716 (N_2716,N_1708,N_1966);
or U2717 (N_2717,N_1120,N_1546);
or U2718 (N_2718,N_1087,N_1458);
and U2719 (N_2719,N_1501,N_1764);
xor U2720 (N_2720,N_1757,N_1145);
nand U2721 (N_2721,N_1495,N_1564);
nor U2722 (N_2722,N_1127,N_1199);
and U2723 (N_2723,N_1357,N_1979);
nand U2724 (N_2724,N_1052,N_1086);
and U2725 (N_2725,N_1291,N_1292);
nor U2726 (N_2726,N_1749,N_1819);
nor U2727 (N_2727,N_1482,N_1323);
nand U2728 (N_2728,N_1341,N_1240);
nand U2729 (N_2729,N_1659,N_1109);
nand U2730 (N_2730,N_1934,N_1506);
nor U2731 (N_2731,N_1819,N_1015);
or U2732 (N_2732,N_1576,N_1536);
or U2733 (N_2733,N_1981,N_1139);
nor U2734 (N_2734,N_1733,N_1956);
or U2735 (N_2735,N_1866,N_1686);
or U2736 (N_2736,N_1938,N_1815);
or U2737 (N_2737,N_1607,N_1472);
and U2738 (N_2738,N_1025,N_1170);
or U2739 (N_2739,N_1875,N_1894);
nor U2740 (N_2740,N_1345,N_1179);
nor U2741 (N_2741,N_1295,N_1141);
nor U2742 (N_2742,N_1343,N_1691);
nand U2743 (N_2743,N_1939,N_1283);
and U2744 (N_2744,N_1359,N_1743);
or U2745 (N_2745,N_1740,N_1710);
nand U2746 (N_2746,N_1456,N_1498);
and U2747 (N_2747,N_1283,N_1716);
nor U2748 (N_2748,N_1704,N_1662);
or U2749 (N_2749,N_1071,N_1047);
and U2750 (N_2750,N_1987,N_1151);
nand U2751 (N_2751,N_1844,N_1546);
nand U2752 (N_2752,N_1248,N_1249);
nand U2753 (N_2753,N_1788,N_1560);
and U2754 (N_2754,N_1017,N_1044);
or U2755 (N_2755,N_1449,N_1095);
or U2756 (N_2756,N_1548,N_1895);
nor U2757 (N_2757,N_1510,N_1372);
or U2758 (N_2758,N_1005,N_1228);
or U2759 (N_2759,N_1190,N_1133);
nand U2760 (N_2760,N_1697,N_1621);
nand U2761 (N_2761,N_1982,N_1886);
xor U2762 (N_2762,N_1755,N_1361);
nor U2763 (N_2763,N_1349,N_1839);
nor U2764 (N_2764,N_1270,N_1922);
or U2765 (N_2765,N_1022,N_1880);
and U2766 (N_2766,N_1906,N_1829);
xor U2767 (N_2767,N_1143,N_1022);
and U2768 (N_2768,N_1631,N_1166);
nand U2769 (N_2769,N_1640,N_1760);
nor U2770 (N_2770,N_1554,N_1046);
or U2771 (N_2771,N_1696,N_1388);
nand U2772 (N_2772,N_1998,N_1007);
and U2773 (N_2773,N_1310,N_1358);
nand U2774 (N_2774,N_1615,N_1529);
or U2775 (N_2775,N_1185,N_1331);
and U2776 (N_2776,N_1003,N_1992);
nand U2777 (N_2777,N_1907,N_1489);
or U2778 (N_2778,N_1801,N_1832);
nand U2779 (N_2779,N_1865,N_1860);
or U2780 (N_2780,N_1452,N_1524);
or U2781 (N_2781,N_1952,N_1522);
nor U2782 (N_2782,N_1655,N_1514);
nor U2783 (N_2783,N_1353,N_1030);
xor U2784 (N_2784,N_1794,N_1038);
nand U2785 (N_2785,N_1811,N_1379);
nor U2786 (N_2786,N_1998,N_1202);
nand U2787 (N_2787,N_1640,N_1083);
nor U2788 (N_2788,N_1141,N_1190);
nand U2789 (N_2789,N_1240,N_1010);
and U2790 (N_2790,N_1742,N_1062);
nand U2791 (N_2791,N_1672,N_1293);
nor U2792 (N_2792,N_1345,N_1143);
xor U2793 (N_2793,N_1719,N_1156);
and U2794 (N_2794,N_1762,N_1014);
nand U2795 (N_2795,N_1193,N_1289);
or U2796 (N_2796,N_1470,N_1821);
and U2797 (N_2797,N_1444,N_1374);
nor U2798 (N_2798,N_1296,N_1405);
nor U2799 (N_2799,N_1498,N_1578);
nand U2800 (N_2800,N_1812,N_1134);
nor U2801 (N_2801,N_1875,N_1734);
and U2802 (N_2802,N_1110,N_1748);
nor U2803 (N_2803,N_1126,N_1870);
or U2804 (N_2804,N_1990,N_1672);
nand U2805 (N_2805,N_1437,N_1197);
nor U2806 (N_2806,N_1207,N_1190);
and U2807 (N_2807,N_1359,N_1419);
and U2808 (N_2808,N_1014,N_1593);
nand U2809 (N_2809,N_1106,N_1483);
nand U2810 (N_2810,N_1449,N_1667);
or U2811 (N_2811,N_1537,N_1005);
nor U2812 (N_2812,N_1695,N_1875);
nand U2813 (N_2813,N_1966,N_1740);
and U2814 (N_2814,N_1581,N_1721);
nand U2815 (N_2815,N_1039,N_1629);
nor U2816 (N_2816,N_1266,N_1359);
nand U2817 (N_2817,N_1485,N_1894);
nor U2818 (N_2818,N_1121,N_1664);
and U2819 (N_2819,N_1405,N_1865);
nand U2820 (N_2820,N_1004,N_1581);
or U2821 (N_2821,N_1156,N_1194);
and U2822 (N_2822,N_1065,N_1190);
and U2823 (N_2823,N_1309,N_1508);
and U2824 (N_2824,N_1913,N_1844);
and U2825 (N_2825,N_1932,N_1871);
nand U2826 (N_2826,N_1421,N_1646);
nor U2827 (N_2827,N_1810,N_1026);
and U2828 (N_2828,N_1713,N_1624);
xor U2829 (N_2829,N_1599,N_1995);
nor U2830 (N_2830,N_1796,N_1030);
nand U2831 (N_2831,N_1252,N_1261);
nand U2832 (N_2832,N_1015,N_1681);
or U2833 (N_2833,N_1592,N_1030);
or U2834 (N_2834,N_1557,N_1086);
and U2835 (N_2835,N_1753,N_1027);
nand U2836 (N_2836,N_1889,N_1643);
nor U2837 (N_2837,N_1848,N_1291);
and U2838 (N_2838,N_1216,N_1655);
nor U2839 (N_2839,N_1391,N_1582);
and U2840 (N_2840,N_1093,N_1102);
or U2841 (N_2841,N_1281,N_1104);
or U2842 (N_2842,N_1010,N_1494);
and U2843 (N_2843,N_1390,N_1071);
and U2844 (N_2844,N_1436,N_1297);
or U2845 (N_2845,N_1664,N_1262);
or U2846 (N_2846,N_1432,N_1953);
and U2847 (N_2847,N_1722,N_1325);
nor U2848 (N_2848,N_1900,N_1904);
and U2849 (N_2849,N_1846,N_1477);
nand U2850 (N_2850,N_1479,N_1195);
nor U2851 (N_2851,N_1172,N_1143);
and U2852 (N_2852,N_1991,N_1472);
nor U2853 (N_2853,N_1795,N_1300);
nand U2854 (N_2854,N_1653,N_1401);
nand U2855 (N_2855,N_1487,N_1758);
or U2856 (N_2856,N_1313,N_1963);
nor U2857 (N_2857,N_1254,N_1982);
or U2858 (N_2858,N_1614,N_1480);
or U2859 (N_2859,N_1643,N_1005);
and U2860 (N_2860,N_1238,N_1080);
or U2861 (N_2861,N_1755,N_1752);
and U2862 (N_2862,N_1594,N_1957);
nor U2863 (N_2863,N_1077,N_1348);
nand U2864 (N_2864,N_1963,N_1775);
or U2865 (N_2865,N_1472,N_1671);
or U2866 (N_2866,N_1897,N_1307);
nand U2867 (N_2867,N_1653,N_1152);
nor U2868 (N_2868,N_1313,N_1950);
or U2869 (N_2869,N_1527,N_1720);
nor U2870 (N_2870,N_1909,N_1648);
nand U2871 (N_2871,N_1997,N_1479);
and U2872 (N_2872,N_1257,N_1213);
or U2873 (N_2873,N_1969,N_1096);
or U2874 (N_2874,N_1006,N_1940);
and U2875 (N_2875,N_1719,N_1292);
nand U2876 (N_2876,N_1813,N_1109);
or U2877 (N_2877,N_1745,N_1082);
and U2878 (N_2878,N_1746,N_1554);
or U2879 (N_2879,N_1098,N_1429);
or U2880 (N_2880,N_1002,N_1987);
nor U2881 (N_2881,N_1176,N_1748);
and U2882 (N_2882,N_1382,N_1930);
nand U2883 (N_2883,N_1023,N_1239);
and U2884 (N_2884,N_1925,N_1108);
nor U2885 (N_2885,N_1999,N_1118);
and U2886 (N_2886,N_1303,N_1113);
and U2887 (N_2887,N_1670,N_1300);
or U2888 (N_2888,N_1236,N_1239);
and U2889 (N_2889,N_1893,N_1089);
or U2890 (N_2890,N_1535,N_1385);
nand U2891 (N_2891,N_1599,N_1780);
nor U2892 (N_2892,N_1478,N_1744);
or U2893 (N_2893,N_1775,N_1981);
nor U2894 (N_2894,N_1088,N_1405);
or U2895 (N_2895,N_1149,N_1228);
and U2896 (N_2896,N_1792,N_1794);
or U2897 (N_2897,N_1841,N_1706);
nand U2898 (N_2898,N_1021,N_1842);
and U2899 (N_2899,N_1973,N_1728);
and U2900 (N_2900,N_1013,N_1231);
or U2901 (N_2901,N_1863,N_1538);
or U2902 (N_2902,N_1532,N_1169);
or U2903 (N_2903,N_1802,N_1064);
nand U2904 (N_2904,N_1463,N_1208);
and U2905 (N_2905,N_1387,N_1936);
nor U2906 (N_2906,N_1149,N_1313);
or U2907 (N_2907,N_1831,N_1665);
and U2908 (N_2908,N_1647,N_1953);
nand U2909 (N_2909,N_1342,N_1698);
nand U2910 (N_2910,N_1606,N_1720);
or U2911 (N_2911,N_1891,N_1089);
and U2912 (N_2912,N_1332,N_1423);
nand U2913 (N_2913,N_1077,N_1967);
nor U2914 (N_2914,N_1165,N_1780);
or U2915 (N_2915,N_1293,N_1952);
nor U2916 (N_2916,N_1925,N_1216);
nand U2917 (N_2917,N_1267,N_1304);
nand U2918 (N_2918,N_1131,N_1727);
nand U2919 (N_2919,N_1666,N_1462);
and U2920 (N_2920,N_1970,N_1433);
xnor U2921 (N_2921,N_1919,N_1921);
nand U2922 (N_2922,N_1862,N_1149);
and U2923 (N_2923,N_1022,N_1821);
or U2924 (N_2924,N_1985,N_1016);
nand U2925 (N_2925,N_1773,N_1541);
and U2926 (N_2926,N_1400,N_1907);
nand U2927 (N_2927,N_1461,N_1733);
nand U2928 (N_2928,N_1688,N_1764);
nor U2929 (N_2929,N_1121,N_1477);
nand U2930 (N_2930,N_1703,N_1175);
nor U2931 (N_2931,N_1119,N_1971);
or U2932 (N_2932,N_1621,N_1819);
nor U2933 (N_2933,N_1999,N_1801);
or U2934 (N_2934,N_1372,N_1906);
nor U2935 (N_2935,N_1626,N_1080);
and U2936 (N_2936,N_1953,N_1750);
nand U2937 (N_2937,N_1241,N_1479);
nor U2938 (N_2938,N_1352,N_1022);
nand U2939 (N_2939,N_1997,N_1427);
and U2940 (N_2940,N_1683,N_1591);
nand U2941 (N_2941,N_1850,N_1584);
and U2942 (N_2942,N_1371,N_1002);
and U2943 (N_2943,N_1673,N_1196);
nor U2944 (N_2944,N_1195,N_1472);
and U2945 (N_2945,N_1777,N_1123);
nand U2946 (N_2946,N_1680,N_1667);
and U2947 (N_2947,N_1014,N_1949);
or U2948 (N_2948,N_1131,N_1881);
nand U2949 (N_2949,N_1254,N_1997);
nand U2950 (N_2950,N_1468,N_1899);
nand U2951 (N_2951,N_1208,N_1874);
nor U2952 (N_2952,N_1741,N_1044);
and U2953 (N_2953,N_1027,N_1211);
or U2954 (N_2954,N_1774,N_1393);
or U2955 (N_2955,N_1855,N_1024);
nor U2956 (N_2956,N_1006,N_1696);
nor U2957 (N_2957,N_1152,N_1200);
nand U2958 (N_2958,N_1090,N_1474);
and U2959 (N_2959,N_1324,N_1864);
nand U2960 (N_2960,N_1469,N_1855);
nor U2961 (N_2961,N_1791,N_1674);
and U2962 (N_2962,N_1236,N_1421);
xor U2963 (N_2963,N_1072,N_1738);
nor U2964 (N_2964,N_1204,N_1514);
nand U2965 (N_2965,N_1102,N_1227);
nand U2966 (N_2966,N_1936,N_1135);
nand U2967 (N_2967,N_1204,N_1617);
nand U2968 (N_2968,N_1035,N_1897);
or U2969 (N_2969,N_1154,N_1774);
or U2970 (N_2970,N_1014,N_1298);
or U2971 (N_2971,N_1493,N_1318);
and U2972 (N_2972,N_1853,N_1114);
nand U2973 (N_2973,N_1655,N_1066);
nand U2974 (N_2974,N_1175,N_1765);
nand U2975 (N_2975,N_1906,N_1230);
or U2976 (N_2976,N_1045,N_1342);
xor U2977 (N_2977,N_1347,N_1848);
or U2978 (N_2978,N_1846,N_1098);
nor U2979 (N_2979,N_1314,N_1034);
or U2980 (N_2980,N_1814,N_1830);
xor U2981 (N_2981,N_1471,N_1885);
nor U2982 (N_2982,N_1644,N_1008);
nand U2983 (N_2983,N_1161,N_1687);
nand U2984 (N_2984,N_1785,N_1538);
nand U2985 (N_2985,N_1239,N_1227);
nand U2986 (N_2986,N_1784,N_1888);
nand U2987 (N_2987,N_1714,N_1740);
nand U2988 (N_2988,N_1874,N_1829);
nor U2989 (N_2989,N_1849,N_1294);
or U2990 (N_2990,N_1170,N_1068);
and U2991 (N_2991,N_1032,N_1268);
nor U2992 (N_2992,N_1916,N_1920);
nor U2993 (N_2993,N_1611,N_1912);
nor U2994 (N_2994,N_1848,N_1336);
nor U2995 (N_2995,N_1179,N_1037);
xnor U2996 (N_2996,N_1602,N_1719);
nand U2997 (N_2997,N_1009,N_1560);
or U2998 (N_2998,N_1939,N_1941);
and U2999 (N_2999,N_1237,N_1014);
and U3000 (N_3000,N_2165,N_2247);
nor U3001 (N_3001,N_2492,N_2632);
xnor U3002 (N_3002,N_2903,N_2219);
nand U3003 (N_3003,N_2383,N_2693);
nor U3004 (N_3004,N_2627,N_2960);
nor U3005 (N_3005,N_2944,N_2140);
nor U3006 (N_3006,N_2063,N_2856);
nand U3007 (N_3007,N_2688,N_2530);
and U3008 (N_3008,N_2723,N_2348);
nand U3009 (N_3009,N_2604,N_2649);
nand U3010 (N_3010,N_2470,N_2394);
nor U3011 (N_3011,N_2204,N_2437);
nand U3012 (N_3012,N_2767,N_2934);
and U3013 (N_3013,N_2188,N_2322);
or U3014 (N_3014,N_2133,N_2123);
or U3015 (N_3015,N_2257,N_2864);
nor U3016 (N_3016,N_2429,N_2045);
nand U3017 (N_3017,N_2240,N_2846);
nor U3018 (N_3018,N_2464,N_2167);
nand U3019 (N_3019,N_2695,N_2738);
or U3020 (N_3020,N_2332,N_2431);
or U3021 (N_3021,N_2516,N_2806);
and U3022 (N_3022,N_2807,N_2430);
or U3023 (N_3023,N_2832,N_2007);
nand U3024 (N_3024,N_2355,N_2619);
and U3025 (N_3025,N_2075,N_2935);
nand U3026 (N_3026,N_2639,N_2117);
nand U3027 (N_3027,N_2377,N_2000);
xor U3028 (N_3028,N_2620,N_2655);
and U3029 (N_3029,N_2783,N_2917);
nor U3030 (N_3030,N_2091,N_2034);
and U3031 (N_3031,N_2652,N_2481);
nand U3032 (N_3032,N_2787,N_2413);
or U3033 (N_3033,N_2284,N_2775);
nand U3034 (N_3034,N_2364,N_2495);
and U3035 (N_3035,N_2291,N_2535);
and U3036 (N_3036,N_2074,N_2904);
or U3037 (N_3037,N_2670,N_2035);
nor U3038 (N_3038,N_2385,N_2040);
or U3039 (N_3039,N_2174,N_2854);
nand U3040 (N_3040,N_2131,N_2511);
nor U3041 (N_3041,N_2786,N_2814);
nand U3042 (N_3042,N_2937,N_2745);
or U3043 (N_3043,N_2606,N_2314);
and U3044 (N_3044,N_2714,N_2451);
nor U3045 (N_3045,N_2093,N_2972);
nor U3046 (N_3046,N_2386,N_2958);
nand U3047 (N_3047,N_2363,N_2641);
nand U3048 (N_3048,N_2466,N_2698);
nand U3049 (N_3049,N_2733,N_2054);
and U3050 (N_3050,N_2577,N_2270);
or U3051 (N_3051,N_2721,N_2319);
xnor U3052 (N_3052,N_2390,N_2462);
nor U3053 (N_3053,N_2845,N_2456);
nor U3054 (N_3054,N_2664,N_2764);
or U3055 (N_3055,N_2229,N_2849);
or U3056 (N_3056,N_2209,N_2740);
nand U3057 (N_3057,N_2378,N_2870);
and U3058 (N_3058,N_2736,N_2907);
nand U3059 (N_3059,N_2153,N_2246);
nand U3060 (N_3060,N_2758,N_2657);
nand U3061 (N_3061,N_2112,N_2942);
xor U3062 (N_3062,N_2605,N_2732);
nor U3063 (N_3063,N_2899,N_2964);
and U3064 (N_3064,N_2803,N_2371);
or U3065 (N_3065,N_2275,N_2752);
or U3066 (N_3066,N_2144,N_2759);
nand U3067 (N_3067,N_2196,N_2599);
and U3068 (N_3068,N_2947,N_2438);
nor U3069 (N_3069,N_2457,N_2003);
or U3070 (N_3070,N_2690,N_2529);
xnor U3071 (N_3071,N_2648,N_2876);
and U3072 (N_3072,N_2614,N_2242);
nand U3073 (N_3073,N_2677,N_2800);
nor U3074 (N_3074,N_2062,N_2598);
nor U3075 (N_3075,N_2997,N_2135);
or U3076 (N_3076,N_2175,N_2354);
and U3077 (N_3077,N_2099,N_2720);
or U3078 (N_3078,N_2742,N_2852);
and U3079 (N_3079,N_2628,N_2223);
and U3080 (N_3080,N_2224,N_2624);
and U3081 (N_3081,N_2556,N_2453);
nor U3082 (N_3082,N_2588,N_2872);
nand U3083 (N_3083,N_2396,N_2743);
or U3084 (N_3084,N_2662,N_2032);
and U3085 (N_3085,N_2881,N_2748);
nor U3086 (N_3086,N_2531,N_2358);
or U3087 (N_3087,N_2602,N_2946);
or U3088 (N_3088,N_2412,N_2191);
nor U3089 (N_3089,N_2900,N_2809);
and U3090 (N_3090,N_2537,N_2791);
nand U3091 (N_3091,N_2879,N_2067);
or U3092 (N_3092,N_2129,N_2966);
or U3093 (N_3093,N_2269,N_2924);
or U3094 (N_3094,N_2799,N_2086);
or U3095 (N_3095,N_2974,N_2716);
or U3096 (N_3096,N_2256,N_2763);
or U3097 (N_3097,N_2667,N_2392);
nand U3098 (N_3098,N_2236,N_2482);
and U3099 (N_3099,N_2812,N_2681);
nor U3100 (N_3100,N_2212,N_2336);
and U3101 (N_3101,N_2414,N_2169);
nand U3102 (N_3102,N_2725,N_2595);
nor U3103 (N_3103,N_2692,N_2747);
nor U3104 (N_3104,N_2558,N_2058);
and U3105 (N_3105,N_2724,N_2940);
nor U3106 (N_3106,N_2887,N_2391);
nand U3107 (N_3107,N_2017,N_2452);
nor U3108 (N_3108,N_2288,N_2327);
or U3109 (N_3109,N_2335,N_2202);
nand U3110 (N_3110,N_2611,N_2633);
or U3111 (N_3111,N_2376,N_2933);
nand U3112 (N_3112,N_2160,N_2147);
nor U3113 (N_3113,N_2976,N_2741);
and U3114 (N_3114,N_2761,N_2936);
nand U3115 (N_3115,N_2410,N_2709);
nor U3116 (N_3116,N_2717,N_2168);
nor U3117 (N_3117,N_2315,N_2861);
or U3118 (N_3118,N_2318,N_2258);
nor U3119 (N_3119,N_2132,N_2389);
or U3120 (N_3120,N_2102,N_2361);
and U3121 (N_3121,N_2417,N_2467);
nor U3122 (N_3122,N_2221,N_2778);
and U3123 (N_3123,N_2066,N_2243);
nor U3124 (N_3124,N_2722,N_2918);
nand U3125 (N_3125,N_2834,N_2894);
or U3126 (N_3126,N_2506,N_2345);
nand U3127 (N_3127,N_2488,N_2827);
nand U3128 (N_3128,N_2965,N_2434);
or U3129 (N_3129,N_2828,N_2163);
nor U3130 (N_3130,N_2645,N_2995);
nor U3131 (N_3131,N_2494,N_2638);
nor U3132 (N_3132,N_2986,N_2514);
xor U3133 (N_3133,N_2475,N_2796);
or U3134 (N_3134,N_2047,N_2938);
nor U3135 (N_3135,N_2612,N_2850);
nor U3136 (N_3136,N_2433,N_2955);
and U3137 (N_3137,N_2730,N_2181);
or U3138 (N_3138,N_2238,N_2959);
nor U3139 (N_3139,N_2836,N_2517);
nor U3140 (N_3140,N_2374,N_2746);
and U3141 (N_3141,N_2211,N_2519);
or U3142 (N_3142,N_2979,N_2218);
nor U3143 (N_3143,N_2427,N_2963);
nand U3144 (N_3144,N_2571,N_2561);
nor U3145 (N_3145,N_2473,N_2715);
xor U3146 (N_3146,N_2267,N_2950);
and U3147 (N_3147,N_2815,N_2625);
nand U3148 (N_3148,N_2014,N_2838);
nand U3149 (N_3149,N_2330,N_2290);
and U3150 (N_3150,N_2309,N_2908);
nand U3151 (N_3151,N_2436,N_2265);
and U3152 (N_3152,N_2992,N_2151);
or U3153 (N_3153,N_2274,N_2948);
nand U3154 (N_3154,N_2909,N_2448);
or U3155 (N_3155,N_2308,N_2210);
and U3156 (N_3156,N_2549,N_2072);
and U3157 (N_3157,N_2603,N_2435);
and U3158 (N_3158,N_2989,N_2663);
or U3159 (N_3159,N_2483,N_2888);
nor U3160 (N_3160,N_2671,N_2932);
xor U3161 (N_3161,N_2418,N_2220);
and U3162 (N_3162,N_2016,N_2981);
and U3163 (N_3163,N_2416,N_2178);
nor U3164 (N_3164,N_2176,N_2923);
nand U3165 (N_3165,N_2768,N_2341);
nor U3166 (N_3166,N_2021,N_2970);
and U3167 (N_3167,N_2712,N_2420);
or U3168 (N_3168,N_2039,N_2277);
nand U3169 (N_3169,N_2630,N_2069);
or U3170 (N_3170,N_2851,N_2208);
or U3171 (N_3171,N_2460,N_2941);
and U3172 (N_3172,N_2772,N_2447);
or U3173 (N_3173,N_2527,N_2037);
or U3174 (N_3174,N_2076,N_2104);
nor U3175 (N_3175,N_2490,N_2750);
and U3176 (N_3176,N_2644,N_2161);
or U3177 (N_3177,N_2073,N_2019);
and U3178 (N_3178,N_2651,N_2214);
or U3179 (N_3179,N_2773,N_2245);
nand U3180 (N_3180,N_2896,N_2610);
or U3181 (N_3181,N_2572,N_2818);
nand U3182 (N_3182,N_2885,N_2889);
and U3183 (N_3183,N_2339,N_2484);
and U3184 (N_3184,N_2111,N_2871);
or U3185 (N_3185,N_2454,N_2329);
nor U3186 (N_3186,N_2911,N_2675);
or U3187 (N_3187,N_2985,N_2225);
nor U3188 (N_3188,N_2468,N_2824);
and U3189 (N_3189,N_2674,N_2281);
nor U3190 (N_3190,N_2756,N_2555);
nor U3191 (N_3191,N_2878,N_2975);
and U3192 (N_3192,N_2043,N_2592);
nor U3193 (N_3193,N_2875,N_2387);
nor U3194 (N_3194,N_2874,N_2026);
nor U3195 (N_3195,N_2668,N_2794);
nand U3196 (N_3196,N_2080,N_2987);
nand U3197 (N_3197,N_2890,N_2926);
or U3198 (N_3198,N_2790,N_2840);
nor U3199 (N_3199,N_2672,N_2449);
and U3200 (N_3200,N_2497,N_2010);
and U3201 (N_3201,N_2347,N_2540);
nor U3202 (N_3202,N_2839,N_2370);
or U3203 (N_3203,N_2152,N_2496);
nor U3204 (N_3204,N_2929,N_2260);
or U3205 (N_3205,N_2423,N_2751);
and U3206 (N_3206,N_2422,N_2106);
nand U3207 (N_3207,N_2868,N_2798);
nor U3208 (N_3208,N_2707,N_2015);
nand U3209 (N_3209,N_2150,N_2182);
or U3210 (N_3210,N_2404,N_2479);
or U3211 (N_3211,N_2835,N_2705);
and U3212 (N_3212,N_2068,N_2008);
nor U3213 (N_3213,N_2248,N_2939);
nor U3214 (N_3214,N_2333,N_2562);
nor U3215 (N_3215,N_2425,N_2119);
nand U3216 (N_3216,N_2568,N_2233);
nand U3217 (N_3217,N_2244,N_2266);
nand U3218 (N_3218,N_2321,N_2542);
or U3219 (N_3219,N_2320,N_2622);
and U3220 (N_3220,N_2646,N_2158);
nor U3221 (N_3221,N_2859,N_2398);
nor U3222 (N_3222,N_2793,N_2678);
or U3223 (N_3223,N_2729,N_2699);
or U3224 (N_3224,N_2115,N_2421);
nand U3225 (N_3225,N_2952,N_2727);
nand U3226 (N_3226,N_2613,N_2538);
nor U3227 (N_3227,N_2754,N_2222);
nand U3228 (N_3228,N_2050,N_2821);
and U3229 (N_3229,N_2125,N_2198);
nand U3230 (N_3230,N_2801,N_2031);
and U3231 (N_3231,N_2190,N_2253);
nor U3232 (N_3232,N_2575,N_2647);
or U3233 (N_3233,N_2951,N_2559);
nor U3234 (N_3234,N_2583,N_2581);
nand U3235 (N_3235,N_2982,N_2597);
and U3236 (N_3236,N_2316,N_2660);
or U3237 (N_3237,N_2276,N_2126);
or U3238 (N_3238,N_2061,N_2465);
nand U3239 (N_3239,N_2795,N_2295);
nor U3240 (N_3240,N_2443,N_2891);
nor U3241 (N_3241,N_2297,N_2411);
and U3242 (N_3242,N_2477,N_2977);
nor U3243 (N_3243,N_2916,N_2428);
or U3244 (N_3244,N_2541,N_2078);
and U3245 (N_3245,N_2910,N_2862);
nor U3246 (N_3246,N_2544,N_2967);
nor U3247 (N_3247,N_2407,N_2501);
nor U3248 (N_3248,N_2819,N_2731);
nand U3249 (N_3249,N_2018,N_2028);
nand U3250 (N_3250,N_2215,N_2842);
nand U3251 (N_3251,N_2869,N_2388);
or U3252 (N_3252,N_2512,N_2493);
nor U3253 (N_3253,N_2401,N_2005);
nand U3254 (N_3254,N_2006,N_2805);
or U3255 (N_3255,N_2817,N_2357);
nor U3256 (N_3256,N_2697,N_2199);
and U3257 (N_3257,N_2122,N_2145);
nor U3258 (N_3258,N_2525,N_2359);
nor U3259 (N_3259,N_2779,N_2521);
or U3260 (N_3260,N_2680,N_2441);
or U3261 (N_3261,N_2925,N_2858);
nor U3262 (N_3262,N_2737,N_2691);
nand U3263 (N_3263,N_2591,N_2187);
nor U3264 (N_3264,N_2088,N_2252);
nand U3265 (N_3265,N_2089,N_2070);
or U3266 (N_3266,N_2439,N_2128);
nor U3267 (N_3267,N_2079,N_2962);
nand U3268 (N_3268,N_2774,N_2480);
or U3269 (N_3269,N_2621,N_2250);
nand U3270 (N_3270,N_2524,N_2584);
and U3271 (N_3271,N_2254,N_2094);
and U3272 (N_3272,N_2656,N_2090);
nand U3273 (N_3273,N_2822,N_2463);
and U3274 (N_3274,N_2957,N_2659);
nand U3275 (N_3275,N_2255,N_2579);
or U3276 (N_3276,N_2405,N_2227);
or U3277 (N_3277,N_2980,N_2121);
and U3278 (N_3278,N_2155,N_2041);
xnor U3279 (N_3279,N_2331,N_2825);
or U3280 (N_3280,N_2409,N_2564);
nor U3281 (N_3281,N_2600,N_2397);
nand U3282 (N_3282,N_2337,N_2287);
or U3283 (N_3283,N_2931,N_2294);
or U3284 (N_3284,N_2543,N_2718);
nand U3285 (N_3285,N_2897,N_2408);
and U3286 (N_3286,N_2503,N_2547);
nor U3287 (N_3287,N_2676,N_2380);
nand U3288 (N_3288,N_2192,N_2164);
nor U3289 (N_3289,N_2450,N_2107);
nand U3290 (N_3290,N_2608,N_2334);
nand U3291 (N_3291,N_2476,N_2682);
or U3292 (N_3292,N_2552,N_2201);
nand U3293 (N_3293,N_2461,N_2753);
and U3294 (N_3294,N_2013,N_2765);
or U3295 (N_3295,N_2193,N_2789);
and U3296 (N_3296,N_2095,N_2306);
and U3297 (N_3297,N_2100,N_2533);
nor U3298 (N_3298,N_2171,N_2317);
nand U3299 (N_3299,N_2661,N_2042);
nand U3300 (N_3300,N_2097,N_2550);
and U3301 (N_3301,N_2713,N_2103);
nor U3302 (N_3302,N_2012,N_2983);
or U3303 (N_3303,N_2719,N_2285);
and U3304 (N_3304,N_2303,N_2235);
and U3305 (N_3305,N_2177,N_2865);
or U3306 (N_3306,N_2816,N_2101);
nand U3307 (N_3307,N_2880,N_2744);
and U3308 (N_3308,N_2084,N_2142);
and U3309 (N_3309,N_2553,N_2343);
nand U3310 (N_3310,N_2653,N_2513);
and U3311 (N_3311,N_2213,N_2352);
nand U3312 (N_3312,N_2059,N_2351);
nand U3313 (N_3313,N_2580,N_2472);
and U3314 (N_3314,N_2771,N_2637);
nand U3315 (N_3315,N_2120,N_2694);
or U3316 (N_3316,N_2082,N_2726);
nor U3317 (N_3317,N_2578,N_2261);
and U3318 (N_3318,N_2237,N_2507);
nor U3319 (N_3319,N_2313,N_2998);
nor U3320 (N_3320,N_2539,N_2673);
nand U3321 (N_3321,N_2049,N_2280);
and U3322 (N_3322,N_2234,N_2528);
nor U3323 (N_3323,N_2346,N_2442);
or U3324 (N_3324,N_2703,N_2136);
nor U3325 (N_3325,N_2011,N_2282);
xnor U3326 (N_3326,N_2813,N_2585);
nor U3327 (N_3327,N_2304,N_2170);
nand U3328 (N_3328,N_2272,N_2502);
and U3329 (N_3329,N_2268,N_2867);
nor U3330 (N_3330,N_2545,N_2696);
nor U3331 (N_3331,N_2704,N_2366);
nand U3332 (N_3332,N_2271,N_2024);
and U3333 (N_3333,N_2804,N_2855);
or U3334 (N_3334,N_2833,N_2993);
and U3335 (N_3335,N_2249,N_2060);
nor U3336 (N_3336,N_2087,N_2487);
and U3337 (N_3337,N_2776,N_2912);
nand U3338 (N_3338,N_2523,N_2994);
nor U3339 (N_3339,N_2350,N_2471);
and U3340 (N_3340,N_2400,N_2892);
or U3341 (N_3341,N_2141,N_2978);
nand U3342 (N_3342,N_2203,N_2996);
and U3343 (N_3343,N_2841,N_2489);
xor U3344 (N_3344,N_2139,N_2642);
nand U3345 (N_3345,N_2373,N_2326);
nand U3346 (N_3346,N_2232,N_2866);
nor U3347 (N_3347,N_2027,N_2251);
xnor U3348 (N_3348,N_2566,N_2340);
and U3349 (N_3349,N_2548,N_2344);
or U3350 (N_3350,N_2643,N_2582);
nor U3351 (N_3351,N_2038,N_2626);
nand U3352 (N_3352,N_2654,N_2991);
nand U3353 (N_3353,N_2857,N_2207);
nor U3354 (N_3354,N_2921,N_2590);
nor U3355 (N_3355,N_2051,N_2446);
nor U3356 (N_3356,N_2185,N_2615);
or U3357 (N_3357,N_2901,N_2711);
xnor U3358 (N_3358,N_2053,N_2546);
nand U3359 (N_3359,N_2296,N_2478);
and U3360 (N_3360,N_2686,N_2444);
and U3361 (N_3361,N_2618,N_2919);
or U3362 (N_3362,N_2226,N_2360);
nand U3363 (N_3363,N_2368,N_2194);
nor U3364 (N_3364,N_2289,N_2307);
nand U3365 (N_3365,N_2381,N_2968);
xnor U3366 (N_3366,N_2109,N_2785);
nor U3367 (N_3367,N_2395,N_2636);
nor U3368 (N_3368,N_2961,N_2298);
nand U3369 (N_3369,N_2781,N_2701);
or U3370 (N_3370,N_2735,N_2206);
nor U3371 (N_3371,N_2338,N_2162);
or U3372 (N_3372,N_2658,N_2324);
nor U3373 (N_3373,N_2491,N_2669);
nand U3374 (N_3374,N_2230,N_2877);
and U3375 (N_3375,N_2369,N_2949);
or U3376 (N_3376,N_2893,N_2666);
and U3377 (N_3377,N_2001,N_2532);
or U3378 (N_3378,N_2403,N_2971);
or U3379 (N_3379,N_2293,N_2382);
nor U3380 (N_3380,N_2052,N_2105);
nor U3381 (N_3381,N_2883,N_2574);
or U3382 (N_3382,N_2943,N_2459);
and U3383 (N_3383,N_2739,N_2157);
or U3384 (N_3384,N_2515,N_2906);
and U3385 (N_3385,N_2486,N_2914);
xor U3386 (N_3386,N_2156,N_2264);
or U3387 (N_3387,N_2797,N_2990);
nand U3388 (N_3388,N_2205,N_2399);
and U3389 (N_3389,N_2913,N_2920);
nand U3390 (N_3390,N_2002,N_2301);
and U3391 (N_3391,N_2510,N_2372);
and U3392 (N_3392,N_2195,N_2033);
and U3393 (N_3393,N_2953,N_2356);
or U3394 (N_3394,N_2057,N_2262);
nor U3395 (N_3395,N_2829,N_2113);
and U3396 (N_3396,N_2044,N_2782);
and U3397 (N_3397,N_2780,N_2402);
or U3398 (N_3398,N_2534,N_2760);
nand U3399 (N_3399,N_2029,N_2004);
or U3400 (N_3400,N_2762,N_2180);
and U3401 (N_3401,N_2848,N_2124);
or U3402 (N_3402,N_2536,N_2077);
xnor U3403 (N_3403,N_2616,N_2166);
nand U3404 (N_3404,N_2820,N_2081);
and U3405 (N_3405,N_2665,N_2945);
xor U3406 (N_3406,N_2922,N_2769);
nor U3407 (N_3407,N_2504,N_2071);
and U3408 (N_3408,N_2365,N_2143);
and U3409 (N_3409,N_2127,N_2689);
nand U3410 (N_3410,N_2096,N_2469);
and U3411 (N_3411,N_2149,N_2172);
and U3412 (N_3412,N_2508,N_2623);
or U3413 (N_3413,N_2183,N_2593);
or U3414 (N_3414,N_2576,N_2036);
and U3415 (N_3415,N_2823,N_2184);
nand U3416 (N_3416,N_2065,N_2179);
or U3417 (N_3417,N_2292,N_2518);
nor U3418 (N_3418,N_2217,N_2116);
and U3419 (N_3419,N_2902,N_2830);
or U3420 (N_3420,N_2323,N_2189);
or U3421 (N_3421,N_2837,N_2586);
or U3422 (N_3422,N_2311,N_2847);
and U3423 (N_3423,N_2216,N_2312);
and U3424 (N_3424,N_2200,N_2895);
nor U3425 (N_3425,N_2310,N_2954);
or U3426 (N_3426,N_2607,N_2898);
nand U3427 (N_3427,N_2342,N_2114);
or U3428 (N_3428,N_2601,N_2565);
nor U3429 (N_3429,N_2025,N_2520);
nand U3430 (N_3430,N_2551,N_2860);
or U3431 (N_3431,N_2046,N_2138);
xnor U3432 (N_3432,N_2810,N_2755);
and U3433 (N_3433,N_2757,N_2009);
and U3434 (N_3434,N_2589,N_2927);
nor U3435 (N_3435,N_2700,N_2259);
nor U3436 (N_3436,N_2419,N_2154);
or U3437 (N_3437,N_2882,N_2505);
nor U3438 (N_3438,N_2134,N_2915);
nor U3439 (N_3439,N_2609,N_2300);
and U3440 (N_3440,N_2474,N_2173);
and U3441 (N_3441,N_2956,N_2239);
or U3442 (N_3442,N_2728,N_2843);
nor U3443 (N_3443,N_2137,N_2279);
and U3444 (N_3444,N_2831,N_2159);
or U3445 (N_3445,N_2424,N_2055);
or U3446 (N_3446,N_2440,N_2415);
nor U3447 (N_3447,N_2905,N_2263);
xnor U3448 (N_3448,N_2393,N_2375);
xor U3449 (N_3449,N_2098,N_2687);
or U3450 (N_3450,N_2873,N_2020);
nor U3451 (N_3451,N_2148,N_2064);
or U3452 (N_3452,N_2999,N_2353);
and U3453 (N_3453,N_2749,N_2766);
or U3454 (N_3454,N_2617,N_2808);
nand U3455 (N_3455,N_2485,N_2587);
or U3456 (N_3456,N_2406,N_2706);
nor U3457 (N_3457,N_2186,N_2973);
nand U3458 (N_3458,N_2278,N_2573);
xor U3459 (N_3459,N_2299,N_2458);
nand U3460 (N_3460,N_2305,N_2563);
or U3461 (N_3461,N_2930,N_2969);
and U3462 (N_3462,N_2792,N_2022);
or U3463 (N_3463,N_2734,N_2629);
or U3464 (N_3464,N_2777,N_2635);
or U3465 (N_3465,N_2455,N_2928);
nand U3466 (N_3466,N_2710,N_2567);
and U3467 (N_3467,N_2325,N_2596);
nor U3468 (N_3468,N_2844,N_2023);
nand U3469 (N_3469,N_2241,N_2826);
nand U3470 (N_3470,N_2560,N_2110);
nand U3471 (N_3471,N_2500,N_2770);
nor U3472 (N_3472,N_2030,N_2594);
and U3473 (N_3473,N_2302,N_2228);
nor U3474 (N_3474,N_2349,N_2853);
or U3475 (N_3475,N_2802,N_2432);
and U3476 (N_3476,N_2108,N_2640);
and U3477 (N_3477,N_2362,N_2286);
nand U3478 (N_3478,N_2685,N_2092);
nor U3479 (N_3479,N_2197,N_2988);
nor U3480 (N_3480,N_2863,N_2886);
or U3481 (N_3481,N_2650,N_2231);
nand U3482 (N_3482,N_2056,N_2498);
and U3483 (N_3483,N_2683,N_2788);
and U3484 (N_3484,N_2273,N_2557);
or U3485 (N_3485,N_2328,N_2708);
and U3486 (N_3486,N_2083,N_2445);
or U3487 (N_3487,N_2631,N_2048);
or U3488 (N_3488,N_2379,N_2085);
and U3489 (N_3489,N_2367,N_2130);
and U3490 (N_3490,N_2526,N_2118);
or U3491 (N_3491,N_2569,N_2811);
or U3492 (N_3492,N_2634,N_2384);
and U3493 (N_3493,N_2884,N_2554);
nor U3494 (N_3494,N_2146,N_2984);
nor U3495 (N_3495,N_2570,N_2702);
nand U3496 (N_3496,N_2784,N_2426);
or U3497 (N_3497,N_2679,N_2684);
and U3498 (N_3498,N_2522,N_2283);
and U3499 (N_3499,N_2509,N_2499);
or U3500 (N_3500,N_2091,N_2658);
xor U3501 (N_3501,N_2901,N_2634);
or U3502 (N_3502,N_2733,N_2068);
nor U3503 (N_3503,N_2679,N_2438);
nand U3504 (N_3504,N_2220,N_2279);
nor U3505 (N_3505,N_2810,N_2553);
or U3506 (N_3506,N_2361,N_2399);
nor U3507 (N_3507,N_2467,N_2390);
nor U3508 (N_3508,N_2634,N_2609);
nand U3509 (N_3509,N_2502,N_2354);
nand U3510 (N_3510,N_2140,N_2684);
nor U3511 (N_3511,N_2577,N_2093);
or U3512 (N_3512,N_2808,N_2171);
xnor U3513 (N_3513,N_2962,N_2231);
nand U3514 (N_3514,N_2867,N_2517);
or U3515 (N_3515,N_2067,N_2071);
nand U3516 (N_3516,N_2902,N_2491);
nand U3517 (N_3517,N_2401,N_2174);
and U3518 (N_3518,N_2414,N_2432);
or U3519 (N_3519,N_2702,N_2862);
nor U3520 (N_3520,N_2236,N_2855);
and U3521 (N_3521,N_2336,N_2415);
nand U3522 (N_3522,N_2116,N_2100);
and U3523 (N_3523,N_2913,N_2232);
and U3524 (N_3524,N_2003,N_2487);
and U3525 (N_3525,N_2257,N_2064);
nor U3526 (N_3526,N_2021,N_2881);
and U3527 (N_3527,N_2172,N_2919);
and U3528 (N_3528,N_2658,N_2243);
and U3529 (N_3529,N_2014,N_2875);
or U3530 (N_3530,N_2786,N_2328);
and U3531 (N_3531,N_2926,N_2327);
nor U3532 (N_3532,N_2428,N_2586);
xor U3533 (N_3533,N_2843,N_2061);
nor U3534 (N_3534,N_2457,N_2122);
and U3535 (N_3535,N_2974,N_2784);
and U3536 (N_3536,N_2973,N_2216);
nand U3537 (N_3537,N_2058,N_2958);
nor U3538 (N_3538,N_2332,N_2123);
nand U3539 (N_3539,N_2932,N_2971);
or U3540 (N_3540,N_2571,N_2643);
and U3541 (N_3541,N_2501,N_2680);
or U3542 (N_3542,N_2955,N_2185);
and U3543 (N_3543,N_2412,N_2428);
nor U3544 (N_3544,N_2171,N_2740);
and U3545 (N_3545,N_2291,N_2356);
xor U3546 (N_3546,N_2841,N_2860);
and U3547 (N_3547,N_2735,N_2387);
or U3548 (N_3548,N_2958,N_2990);
nand U3549 (N_3549,N_2697,N_2756);
or U3550 (N_3550,N_2292,N_2044);
and U3551 (N_3551,N_2170,N_2676);
nand U3552 (N_3552,N_2759,N_2474);
nor U3553 (N_3553,N_2035,N_2936);
nand U3554 (N_3554,N_2609,N_2718);
or U3555 (N_3555,N_2855,N_2360);
nor U3556 (N_3556,N_2438,N_2848);
or U3557 (N_3557,N_2848,N_2879);
and U3558 (N_3558,N_2123,N_2748);
nand U3559 (N_3559,N_2498,N_2267);
nand U3560 (N_3560,N_2996,N_2395);
nor U3561 (N_3561,N_2628,N_2644);
nor U3562 (N_3562,N_2478,N_2857);
and U3563 (N_3563,N_2273,N_2326);
xor U3564 (N_3564,N_2394,N_2835);
nand U3565 (N_3565,N_2127,N_2669);
or U3566 (N_3566,N_2946,N_2397);
and U3567 (N_3567,N_2893,N_2906);
and U3568 (N_3568,N_2565,N_2009);
xor U3569 (N_3569,N_2899,N_2225);
xnor U3570 (N_3570,N_2054,N_2853);
nor U3571 (N_3571,N_2280,N_2982);
nor U3572 (N_3572,N_2204,N_2898);
or U3573 (N_3573,N_2661,N_2462);
nand U3574 (N_3574,N_2568,N_2472);
nor U3575 (N_3575,N_2285,N_2482);
nor U3576 (N_3576,N_2851,N_2041);
and U3577 (N_3577,N_2639,N_2709);
nor U3578 (N_3578,N_2615,N_2381);
nand U3579 (N_3579,N_2882,N_2326);
and U3580 (N_3580,N_2149,N_2617);
and U3581 (N_3581,N_2150,N_2553);
and U3582 (N_3582,N_2237,N_2797);
and U3583 (N_3583,N_2907,N_2136);
nand U3584 (N_3584,N_2486,N_2934);
nor U3585 (N_3585,N_2847,N_2205);
and U3586 (N_3586,N_2368,N_2059);
nand U3587 (N_3587,N_2484,N_2759);
nor U3588 (N_3588,N_2488,N_2624);
or U3589 (N_3589,N_2052,N_2043);
xor U3590 (N_3590,N_2289,N_2218);
xnor U3591 (N_3591,N_2129,N_2302);
and U3592 (N_3592,N_2457,N_2117);
and U3593 (N_3593,N_2655,N_2987);
xnor U3594 (N_3594,N_2179,N_2556);
or U3595 (N_3595,N_2775,N_2408);
and U3596 (N_3596,N_2585,N_2270);
or U3597 (N_3597,N_2446,N_2239);
and U3598 (N_3598,N_2110,N_2551);
and U3599 (N_3599,N_2431,N_2617);
nand U3600 (N_3600,N_2063,N_2328);
or U3601 (N_3601,N_2899,N_2890);
nand U3602 (N_3602,N_2118,N_2949);
and U3603 (N_3603,N_2378,N_2103);
or U3604 (N_3604,N_2434,N_2154);
and U3605 (N_3605,N_2073,N_2732);
nor U3606 (N_3606,N_2975,N_2143);
nand U3607 (N_3607,N_2813,N_2308);
and U3608 (N_3608,N_2704,N_2964);
xnor U3609 (N_3609,N_2893,N_2410);
and U3610 (N_3610,N_2474,N_2833);
nand U3611 (N_3611,N_2928,N_2577);
and U3612 (N_3612,N_2481,N_2616);
or U3613 (N_3613,N_2979,N_2673);
nand U3614 (N_3614,N_2783,N_2513);
nor U3615 (N_3615,N_2578,N_2783);
nor U3616 (N_3616,N_2062,N_2709);
xnor U3617 (N_3617,N_2358,N_2595);
or U3618 (N_3618,N_2665,N_2800);
nor U3619 (N_3619,N_2002,N_2324);
and U3620 (N_3620,N_2027,N_2109);
nand U3621 (N_3621,N_2151,N_2436);
or U3622 (N_3622,N_2019,N_2294);
nor U3623 (N_3623,N_2977,N_2804);
or U3624 (N_3624,N_2761,N_2067);
nor U3625 (N_3625,N_2133,N_2182);
nor U3626 (N_3626,N_2722,N_2226);
and U3627 (N_3627,N_2608,N_2307);
or U3628 (N_3628,N_2959,N_2369);
nor U3629 (N_3629,N_2808,N_2868);
or U3630 (N_3630,N_2003,N_2325);
or U3631 (N_3631,N_2121,N_2810);
nor U3632 (N_3632,N_2082,N_2107);
and U3633 (N_3633,N_2386,N_2425);
and U3634 (N_3634,N_2689,N_2269);
or U3635 (N_3635,N_2439,N_2116);
and U3636 (N_3636,N_2978,N_2322);
or U3637 (N_3637,N_2153,N_2417);
xnor U3638 (N_3638,N_2319,N_2918);
nand U3639 (N_3639,N_2586,N_2405);
nand U3640 (N_3640,N_2778,N_2745);
nor U3641 (N_3641,N_2737,N_2286);
nand U3642 (N_3642,N_2939,N_2558);
and U3643 (N_3643,N_2374,N_2186);
xor U3644 (N_3644,N_2220,N_2594);
nand U3645 (N_3645,N_2322,N_2518);
nand U3646 (N_3646,N_2860,N_2481);
nand U3647 (N_3647,N_2172,N_2861);
nand U3648 (N_3648,N_2279,N_2588);
or U3649 (N_3649,N_2314,N_2400);
nand U3650 (N_3650,N_2678,N_2192);
nor U3651 (N_3651,N_2925,N_2125);
nand U3652 (N_3652,N_2504,N_2723);
nand U3653 (N_3653,N_2073,N_2054);
or U3654 (N_3654,N_2795,N_2283);
and U3655 (N_3655,N_2162,N_2296);
or U3656 (N_3656,N_2791,N_2031);
nand U3657 (N_3657,N_2490,N_2331);
or U3658 (N_3658,N_2550,N_2531);
and U3659 (N_3659,N_2948,N_2456);
and U3660 (N_3660,N_2430,N_2688);
nor U3661 (N_3661,N_2799,N_2924);
and U3662 (N_3662,N_2546,N_2933);
or U3663 (N_3663,N_2735,N_2664);
or U3664 (N_3664,N_2255,N_2722);
nor U3665 (N_3665,N_2039,N_2813);
nor U3666 (N_3666,N_2889,N_2507);
and U3667 (N_3667,N_2061,N_2335);
and U3668 (N_3668,N_2489,N_2845);
and U3669 (N_3669,N_2602,N_2194);
nor U3670 (N_3670,N_2733,N_2421);
nand U3671 (N_3671,N_2267,N_2472);
and U3672 (N_3672,N_2613,N_2183);
and U3673 (N_3673,N_2360,N_2085);
nand U3674 (N_3674,N_2155,N_2374);
nor U3675 (N_3675,N_2727,N_2625);
or U3676 (N_3676,N_2138,N_2174);
nand U3677 (N_3677,N_2959,N_2171);
or U3678 (N_3678,N_2864,N_2644);
nor U3679 (N_3679,N_2690,N_2073);
and U3680 (N_3680,N_2063,N_2190);
and U3681 (N_3681,N_2868,N_2946);
nand U3682 (N_3682,N_2859,N_2092);
nand U3683 (N_3683,N_2681,N_2349);
and U3684 (N_3684,N_2506,N_2525);
or U3685 (N_3685,N_2848,N_2639);
nand U3686 (N_3686,N_2674,N_2659);
nand U3687 (N_3687,N_2674,N_2099);
nand U3688 (N_3688,N_2305,N_2053);
and U3689 (N_3689,N_2361,N_2445);
and U3690 (N_3690,N_2689,N_2734);
and U3691 (N_3691,N_2815,N_2233);
or U3692 (N_3692,N_2427,N_2576);
or U3693 (N_3693,N_2445,N_2257);
or U3694 (N_3694,N_2963,N_2145);
or U3695 (N_3695,N_2966,N_2930);
or U3696 (N_3696,N_2083,N_2753);
or U3697 (N_3697,N_2446,N_2646);
and U3698 (N_3698,N_2593,N_2755);
or U3699 (N_3699,N_2621,N_2195);
and U3700 (N_3700,N_2528,N_2901);
and U3701 (N_3701,N_2294,N_2240);
nor U3702 (N_3702,N_2943,N_2583);
or U3703 (N_3703,N_2504,N_2710);
or U3704 (N_3704,N_2073,N_2839);
nand U3705 (N_3705,N_2769,N_2578);
nor U3706 (N_3706,N_2981,N_2861);
nor U3707 (N_3707,N_2979,N_2079);
xor U3708 (N_3708,N_2851,N_2616);
nor U3709 (N_3709,N_2189,N_2531);
or U3710 (N_3710,N_2261,N_2641);
or U3711 (N_3711,N_2667,N_2329);
and U3712 (N_3712,N_2773,N_2876);
nand U3713 (N_3713,N_2267,N_2401);
or U3714 (N_3714,N_2182,N_2279);
and U3715 (N_3715,N_2998,N_2043);
xor U3716 (N_3716,N_2992,N_2167);
nor U3717 (N_3717,N_2620,N_2299);
nand U3718 (N_3718,N_2452,N_2683);
nand U3719 (N_3719,N_2357,N_2500);
nand U3720 (N_3720,N_2278,N_2810);
nand U3721 (N_3721,N_2752,N_2665);
nor U3722 (N_3722,N_2832,N_2176);
nor U3723 (N_3723,N_2723,N_2154);
and U3724 (N_3724,N_2917,N_2408);
or U3725 (N_3725,N_2696,N_2806);
or U3726 (N_3726,N_2508,N_2299);
nor U3727 (N_3727,N_2821,N_2194);
and U3728 (N_3728,N_2681,N_2473);
and U3729 (N_3729,N_2866,N_2905);
xor U3730 (N_3730,N_2762,N_2620);
and U3731 (N_3731,N_2135,N_2527);
nand U3732 (N_3732,N_2201,N_2777);
nand U3733 (N_3733,N_2801,N_2491);
or U3734 (N_3734,N_2190,N_2955);
and U3735 (N_3735,N_2661,N_2229);
nand U3736 (N_3736,N_2968,N_2621);
or U3737 (N_3737,N_2084,N_2178);
and U3738 (N_3738,N_2644,N_2669);
nand U3739 (N_3739,N_2495,N_2703);
xnor U3740 (N_3740,N_2450,N_2612);
nor U3741 (N_3741,N_2525,N_2171);
or U3742 (N_3742,N_2570,N_2541);
nand U3743 (N_3743,N_2552,N_2861);
nand U3744 (N_3744,N_2238,N_2800);
nor U3745 (N_3745,N_2609,N_2583);
or U3746 (N_3746,N_2922,N_2172);
or U3747 (N_3747,N_2678,N_2391);
and U3748 (N_3748,N_2016,N_2810);
xor U3749 (N_3749,N_2564,N_2457);
nand U3750 (N_3750,N_2211,N_2462);
xor U3751 (N_3751,N_2582,N_2912);
nand U3752 (N_3752,N_2297,N_2410);
xor U3753 (N_3753,N_2296,N_2856);
or U3754 (N_3754,N_2218,N_2718);
nand U3755 (N_3755,N_2684,N_2183);
and U3756 (N_3756,N_2638,N_2648);
nor U3757 (N_3757,N_2070,N_2492);
or U3758 (N_3758,N_2352,N_2691);
and U3759 (N_3759,N_2362,N_2810);
and U3760 (N_3760,N_2275,N_2923);
nor U3761 (N_3761,N_2486,N_2218);
nand U3762 (N_3762,N_2223,N_2458);
nand U3763 (N_3763,N_2770,N_2830);
nor U3764 (N_3764,N_2815,N_2117);
and U3765 (N_3765,N_2011,N_2971);
nand U3766 (N_3766,N_2667,N_2965);
or U3767 (N_3767,N_2601,N_2057);
and U3768 (N_3768,N_2348,N_2651);
and U3769 (N_3769,N_2480,N_2428);
nor U3770 (N_3770,N_2583,N_2743);
or U3771 (N_3771,N_2173,N_2328);
nor U3772 (N_3772,N_2523,N_2194);
or U3773 (N_3773,N_2987,N_2359);
nand U3774 (N_3774,N_2013,N_2927);
and U3775 (N_3775,N_2520,N_2368);
and U3776 (N_3776,N_2370,N_2271);
nand U3777 (N_3777,N_2880,N_2774);
xnor U3778 (N_3778,N_2931,N_2494);
nor U3779 (N_3779,N_2923,N_2215);
nor U3780 (N_3780,N_2594,N_2647);
and U3781 (N_3781,N_2842,N_2971);
and U3782 (N_3782,N_2062,N_2422);
nor U3783 (N_3783,N_2543,N_2598);
xnor U3784 (N_3784,N_2356,N_2842);
nand U3785 (N_3785,N_2016,N_2538);
or U3786 (N_3786,N_2542,N_2002);
and U3787 (N_3787,N_2501,N_2199);
nand U3788 (N_3788,N_2344,N_2973);
or U3789 (N_3789,N_2890,N_2695);
nand U3790 (N_3790,N_2210,N_2868);
nor U3791 (N_3791,N_2985,N_2696);
and U3792 (N_3792,N_2437,N_2571);
nand U3793 (N_3793,N_2477,N_2816);
and U3794 (N_3794,N_2068,N_2495);
or U3795 (N_3795,N_2874,N_2849);
nand U3796 (N_3796,N_2171,N_2818);
and U3797 (N_3797,N_2125,N_2611);
nand U3798 (N_3798,N_2653,N_2586);
and U3799 (N_3799,N_2819,N_2471);
nor U3800 (N_3800,N_2409,N_2362);
or U3801 (N_3801,N_2797,N_2040);
and U3802 (N_3802,N_2302,N_2100);
nand U3803 (N_3803,N_2420,N_2827);
or U3804 (N_3804,N_2016,N_2365);
and U3805 (N_3805,N_2137,N_2216);
and U3806 (N_3806,N_2524,N_2144);
and U3807 (N_3807,N_2067,N_2677);
or U3808 (N_3808,N_2402,N_2351);
and U3809 (N_3809,N_2478,N_2725);
or U3810 (N_3810,N_2873,N_2249);
nor U3811 (N_3811,N_2592,N_2760);
or U3812 (N_3812,N_2346,N_2539);
nand U3813 (N_3813,N_2315,N_2755);
or U3814 (N_3814,N_2953,N_2831);
and U3815 (N_3815,N_2184,N_2407);
or U3816 (N_3816,N_2718,N_2584);
or U3817 (N_3817,N_2825,N_2706);
nand U3818 (N_3818,N_2740,N_2911);
xnor U3819 (N_3819,N_2302,N_2598);
and U3820 (N_3820,N_2080,N_2084);
nand U3821 (N_3821,N_2296,N_2270);
and U3822 (N_3822,N_2918,N_2630);
nor U3823 (N_3823,N_2510,N_2450);
or U3824 (N_3824,N_2964,N_2520);
nand U3825 (N_3825,N_2846,N_2108);
or U3826 (N_3826,N_2801,N_2408);
nor U3827 (N_3827,N_2129,N_2911);
nand U3828 (N_3828,N_2600,N_2798);
nand U3829 (N_3829,N_2139,N_2174);
or U3830 (N_3830,N_2132,N_2754);
and U3831 (N_3831,N_2257,N_2039);
nor U3832 (N_3832,N_2691,N_2249);
and U3833 (N_3833,N_2761,N_2598);
and U3834 (N_3834,N_2678,N_2207);
and U3835 (N_3835,N_2432,N_2452);
nand U3836 (N_3836,N_2129,N_2287);
or U3837 (N_3837,N_2596,N_2844);
nor U3838 (N_3838,N_2137,N_2568);
xnor U3839 (N_3839,N_2667,N_2814);
nor U3840 (N_3840,N_2238,N_2752);
nand U3841 (N_3841,N_2757,N_2649);
nor U3842 (N_3842,N_2346,N_2828);
nand U3843 (N_3843,N_2650,N_2267);
nor U3844 (N_3844,N_2977,N_2774);
nor U3845 (N_3845,N_2121,N_2961);
or U3846 (N_3846,N_2772,N_2830);
xor U3847 (N_3847,N_2988,N_2162);
nor U3848 (N_3848,N_2176,N_2462);
and U3849 (N_3849,N_2189,N_2959);
or U3850 (N_3850,N_2302,N_2404);
nand U3851 (N_3851,N_2785,N_2978);
nand U3852 (N_3852,N_2849,N_2064);
or U3853 (N_3853,N_2116,N_2816);
and U3854 (N_3854,N_2446,N_2935);
or U3855 (N_3855,N_2518,N_2496);
and U3856 (N_3856,N_2680,N_2275);
and U3857 (N_3857,N_2502,N_2269);
nor U3858 (N_3858,N_2331,N_2530);
nand U3859 (N_3859,N_2774,N_2263);
or U3860 (N_3860,N_2700,N_2185);
nor U3861 (N_3861,N_2397,N_2010);
or U3862 (N_3862,N_2803,N_2724);
or U3863 (N_3863,N_2943,N_2669);
or U3864 (N_3864,N_2085,N_2528);
nand U3865 (N_3865,N_2317,N_2518);
and U3866 (N_3866,N_2792,N_2750);
or U3867 (N_3867,N_2640,N_2229);
xnor U3868 (N_3868,N_2832,N_2235);
and U3869 (N_3869,N_2036,N_2939);
nor U3870 (N_3870,N_2685,N_2132);
and U3871 (N_3871,N_2803,N_2347);
nor U3872 (N_3872,N_2229,N_2695);
or U3873 (N_3873,N_2516,N_2488);
and U3874 (N_3874,N_2691,N_2879);
or U3875 (N_3875,N_2343,N_2640);
nor U3876 (N_3876,N_2517,N_2608);
xnor U3877 (N_3877,N_2703,N_2759);
and U3878 (N_3878,N_2554,N_2156);
nand U3879 (N_3879,N_2096,N_2037);
or U3880 (N_3880,N_2428,N_2382);
or U3881 (N_3881,N_2857,N_2814);
and U3882 (N_3882,N_2720,N_2028);
nand U3883 (N_3883,N_2223,N_2093);
nand U3884 (N_3884,N_2547,N_2400);
nor U3885 (N_3885,N_2324,N_2891);
nand U3886 (N_3886,N_2338,N_2204);
nor U3887 (N_3887,N_2161,N_2737);
and U3888 (N_3888,N_2511,N_2243);
nand U3889 (N_3889,N_2635,N_2236);
and U3890 (N_3890,N_2322,N_2362);
and U3891 (N_3891,N_2038,N_2458);
nand U3892 (N_3892,N_2192,N_2871);
nor U3893 (N_3893,N_2235,N_2288);
and U3894 (N_3894,N_2139,N_2470);
or U3895 (N_3895,N_2717,N_2413);
nor U3896 (N_3896,N_2695,N_2391);
and U3897 (N_3897,N_2200,N_2074);
xnor U3898 (N_3898,N_2421,N_2420);
or U3899 (N_3899,N_2266,N_2422);
nor U3900 (N_3900,N_2684,N_2922);
and U3901 (N_3901,N_2856,N_2875);
nor U3902 (N_3902,N_2863,N_2118);
nand U3903 (N_3903,N_2374,N_2258);
nand U3904 (N_3904,N_2986,N_2030);
or U3905 (N_3905,N_2514,N_2360);
or U3906 (N_3906,N_2836,N_2970);
or U3907 (N_3907,N_2272,N_2069);
or U3908 (N_3908,N_2366,N_2367);
nand U3909 (N_3909,N_2877,N_2458);
or U3910 (N_3910,N_2058,N_2590);
or U3911 (N_3911,N_2799,N_2609);
nand U3912 (N_3912,N_2531,N_2911);
and U3913 (N_3913,N_2036,N_2966);
nand U3914 (N_3914,N_2550,N_2688);
nor U3915 (N_3915,N_2737,N_2209);
and U3916 (N_3916,N_2000,N_2536);
nor U3917 (N_3917,N_2163,N_2938);
or U3918 (N_3918,N_2100,N_2597);
nand U3919 (N_3919,N_2339,N_2707);
nor U3920 (N_3920,N_2796,N_2648);
and U3921 (N_3921,N_2595,N_2843);
nand U3922 (N_3922,N_2695,N_2497);
or U3923 (N_3923,N_2641,N_2665);
nand U3924 (N_3924,N_2455,N_2274);
nor U3925 (N_3925,N_2512,N_2202);
nand U3926 (N_3926,N_2298,N_2401);
nor U3927 (N_3927,N_2583,N_2875);
nor U3928 (N_3928,N_2667,N_2726);
nand U3929 (N_3929,N_2165,N_2770);
and U3930 (N_3930,N_2714,N_2742);
and U3931 (N_3931,N_2563,N_2632);
or U3932 (N_3932,N_2933,N_2387);
or U3933 (N_3933,N_2789,N_2644);
nor U3934 (N_3934,N_2803,N_2129);
or U3935 (N_3935,N_2034,N_2646);
nand U3936 (N_3936,N_2098,N_2369);
nand U3937 (N_3937,N_2001,N_2764);
nor U3938 (N_3938,N_2383,N_2692);
nor U3939 (N_3939,N_2674,N_2938);
or U3940 (N_3940,N_2600,N_2534);
nor U3941 (N_3941,N_2725,N_2538);
or U3942 (N_3942,N_2082,N_2235);
nand U3943 (N_3943,N_2154,N_2908);
nor U3944 (N_3944,N_2309,N_2952);
nand U3945 (N_3945,N_2981,N_2832);
or U3946 (N_3946,N_2369,N_2950);
or U3947 (N_3947,N_2707,N_2924);
or U3948 (N_3948,N_2951,N_2583);
and U3949 (N_3949,N_2324,N_2272);
and U3950 (N_3950,N_2169,N_2147);
nand U3951 (N_3951,N_2241,N_2120);
nand U3952 (N_3952,N_2043,N_2552);
nor U3953 (N_3953,N_2942,N_2375);
or U3954 (N_3954,N_2249,N_2840);
nand U3955 (N_3955,N_2688,N_2310);
nand U3956 (N_3956,N_2944,N_2460);
or U3957 (N_3957,N_2909,N_2898);
and U3958 (N_3958,N_2976,N_2176);
nand U3959 (N_3959,N_2734,N_2727);
or U3960 (N_3960,N_2813,N_2494);
or U3961 (N_3961,N_2921,N_2855);
nor U3962 (N_3962,N_2249,N_2689);
or U3963 (N_3963,N_2176,N_2124);
or U3964 (N_3964,N_2264,N_2150);
or U3965 (N_3965,N_2936,N_2747);
nand U3966 (N_3966,N_2865,N_2866);
nor U3967 (N_3967,N_2213,N_2109);
nor U3968 (N_3968,N_2721,N_2152);
nor U3969 (N_3969,N_2179,N_2118);
nor U3970 (N_3970,N_2766,N_2930);
and U3971 (N_3971,N_2130,N_2155);
or U3972 (N_3972,N_2605,N_2978);
nand U3973 (N_3973,N_2471,N_2280);
nand U3974 (N_3974,N_2469,N_2189);
nand U3975 (N_3975,N_2412,N_2835);
and U3976 (N_3976,N_2958,N_2029);
or U3977 (N_3977,N_2938,N_2987);
nand U3978 (N_3978,N_2521,N_2315);
or U3979 (N_3979,N_2939,N_2227);
and U3980 (N_3980,N_2716,N_2719);
nor U3981 (N_3981,N_2678,N_2866);
nand U3982 (N_3982,N_2101,N_2062);
nand U3983 (N_3983,N_2609,N_2598);
nand U3984 (N_3984,N_2789,N_2778);
xnor U3985 (N_3985,N_2599,N_2345);
nand U3986 (N_3986,N_2661,N_2782);
and U3987 (N_3987,N_2029,N_2288);
and U3988 (N_3988,N_2038,N_2290);
nor U3989 (N_3989,N_2314,N_2496);
nand U3990 (N_3990,N_2625,N_2607);
and U3991 (N_3991,N_2317,N_2592);
or U3992 (N_3992,N_2555,N_2926);
nor U3993 (N_3993,N_2126,N_2966);
and U3994 (N_3994,N_2113,N_2465);
or U3995 (N_3995,N_2515,N_2443);
and U3996 (N_3996,N_2075,N_2146);
and U3997 (N_3997,N_2682,N_2839);
and U3998 (N_3998,N_2665,N_2722);
nor U3999 (N_3999,N_2327,N_2603);
and U4000 (N_4000,N_3394,N_3661);
nand U4001 (N_4001,N_3400,N_3033);
or U4002 (N_4002,N_3318,N_3582);
and U4003 (N_4003,N_3561,N_3377);
and U4004 (N_4004,N_3922,N_3387);
nor U4005 (N_4005,N_3460,N_3032);
nand U4006 (N_4006,N_3636,N_3774);
or U4007 (N_4007,N_3771,N_3803);
and U4008 (N_4008,N_3601,N_3980);
nand U4009 (N_4009,N_3305,N_3877);
nor U4010 (N_4010,N_3551,N_3874);
or U4011 (N_4011,N_3448,N_3993);
or U4012 (N_4012,N_3667,N_3543);
and U4013 (N_4013,N_3587,N_3221);
and U4014 (N_4014,N_3853,N_3795);
and U4015 (N_4015,N_3609,N_3101);
and U4016 (N_4016,N_3693,N_3258);
nand U4017 (N_4017,N_3140,N_3899);
nand U4018 (N_4018,N_3492,N_3003);
or U4019 (N_4019,N_3674,N_3982);
and U4020 (N_4020,N_3904,N_3730);
or U4021 (N_4021,N_3230,N_3638);
nand U4022 (N_4022,N_3536,N_3040);
nor U4023 (N_4023,N_3580,N_3896);
nor U4024 (N_4024,N_3079,N_3145);
nor U4025 (N_4025,N_3379,N_3490);
nand U4026 (N_4026,N_3268,N_3312);
and U4027 (N_4027,N_3051,N_3444);
nand U4028 (N_4028,N_3298,N_3016);
nand U4029 (N_4029,N_3664,N_3245);
and U4030 (N_4030,N_3184,N_3441);
or U4031 (N_4031,N_3926,N_3030);
and U4032 (N_4032,N_3930,N_3384);
nor U4033 (N_4033,N_3012,N_3205);
or U4034 (N_4034,N_3590,N_3951);
nor U4035 (N_4035,N_3626,N_3341);
nor U4036 (N_4036,N_3246,N_3645);
nand U4037 (N_4037,N_3973,N_3628);
and U4038 (N_4038,N_3884,N_3810);
and U4039 (N_4039,N_3672,N_3261);
or U4040 (N_4040,N_3337,N_3373);
and U4041 (N_4041,N_3871,N_3272);
nor U4042 (N_4042,N_3494,N_3333);
nand U4043 (N_4043,N_3046,N_3112);
and U4044 (N_4044,N_3635,N_3090);
nor U4045 (N_4045,N_3142,N_3686);
nor U4046 (N_4046,N_3928,N_3598);
and U4047 (N_4047,N_3128,N_3507);
or U4048 (N_4048,N_3282,N_3855);
or U4049 (N_4049,N_3329,N_3734);
nor U4050 (N_4050,N_3193,N_3326);
and U4051 (N_4051,N_3447,N_3083);
xnor U4052 (N_4052,N_3866,N_3009);
nand U4053 (N_4053,N_3331,N_3669);
or U4054 (N_4054,N_3278,N_3560);
and U4055 (N_4055,N_3201,N_3036);
nor U4056 (N_4056,N_3822,N_3470);
nand U4057 (N_4057,N_3025,N_3443);
nand U4058 (N_4058,N_3388,N_3087);
or U4059 (N_4059,N_3613,N_3354);
or U4060 (N_4060,N_3809,N_3027);
or U4061 (N_4061,N_3653,N_3017);
nand U4062 (N_4062,N_3089,N_3624);
and U4063 (N_4063,N_3817,N_3961);
or U4064 (N_4064,N_3204,N_3563);
or U4065 (N_4065,N_3621,N_3954);
nor U4066 (N_4066,N_3721,N_3709);
and U4067 (N_4067,N_3405,N_3262);
and U4068 (N_4068,N_3022,N_3981);
nor U4069 (N_4069,N_3106,N_3911);
or U4070 (N_4070,N_3646,N_3562);
and U4071 (N_4071,N_3727,N_3210);
nand U4072 (N_4072,N_3241,N_3066);
and U4073 (N_4073,N_3121,N_3691);
or U4074 (N_4074,N_3117,N_3620);
nor U4075 (N_4075,N_3239,N_3712);
or U4076 (N_4076,N_3720,N_3830);
nand U4077 (N_4077,N_3992,N_3048);
nand U4078 (N_4078,N_3705,N_3081);
and U4079 (N_4079,N_3538,N_3589);
nand U4080 (N_4080,N_3356,N_3419);
nor U4081 (N_4081,N_3486,N_3794);
nor U4082 (N_4082,N_3700,N_3584);
nand U4083 (N_4083,N_3034,N_3556);
or U4084 (N_4084,N_3445,N_3449);
nand U4085 (N_4085,N_3959,N_3429);
xnor U4086 (N_4086,N_3348,N_3127);
nand U4087 (N_4087,N_3599,N_3537);
and U4088 (N_4088,N_3019,N_3767);
or U4089 (N_4089,N_3119,N_3828);
nand U4090 (N_4090,N_3300,N_3832);
or U4091 (N_4091,N_3149,N_3313);
nor U4092 (N_4092,N_3113,N_3276);
or U4093 (N_4093,N_3752,N_3579);
or U4094 (N_4094,N_3895,N_3632);
and U4095 (N_4095,N_3513,N_3948);
and U4096 (N_4096,N_3708,N_3849);
nor U4097 (N_4097,N_3190,N_3931);
or U4098 (N_4098,N_3846,N_3029);
nor U4099 (N_4099,N_3013,N_3857);
nand U4100 (N_4100,N_3126,N_3364);
nor U4101 (N_4101,N_3612,N_3649);
and U4102 (N_4102,N_3411,N_3530);
or U4103 (N_4103,N_3921,N_3330);
nor U4104 (N_4104,N_3963,N_3323);
and U4105 (N_4105,N_3478,N_3055);
or U4106 (N_4106,N_3737,N_3196);
or U4107 (N_4107,N_3296,N_3011);
and U4108 (N_4108,N_3479,N_3656);
and U4109 (N_4109,N_3657,N_3269);
nor U4110 (N_4110,N_3914,N_3380);
and U4111 (N_4111,N_3906,N_3365);
nor U4112 (N_4112,N_3511,N_3283);
xor U4113 (N_4113,N_3985,N_3662);
nand U4114 (N_4114,N_3541,N_3195);
or U4115 (N_4115,N_3988,N_3247);
and U4116 (N_4116,N_3450,N_3726);
nand U4117 (N_4117,N_3848,N_3021);
nor U4118 (N_4118,N_3887,N_3116);
and U4119 (N_4119,N_3728,N_3989);
nor U4120 (N_4120,N_3160,N_3633);
or U4121 (N_4121,N_3243,N_3058);
nand U4122 (N_4122,N_3223,N_3927);
nand U4123 (N_4123,N_3938,N_3177);
or U4124 (N_4124,N_3965,N_3352);
nand U4125 (N_4125,N_3392,N_3234);
or U4126 (N_4126,N_3796,N_3683);
nand U4127 (N_4127,N_3039,N_3173);
nor U4128 (N_4128,N_3566,N_3671);
nand U4129 (N_4129,N_3052,N_3236);
and U4130 (N_4130,N_3153,N_3362);
nor U4131 (N_4131,N_3870,N_3309);
or U4132 (N_4132,N_3383,N_3008);
nor U4133 (N_4133,N_3465,N_3650);
nand U4134 (N_4134,N_3840,N_3607);
nand U4135 (N_4135,N_3968,N_3398);
and U4136 (N_4136,N_3838,N_3781);
nand U4137 (N_4137,N_3357,N_3426);
and U4138 (N_4138,N_3452,N_3102);
xnor U4139 (N_4139,N_3824,N_3964);
nand U4140 (N_4140,N_3756,N_3099);
nor U4141 (N_4141,N_3274,N_3468);
or U4142 (N_4142,N_3944,N_3814);
xor U4143 (N_4143,N_3457,N_3924);
nor U4144 (N_4144,N_3542,N_3422);
or U4145 (N_4145,N_3271,N_3932);
and U4146 (N_4146,N_3018,N_3666);
and U4147 (N_4147,N_3002,N_3403);
and U4148 (N_4148,N_3484,N_3421);
nor U4149 (N_4149,N_3610,N_3835);
or U4150 (N_4150,N_3427,N_3876);
or U4151 (N_4151,N_3044,N_3045);
nand U4152 (N_4152,N_3630,N_3557);
nor U4153 (N_4153,N_3334,N_3361);
and U4154 (N_4154,N_3605,N_3570);
nor U4155 (N_4155,N_3191,N_3676);
nand U4156 (N_4156,N_3049,N_3163);
or U4157 (N_4157,N_3859,N_3792);
nor U4158 (N_4158,N_3120,N_3375);
and U4159 (N_4159,N_3881,N_3094);
nand U4160 (N_4160,N_3722,N_3186);
nand U4161 (N_4161,N_3413,N_3529);
or U4162 (N_4162,N_3769,N_3936);
and U4163 (N_4163,N_3151,N_3496);
nor U4164 (N_4164,N_3521,N_3696);
and U4165 (N_4165,N_3080,N_3885);
and U4166 (N_4166,N_3459,N_3061);
or U4167 (N_4167,N_3138,N_3684);
nor U4168 (N_4168,N_3716,N_3783);
or U4169 (N_4169,N_3615,N_3369);
nand U4170 (N_4170,N_3303,N_3284);
and U4171 (N_4171,N_3606,N_3692);
nand U4172 (N_4172,N_3131,N_3869);
nand U4173 (N_4173,N_3670,N_3146);
or U4174 (N_4174,N_3575,N_3604);
or U4175 (N_4175,N_3368,N_3042);
nand U4176 (N_4176,N_3335,N_3984);
xor U4177 (N_4177,N_3839,N_3436);
or U4178 (N_4178,N_3107,N_3995);
and U4179 (N_4179,N_3719,N_3439);
nor U4180 (N_4180,N_3934,N_3843);
nor U4181 (N_4181,N_3360,N_3169);
xor U4182 (N_4182,N_3353,N_3041);
xnor U4183 (N_4183,N_3808,N_3004);
nand U4184 (N_4184,N_3837,N_3510);
nand U4185 (N_4185,N_3028,N_3209);
nand U4186 (N_4186,N_3109,N_3742);
nand U4187 (N_4187,N_3172,N_3784);
nand U4188 (N_4188,N_3523,N_3553);
nand U4189 (N_4189,N_3315,N_3182);
or U4190 (N_4190,N_3785,N_3732);
or U4191 (N_4191,N_3997,N_3324);
xor U4192 (N_4192,N_3139,N_3455);
and U4193 (N_4193,N_3493,N_3020);
or U4194 (N_4194,N_3372,N_3717);
and U4195 (N_4195,N_3322,N_3873);
and U4196 (N_4196,N_3349,N_3996);
or U4197 (N_4197,N_3043,N_3761);
or U4198 (N_4198,N_3559,N_3949);
and U4199 (N_4199,N_3788,N_3135);
nor U4200 (N_4200,N_3875,N_3897);
nor U4201 (N_4201,N_3189,N_3317);
nor U4202 (N_4202,N_3111,N_3347);
nor U4203 (N_4203,N_3147,N_3483);
nand U4204 (N_4204,N_3277,N_3548);
and U4205 (N_4205,N_3891,N_3180);
nor U4206 (N_4206,N_3962,N_3495);
nand U4207 (N_4207,N_3945,N_3974);
or U4208 (N_4208,N_3156,N_3572);
nand U4209 (N_4209,N_3603,N_3371);
or U4210 (N_4210,N_3110,N_3285);
nor U4211 (N_4211,N_3505,N_3816);
or U4212 (N_4212,N_3807,N_3497);
nor U4213 (N_4213,N_3084,N_3654);
and U4214 (N_4214,N_3697,N_3618);
and U4215 (N_4215,N_3199,N_3161);
or U4216 (N_4216,N_3908,N_3381);
nor U4217 (N_4217,N_3144,N_3047);
and U4218 (N_4218,N_3213,N_3760);
xnor U4219 (N_4219,N_3321,N_3634);
and U4220 (N_4220,N_3759,N_3150);
xor U4221 (N_4221,N_3007,N_3037);
or U4222 (N_4222,N_3917,N_3342);
nor U4223 (N_4223,N_3658,N_3539);
or U4224 (N_4224,N_3202,N_3898);
or U4225 (N_4225,N_3216,N_3753);
nand U4226 (N_4226,N_3776,N_3214);
nand U4227 (N_4227,N_3990,N_3220);
or U4228 (N_4228,N_3772,N_3865);
nand U4229 (N_4229,N_3446,N_3137);
or U4230 (N_4230,N_3533,N_3549);
or U4231 (N_4231,N_3279,N_3660);
nor U4232 (N_4232,N_3229,N_3925);
or U4233 (N_4233,N_3733,N_3095);
and U4234 (N_4234,N_3801,N_3056);
nor U4235 (N_4235,N_3790,N_3332);
and U4236 (N_4236,N_3010,N_3006);
or U4237 (N_4237,N_3291,N_3132);
and U4238 (N_4238,N_3069,N_3763);
nand U4239 (N_4239,N_3292,N_3703);
nor U4240 (N_4240,N_3967,N_3024);
or U4241 (N_4241,N_3585,N_3953);
nand U4242 (N_4242,N_3819,N_3578);
xnor U4243 (N_4243,N_3129,N_3577);
and U4244 (N_4244,N_3503,N_3344);
nor U4245 (N_4245,N_3076,N_3224);
and U4246 (N_4246,N_3860,N_3544);
nand U4247 (N_4247,N_3583,N_3168);
xnor U4248 (N_4248,N_3154,N_3687);
nand U4249 (N_4249,N_3520,N_3892);
nor U4250 (N_4250,N_3273,N_3386);
or U4251 (N_4251,N_3183,N_3937);
nand U4252 (N_4252,N_3957,N_3913);
nor U4253 (N_4253,N_3608,N_3912);
xor U4254 (N_4254,N_3152,N_3404);
or U4255 (N_4255,N_3136,N_3355);
and U4256 (N_4256,N_3569,N_3746);
and U4257 (N_4257,N_3829,N_3251);
nor U4258 (N_4258,N_3237,N_3762);
and U4259 (N_4259,N_3454,N_3038);
or U4260 (N_4260,N_3327,N_3133);
nor U4261 (N_4261,N_3212,N_3339);
nand U4262 (N_4262,N_3698,N_3826);
or U4263 (N_4263,N_3909,N_3690);
and U4264 (N_4264,N_3555,N_3594);
nand U4265 (N_4265,N_3531,N_3242);
nor U4266 (N_4266,N_3304,N_3407);
or U4267 (N_4267,N_3611,N_3713);
nor U4268 (N_4268,N_3438,N_3415);
nor U4269 (N_4269,N_3841,N_3714);
and U4270 (N_4270,N_3155,N_3623);
and U4271 (N_4271,N_3082,N_3588);
and U4272 (N_4272,N_3085,N_3867);
nor U4273 (N_4273,N_3886,N_3310);
nand U4274 (N_4274,N_3343,N_3275);
or U4275 (N_4275,N_3178,N_3677);
and U4276 (N_4276,N_3900,N_3681);
nand U4277 (N_4277,N_3519,N_3975);
and U4278 (N_4278,N_3745,N_3527);
or U4279 (N_4279,N_3319,N_3328);
and U4280 (N_4280,N_3504,N_3652);
and U4281 (N_4281,N_3804,N_3888);
xnor U4282 (N_4282,N_3389,N_3836);
nand U4283 (N_4283,N_3458,N_3882);
nor U4284 (N_4284,N_3518,N_3500);
nor U4285 (N_4285,N_3969,N_3280);
nor U4286 (N_4286,N_3787,N_3098);
or U4287 (N_4287,N_3862,N_3651);
nand U4288 (N_4288,N_3031,N_3971);
nand U4289 (N_4289,N_3092,N_3738);
nand U4290 (N_4290,N_3847,N_3424);
nand U4291 (N_4291,N_3747,N_3266);
nor U4292 (N_4292,N_3983,N_3910);
nand U4293 (N_4293,N_3994,N_3573);
nand U4294 (N_4294,N_3694,N_3440);
and U4295 (N_4295,N_3525,N_3431);
nand U4296 (N_4296,N_3665,N_3167);
nand U4297 (N_4297,N_3782,N_3564);
or U4298 (N_4298,N_3023,N_3831);
or U4299 (N_4299,N_3648,N_3540);
or U4300 (N_4300,N_3907,N_3778);
or U4301 (N_4301,N_3397,N_3935);
nand U4302 (N_4302,N_3616,N_3207);
nand U4303 (N_4303,N_3314,N_3346);
or U4304 (N_4304,N_3073,N_3627);
and U4305 (N_4305,N_3915,N_3845);
or U4306 (N_4306,N_3851,N_3170);
nor U4307 (N_4307,N_3868,N_3554);
nand U4308 (N_4308,N_3115,N_3735);
nor U4309 (N_4309,N_3820,N_3522);
or U4310 (N_4310,N_3487,N_3456);
nor U4311 (N_4311,N_3288,N_3534);
and U4312 (N_4312,N_3200,N_3286);
and U4313 (N_4313,N_3821,N_3729);
nor U4314 (N_4314,N_3358,N_3863);
nand U4315 (N_4315,N_3463,N_3923);
and U4316 (N_4316,N_3192,N_3707);
xnor U4317 (N_4317,N_3059,N_3780);
or U4318 (N_4318,N_3134,N_3679);
nor U4319 (N_4319,N_3515,N_3476);
nor U4320 (N_4320,N_3749,N_3114);
or U4321 (N_4321,N_3395,N_3799);
nor U4322 (N_4322,N_3185,N_3701);
and U4323 (N_4323,N_3015,N_3054);
nand U4324 (N_4324,N_3933,N_3710);
nor U4325 (N_4325,N_3162,N_3471);
nand U4326 (N_4326,N_3755,N_3157);
nor U4327 (N_4327,N_3068,N_3481);
nand U4328 (N_4328,N_3797,N_3402);
or U4329 (N_4329,N_3545,N_3451);
nand U4330 (N_4330,N_3568,N_3437);
nand U4331 (N_4331,N_3420,N_3078);
nor U4332 (N_4332,N_3297,N_3706);
or U4333 (N_4333,N_3225,N_3122);
nand U4334 (N_4334,N_3524,N_3070);
and U4335 (N_4335,N_3528,N_3433);
xnor U4336 (N_4336,N_3725,N_3259);
nor U4337 (N_4337,N_3757,N_3340);
or U4338 (N_4338,N_3077,N_3086);
and U4339 (N_4339,N_3736,N_3668);
nand U4340 (N_4340,N_3567,N_3475);
nand U4341 (N_4341,N_3592,N_3453);
nor U4342 (N_4342,N_3902,N_3754);
nand U4343 (N_4343,N_3104,N_3100);
or U4344 (N_4344,N_3800,N_3485);
xnor U4345 (N_4345,N_3637,N_3806);
or U4346 (N_4346,N_3711,N_3956);
and U4347 (N_4347,N_3724,N_3663);
nor U4348 (N_4348,N_3659,N_3643);
or U4349 (N_4349,N_3072,N_3417);
xnor U4350 (N_4350,N_3267,N_3976);
and U4351 (N_4351,N_3345,N_3103);
and U4352 (N_4352,N_3942,N_3188);
xor U4353 (N_4353,N_3940,N_3219);
and U4354 (N_4354,N_3673,N_3939);
or U4355 (N_4355,N_3593,N_3075);
nand U4356 (N_4356,N_3316,N_3434);
and U4357 (N_4357,N_3978,N_3532);
and U4358 (N_4358,N_3320,N_3215);
nor U4359 (N_4359,N_3743,N_3929);
or U4360 (N_4360,N_3766,N_3306);
nand U4361 (N_4361,N_3057,N_3255);
and U4362 (N_4362,N_3641,N_3695);
or U4363 (N_4363,N_3508,N_3063);
and U4364 (N_4364,N_3864,N_3854);
nand U4365 (N_4365,N_3617,N_3062);
nand U4366 (N_4366,N_3165,N_3217);
nor U4367 (N_4367,N_3702,N_3748);
nand U4368 (N_4368,N_3308,N_3093);
nor U4369 (N_4369,N_3432,N_3805);
or U4370 (N_4370,N_3174,N_3370);
and U4371 (N_4371,N_3442,N_3642);
and U4372 (N_4372,N_3416,N_3802);
nand U4373 (N_4373,N_3770,N_3890);
and U4374 (N_4374,N_3744,N_3249);
or U4375 (N_4375,N_3889,N_3689);
nor U4376 (N_4376,N_3833,N_3464);
and U4377 (N_4377,N_3883,N_3108);
nor U4378 (N_4378,N_3488,N_3194);
nor U4379 (N_4379,N_3685,N_3571);
or U4380 (N_4380,N_3480,N_3252);
nor U4381 (N_4381,N_3960,N_3526);
xnor U4382 (N_4382,N_3894,N_3385);
or U4383 (N_4383,N_3768,N_3629);
nand U4384 (N_4384,N_3901,N_3311);
and U4385 (N_4385,N_3260,N_3461);
nor U4386 (N_4386,N_3430,N_3005);
or U4387 (N_4387,N_3576,N_3655);
nand U4388 (N_4388,N_3158,N_3970);
nand U4389 (N_4389,N_3998,N_3265);
and U4390 (N_4390,N_3740,N_3143);
xnor U4391 (N_4391,N_3105,N_3097);
nor U4392 (N_4392,N_3164,N_3773);
or U4393 (N_4393,N_3903,N_3001);
or U4394 (N_4394,N_3893,N_3823);
nand U4395 (N_4395,N_3071,N_3425);
nand U4396 (N_4396,N_3208,N_3946);
and U4397 (N_4397,N_3535,N_3777);
nand U4398 (N_4398,N_3123,N_3509);
and U4399 (N_4399,N_3999,N_3842);
nand U4400 (N_4400,N_3779,N_3435);
nand U4401 (N_4401,N_3644,N_3264);
and U4402 (N_4402,N_3466,N_3552);
or U4403 (N_4403,N_3197,N_3240);
nand U4404 (N_4404,N_3467,N_3232);
nor U4405 (N_4405,N_3060,N_3293);
nand U4406 (N_4406,N_3250,N_3382);
or U4407 (N_4407,N_3181,N_3401);
nand U4408 (N_4408,N_3764,N_3226);
or U4409 (N_4409,N_3918,N_3235);
and U4410 (N_4410,N_3789,N_3423);
or U4411 (N_4411,N_3558,N_3966);
and U4412 (N_4412,N_3474,N_3750);
nand U4413 (N_4413,N_3299,N_3124);
and U4414 (N_4414,N_3091,N_3813);
nand U4415 (N_4415,N_3675,N_3414);
or U4416 (N_4416,N_3986,N_3614);
nor U4417 (N_4417,N_3597,N_3166);
and U4418 (N_4418,N_3159,N_3639);
and U4419 (N_4419,N_3501,N_3428);
nor U4420 (N_4420,N_3682,N_3281);
nor U4421 (N_4421,N_3253,N_3231);
and U4422 (N_4422,N_3263,N_3919);
and U4423 (N_4423,N_3256,N_3035);
nand U4424 (N_4424,N_3798,N_3818);
and U4425 (N_4425,N_3294,N_3141);
nand U4426 (N_4426,N_3850,N_3053);
nor U4427 (N_4427,N_3491,N_3872);
nand U4428 (N_4428,N_3878,N_3815);
nand U4429 (N_4429,N_3506,N_3751);
or U4430 (N_4430,N_3290,N_3171);
xnor U4431 (N_4431,N_3565,N_3812);
nor U4432 (N_4432,N_3793,N_3958);
nand U4433 (N_4433,N_3574,N_3977);
nor U4434 (N_4434,N_3130,N_3499);
and U4435 (N_4435,N_3858,N_3238);
and U4436 (N_4436,N_3699,N_3410);
or U4437 (N_4437,N_3625,N_3987);
nor U4438 (N_4438,N_3920,N_3880);
nor U4439 (N_4439,N_3739,N_3825);
nor U4440 (N_4440,N_3680,N_3905);
and U4441 (N_4441,N_3175,N_3148);
or U4442 (N_4442,N_3775,N_3391);
nand U4443 (N_4443,N_3363,N_3014);
or U4444 (N_4444,N_3514,N_3955);
or U4445 (N_4445,N_3096,N_3834);
and U4446 (N_4446,N_3118,N_3502);
nor U4447 (N_4447,N_3359,N_3546);
and U4448 (N_4448,N_3991,N_3295);
and U4449 (N_4449,N_3943,N_3254);
and U4450 (N_4450,N_3852,N_3622);
and U4451 (N_4451,N_3301,N_3418);
nand U4452 (N_4452,N_3586,N_3396);
nor U4453 (N_4453,N_3336,N_3489);
or U4454 (N_4454,N_3704,N_3000);
and U4455 (N_4455,N_3947,N_3602);
xor U4456 (N_4456,N_3547,N_3972);
or U4457 (N_4457,N_3325,N_3879);
or U4458 (N_4458,N_3469,N_3950);
nand U4459 (N_4459,N_3600,N_3026);
nor U4460 (N_4460,N_3307,N_3591);
and U4461 (N_4461,N_3856,N_3477);
and U4462 (N_4462,N_3498,N_3257);
and U4463 (N_4463,N_3393,N_3941);
nand U4464 (N_4464,N_3688,N_3064);
or U4465 (N_4465,N_3861,N_3198);
or U4466 (N_4466,N_3203,N_3718);
and U4467 (N_4467,N_3723,N_3916);
nor U4468 (N_4468,N_3065,N_3473);
nand U4469 (N_4469,N_3270,N_3287);
nor U4470 (N_4470,N_3516,N_3376);
and U4471 (N_4471,N_3176,N_3125);
or U4472 (N_4472,N_3179,N_3244);
or U4473 (N_4473,N_3581,N_3765);
and U4474 (N_4474,N_3482,N_3050);
and U4475 (N_4475,N_3222,N_3067);
nand U4476 (N_4476,N_3350,N_3218);
nor U4477 (N_4477,N_3640,N_3302);
nand U4478 (N_4478,N_3399,N_3206);
or U4479 (N_4479,N_3367,N_3731);
nand U4480 (N_4480,N_3517,N_3406);
or U4481 (N_4481,N_3827,N_3619);
and U4482 (N_4482,N_3351,N_3289);
or U4483 (N_4483,N_3472,N_3715);
or U4484 (N_4484,N_3338,N_3390);
nand U4485 (N_4485,N_3550,N_3187);
nor U4486 (N_4486,N_3791,N_3412);
or U4487 (N_4487,N_3647,N_3631);
or U4488 (N_4488,N_3233,N_3366);
or U4489 (N_4489,N_3409,N_3758);
and U4490 (N_4490,N_3512,N_3228);
or U4491 (N_4491,N_3952,N_3088);
or U4492 (N_4492,N_3248,N_3786);
nand U4493 (N_4493,N_3378,N_3811);
nor U4494 (N_4494,N_3227,N_3595);
and U4495 (N_4495,N_3596,N_3074);
nand U4496 (N_4496,N_3741,N_3211);
nand U4497 (N_4497,N_3408,N_3374);
or U4498 (N_4498,N_3678,N_3979);
nor U4499 (N_4499,N_3844,N_3462);
nor U4500 (N_4500,N_3936,N_3948);
nand U4501 (N_4501,N_3584,N_3945);
nand U4502 (N_4502,N_3349,N_3359);
or U4503 (N_4503,N_3848,N_3706);
xnor U4504 (N_4504,N_3002,N_3229);
nand U4505 (N_4505,N_3415,N_3003);
or U4506 (N_4506,N_3338,N_3068);
and U4507 (N_4507,N_3993,N_3144);
nor U4508 (N_4508,N_3234,N_3723);
or U4509 (N_4509,N_3355,N_3351);
nor U4510 (N_4510,N_3382,N_3814);
or U4511 (N_4511,N_3533,N_3269);
or U4512 (N_4512,N_3929,N_3623);
or U4513 (N_4513,N_3810,N_3408);
nor U4514 (N_4514,N_3941,N_3691);
or U4515 (N_4515,N_3055,N_3588);
or U4516 (N_4516,N_3726,N_3363);
or U4517 (N_4517,N_3467,N_3276);
and U4518 (N_4518,N_3428,N_3041);
nand U4519 (N_4519,N_3926,N_3014);
nor U4520 (N_4520,N_3481,N_3776);
and U4521 (N_4521,N_3438,N_3564);
nand U4522 (N_4522,N_3164,N_3071);
nor U4523 (N_4523,N_3390,N_3707);
nand U4524 (N_4524,N_3013,N_3357);
and U4525 (N_4525,N_3130,N_3090);
or U4526 (N_4526,N_3962,N_3666);
nand U4527 (N_4527,N_3295,N_3998);
nand U4528 (N_4528,N_3674,N_3068);
xor U4529 (N_4529,N_3350,N_3513);
and U4530 (N_4530,N_3139,N_3700);
or U4531 (N_4531,N_3897,N_3844);
nand U4532 (N_4532,N_3648,N_3702);
or U4533 (N_4533,N_3169,N_3720);
nor U4534 (N_4534,N_3400,N_3120);
nor U4535 (N_4535,N_3077,N_3537);
nor U4536 (N_4536,N_3711,N_3791);
and U4537 (N_4537,N_3135,N_3074);
nor U4538 (N_4538,N_3947,N_3523);
nand U4539 (N_4539,N_3263,N_3083);
or U4540 (N_4540,N_3492,N_3615);
nand U4541 (N_4541,N_3248,N_3157);
or U4542 (N_4542,N_3903,N_3551);
nand U4543 (N_4543,N_3695,N_3815);
and U4544 (N_4544,N_3775,N_3933);
nand U4545 (N_4545,N_3857,N_3036);
nor U4546 (N_4546,N_3879,N_3459);
or U4547 (N_4547,N_3558,N_3249);
nor U4548 (N_4548,N_3064,N_3800);
nand U4549 (N_4549,N_3868,N_3665);
nand U4550 (N_4550,N_3149,N_3022);
nor U4551 (N_4551,N_3164,N_3343);
nand U4552 (N_4552,N_3566,N_3210);
nand U4553 (N_4553,N_3313,N_3668);
or U4554 (N_4554,N_3665,N_3854);
or U4555 (N_4555,N_3532,N_3419);
and U4556 (N_4556,N_3424,N_3673);
nand U4557 (N_4557,N_3491,N_3970);
or U4558 (N_4558,N_3374,N_3842);
nor U4559 (N_4559,N_3237,N_3455);
and U4560 (N_4560,N_3200,N_3092);
or U4561 (N_4561,N_3809,N_3387);
nand U4562 (N_4562,N_3371,N_3942);
nand U4563 (N_4563,N_3196,N_3286);
or U4564 (N_4564,N_3669,N_3473);
or U4565 (N_4565,N_3690,N_3309);
or U4566 (N_4566,N_3734,N_3272);
or U4567 (N_4567,N_3167,N_3055);
or U4568 (N_4568,N_3097,N_3609);
nor U4569 (N_4569,N_3757,N_3587);
nand U4570 (N_4570,N_3518,N_3480);
nor U4571 (N_4571,N_3248,N_3487);
nor U4572 (N_4572,N_3357,N_3037);
nand U4573 (N_4573,N_3829,N_3296);
nand U4574 (N_4574,N_3076,N_3676);
nor U4575 (N_4575,N_3120,N_3569);
nand U4576 (N_4576,N_3235,N_3168);
and U4577 (N_4577,N_3356,N_3778);
or U4578 (N_4578,N_3864,N_3838);
nor U4579 (N_4579,N_3716,N_3110);
or U4580 (N_4580,N_3818,N_3521);
or U4581 (N_4581,N_3007,N_3253);
nand U4582 (N_4582,N_3593,N_3810);
nand U4583 (N_4583,N_3146,N_3791);
and U4584 (N_4584,N_3929,N_3266);
or U4585 (N_4585,N_3377,N_3911);
xor U4586 (N_4586,N_3842,N_3142);
nand U4587 (N_4587,N_3651,N_3168);
or U4588 (N_4588,N_3221,N_3168);
nand U4589 (N_4589,N_3781,N_3483);
and U4590 (N_4590,N_3642,N_3268);
nand U4591 (N_4591,N_3833,N_3011);
xor U4592 (N_4592,N_3731,N_3835);
nor U4593 (N_4593,N_3728,N_3410);
or U4594 (N_4594,N_3185,N_3394);
or U4595 (N_4595,N_3801,N_3658);
nand U4596 (N_4596,N_3117,N_3005);
nand U4597 (N_4597,N_3900,N_3082);
and U4598 (N_4598,N_3849,N_3641);
and U4599 (N_4599,N_3432,N_3425);
nor U4600 (N_4600,N_3087,N_3352);
nor U4601 (N_4601,N_3912,N_3807);
nand U4602 (N_4602,N_3073,N_3888);
nor U4603 (N_4603,N_3325,N_3551);
and U4604 (N_4604,N_3608,N_3173);
or U4605 (N_4605,N_3161,N_3119);
nand U4606 (N_4606,N_3117,N_3023);
nor U4607 (N_4607,N_3755,N_3807);
and U4608 (N_4608,N_3525,N_3888);
nor U4609 (N_4609,N_3405,N_3072);
nand U4610 (N_4610,N_3287,N_3593);
or U4611 (N_4611,N_3597,N_3850);
and U4612 (N_4612,N_3258,N_3620);
nor U4613 (N_4613,N_3071,N_3373);
or U4614 (N_4614,N_3337,N_3527);
and U4615 (N_4615,N_3114,N_3639);
nand U4616 (N_4616,N_3274,N_3610);
and U4617 (N_4617,N_3552,N_3063);
and U4618 (N_4618,N_3010,N_3571);
nor U4619 (N_4619,N_3015,N_3532);
or U4620 (N_4620,N_3805,N_3240);
xor U4621 (N_4621,N_3828,N_3718);
or U4622 (N_4622,N_3348,N_3479);
nor U4623 (N_4623,N_3438,N_3625);
and U4624 (N_4624,N_3212,N_3817);
and U4625 (N_4625,N_3241,N_3437);
or U4626 (N_4626,N_3501,N_3338);
or U4627 (N_4627,N_3156,N_3044);
nand U4628 (N_4628,N_3021,N_3888);
nand U4629 (N_4629,N_3158,N_3047);
nor U4630 (N_4630,N_3449,N_3588);
nor U4631 (N_4631,N_3999,N_3382);
nor U4632 (N_4632,N_3778,N_3348);
and U4633 (N_4633,N_3565,N_3837);
and U4634 (N_4634,N_3910,N_3970);
or U4635 (N_4635,N_3588,N_3503);
nor U4636 (N_4636,N_3051,N_3048);
nor U4637 (N_4637,N_3103,N_3497);
nand U4638 (N_4638,N_3710,N_3023);
nor U4639 (N_4639,N_3598,N_3594);
and U4640 (N_4640,N_3059,N_3278);
nand U4641 (N_4641,N_3615,N_3240);
nor U4642 (N_4642,N_3102,N_3523);
xnor U4643 (N_4643,N_3916,N_3806);
or U4644 (N_4644,N_3088,N_3685);
or U4645 (N_4645,N_3679,N_3489);
nand U4646 (N_4646,N_3478,N_3162);
or U4647 (N_4647,N_3253,N_3720);
nor U4648 (N_4648,N_3325,N_3186);
or U4649 (N_4649,N_3536,N_3985);
or U4650 (N_4650,N_3377,N_3843);
or U4651 (N_4651,N_3272,N_3835);
nor U4652 (N_4652,N_3742,N_3714);
and U4653 (N_4653,N_3795,N_3021);
nand U4654 (N_4654,N_3734,N_3978);
or U4655 (N_4655,N_3738,N_3937);
nor U4656 (N_4656,N_3653,N_3938);
and U4657 (N_4657,N_3482,N_3737);
and U4658 (N_4658,N_3300,N_3386);
nor U4659 (N_4659,N_3185,N_3730);
and U4660 (N_4660,N_3060,N_3778);
and U4661 (N_4661,N_3087,N_3206);
nor U4662 (N_4662,N_3626,N_3525);
nand U4663 (N_4663,N_3575,N_3795);
nor U4664 (N_4664,N_3571,N_3687);
nor U4665 (N_4665,N_3976,N_3679);
nor U4666 (N_4666,N_3895,N_3253);
nor U4667 (N_4667,N_3086,N_3585);
nand U4668 (N_4668,N_3818,N_3218);
nor U4669 (N_4669,N_3197,N_3597);
or U4670 (N_4670,N_3855,N_3632);
or U4671 (N_4671,N_3059,N_3329);
nor U4672 (N_4672,N_3410,N_3237);
nor U4673 (N_4673,N_3483,N_3008);
nand U4674 (N_4674,N_3345,N_3042);
and U4675 (N_4675,N_3761,N_3171);
or U4676 (N_4676,N_3210,N_3951);
and U4677 (N_4677,N_3881,N_3713);
xor U4678 (N_4678,N_3518,N_3935);
nand U4679 (N_4679,N_3366,N_3866);
nand U4680 (N_4680,N_3911,N_3576);
and U4681 (N_4681,N_3846,N_3082);
or U4682 (N_4682,N_3360,N_3083);
nand U4683 (N_4683,N_3746,N_3518);
nand U4684 (N_4684,N_3254,N_3627);
nor U4685 (N_4685,N_3155,N_3637);
nand U4686 (N_4686,N_3171,N_3585);
nand U4687 (N_4687,N_3166,N_3001);
nor U4688 (N_4688,N_3709,N_3285);
nor U4689 (N_4689,N_3700,N_3776);
or U4690 (N_4690,N_3204,N_3388);
or U4691 (N_4691,N_3578,N_3187);
nor U4692 (N_4692,N_3276,N_3908);
xnor U4693 (N_4693,N_3402,N_3642);
nor U4694 (N_4694,N_3342,N_3118);
or U4695 (N_4695,N_3420,N_3875);
and U4696 (N_4696,N_3443,N_3561);
nor U4697 (N_4697,N_3258,N_3051);
nor U4698 (N_4698,N_3576,N_3992);
or U4699 (N_4699,N_3977,N_3313);
and U4700 (N_4700,N_3356,N_3418);
nor U4701 (N_4701,N_3602,N_3095);
or U4702 (N_4702,N_3810,N_3245);
nor U4703 (N_4703,N_3298,N_3012);
nand U4704 (N_4704,N_3067,N_3317);
nor U4705 (N_4705,N_3428,N_3926);
and U4706 (N_4706,N_3158,N_3653);
nor U4707 (N_4707,N_3646,N_3701);
nor U4708 (N_4708,N_3292,N_3743);
nor U4709 (N_4709,N_3682,N_3878);
nor U4710 (N_4710,N_3209,N_3632);
nand U4711 (N_4711,N_3253,N_3746);
or U4712 (N_4712,N_3351,N_3317);
nor U4713 (N_4713,N_3974,N_3007);
nor U4714 (N_4714,N_3842,N_3324);
or U4715 (N_4715,N_3080,N_3886);
and U4716 (N_4716,N_3076,N_3854);
or U4717 (N_4717,N_3613,N_3696);
nand U4718 (N_4718,N_3264,N_3389);
or U4719 (N_4719,N_3895,N_3550);
nor U4720 (N_4720,N_3280,N_3738);
and U4721 (N_4721,N_3331,N_3037);
nand U4722 (N_4722,N_3068,N_3226);
and U4723 (N_4723,N_3595,N_3114);
or U4724 (N_4724,N_3627,N_3146);
and U4725 (N_4725,N_3981,N_3412);
or U4726 (N_4726,N_3281,N_3878);
and U4727 (N_4727,N_3513,N_3091);
nor U4728 (N_4728,N_3935,N_3762);
or U4729 (N_4729,N_3869,N_3051);
xor U4730 (N_4730,N_3728,N_3898);
and U4731 (N_4731,N_3971,N_3346);
and U4732 (N_4732,N_3836,N_3151);
nand U4733 (N_4733,N_3545,N_3685);
or U4734 (N_4734,N_3693,N_3076);
nor U4735 (N_4735,N_3544,N_3055);
and U4736 (N_4736,N_3135,N_3416);
and U4737 (N_4737,N_3931,N_3519);
xor U4738 (N_4738,N_3136,N_3001);
nand U4739 (N_4739,N_3245,N_3329);
or U4740 (N_4740,N_3044,N_3327);
and U4741 (N_4741,N_3988,N_3689);
and U4742 (N_4742,N_3916,N_3261);
nand U4743 (N_4743,N_3399,N_3104);
nor U4744 (N_4744,N_3704,N_3342);
or U4745 (N_4745,N_3053,N_3003);
nand U4746 (N_4746,N_3049,N_3238);
and U4747 (N_4747,N_3878,N_3139);
nand U4748 (N_4748,N_3254,N_3777);
nand U4749 (N_4749,N_3720,N_3958);
nand U4750 (N_4750,N_3565,N_3550);
nand U4751 (N_4751,N_3400,N_3677);
nor U4752 (N_4752,N_3819,N_3525);
nand U4753 (N_4753,N_3221,N_3445);
nand U4754 (N_4754,N_3920,N_3128);
and U4755 (N_4755,N_3526,N_3332);
nand U4756 (N_4756,N_3547,N_3237);
or U4757 (N_4757,N_3830,N_3431);
nand U4758 (N_4758,N_3596,N_3267);
nand U4759 (N_4759,N_3904,N_3537);
and U4760 (N_4760,N_3779,N_3467);
or U4761 (N_4761,N_3580,N_3543);
and U4762 (N_4762,N_3518,N_3017);
or U4763 (N_4763,N_3847,N_3611);
and U4764 (N_4764,N_3411,N_3101);
nor U4765 (N_4765,N_3616,N_3885);
or U4766 (N_4766,N_3883,N_3534);
and U4767 (N_4767,N_3458,N_3991);
or U4768 (N_4768,N_3004,N_3490);
or U4769 (N_4769,N_3659,N_3720);
nor U4770 (N_4770,N_3302,N_3875);
or U4771 (N_4771,N_3167,N_3428);
nor U4772 (N_4772,N_3851,N_3480);
nor U4773 (N_4773,N_3460,N_3860);
and U4774 (N_4774,N_3639,N_3433);
nand U4775 (N_4775,N_3904,N_3281);
nand U4776 (N_4776,N_3732,N_3667);
nand U4777 (N_4777,N_3176,N_3382);
and U4778 (N_4778,N_3221,N_3273);
or U4779 (N_4779,N_3691,N_3332);
nor U4780 (N_4780,N_3341,N_3507);
and U4781 (N_4781,N_3626,N_3302);
nand U4782 (N_4782,N_3415,N_3693);
and U4783 (N_4783,N_3798,N_3571);
or U4784 (N_4784,N_3457,N_3850);
nand U4785 (N_4785,N_3728,N_3797);
nor U4786 (N_4786,N_3502,N_3072);
or U4787 (N_4787,N_3462,N_3355);
or U4788 (N_4788,N_3755,N_3054);
xor U4789 (N_4789,N_3107,N_3985);
or U4790 (N_4790,N_3446,N_3988);
nor U4791 (N_4791,N_3023,N_3753);
or U4792 (N_4792,N_3476,N_3437);
nor U4793 (N_4793,N_3344,N_3163);
or U4794 (N_4794,N_3717,N_3157);
or U4795 (N_4795,N_3361,N_3179);
and U4796 (N_4796,N_3214,N_3034);
and U4797 (N_4797,N_3583,N_3013);
nand U4798 (N_4798,N_3949,N_3398);
nor U4799 (N_4799,N_3754,N_3711);
nand U4800 (N_4800,N_3920,N_3672);
and U4801 (N_4801,N_3778,N_3282);
nand U4802 (N_4802,N_3245,N_3976);
and U4803 (N_4803,N_3952,N_3810);
nor U4804 (N_4804,N_3487,N_3313);
nor U4805 (N_4805,N_3498,N_3483);
and U4806 (N_4806,N_3592,N_3443);
nor U4807 (N_4807,N_3856,N_3521);
xor U4808 (N_4808,N_3538,N_3084);
and U4809 (N_4809,N_3643,N_3424);
or U4810 (N_4810,N_3088,N_3441);
nor U4811 (N_4811,N_3902,N_3056);
nor U4812 (N_4812,N_3794,N_3962);
nand U4813 (N_4813,N_3295,N_3173);
nand U4814 (N_4814,N_3823,N_3444);
nand U4815 (N_4815,N_3404,N_3073);
or U4816 (N_4816,N_3126,N_3209);
nor U4817 (N_4817,N_3317,N_3749);
and U4818 (N_4818,N_3901,N_3832);
and U4819 (N_4819,N_3407,N_3262);
and U4820 (N_4820,N_3054,N_3831);
nand U4821 (N_4821,N_3546,N_3396);
nand U4822 (N_4822,N_3026,N_3929);
or U4823 (N_4823,N_3087,N_3083);
nand U4824 (N_4824,N_3697,N_3582);
and U4825 (N_4825,N_3171,N_3292);
nand U4826 (N_4826,N_3814,N_3533);
nor U4827 (N_4827,N_3251,N_3432);
and U4828 (N_4828,N_3810,N_3838);
nand U4829 (N_4829,N_3482,N_3315);
and U4830 (N_4830,N_3337,N_3244);
nor U4831 (N_4831,N_3672,N_3609);
and U4832 (N_4832,N_3950,N_3197);
xnor U4833 (N_4833,N_3591,N_3149);
or U4834 (N_4834,N_3046,N_3457);
and U4835 (N_4835,N_3576,N_3384);
and U4836 (N_4836,N_3696,N_3035);
nand U4837 (N_4837,N_3718,N_3239);
nand U4838 (N_4838,N_3731,N_3851);
nor U4839 (N_4839,N_3253,N_3101);
nor U4840 (N_4840,N_3154,N_3649);
nand U4841 (N_4841,N_3092,N_3762);
and U4842 (N_4842,N_3739,N_3468);
nand U4843 (N_4843,N_3816,N_3671);
nand U4844 (N_4844,N_3825,N_3282);
nor U4845 (N_4845,N_3442,N_3667);
or U4846 (N_4846,N_3932,N_3803);
and U4847 (N_4847,N_3309,N_3448);
nor U4848 (N_4848,N_3635,N_3342);
nand U4849 (N_4849,N_3593,N_3920);
xnor U4850 (N_4850,N_3668,N_3325);
or U4851 (N_4851,N_3060,N_3124);
nor U4852 (N_4852,N_3491,N_3893);
nand U4853 (N_4853,N_3900,N_3370);
nor U4854 (N_4854,N_3305,N_3446);
and U4855 (N_4855,N_3652,N_3936);
xor U4856 (N_4856,N_3779,N_3849);
nor U4857 (N_4857,N_3781,N_3720);
or U4858 (N_4858,N_3554,N_3557);
or U4859 (N_4859,N_3586,N_3795);
nand U4860 (N_4860,N_3529,N_3679);
or U4861 (N_4861,N_3853,N_3367);
and U4862 (N_4862,N_3037,N_3320);
nor U4863 (N_4863,N_3255,N_3496);
nor U4864 (N_4864,N_3596,N_3445);
and U4865 (N_4865,N_3581,N_3552);
nor U4866 (N_4866,N_3040,N_3057);
nor U4867 (N_4867,N_3607,N_3426);
nor U4868 (N_4868,N_3254,N_3119);
nand U4869 (N_4869,N_3984,N_3322);
and U4870 (N_4870,N_3687,N_3955);
or U4871 (N_4871,N_3306,N_3096);
xor U4872 (N_4872,N_3441,N_3593);
and U4873 (N_4873,N_3229,N_3868);
nor U4874 (N_4874,N_3676,N_3630);
or U4875 (N_4875,N_3724,N_3690);
or U4876 (N_4876,N_3582,N_3093);
nor U4877 (N_4877,N_3135,N_3109);
nand U4878 (N_4878,N_3663,N_3524);
nor U4879 (N_4879,N_3571,N_3290);
nand U4880 (N_4880,N_3547,N_3721);
nand U4881 (N_4881,N_3940,N_3053);
xor U4882 (N_4882,N_3297,N_3692);
nand U4883 (N_4883,N_3911,N_3279);
nor U4884 (N_4884,N_3113,N_3185);
and U4885 (N_4885,N_3117,N_3368);
xor U4886 (N_4886,N_3988,N_3570);
nand U4887 (N_4887,N_3951,N_3393);
nand U4888 (N_4888,N_3353,N_3134);
nand U4889 (N_4889,N_3982,N_3132);
or U4890 (N_4890,N_3132,N_3953);
or U4891 (N_4891,N_3359,N_3883);
and U4892 (N_4892,N_3899,N_3684);
and U4893 (N_4893,N_3899,N_3574);
nor U4894 (N_4894,N_3259,N_3535);
and U4895 (N_4895,N_3225,N_3535);
and U4896 (N_4896,N_3353,N_3795);
and U4897 (N_4897,N_3235,N_3723);
nand U4898 (N_4898,N_3499,N_3810);
nand U4899 (N_4899,N_3283,N_3838);
nor U4900 (N_4900,N_3907,N_3263);
nor U4901 (N_4901,N_3302,N_3227);
and U4902 (N_4902,N_3879,N_3599);
nand U4903 (N_4903,N_3654,N_3018);
and U4904 (N_4904,N_3524,N_3913);
xnor U4905 (N_4905,N_3650,N_3822);
nand U4906 (N_4906,N_3089,N_3908);
nor U4907 (N_4907,N_3963,N_3732);
and U4908 (N_4908,N_3101,N_3997);
nor U4909 (N_4909,N_3500,N_3745);
or U4910 (N_4910,N_3043,N_3063);
and U4911 (N_4911,N_3394,N_3983);
nor U4912 (N_4912,N_3429,N_3075);
and U4913 (N_4913,N_3284,N_3445);
and U4914 (N_4914,N_3135,N_3063);
and U4915 (N_4915,N_3734,N_3771);
or U4916 (N_4916,N_3583,N_3982);
nand U4917 (N_4917,N_3729,N_3355);
nand U4918 (N_4918,N_3423,N_3572);
xnor U4919 (N_4919,N_3142,N_3809);
or U4920 (N_4920,N_3910,N_3229);
or U4921 (N_4921,N_3439,N_3805);
or U4922 (N_4922,N_3941,N_3952);
nor U4923 (N_4923,N_3571,N_3124);
or U4924 (N_4924,N_3008,N_3917);
nor U4925 (N_4925,N_3395,N_3896);
and U4926 (N_4926,N_3629,N_3101);
and U4927 (N_4927,N_3221,N_3644);
nor U4928 (N_4928,N_3062,N_3426);
or U4929 (N_4929,N_3004,N_3566);
xor U4930 (N_4930,N_3134,N_3368);
and U4931 (N_4931,N_3336,N_3763);
nor U4932 (N_4932,N_3059,N_3889);
nand U4933 (N_4933,N_3768,N_3024);
and U4934 (N_4934,N_3411,N_3365);
nor U4935 (N_4935,N_3030,N_3063);
nand U4936 (N_4936,N_3606,N_3718);
nor U4937 (N_4937,N_3138,N_3947);
nand U4938 (N_4938,N_3191,N_3932);
nor U4939 (N_4939,N_3754,N_3088);
nand U4940 (N_4940,N_3838,N_3969);
nand U4941 (N_4941,N_3947,N_3605);
nand U4942 (N_4942,N_3184,N_3293);
nand U4943 (N_4943,N_3644,N_3620);
or U4944 (N_4944,N_3269,N_3806);
and U4945 (N_4945,N_3950,N_3115);
or U4946 (N_4946,N_3275,N_3902);
nand U4947 (N_4947,N_3631,N_3825);
nor U4948 (N_4948,N_3623,N_3036);
or U4949 (N_4949,N_3554,N_3454);
nand U4950 (N_4950,N_3092,N_3356);
or U4951 (N_4951,N_3682,N_3902);
and U4952 (N_4952,N_3595,N_3752);
nand U4953 (N_4953,N_3665,N_3301);
nand U4954 (N_4954,N_3424,N_3369);
nand U4955 (N_4955,N_3266,N_3873);
nand U4956 (N_4956,N_3844,N_3893);
nand U4957 (N_4957,N_3475,N_3371);
nand U4958 (N_4958,N_3277,N_3862);
nand U4959 (N_4959,N_3785,N_3817);
or U4960 (N_4960,N_3316,N_3857);
nor U4961 (N_4961,N_3257,N_3473);
xor U4962 (N_4962,N_3820,N_3831);
nor U4963 (N_4963,N_3974,N_3890);
and U4964 (N_4964,N_3115,N_3972);
nor U4965 (N_4965,N_3076,N_3970);
or U4966 (N_4966,N_3671,N_3467);
nor U4967 (N_4967,N_3544,N_3172);
or U4968 (N_4968,N_3236,N_3554);
or U4969 (N_4969,N_3957,N_3520);
nand U4970 (N_4970,N_3179,N_3293);
or U4971 (N_4971,N_3959,N_3815);
nand U4972 (N_4972,N_3037,N_3172);
nand U4973 (N_4973,N_3224,N_3699);
and U4974 (N_4974,N_3284,N_3340);
or U4975 (N_4975,N_3017,N_3254);
nand U4976 (N_4976,N_3505,N_3422);
and U4977 (N_4977,N_3766,N_3747);
xnor U4978 (N_4978,N_3506,N_3568);
and U4979 (N_4979,N_3079,N_3059);
nor U4980 (N_4980,N_3619,N_3873);
or U4981 (N_4981,N_3442,N_3904);
nor U4982 (N_4982,N_3113,N_3722);
and U4983 (N_4983,N_3911,N_3817);
or U4984 (N_4984,N_3774,N_3623);
nand U4985 (N_4985,N_3796,N_3190);
nand U4986 (N_4986,N_3470,N_3477);
nand U4987 (N_4987,N_3685,N_3001);
nand U4988 (N_4988,N_3499,N_3764);
or U4989 (N_4989,N_3622,N_3292);
xnor U4990 (N_4990,N_3762,N_3362);
nor U4991 (N_4991,N_3750,N_3343);
and U4992 (N_4992,N_3543,N_3508);
nor U4993 (N_4993,N_3698,N_3444);
nor U4994 (N_4994,N_3141,N_3057);
nor U4995 (N_4995,N_3959,N_3795);
nor U4996 (N_4996,N_3558,N_3496);
nand U4997 (N_4997,N_3807,N_3842);
nor U4998 (N_4998,N_3757,N_3439);
and U4999 (N_4999,N_3624,N_3195);
nand UO_0 (O_0,N_4377,N_4712);
and UO_1 (O_1,N_4122,N_4514);
or UO_2 (O_2,N_4996,N_4944);
nand UO_3 (O_3,N_4287,N_4715);
or UO_4 (O_4,N_4913,N_4663);
or UO_5 (O_5,N_4928,N_4704);
or UO_6 (O_6,N_4464,N_4972);
or UO_7 (O_7,N_4261,N_4963);
nor UO_8 (O_8,N_4306,N_4193);
nand UO_9 (O_9,N_4606,N_4628);
nand UO_10 (O_10,N_4025,N_4175);
nor UO_11 (O_11,N_4503,N_4599);
or UO_12 (O_12,N_4524,N_4227);
or UO_13 (O_13,N_4086,N_4338);
nand UO_14 (O_14,N_4619,N_4866);
xor UO_15 (O_15,N_4266,N_4666);
or UO_16 (O_16,N_4404,N_4310);
or UO_17 (O_17,N_4724,N_4490);
xnor UO_18 (O_18,N_4238,N_4476);
and UO_19 (O_19,N_4284,N_4861);
and UO_20 (O_20,N_4615,N_4991);
or UO_21 (O_21,N_4333,N_4806);
or UO_22 (O_22,N_4090,N_4067);
nand UO_23 (O_23,N_4643,N_4255);
and UO_24 (O_24,N_4061,N_4573);
nor UO_25 (O_25,N_4818,N_4368);
or UO_26 (O_26,N_4700,N_4716);
and UO_27 (O_27,N_4190,N_4066);
nor UO_28 (O_28,N_4869,N_4384);
and UO_29 (O_29,N_4118,N_4096);
and UO_30 (O_30,N_4920,N_4785);
nand UO_31 (O_31,N_4760,N_4722);
xnor UO_32 (O_32,N_4985,N_4537);
or UO_33 (O_33,N_4016,N_4923);
xor UO_34 (O_34,N_4951,N_4426);
nand UO_35 (O_35,N_4520,N_4626);
and UO_36 (O_36,N_4607,N_4932);
or UO_37 (O_37,N_4186,N_4660);
or UO_38 (O_38,N_4301,N_4917);
and UO_39 (O_39,N_4883,N_4587);
nand UO_40 (O_40,N_4059,N_4511);
and UO_41 (O_41,N_4056,N_4269);
and UO_42 (O_42,N_4813,N_4640);
and UO_43 (O_43,N_4735,N_4062);
and UO_44 (O_44,N_4082,N_4801);
nor UO_45 (O_45,N_4814,N_4230);
nand UO_46 (O_46,N_4406,N_4938);
nor UO_47 (O_47,N_4205,N_4480);
or UO_48 (O_48,N_4455,N_4325);
or UO_49 (O_49,N_4459,N_4671);
nand UO_50 (O_50,N_4054,N_4342);
or UO_51 (O_51,N_4177,N_4199);
and UO_52 (O_52,N_4746,N_4627);
and UO_53 (O_53,N_4576,N_4994);
and UO_54 (O_54,N_4579,N_4945);
nor UO_55 (O_55,N_4931,N_4609);
and UO_56 (O_56,N_4100,N_4302);
nor UO_57 (O_57,N_4577,N_4827);
nand UO_58 (O_58,N_4611,N_4113);
and UO_59 (O_59,N_4151,N_4367);
and UO_60 (O_60,N_4967,N_4895);
and UO_61 (O_61,N_4303,N_4437);
and UO_62 (O_62,N_4389,N_4027);
nor UO_63 (O_63,N_4852,N_4934);
nor UO_64 (O_64,N_4892,N_4010);
nand UO_65 (O_65,N_4973,N_4800);
and UO_66 (O_66,N_4851,N_4115);
or UO_67 (O_67,N_4204,N_4231);
nor UO_68 (O_68,N_4905,N_4574);
or UO_69 (O_69,N_4992,N_4962);
and UO_70 (O_70,N_4557,N_4784);
or UO_71 (O_71,N_4629,N_4262);
nor UO_72 (O_72,N_4946,N_4289);
or UO_73 (O_73,N_4327,N_4335);
nand UO_74 (O_74,N_4085,N_4670);
and UO_75 (O_75,N_4645,N_4114);
and UO_76 (O_76,N_4634,N_4353);
nand UO_77 (O_77,N_4295,N_4949);
or UO_78 (O_78,N_4065,N_4652);
or UO_79 (O_79,N_4947,N_4469);
nand UO_80 (O_80,N_4228,N_4064);
nor UO_81 (O_81,N_4235,N_4635);
and UO_82 (O_82,N_4694,N_4549);
xnor UO_83 (O_83,N_4942,N_4309);
or UO_84 (O_84,N_4154,N_4969);
nand UO_85 (O_85,N_4271,N_4641);
or UO_86 (O_86,N_4896,N_4134);
nor UO_87 (O_87,N_4446,N_4732);
or UO_88 (O_88,N_4349,N_4457);
and UO_89 (O_89,N_4174,N_4103);
nor UO_90 (O_90,N_4968,N_4201);
nand UO_91 (O_91,N_4270,N_4378);
or UO_92 (O_92,N_4790,N_4195);
nand UO_93 (O_93,N_4868,N_4570);
xnor UO_94 (O_94,N_4127,N_4144);
and UO_95 (O_95,N_4173,N_4246);
or UO_96 (O_96,N_4959,N_4636);
and UO_97 (O_97,N_4534,N_4850);
and UO_98 (O_98,N_4493,N_4372);
nand UO_99 (O_99,N_4362,N_4374);
nand UO_100 (O_100,N_4559,N_4849);
nor UO_101 (O_101,N_4009,N_4902);
nor UO_102 (O_102,N_4546,N_4754);
nand UO_103 (O_103,N_4621,N_4239);
or UO_104 (O_104,N_4111,N_4854);
nand UO_105 (O_105,N_4075,N_4717);
nor UO_106 (O_106,N_4624,N_4099);
and UO_107 (O_107,N_4728,N_4145);
nor UO_108 (O_108,N_4128,N_4202);
nor UO_109 (O_109,N_4657,N_4795);
xnor UO_110 (O_110,N_4882,N_4763);
and UO_111 (O_111,N_4681,N_4598);
or UO_112 (O_112,N_4444,N_4799);
nor UO_113 (O_113,N_4453,N_4815);
or UO_114 (O_114,N_4729,N_4108);
or UO_115 (O_115,N_4220,N_4417);
nor UO_116 (O_116,N_4519,N_4502);
nand UO_117 (O_117,N_4523,N_4345);
nor UO_118 (O_118,N_4069,N_4981);
or UO_119 (O_119,N_4304,N_4460);
xor UO_120 (O_120,N_4176,N_4680);
or UO_121 (O_121,N_4679,N_4562);
and UO_122 (O_122,N_4727,N_4730);
nor UO_123 (O_123,N_4178,N_4780);
or UO_124 (O_124,N_4165,N_4129);
nand UO_125 (O_125,N_4567,N_4209);
and UO_126 (O_126,N_4617,N_4846);
nand UO_127 (O_127,N_4839,N_4288);
and UO_128 (O_128,N_4792,N_4102);
or UO_129 (O_129,N_4881,N_4402);
nor UO_130 (O_130,N_4263,N_4560);
nand UO_131 (O_131,N_4131,N_4019);
nor UO_132 (O_132,N_4070,N_4646);
nor UO_133 (O_133,N_4488,N_4484);
xor UO_134 (O_134,N_4221,N_4467);
and UO_135 (O_135,N_4112,N_4168);
and UO_136 (O_136,N_4419,N_4192);
nor UO_137 (O_137,N_4862,N_4995);
nand UO_138 (O_138,N_4157,N_4907);
nor UO_139 (O_139,N_4369,N_4012);
nor UO_140 (O_140,N_4498,N_4471);
nand UO_141 (O_141,N_4136,N_4911);
or UO_142 (O_142,N_4890,N_4217);
nand UO_143 (O_143,N_4508,N_4653);
or UO_144 (O_144,N_4473,N_4757);
or UO_145 (O_145,N_4743,N_4358);
nand UO_146 (O_146,N_4448,N_4739);
or UO_147 (O_147,N_4501,N_4361);
xor UO_148 (O_148,N_4713,N_4485);
or UO_149 (O_149,N_4966,N_4738);
nand UO_150 (O_150,N_4030,N_4472);
nor UO_151 (O_151,N_4400,N_4871);
or UO_152 (O_152,N_4328,N_4590);
or UO_153 (O_153,N_4161,N_4989);
and UO_154 (O_154,N_4407,N_4443);
and UO_155 (O_155,N_4535,N_4873);
and UO_156 (O_156,N_4495,N_4420);
nor UO_157 (O_157,N_4410,N_4006);
and UO_158 (O_158,N_4999,N_4647);
and UO_159 (O_159,N_4935,N_4505);
or UO_160 (O_160,N_4053,N_4462);
or UO_161 (O_161,N_4213,N_4433);
or UO_162 (O_162,N_4551,N_4036);
and UO_163 (O_163,N_4139,N_4983);
nor UO_164 (O_164,N_4847,N_4399);
nor UO_165 (O_165,N_4817,N_4380);
nor UO_166 (O_166,N_4774,N_4661);
and UO_167 (O_167,N_4656,N_4980);
or UO_168 (O_168,N_4897,N_4838);
nand UO_169 (O_169,N_4334,N_4805);
nand UO_170 (O_170,N_4564,N_4770);
or UO_171 (O_171,N_4719,N_4418);
nand UO_172 (O_172,N_4918,N_4809);
or UO_173 (O_173,N_4084,N_4642);
and UO_174 (O_174,N_4702,N_4563);
or UO_175 (O_175,N_4997,N_4341);
nor UO_176 (O_176,N_4572,N_4241);
nor UO_177 (O_177,N_4783,N_4842);
nor UO_178 (O_178,N_4547,N_4058);
or UO_179 (O_179,N_4180,N_4987);
or UO_180 (O_180,N_4299,N_4648);
and UO_181 (O_181,N_4143,N_4941);
and UO_182 (O_182,N_4394,N_4939);
or UO_183 (O_183,N_4740,N_4706);
nor UO_184 (O_184,N_4900,N_4366);
or UO_185 (O_185,N_4509,N_4046);
or UO_186 (O_186,N_4028,N_4899);
or UO_187 (O_187,N_4593,N_4474);
and UO_188 (O_188,N_4592,N_4222);
and UO_189 (O_189,N_4252,N_4610);
or UO_190 (O_190,N_4290,N_4786);
or UO_191 (O_191,N_4167,N_4580);
and UO_192 (O_192,N_4893,N_4605);
or UO_193 (O_193,N_4080,N_4015);
nand UO_194 (O_194,N_4424,N_4856);
and UO_195 (O_195,N_4933,N_4211);
or UO_196 (O_196,N_4033,N_4014);
nand UO_197 (O_197,N_4050,N_4658);
nor UO_198 (O_198,N_4575,N_4521);
nor UO_199 (O_199,N_4264,N_4007);
and UO_200 (O_200,N_4477,N_4747);
nor UO_201 (O_201,N_4737,N_4240);
nand UO_202 (O_202,N_4285,N_4098);
nor UO_203 (O_203,N_4398,N_4779);
nand UO_204 (O_204,N_4595,N_4874);
nand UO_205 (O_205,N_4820,N_4614);
nor UO_206 (O_206,N_4319,N_4764);
nand UO_207 (O_207,N_4164,N_4215);
nor UO_208 (O_208,N_4278,N_4330);
or UO_209 (O_209,N_4482,N_4692);
and UO_210 (O_210,N_4990,N_4736);
or UO_211 (O_211,N_4507,N_4216);
nand UO_212 (O_212,N_4499,N_4245);
nor UO_213 (O_213,N_4170,N_4206);
nor UO_214 (O_214,N_4860,N_4365);
or UO_215 (O_215,N_4031,N_4710);
and UO_216 (O_216,N_4583,N_4940);
nand UO_217 (O_217,N_4068,N_4669);
and UO_218 (O_218,N_4916,N_4582);
and UO_219 (O_219,N_4773,N_4589);
nand UO_220 (O_220,N_4396,N_4588);
nand UO_221 (O_221,N_4275,N_4376);
or UO_222 (O_222,N_4352,N_4359);
or UO_223 (O_223,N_4516,N_4682);
nor UO_224 (O_224,N_4872,N_4123);
nand UO_225 (O_225,N_4234,N_4057);
nor UO_226 (O_226,N_4711,N_4863);
or UO_227 (O_227,N_4789,N_4355);
and UO_228 (O_228,N_4357,N_4542);
or UO_229 (O_229,N_4055,N_4531);
nor UO_230 (O_230,N_4777,N_4385);
and UO_231 (O_231,N_4875,N_4162);
nor UO_232 (O_232,N_4137,N_4859);
nand UO_233 (O_233,N_4494,N_4117);
or UO_234 (O_234,N_4841,N_4320);
or UO_235 (O_235,N_4707,N_4052);
or UO_236 (O_236,N_4926,N_4581);
and UO_237 (O_237,N_4458,N_4930);
nor UO_238 (O_238,N_4370,N_4725);
nand UO_239 (O_239,N_4533,N_4836);
nor UO_240 (O_240,N_4884,N_4898);
or UO_241 (O_241,N_4919,N_4078);
and UO_242 (O_242,N_4155,N_4925);
nand UO_243 (O_243,N_4116,N_4004);
and UO_244 (O_244,N_4639,N_4037);
or UO_245 (O_245,N_4512,N_4133);
nand UO_246 (O_246,N_4927,N_4705);
and UO_247 (O_247,N_4011,N_4260);
and UO_248 (O_248,N_4522,N_4771);
nand UO_249 (O_249,N_4960,N_4584);
or UO_250 (O_250,N_4699,N_4237);
nand UO_251 (O_251,N_4936,N_4314);
and UO_252 (O_252,N_4796,N_4254);
and UO_253 (O_253,N_4687,N_4423);
or UO_254 (O_254,N_4431,N_4421);
nor UO_255 (O_255,N_4432,N_4776);
nand UO_256 (O_256,N_4553,N_4486);
nand UO_257 (O_257,N_4879,N_4819);
nor UO_258 (O_258,N_4544,N_4038);
or UO_259 (O_259,N_4637,N_4071);
nor UO_260 (O_260,N_4908,N_4701);
and UO_261 (O_261,N_4409,N_4929);
or UO_262 (O_262,N_4219,N_4998);
and UO_263 (O_263,N_4293,N_4076);
nand UO_264 (O_264,N_4625,N_4447);
nor UO_265 (O_265,N_4974,N_4571);
and UO_266 (O_266,N_4844,N_4371);
or UO_267 (O_267,N_4840,N_4673);
nand UO_268 (O_268,N_4184,N_4346);
nor UO_269 (O_269,N_4307,N_4708);
nor UO_270 (O_270,N_4022,N_4121);
or UO_271 (O_271,N_4709,N_4388);
nor UO_272 (O_272,N_4977,N_4802);
nand UO_273 (O_273,N_4984,N_4250);
and UO_274 (O_274,N_4104,N_4650);
and UO_275 (O_275,N_4752,N_4953);
nand UO_276 (O_276,N_4318,N_4470);
or UO_277 (O_277,N_4718,N_4315);
xnor UO_278 (O_278,N_4042,N_4449);
nand UO_279 (O_279,N_4665,N_4568);
or UO_280 (O_280,N_4837,N_4001);
or UO_281 (O_281,N_4343,N_4613);
or UO_282 (O_282,N_4397,N_4183);
or UO_283 (O_283,N_4094,N_4914);
or UO_284 (O_284,N_4405,N_4703);
nand UO_285 (O_285,N_4363,N_4691);
or UO_286 (O_286,N_4922,N_4768);
nor UO_287 (O_287,N_4630,N_4158);
or UO_288 (O_288,N_4224,N_4878);
and UO_289 (O_289,N_4045,N_4829);
and UO_290 (O_290,N_4734,N_4294);
nand UO_291 (O_291,N_4857,N_4350);
and UO_292 (O_292,N_4616,N_4159);
nor UO_293 (O_293,N_4281,N_4243);
nor UO_294 (O_294,N_4552,N_4268);
and UO_295 (O_295,N_4889,N_4283);
or UO_296 (O_296,N_4412,N_4324);
or UO_297 (O_297,N_4244,N_4257);
and UO_298 (O_298,N_4620,N_4688);
nor UO_299 (O_299,N_4504,N_4020);
nand UO_300 (O_300,N_4379,N_4487);
nand UO_301 (O_301,N_4638,N_4955);
or UO_302 (O_302,N_4748,N_4525);
or UO_303 (O_303,N_4169,N_4539);
nand UO_304 (O_304,N_4769,N_4182);
or UO_305 (O_305,N_4690,N_4608);
and UO_306 (O_306,N_4612,N_4017);
nand UO_307 (O_307,N_4513,N_4744);
nand UO_308 (O_308,N_4714,N_4408);
or UO_309 (O_309,N_4329,N_4074);
and UO_310 (O_310,N_4340,N_4381);
nor UO_311 (O_311,N_4903,N_4877);
nand UO_312 (O_312,N_4492,N_4282);
nand UO_313 (O_313,N_4695,N_4781);
and UO_314 (O_314,N_4259,N_4092);
nor UO_315 (O_315,N_4073,N_4021);
nand UO_316 (O_316,N_4043,N_4142);
and UO_317 (O_317,N_4886,N_4256);
or UO_318 (O_318,N_4870,N_4978);
and UO_319 (O_319,N_4454,N_4957);
or UO_320 (O_320,N_4354,N_4596);
nor UO_321 (O_321,N_4632,N_4803);
and UO_322 (O_322,N_4496,N_4876);
or UO_323 (O_323,N_4326,N_4292);
or UO_324 (O_324,N_4489,N_4152);
nor UO_325 (O_325,N_4214,N_4047);
nand UO_326 (O_326,N_4697,N_4880);
and UO_327 (O_327,N_4600,N_4003);
or UO_328 (O_328,N_4060,N_4272);
or UO_329 (O_329,N_4253,N_4988);
or UO_330 (O_330,N_4664,N_4654);
and UO_331 (O_331,N_4440,N_4438);
nor UO_332 (O_332,N_4644,N_4604);
and UO_333 (O_333,N_4591,N_4811);
or UO_334 (O_334,N_4415,N_4950);
and UO_335 (O_335,N_4382,N_4517);
and UO_336 (O_336,N_4149,N_4403);
xor UO_337 (O_337,N_4226,N_4478);
nand UO_338 (O_338,N_4236,N_4207);
nor UO_339 (O_339,N_4348,N_4723);
or UO_340 (O_340,N_4312,N_4291);
nor UO_341 (O_341,N_4203,N_4982);
and UO_342 (O_342,N_4594,N_4762);
or UO_343 (O_343,N_4297,N_4197);
nor UO_344 (O_344,N_4126,N_4441);
nand UO_345 (O_345,N_4035,N_4364);
and UO_346 (O_346,N_4427,N_4623);
and UO_347 (O_347,N_4798,N_4585);
nor UO_348 (O_348,N_4466,N_4434);
or UO_349 (O_349,N_4566,N_4156);
and UO_350 (O_350,N_4993,N_4778);
nor UO_351 (O_351,N_4049,N_4249);
nor UO_352 (O_352,N_4891,N_4565);
nand UO_353 (O_353,N_4451,N_4845);
nand UO_354 (O_354,N_4834,N_4888);
or UO_355 (O_355,N_4649,N_4824);
nand UO_356 (O_356,N_4087,N_4097);
nand UO_357 (O_357,N_4414,N_4631);
nand UO_358 (O_358,N_4541,N_4185);
xnor UO_359 (O_359,N_4475,N_4924);
xor UO_360 (O_360,N_4825,N_4586);
or UO_361 (O_361,N_4425,N_4251);
nand UO_362 (O_362,N_4741,N_4767);
or UO_363 (O_363,N_4005,N_4428);
nand UO_364 (O_364,N_4390,N_4558);
and UO_365 (O_365,N_4810,N_4088);
and UO_366 (O_366,N_4435,N_4543);
or UO_367 (O_367,N_4360,N_4279);
and UO_368 (O_368,N_4233,N_4976);
nand UO_369 (O_369,N_4336,N_4393);
nor UO_370 (O_370,N_4450,N_4826);
nand UO_371 (O_371,N_4305,N_4041);
xnor UO_372 (O_372,N_4667,N_4659);
nor UO_373 (O_373,N_4160,N_4051);
or UO_374 (O_374,N_4759,N_4823);
nand UO_375 (O_375,N_4677,N_4797);
and UO_376 (O_376,N_4461,N_4756);
or UO_377 (O_377,N_4110,N_4830);
nand UO_378 (O_378,N_4528,N_4300);
nand UO_379 (O_379,N_4242,N_4812);
or UO_380 (O_380,N_4698,N_4506);
or UO_381 (O_381,N_4039,N_4124);
and UO_382 (O_382,N_4411,N_4497);
and UO_383 (O_383,N_4029,N_4316);
or UO_384 (O_384,N_4855,N_4527);
nand UO_385 (O_385,N_4848,N_4791);
or UO_386 (O_386,N_4150,N_4597);
nor UO_387 (O_387,N_4745,N_4675);
nand UO_388 (O_388,N_4970,N_4008);
nand UO_389 (O_389,N_4858,N_4678);
or UO_390 (O_390,N_4548,N_4132);
xnor UO_391 (O_391,N_4761,N_4954);
nor UO_392 (O_392,N_4794,N_4463);
nor UO_393 (O_393,N_4120,N_4906);
and UO_394 (O_394,N_4172,N_4821);
or UO_395 (O_395,N_4040,N_4072);
and UO_396 (O_396,N_4089,N_4833);
and UO_397 (O_397,N_4693,N_4672);
and UO_398 (O_398,N_4422,N_4550);
nand UO_399 (O_399,N_4832,N_4750);
nor UO_400 (O_400,N_4171,N_4212);
and UO_401 (O_401,N_4958,N_4146);
and UO_402 (O_402,N_4948,N_4188);
nor UO_403 (O_403,N_4018,N_4223);
nand UO_404 (O_404,N_4835,N_4296);
xnor UO_405 (O_405,N_4375,N_4483);
and UO_406 (O_406,N_4179,N_4141);
nor UO_407 (O_407,N_4952,N_4187);
and UO_408 (O_408,N_4742,N_4125);
or UO_409 (O_409,N_4383,N_4332);
nor UO_410 (O_410,N_4258,N_4696);
nor UO_411 (O_411,N_4265,N_4442);
or UO_412 (O_412,N_4048,N_4273);
or UO_413 (O_413,N_4119,N_4392);
nor UO_414 (O_414,N_4445,N_4232);
nor UO_415 (O_415,N_4063,N_4532);
or UO_416 (O_416,N_4194,N_4210);
or UO_417 (O_417,N_4721,N_4726);
nand UO_418 (O_418,N_4965,N_4106);
nand UO_419 (O_419,N_4676,N_4196);
nand UO_420 (O_420,N_4308,N_4788);
nand UO_421 (O_421,N_4248,N_4822);
nand UO_422 (O_422,N_4356,N_4387);
or UO_423 (O_423,N_4655,N_4468);
nand UO_424 (O_424,N_4023,N_4865);
nor UO_425 (O_425,N_4000,N_4910);
and UO_426 (O_426,N_4373,N_4828);
or UO_427 (O_427,N_4083,N_4135);
and UO_428 (O_428,N_4943,N_4733);
or UO_429 (O_429,N_4816,N_4554);
and UO_430 (O_430,N_4218,N_4286);
and UO_431 (O_431,N_4166,N_4140);
nand UO_432 (O_432,N_4191,N_4843);
or UO_433 (O_433,N_4569,N_4130);
nor UO_434 (O_434,N_4321,N_4298);
or UO_435 (O_435,N_4093,N_4685);
or UO_436 (O_436,N_4530,N_4971);
or UO_437 (O_437,N_4602,N_4720);
nor UO_438 (O_438,N_4351,N_4322);
nor UO_439 (O_439,N_4429,N_4515);
and UO_440 (O_440,N_4684,N_4200);
nand UO_441 (O_441,N_4979,N_4456);
or UO_442 (O_442,N_4311,N_4079);
nor UO_443 (O_443,N_4081,N_4651);
nand UO_444 (O_444,N_4975,N_4904);
or UO_445 (O_445,N_4526,N_4793);
nand UO_446 (O_446,N_4095,N_4561);
or UO_447 (O_447,N_4804,N_4555);
and UO_448 (O_448,N_4339,N_4853);
nand UO_449 (O_449,N_4107,N_4344);
nand UO_450 (O_450,N_4961,N_4208);
nor UO_451 (O_451,N_4772,N_4109);
and UO_452 (O_452,N_4765,N_4864);
and UO_453 (O_453,N_4831,N_4901);
nand UO_454 (O_454,N_4578,N_4956);
nor UO_455 (O_455,N_4668,N_4163);
nor UO_456 (O_456,N_4758,N_4481);
xor UO_457 (O_457,N_4937,N_4686);
nand UO_458 (O_458,N_4401,N_4545);
or UO_459 (O_459,N_4518,N_4807);
nand UO_460 (O_460,N_4229,N_4683);
or UO_461 (O_461,N_4337,N_4491);
and UO_462 (O_462,N_4138,N_4077);
nor UO_463 (O_463,N_4618,N_4500);
nor UO_464 (O_464,N_4386,N_4601);
or UO_465 (O_465,N_4013,N_4749);
nor UO_466 (O_466,N_4465,N_4024);
nand UO_467 (O_467,N_4181,N_4331);
nand UO_468 (O_468,N_4101,N_4002);
and UO_469 (O_469,N_4894,N_4479);
nand UO_470 (O_470,N_4867,N_4277);
or UO_471 (O_471,N_4267,N_4416);
nor UO_472 (O_472,N_4766,N_4536);
and UO_473 (O_473,N_4280,N_4044);
nor UO_474 (O_474,N_4436,N_4775);
nor UO_475 (O_475,N_4603,N_4189);
nor UO_476 (O_476,N_4391,N_4662);
or UO_477 (O_477,N_4909,N_4276);
nor UO_478 (O_478,N_4787,N_4529);
nor UO_479 (O_479,N_4689,N_4032);
nand UO_480 (O_480,N_4912,N_4755);
nand UO_481 (O_481,N_4153,N_4887);
or UO_482 (O_482,N_4198,N_4395);
and UO_483 (O_483,N_4986,N_4026);
or UO_484 (O_484,N_4622,N_4317);
nor UO_485 (O_485,N_4921,N_4452);
or UO_486 (O_486,N_4915,N_4808);
nand UO_487 (O_487,N_4430,N_4439);
nor UO_488 (O_488,N_4538,N_4885);
nor UO_489 (O_489,N_4751,N_4674);
or UO_490 (O_490,N_4313,N_4323);
and UO_491 (O_491,N_4964,N_4413);
nor UO_492 (O_492,N_4731,N_4148);
and UO_493 (O_493,N_4510,N_4347);
nor UO_494 (O_494,N_4753,N_4633);
nor UO_495 (O_495,N_4247,N_4274);
and UO_496 (O_496,N_4556,N_4147);
nor UO_497 (O_497,N_4225,N_4105);
or UO_498 (O_498,N_4034,N_4091);
nor UO_499 (O_499,N_4782,N_4540);
nand UO_500 (O_500,N_4908,N_4648);
or UO_501 (O_501,N_4116,N_4607);
or UO_502 (O_502,N_4364,N_4119);
nor UO_503 (O_503,N_4373,N_4352);
and UO_504 (O_504,N_4066,N_4392);
nand UO_505 (O_505,N_4565,N_4839);
and UO_506 (O_506,N_4221,N_4967);
nand UO_507 (O_507,N_4816,N_4693);
or UO_508 (O_508,N_4954,N_4021);
nand UO_509 (O_509,N_4165,N_4632);
nand UO_510 (O_510,N_4155,N_4453);
nor UO_511 (O_511,N_4634,N_4799);
nand UO_512 (O_512,N_4105,N_4069);
or UO_513 (O_513,N_4688,N_4390);
nand UO_514 (O_514,N_4071,N_4617);
nand UO_515 (O_515,N_4806,N_4850);
and UO_516 (O_516,N_4554,N_4297);
nand UO_517 (O_517,N_4925,N_4246);
or UO_518 (O_518,N_4748,N_4164);
nand UO_519 (O_519,N_4240,N_4060);
nor UO_520 (O_520,N_4660,N_4869);
nor UO_521 (O_521,N_4074,N_4660);
nand UO_522 (O_522,N_4853,N_4189);
nor UO_523 (O_523,N_4333,N_4673);
nor UO_524 (O_524,N_4403,N_4861);
or UO_525 (O_525,N_4743,N_4147);
or UO_526 (O_526,N_4657,N_4218);
and UO_527 (O_527,N_4711,N_4496);
nand UO_528 (O_528,N_4038,N_4750);
nand UO_529 (O_529,N_4213,N_4773);
nand UO_530 (O_530,N_4065,N_4359);
and UO_531 (O_531,N_4368,N_4474);
nand UO_532 (O_532,N_4426,N_4343);
or UO_533 (O_533,N_4411,N_4080);
nand UO_534 (O_534,N_4310,N_4940);
nor UO_535 (O_535,N_4010,N_4438);
nand UO_536 (O_536,N_4590,N_4388);
and UO_537 (O_537,N_4971,N_4114);
nor UO_538 (O_538,N_4115,N_4036);
and UO_539 (O_539,N_4943,N_4197);
nor UO_540 (O_540,N_4777,N_4298);
nor UO_541 (O_541,N_4233,N_4739);
nand UO_542 (O_542,N_4659,N_4711);
or UO_543 (O_543,N_4748,N_4889);
nor UO_544 (O_544,N_4324,N_4233);
and UO_545 (O_545,N_4183,N_4146);
or UO_546 (O_546,N_4492,N_4153);
and UO_547 (O_547,N_4980,N_4495);
and UO_548 (O_548,N_4658,N_4708);
nand UO_549 (O_549,N_4020,N_4432);
or UO_550 (O_550,N_4140,N_4420);
and UO_551 (O_551,N_4132,N_4620);
xor UO_552 (O_552,N_4408,N_4765);
nand UO_553 (O_553,N_4521,N_4824);
and UO_554 (O_554,N_4078,N_4651);
nand UO_555 (O_555,N_4093,N_4443);
nand UO_556 (O_556,N_4473,N_4325);
nor UO_557 (O_557,N_4458,N_4830);
or UO_558 (O_558,N_4306,N_4377);
nand UO_559 (O_559,N_4379,N_4183);
or UO_560 (O_560,N_4125,N_4826);
or UO_561 (O_561,N_4011,N_4710);
and UO_562 (O_562,N_4859,N_4645);
nand UO_563 (O_563,N_4648,N_4220);
xor UO_564 (O_564,N_4213,N_4171);
nor UO_565 (O_565,N_4007,N_4195);
xor UO_566 (O_566,N_4966,N_4643);
nand UO_567 (O_567,N_4915,N_4057);
nand UO_568 (O_568,N_4190,N_4316);
nand UO_569 (O_569,N_4554,N_4272);
nand UO_570 (O_570,N_4266,N_4072);
or UO_571 (O_571,N_4325,N_4163);
nor UO_572 (O_572,N_4296,N_4743);
and UO_573 (O_573,N_4819,N_4461);
or UO_574 (O_574,N_4490,N_4249);
nor UO_575 (O_575,N_4550,N_4893);
or UO_576 (O_576,N_4109,N_4686);
or UO_577 (O_577,N_4990,N_4105);
or UO_578 (O_578,N_4063,N_4462);
and UO_579 (O_579,N_4315,N_4747);
nor UO_580 (O_580,N_4227,N_4982);
nand UO_581 (O_581,N_4467,N_4055);
nand UO_582 (O_582,N_4314,N_4480);
and UO_583 (O_583,N_4027,N_4490);
nor UO_584 (O_584,N_4158,N_4717);
nor UO_585 (O_585,N_4428,N_4529);
nand UO_586 (O_586,N_4604,N_4887);
nand UO_587 (O_587,N_4099,N_4987);
nor UO_588 (O_588,N_4746,N_4889);
and UO_589 (O_589,N_4183,N_4948);
and UO_590 (O_590,N_4174,N_4681);
or UO_591 (O_591,N_4222,N_4627);
or UO_592 (O_592,N_4624,N_4061);
or UO_593 (O_593,N_4261,N_4550);
nor UO_594 (O_594,N_4234,N_4198);
or UO_595 (O_595,N_4502,N_4358);
and UO_596 (O_596,N_4188,N_4310);
nor UO_597 (O_597,N_4260,N_4190);
or UO_598 (O_598,N_4561,N_4840);
or UO_599 (O_599,N_4054,N_4165);
and UO_600 (O_600,N_4761,N_4012);
nor UO_601 (O_601,N_4939,N_4043);
or UO_602 (O_602,N_4600,N_4006);
xnor UO_603 (O_603,N_4729,N_4588);
or UO_604 (O_604,N_4873,N_4298);
nor UO_605 (O_605,N_4037,N_4780);
nand UO_606 (O_606,N_4805,N_4758);
nand UO_607 (O_607,N_4783,N_4634);
nand UO_608 (O_608,N_4012,N_4791);
or UO_609 (O_609,N_4816,N_4613);
or UO_610 (O_610,N_4414,N_4320);
nand UO_611 (O_611,N_4315,N_4647);
or UO_612 (O_612,N_4798,N_4639);
and UO_613 (O_613,N_4592,N_4731);
or UO_614 (O_614,N_4838,N_4666);
or UO_615 (O_615,N_4754,N_4611);
nor UO_616 (O_616,N_4144,N_4168);
nor UO_617 (O_617,N_4987,N_4507);
and UO_618 (O_618,N_4927,N_4237);
nand UO_619 (O_619,N_4853,N_4683);
and UO_620 (O_620,N_4454,N_4748);
or UO_621 (O_621,N_4768,N_4796);
or UO_622 (O_622,N_4000,N_4539);
and UO_623 (O_623,N_4211,N_4489);
nor UO_624 (O_624,N_4137,N_4663);
and UO_625 (O_625,N_4102,N_4684);
nand UO_626 (O_626,N_4523,N_4627);
and UO_627 (O_627,N_4652,N_4152);
nor UO_628 (O_628,N_4144,N_4209);
nand UO_629 (O_629,N_4826,N_4344);
nand UO_630 (O_630,N_4421,N_4410);
and UO_631 (O_631,N_4826,N_4804);
nor UO_632 (O_632,N_4697,N_4919);
or UO_633 (O_633,N_4926,N_4481);
and UO_634 (O_634,N_4970,N_4053);
nor UO_635 (O_635,N_4959,N_4909);
and UO_636 (O_636,N_4766,N_4112);
nor UO_637 (O_637,N_4230,N_4792);
nand UO_638 (O_638,N_4116,N_4032);
and UO_639 (O_639,N_4732,N_4251);
nor UO_640 (O_640,N_4751,N_4011);
nand UO_641 (O_641,N_4881,N_4333);
and UO_642 (O_642,N_4645,N_4224);
and UO_643 (O_643,N_4978,N_4029);
nand UO_644 (O_644,N_4712,N_4332);
nor UO_645 (O_645,N_4586,N_4974);
nor UO_646 (O_646,N_4137,N_4182);
nand UO_647 (O_647,N_4205,N_4867);
or UO_648 (O_648,N_4098,N_4961);
nor UO_649 (O_649,N_4583,N_4436);
nor UO_650 (O_650,N_4610,N_4553);
and UO_651 (O_651,N_4766,N_4826);
and UO_652 (O_652,N_4904,N_4065);
or UO_653 (O_653,N_4520,N_4366);
or UO_654 (O_654,N_4230,N_4531);
nor UO_655 (O_655,N_4659,N_4744);
nor UO_656 (O_656,N_4469,N_4111);
nor UO_657 (O_657,N_4208,N_4354);
or UO_658 (O_658,N_4594,N_4161);
nor UO_659 (O_659,N_4491,N_4311);
or UO_660 (O_660,N_4233,N_4490);
xnor UO_661 (O_661,N_4580,N_4249);
and UO_662 (O_662,N_4200,N_4489);
nand UO_663 (O_663,N_4483,N_4322);
and UO_664 (O_664,N_4966,N_4138);
and UO_665 (O_665,N_4472,N_4637);
nor UO_666 (O_666,N_4810,N_4056);
and UO_667 (O_667,N_4638,N_4386);
nor UO_668 (O_668,N_4579,N_4188);
or UO_669 (O_669,N_4533,N_4854);
xnor UO_670 (O_670,N_4444,N_4208);
or UO_671 (O_671,N_4322,N_4458);
and UO_672 (O_672,N_4485,N_4478);
or UO_673 (O_673,N_4175,N_4897);
and UO_674 (O_674,N_4916,N_4976);
nand UO_675 (O_675,N_4385,N_4603);
or UO_676 (O_676,N_4677,N_4073);
or UO_677 (O_677,N_4352,N_4534);
xor UO_678 (O_678,N_4136,N_4529);
nor UO_679 (O_679,N_4664,N_4105);
or UO_680 (O_680,N_4273,N_4820);
and UO_681 (O_681,N_4015,N_4344);
and UO_682 (O_682,N_4829,N_4079);
or UO_683 (O_683,N_4460,N_4912);
nand UO_684 (O_684,N_4983,N_4716);
and UO_685 (O_685,N_4559,N_4416);
or UO_686 (O_686,N_4079,N_4414);
nor UO_687 (O_687,N_4976,N_4415);
and UO_688 (O_688,N_4787,N_4595);
and UO_689 (O_689,N_4609,N_4848);
and UO_690 (O_690,N_4998,N_4130);
or UO_691 (O_691,N_4816,N_4027);
nand UO_692 (O_692,N_4740,N_4799);
nand UO_693 (O_693,N_4309,N_4914);
nand UO_694 (O_694,N_4096,N_4736);
nand UO_695 (O_695,N_4990,N_4236);
xor UO_696 (O_696,N_4387,N_4859);
nand UO_697 (O_697,N_4009,N_4189);
and UO_698 (O_698,N_4486,N_4973);
nand UO_699 (O_699,N_4892,N_4917);
nor UO_700 (O_700,N_4749,N_4218);
and UO_701 (O_701,N_4256,N_4050);
or UO_702 (O_702,N_4272,N_4371);
or UO_703 (O_703,N_4731,N_4187);
and UO_704 (O_704,N_4254,N_4603);
or UO_705 (O_705,N_4690,N_4907);
and UO_706 (O_706,N_4459,N_4081);
nor UO_707 (O_707,N_4408,N_4785);
or UO_708 (O_708,N_4663,N_4198);
nand UO_709 (O_709,N_4862,N_4543);
nor UO_710 (O_710,N_4892,N_4234);
and UO_711 (O_711,N_4793,N_4575);
nand UO_712 (O_712,N_4213,N_4499);
nor UO_713 (O_713,N_4054,N_4161);
nor UO_714 (O_714,N_4314,N_4441);
nor UO_715 (O_715,N_4804,N_4687);
and UO_716 (O_716,N_4182,N_4586);
and UO_717 (O_717,N_4633,N_4270);
nand UO_718 (O_718,N_4739,N_4912);
or UO_719 (O_719,N_4299,N_4284);
or UO_720 (O_720,N_4075,N_4771);
or UO_721 (O_721,N_4907,N_4384);
nand UO_722 (O_722,N_4530,N_4322);
and UO_723 (O_723,N_4024,N_4291);
or UO_724 (O_724,N_4085,N_4462);
or UO_725 (O_725,N_4847,N_4122);
nor UO_726 (O_726,N_4810,N_4693);
nand UO_727 (O_727,N_4146,N_4376);
nand UO_728 (O_728,N_4106,N_4105);
nand UO_729 (O_729,N_4855,N_4439);
nand UO_730 (O_730,N_4590,N_4841);
nand UO_731 (O_731,N_4554,N_4844);
nand UO_732 (O_732,N_4891,N_4045);
and UO_733 (O_733,N_4227,N_4818);
nor UO_734 (O_734,N_4484,N_4592);
and UO_735 (O_735,N_4338,N_4355);
and UO_736 (O_736,N_4782,N_4700);
or UO_737 (O_737,N_4701,N_4430);
or UO_738 (O_738,N_4603,N_4216);
and UO_739 (O_739,N_4785,N_4559);
or UO_740 (O_740,N_4976,N_4934);
nor UO_741 (O_741,N_4134,N_4113);
or UO_742 (O_742,N_4793,N_4445);
nand UO_743 (O_743,N_4100,N_4904);
nand UO_744 (O_744,N_4377,N_4249);
or UO_745 (O_745,N_4630,N_4303);
or UO_746 (O_746,N_4277,N_4574);
nor UO_747 (O_747,N_4161,N_4625);
or UO_748 (O_748,N_4073,N_4623);
or UO_749 (O_749,N_4882,N_4627);
and UO_750 (O_750,N_4470,N_4798);
nor UO_751 (O_751,N_4951,N_4744);
nor UO_752 (O_752,N_4339,N_4302);
nor UO_753 (O_753,N_4342,N_4049);
xnor UO_754 (O_754,N_4412,N_4528);
nor UO_755 (O_755,N_4748,N_4519);
or UO_756 (O_756,N_4279,N_4017);
nand UO_757 (O_757,N_4733,N_4923);
nor UO_758 (O_758,N_4474,N_4838);
nand UO_759 (O_759,N_4499,N_4555);
nor UO_760 (O_760,N_4178,N_4344);
xor UO_761 (O_761,N_4353,N_4080);
nor UO_762 (O_762,N_4071,N_4015);
nand UO_763 (O_763,N_4198,N_4154);
or UO_764 (O_764,N_4383,N_4752);
nand UO_765 (O_765,N_4756,N_4383);
nand UO_766 (O_766,N_4051,N_4935);
nand UO_767 (O_767,N_4852,N_4780);
and UO_768 (O_768,N_4642,N_4331);
nand UO_769 (O_769,N_4651,N_4156);
or UO_770 (O_770,N_4486,N_4925);
or UO_771 (O_771,N_4363,N_4785);
nand UO_772 (O_772,N_4693,N_4145);
nor UO_773 (O_773,N_4787,N_4471);
or UO_774 (O_774,N_4692,N_4413);
or UO_775 (O_775,N_4811,N_4034);
and UO_776 (O_776,N_4547,N_4676);
or UO_777 (O_777,N_4175,N_4253);
nor UO_778 (O_778,N_4475,N_4582);
nand UO_779 (O_779,N_4938,N_4622);
nor UO_780 (O_780,N_4664,N_4759);
nand UO_781 (O_781,N_4891,N_4572);
nand UO_782 (O_782,N_4442,N_4978);
nand UO_783 (O_783,N_4079,N_4288);
and UO_784 (O_784,N_4836,N_4195);
nand UO_785 (O_785,N_4114,N_4157);
nand UO_786 (O_786,N_4854,N_4589);
and UO_787 (O_787,N_4325,N_4269);
nor UO_788 (O_788,N_4375,N_4843);
nor UO_789 (O_789,N_4480,N_4630);
nand UO_790 (O_790,N_4926,N_4781);
nand UO_791 (O_791,N_4211,N_4017);
nor UO_792 (O_792,N_4948,N_4395);
nor UO_793 (O_793,N_4508,N_4708);
or UO_794 (O_794,N_4795,N_4681);
and UO_795 (O_795,N_4372,N_4123);
and UO_796 (O_796,N_4082,N_4234);
and UO_797 (O_797,N_4888,N_4436);
nand UO_798 (O_798,N_4070,N_4972);
nand UO_799 (O_799,N_4967,N_4314);
nor UO_800 (O_800,N_4350,N_4558);
or UO_801 (O_801,N_4904,N_4733);
nor UO_802 (O_802,N_4155,N_4803);
nor UO_803 (O_803,N_4766,N_4829);
nand UO_804 (O_804,N_4203,N_4381);
nand UO_805 (O_805,N_4097,N_4993);
nand UO_806 (O_806,N_4823,N_4036);
nand UO_807 (O_807,N_4272,N_4527);
xor UO_808 (O_808,N_4973,N_4678);
nand UO_809 (O_809,N_4070,N_4420);
and UO_810 (O_810,N_4649,N_4024);
xnor UO_811 (O_811,N_4666,N_4606);
nor UO_812 (O_812,N_4684,N_4483);
and UO_813 (O_813,N_4360,N_4389);
and UO_814 (O_814,N_4957,N_4163);
or UO_815 (O_815,N_4448,N_4617);
or UO_816 (O_816,N_4331,N_4509);
and UO_817 (O_817,N_4435,N_4836);
and UO_818 (O_818,N_4164,N_4281);
xor UO_819 (O_819,N_4612,N_4322);
and UO_820 (O_820,N_4225,N_4765);
nand UO_821 (O_821,N_4416,N_4849);
nor UO_822 (O_822,N_4201,N_4450);
nand UO_823 (O_823,N_4614,N_4744);
nand UO_824 (O_824,N_4926,N_4393);
nand UO_825 (O_825,N_4444,N_4450);
nand UO_826 (O_826,N_4536,N_4656);
nand UO_827 (O_827,N_4215,N_4234);
or UO_828 (O_828,N_4015,N_4408);
nand UO_829 (O_829,N_4608,N_4899);
nor UO_830 (O_830,N_4345,N_4791);
nor UO_831 (O_831,N_4791,N_4578);
nand UO_832 (O_832,N_4432,N_4530);
nor UO_833 (O_833,N_4578,N_4912);
or UO_834 (O_834,N_4929,N_4962);
or UO_835 (O_835,N_4789,N_4189);
nand UO_836 (O_836,N_4565,N_4577);
nand UO_837 (O_837,N_4640,N_4437);
and UO_838 (O_838,N_4874,N_4833);
nand UO_839 (O_839,N_4775,N_4717);
nand UO_840 (O_840,N_4988,N_4238);
or UO_841 (O_841,N_4348,N_4180);
nor UO_842 (O_842,N_4139,N_4236);
nor UO_843 (O_843,N_4107,N_4833);
or UO_844 (O_844,N_4553,N_4934);
or UO_845 (O_845,N_4312,N_4975);
nor UO_846 (O_846,N_4072,N_4808);
nand UO_847 (O_847,N_4346,N_4585);
nand UO_848 (O_848,N_4411,N_4961);
nand UO_849 (O_849,N_4164,N_4396);
nand UO_850 (O_850,N_4704,N_4933);
and UO_851 (O_851,N_4400,N_4200);
or UO_852 (O_852,N_4411,N_4021);
and UO_853 (O_853,N_4423,N_4003);
nand UO_854 (O_854,N_4643,N_4926);
and UO_855 (O_855,N_4472,N_4960);
nor UO_856 (O_856,N_4657,N_4174);
and UO_857 (O_857,N_4183,N_4171);
nand UO_858 (O_858,N_4500,N_4643);
nand UO_859 (O_859,N_4220,N_4479);
and UO_860 (O_860,N_4828,N_4764);
nand UO_861 (O_861,N_4113,N_4548);
nand UO_862 (O_862,N_4732,N_4570);
nand UO_863 (O_863,N_4913,N_4472);
or UO_864 (O_864,N_4567,N_4118);
or UO_865 (O_865,N_4475,N_4022);
nor UO_866 (O_866,N_4246,N_4501);
and UO_867 (O_867,N_4232,N_4971);
nor UO_868 (O_868,N_4151,N_4899);
or UO_869 (O_869,N_4883,N_4346);
nor UO_870 (O_870,N_4241,N_4856);
nor UO_871 (O_871,N_4956,N_4007);
nor UO_872 (O_872,N_4780,N_4552);
or UO_873 (O_873,N_4221,N_4243);
nor UO_874 (O_874,N_4337,N_4371);
and UO_875 (O_875,N_4430,N_4844);
or UO_876 (O_876,N_4050,N_4187);
nand UO_877 (O_877,N_4976,N_4876);
and UO_878 (O_878,N_4244,N_4129);
and UO_879 (O_879,N_4932,N_4057);
or UO_880 (O_880,N_4966,N_4721);
nor UO_881 (O_881,N_4541,N_4627);
and UO_882 (O_882,N_4921,N_4735);
and UO_883 (O_883,N_4749,N_4144);
nor UO_884 (O_884,N_4373,N_4241);
nor UO_885 (O_885,N_4834,N_4628);
nand UO_886 (O_886,N_4025,N_4376);
nor UO_887 (O_887,N_4851,N_4419);
nand UO_888 (O_888,N_4041,N_4937);
nand UO_889 (O_889,N_4670,N_4833);
and UO_890 (O_890,N_4467,N_4286);
nand UO_891 (O_891,N_4319,N_4787);
and UO_892 (O_892,N_4850,N_4439);
or UO_893 (O_893,N_4671,N_4325);
and UO_894 (O_894,N_4589,N_4739);
or UO_895 (O_895,N_4455,N_4954);
or UO_896 (O_896,N_4132,N_4976);
and UO_897 (O_897,N_4881,N_4204);
nand UO_898 (O_898,N_4814,N_4596);
nand UO_899 (O_899,N_4659,N_4884);
and UO_900 (O_900,N_4708,N_4551);
or UO_901 (O_901,N_4167,N_4074);
nor UO_902 (O_902,N_4075,N_4001);
nor UO_903 (O_903,N_4004,N_4563);
nand UO_904 (O_904,N_4018,N_4938);
and UO_905 (O_905,N_4566,N_4889);
and UO_906 (O_906,N_4232,N_4977);
and UO_907 (O_907,N_4039,N_4803);
or UO_908 (O_908,N_4594,N_4505);
nor UO_909 (O_909,N_4898,N_4590);
nand UO_910 (O_910,N_4092,N_4404);
xor UO_911 (O_911,N_4103,N_4913);
nand UO_912 (O_912,N_4900,N_4825);
nor UO_913 (O_913,N_4315,N_4891);
and UO_914 (O_914,N_4616,N_4701);
or UO_915 (O_915,N_4820,N_4928);
nand UO_916 (O_916,N_4814,N_4380);
and UO_917 (O_917,N_4651,N_4856);
or UO_918 (O_918,N_4305,N_4499);
or UO_919 (O_919,N_4444,N_4735);
nand UO_920 (O_920,N_4443,N_4192);
or UO_921 (O_921,N_4981,N_4396);
nor UO_922 (O_922,N_4171,N_4426);
nand UO_923 (O_923,N_4091,N_4139);
and UO_924 (O_924,N_4761,N_4189);
and UO_925 (O_925,N_4787,N_4260);
nor UO_926 (O_926,N_4082,N_4459);
or UO_927 (O_927,N_4003,N_4228);
nand UO_928 (O_928,N_4575,N_4934);
nand UO_929 (O_929,N_4628,N_4683);
nand UO_930 (O_930,N_4233,N_4754);
nor UO_931 (O_931,N_4373,N_4688);
and UO_932 (O_932,N_4060,N_4974);
xnor UO_933 (O_933,N_4817,N_4776);
or UO_934 (O_934,N_4008,N_4494);
nor UO_935 (O_935,N_4413,N_4211);
nand UO_936 (O_936,N_4203,N_4901);
nand UO_937 (O_937,N_4476,N_4719);
nand UO_938 (O_938,N_4833,N_4376);
nor UO_939 (O_939,N_4451,N_4241);
nand UO_940 (O_940,N_4834,N_4316);
and UO_941 (O_941,N_4274,N_4759);
or UO_942 (O_942,N_4528,N_4380);
nor UO_943 (O_943,N_4672,N_4846);
nor UO_944 (O_944,N_4922,N_4891);
or UO_945 (O_945,N_4551,N_4083);
nand UO_946 (O_946,N_4358,N_4145);
and UO_947 (O_947,N_4127,N_4248);
nand UO_948 (O_948,N_4159,N_4931);
or UO_949 (O_949,N_4616,N_4711);
nand UO_950 (O_950,N_4104,N_4799);
and UO_951 (O_951,N_4302,N_4780);
nor UO_952 (O_952,N_4062,N_4793);
and UO_953 (O_953,N_4585,N_4492);
nand UO_954 (O_954,N_4775,N_4420);
nor UO_955 (O_955,N_4350,N_4369);
nor UO_956 (O_956,N_4441,N_4109);
or UO_957 (O_957,N_4410,N_4850);
xor UO_958 (O_958,N_4448,N_4778);
or UO_959 (O_959,N_4623,N_4403);
nor UO_960 (O_960,N_4323,N_4907);
and UO_961 (O_961,N_4561,N_4537);
or UO_962 (O_962,N_4573,N_4864);
nand UO_963 (O_963,N_4182,N_4159);
nor UO_964 (O_964,N_4871,N_4035);
and UO_965 (O_965,N_4980,N_4124);
and UO_966 (O_966,N_4890,N_4524);
nor UO_967 (O_967,N_4728,N_4565);
nand UO_968 (O_968,N_4277,N_4528);
nor UO_969 (O_969,N_4908,N_4979);
xor UO_970 (O_970,N_4885,N_4406);
and UO_971 (O_971,N_4835,N_4967);
and UO_972 (O_972,N_4902,N_4380);
nor UO_973 (O_973,N_4727,N_4028);
and UO_974 (O_974,N_4339,N_4515);
or UO_975 (O_975,N_4709,N_4713);
and UO_976 (O_976,N_4580,N_4981);
nor UO_977 (O_977,N_4181,N_4293);
and UO_978 (O_978,N_4752,N_4433);
and UO_979 (O_979,N_4308,N_4113);
nor UO_980 (O_980,N_4238,N_4109);
nor UO_981 (O_981,N_4762,N_4613);
nand UO_982 (O_982,N_4670,N_4596);
and UO_983 (O_983,N_4722,N_4567);
or UO_984 (O_984,N_4017,N_4189);
nand UO_985 (O_985,N_4920,N_4793);
or UO_986 (O_986,N_4801,N_4917);
or UO_987 (O_987,N_4919,N_4096);
nand UO_988 (O_988,N_4499,N_4913);
xnor UO_989 (O_989,N_4105,N_4076);
and UO_990 (O_990,N_4192,N_4969);
xor UO_991 (O_991,N_4511,N_4127);
and UO_992 (O_992,N_4735,N_4514);
nor UO_993 (O_993,N_4420,N_4242);
nand UO_994 (O_994,N_4905,N_4684);
or UO_995 (O_995,N_4348,N_4067);
nor UO_996 (O_996,N_4483,N_4536);
nor UO_997 (O_997,N_4209,N_4381);
nand UO_998 (O_998,N_4094,N_4413);
or UO_999 (O_999,N_4252,N_4343);
endmodule