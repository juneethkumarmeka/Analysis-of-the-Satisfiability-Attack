module basic_1500_15000_2000_120_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_539,In_341);
xor U1 (N_1,In_878,In_491);
or U2 (N_2,In_1442,In_413);
nor U3 (N_3,In_1468,In_786);
nand U4 (N_4,In_1285,In_774);
and U5 (N_5,In_829,In_1276);
and U6 (N_6,In_1294,In_689);
xor U7 (N_7,In_1232,In_1281);
nor U8 (N_8,In_1224,In_452);
or U9 (N_9,In_486,In_1209);
xor U10 (N_10,In_783,In_143);
nor U11 (N_11,In_335,In_494);
or U12 (N_12,In_65,In_986);
nand U13 (N_13,In_831,In_771);
and U14 (N_14,In_227,In_408);
nor U15 (N_15,In_321,In_320);
or U16 (N_16,In_740,In_392);
nor U17 (N_17,In_344,In_924);
xnor U18 (N_18,In_850,In_205);
xor U19 (N_19,In_1101,In_1445);
nor U20 (N_20,In_197,In_456);
nand U21 (N_21,In_317,In_1356);
nand U22 (N_22,In_1251,In_93);
and U23 (N_23,In_378,In_985);
and U24 (N_24,In_1187,In_1018);
or U25 (N_25,In_241,In_707);
nor U26 (N_26,In_654,In_1078);
and U27 (N_27,In_1343,In_1299);
xnor U28 (N_28,In_1186,In_1047);
nand U29 (N_29,In_386,In_168);
and U30 (N_30,In_798,In_659);
nor U31 (N_31,In_1165,In_222);
nor U32 (N_32,In_379,In_834);
or U33 (N_33,In_1094,In_588);
xnor U34 (N_34,In_279,In_810);
or U35 (N_35,In_1042,In_1496);
xor U36 (N_36,In_1036,In_109);
xor U37 (N_37,In_474,In_789);
nor U38 (N_38,In_1336,In_936);
or U39 (N_39,In_807,In_116);
nand U40 (N_40,In_663,In_1338);
xnor U41 (N_41,In_285,In_504);
or U42 (N_42,In_1002,In_984);
xnor U43 (N_43,In_943,In_1210);
and U44 (N_44,In_395,In_1071);
nand U45 (N_45,In_409,In_202);
nand U46 (N_46,In_1172,In_356);
nand U47 (N_47,In_80,In_181);
nand U48 (N_48,In_447,In_1325);
and U49 (N_49,In_477,In_399);
xnor U50 (N_50,In_195,In_1481);
xnor U51 (N_51,In_1200,In_290);
and U52 (N_52,In_581,In_544);
nand U53 (N_53,In_1215,In_1463);
nand U54 (N_54,In_684,In_120);
and U55 (N_55,In_639,In_235);
nor U56 (N_56,In_180,In_1167);
xnor U57 (N_57,In_1374,In_1246);
nand U58 (N_58,In_1008,In_1168);
or U59 (N_59,In_348,In_609);
and U60 (N_60,In_1024,In_1271);
xnor U61 (N_61,In_1323,In_1064);
or U62 (N_62,In_816,In_621);
or U63 (N_63,In_246,In_644);
xnor U64 (N_64,In_294,In_459);
and U65 (N_65,In_1406,In_1128);
or U66 (N_66,In_1181,In_914);
nor U67 (N_67,In_1477,In_144);
xnor U68 (N_68,In_1196,In_94);
and U69 (N_69,In_211,In_510);
nand U70 (N_70,In_342,In_618);
xor U71 (N_71,In_1169,In_697);
nand U72 (N_72,In_425,In_763);
nor U73 (N_73,In_655,In_855);
nor U74 (N_74,In_1283,In_590);
nor U75 (N_75,In_377,In_999);
or U76 (N_76,In_90,In_809);
nor U77 (N_77,In_72,In_1194);
nand U78 (N_78,In_1301,In_137);
and U79 (N_79,In_687,In_1397);
and U80 (N_80,In_499,In_46);
and U81 (N_81,In_201,In_860);
nand U82 (N_82,In_801,In_1157);
and U83 (N_83,In_1160,In_20);
nor U84 (N_84,In_1471,In_1004);
and U85 (N_85,In_1459,In_1351);
or U86 (N_86,In_398,In_1487);
or U87 (N_87,In_592,In_1121);
nor U88 (N_88,In_1309,In_1377);
xor U89 (N_89,In_569,In_752);
xor U90 (N_90,In_135,In_1082);
or U91 (N_91,In_974,In_983);
nand U92 (N_92,In_226,In_1393);
nor U93 (N_93,In_558,In_1162);
and U94 (N_94,In_533,In_393);
and U95 (N_95,In_126,In_637);
or U96 (N_96,In_819,In_10);
xor U97 (N_97,In_1049,In_957);
nor U98 (N_98,In_1131,In_1013);
nor U99 (N_99,In_1120,In_263);
xor U100 (N_100,In_694,In_726);
and U101 (N_101,In_928,In_704);
nor U102 (N_102,In_11,In_402);
xnor U103 (N_103,In_1416,In_318);
or U104 (N_104,In_910,In_715);
and U105 (N_105,In_74,In_1006);
nor U106 (N_106,In_273,In_147);
xor U107 (N_107,In_1054,In_1300);
nor U108 (N_108,In_476,In_1478);
nand U109 (N_109,In_1414,In_1225);
nand U110 (N_110,In_207,In_63);
xor U111 (N_111,In_958,In_138);
and U112 (N_112,In_1352,In_1217);
nand U113 (N_113,In_1443,In_753);
nand U114 (N_114,In_362,In_417);
nand U115 (N_115,In_1365,In_1080);
nand U116 (N_116,In_708,In_1012);
nand U117 (N_117,In_1439,In_847);
nor U118 (N_118,In_475,In_259);
nor U119 (N_119,In_719,In_997);
and U120 (N_120,In_1129,In_555);
and U121 (N_121,In_1124,In_230);
and U122 (N_122,In_653,In_433);
nand U123 (N_123,In_822,In_306);
or U124 (N_124,In_372,In_365);
xnor U125 (N_125,In_779,In_9);
nor U126 (N_126,In_1424,In_160);
nand U127 (N_127,N_42,In_1432);
xnor U128 (N_128,In_1243,In_620);
nor U129 (N_129,In_665,In_307);
and U130 (N_130,N_100,In_849);
nor U131 (N_131,In_781,In_755);
or U132 (N_132,In_946,In_165);
nor U133 (N_133,In_623,In_815);
and U134 (N_134,N_121,N_120);
nor U135 (N_135,In_38,In_1378);
xor U136 (N_136,In_1206,In_612);
nor U137 (N_137,In_1482,In_1122);
or U138 (N_138,N_6,In_531);
or U139 (N_139,In_1237,In_1110);
xor U140 (N_140,In_337,In_778);
and U141 (N_141,In_1093,In_703);
nor U142 (N_142,In_336,In_1239);
or U143 (N_143,In_1041,N_122);
and U144 (N_144,In_125,In_71);
xnor U145 (N_145,In_1292,In_376);
or U146 (N_146,In_595,In_537);
or U147 (N_147,In_1428,In_1188);
or U148 (N_148,N_34,In_328);
nand U149 (N_149,N_106,In_1058);
nand U150 (N_150,In_1405,In_1372);
nor U151 (N_151,In_870,In_596);
or U152 (N_152,In_909,In_705);
and U153 (N_153,In_407,In_791);
or U154 (N_154,In_113,In_700);
or U155 (N_155,In_481,In_1211);
xor U156 (N_156,N_19,In_1025);
and U157 (N_157,In_680,In_131);
and U158 (N_158,In_613,In_671);
or U159 (N_159,In_625,In_1458);
nand U160 (N_160,In_1083,In_35);
nand U161 (N_161,In_45,In_280);
xnor U162 (N_162,In_296,In_370);
nor U163 (N_163,In_432,In_1052);
and U164 (N_164,In_1197,In_1460);
nand U165 (N_165,In_628,N_31);
nand U166 (N_166,In_1087,In_978);
or U167 (N_167,In_1256,In_39);
xnor U168 (N_168,In_701,In_992);
nor U169 (N_169,In_1112,In_495);
or U170 (N_170,In_820,In_769);
xor U171 (N_171,In_360,In_208);
nand U172 (N_172,In_213,In_553);
nand U173 (N_173,N_87,In_1180);
and U174 (N_174,In_964,In_519);
or U175 (N_175,In_940,In_567);
and U176 (N_176,In_1193,In_7);
nand U177 (N_177,In_502,In_1067);
xor U178 (N_178,In_584,In_954);
or U179 (N_179,In_119,In_237);
xnor U180 (N_180,N_79,In_445);
or U181 (N_181,In_411,In_1177);
and U182 (N_182,In_128,In_394);
nor U183 (N_183,N_63,In_721);
nor U184 (N_184,In_480,In_1044);
or U185 (N_185,In_1244,In_1408);
nand U186 (N_186,In_518,In_1248);
nand U187 (N_187,In_1274,In_1486);
nand U188 (N_188,In_384,In_134);
xnor U189 (N_189,In_151,In_146);
xor U190 (N_190,In_1231,In_286);
xnor U191 (N_191,In_367,In_728);
nor U192 (N_192,N_86,In_571);
or U193 (N_193,In_439,In_514);
or U194 (N_194,In_1390,In_839);
and U195 (N_195,In_1137,In_1003);
or U196 (N_196,In_686,In_124);
or U197 (N_197,In_1060,In_239);
xnor U198 (N_198,In_1347,In_450);
and U199 (N_199,In_513,In_496);
xor U200 (N_200,In_1056,In_303);
nor U201 (N_201,N_37,In_966);
and U202 (N_202,N_46,In_890);
nor U203 (N_203,In_267,In_354);
and U204 (N_204,In_617,In_1322);
and U205 (N_205,In_47,N_67);
or U206 (N_206,In_174,In_1100);
xor U207 (N_207,In_1389,In_437);
xnor U208 (N_208,N_12,In_908);
nor U209 (N_209,In_258,In_1423);
xnor U210 (N_210,In_599,In_1409);
or U211 (N_211,In_58,In_1297);
nor U212 (N_212,N_108,In_1119);
nand U213 (N_213,In_111,In_552);
nand U214 (N_214,In_123,In_1005);
nand U215 (N_215,In_685,In_973);
xnor U216 (N_216,In_879,In_1220);
and U217 (N_217,In_852,In_866);
nand U218 (N_218,In_380,In_811);
nand U219 (N_219,In_1203,In_1022);
xor U220 (N_220,N_33,In_383);
or U221 (N_221,In_189,In_436);
xor U222 (N_222,In_785,In_359);
or U223 (N_223,In_915,In_1250);
nor U224 (N_224,N_92,In_875);
xnor U225 (N_225,In_1306,In_42);
nand U226 (N_226,In_522,In_219);
xor U227 (N_227,In_920,In_1035);
xnor U228 (N_228,N_84,In_2);
nor U229 (N_229,In_81,In_698);
nand U230 (N_230,N_98,In_534);
or U231 (N_231,In_214,In_892);
or U232 (N_232,In_767,In_1046);
nand U233 (N_233,In_1163,In_470);
and U234 (N_234,In_720,In_300);
xor U235 (N_235,In_509,In_526);
nor U236 (N_236,N_75,In_632);
nand U237 (N_237,N_32,N_65);
and U238 (N_238,In_465,In_883);
or U239 (N_239,In_594,N_80);
xor U240 (N_240,In_1411,In_68);
nor U241 (N_241,In_1114,In_21);
nor U242 (N_242,In_1033,N_35);
and U243 (N_243,In_1303,In_742);
nand U244 (N_244,N_52,In_672);
nor U245 (N_245,In_517,In_1434);
nand U246 (N_246,In_563,N_107);
nor U247 (N_247,In_265,In_345);
or U248 (N_248,In_570,In_1464);
xnor U249 (N_249,N_113,In_930);
or U250 (N_250,In_1291,In_787);
nand U251 (N_251,N_184,N_209);
or U252 (N_252,In_1495,In_1);
xnor U253 (N_253,In_813,N_149);
and U254 (N_254,In_177,In_56);
xnor U255 (N_255,In_224,N_85);
and U256 (N_256,N_226,In_1295);
and U257 (N_257,In_505,In_492);
and U258 (N_258,In_1339,N_193);
and U259 (N_259,In_926,In_746);
nand U260 (N_260,In_57,In_1407);
nor U261 (N_261,In_287,N_102);
xor U262 (N_262,In_876,In_466);
xnor U263 (N_263,In_1360,In_955);
nor U264 (N_264,In_261,N_127);
nand U265 (N_265,N_110,N_1);
nand U266 (N_266,In_405,In_77);
xnor U267 (N_267,In_190,In_770);
and U268 (N_268,In_754,In_1312);
or U269 (N_269,N_41,In_833);
xor U270 (N_270,In_311,N_214);
nand U271 (N_271,In_414,In_489);
nand U272 (N_272,In_1099,In_765);
xor U273 (N_273,In_289,In_4);
and U274 (N_274,In_25,In_1258);
and U275 (N_275,In_1453,In_350);
nor U276 (N_276,N_233,N_73);
nor U277 (N_277,In_1192,In_22);
nor U278 (N_278,N_70,In_1133);
nand U279 (N_279,N_146,In_757);
nor U280 (N_280,In_1418,N_195);
xnor U281 (N_281,In_727,In_699);
and U282 (N_282,In_212,In_196);
nor U283 (N_283,In_650,N_229);
nand U284 (N_284,N_99,In_1331);
nand U285 (N_285,In_153,In_149);
nand U286 (N_286,In_54,In_387);
nor U287 (N_287,In_52,In_87);
nand U288 (N_288,In_861,In_369);
xor U289 (N_289,In_1394,In_987);
xor U290 (N_290,In_1402,In_817);
xor U291 (N_291,In_1334,In_1324);
nand U292 (N_292,N_185,In_1214);
nor U293 (N_293,In_1433,In_607);
xor U294 (N_294,N_24,In_739);
and U295 (N_295,In_1342,In_1465);
nand U296 (N_296,In_347,N_118);
and U297 (N_297,In_479,In_430);
xor U298 (N_298,In_1399,N_216);
or U299 (N_299,In_1249,In_1176);
or U300 (N_300,In_1233,In_1227);
or U301 (N_301,In_990,In_679);
xnor U302 (N_302,In_150,In_1391);
nand U303 (N_303,N_167,In_269);
or U304 (N_304,In_640,In_423);
and U305 (N_305,In_1102,N_145);
nor U306 (N_306,In_83,In_431);
nor U307 (N_307,In_1494,In_389);
or U308 (N_308,In_1095,In_587);
nand U309 (N_309,N_39,N_129);
nor U310 (N_310,In_877,In_709);
xnor U311 (N_311,In_349,In_493);
and U312 (N_312,In_175,In_23);
nand U313 (N_313,In_506,In_1057);
nor U314 (N_314,In_961,In_1375);
and U315 (N_315,In_8,In_1107);
nand U316 (N_316,In_1272,N_128);
or U317 (N_317,In_925,In_472);
or U318 (N_318,In_1440,N_132);
and U319 (N_319,N_156,In_541);
nor U320 (N_320,In_33,In_251);
and U321 (N_321,In_451,In_988);
or U322 (N_322,In_1387,In_1497);
nand U323 (N_323,N_4,In_716);
or U324 (N_324,In_1084,In_215);
nor U325 (N_325,In_963,In_1261);
nand U326 (N_326,In_714,In_1255);
nor U327 (N_327,In_48,In_950);
or U328 (N_328,In_304,In_556);
and U329 (N_329,In_803,N_235);
nand U330 (N_330,In_645,In_1175);
and U331 (N_331,In_164,N_135);
and U332 (N_332,In_1259,In_758);
xnor U333 (N_333,In_1470,In_1127);
nand U334 (N_334,In_911,In_1308);
and U335 (N_335,In_965,In_1048);
and U336 (N_336,In_136,In_1016);
xnor U337 (N_337,In_217,In_1316);
xor U338 (N_338,In_1030,In_322);
and U339 (N_339,In_1370,In_947);
and U340 (N_340,In_1436,In_96);
nor U341 (N_341,N_228,N_213);
xnor U342 (N_342,In_1412,In_1069);
nor U343 (N_343,In_808,In_976);
nor U344 (N_344,In_315,In_871);
xnor U345 (N_345,In_406,In_1065);
xor U346 (N_346,In_1269,N_54);
or U347 (N_347,In_1268,In_667);
nand U348 (N_348,N_143,In_887);
or U349 (N_349,In_585,N_14);
or U350 (N_350,N_222,N_186);
xor U351 (N_351,In_636,In_1135);
nand U352 (N_352,In_604,In_568);
and U353 (N_353,N_27,In_1469);
nor U354 (N_354,N_28,In_18);
nor U355 (N_355,In_457,In_788);
xor U356 (N_356,In_615,In_163);
and U357 (N_357,In_82,In_827);
and U358 (N_358,In_385,N_243);
or U359 (N_359,In_99,In_741);
and U360 (N_360,N_104,In_1426);
nor U361 (N_361,In_253,N_240);
or U362 (N_362,N_111,In_1179);
or U363 (N_363,In_242,In_856);
nor U364 (N_364,In_1247,In_1457);
xnor U365 (N_365,In_666,In_841);
nor U366 (N_366,In_766,In_1147);
nand U367 (N_367,In_1310,In_40);
nand U368 (N_368,In_1159,In_589);
xnor U369 (N_369,In_1350,In_900);
nand U370 (N_370,N_151,In_1381);
or U371 (N_371,In_62,In_916);
nand U372 (N_372,In_648,In_873);
xor U373 (N_373,In_591,N_133);
nand U374 (N_374,In_371,In_102);
nor U375 (N_375,In_1222,In_882);
nand U376 (N_376,In_1346,In_1320);
and U377 (N_377,In_793,N_322);
nand U378 (N_378,N_257,In_762);
nand U379 (N_379,In_1241,In_790);
and U380 (N_380,In_1189,In_1104);
and U381 (N_381,N_13,In_50);
and U382 (N_382,In_1483,In_837);
nor U383 (N_383,In_464,In_772);
nor U384 (N_384,N_159,N_55);
xnor U385 (N_385,In_863,In_927);
and U386 (N_386,In_935,In_1236);
nor U387 (N_387,In_660,In_1435);
and U388 (N_388,In_843,In_262);
xor U389 (N_389,In_220,In_1021);
and U390 (N_390,In_1447,In_1344);
xnor U391 (N_391,N_155,N_335);
xor U392 (N_392,In_980,In_1371);
and U393 (N_393,In_37,In_743);
or U394 (N_394,N_292,In_130);
nor U395 (N_395,In_503,In_283);
xor U396 (N_396,In_748,In_874);
and U397 (N_397,N_194,In_101);
xnor U398 (N_398,In_904,In_1205);
nand U399 (N_399,In_784,In_108);
nor U400 (N_400,In_1155,In_1116);
nor U401 (N_401,N_350,N_196);
nor U402 (N_402,N_191,N_334);
nand U403 (N_403,In_204,N_21);
and U404 (N_404,In_917,N_90);
nor U405 (N_405,In_117,In_1386);
xnor U406 (N_406,N_97,N_299);
nand U407 (N_407,In_989,N_50);
xor U408 (N_408,In_188,In_918);
or U409 (N_409,In_92,In_112);
nand U410 (N_410,In_1280,In_845);
nand U411 (N_411,In_234,N_227);
nand U412 (N_412,In_396,In_546);
or U413 (N_413,In_551,In_566);
nand U414 (N_414,In_934,N_252);
nor U415 (N_415,N_74,N_183);
or U416 (N_416,In_141,In_1484);
and U417 (N_417,In_603,N_269);
or U418 (N_418,In_338,In_418);
or U419 (N_419,In_352,In_610);
and U420 (N_420,In_24,In_1430);
or U421 (N_421,In_1466,In_233);
or U422 (N_422,In_806,N_288);
or U423 (N_423,In_1072,In_184);
or U424 (N_424,In_962,In_1051);
or U425 (N_425,In_314,N_273);
xnor U426 (N_426,N_175,N_215);
xor U427 (N_427,In_231,N_370);
and U428 (N_428,In_1368,In_601);
or U429 (N_429,N_224,In_664);
or U430 (N_430,In_1345,N_336);
and U431 (N_431,In_1395,In_429);
xnor U432 (N_432,N_357,N_48);
nor U433 (N_433,N_312,In_435);
nor U434 (N_434,In_19,In_718);
nor U435 (N_435,In_1260,In_85);
and U436 (N_436,N_307,In_404);
xnor U437 (N_437,N_189,N_302);
and U438 (N_438,In_1396,In_14);
nand U439 (N_439,N_172,In_434);
nand U440 (N_440,In_291,In_1096);
nor U441 (N_441,In_886,In_331);
xnor U442 (N_442,In_1014,In_674);
nand U443 (N_443,In_257,In_170);
xnor U444 (N_444,In_724,N_140);
xor U445 (N_445,N_241,N_300);
and U446 (N_446,In_832,In_1449);
nand U447 (N_447,In_562,In_1366);
nor U448 (N_448,In_5,In_182);
and U449 (N_449,N_303,In_1098);
nor U450 (N_450,In_670,In_1050);
nor U451 (N_451,In_525,In_661);
xor U452 (N_452,In_629,In_366);
xor U453 (N_453,In_1111,In_775);
or U454 (N_454,In_1242,N_279);
and U455 (N_455,In_1229,In_516);
xnor U456 (N_456,In_865,In_899);
and U457 (N_457,In_884,In_630);
nand U458 (N_458,In_582,N_115);
nand U459 (N_459,In_107,In_897);
nor U460 (N_460,In_545,N_147);
or U461 (N_461,In_717,In_3);
xnor U462 (N_462,In_326,In_268);
xnor U463 (N_463,N_321,In_1473);
xnor U464 (N_464,N_266,In_1109);
nor U465 (N_465,In_487,In_1431);
nor U466 (N_466,In_478,In_862);
or U467 (N_467,N_3,In_327);
and U468 (N_468,In_75,N_8);
xor U469 (N_469,In_458,N_276);
or U470 (N_470,In_240,In_919);
and U471 (N_471,In_30,In_658);
xor U472 (N_472,In_309,In_635);
nand U473 (N_473,In_1328,N_210);
nand U474 (N_474,N_255,In_293);
nand U475 (N_475,N_198,In_390);
nand U476 (N_476,N_53,In_608);
xor U477 (N_477,N_38,In_633);
and U478 (N_478,In_768,In_794);
xnor U479 (N_479,In_1141,N_271);
or U480 (N_480,N_373,In_1448);
xnor U481 (N_481,In_1373,In_932);
or U482 (N_482,N_242,N_187);
nor U483 (N_483,In_64,In_455);
nor U484 (N_484,In_1178,In_854);
nor U485 (N_485,N_264,In_1149);
nor U486 (N_486,In_1208,N_165);
xnor U487 (N_487,In_764,N_153);
and U488 (N_488,In_277,N_188);
xor U489 (N_489,In_804,N_262);
or U490 (N_490,N_328,N_5);
xnor U491 (N_491,In_521,N_161);
and U492 (N_492,N_283,In_363);
nor U493 (N_493,N_23,In_316);
or U494 (N_494,In_975,N_359);
nand U495 (N_495,In_1066,N_76);
or U496 (N_496,In_167,In_1139);
and U497 (N_497,In_1425,In_462);
and U498 (N_498,In_548,In_1314);
nand U499 (N_499,In_577,In_729);
xnor U500 (N_500,N_88,In_51);
nor U501 (N_501,In_70,N_305);
nand U502 (N_502,N_296,N_51);
nand U503 (N_503,In_1491,In_1031);
xnor U504 (N_504,In_792,In_605);
nor U505 (N_505,In_614,In_334);
nand U506 (N_506,N_458,In_1462);
and U507 (N_507,In_1353,In_1228);
nor U508 (N_508,In_1138,In_256);
or U509 (N_509,In_1103,In_795);
xor U510 (N_510,In_642,In_1090);
nor U511 (N_511,In_78,N_22);
xnor U512 (N_512,N_96,In_970);
nand U513 (N_513,N_470,In_1266);
xor U514 (N_514,In_210,N_139);
nor U515 (N_515,In_66,In_711);
nor U516 (N_516,In_152,N_492);
nand U517 (N_517,In_646,In_1240);
nand U518 (N_518,In_1296,N_417);
nor U519 (N_519,N_383,N_412);
nor U520 (N_520,N_317,In_1158);
nand U521 (N_521,In_857,In_1174);
and U522 (N_522,In_461,N_401);
nor U523 (N_523,N_319,N_91);
nor U524 (N_524,In_1166,N_58);
nor U525 (N_525,In_28,In_375);
nor U526 (N_526,In_737,In_43);
xor U527 (N_527,In_17,In_1226);
xnor U528 (N_528,N_406,In_401);
nor U529 (N_529,N_49,In_800);
or U530 (N_530,N_407,In_266);
or U531 (N_531,In_1262,In_600);
or U532 (N_532,In_692,N_134);
xnor U533 (N_533,In_1106,In_49);
or U534 (N_534,In_944,In_249);
and U535 (N_535,In_357,In_421);
nand U536 (N_536,N_475,In_497);
and U537 (N_537,N_331,In_508);
and U538 (N_538,In_1097,In_368);
nor U539 (N_539,In_114,In_98);
xnor U540 (N_540,In_271,N_0);
or U541 (N_541,N_116,In_1212);
nand U542 (N_542,In_780,N_313);
or U543 (N_543,In_657,In_1245);
or U544 (N_544,In_1293,In_140);
nand U545 (N_545,In_1437,N_286);
xor U546 (N_546,In_937,In_346);
and U547 (N_547,N_16,N_481);
nand U548 (N_548,N_206,N_418);
nand U549 (N_549,N_441,In_122);
nand U550 (N_550,In_891,In_1361);
nand U551 (N_551,In_1199,In_420);
nor U552 (N_552,In_448,In_1230);
or U553 (N_553,N_374,In_332);
and U554 (N_554,In_1039,In_1493);
nand U555 (N_555,In_127,N_329);
nor U556 (N_556,In_374,In_1038);
nor U557 (N_557,In_529,N_30);
nor U558 (N_558,In_416,N_455);
nor U559 (N_559,In_1485,In_31);
xor U560 (N_560,In_187,N_274);
or U561 (N_561,In_1182,In_1273);
and U562 (N_562,In_1221,In_696);
and U563 (N_563,N_69,N_36);
nor U564 (N_564,N_341,In_1441);
or U565 (N_565,In_488,In_32);
nor U566 (N_566,In_869,N_436);
and U567 (N_567,In_172,In_248);
nand U568 (N_568,In_118,In_1315);
xor U569 (N_569,N_497,In_512);
and U570 (N_570,N_392,In_206);
or U571 (N_571,In_364,In_515);
nor U572 (N_572,In_1488,In_1337);
or U573 (N_573,N_212,In_232);
or U574 (N_574,In_851,N_289);
nor U575 (N_575,N_260,N_413);
nand U576 (N_576,In_55,In_756);
nor U577 (N_577,In_340,N_326);
nand U578 (N_578,In_1079,In_641);
and U579 (N_579,In_1253,N_168);
nand U580 (N_580,In_773,In_176);
and U581 (N_581,In_1382,N_342);
nor U582 (N_582,In_1207,In_826);
or U583 (N_583,In_690,N_254);
xnor U584 (N_584,In_225,In_1384);
and U585 (N_585,N_95,In_669);
and U586 (N_586,N_171,N_442);
or U587 (N_587,In_97,N_496);
or U588 (N_588,In_1489,N_384);
nand U589 (N_589,N_450,N_192);
xor U590 (N_590,N_333,In_209);
and U591 (N_591,In_777,N_82);
xnor U592 (N_592,In_186,N_221);
or U593 (N_593,N_314,In_1263);
and U594 (N_594,In_1146,N_114);
and U595 (N_595,In_166,In_1045);
and U596 (N_596,In_1195,In_255);
nor U597 (N_597,In_723,N_379);
and U598 (N_598,In_388,In_1498);
nand U599 (N_599,In_1313,N_179);
nand U600 (N_600,N_422,In_1475);
and U601 (N_601,In_1092,N_308);
nand U602 (N_602,In_484,N_498);
xnor U603 (N_603,N_390,N_256);
xnor U604 (N_604,In_1201,In_981);
and U605 (N_605,N_354,In_616);
xor U606 (N_606,In_1086,N_125);
and U607 (N_607,N_29,N_287);
nand U608 (N_608,N_376,In_221);
or U609 (N_609,In_889,N_468);
and U610 (N_610,In_199,In_442);
nand U611 (N_611,In_154,In_799);
xor U612 (N_612,N_174,N_394);
nor U613 (N_613,In_158,In_1383);
and U614 (N_614,N_494,In_830);
xnor U615 (N_615,In_319,In_933);
nor U616 (N_616,In_1354,In_812);
nor U617 (N_617,In_469,In_1410);
nor U618 (N_618,In_583,In_953);
xnor U619 (N_619,In_823,In_60);
and U620 (N_620,In_36,N_490);
xnor U621 (N_621,In_941,N_361);
nand U622 (N_622,In_1091,In_574);
and U623 (N_623,N_20,In_1173);
nand U624 (N_624,N_369,In_1357);
nor U625 (N_625,N_595,In_1043);
xor U626 (N_626,In_1358,In_88);
and U627 (N_627,N_421,In_382);
or U628 (N_628,N_119,In_1023);
xor U629 (N_629,In_624,In_913);
nand U630 (N_630,In_938,In_483);
and U631 (N_631,In_1053,In_228);
or U632 (N_632,N_531,N_573);
xnor U633 (N_633,N_591,N_45);
xor U634 (N_634,In_1326,N_440);
nand U635 (N_635,N_208,In_1298);
nand U636 (N_636,In_278,N_429);
nor U637 (N_637,N_517,In_1252);
nor U638 (N_638,N_306,N_81);
and U639 (N_639,In_73,N_395);
nor U640 (N_640,N_397,In_440);
or U641 (N_641,N_589,In_1364);
nand U642 (N_642,In_446,In_929);
nand U643 (N_643,In_649,N_563);
or U644 (N_644,In_725,N_414);
or U645 (N_645,In_896,In_157);
or U646 (N_646,N_515,In_538);
nand U647 (N_647,In_557,N_544);
xor U648 (N_648,N_47,N_602);
and U649 (N_649,N_499,In_710);
nor U650 (N_650,In_292,In_905);
nand U651 (N_651,N_600,In_1380);
or U652 (N_652,In_84,In_713);
and U653 (N_653,In_643,In_951);
and U654 (N_654,In_530,N_249);
and U655 (N_655,In_972,In_312);
or U656 (N_656,In_1183,N_377);
and U657 (N_657,In_1073,In_1185);
nand U658 (N_658,In_95,In_921);
and U659 (N_659,N_83,In_148);
and U660 (N_660,N_343,N_340);
nor U661 (N_661,N_339,N_410);
and U662 (N_662,N_597,N_451);
or U663 (N_663,N_530,N_557);
and U664 (N_664,In_1403,In_693);
xnor U665 (N_665,In_29,N_540);
or U666 (N_666,In_524,N_448);
and U667 (N_667,In_712,In_561);
and U668 (N_668,In_853,In_1490);
nand U669 (N_669,N_447,N_574);
nand U670 (N_670,In_281,N_144);
and U671 (N_671,In_1151,In_942);
or U672 (N_672,In_907,N_378);
nor U673 (N_673,N_488,N_613);
nor U674 (N_674,In_945,In_846);
and U675 (N_675,N_603,In_1404);
and U676 (N_676,N_385,In_89);
or U677 (N_677,In_893,In_162);
xnor U678 (N_678,In_894,N_516);
or U679 (N_679,N_491,N_138);
nor U680 (N_680,In_313,In_254);
nor U681 (N_681,In_1115,N_500);
or U682 (N_682,In_1419,N_587);
and U683 (N_683,N_464,N_509);
or U684 (N_684,In_1213,In_722);
nand U685 (N_685,N_553,N_251);
or U686 (N_686,N_566,In_838);
nand U687 (N_687,N_569,N_380);
nand U688 (N_688,In_276,N_211);
xnor U689 (N_689,N_137,In_880);
xor U690 (N_690,In_864,In_673);
or U691 (N_691,In_454,In_76);
nand U692 (N_692,In_1027,In_902);
nor U693 (N_693,N_493,In_295);
xor U694 (N_694,N_576,In_415);
nand U695 (N_695,N_467,N_482);
or U696 (N_696,N_154,N_608);
or U697 (N_697,N_560,In_27);
or U698 (N_698,In_1132,In_735);
nor U699 (N_699,N_382,N_471);
nor U700 (N_700,N_529,In_1264);
and U701 (N_701,N_105,N_217);
and U702 (N_702,N_248,In_828);
xor U703 (N_703,N_614,N_259);
nor U704 (N_704,N_346,In_1134);
and U705 (N_705,In_1085,N_405);
xor U706 (N_706,In_683,In_156);
nand U707 (N_707,In_1034,In_859);
xor U708 (N_708,In_1037,In_1362);
nand U709 (N_709,In_912,In_1284);
nand U710 (N_710,In_1355,In_586);
and U711 (N_711,N_59,In_979);
and U712 (N_712,N_444,N_393);
nand U713 (N_713,In_814,N_427);
xnor U714 (N_714,In_782,In_872);
nand U715 (N_715,N_265,In_361);
nand U716 (N_716,In_1289,In_155);
or U717 (N_717,In_702,N_232);
nand U718 (N_718,In_1367,In_86);
and U719 (N_719,N_207,In_598);
or U720 (N_720,In_631,In_191);
nand U721 (N_721,In_301,N_505);
or U722 (N_722,N_585,In_1348);
nor U723 (N_723,N_570,In_532);
xor U724 (N_724,N_219,In_419);
or U725 (N_725,N_26,N_176);
and U726 (N_726,N_409,N_571);
nor U727 (N_727,In_467,N_351);
and U728 (N_728,In_1288,N_163);
nor U729 (N_729,In_1429,In_564);
and U730 (N_730,In_133,N_443);
nand U731 (N_731,In_959,N_415);
or U732 (N_732,N_363,N_575);
nor U733 (N_733,In_482,In_691);
nor U734 (N_734,N_541,N_431);
or U735 (N_735,In_895,N_230);
or U736 (N_736,In_178,In_611);
nand U737 (N_737,N_316,In_523);
or U738 (N_738,N_518,N_290);
and U739 (N_739,In_61,N_275);
and U740 (N_740,In_1140,In_1144);
nand U741 (N_741,N_126,In_260);
nand U742 (N_742,In_218,In_15);
nor U743 (N_743,N_424,In_1307);
or U744 (N_744,In_652,In_412);
or U745 (N_745,N_398,In_1492);
xor U746 (N_746,In_1070,In_675);
nand U747 (N_747,N_352,In_1088);
nor U748 (N_748,N_270,N_320);
xor U749 (N_749,N_281,N_521);
nor U750 (N_750,N_619,N_651);
or U751 (N_751,N_736,N_606);
and U752 (N_752,N_568,In_682);
and U753 (N_753,In_1286,N_565);
or U754 (N_754,In_842,N_723);
nand U755 (N_755,N_667,N_477);
nor U756 (N_756,In_560,In_573);
xnor U757 (N_757,N_643,N_170);
and U758 (N_758,In_302,In_1398);
nand U759 (N_759,N_624,N_463);
nor U760 (N_760,N_109,In_1420);
xnor U761 (N_761,N_44,N_749);
or U762 (N_762,In_1061,In_1417);
and U763 (N_763,In_485,N_453);
or U764 (N_764,In_536,In_747);
or U765 (N_765,N_483,In_1461);
xnor U766 (N_766,N_725,N_150);
nand U767 (N_767,N_452,In_744);
nor U768 (N_768,N_349,In_662);
xnor U769 (N_769,N_716,N_244);
nand U770 (N_770,In_593,In_26);
or U771 (N_771,N_648,N_735);
and U772 (N_772,N_598,N_446);
xor U773 (N_773,N_709,N_148);
nand U774 (N_774,In_67,N_131);
and U775 (N_775,In_490,N_702);
nor U776 (N_776,In_1329,In_1413);
xnor U777 (N_777,In_1068,N_546);
and U778 (N_778,N_358,N_681);
and U779 (N_779,In_183,N_291);
xor U780 (N_780,In_922,N_435);
nor U781 (N_781,In_1202,N_672);
nand U782 (N_782,N_368,In_1015);
nand U783 (N_783,N_425,In_1302);
nor U784 (N_784,N_522,In_1421);
or U785 (N_785,N_742,N_57);
or U786 (N_786,In_16,N_607);
nor U787 (N_787,In_676,In_967);
nor U788 (N_788,In_1349,In_463);
xor U789 (N_789,N_130,N_484);
nor U790 (N_790,In_298,In_1171);
or U791 (N_791,N_124,In_576);
and U792 (N_792,N_495,N_616);
xnor U793 (N_793,N_630,In_355);
nor U794 (N_794,In_797,N_578);
xor U795 (N_795,N_93,In_1317);
nand U796 (N_796,In_325,In_1076);
nor U797 (N_797,N_117,In_139);
xor U798 (N_798,In_1446,N_375);
and U799 (N_799,In_1117,N_386);
xnor U800 (N_800,N_534,N_519);
nor U801 (N_801,In_511,In_706);
or U802 (N_802,N_190,In_1105);
or U803 (N_803,In_734,In_100);
nand U804 (N_804,In_1234,N_732);
nor U805 (N_805,N_701,In_923);
xnor U806 (N_806,In_730,In_867);
or U807 (N_807,N_318,In_1126);
and U808 (N_808,N_638,In_1388);
nand U809 (N_809,N_204,N_201);
and U810 (N_810,N_180,In_1456);
or U811 (N_811,In_881,In_274);
xnor U812 (N_812,In_339,In_1333);
or U813 (N_813,In_1422,In_1392);
or U814 (N_814,In_252,N_439);
and U815 (N_815,N_103,In_264);
and U816 (N_816,N_236,In_308);
or U817 (N_817,N_707,N_347);
nand U818 (N_818,N_712,N_400);
xor U819 (N_819,N_508,In_1278);
nor U820 (N_820,N_572,In_333);
nand U821 (N_821,In_656,N_267);
nor U822 (N_822,N_549,N_579);
xnor U823 (N_823,N_640,N_237);
and U824 (N_824,N_641,N_599);
and U825 (N_825,N_620,N_310);
nor U826 (N_826,N_739,In_647);
or U827 (N_827,N_456,N_420);
nor U828 (N_828,N_617,In_1204);
xnor U829 (N_829,N_348,N_520);
nand U830 (N_830,In_161,In_6);
xor U831 (N_831,N_66,In_129);
or U832 (N_832,N_11,In_179);
or U833 (N_833,N_152,N_666);
nor U834 (N_834,N_586,In_282);
and U835 (N_835,In_198,N_523);
nor U836 (N_836,In_745,In_203);
and U837 (N_837,In_1118,In_547);
nand U838 (N_838,N_367,In_952);
or U839 (N_839,In_1341,N_652);
and U840 (N_840,N_199,N_433);
and U841 (N_841,N_545,N_669);
and U842 (N_842,In_559,In_1476);
nor U843 (N_843,N_462,In_500);
nor U844 (N_844,N_710,N_173);
and U845 (N_845,In_1164,N_526);
xor U846 (N_846,N_621,In_977);
nand U847 (N_847,In_1000,In_1218);
or U848 (N_848,In_272,In_185);
nor U849 (N_849,N_703,N_325);
nand U850 (N_850,N_10,N_454);
and U851 (N_851,In_353,In_449);
nand U852 (N_852,In_236,N_78);
and U853 (N_853,N_60,In_1011);
xnor U854 (N_854,In_275,N_416);
nor U855 (N_855,In_1089,In_971);
xor U856 (N_856,N_659,N_503);
xnor U857 (N_857,N_278,N_513);
nor U858 (N_858,In_1401,In_323);
nor U859 (N_859,N_158,In_1113);
nand U860 (N_860,N_636,In_1400);
nor U861 (N_861,In_520,In_373);
nor U862 (N_862,N_524,N_525);
xor U863 (N_863,In_132,N_697);
and U864 (N_864,N_9,N_564);
xor U865 (N_865,In_1184,N_609);
or U866 (N_866,In_444,N_501);
nor U867 (N_867,N_337,N_605);
nor U868 (N_868,In_898,In_1154);
and U869 (N_869,N_647,N_733);
or U870 (N_870,N_592,N_182);
or U871 (N_871,N_411,N_649);
and U872 (N_872,In_824,In_736);
nor U873 (N_873,In_805,In_1062);
xor U874 (N_874,N_112,In_1190);
nor U875 (N_875,N_472,In_1170);
xnor U876 (N_876,N_704,N_727);
nand U877 (N_877,N_671,N_40);
and U878 (N_878,N_590,N_837);
nor U879 (N_879,N_770,In_796);
and U880 (N_880,In_1028,N_626);
xor U881 (N_881,N_686,N_744);
xnor U882 (N_882,In_1304,N_673);
or U883 (N_883,N_668,In_1451);
and U884 (N_884,In_695,In_1007);
nor U885 (N_885,In_1385,In_351);
nand U886 (N_886,N_695,N_836);
nand U887 (N_887,N_486,N_761);
xor U888 (N_888,N_543,N_844);
nand U889 (N_889,N_786,In_956);
xnor U890 (N_890,N_816,N_746);
nor U891 (N_891,In_223,N_774);
xnor U892 (N_892,N_828,N_218);
or U893 (N_893,In_996,N_611);
and U894 (N_894,N_745,In_1438);
nand U895 (N_895,In_44,N_381);
or U896 (N_896,N_776,In_1152);
nor U897 (N_897,N_389,In_1156);
nand U898 (N_898,In_668,In_651);
and U899 (N_899,N_366,N_502);
nor U900 (N_900,In_460,N_855);
nor U901 (N_901,N_860,N_806);
xnor U902 (N_902,N_465,N_231);
nand U903 (N_903,N_404,N_741);
and U904 (N_904,N_789,In_681);
or U905 (N_905,N_677,N_282);
xor U906 (N_906,N_253,In_678);
nor U907 (N_907,N_89,N_740);
nand U908 (N_908,N_824,In_194);
and U909 (N_909,N_773,N_682);
or U910 (N_910,In_1455,N_327);
xnor U911 (N_911,N_532,N_330);
xnor U912 (N_912,N_556,In_738);
nand U913 (N_913,N_699,In_995);
or U914 (N_914,N_863,N_555);
or U915 (N_915,N_657,N_775);
nand U916 (N_916,N_788,N_17);
and U917 (N_917,N_752,N_852);
and U918 (N_918,In_13,In_1108);
nand U919 (N_919,N_459,N_7);
xnor U920 (N_920,N_506,N_840);
and U921 (N_921,N_756,In_1029);
xnor U922 (N_922,In_438,In_142);
or U923 (N_923,In_330,N_757);
nand U924 (N_924,N_166,N_345);
and U925 (N_925,N_711,N_528);
and U926 (N_926,N_101,N_653);
nand U927 (N_927,In_1290,N_815);
xor U928 (N_928,N_567,In_554);
nor U929 (N_929,N_250,In_1369);
nor U930 (N_930,N_539,In_310);
xnor U931 (N_931,In_1282,N_466);
and U932 (N_932,N_793,N_848);
nor U933 (N_933,N_698,In_193);
nor U934 (N_934,N_737,N_683);
nor U935 (N_935,In_731,In_12);
or U936 (N_936,N_268,In_91);
or U937 (N_937,In_579,N_684);
xnor U938 (N_938,N_438,N_845);
and U939 (N_939,In_688,N_449);
and U940 (N_940,N_618,N_371);
nand U941 (N_941,N_817,N_141);
and U942 (N_942,N_796,N_646);
xor U943 (N_943,In_1026,In_103);
nor U944 (N_944,In_1040,In_1235);
or U945 (N_945,N_593,N_759);
or U946 (N_946,In_602,N_720);
nor U947 (N_947,N_536,In_305);
xor U948 (N_948,In_885,In_1143);
nand U949 (N_949,N_859,N_718);
nor U950 (N_950,In_626,In_528);
or U951 (N_951,N_72,In_428);
nand U952 (N_952,N_512,N_419);
nor U953 (N_953,N_315,N_691);
nor U954 (N_954,N_706,N_751);
nor U955 (N_955,N_293,In_104);
nor U956 (N_956,N_507,In_106);
xnor U957 (N_957,N_301,N_758);
xor U958 (N_958,N_868,N_696);
and U959 (N_959,N_62,N_445);
or U960 (N_960,N_854,In_549);
or U961 (N_961,In_422,In_627);
nand U962 (N_962,In_565,N_838);
and U963 (N_963,N_391,In_761);
and U964 (N_964,N_784,N_362);
or U965 (N_965,In_1125,In_1472);
nor U966 (N_966,In_427,N_297);
or U967 (N_967,In_173,N_825);
nor U968 (N_968,N_835,In_471);
or U969 (N_969,N_777,N_856);
xnor U970 (N_970,N_510,In_1311);
xnor U971 (N_971,In_1340,N_247);
nor U972 (N_972,In_991,N_791);
xnor U973 (N_973,N_785,N_263);
nor U974 (N_974,N_461,N_487);
nand U975 (N_975,N_332,In_498);
xnor U976 (N_976,N_511,In_115);
nor U977 (N_977,In_527,N_820);
xor U978 (N_978,In_426,In_535);
and U979 (N_979,N_581,In_159);
nor U980 (N_980,In_1150,N_867);
and U981 (N_981,N_548,In_400);
xor U982 (N_982,In_821,N_402);
or U983 (N_983,N_870,N_715);
nand U984 (N_984,N_850,In_597);
xnor U985 (N_985,N_437,In_1017);
xor U986 (N_986,In_998,N_277);
nor U987 (N_987,N_680,N_399);
xor U988 (N_988,N_43,N_851);
nor U989 (N_989,N_181,In_1415);
and U990 (N_990,N_713,N_527);
or U991 (N_991,N_692,In_1335);
xor U992 (N_992,N_804,N_678);
or U993 (N_993,N_403,N_284);
and U994 (N_994,N_782,N_311);
and U995 (N_995,In_453,N_61);
and U996 (N_996,N_434,In_1219);
xor U997 (N_997,In_1148,N_679);
xnor U998 (N_998,N_762,N_627);
and U999 (N_999,In_1238,N_753);
or U1000 (N_1000,In_836,N_877);
nand U1001 (N_1001,N_908,N_853);
nand U1002 (N_1002,N_931,N_768);
nand U1003 (N_1003,N_665,N_552);
or U1004 (N_1004,In_1265,N_996);
xnor U1005 (N_1005,In_1216,N_974);
and U1006 (N_1006,In_1499,N_821);
and U1007 (N_1007,In_776,N_705);
nand U1008 (N_1008,N_604,N_950);
xor U1009 (N_1009,N_919,In_324);
or U1010 (N_1010,In_41,N_798);
nor U1011 (N_1011,N_623,N_730);
or U1012 (N_1012,N_955,N_309);
nand U1013 (N_1013,N_968,In_901);
nand U1014 (N_1014,N_901,In_1379);
xnor U1015 (N_1015,N_926,N_792);
or U1016 (N_1016,N_246,N_993);
nor U1017 (N_1017,N_960,In_1363);
nand U1018 (N_1018,N_360,N_797);
nor U1019 (N_1019,In_1142,In_1059);
nand U1020 (N_1020,N_780,N_790);
nor U1021 (N_1021,N_846,N_989);
nand U1022 (N_1022,N_779,In_1305);
nor U1023 (N_1023,N_862,In_1330);
or U1024 (N_1024,In_906,N_822);
and U1025 (N_1025,N_675,N_934);
nor U1026 (N_1026,In_507,N_584);
nand U1027 (N_1027,N_930,In_243);
and U1028 (N_1028,N_750,In_1450);
xnor U1029 (N_1029,N_808,In_750);
nor U1030 (N_1030,In_0,In_34);
or U1031 (N_1031,N_661,N_582);
or U1032 (N_1032,N_726,N_830);
nor U1033 (N_1033,N_304,N_771);
or U1034 (N_1034,N_805,N_355);
and U1035 (N_1035,In_1009,In_1136);
nor U1036 (N_1036,In_840,In_606);
and U1037 (N_1037,In_1332,N_964);
and U1038 (N_1038,N_970,N_879);
xor U1039 (N_1039,N_940,N_906);
or U1040 (N_1040,In_1123,In_105);
and U1041 (N_1041,N_489,N_766);
xnor U1042 (N_1042,N_396,In_619);
nor U1043 (N_1043,N_205,N_864);
nand U1044 (N_1044,N_829,N_162);
nand U1045 (N_1045,In_245,In_424);
or U1046 (N_1046,N_928,N_980);
nand U1047 (N_1047,N_688,N_975);
nor U1048 (N_1048,N_734,N_887);
xnor U1049 (N_1049,N_947,N_935);
and U1050 (N_1050,In_868,N_457);
xnor U1051 (N_1051,N_832,N_984);
or U1052 (N_1052,In_638,N_801);
nor U1053 (N_1053,N_842,N_760);
nand U1054 (N_1054,N_834,N_615);
nor U1055 (N_1055,N_662,In_939);
or U1056 (N_1056,N_878,N_504);
xor U1057 (N_1057,N_802,N_430);
or U1058 (N_1058,N_841,N_478);
nor U1059 (N_1059,N_663,N_239);
xor U1060 (N_1060,N_694,In_1287);
nand U1061 (N_1061,In_229,N_897);
and U1062 (N_1062,N_537,In_1001);
xor U1063 (N_1063,N_344,In_575);
xnor U1064 (N_1064,N_910,In_1321);
and U1065 (N_1065,In_578,N_889);
xor U1066 (N_1066,In_858,In_329);
and U1067 (N_1067,N_474,N_872);
or U1068 (N_1068,N_833,N_823);
nand U1069 (N_1069,N_767,N_861);
and U1070 (N_1070,N_812,N_818);
nand U1071 (N_1071,In_238,In_1161);
or U1072 (N_1072,N_976,N_408);
nand U1073 (N_1073,N_476,N_550);
nand U1074 (N_1074,N_225,In_543);
nand U1075 (N_1075,N_977,N_943);
or U1076 (N_1076,N_714,N_670);
nor U1077 (N_1077,In_200,N_900);
nor U1078 (N_1078,In_1145,N_238);
nand U1079 (N_1079,In_732,N_728);
or U1080 (N_1080,N_982,In_1480);
and U1081 (N_1081,N_942,N_365);
xnor U1082 (N_1082,N_987,N_622);
nand U1083 (N_1083,In_270,N_874);
or U1084 (N_1084,N_986,N_927);
or U1085 (N_1085,N_324,N_432);
or U1086 (N_1086,N_952,In_540);
nand U1087 (N_1087,N_722,N_921);
and U1088 (N_1088,In_1063,In_634);
nor U1089 (N_1089,In_1257,N_883);
or U1090 (N_1090,In_1454,N_200);
or U1091 (N_1091,N_280,In_994);
and U1092 (N_1092,N_915,In_69);
nor U1093 (N_1093,In_1020,N_690);
xor U1094 (N_1094,In_1279,N_2);
or U1095 (N_1095,N_634,N_558);
nand U1096 (N_1096,N_693,N_787);
and U1097 (N_1097,In_358,N_876);
and U1098 (N_1098,In_410,N_895);
nand U1099 (N_1099,In_1032,N_764);
nand U1100 (N_1100,N_25,N_577);
or U1101 (N_1101,N_810,N_925);
nand U1102 (N_1102,N_729,N_272);
nor U1103 (N_1103,N_932,In_145);
or U1104 (N_1104,N_847,N_685);
nor U1105 (N_1105,In_501,In_969);
xnor U1106 (N_1106,N_769,In_1130);
and U1107 (N_1107,N_891,In_948);
nand U1108 (N_1108,N_142,N_708);
nand U1109 (N_1109,N_933,N_916);
and U1110 (N_1110,N_966,N_988);
xnor U1111 (N_1111,N_999,N_914);
nor U1112 (N_1112,N_807,N_387);
xnor U1113 (N_1113,N_650,N_936);
nor U1114 (N_1114,N_644,N_763);
xnor U1115 (N_1115,N_654,N_898);
nand U1116 (N_1116,N_295,In_288);
and U1117 (N_1117,N_951,N_994);
or U1118 (N_1118,In_982,N_985);
xnor U1119 (N_1119,In_1153,N_866);
or U1120 (N_1120,In_760,N_157);
nor U1121 (N_1121,N_896,N_583);
xor U1122 (N_1122,N_77,In_343);
xnor U1123 (N_1123,N_857,N_962);
xnor U1124 (N_1124,N_965,N_473);
and U1125 (N_1125,In_1010,N_1120);
or U1126 (N_1126,In_297,In_572);
or U1127 (N_1127,N_731,N_1068);
and U1128 (N_1128,N_178,N_814);
or U1129 (N_1129,N_783,N_559);
and U1130 (N_1130,N_1054,N_1084);
nor U1131 (N_1131,In_802,In_1452);
xnor U1132 (N_1132,N_748,N_1081);
or U1133 (N_1133,N_1056,N_1052);
nor U1134 (N_1134,N_1048,N_1014);
or U1135 (N_1135,In_1444,N_871);
xnor U1136 (N_1136,N_197,In_441);
xor U1137 (N_1137,N_1106,N_1003);
and U1138 (N_1138,N_485,N_1079);
or U1139 (N_1139,In_1319,N_827);
xnor U1140 (N_1140,N_1102,N_388);
xor U1141 (N_1141,N_596,N_1118);
xnor U1142 (N_1142,In_622,In_468);
xnor U1143 (N_1143,N_1002,N_1123);
nand U1144 (N_1144,N_813,N_918);
nor U1145 (N_1145,N_547,In_121);
nand U1146 (N_1146,N_1031,In_381);
nor U1147 (N_1147,N_886,N_997);
and U1148 (N_1148,N_967,N_1093);
xnor U1149 (N_1149,N_1059,In_1254);
xor U1150 (N_1150,N_1089,N_719);
nand U1151 (N_1151,N_849,N_911);
nor U1152 (N_1152,N_875,N_1096);
nor U1153 (N_1153,N_972,N_1122);
xor U1154 (N_1154,N_551,N_372);
xor U1155 (N_1155,N_1070,N_958);
or U1156 (N_1156,N_561,N_1001);
and U1157 (N_1157,N_71,In_1074);
or U1158 (N_1158,N_136,In_677);
nand U1159 (N_1159,N_1075,N_535);
xnor U1160 (N_1160,In_391,In_1318);
xnor U1161 (N_1161,N_298,N_1022);
nand U1162 (N_1162,N_601,N_924);
or U1163 (N_1163,N_1078,N_700);
and U1164 (N_1164,N_979,N_258);
and U1165 (N_1165,N_542,N_479);
xnor U1166 (N_1166,N_1083,N_1107);
nand U1167 (N_1167,N_948,N_1063);
nand U1168 (N_1168,N_1029,N_1038);
or U1169 (N_1169,N_755,N_1119);
or U1170 (N_1170,N_1097,N_956);
nor U1171 (N_1171,N_689,N_1042);
nor U1172 (N_1172,N_922,N_469);
xnor U1173 (N_1173,N_1039,N_1017);
nor U1174 (N_1174,N_907,N_880);
or U1175 (N_1175,N_941,N_839);
nor U1176 (N_1176,N_164,N_645);
nand U1177 (N_1177,N_1064,N_1000);
nor U1178 (N_1178,N_610,In_473);
nor U1179 (N_1179,N_949,N_580);
and U1180 (N_1180,N_202,In_1376);
and U1181 (N_1181,N_1104,N_364);
or U1182 (N_1182,N_245,N_899);
or U1183 (N_1183,In_1467,N_674);
nor U1184 (N_1184,N_1032,N_1036);
and U1185 (N_1185,In_1055,N_717);
or U1186 (N_1186,N_905,N_1086);
or U1187 (N_1187,N_1105,N_917);
xnor U1188 (N_1188,N_743,N_843);
and U1189 (N_1189,N_428,N_177);
xnor U1190 (N_1190,N_1037,In_751);
xor U1191 (N_1191,In_844,N_1111);
nand U1192 (N_1192,N_68,N_1094);
and U1193 (N_1193,N_873,N_938);
nor U1194 (N_1194,N_778,N_894);
nand U1195 (N_1195,N_338,N_920);
and U1196 (N_1196,N_971,N_203);
nor U1197 (N_1197,N_1114,N_865);
nor U1198 (N_1198,N_800,N_639);
or U1199 (N_1199,In_1081,N_220);
nand U1200 (N_1200,In_825,N_961);
and U1201 (N_1201,N_959,N_426);
nand U1202 (N_1202,N_594,N_893);
or U1203 (N_1203,In_733,N_1085);
nor U1204 (N_1204,N_1072,In_53);
or U1205 (N_1205,N_747,N_892);
and U1206 (N_1206,N_64,N_1008);
xnor U1207 (N_1207,N_923,N_1100);
or U1208 (N_1208,N_995,N_1099);
nand U1209 (N_1209,N_1047,N_969);
nor U1210 (N_1210,N_881,N_946);
or U1211 (N_1211,N_1091,N_1103);
nand U1212 (N_1212,N_1098,In_1019);
nand U1213 (N_1213,N_885,N_963);
and U1214 (N_1214,N_658,In_818);
nor U1215 (N_1215,N_1061,In_1191);
nand U1216 (N_1216,N_1053,N_1007);
nor U1217 (N_1217,In_403,N_1016);
nor U1218 (N_1218,N_1050,N_772);
nor U1219 (N_1219,N_1033,N_811);
nand U1220 (N_1220,N_795,In_1479);
nor U1221 (N_1221,In_1198,N_1049);
nand U1222 (N_1222,N_294,N_939);
nand U1223 (N_1223,N_913,N_1090);
nor U1224 (N_1224,N_562,N_944);
xnor U1225 (N_1225,N_1076,N_423);
xnor U1226 (N_1226,N_1045,N_94);
and U1227 (N_1227,N_799,N_957);
and U1228 (N_1228,N_781,In_1277);
xor U1229 (N_1229,N_1124,N_1028);
xnor U1230 (N_1230,In_169,N_909);
and U1231 (N_1231,N_635,N_1067);
nand U1232 (N_1232,N_15,N_809);
and U1233 (N_1233,N_1021,In_1075);
nor U1234 (N_1234,N_831,N_687);
nor U1235 (N_1235,N_169,N_1010);
nand U1236 (N_1236,N_1030,N_664);
and U1237 (N_1237,In_284,N_223);
and U1238 (N_1238,In_580,N_612);
and U1239 (N_1239,N_1046,N_1115);
nor U1240 (N_1240,In_79,N_1025);
nor U1241 (N_1241,N_1088,N_1057);
or U1242 (N_1242,N_981,N_1060);
xor U1243 (N_1243,N_902,N_642);
xnor U1244 (N_1244,N_1026,In_171);
nand U1245 (N_1245,In_542,In_1077);
nor U1246 (N_1246,N_884,N_625);
xnor U1247 (N_1247,N_637,In_949);
nor U1248 (N_1248,N_912,N_629);
and U1249 (N_1249,N_285,N_1112);
or U1250 (N_1250,In_835,In_247);
or U1251 (N_1251,N_1149,N_1218);
nor U1252 (N_1252,In_888,N_1147);
xnor U1253 (N_1253,N_1182,N_990);
nand U1254 (N_1254,N_1020,N_353);
and U1255 (N_1255,N_234,N_1035);
and U1256 (N_1256,N_1233,N_1196);
and U1257 (N_1257,N_1205,N_1171);
nand U1258 (N_1258,N_1176,In_903);
nor U1259 (N_1259,N_1141,N_1209);
and U1260 (N_1260,N_633,N_1129);
or U1261 (N_1261,In_397,In_110);
and U1262 (N_1262,N_1126,N_1136);
and U1263 (N_1263,N_929,N_983);
xnor U1264 (N_1264,In_250,N_1069);
or U1265 (N_1265,In_960,N_954);
or U1266 (N_1266,N_660,N_123);
or U1267 (N_1267,In_968,N_724);
or U1268 (N_1268,N_1202,N_1197);
and U1269 (N_1269,N_261,N_1101);
xnor U1270 (N_1270,In_1275,N_1154);
nor U1271 (N_1271,N_18,N_1128);
or U1272 (N_1272,N_1121,N_1234);
nor U1273 (N_1273,N_1095,N_1221);
or U1274 (N_1274,N_1242,N_656);
and U1275 (N_1275,In_1327,N_1236);
nor U1276 (N_1276,N_1212,N_1181);
nor U1277 (N_1277,N_937,N_1201);
or U1278 (N_1278,In_1267,N_1133);
and U1279 (N_1279,N_826,N_1164);
and U1280 (N_1280,In_1359,N_1051);
nor U1281 (N_1281,N_1130,N_1208);
or U1282 (N_1282,N_1240,N_1206);
xnor U1283 (N_1283,N_1011,N_533);
nand U1284 (N_1284,N_676,N_754);
xor U1285 (N_1285,N_1148,N_1169);
or U1286 (N_1286,N_480,N_1157);
and U1287 (N_1287,N_1082,N_1155);
xor U1288 (N_1288,N_1023,N_1195);
or U1289 (N_1289,N_1204,In_1474);
xor U1290 (N_1290,N_1138,N_1062);
nor U1291 (N_1291,N_1214,N_1249);
or U1292 (N_1292,N_1170,N_1151);
xor U1293 (N_1293,N_1211,N_858);
and U1294 (N_1294,N_1243,N_1006);
and U1295 (N_1295,N_1220,N_973);
xnor U1296 (N_1296,N_1188,N_460);
nor U1297 (N_1297,N_56,N_1139);
nand U1298 (N_1298,N_1230,N_1232);
or U1299 (N_1299,N_1215,N_1179);
and U1300 (N_1300,In_759,N_655);
xnor U1301 (N_1301,N_1241,N_869);
and U1302 (N_1302,In_749,N_356);
nor U1303 (N_1303,N_1018,N_1077);
nand U1304 (N_1304,N_1041,N_904);
or U1305 (N_1305,N_1127,N_1116);
xnor U1306 (N_1306,N_1131,N_1237);
nand U1307 (N_1307,N_992,N_998);
and U1308 (N_1308,In_848,N_1175);
nand U1309 (N_1309,N_1192,N_882);
xor U1310 (N_1310,N_1013,N_1012);
nor U1311 (N_1311,N_1183,N_1189);
nor U1312 (N_1312,N_1108,N_628);
or U1313 (N_1313,N_888,N_1140);
nor U1314 (N_1314,N_794,N_1113);
nor U1315 (N_1315,N_1247,N_1224);
xor U1316 (N_1316,N_1024,N_1027);
xnor U1317 (N_1317,N_1199,N_1225);
or U1318 (N_1318,In_550,N_1172);
and U1319 (N_1319,N_631,N_1227);
nand U1320 (N_1320,In_59,N_1087);
nor U1321 (N_1321,N_1207,N_1226);
nand U1322 (N_1322,N_890,N_1040);
xnor U1323 (N_1323,N_1210,In_299);
nand U1324 (N_1324,N_1117,N_1159);
nor U1325 (N_1325,N_1137,N_1167);
nand U1326 (N_1326,N_953,N_1173);
nor U1327 (N_1327,N_1055,In_1223);
xor U1328 (N_1328,N_1191,N_538);
and U1329 (N_1329,N_1019,N_1193);
nor U1330 (N_1330,N_1248,N_1066);
nor U1331 (N_1331,In_993,N_1216);
and U1332 (N_1332,N_1213,N_632);
nor U1333 (N_1333,N_1160,N_1244);
and U1334 (N_1334,N_1246,N_1198);
or U1335 (N_1335,N_1200,N_1142);
nor U1336 (N_1336,N_1110,N_1150);
nor U1337 (N_1337,In_192,N_1080);
or U1338 (N_1338,In_443,N_1239);
and U1339 (N_1339,In_931,N_1229);
xnor U1340 (N_1340,N_1009,N_1174);
nand U1341 (N_1341,N_1144,N_1168);
nor U1342 (N_1342,N_1235,N_1222);
xnor U1343 (N_1343,N_991,N_1165);
xnor U1344 (N_1344,N_160,N_1158);
xnor U1345 (N_1345,N_803,N_1109);
nor U1346 (N_1346,N_1005,N_1043);
nand U1347 (N_1347,N_1146,N_738);
nor U1348 (N_1348,N_1223,N_1162);
or U1349 (N_1349,N_1073,N_1152);
nand U1350 (N_1350,N_1245,N_1135);
nand U1351 (N_1351,N_1219,N_1004);
or U1352 (N_1352,N_1163,N_1132);
nand U1353 (N_1353,N_514,In_1427);
nand U1354 (N_1354,N_721,In_1270);
and U1355 (N_1355,In_216,N_1190);
nor U1356 (N_1356,N_1187,N_1231);
nand U1357 (N_1357,N_323,N_1180);
nand U1358 (N_1358,N_1044,N_978);
nand U1359 (N_1359,N_945,N_1156);
or U1360 (N_1360,N_903,N_1153);
xnor U1361 (N_1361,N_765,N_1166);
nor U1362 (N_1362,In_244,N_1185);
nand U1363 (N_1363,N_1145,N_1203);
xor U1364 (N_1364,N_1065,N_1134);
xnor U1365 (N_1365,N_1034,N_1143);
xnor U1366 (N_1366,N_1178,N_819);
nor U1367 (N_1367,N_1238,N_1074);
or U1368 (N_1368,N_1177,N_1161);
nor U1369 (N_1369,N_1125,N_1184);
xor U1370 (N_1370,N_1071,N_1092);
and U1371 (N_1371,N_1186,N_554);
and U1372 (N_1372,N_1228,N_1217);
xnor U1373 (N_1373,N_1058,N_588);
or U1374 (N_1374,N_1015,N_1194);
or U1375 (N_1375,N_1273,N_1291);
xnor U1376 (N_1376,N_1257,N_1353);
nor U1377 (N_1377,N_1347,N_1290);
xnor U1378 (N_1378,N_1306,N_1331);
xor U1379 (N_1379,N_1364,N_1345);
nor U1380 (N_1380,N_1368,N_1318);
nor U1381 (N_1381,N_1283,N_1262);
and U1382 (N_1382,N_1374,N_1354);
or U1383 (N_1383,N_1363,N_1281);
or U1384 (N_1384,N_1298,N_1282);
and U1385 (N_1385,N_1315,N_1277);
and U1386 (N_1386,N_1333,N_1320);
xnor U1387 (N_1387,N_1335,N_1324);
and U1388 (N_1388,N_1362,N_1373);
nor U1389 (N_1389,N_1321,N_1254);
nor U1390 (N_1390,N_1270,N_1356);
nor U1391 (N_1391,N_1312,N_1371);
nor U1392 (N_1392,N_1302,N_1310);
and U1393 (N_1393,N_1292,N_1288);
nor U1394 (N_1394,N_1266,N_1342);
nor U1395 (N_1395,N_1369,N_1326);
and U1396 (N_1396,N_1286,N_1336);
or U1397 (N_1397,N_1264,N_1260);
nand U1398 (N_1398,N_1349,N_1276);
nand U1399 (N_1399,N_1337,N_1329);
nor U1400 (N_1400,N_1304,N_1370);
and U1401 (N_1401,N_1278,N_1358);
and U1402 (N_1402,N_1268,N_1322);
and U1403 (N_1403,N_1250,N_1359);
xnor U1404 (N_1404,N_1305,N_1280);
xor U1405 (N_1405,N_1323,N_1297);
and U1406 (N_1406,N_1293,N_1267);
nor U1407 (N_1407,N_1272,N_1372);
nand U1408 (N_1408,N_1301,N_1279);
and U1409 (N_1409,N_1289,N_1299);
xnor U1410 (N_1410,N_1346,N_1367);
and U1411 (N_1411,N_1316,N_1355);
or U1412 (N_1412,N_1309,N_1338);
or U1413 (N_1413,N_1259,N_1339);
or U1414 (N_1414,N_1319,N_1303);
or U1415 (N_1415,N_1296,N_1317);
and U1416 (N_1416,N_1307,N_1311);
and U1417 (N_1417,N_1366,N_1357);
and U1418 (N_1418,N_1334,N_1365);
nor U1419 (N_1419,N_1344,N_1325);
xor U1420 (N_1420,N_1251,N_1255);
and U1421 (N_1421,N_1275,N_1327);
nand U1422 (N_1422,N_1352,N_1253);
and U1423 (N_1423,N_1265,N_1343);
and U1424 (N_1424,N_1287,N_1314);
or U1425 (N_1425,N_1351,N_1294);
xnor U1426 (N_1426,N_1332,N_1274);
xor U1427 (N_1427,N_1269,N_1300);
xor U1428 (N_1428,N_1252,N_1271);
nand U1429 (N_1429,N_1258,N_1360);
xor U1430 (N_1430,N_1328,N_1285);
xor U1431 (N_1431,N_1295,N_1350);
nor U1432 (N_1432,N_1330,N_1263);
nor U1433 (N_1433,N_1340,N_1308);
or U1434 (N_1434,N_1261,N_1348);
or U1435 (N_1435,N_1313,N_1256);
and U1436 (N_1436,N_1341,N_1361);
xnor U1437 (N_1437,N_1284,N_1255);
xor U1438 (N_1438,N_1264,N_1354);
nor U1439 (N_1439,N_1334,N_1368);
nand U1440 (N_1440,N_1281,N_1293);
xnor U1441 (N_1441,N_1257,N_1306);
nor U1442 (N_1442,N_1299,N_1286);
or U1443 (N_1443,N_1353,N_1337);
xnor U1444 (N_1444,N_1342,N_1334);
nor U1445 (N_1445,N_1282,N_1250);
xor U1446 (N_1446,N_1265,N_1272);
xor U1447 (N_1447,N_1349,N_1304);
nor U1448 (N_1448,N_1311,N_1368);
xnor U1449 (N_1449,N_1341,N_1372);
and U1450 (N_1450,N_1292,N_1265);
nor U1451 (N_1451,N_1291,N_1365);
or U1452 (N_1452,N_1358,N_1357);
and U1453 (N_1453,N_1359,N_1373);
and U1454 (N_1454,N_1357,N_1287);
or U1455 (N_1455,N_1303,N_1269);
xor U1456 (N_1456,N_1358,N_1270);
nor U1457 (N_1457,N_1272,N_1359);
and U1458 (N_1458,N_1325,N_1251);
nand U1459 (N_1459,N_1293,N_1366);
nor U1460 (N_1460,N_1334,N_1270);
nand U1461 (N_1461,N_1287,N_1313);
xor U1462 (N_1462,N_1335,N_1264);
nand U1463 (N_1463,N_1261,N_1319);
or U1464 (N_1464,N_1330,N_1370);
xnor U1465 (N_1465,N_1359,N_1361);
or U1466 (N_1466,N_1331,N_1302);
nor U1467 (N_1467,N_1302,N_1333);
nor U1468 (N_1468,N_1355,N_1305);
nand U1469 (N_1469,N_1358,N_1306);
or U1470 (N_1470,N_1305,N_1353);
nor U1471 (N_1471,N_1310,N_1263);
or U1472 (N_1472,N_1305,N_1266);
nor U1473 (N_1473,N_1304,N_1310);
nand U1474 (N_1474,N_1258,N_1334);
xnor U1475 (N_1475,N_1346,N_1310);
xor U1476 (N_1476,N_1259,N_1250);
or U1477 (N_1477,N_1367,N_1270);
and U1478 (N_1478,N_1366,N_1308);
nand U1479 (N_1479,N_1323,N_1287);
or U1480 (N_1480,N_1367,N_1332);
xnor U1481 (N_1481,N_1285,N_1345);
nand U1482 (N_1482,N_1347,N_1315);
nor U1483 (N_1483,N_1316,N_1250);
nor U1484 (N_1484,N_1261,N_1332);
nand U1485 (N_1485,N_1302,N_1297);
or U1486 (N_1486,N_1270,N_1316);
and U1487 (N_1487,N_1367,N_1311);
nand U1488 (N_1488,N_1344,N_1307);
or U1489 (N_1489,N_1357,N_1276);
nor U1490 (N_1490,N_1305,N_1371);
and U1491 (N_1491,N_1312,N_1313);
nor U1492 (N_1492,N_1305,N_1336);
nand U1493 (N_1493,N_1291,N_1309);
xor U1494 (N_1494,N_1336,N_1311);
or U1495 (N_1495,N_1279,N_1254);
nand U1496 (N_1496,N_1365,N_1301);
and U1497 (N_1497,N_1288,N_1356);
xnor U1498 (N_1498,N_1350,N_1254);
xor U1499 (N_1499,N_1284,N_1294);
nand U1500 (N_1500,N_1495,N_1375);
and U1501 (N_1501,N_1383,N_1405);
and U1502 (N_1502,N_1435,N_1494);
and U1503 (N_1503,N_1473,N_1421);
xor U1504 (N_1504,N_1396,N_1482);
xor U1505 (N_1505,N_1417,N_1378);
and U1506 (N_1506,N_1377,N_1387);
nor U1507 (N_1507,N_1457,N_1449);
xnor U1508 (N_1508,N_1413,N_1477);
and U1509 (N_1509,N_1462,N_1474);
or U1510 (N_1510,N_1490,N_1382);
nor U1511 (N_1511,N_1437,N_1480);
or U1512 (N_1512,N_1426,N_1386);
or U1513 (N_1513,N_1436,N_1452);
nand U1514 (N_1514,N_1418,N_1476);
nor U1515 (N_1515,N_1468,N_1401);
or U1516 (N_1516,N_1407,N_1428);
nand U1517 (N_1517,N_1464,N_1486);
xnor U1518 (N_1518,N_1489,N_1433);
xnor U1519 (N_1519,N_1414,N_1499);
xnor U1520 (N_1520,N_1496,N_1458);
nand U1521 (N_1521,N_1424,N_1429);
nand U1522 (N_1522,N_1438,N_1451);
or U1523 (N_1523,N_1453,N_1397);
xnor U1524 (N_1524,N_1445,N_1446);
nand U1525 (N_1525,N_1393,N_1406);
xnor U1526 (N_1526,N_1427,N_1416);
xnor U1527 (N_1527,N_1402,N_1487);
and U1528 (N_1528,N_1450,N_1390);
nand U1529 (N_1529,N_1432,N_1465);
nor U1530 (N_1530,N_1442,N_1481);
and U1531 (N_1531,N_1431,N_1485);
or U1532 (N_1532,N_1392,N_1430);
xnor U1533 (N_1533,N_1471,N_1479);
or U1534 (N_1534,N_1423,N_1381);
nor U1535 (N_1535,N_1439,N_1394);
nand U1536 (N_1536,N_1475,N_1420);
and U1537 (N_1537,N_1440,N_1409);
or U1538 (N_1538,N_1376,N_1408);
and U1539 (N_1539,N_1460,N_1410);
xnor U1540 (N_1540,N_1443,N_1498);
xnor U1541 (N_1541,N_1455,N_1472);
nand U1542 (N_1542,N_1447,N_1483);
or U1543 (N_1543,N_1384,N_1456);
xor U1544 (N_1544,N_1415,N_1461);
xnor U1545 (N_1545,N_1478,N_1484);
nor U1546 (N_1546,N_1389,N_1463);
and U1547 (N_1547,N_1493,N_1441);
or U1548 (N_1548,N_1391,N_1422);
xor U1549 (N_1549,N_1492,N_1497);
nor U1550 (N_1550,N_1403,N_1385);
nand U1551 (N_1551,N_1425,N_1448);
or U1552 (N_1552,N_1488,N_1466);
and U1553 (N_1553,N_1380,N_1459);
nand U1554 (N_1554,N_1399,N_1379);
nor U1555 (N_1555,N_1411,N_1469);
and U1556 (N_1556,N_1388,N_1454);
xor U1557 (N_1557,N_1395,N_1434);
nand U1558 (N_1558,N_1398,N_1412);
nand U1559 (N_1559,N_1470,N_1444);
nand U1560 (N_1560,N_1467,N_1400);
nand U1561 (N_1561,N_1404,N_1419);
xor U1562 (N_1562,N_1491,N_1486);
or U1563 (N_1563,N_1376,N_1420);
nor U1564 (N_1564,N_1407,N_1449);
xnor U1565 (N_1565,N_1409,N_1464);
nor U1566 (N_1566,N_1485,N_1419);
nor U1567 (N_1567,N_1436,N_1402);
xnor U1568 (N_1568,N_1419,N_1493);
or U1569 (N_1569,N_1456,N_1399);
or U1570 (N_1570,N_1409,N_1395);
nor U1571 (N_1571,N_1455,N_1383);
and U1572 (N_1572,N_1383,N_1498);
nand U1573 (N_1573,N_1375,N_1438);
xor U1574 (N_1574,N_1420,N_1411);
and U1575 (N_1575,N_1406,N_1381);
xor U1576 (N_1576,N_1399,N_1455);
nand U1577 (N_1577,N_1397,N_1386);
or U1578 (N_1578,N_1458,N_1396);
xnor U1579 (N_1579,N_1482,N_1450);
nor U1580 (N_1580,N_1387,N_1404);
xor U1581 (N_1581,N_1460,N_1491);
xor U1582 (N_1582,N_1426,N_1473);
and U1583 (N_1583,N_1407,N_1416);
nor U1584 (N_1584,N_1459,N_1458);
xor U1585 (N_1585,N_1443,N_1493);
and U1586 (N_1586,N_1449,N_1434);
nor U1587 (N_1587,N_1484,N_1459);
nor U1588 (N_1588,N_1498,N_1445);
or U1589 (N_1589,N_1430,N_1405);
or U1590 (N_1590,N_1493,N_1457);
xnor U1591 (N_1591,N_1497,N_1493);
xnor U1592 (N_1592,N_1475,N_1473);
xor U1593 (N_1593,N_1388,N_1399);
nand U1594 (N_1594,N_1375,N_1382);
and U1595 (N_1595,N_1442,N_1424);
nor U1596 (N_1596,N_1399,N_1384);
and U1597 (N_1597,N_1395,N_1412);
xor U1598 (N_1598,N_1495,N_1419);
nor U1599 (N_1599,N_1425,N_1469);
nor U1600 (N_1600,N_1429,N_1438);
nand U1601 (N_1601,N_1412,N_1481);
and U1602 (N_1602,N_1436,N_1489);
nand U1603 (N_1603,N_1444,N_1436);
nor U1604 (N_1604,N_1420,N_1429);
and U1605 (N_1605,N_1456,N_1417);
nor U1606 (N_1606,N_1436,N_1445);
and U1607 (N_1607,N_1414,N_1429);
xor U1608 (N_1608,N_1451,N_1454);
nor U1609 (N_1609,N_1455,N_1445);
xnor U1610 (N_1610,N_1454,N_1466);
nor U1611 (N_1611,N_1492,N_1384);
nand U1612 (N_1612,N_1426,N_1395);
nand U1613 (N_1613,N_1378,N_1416);
nor U1614 (N_1614,N_1473,N_1498);
or U1615 (N_1615,N_1492,N_1464);
nor U1616 (N_1616,N_1382,N_1457);
nor U1617 (N_1617,N_1391,N_1491);
xor U1618 (N_1618,N_1418,N_1402);
nor U1619 (N_1619,N_1486,N_1446);
or U1620 (N_1620,N_1419,N_1413);
nand U1621 (N_1621,N_1466,N_1400);
and U1622 (N_1622,N_1457,N_1435);
nor U1623 (N_1623,N_1436,N_1427);
xnor U1624 (N_1624,N_1451,N_1480);
xor U1625 (N_1625,N_1516,N_1604);
and U1626 (N_1626,N_1595,N_1523);
nand U1627 (N_1627,N_1588,N_1501);
nand U1628 (N_1628,N_1589,N_1561);
nand U1629 (N_1629,N_1544,N_1521);
and U1630 (N_1630,N_1616,N_1584);
nor U1631 (N_1631,N_1507,N_1526);
nor U1632 (N_1632,N_1570,N_1509);
and U1633 (N_1633,N_1567,N_1510);
nand U1634 (N_1634,N_1573,N_1527);
nand U1635 (N_1635,N_1624,N_1529);
nor U1636 (N_1636,N_1512,N_1586);
and U1637 (N_1637,N_1543,N_1608);
and U1638 (N_1638,N_1623,N_1505);
and U1639 (N_1639,N_1539,N_1541);
and U1640 (N_1640,N_1576,N_1525);
nor U1641 (N_1641,N_1552,N_1532);
nand U1642 (N_1642,N_1577,N_1592);
nor U1643 (N_1643,N_1599,N_1620);
or U1644 (N_1644,N_1585,N_1538);
and U1645 (N_1645,N_1502,N_1517);
xor U1646 (N_1646,N_1542,N_1563);
and U1647 (N_1647,N_1603,N_1609);
nor U1648 (N_1648,N_1601,N_1550);
nor U1649 (N_1649,N_1515,N_1602);
nand U1650 (N_1650,N_1613,N_1606);
nand U1651 (N_1651,N_1574,N_1607);
nand U1652 (N_1652,N_1564,N_1508);
nand U1653 (N_1653,N_1559,N_1503);
and U1654 (N_1654,N_1571,N_1534);
or U1655 (N_1655,N_1554,N_1513);
or U1656 (N_1656,N_1610,N_1611);
and U1657 (N_1657,N_1518,N_1560);
nor U1658 (N_1658,N_1533,N_1565);
nand U1659 (N_1659,N_1504,N_1583);
xor U1660 (N_1660,N_1617,N_1558);
nand U1661 (N_1661,N_1511,N_1580);
and U1662 (N_1662,N_1528,N_1522);
xnor U1663 (N_1663,N_1596,N_1612);
nand U1664 (N_1664,N_1535,N_1621);
nand U1665 (N_1665,N_1622,N_1591);
or U1666 (N_1666,N_1557,N_1569);
xnor U1667 (N_1667,N_1578,N_1594);
xor U1668 (N_1668,N_1562,N_1587);
xor U1669 (N_1669,N_1566,N_1537);
and U1670 (N_1670,N_1549,N_1545);
nand U1671 (N_1671,N_1520,N_1600);
and U1672 (N_1672,N_1514,N_1579);
or U1673 (N_1673,N_1619,N_1618);
xor U1674 (N_1674,N_1530,N_1575);
and U1675 (N_1675,N_1605,N_1546);
xor U1676 (N_1676,N_1531,N_1555);
nand U1677 (N_1677,N_1614,N_1524);
or U1678 (N_1678,N_1556,N_1536);
nand U1679 (N_1679,N_1582,N_1551);
nor U1680 (N_1680,N_1540,N_1506);
or U1681 (N_1681,N_1568,N_1581);
nor U1682 (N_1682,N_1553,N_1598);
or U1683 (N_1683,N_1593,N_1548);
and U1684 (N_1684,N_1615,N_1500);
nor U1685 (N_1685,N_1590,N_1519);
nand U1686 (N_1686,N_1572,N_1597);
nor U1687 (N_1687,N_1547,N_1581);
xnor U1688 (N_1688,N_1545,N_1560);
nand U1689 (N_1689,N_1621,N_1545);
and U1690 (N_1690,N_1607,N_1593);
nor U1691 (N_1691,N_1510,N_1575);
and U1692 (N_1692,N_1580,N_1602);
or U1693 (N_1693,N_1601,N_1622);
or U1694 (N_1694,N_1501,N_1605);
or U1695 (N_1695,N_1565,N_1613);
and U1696 (N_1696,N_1608,N_1540);
nand U1697 (N_1697,N_1561,N_1595);
nor U1698 (N_1698,N_1536,N_1590);
nand U1699 (N_1699,N_1563,N_1536);
or U1700 (N_1700,N_1545,N_1596);
nor U1701 (N_1701,N_1549,N_1564);
nand U1702 (N_1702,N_1575,N_1590);
xor U1703 (N_1703,N_1547,N_1568);
xor U1704 (N_1704,N_1504,N_1578);
or U1705 (N_1705,N_1600,N_1577);
nand U1706 (N_1706,N_1513,N_1548);
or U1707 (N_1707,N_1501,N_1612);
xor U1708 (N_1708,N_1512,N_1542);
nor U1709 (N_1709,N_1555,N_1521);
nand U1710 (N_1710,N_1583,N_1612);
xnor U1711 (N_1711,N_1624,N_1615);
and U1712 (N_1712,N_1593,N_1544);
nor U1713 (N_1713,N_1605,N_1603);
or U1714 (N_1714,N_1524,N_1577);
nor U1715 (N_1715,N_1593,N_1620);
xor U1716 (N_1716,N_1558,N_1555);
or U1717 (N_1717,N_1608,N_1565);
nor U1718 (N_1718,N_1502,N_1602);
or U1719 (N_1719,N_1624,N_1581);
nand U1720 (N_1720,N_1571,N_1513);
nand U1721 (N_1721,N_1500,N_1531);
nor U1722 (N_1722,N_1554,N_1585);
and U1723 (N_1723,N_1551,N_1549);
nor U1724 (N_1724,N_1542,N_1620);
nand U1725 (N_1725,N_1568,N_1595);
and U1726 (N_1726,N_1567,N_1558);
nand U1727 (N_1727,N_1562,N_1566);
nor U1728 (N_1728,N_1619,N_1588);
or U1729 (N_1729,N_1563,N_1569);
nand U1730 (N_1730,N_1614,N_1576);
or U1731 (N_1731,N_1563,N_1556);
nor U1732 (N_1732,N_1536,N_1611);
nand U1733 (N_1733,N_1610,N_1595);
and U1734 (N_1734,N_1587,N_1585);
nor U1735 (N_1735,N_1597,N_1595);
xnor U1736 (N_1736,N_1597,N_1536);
or U1737 (N_1737,N_1572,N_1613);
nor U1738 (N_1738,N_1554,N_1508);
and U1739 (N_1739,N_1503,N_1500);
nand U1740 (N_1740,N_1566,N_1589);
xor U1741 (N_1741,N_1552,N_1616);
or U1742 (N_1742,N_1554,N_1507);
or U1743 (N_1743,N_1605,N_1512);
xor U1744 (N_1744,N_1594,N_1603);
xnor U1745 (N_1745,N_1608,N_1606);
xnor U1746 (N_1746,N_1515,N_1605);
nand U1747 (N_1747,N_1506,N_1608);
nor U1748 (N_1748,N_1500,N_1607);
or U1749 (N_1749,N_1514,N_1563);
or U1750 (N_1750,N_1641,N_1733);
and U1751 (N_1751,N_1731,N_1643);
or U1752 (N_1752,N_1693,N_1628);
and U1753 (N_1753,N_1721,N_1640);
nor U1754 (N_1754,N_1743,N_1725);
xor U1755 (N_1755,N_1635,N_1708);
or U1756 (N_1756,N_1688,N_1707);
nand U1757 (N_1757,N_1703,N_1726);
and U1758 (N_1758,N_1696,N_1626);
xnor U1759 (N_1759,N_1709,N_1748);
xor U1760 (N_1760,N_1682,N_1702);
and U1761 (N_1761,N_1657,N_1684);
xor U1762 (N_1762,N_1716,N_1712);
xor U1763 (N_1763,N_1711,N_1625);
nand U1764 (N_1764,N_1705,N_1699);
or U1765 (N_1765,N_1692,N_1660);
or U1766 (N_1766,N_1663,N_1737);
and U1767 (N_1767,N_1666,N_1740);
xor U1768 (N_1768,N_1720,N_1686);
or U1769 (N_1769,N_1741,N_1706);
nand U1770 (N_1770,N_1713,N_1632);
and U1771 (N_1771,N_1749,N_1727);
nor U1772 (N_1772,N_1649,N_1656);
or U1773 (N_1773,N_1667,N_1664);
nor U1774 (N_1774,N_1668,N_1665);
or U1775 (N_1775,N_1734,N_1652);
nand U1776 (N_1776,N_1669,N_1655);
and U1777 (N_1777,N_1698,N_1654);
nand U1778 (N_1778,N_1647,N_1627);
or U1779 (N_1779,N_1630,N_1650);
nand U1780 (N_1780,N_1680,N_1633);
or U1781 (N_1781,N_1658,N_1639);
or U1782 (N_1782,N_1746,N_1637);
nand U1783 (N_1783,N_1638,N_1739);
or U1784 (N_1784,N_1644,N_1670);
or U1785 (N_1785,N_1747,N_1697);
xnor U1786 (N_1786,N_1672,N_1719);
and U1787 (N_1787,N_1714,N_1744);
nand U1788 (N_1788,N_1675,N_1673);
and U1789 (N_1789,N_1631,N_1634);
xnor U1790 (N_1790,N_1642,N_1723);
xnor U1791 (N_1791,N_1653,N_1690);
and U1792 (N_1792,N_1645,N_1676);
xnor U1793 (N_1793,N_1636,N_1729);
xor U1794 (N_1794,N_1678,N_1674);
nor U1795 (N_1795,N_1687,N_1700);
nor U1796 (N_1796,N_1671,N_1722);
or U1797 (N_1797,N_1728,N_1718);
and U1798 (N_1798,N_1695,N_1710);
nor U1799 (N_1799,N_1732,N_1691);
nor U1800 (N_1800,N_1679,N_1689);
nand U1801 (N_1801,N_1742,N_1694);
nand U1802 (N_1802,N_1646,N_1704);
and U1803 (N_1803,N_1659,N_1683);
or U1804 (N_1804,N_1715,N_1717);
nand U1805 (N_1805,N_1730,N_1629);
nand U1806 (N_1806,N_1735,N_1681);
and U1807 (N_1807,N_1661,N_1651);
xor U1808 (N_1808,N_1662,N_1685);
and U1809 (N_1809,N_1648,N_1736);
and U1810 (N_1810,N_1701,N_1724);
xor U1811 (N_1811,N_1677,N_1745);
nor U1812 (N_1812,N_1738,N_1646);
nand U1813 (N_1813,N_1740,N_1656);
xnor U1814 (N_1814,N_1670,N_1655);
nor U1815 (N_1815,N_1676,N_1669);
nor U1816 (N_1816,N_1720,N_1732);
xnor U1817 (N_1817,N_1647,N_1742);
nand U1818 (N_1818,N_1645,N_1721);
nand U1819 (N_1819,N_1728,N_1706);
xor U1820 (N_1820,N_1734,N_1730);
nand U1821 (N_1821,N_1696,N_1662);
nand U1822 (N_1822,N_1727,N_1742);
or U1823 (N_1823,N_1729,N_1735);
and U1824 (N_1824,N_1726,N_1739);
or U1825 (N_1825,N_1726,N_1731);
nand U1826 (N_1826,N_1708,N_1732);
nand U1827 (N_1827,N_1700,N_1697);
and U1828 (N_1828,N_1644,N_1689);
or U1829 (N_1829,N_1659,N_1649);
xnor U1830 (N_1830,N_1698,N_1707);
and U1831 (N_1831,N_1700,N_1673);
nand U1832 (N_1832,N_1664,N_1704);
and U1833 (N_1833,N_1678,N_1698);
nand U1834 (N_1834,N_1639,N_1637);
and U1835 (N_1835,N_1686,N_1625);
xor U1836 (N_1836,N_1684,N_1637);
nor U1837 (N_1837,N_1664,N_1693);
nor U1838 (N_1838,N_1686,N_1707);
nor U1839 (N_1839,N_1629,N_1649);
xnor U1840 (N_1840,N_1641,N_1697);
nand U1841 (N_1841,N_1646,N_1749);
nand U1842 (N_1842,N_1720,N_1659);
xor U1843 (N_1843,N_1699,N_1714);
nand U1844 (N_1844,N_1639,N_1741);
xor U1845 (N_1845,N_1727,N_1655);
and U1846 (N_1846,N_1654,N_1630);
nand U1847 (N_1847,N_1654,N_1718);
and U1848 (N_1848,N_1640,N_1683);
xor U1849 (N_1849,N_1674,N_1686);
nand U1850 (N_1850,N_1705,N_1730);
and U1851 (N_1851,N_1671,N_1724);
and U1852 (N_1852,N_1626,N_1682);
or U1853 (N_1853,N_1672,N_1739);
xnor U1854 (N_1854,N_1674,N_1639);
nor U1855 (N_1855,N_1636,N_1675);
or U1856 (N_1856,N_1688,N_1637);
nand U1857 (N_1857,N_1740,N_1660);
or U1858 (N_1858,N_1684,N_1626);
or U1859 (N_1859,N_1684,N_1687);
nand U1860 (N_1860,N_1636,N_1655);
nor U1861 (N_1861,N_1681,N_1651);
nor U1862 (N_1862,N_1655,N_1672);
nand U1863 (N_1863,N_1637,N_1647);
xor U1864 (N_1864,N_1664,N_1748);
or U1865 (N_1865,N_1625,N_1673);
and U1866 (N_1866,N_1657,N_1649);
nand U1867 (N_1867,N_1738,N_1713);
and U1868 (N_1868,N_1685,N_1705);
xnor U1869 (N_1869,N_1749,N_1668);
nor U1870 (N_1870,N_1663,N_1635);
xnor U1871 (N_1871,N_1745,N_1681);
or U1872 (N_1872,N_1692,N_1702);
nor U1873 (N_1873,N_1659,N_1721);
and U1874 (N_1874,N_1702,N_1722);
and U1875 (N_1875,N_1839,N_1760);
xor U1876 (N_1876,N_1802,N_1849);
nor U1877 (N_1877,N_1751,N_1775);
or U1878 (N_1878,N_1830,N_1753);
nand U1879 (N_1879,N_1829,N_1758);
nor U1880 (N_1880,N_1812,N_1784);
nand U1881 (N_1881,N_1823,N_1864);
nor U1882 (N_1882,N_1790,N_1773);
nor U1883 (N_1883,N_1863,N_1844);
xnor U1884 (N_1884,N_1789,N_1845);
nand U1885 (N_1885,N_1800,N_1759);
nand U1886 (N_1886,N_1810,N_1873);
xor U1887 (N_1887,N_1815,N_1861);
nor U1888 (N_1888,N_1846,N_1862);
nor U1889 (N_1889,N_1872,N_1827);
nor U1890 (N_1890,N_1824,N_1836);
and U1891 (N_1891,N_1762,N_1848);
and U1892 (N_1892,N_1780,N_1787);
xor U1893 (N_1893,N_1786,N_1799);
nand U1894 (N_1894,N_1806,N_1819);
and U1895 (N_1895,N_1811,N_1779);
and U1896 (N_1896,N_1854,N_1757);
nor U1897 (N_1897,N_1756,N_1852);
nor U1898 (N_1898,N_1826,N_1755);
nor U1899 (N_1899,N_1754,N_1814);
xor U1900 (N_1900,N_1870,N_1809);
or U1901 (N_1901,N_1788,N_1769);
xor U1902 (N_1902,N_1791,N_1856);
nand U1903 (N_1903,N_1767,N_1794);
nand U1904 (N_1904,N_1752,N_1853);
xnor U1905 (N_1905,N_1792,N_1813);
nor U1906 (N_1906,N_1777,N_1785);
nor U1907 (N_1907,N_1774,N_1803);
or U1908 (N_1908,N_1764,N_1866);
nand U1909 (N_1909,N_1822,N_1765);
nor U1910 (N_1910,N_1797,N_1818);
nand U1911 (N_1911,N_1763,N_1772);
and U1912 (N_1912,N_1842,N_1857);
or U1913 (N_1913,N_1835,N_1874);
nand U1914 (N_1914,N_1801,N_1778);
nand U1915 (N_1915,N_1796,N_1770);
xnor U1916 (N_1916,N_1871,N_1867);
or U1917 (N_1917,N_1865,N_1795);
nor U1918 (N_1918,N_1869,N_1847);
or U1919 (N_1919,N_1821,N_1805);
xnor U1920 (N_1920,N_1838,N_1776);
nor U1921 (N_1921,N_1816,N_1840);
xor U1922 (N_1922,N_1860,N_1793);
nor U1923 (N_1923,N_1837,N_1771);
or U1924 (N_1924,N_1868,N_1833);
nor U1925 (N_1925,N_1831,N_1851);
nor U1926 (N_1926,N_1781,N_1783);
or U1927 (N_1927,N_1828,N_1804);
xnor U1928 (N_1928,N_1798,N_1766);
nor U1929 (N_1929,N_1782,N_1843);
nor U1930 (N_1930,N_1859,N_1808);
nor U1931 (N_1931,N_1761,N_1768);
nor U1932 (N_1932,N_1858,N_1850);
nor U1933 (N_1933,N_1807,N_1825);
nor U1934 (N_1934,N_1750,N_1817);
and U1935 (N_1935,N_1841,N_1855);
or U1936 (N_1936,N_1834,N_1820);
or U1937 (N_1937,N_1832,N_1869);
nor U1938 (N_1938,N_1806,N_1874);
or U1939 (N_1939,N_1817,N_1814);
nand U1940 (N_1940,N_1830,N_1835);
xor U1941 (N_1941,N_1832,N_1841);
xnor U1942 (N_1942,N_1862,N_1768);
or U1943 (N_1943,N_1811,N_1842);
and U1944 (N_1944,N_1854,N_1787);
or U1945 (N_1945,N_1790,N_1800);
xor U1946 (N_1946,N_1766,N_1799);
xor U1947 (N_1947,N_1793,N_1813);
and U1948 (N_1948,N_1858,N_1801);
or U1949 (N_1949,N_1760,N_1859);
nor U1950 (N_1950,N_1759,N_1853);
nand U1951 (N_1951,N_1841,N_1871);
or U1952 (N_1952,N_1817,N_1765);
or U1953 (N_1953,N_1803,N_1770);
nand U1954 (N_1954,N_1800,N_1813);
or U1955 (N_1955,N_1794,N_1783);
or U1956 (N_1956,N_1758,N_1811);
xnor U1957 (N_1957,N_1794,N_1852);
and U1958 (N_1958,N_1764,N_1792);
nand U1959 (N_1959,N_1826,N_1773);
nand U1960 (N_1960,N_1753,N_1758);
or U1961 (N_1961,N_1762,N_1808);
and U1962 (N_1962,N_1772,N_1869);
or U1963 (N_1963,N_1807,N_1828);
and U1964 (N_1964,N_1786,N_1835);
and U1965 (N_1965,N_1753,N_1834);
nor U1966 (N_1966,N_1769,N_1789);
xor U1967 (N_1967,N_1864,N_1798);
or U1968 (N_1968,N_1813,N_1762);
xor U1969 (N_1969,N_1753,N_1851);
nand U1970 (N_1970,N_1756,N_1812);
or U1971 (N_1971,N_1866,N_1771);
and U1972 (N_1972,N_1791,N_1873);
nand U1973 (N_1973,N_1866,N_1775);
and U1974 (N_1974,N_1783,N_1773);
nand U1975 (N_1975,N_1856,N_1841);
xor U1976 (N_1976,N_1781,N_1755);
nand U1977 (N_1977,N_1824,N_1858);
nor U1978 (N_1978,N_1839,N_1854);
and U1979 (N_1979,N_1812,N_1846);
xor U1980 (N_1980,N_1856,N_1818);
nor U1981 (N_1981,N_1804,N_1856);
xnor U1982 (N_1982,N_1771,N_1756);
and U1983 (N_1983,N_1822,N_1795);
nor U1984 (N_1984,N_1805,N_1840);
or U1985 (N_1985,N_1793,N_1836);
or U1986 (N_1986,N_1840,N_1844);
xnor U1987 (N_1987,N_1834,N_1762);
nor U1988 (N_1988,N_1763,N_1843);
or U1989 (N_1989,N_1752,N_1834);
and U1990 (N_1990,N_1781,N_1803);
nand U1991 (N_1991,N_1822,N_1771);
xor U1992 (N_1992,N_1820,N_1784);
xnor U1993 (N_1993,N_1770,N_1860);
xor U1994 (N_1994,N_1861,N_1867);
nor U1995 (N_1995,N_1816,N_1866);
xnor U1996 (N_1996,N_1772,N_1821);
and U1997 (N_1997,N_1760,N_1852);
or U1998 (N_1998,N_1855,N_1787);
or U1999 (N_1999,N_1795,N_1833);
nand U2000 (N_2000,N_1950,N_1889);
or U2001 (N_2001,N_1948,N_1936);
and U2002 (N_2002,N_1941,N_1896);
or U2003 (N_2003,N_1980,N_1903);
and U2004 (N_2004,N_1892,N_1884);
xnor U2005 (N_2005,N_1931,N_1909);
or U2006 (N_2006,N_1891,N_1984);
and U2007 (N_2007,N_1910,N_1929);
or U2008 (N_2008,N_1912,N_1901);
nand U2009 (N_2009,N_1922,N_1881);
nor U2010 (N_2010,N_1930,N_1888);
and U2011 (N_2011,N_1998,N_1959);
or U2012 (N_2012,N_1895,N_1900);
nand U2013 (N_2013,N_1978,N_1920);
and U2014 (N_2014,N_1887,N_1951);
and U2015 (N_2015,N_1878,N_1907);
and U2016 (N_2016,N_1994,N_1995);
xnor U2017 (N_2017,N_1971,N_1992);
or U2018 (N_2018,N_1924,N_1964);
and U2019 (N_2019,N_1976,N_1933);
and U2020 (N_2020,N_1989,N_1905);
xor U2021 (N_2021,N_1990,N_1897);
xor U2022 (N_2022,N_1882,N_1885);
nand U2023 (N_2023,N_1915,N_1916);
nor U2024 (N_2024,N_1982,N_1952);
nand U2025 (N_2025,N_1974,N_1925);
or U2026 (N_2026,N_1939,N_1906);
nand U2027 (N_2027,N_1957,N_1945);
nand U2028 (N_2028,N_1960,N_1965);
nand U2029 (N_2029,N_1926,N_1918);
nand U2030 (N_2030,N_1899,N_1911);
xor U2031 (N_2031,N_1968,N_1997);
nand U2032 (N_2032,N_1908,N_1988);
nor U2033 (N_2033,N_1983,N_1953);
nand U2034 (N_2034,N_1880,N_1877);
nand U2035 (N_2035,N_1967,N_1993);
nor U2036 (N_2036,N_1913,N_1928);
xor U2037 (N_2037,N_1919,N_1966);
nand U2038 (N_2038,N_1956,N_1955);
and U2039 (N_2039,N_1927,N_1962);
nor U2040 (N_2040,N_1876,N_1975);
and U2041 (N_2041,N_1954,N_1923);
and U2042 (N_2042,N_1981,N_1999);
nor U2043 (N_2043,N_1985,N_1875);
nor U2044 (N_2044,N_1943,N_1977);
nor U2045 (N_2045,N_1946,N_1944);
nor U2046 (N_2046,N_1883,N_1917);
xor U2047 (N_2047,N_1938,N_1898);
nor U2048 (N_2048,N_1942,N_1996);
nor U2049 (N_2049,N_1932,N_1902);
and U2050 (N_2050,N_1979,N_1961);
nand U2051 (N_2051,N_1940,N_1886);
or U2052 (N_2052,N_1935,N_1963);
nor U2053 (N_2053,N_1969,N_1986);
and U2054 (N_2054,N_1921,N_1893);
nand U2055 (N_2055,N_1991,N_1973);
or U2056 (N_2056,N_1879,N_1890);
xor U2057 (N_2057,N_1949,N_1904);
or U2058 (N_2058,N_1894,N_1937);
nor U2059 (N_2059,N_1914,N_1972);
nand U2060 (N_2060,N_1947,N_1987);
xnor U2061 (N_2061,N_1934,N_1970);
nand U2062 (N_2062,N_1958,N_1993);
nor U2063 (N_2063,N_1986,N_1999);
and U2064 (N_2064,N_1923,N_1922);
and U2065 (N_2065,N_1954,N_1926);
nor U2066 (N_2066,N_1927,N_1966);
xor U2067 (N_2067,N_1990,N_1886);
nor U2068 (N_2068,N_1877,N_1973);
nor U2069 (N_2069,N_1994,N_1959);
nor U2070 (N_2070,N_1969,N_1984);
nor U2071 (N_2071,N_1993,N_1989);
xor U2072 (N_2072,N_1965,N_1879);
nor U2073 (N_2073,N_1896,N_1906);
and U2074 (N_2074,N_1974,N_1880);
nand U2075 (N_2075,N_1987,N_1967);
xnor U2076 (N_2076,N_1935,N_1953);
or U2077 (N_2077,N_1914,N_1879);
nor U2078 (N_2078,N_1927,N_1878);
or U2079 (N_2079,N_1921,N_1931);
or U2080 (N_2080,N_1964,N_1911);
nor U2081 (N_2081,N_1943,N_1965);
nor U2082 (N_2082,N_1887,N_1997);
nand U2083 (N_2083,N_1885,N_1939);
xnor U2084 (N_2084,N_1901,N_1944);
xnor U2085 (N_2085,N_1899,N_1940);
or U2086 (N_2086,N_1887,N_1993);
nor U2087 (N_2087,N_1945,N_1915);
nor U2088 (N_2088,N_1893,N_1930);
nand U2089 (N_2089,N_1899,N_1881);
nor U2090 (N_2090,N_1890,N_1898);
xnor U2091 (N_2091,N_1907,N_1987);
nand U2092 (N_2092,N_1898,N_1948);
or U2093 (N_2093,N_1905,N_1888);
xor U2094 (N_2094,N_1967,N_1966);
xnor U2095 (N_2095,N_1891,N_1922);
xnor U2096 (N_2096,N_1994,N_1934);
nand U2097 (N_2097,N_1945,N_1993);
nand U2098 (N_2098,N_1881,N_1977);
xnor U2099 (N_2099,N_1897,N_1887);
nor U2100 (N_2100,N_1937,N_1985);
xor U2101 (N_2101,N_1964,N_1892);
and U2102 (N_2102,N_1951,N_1891);
xor U2103 (N_2103,N_1944,N_1964);
or U2104 (N_2104,N_1985,N_1876);
xor U2105 (N_2105,N_1883,N_1947);
nand U2106 (N_2106,N_1945,N_1907);
nand U2107 (N_2107,N_1901,N_1986);
or U2108 (N_2108,N_1929,N_1896);
nand U2109 (N_2109,N_1984,N_1941);
and U2110 (N_2110,N_1932,N_1929);
and U2111 (N_2111,N_1955,N_1996);
or U2112 (N_2112,N_1968,N_1885);
nand U2113 (N_2113,N_1953,N_1987);
xnor U2114 (N_2114,N_1913,N_1948);
nor U2115 (N_2115,N_1994,N_1896);
xnor U2116 (N_2116,N_1914,N_1993);
nand U2117 (N_2117,N_1990,N_1969);
and U2118 (N_2118,N_1880,N_1991);
xor U2119 (N_2119,N_1905,N_1953);
or U2120 (N_2120,N_1991,N_1923);
nor U2121 (N_2121,N_1893,N_1925);
and U2122 (N_2122,N_1912,N_1930);
nor U2123 (N_2123,N_1958,N_1884);
xnor U2124 (N_2124,N_1902,N_1963);
and U2125 (N_2125,N_2049,N_2010);
nand U2126 (N_2126,N_2120,N_2089);
and U2127 (N_2127,N_2035,N_2013);
or U2128 (N_2128,N_2090,N_2063);
nor U2129 (N_2129,N_2041,N_2042);
or U2130 (N_2130,N_2018,N_2102);
nand U2131 (N_2131,N_2060,N_2012);
and U2132 (N_2132,N_2074,N_2119);
or U2133 (N_2133,N_2075,N_2053);
xor U2134 (N_2134,N_2083,N_2023);
or U2135 (N_2135,N_2122,N_2043);
xor U2136 (N_2136,N_2028,N_2069);
or U2137 (N_2137,N_2052,N_2124);
xnor U2138 (N_2138,N_2088,N_2025);
xor U2139 (N_2139,N_2026,N_2007);
and U2140 (N_2140,N_2044,N_2115);
xnor U2141 (N_2141,N_2011,N_2095);
xor U2142 (N_2142,N_2117,N_2091);
nand U2143 (N_2143,N_2070,N_2033);
nand U2144 (N_2144,N_2019,N_2098);
xnor U2145 (N_2145,N_2045,N_2108);
nand U2146 (N_2146,N_2058,N_2066);
or U2147 (N_2147,N_2077,N_2079);
nand U2148 (N_2148,N_2014,N_2032);
or U2149 (N_2149,N_2085,N_2104);
or U2150 (N_2150,N_2123,N_2038);
nor U2151 (N_2151,N_2051,N_2116);
and U2152 (N_2152,N_2110,N_2103);
or U2153 (N_2153,N_2111,N_2109);
xor U2154 (N_2154,N_2029,N_2105);
xnor U2155 (N_2155,N_2073,N_2002);
nor U2156 (N_2156,N_2087,N_2068);
xor U2157 (N_2157,N_2027,N_2024);
nand U2158 (N_2158,N_2016,N_2076);
nor U2159 (N_2159,N_2061,N_2001);
or U2160 (N_2160,N_2004,N_2112);
and U2161 (N_2161,N_2006,N_2071);
and U2162 (N_2162,N_2021,N_2009);
nand U2163 (N_2163,N_2086,N_2000);
nor U2164 (N_2164,N_2022,N_2106);
nor U2165 (N_2165,N_2017,N_2101);
or U2166 (N_2166,N_2055,N_2118);
nor U2167 (N_2167,N_2100,N_2081);
or U2168 (N_2168,N_2097,N_2005);
nand U2169 (N_2169,N_2113,N_2046);
nand U2170 (N_2170,N_2080,N_2031);
nand U2171 (N_2171,N_2003,N_2047);
nor U2172 (N_2172,N_2093,N_2057);
nor U2173 (N_2173,N_2114,N_2099);
or U2174 (N_2174,N_2067,N_2020);
and U2175 (N_2175,N_2050,N_2082);
and U2176 (N_2176,N_2092,N_2030);
and U2177 (N_2177,N_2008,N_2062);
nand U2178 (N_2178,N_2054,N_2094);
or U2179 (N_2179,N_2072,N_2121);
nand U2180 (N_2180,N_2048,N_2036);
and U2181 (N_2181,N_2040,N_2064);
and U2182 (N_2182,N_2059,N_2065);
xnor U2183 (N_2183,N_2078,N_2107);
nand U2184 (N_2184,N_2096,N_2037);
or U2185 (N_2185,N_2039,N_2015);
nor U2186 (N_2186,N_2084,N_2056);
nor U2187 (N_2187,N_2034,N_2109);
xnor U2188 (N_2188,N_2123,N_2041);
nand U2189 (N_2189,N_2070,N_2016);
and U2190 (N_2190,N_2107,N_2091);
nor U2191 (N_2191,N_2055,N_2008);
or U2192 (N_2192,N_2062,N_2002);
and U2193 (N_2193,N_2109,N_2027);
nor U2194 (N_2194,N_2081,N_2011);
xor U2195 (N_2195,N_2118,N_2124);
nor U2196 (N_2196,N_2023,N_2033);
nor U2197 (N_2197,N_2000,N_2066);
nand U2198 (N_2198,N_2012,N_2071);
nand U2199 (N_2199,N_2022,N_2123);
nand U2200 (N_2200,N_2083,N_2057);
and U2201 (N_2201,N_2018,N_2009);
and U2202 (N_2202,N_2043,N_2050);
or U2203 (N_2203,N_2079,N_2035);
nand U2204 (N_2204,N_2092,N_2088);
nor U2205 (N_2205,N_2068,N_2065);
nand U2206 (N_2206,N_2020,N_2115);
or U2207 (N_2207,N_2073,N_2017);
and U2208 (N_2208,N_2006,N_2020);
nor U2209 (N_2209,N_2092,N_2051);
or U2210 (N_2210,N_2035,N_2055);
nor U2211 (N_2211,N_2072,N_2053);
xor U2212 (N_2212,N_2001,N_2033);
xor U2213 (N_2213,N_2005,N_2001);
and U2214 (N_2214,N_2031,N_2103);
and U2215 (N_2215,N_2097,N_2007);
and U2216 (N_2216,N_2046,N_2064);
and U2217 (N_2217,N_2079,N_2113);
or U2218 (N_2218,N_2032,N_2068);
or U2219 (N_2219,N_2084,N_2075);
or U2220 (N_2220,N_2075,N_2089);
and U2221 (N_2221,N_2041,N_2048);
and U2222 (N_2222,N_2114,N_2086);
nor U2223 (N_2223,N_2043,N_2083);
and U2224 (N_2224,N_2000,N_2118);
nand U2225 (N_2225,N_2059,N_2082);
nand U2226 (N_2226,N_2082,N_2028);
nand U2227 (N_2227,N_2109,N_2088);
nor U2228 (N_2228,N_2048,N_2057);
xnor U2229 (N_2229,N_2027,N_2107);
or U2230 (N_2230,N_2006,N_2044);
nand U2231 (N_2231,N_2010,N_2015);
or U2232 (N_2232,N_2097,N_2045);
xnor U2233 (N_2233,N_2006,N_2021);
nand U2234 (N_2234,N_2085,N_2103);
nor U2235 (N_2235,N_2073,N_2041);
nor U2236 (N_2236,N_2075,N_2114);
nand U2237 (N_2237,N_2067,N_2022);
nand U2238 (N_2238,N_2099,N_2030);
xnor U2239 (N_2239,N_2045,N_2081);
xnor U2240 (N_2240,N_2062,N_2095);
or U2241 (N_2241,N_2050,N_2080);
and U2242 (N_2242,N_2097,N_2003);
or U2243 (N_2243,N_2071,N_2016);
xor U2244 (N_2244,N_2083,N_2025);
xnor U2245 (N_2245,N_2023,N_2124);
or U2246 (N_2246,N_2080,N_2003);
and U2247 (N_2247,N_2092,N_2109);
nor U2248 (N_2248,N_2013,N_2062);
nor U2249 (N_2249,N_2090,N_2040);
xnor U2250 (N_2250,N_2197,N_2166);
and U2251 (N_2251,N_2228,N_2208);
xnor U2252 (N_2252,N_2209,N_2161);
xor U2253 (N_2253,N_2183,N_2226);
xor U2254 (N_2254,N_2225,N_2221);
nor U2255 (N_2255,N_2187,N_2165);
and U2256 (N_2256,N_2206,N_2235);
and U2257 (N_2257,N_2142,N_2134);
nand U2258 (N_2258,N_2216,N_2178);
nor U2259 (N_2259,N_2131,N_2169);
xor U2260 (N_2260,N_2143,N_2170);
and U2261 (N_2261,N_2214,N_2229);
nand U2262 (N_2262,N_2151,N_2147);
or U2263 (N_2263,N_2173,N_2158);
xor U2264 (N_2264,N_2210,N_2141);
nor U2265 (N_2265,N_2242,N_2185);
nor U2266 (N_2266,N_2247,N_2241);
and U2267 (N_2267,N_2144,N_2138);
nand U2268 (N_2268,N_2139,N_2159);
nand U2269 (N_2269,N_2237,N_2201);
and U2270 (N_2270,N_2204,N_2203);
and U2271 (N_2271,N_2233,N_2163);
nor U2272 (N_2272,N_2150,N_2231);
xnor U2273 (N_2273,N_2156,N_2130);
or U2274 (N_2274,N_2227,N_2194);
nor U2275 (N_2275,N_2249,N_2145);
xor U2276 (N_2276,N_2244,N_2192);
and U2277 (N_2277,N_2193,N_2167);
and U2278 (N_2278,N_2177,N_2219);
and U2279 (N_2279,N_2196,N_2190);
and U2280 (N_2280,N_2146,N_2129);
nor U2281 (N_2281,N_2205,N_2184);
and U2282 (N_2282,N_2245,N_2236);
nand U2283 (N_2283,N_2176,N_2174);
and U2284 (N_2284,N_2137,N_2238);
or U2285 (N_2285,N_2148,N_2195);
nor U2286 (N_2286,N_2202,N_2180);
and U2287 (N_2287,N_2135,N_2200);
or U2288 (N_2288,N_2136,N_2188);
nand U2289 (N_2289,N_2160,N_2127);
xor U2290 (N_2290,N_2125,N_2155);
xnor U2291 (N_2291,N_2199,N_2181);
nor U2292 (N_2292,N_2153,N_2179);
or U2293 (N_2293,N_2223,N_2232);
nor U2294 (N_2294,N_2217,N_2152);
xnor U2295 (N_2295,N_2246,N_2191);
or U2296 (N_2296,N_2230,N_2149);
nor U2297 (N_2297,N_2218,N_2224);
and U2298 (N_2298,N_2126,N_2207);
or U2299 (N_2299,N_2171,N_2212);
or U2300 (N_2300,N_2162,N_2186);
nand U2301 (N_2301,N_2240,N_2243);
nand U2302 (N_2302,N_2222,N_2198);
nand U2303 (N_2303,N_2211,N_2128);
and U2304 (N_2304,N_2234,N_2175);
nand U2305 (N_2305,N_2140,N_2168);
and U2306 (N_2306,N_2215,N_2154);
nand U2307 (N_2307,N_2157,N_2248);
and U2308 (N_2308,N_2189,N_2133);
xor U2309 (N_2309,N_2239,N_2220);
nand U2310 (N_2310,N_2164,N_2172);
nand U2311 (N_2311,N_2132,N_2182);
nor U2312 (N_2312,N_2213,N_2214);
and U2313 (N_2313,N_2150,N_2140);
xor U2314 (N_2314,N_2185,N_2201);
nand U2315 (N_2315,N_2178,N_2245);
xnor U2316 (N_2316,N_2204,N_2150);
nor U2317 (N_2317,N_2129,N_2128);
xnor U2318 (N_2318,N_2140,N_2249);
or U2319 (N_2319,N_2219,N_2240);
nand U2320 (N_2320,N_2140,N_2217);
and U2321 (N_2321,N_2196,N_2180);
nand U2322 (N_2322,N_2218,N_2225);
or U2323 (N_2323,N_2144,N_2196);
nand U2324 (N_2324,N_2135,N_2182);
nor U2325 (N_2325,N_2145,N_2156);
and U2326 (N_2326,N_2236,N_2151);
and U2327 (N_2327,N_2190,N_2240);
nor U2328 (N_2328,N_2238,N_2193);
or U2329 (N_2329,N_2146,N_2184);
nor U2330 (N_2330,N_2229,N_2217);
and U2331 (N_2331,N_2231,N_2226);
or U2332 (N_2332,N_2216,N_2221);
xor U2333 (N_2333,N_2125,N_2231);
or U2334 (N_2334,N_2210,N_2231);
or U2335 (N_2335,N_2181,N_2174);
nor U2336 (N_2336,N_2163,N_2185);
or U2337 (N_2337,N_2234,N_2176);
nor U2338 (N_2338,N_2125,N_2194);
nand U2339 (N_2339,N_2208,N_2151);
nand U2340 (N_2340,N_2141,N_2228);
nand U2341 (N_2341,N_2190,N_2247);
or U2342 (N_2342,N_2132,N_2175);
nor U2343 (N_2343,N_2221,N_2193);
xnor U2344 (N_2344,N_2213,N_2196);
or U2345 (N_2345,N_2183,N_2150);
nand U2346 (N_2346,N_2225,N_2172);
and U2347 (N_2347,N_2163,N_2179);
xnor U2348 (N_2348,N_2222,N_2152);
nand U2349 (N_2349,N_2213,N_2181);
nand U2350 (N_2350,N_2225,N_2191);
xnor U2351 (N_2351,N_2238,N_2135);
nand U2352 (N_2352,N_2158,N_2161);
or U2353 (N_2353,N_2183,N_2161);
nor U2354 (N_2354,N_2129,N_2162);
or U2355 (N_2355,N_2143,N_2216);
xnor U2356 (N_2356,N_2156,N_2133);
or U2357 (N_2357,N_2212,N_2165);
and U2358 (N_2358,N_2177,N_2125);
nor U2359 (N_2359,N_2143,N_2217);
xor U2360 (N_2360,N_2171,N_2241);
or U2361 (N_2361,N_2194,N_2191);
nor U2362 (N_2362,N_2230,N_2187);
and U2363 (N_2363,N_2179,N_2144);
or U2364 (N_2364,N_2219,N_2195);
and U2365 (N_2365,N_2148,N_2184);
nand U2366 (N_2366,N_2133,N_2231);
nor U2367 (N_2367,N_2235,N_2201);
nor U2368 (N_2368,N_2171,N_2180);
nand U2369 (N_2369,N_2217,N_2246);
or U2370 (N_2370,N_2228,N_2130);
and U2371 (N_2371,N_2224,N_2134);
and U2372 (N_2372,N_2189,N_2229);
nor U2373 (N_2373,N_2181,N_2214);
nor U2374 (N_2374,N_2218,N_2214);
xnor U2375 (N_2375,N_2264,N_2297);
nand U2376 (N_2376,N_2274,N_2366);
or U2377 (N_2377,N_2273,N_2277);
nor U2378 (N_2378,N_2279,N_2353);
or U2379 (N_2379,N_2299,N_2369);
nand U2380 (N_2380,N_2271,N_2269);
nand U2381 (N_2381,N_2255,N_2260);
and U2382 (N_2382,N_2372,N_2275);
or U2383 (N_2383,N_2365,N_2310);
xnor U2384 (N_2384,N_2252,N_2312);
nor U2385 (N_2385,N_2281,N_2316);
nand U2386 (N_2386,N_2250,N_2280);
or U2387 (N_2387,N_2315,N_2323);
nor U2388 (N_2388,N_2278,N_2289);
and U2389 (N_2389,N_2295,N_2256);
xor U2390 (N_2390,N_2346,N_2347);
nand U2391 (N_2391,N_2322,N_2341);
xnor U2392 (N_2392,N_2263,N_2298);
or U2393 (N_2393,N_2304,N_2259);
nand U2394 (N_2394,N_2305,N_2272);
xnor U2395 (N_2395,N_2370,N_2330);
nor U2396 (N_2396,N_2267,N_2368);
or U2397 (N_2397,N_2268,N_2261);
nand U2398 (N_2398,N_2287,N_2284);
or U2399 (N_2399,N_2342,N_2296);
xor U2400 (N_2400,N_2350,N_2321);
nand U2401 (N_2401,N_2282,N_2328);
xnor U2402 (N_2402,N_2340,N_2336);
and U2403 (N_2403,N_2292,N_2302);
xnor U2404 (N_2404,N_2334,N_2358);
and U2405 (N_2405,N_2300,N_2363);
or U2406 (N_2406,N_2327,N_2262);
nand U2407 (N_2407,N_2331,N_2355);
xnor U2408 (N_2408,N_2301,N_2337);
nor U2409 (N_2409,N_2319,N_2254);
xnor U2410 (N_2410,N_2345,N_2360);
and U2411 (N_2411,N_2314,N_2326);
and U2412 (N_2412,N_2324,N_2276);
and U2413 (N_2413,N_2352,N_2339);
xor U2414 (N_2414,N_2335,N_2351);
nand U2415 (N_2415,N_2343,N_2313);
xor U2416 (N_2416,N_2303,N_2359);
or U2417 (N_2417,N_2371,N_2290);
nor U2418 (N_2418,N_2318,N_2257);
nand U2419 (N_2419,N_2286,N_2332);
xnor U2420 (N_2420,N_2291,N_2348);
xor U2421 (N_2421,N_2333,N_2306);
xor U2422 (N_2422,N_2288,N_2349);
nand U2423 (N_2423,N_2356,N_2307);
xor U2424 (N_2424,N_2317,N_2367);
nand U2425 (N_2425,N_2374,N_2357);
xnor U2426 (N_2426,N_2362,N_2265);
and U2427 (N_2427,N_2270,N_2338);
or U2428 (N_2428,N_2251,N_2294);
and U2429 (N_2429,N_2293,N_2253);
or U2430 (N_2430,N_2308,N_2325);
or U2431 (N_2431,N_2309,N_2329);
or U2432 (N_2432,N_2266,N_2354);
xnor U2433 (N_2433,N_2283,N_2285);
nor U2434 (N_2434,N_2373,N_2364);
nand U2435 (N_2435,N_2361,N_2320);
and U2436 (N_2436,N_2344,N_2258);
or U2437 (N_2437,N_2311,N_2250);
nor U2438 (N_2438,N_2262,N_2337);
or U2439 (N_2439,N_2342,N_2310);
xnor U2440 (N_2440,N_2290,N_2306);
or U2441 (N_2441,N_2355,N_2291);
nand U2442 (N_2442,N_2314,N_2255);
nor U2443 (N_2443,N_2335,N_2310);
or U2444 (N_2444,N_2343,N_2289);
and U2445 (N_2445,N_2363,N_2293);
and U2446 (N_2446,N_2272,N_2329);
or U2447 (N_2447,N_2324,N_2344);
and U2448 (N_2448,N_2262,N_2261);
nor U2449 (N_2449,N_2268,N_2373);
nor U2450 (N_2450,N_2359,N_2344);
nand U2451 (N_2451,N_2323,N_2310);
nor U2452 (N_2452,N_2364,N_2280);
nor U2453 (N_2453,N_2331,N_2338);
and U2454 (N_2454,N_2354,N_2294);
nand U2455 (N_2455,N_2294,N_2290);
xor U2456 (N_2456,N_2356,N_2250);
and U2457 (N_2457,N_2347,N_2261);
nand U2458 (N_2458,N_2291,N_2332);
and U2459 (N_2459,N_2359,N_2277);
or U2460 (N_2460,N_2290,N_2295);
nand U2461 (N_2461,N_2309,N_2317);
and U2462 (N_2462,N_2278,N_2292);
or U2463 (N_2463,N_2289,N_2354);
nor U2464 (N_2464,N_2296,N_2251);
or U2465 (N_2465,N_2290,N_2289);
or U2466 (N_2466,N_2371,N_2364);
and U2467 (N_2467,N_2373,N_2336);
xor U2468 (N_2468,N_2298,N_2330);
nand U2469 (N_2469,N_2348,N_2320);
nand U2470 (N_2470,N_2313,N_2282);
or U2471 (N_2471,N_2279,N_2339);
nand U2472 (N_2472,N_2357,N_2349);
nor U2473 (N_2473,N_2271,N_2261);
nor U2474 (N_2474,N_2272,N_2256);
xor U2475 (N_2475,N_2313,N_2271);
or U2476 (N_2476,N_2311,N_2274);
xor U2477 (N_2477,N_2328,N_2252);
nand U2478 (N_2478,N_2315,N_2256);
nand U2479 (N_2479,N_2363,N_2279);
nand U2480 (N_2480,N_2282,N_2307);
and U2481 (N_2481,N_2292,N_2341);
and U2482 (N_2482,N_2318,N_2294);
nor U2483 (N_2483,N_2290,N_2370);
nand U2484 (N_2484,N_2302,N_2275);
xor U2485 (N_2485,N_2373,N_2368);
and U2486 (N_2486,N_2371,N_2299);
xnor U2487 (N_2487,N_2374,N_2293);
xor U2488 (N_2488,N_2309,N_2369);
or U2489 (N_2489,N_2253,N_2318);
xor U2490 (N_2490,N_2329,N_2353);
nand U2491 (N_2491,N_2327,N_2311);
nor U2492 (N_2492,N_2362,N_2252);
nand U2493 (N_2493,N_2341,N_2333);
xnor U2494 (N_2494,N_2278,N_2270);
nor U2495 (N_2495,N_2345,N_2274);
and U2496 (N_2496,N_2311,N_2336);
nor U2497 (N_2497,N_2308,N_2290);
nor U2498 (N_2498,N_2352,N_2322);
and U2499 (N_2499,N_2368,N_2265);
nand U2500 (N_2500,N_2404,N_2469);
nor U2501 (N_2501,N_2452,N_2409);
xnor U2502 (N_2502,N_2397,N_2418);
nand U2503 (N_2503,N_2447,N_2480);
nand U2504 (N_2504,N_2382,N_2392);
xor U2505 (N_2505,N_2462,N_2408);
or U2506 (N_2506,N_2431,N_2394);
nand U2507 (N_2507,N_2490,N_2437);
nand U2508 (N_2508,N_2495,N_2391);
and U2509 (N_2509,N_2375,N_2470);
nand U2510 (N_2510,N_2402,N_2428);
and U2511 (N_2511,N_2379,N_2396);
and U2512 (N_2512,N_2411,N_2453);
nor U2513 (N_2513,N_2487,N_2460);
or U2514 (N_2514,N_2496,N_2421);
nor U2515 (N_2515,N_2483,N_2430);
and U2516 (N_2516,N_2491,N_2414);
nor U2517 (N_2517,N_2486,N_2420);
or U2518 (N_2518,N_2429,N_2489);
nand U2519 (N_2519,N_2376,N_2381);
or U2520 (N_2520,N_2450,N_2398);
nand U2521 (N_2521,N_2434,N_2454);
nand U2522 (N_2522,N_2481,N_2467);
and U2523 (N_2523,N_2444,N_2406);
and U2524 (N_2524,N_2390,N_2493);
nor U2525 (N_2525,N_2426,N_2463);
xnor U2526 (N_2526,N_2488,N_2464);
nand U2527 (N_2527,N_2419,N_2427);
nor U2528 (N_2528,N_2446,N_2477);
xnor U2529 (N_2529,N_2494,N_2461);
and U2530 (N_2530,N_2478,N_2433);
or U2531 (N_2531,N_2442,N_2498);
xnor U2532 (N_2532,N_2425,N_2466);
nor U2533 (N_2533,N_2378,N_2474);
xnor U2534 (N_2534,N_2440,N_2412);
nor U2535 (N_2535,N_2380,N_2482);
and U2536 (N_2536,N_2417,N_2445);
or U2537 (N_2537,N_2436,N_2422);
nor U2538 (N_2538,N_2497,N_2499);
or U2539 (N_2539,N_2485,N_2472);
xnor U2540 (N_2540,N_2403,N_2388);
and U2541 (N_2541,N_2448,N_2386);
nand U2542 (N_2542,N_2395,N_2439);
nor U2543 (N_2543,N_2473,N_2407);
nor U2544 (N_2544,N_2432,N_2383);
nand U2545 (N_2545,N_2393,N_2401);
and U2546 (N_2546,N_2492,N_2457);
xor U2547 (N_2547,N_2455,N_2438);
nor U2548 (N_2548,N_2405,N_2389);
and U2549 (N_2549,N_2410,N_2476);
nor U2550 (N_2550,N_2399,N_2456);
or U2551 (N_2551,N_2435,N_2416);
xor U2552 (N_2552,N_2468,N_2423);
and U2553 (N_2553,N_2413,N_2424);
xnor U2554 (N_2554,N_2415,N_2377);
xnor U2555 (N_2555,N_2385,N_2400);
xor U2556 (N_2556,N_2451,N_2384);
xor U2557 (N_2557,N_2443,N_2387);
nand U2558 (N_2558,N_2449,N_2471);
and U2559 (N_2559,N_2459,N_2475);
and U2560 (N_2560,N_2479,N_2465);
xor U2561 (N_2561,N_2458,N_2441);
nor U2562 (N_2562,N_2484,N_2408);
nand U2563 (N_2563,N_2412,N_2430);
nand U2564 (N_2564,N_2456,N_2496);
xnor U2565 (N_2565,N_2400,N_2427);
nor U2566 (N_2566,N_2496,N_2471);
xnor U2567 (N_2567,N_2408,N_2389);
nor U2568 (N_2568,N_2382,N_2385);
nor U2569 (N_2569,N_2438,N_2458);
nand U2570 (N_2570,N_2476,N_2457);
nor U2571 (N_2571,N_2394,N_2444);
xor U2572 (N_2572,N_2385,N_2498);
nor U2573 (N_2573,N_2457,N_2456);
and U2574 (N_2574,N_2471,N_2481);
and U2575 (N_2575,N_2463,N_2443);
xor U2576 (N_2576,N_2462,N_2451);
nand U2577 (N_2577,N_2409,N_2418);
nand U2578 (N_2578,N_2469,N_2481);
and U2579 (N_2579,N_2477,N_2436);
xnor U2580 (N_2580,N_2404,N_2380);
nand U2581 (N_2581,N_2442,N_2434);
or U2582 (N_2582,N_2375,N_2405);
nand U2583 (N_2583,N_2409,N_2439);
xnor U2584 (N_2584,N_2448,N_2428);
nor U2585 (N_2585,N_2438,N_2451);
nand U2586 (N_2586,N_2465,N_2467);
nand U2587 (N_2587,N_2459,N_2411);
nor U2588 (N_2588,N_2442,N_2451);
nor U2589 (N_2589,N_2486,N_2414);
or U2590 (N_2590,N_2406,N_2394);
and U2591 (N_2591,N_2382,N_2484);
nand U2592 (N_2592,N_2460,N_2482);
nand U2593 (N_2593,N_2383,N_2487);
xor U2594 (N_2594,N_2400,N_2482);
and U2595 (N_2595,N_2429,N_2483);
or U2596 (N_2596,N_2498,N_2401);
nor U2597 (N_2597,N_2460,N_2447);
and U2598 (N_2598,N_2469,N_2464);
xor U2599 (N_2599,N_2450,N_2431);
or U2600 (N_2600,N_2384,N_2476);
and U2601 (N_2601,N_2497,N_2395);
and U2602 (N_2602,N_2478,N_2450);
and U2603 (N_2603,N_2468,N_2377);
nand U2604 (N_2604,N_2418,N_2445);
nand U2605 (N_2605,N_2402,N_2451);
nand U2606 (N_2606,N_2449,N_2494);
or U2607 (N_2607,N_2450,N_2453);
nand U2608 (N_2608,N_2444,N_2474);
nor U2609 (N_2609,N_2375,N_2427);
nand U2610 (N_2610,N_2413,N_2490);
or U2611 (N_2611,N_2450,N_2440);
or U2612 (N_2612,N_2471,N_2458);
nor U2613 (N_2613,N_2410,N_2475);
nor U2614 (N_2614,N_2405,N_2398);
and U2615 (N_2615,N_2380,N_2474);
xnor U2616 (N_2616,N_2489,N_2470);
or U2617 (N_2617,N_2490,N_2488);
or U2618 (N_2618,N_2409,N_2415);
and U2619 (N_2619,N_2493,N_2484);
nand U2620 (N_2620,N_2449,N_2459);
xor U2621 (N_2621,N_2444,N_2385);
nand U2622 (N_2622,N_2397,N_2404);
xnor U2623 (N_2623,N_2440,N_2443);
xor U2624 (N_2624,N_2379,N_2454);
or U2625 (N_2625,N_2614,N_2553);
nor U2626 (N_2626,N_2581,N_2511);
or U2627 (N_2627,N_2622,N_2595);
or U2628 (N_2628,N_2576,N_2543);
nor U2629 (N_2629,N_2609,N_2551);
or U2630 (N_2630,N_2522,N_2577);
or U2631 (N_2631,N_2601,N_2503);
and U2632 (N_2632,N_2545,N_2607);
xor U2633 (N_2633,N_2570,N_2538);
and U2634 (N_2634,N_2500,N_2572);
and U2635 (N_2635,N_2573,N_2539);
or U2636 (N_2636,N_2535,N_2563);
nand U2637 (N_2637,N_2586,N_2624);
nor U2638 (N_2638,N_2571,N_2596);
and U2639 (N_2639,N_2575,N_2527);
or U2640 (N_2640,N_2517,N_2598);
nand U2641 (N_2641,N_2618,N_2506);
nand U2642 (N_2642,N_2556,N_2608);
nand U2643 (N_2643,N_2593,N_2617);
and U2644 (N_2644,N_2588,N_2557);
nand U2645 (N_2645,N_2621,N_2574);
nor U2646 (N_2646,N_2584,N_2569);
nor U2647 (N_2647,N_2568,N_2565);
nand U2648 (N_2648,N_2532,N_2585);
nor U2649 (N_2649,N_2620,N_2520);
or U2650 (N_2650,N_2513,N_2518);
or U2651 (N_2651,N_2610,N_2619);
xnor U2652 (N_2652,N_2602,N_2550);
or U2653 (N_2653,N_2526,N_2597);
xor U2654 (N_2654,N_2605,N_2583);
nand U2655 (N_2655,N_2566,N_2567);
nor U2656 (N_2656,N_2623,N_2509);
xor U2657 (N_2657,N_2541,N_2615);
and U2658 (N_2658,N_2606,N_2560);
nand U2659 (N_2659,N_2555,N_2504);
nand U2660 (N_2660,N_2536,N_2599);
xor U2661 (N_2661,N_2502,N_2534);
xnor U2662 (N_2662,N_2531,N_2552);
nor U2663 (N_2663,N_2521,N_2529);
nor U2664 (N_2664,N_2559,N_2612);
xnor U2665 (N_2665,N_2505,N_2603);
xnor U2666 (N_2666,N_2611,N_2547);
xnor U2667 (N_2667,N_2594,N_2523);
nor U2668 (N_2668,N_2516,N_2514);
or U2669 (N_2669,N_2537,N_2591);
xor U2670 (N_2670,N_2579,N_2558);
nor U2671 (N_2671,N_2616,N_2554);
xor U2672 (N_2672,N_2544,N_2580);
and U2673 (N_2673,N_2528,N_2562);
nor U2674 (N_2674,N_2587,N_2582);
xor U2675 (N_2675,N_2512,N_2561);
xnor U2676 (N_2676,N_2501,N_2533);
or U2677 (N_2677,N_2548,N_2525);
or U2678 (N_2678,N_2507,N_2510);
nand U2679 (N_2679,N_2600,N_2519);
or U2680 (N_2680,N_2542,N_2564);
xor U2681 (N_2681,N_2613,N_2546);
nor U2682 (N_2682,N_2540,N_2530);
xnor U2683 (N_2683,N_2524,N_2589);
and U2684 (N_2684,N_2549,N_2578);
nand U2685 (N_2685,N_2592,N_2604);
xor U2686 (N_2686,N_2590,N_2508);
or U2687 (N_2687,N_2515,N_2511);
nand U2688 (N_2688,N_2551,N_2508);
or U2689 (N_2689,N_2529,N_2598);
nor U2690 (N_2690,N_2572,N_2507);
nor U2691 (N_2691,N_2587,N_2538);
nand U2692 (N_2692,N_2528,N_2609);
nor U2693 (N_2693,N_2511,N_2596);
and U2694 (N_2694,N_2613,N_2616);
nor U2695 (N_2695,N_2621,N_2616);
or U2696 (N_2696,N_2562,N_2545);
nor U2697 (N_2697,N_2525,N_2596);
nand U2698 (N_2698,N_2515,N_2529);
and U2699 (N_2699,N_2538,N_2575);
and U2700 (N_2700,N_2524,N_2507);
nor U2701 (N_2701,N_2557,N_2504);
xnor U2702 (N_2702,N_2546,N_2579);
and U2703 (N_2703,N_2622,N_2541);
nand U2704 (N_2704,N_2605,N_2565);
nor U2705 (N_2705,N_2605,N_2512);
nor U2706 (N_2706,N_2555,N_2521);
nor U2707 (N_2707,N_2580,N_2611);
and U2708 (N_2708,N_2536,N_2515);
or U2709 (N_2709,N_2521,N_2564);
nand U2710 (N_2710,N_2573,N_2575);
nor U2711 (N_2711,N_2583,N_2579);
xor U2712 (N_2712,N_2617,N_2505);
and U2713 (N_2713,N_2571,N_2610);
or U2714 (N_2714,N_2501,N_2527);
nand U2715 (N_2715,N_2550,N_2544);
xnor U2716 (N_2716,N_2591,N_2612);
and U2717 (N_2717,N_2542,N_2524);
xnor U2718 (N_2718,N_2568,N_2615);
nor U2719 (N_2719,N_2547,N_2608);
nand U2720 (N_2720,N_2521,N_2621);
nand U2721 (N_2721,N_2595,N_2577);
nor U2722 (N_2722,N_2586,N_2576);
nor U2723 (N_2723,N_2526,N_2580);
nor U2724 (N_2724,N_2575,N_2609);
nor U2725 (N_2725,N_2558,N_2512);
nor U2726 (N_2726,N_2594,N_2534);
nand U2727 (N_2727,N_2605,N_2579);
and U2728 (N_2728,N_2549,N_2506);
nand U2729 (N_2729,N_2575,N_2557);
nor U2730 (N_2730,N_2537,N_2511);
xor U2731 (N_2731,N_2620,N_2592);
and U2732 (N_2732,N_2591,N_2522);
and U2733 (N_2733,N_2610,N_2578);
and U2734 (N_2734,N_2592,N_2618);
nand U2735 (N_2735,N_2538,N_2565);
nor U2736 (N_2736,N_2598,N_2611);
nor U2737 (N_2737,N_2530,N_2623);
xnor U2738 (N_2738,N_2510,N_2594);
nor U2739 (N_2739,N_2622,N_2509);
and U2740 (N_2740,N_2613,N_2555);
and U2741 (N_2741,N_2561,N_2577);
and U2742 (N_2742,N_2615,N_2572);
or U2743 (N_2743,N_2562,N_2609);
xnor U2744 (N_2744,N_2511,N_2603);
or U2745 (N_2745,N_2502,N_2595);
nand U2746 (N_2746,N_2616,N_2575);
nand U2747 (N_2747,N_2582,N_2570);
nor U2748 (N_2748,N_2527,N_2538);
xor U2749 (N_2749,N_2570,N_2512);
nand U2750 (N_2750,N_2724,N_2695);
xnor U2751 (N_2751,N_2701,N_2698);
nand U2752 (N_2752,N_2672,N_2749);
nor U2753 (N_2753,N_2638,N_2737);
and U2754 (N_2754,N_2630,N_2697);
xor U2755 (N_2755,N_2625,N_2626);
nor U2756 (N_2756,N_2746,N_2689);
and U2757 (N_2757,N_2738,N_2735);
nand U2758 (N_2758,N_2692,N_2667);
or U2759 (N_2759,N_2693,N_2706);
or U2760 (N_2760,N_2669,N_2703);
or U2761 (N_2761,N_2690,N_2726);
nor U2762 (N_2762,N_2632,N_2688);
xnor U2763 (N_2763,N_2739,N_2700);
xor U2764 (N_2764,N_2666,N_2641);
xor U2765 (N_2765,N_2637,N_2671);
or U2766 (N_2766,N_2660,N_2646);
xnor U2767 (N_2767,N_2723,N_2714);
or U2768 (N_2768,N_2694,N_2687);
and U2769 (N_2769,N_2643,N_2634);
or U2770 (N_2770,N_2730,N_2691);
and U2771 (N_2771,N_2633,N_2685);
and U2772 (N_2772,N_2742,N_2705);
and U2773 (N_2773,N_2748,N_2718);
and U2774 (N_2774,N_2716,N_2673);
nand U2775 (N_2775,N_2657,N_2704);
nand U2776 (N_2776,N_2658,N_2713);
or U2777 (N_2777,N_2732,N_2731);
or U2778 (N_2778,N_2711,N_2644);
or U2779 (N_2779,N_2696,N_2715);
nand U2780 (N_2780,N_2654,N_2699);
and U2781 (N_2781,N_2642,N_2651);
and U2782 (N_2782,N_2659,N_2639);
and U2783 (N_2783,N_2710,N_2670);
nor U2784 (N_2784,N_2627,N_2647);
nand U2785 (N_2785,N_2719,N_2649);
or U2786 (N_2786,N_2680,N_2648);
and U2787 (N_2787,N_2650,N_2663);
and U2788 (N_2788,N_2717,N_2645);
and U2789 (N_2789,N_2727,N_2636);
nor U2790 (N_2790,N_2686,N_2744);
nor U2791 (N_2791,N_2684,N_2631);
nor U2792 (N_2792,N_2747,N_2652);
and U2793 (N_2793,N_2733,N_2702);
nand U2794 (N_2794,N_2729,N_2721);
or U2795 (N_2795,N_2640,N_2725);
nand U2796 (N_2796,N_2720,N_2683);
or U2797 (N_2797,N_2662,N_2745);
and U2798 (N_2798,N_2675,N_2653);
or U2799 (N_2799,N_2708,N_2635);
nor U2800 (N_2800,N_2676,N_2709);
xor U2801 (N_2801,N_2728,N_2665);
nor U2802 (N_2802,N_2681,N_2656);
xor U2803 (N_2803,N_2677,N_2661);
nand U2804 (N_2804,N_2741,N_2674);
or U2805 (N_2805,N_2736,N_2628);
xnor U2806 (N_2806,N_2679,N_2707);
xnor U2807 (N_2807,N_2740,N_2682);
nand U2808 (N_2808,N_2678,N_2629);
nand U2809 (N_2809,N_2664,N_2712);
xnor U2810 (N_2810,N_2734,N_2668);
or U2811 (N_2811,N_2743,N_2722);
or U2812 (N_2812,N_2655,N_2652);
and U2813 (N_2813,N_2727,N_2642);
xor U2814 (N_2814,N_2746,N_2711);
nor U2815 (N_2815,N_2663,N_2653);
and U2816 (N_2816,N_2638,N_2652);
or U2817 (N_2817,N_2650,N_2706);
nand U2818 (N_2818,N_2746,N_2630);
xor U2819 (N_2819,N_2657,N_2716);
or U2820 (N_2820,N_2684,N_2669);
nand U2821 (N_2821,N_2734,N_2704);
xor U2822 (N_2822,N_2625,N_2713);
nor U2823 (N_2823,N_2741,N_2689);
xnor U2824 (N_2824,N_2731,N_2678);
nand U2825 (N_2825,N_2724,N_2638);
and U2826 (N_2826,N_2664,N_2658);
xor U2827 (N_2827,N_2738,N_2639);
and U2828 (N_2828,N_2677,N_2673);
or U2829 (N_2829,N_2679,N_2644);
xor U2830 (N_2830,N_2653,N_2692);
or U2831 (N_2831,N_2680,N_2661);
nand U2832 (N_2832,N_2710,N_2701);
nand U2833 (N_2833,N_2702,N_2662);
nand U2834 (N_2834,N_2633,N_2679);
and U2835 (N_2835,N_2699,N_2714);
nor U2836 (N_2836,N_2656,N_2686);
or U2837 (N_2837,N_2631,N_2697);
nand U2838 (N_2838,N_2681,N_2720);
xnor U2839 (N_2839,N_2638,N_2704);
nor U2840 (N_2840,N_2723,N_2637);
xor U2841 (N_2841,N_2709,N_2717);
or U2842 (N_2842,N_2749,N_2721);
nand U2843 (N_2843,N_2680,N_2637);
nor U2844 (N_2844,N_2702,N_2742);
xor U2845 (N_2845,N_2696,N_2749);
nor U2846 (N_2846,N_2630,N_2714);
and U2847 (N_2847,N_2638,N_2692);
nor U2848 (N_2848,N_2670,N_2738);
xor U2849 (N_2849,N_2679,N_2687);
or U2850 (N_2850,N_2724,N_2641);
or U2851 (N_2851,N_2660,N_2647);
or U2852 (N_2852,N_2739,N_2707);
or U2853 (N_2853,N_2725,N_2635);
or U2854 (N_2854,N_2727,N_2663);
xnor U2855 (N_2855,N_2738,N_2648);
nor U2856 (N_2856,N_2673,N_2682);
or U2857 (N_2857,N_2734,N_2659);
nand U2858 (N_2858,N_2736,N_2667);
xor U2859 (N_2859,N_2661,N_2697);
or U2860 (N_2860,N_2673,N_2741);
nor U2861 (N_2861,N_2626,N_2698);
xnor U2862 (N_2862,N_2673,N_2706);
or U2863 (N_2863,N_2696,N_2747);
or U2864 (N_2864,N_2633,N_2731);
nand U2865 (N_2865,N_2651,N_2652);
or U2866 (N_2866,N_2650,N_2716);
nand U2867 (N_2867,N_2704,N_2729);
nand U2868 (N_2868,N_2733,N_2692);
nor U2869 (N_2869,N_2728,N_2629);
or U2870 (N_2870,N_2712,N_2688);
nor U2871 (N_2871,N_2680,N_2735);
xor U2872 (N_2872,N_2739,N_2667);
and U2873 (N_2873,N_2685,N_2738);
or U2874 (N_2874,N_2632,N_2636);
xor U2875 (N_2875,N_2793,N_2859);
nand U2876 (N_2876,N_2813,N_2869);
xor U2877 (N_2877,N_2824,N_2840);
xnor U2878 (N_2878,N_2767,N_2865);
nor U2879 (N_2879,N_2848,N_2831);
nor U2880 (N_2880,N_2863,N_2750);
and U2881 (N_2881,N_2784,N_2787);
nor U2882 (N_2882,N_2794,N_2776);
nor U2883 (N_2883,N_2760,N_2817);
nor U2884 (N_2884,N_2758,N_2756);
xor U2885 (N_2885,N_2775,N_2801);
xnor U2886 (N_2886,N_2764,N_2851);
and U2887 (N_2887,N_2862,N_2872);
nor U2888 (N_2888,N_2816,N_2781);
or U2889 (N_2889,N_2792,N_2818);
nor U2890 (N_2890,N_2812,N_2815);
or U2891 (N_2891,N_2828,N_2834);
nand U2892 (N_2892,N_2778,N_2796);
xnor U2893 (N_2893,N_2838,N_2762);
nand U2894 (N_2894,N_2821,N_2871);
nand U2895 (N_2895,N_2829,N_2805);
and U2896 (N_2896,N_2783,N_2809);
and U2897 (N_2897,N_2861,N_2779);
nor U2898 (N_2898,N_2833,N_2769);
xor U2899 (N_2899,N_2845,N_2759);
or U2900 (N_2900,N_2811,N_2823);
nand U2901 (N_2901,N_2804,N_2856);
or U2902 (N_2902,N_2826,N_2772);
nor U2903 (N_2903,N_2790,N_2777);
nor U2904 (N_2904,N_2867,N_2780);
or U2905 (N_2905,N_2860,N_2852);
xor U2906 (N_2906,N_2819,N_2752);
xor U2907 (N_2907,N_2827,N_2765);
and U2908 (N_2908,N_2843,N_2873);
or U2909 (N_2909,N_2763,N_2832);
xnor U2910 (N_2910,N_2830,N_2797);
or U2911 (N_2911,N_2841,N_2810);
nor U2912 (N_2912,N_2808,N_2761);
nand U2913 (N_2913,N_2837,N_2799);
nor U2914 (N_2914,N_2798,N_2757);
and U2915 (N_2915,N_2766,N_2754);
xnor U2916 (N_2916,N_2807,N_2822);
or U2917 (N_2917,N_2850,N_2857);
nor U2918 (N_2918,N_2814,N_2789);
xor U2919 (N_2919,N_2786,N_2802);
nor U2920 (N_2920,N_2849,N_2825);
nand U2921 (N_2921,N_2846,N_2788);
and U2922 (N_2922,N_2782,N_2864);
xnor U2923 (N_2923,N_2751,N_2874);
nor U2924 (N_2924,N_2839,N_2774);
nor U2925 (N_2925,N_2791,N_2768);
nor U2926 (N_2926,N_2806,N_2870);
or U2927 (N_2927,N_2835,N_2847);
and U2928 (N_2928,N_2844,N_2785);
xor U2929 (N_2929,N_2855,N_2836);
or U2930 (N_2930,N_2755,N_2800);
nand U2931 (N_2931,N_2753,N_2842);
nand U2932 (N_2932,N_2771,N_2853);
nand U2933 (N_2933,N_2795,N_2803);
or U2934 (N_2934,N_2868,N_2866);
xor U2935 (N_2935,N_2858,N_2773);
nor U2936 (N_2936,N_2770,N_2820);
and U2937 (N_2937,N_2854,N_2804);
xnor U2938 (N_2938,N_2769,N_2802);
or U2939 (N_2939,N_2777,N_2809);
nor U2940 (N_2940,N_2767,N_2868);
or U2941 (N_2941,N_2866,N_2854);
or U2942 (N_2942,N_2820,N_2865);
or U2943 (N_2943,N_2796,N_2773);
and U2944 (N_2944,N_2779,N_2802);
nor U2945 (N_2945,N_2874,N_2807);
and U2946 (N_2946,N_2852,N_2788);
or U2947 (N_2947,N_2760,N_2777);
or U2948 (N_2948,N_2819,N_2817);
nor U2949 (N_2949,N_2838,N_2867);
or U2950 (N_2950,N_2826,N_2854);
xnor U2951 (N_2951,N_2872,N_2751);
nand U2952 (N_2952,N_2847,N_2750);
nand U2953 (N_2953,N_2783,N_2854);
and U2954 (N_2954,N_2835,N_2806);
nand U2955 (N_2955,N_2824,N_2805);
nor U2956 (N_2956,N_2819,N_2847);
nor U2957 (N_2957,N_2838,N_2857);
nand U2958 (N_2958,N_2794,N_2827);
and U2959 (N_2959,N_2752,N_2770);
nor U2960 (N_2960,N_2760,N_2791);
and U2961 (N_2961,N_2852,N_2834);
or U2962 (N_2962,N_2861,N_2801);
xor U2963 (N_2963,N_2782,N_2867);
or U2964 (N_2964,N_2782,N_2824);
xor U2965 (N_2965,N_2759,N_2784);
xor U2966 (N_2966,N_2779,N_2803);
xnor U2967 (N_2967,N_2871,N_2815);
nand U2968 (N_2968,N_2869,N_2776);
xnor U2969 (N_2969,N_2797,N_2763);
nand U2970 (N_2970,N_2816,N_2856);
or U2971 (N_2971,N_2841,N_2858);
or U2972 (N_2972,N_2825,N_2846);
nand U2973 (N_2973,N_2760,N_2836);
and U2974 (N_2974,N_2870,N_2847);
and U2975 (N_2975,N_2856,N_2777);
or U2976 (N_2976,N_2796,N_2812);
and U2977 (N_2977,N_2806,N_2783);
nand U2978 (N_2978,N_2818,N_2832);
nand U2979 (N_2979,N_2834,N_2846);
or U2980 (N_2980,N_2778,N_2836);
or U2981 (N_2981,N_2805,N_2863);
and U2982 (N_2982,N_2760,N_2809);
or U2983 (N_2983,N_2871,N_2800);
or U2984 (N_2984,N_2752,N_2815);
and U2985 (N_2985,N_2868,N_2853);
or U2986 (N_2986,N_2852,N_2759);
xor U2987 (N_2987,N_2772,N_2858);
xor U2988 (N_2988,N_2823,N_2807);
nor U2989 (N_2989,N_2869,N_2752);
xor U2990 (N_2990,N_2756,N_2832);
xor U2991 (N_2991,N_2840,N_2831);
and U2992 (N_2992,N_2857,N_2755);
nor U2993 (N_2993,N_2808,N_2804);
or U2994 (N_2994,N_2869,N_2757);
and U2995 (N_2995,N_2787,N_2801);
and U2996 (N_2996,N_2774,N_2866);
nand U2997 (N_2997,N_2802,N_2869);
and U2998 (N_2998,N_2752,N_2810);
nor U2999 (N_2999,N_2812,N_2786);
xnor U3000 (N_3000,N_2945,N_2942);
nor U3001 (N_3001,N_2971,N_2974);
and U3002 (N_3002,N_2998,N_2935);
nor U3003 (N_3003,N_2887,N_2928);
nor U3004 (N_3004,N_2947,N_2984);
nand U3005 (N_3005,N_2890,N_2885);
xor U3006 (N_3006,N_2975,N_2976);
xnor U3007 (N_3007,N_2899,N_2962);
and U3008 (N_3008,N_2954,N_2967);
and U3009 (N_3009,N_2878,N_2991);
nand U3010 (N_3010,N_2934,N_2925);
nor U3011 (N_3011,N_2988,N_2972);
xor U3012 (N_3012,N_2985,N_2886);
or U3013 (N_3013,N_2875,N_2939);
nand U3014 (N_3014,N_2959,N_2970);
nand U3015 (N_3015,N_2948,N_2903);
and U3016 (N_3016,N_2904,N_2968);
xor U3017 (N_3017,N_2986,N_2880);
and U3018 (N_3018,N_2940,N_2977);
nor U3019 (N_3019,N_2881,N_2891);
nand U3020 (N_3020,N_2938,N_2882);
xor U3021 (N_3021,N_2907,N_2983);
or U3022 (N_3022,N_2981,N_2941);
nor U3023 (N_3023,N_2946,N_2910);
or U3024 (N_3024,N_2924,N_2933);
nand U3025 (N_3025,N_2990,N_2978);
nand U3026 (N_3026,N_2879,N_2895);
and U3027 (N_3027,N_2996,N_2921);
and U3028 (N_3028,N_2953,N_2961);
nor U3029 (N_3029,N_2969,N_2963);
nor U3030 (N_3030,N_2884,N_2909);
nand U3031 (N_3031,N_2966,N_2914);
nand U3032 (N_3032,N_2932,N_2936);
nand U3033 (N_3033,N_2913,N_2908);
or U3034 (N_3034,N_2927,N_2929);
nor U3035 (N_3035,N_2982,N_2992);
nand U3036 (N_3036,N_2916,N_2979);
and U3037 (N_3037,N_2958,N_2957);
nor U3038 (N_3038,N_2920,N_2956);
nor U3039 (N_3039,N_2922,N_2900);
nor U3040 (N_3040,N_2883,N_2926);
nor U3041 (N_3041,N_2912,N_2892);
nor U3042 (N_3042,N_2993,N_2964);
or U3043 (N_3043,N_2987,N_2898);
xnor U3044 (N_3044,N_2930,N_2951);
nand U3045 (N_3045,N_2923,N_2896);
nor U3046 (N_3046,N_2989,N_2949);
and U3047 (N_3047,N_2955,N_2960);
and U3048 (N_3048,N_2905,N_2937);
xnor U3049 (N_3049,N_2952,N_2889);
and U3050 (N_3050,N_2876,N_2943);
nor U3051 (N_3051,N_2897,N_2915);
nand U3052 (N_3052,N_2931,N_2965);
nand U3053 (N_3053,N_2901,N_2973);
nand U3054 (N_3054,N_2994,N_2997);
or U3055 (N_3055,N_2877,N_2950);
and U3056 (N_3056,N_2944,N_2888);
and U3057 (N_3057,N_2902,N_2919);
nor U3058 (N_3058,N_2893,N_2894);
xor U3059 (N_3059,N_2917,N_2980);
xnor U3060 (N_3060,N_2995,N_2918);
xnor U3061 (N_3061,N_2999,N_2911);
and U3062 (N_3062,N_2906,N_2922);
xor U3063 (N_3063,N_2909,N_2958);
nor U3064 (N_3064,N_2980,N_2940);
or U3065 (N_3065,N_2953,N_2938);
or U3066 (N_3066,N_2950,N_2967);
nand U3067 (N_3067,N_2913,N_2994);
nor U3068 (N_3068,N_2875,N_2953);
xor U3069 (N_3069,N_2955,N_2928);
nand U3070 (N_3070,N_2953,N_2965);
nor U3071 (N_3071,N_2970,N_2979);
xor U3072 (N_3072,N_2940,N_2969);
xnor U3073 (N_3073,N_2997,N_2887);
or U3074 (N_3074,N_2972,N_2918);
and U3075 (N_3075,N_2970,N_2963);
nand U3076 (N_3076,N_2946,N_2914);
and U3077 (N_3077,N_2900,N_2966);
xor U3078 (N_3078,N_2973,N_2883);
xnor U3079 (N_3079,N_2929,N_2907);
or U3080 (N_3080,N_2943,N_2904);
nand U3081 (N_3081,N_2936,N_2903);
and U3082 (N_3082,N_2984,N_2884);
nor U3083 (N_3083,N_2930,N_2921);
or U3084 (N_3084,N_2920,N_2988);
xor U3085 (N_3085,N_2966,N_2887);
nand U3086 (N_3086,N_2926,N_2942);
nand U3087 (N_3087,N_2945,N_2982);
xor U3088 (N_3088,N_2916,N_2919);
and U3089 (N_3089,N_2925,N_2882);
nand U3090 (N_3090,N_2985,N_2973);
or U3091 (N_3091,N_2902,N_2941);
nand U3092 (N_3092,N_2926,N_2987);
nand U3093 (N_3093,N_2956,N_2990);
or U3094 (N_3094,N_2970,N_2887);
or U3095 (N_3095,N_2944,N_2999);
xnor U3096 (N_3096,N_2984,N_2918);
nor U3097 (N_3097,N_2986,N_2991);
or U3098 (N_3098,N_2912,N_2949);
xnor U3099 (N_3099,N_2928,N_2940);
xnor U3100 (N_3100,N_2928,N_2909);
xor U3101 (N_3101,N_2916,N_2881);
nor U3102 (N_3102,N_2891,N_2955);
nand U3103 (N_3103,N_2936,N_2941);
xor U3104 (N_3104,N_2998,N_2961);
nor U3105 (N_3105,N_2911,N_2919);
nor U3106 (N_3106,N_2937,N_2951);
xnor U3107 (N_3107,N_2931,N_2919);
nand U3108 (N_3108,N_2990,N_2969);
xnor U3109 (N_3109,N_2918,N_2980);
xnor U3110 (N_3110,N_2928,N_2994);
or U3111 (N_3111,N_2899,N_2903);
or U3112 (N_3112,N_2969,N_2883);
and U3113 (N_3113,N_2921,N_2983);
and U3114 (N_3114,N_2962,N_2900);
xor U3115 (N_3115,N_2913,N_2991);
xnor U3116 (N_3116,N_2936,N_2924);
or U3117 (N_3117,N_2883,N_2983);
xnor U3118 (N_3118,N_2976,N_2886);
and U3119 (N_3119,N_2971,N_2900);
and U3120 (N_3120,N_2949,N_2930);
nor U3121 (N_3121,N_2928,N_2979);
xnor U3122 (N_3122,N_2910,N_2973);
nand U3123 (N_3123,N_2883,N_2895);
and U3124 (N_3124,N_2886,N_2923);
and U3125 (N_3125,N_3010,N_3122);
xnor U3126 (N_3126,N_3061,N_3085);
nor U3127 (N_3127,N_3081,N_3123);
or U3128 (N_3128,N_3065,N_3025);
xnor U3129 (N_3129,N_3056,N_3066);
and U3130 (N_3130,N_3024,N_3075);
nor U3131 (N_3131,N_3014,N_3060);
xor U3132 (N_3132,N_3041,N_3016);
xor U3133 (N_3133,N_3048,N_3007);
nand U3134 (N_3134,N_3057,N_3110);
xnor U3135 (N_3135,N_3036,N_3071);
nand U3136 (N_3136,N_3062,N_3051);
nor U3137 (N_3137,N_3118,N_3070);
nand U3138 (N_3138,N_3019,N_3073);
and U3139 (N_3139,N_3023,N_3052);
nor U3140 (N_3140,N_3124,N_3043);
xnor U3141 (N_3141,N_3084,N_3015);
or U3142 (N_3142,N_3058,N_3077);
or U3143 (N_3143,N_3018,N_3034);
and U3144 (N_3144,N_3109,N_3047);
nor U3145 (N_3145,N_3026,N_3106);
nor U3146 (N_3146,N_3101,N_3074);
or U3147 (N_3147,N_3092,N_3030);
or U3148 (N_3148,N_3102,N_3063);
and U3149 (N_3149,N_3055,N_3029);
xor U3150 (N_3150,N_3120,N_3094);
xor U3151 (N_3151,N_3076,N_3098);
nor U3152 (N_3152,N_3012,N_3103);
and U3153 (N_3153,N_3003,N_3013);
xor U3154 (N_3154,N_3097,N_3045);
nand U3155 (N_3155,N_3040,N_3049);
nand U3156 (N_3156,N_3044,N_3027);
or U3157 (N_3157,N_3089,N_3087);
or U3158 (N_3158,N_3108,N_3114);
or U3159 (N_3159,N_3080,N_3028);
xnor U3160 (N_3160,N_3107,N_3096);
or U3161 (N_3161,N_3035,N_3068);
nand U3162 (N_3162,N_3017,N_3083);
xor U3163 (N_3163,N_3067,N_3001);
or U3164 (N_3164,N_3005,N_3116);
xor U3165 (N_3165,N_3072,N_3046);
nand U3166 (N_3166,N_3093,N_3054);
nor U3167 (N_3167,N_3090,N_3021);
or U3168 (N_3168,N_3032,N_3078);
nor U3169 (N_3169,N_3095,N_3053);
or U3170 (N_3170,N_3031,N_3022);
or U3171 (N_3171,N_3100,N_3039);
or U3172 (N_3172,N_3011,N_3038);
nor U3173 (N_3173,N_3042,N_3002);
nand U3174 (N_3174,N_3059,N_3050);
or U3175 (N_3175,N_3105,N_3113);
nor U3176 (N_3176,N_3121,N_3064);
xor U3177 (N_3177,N_3117,N_3004);
and U3178 (N_3178,N_3033,N_3008);
or U3179 (N_3179,N_3037,N_3099);
nor U3180 (N_3180,N_3086,N_3009);
xor U3181 (N_3181,N_3000,N_3088);
or U3182 (N_3182,N_3006,N_3119);
nor U3183 (N_3183,N_3082,N_3112);
and U3184 (N_3184,N_3091,N_3104);
nor U3185 (N_3185,N_3115,N_3079);
or U3186 (N_3186,N_3020,N_3111);
xor U3187 (N_3187,N_3069,N_3071);
and U3188 (N_3188,N_3035,N_3003);
nor U3189 (N_3189,N_3049,N_3101);
nor U3190 (N_3190,N_3019,N_3112);
and U3191 (N_3191,N_3060,N_3087);
xnor U3192 (N_3192,N_3005,N_3111);
nand U3193 (N_3193,N_3106,N_3124);
xor U3194 (N_3194,N_3093,N_3045);
nand U3195 (N_3195,N_3069,N_3009);
nand U3196 (N_3196,N_3064,N_3020);
or U3197 (N_3197,N_3036,N_3084);
nand U3198 (N_3198,N_3097,N_3049);
and U3199 (N_3199,N_3061,N_3021);
or U3200 (N_3200,N_3031,N_3091);
and U3201 (N_3201,N_3088,N_3076);
xnor U3202 (N_3202,N_3056,N_3095);
nand U3203 (N_3203,N_3007,N_3124);
xnor U3204 (N_3204,N_3097,N_3079);
or U3205 (N_3205,N_3083,N_3103);
nand U3206 (N_3206,N_3064,N_3108);
nand U3207 (N_3207,N_3053,N_3004);
nor U3208 (N_3208,N_3052,N_3044);
nor U3209 (N_3209,N_3097,N_3053);
or U3210 (N_3210,N_3101,N_3052);
nor U3211 (N_3211,N_3122,N_3123);
nand U3212 (N_3212,N_3083,N_3051);
or U3213 (N_3213,N_3063,N_3054);
or U3214 (N_3214,N_3020,N_3091);
xnor U3215 (N_3215,N_3001,N_3037);
and U3216 (N_3216,N_3042,N_3025);
nand U3217 (N_3217,N_3084,N_3097);
and U3218 (N_3218,N_3098,N_3062);
or U3219 (N_3219,N_3068,N_3092);
and U3220 (N_3220,N_3060,N_3038);
or U3221 (N_3221,N_3069,N_3034);
nand U3222 (N_3222,N_3017,N_3063);
nor U3223 (N_3223,N_3063,N_3114);
nand U3224 (N_3224,N_3009,N_3051);
and U3225 (N_3225,N_3073,N_3066);
and U3226 (N_3226,N_3122,N_3097);
and U3227 (N_3227,N_3067,N_3000);
and U3228 (N_3228,N_3073,N_3064);
or U3229 (N_3229,N_3059,N_3057);
xor U3230 (N_3230,N_3006,N_3021);
xnor U3231 (N_3231,N_3095,N_3033);
and U3232 (N_3232,N_3051,N_3122);
and U3233 (N_3233,N_3028,N_3094);
and U3234 (N_3234,N_3072,N_3064);
and U3235 (N_3235,N_3052,N_3010);
or U3236 (N_3236,N_3014,N_3080);
xnor U3237 (N_3237,N_3007,N_3083);
and U3238 (N_3238,N_3117,N_3082);
and U3239 (N_3239,N_3086,N_3011);
and U3240 (N_3240,N_3067,N_3064);
nand U3241 (N_3241,N_3027,N_3017);
or U3242 (N_3242,N_3070,N_3060);
nor U3243 (N_3243,N_3007,N_3088);
nor U3244 (N_3244,N_3003,N_3016);
nand U3245 (N_3245,N_3108,N_3106);
nor U3246 (N_3246,N_3061,N_3074);
xor U3247 (N_3247,N_3035,N_3057);
and U3248 (N_3248,N_3108,N_3086);
xnor U3249 (N_3249,N_3120,N_3050);
nand U3250 (N_3250,N_3192,N_3229);
nand U3251 (N_3251,N_3138,N_3175);
and U3252 (N_3252,N_3186,N_3159);
xor U3253 (N_3253,N_3197,N_3127);
xor U3254 (N_3254,N_3179,N_3209);
or U3255 (N_3255,N_3219,N_3128);
nand U3256 (N_3256,N_3239,N_3233);
nor U3257 (N_3257,N_3167,N_3243);
or U3258 (N_3258,N_3245,N_3135);
and U3259 (N_3259,N_3149,N_3136);
xor U3260 (N_3260,N_3210,N_3178);
nor U3261 (N_3261,N_3129,N_3247);
or U3262 (N_3262,N_3168,N_3207);
xnor U3263 (N_3263,N_3150,N_3162);
nand U3264 (N_3264,N_3148,N_3173);
or U3265 (N_3265,N_3189,N_3188);
or U3266 (N_3266,N_3170,N_3195);
xor U3267 (N_3267,N_3208,N_3194);
nand U3268 (N_3268,N_3139,N_3137);
xor U3269 (N_3269,N_3153,N_3196);
nor U3270 (N_3270,N_3232,N_3140);
xor U3271 (N_3271,N_3226,N_3241);
nand U3272 (N_3272,N_3152,N_3201);
and U3273 (N_3273,N_3177,N_3214);
nand U3274 (N_3274,N_3211,N_3160);
nor U3275 (N_3275,N_3155,N_3228);
or U3276 (N_3276,N_3236,N_3204);
nor U3277 (N_3277,N_3169,N_3174);
nand U3278 (N_3278,N_3240,N_3130);
xor U3279 (N_3279,N_3193,N_3165);
or U3280 (N_3280,N_3180,N_3143);
nor U3281 (N_3281,N_3230,N_3144);
nor U3282 (N_3282,N_3141,N_3215);
xor U3283 (N_3283,N_3227,N_3125);
nand U3284 (N_3284,N_3132,N_3172);
nand U3285 (N_3285,N_3212,N_3146);
and U3286 (N_3286,N_3200,N_3225);
or U3287 (N_3287,N_3164,N_3248);
or U3288 (N_3288,N_3216,N_3133);
nand U3289 (N_3289,N_3199,N_3151);
and U3290 (N_3290,N_3171,N_3126);
nor U3291 (N_3291,N_3202,N_3161);
and U3292 (N_3292,N_3218,N_3145);
nor U3293 (N_3293,N_3191,N_3181);
xor U3294 (N_3294,N_3183,N_3131);
nand U3295 (N_3295,N_3187,N_3234);
nor U3296 (N_3296,N_3242,N_3249);
xor U3297 (N_3297,N_3158,N_3203);
and U3298 (N_3298,N_3246,N_3238);
and U3299 (N_3299,N_3221,N_3182);
or U3300 (N_3300,N_3222,N_3217);
and U3301 (N_3301,N_3223,N_3184);
and U3302 (N_3302,N_3176,N_3213);
nand U3303 (N_3303,N_3156,N_3205);
nor U3304 (N_3304,N_3163,N_3237);
nor U3305 (N_3305,N_3231,N_3220);
and U3306 (N_3306,N_3235,N_3157);
xnor U3307 (N_3307,N_3190,N_3198);
nand U3308 (N_3308,N_3142,N_3147);
and U3309 (N_3309,N_3244,N_3154);
nand U3310 (N_3310,N_3206,N_3166);
nand U3311 (N_3311,N_3224,N_3185);
and U3312 (N_3312,N_3134,N_3158);
nand U3313 (N_3313,N_3237,N_3133);
nor U3314 (N_3314,N_3167,N_3149);
xnor U3315 (N_3315,N_3197,N_3214);
nand U3316 (N_3316,N_3219,N_3232);
xnor U3317 (N_3317,N_3160,N_3198);
nor U3318 (N_3318,N_3187,N_3165);
and U3319 (N_3319,N_3169,N_3164);
xor U3320 (N_3320,N_3211,N_3221);
nor U3321 (N_3321,N_3213,N_3205);
or U3322 (N_3322,N_3194,N_3144);
nand U3323 (N_3323,N_3199,N_3232);
or U3324 (N_3324,N_3215,N_3185);
or U3325 (N_3325,N_3151,N_3241);
and U3326 (N_3326,N_3131,N_3245);
xnor U3327 (N_3327,N_3232,N_3225);
or U3328 (N_3328,N_3139,N_3245);
and U3329 (N_3329,N_3241,N_3193);
nand U3330 (N_3330,N_3223,N_3156);
and U3331 (N_3331,N_3225,N_3191);
xor U3332 (N_3332,N_3200,N_3202);
nand U3333 (N_3333,N_3232,N_3221);
xnor U3334 (N_3334,N_3172,N_3137);
and U3335 (N_3335,N_3222,N_3144);
nand U3336 (N_3336,N_3226,N_3173);
nor U3337 (N_3337,N_3162,N_3129);
xnor U3338 (N_3338,N_3203,N_3205);
xor U3339 (N_3339,N_3223,N_3137);
nor U3340 (N_3340,N_3197,N_3194);
xor U3341 (N_3341,N_3213,N_3189);
and U3342 (N_3342,N_3173,N_3244);
or U3343 (N_3343,N_3244,N_3169);
or U3344 (N_3344,N_3129,N_3238);
or U3345 (N_3345,N_3240,N_3226);
nor U3346 (N_3346,N_3174,N_3179);
or U3347 (N_3347,N_3205,N_3153);
or U3348 (N_3348,N_3200,N_3235);
or U3349 (N_3349,N_3226,N_3216);
nand U3350 (N_3350,N_3228,N_3153);
xnor U3351 (N_3351,N_3177,N_3182);
nand U3352 (N_3352,N_3212,N_3161);
xor U3353 (N_3353,N_3226,N_3175);
or U3354 (N_3354,N_3128,N_3197);
nand U3355 (N_3355,N_3163,N_3170);
or U3356 (N_3356,N_3183,N_3179);
xnor U3357 (N_3357,N_3236,N_3246);
nor U3358 (N_3358,N_3243,N_3234);
nand U3359 (N_3359,N_3236,N_3196);
or U3360 (N_3360,N_3196,N_3223);
and U3361 (N_3361,N_3195,N_3211);
and U3362 (N_3362,N_3191,N_3211);
or U3363 (N_3363,N_3239,N_3220);
nor U3364 (N_3364,N_3135,N_3192);
xnor U3365 (N_3365,N_3159,N_3231);
nor U3366 (N_3366,N_3225,N_3207);
and U3367 (N_3367,N_3144,N_3190);
nor U3368 (N_3368,N_3140,N_3246);
nand U3369 (N_3369,N_3165,N_3189);
nand U3370 (N_3370,N_3188,N_3165);
or U3371 (N_3371,N_3196,N_3165);
xnor U3372 (N_3372,N_3230,N_3225);
xnor U3373 (N_3373,N_3225,N_3174);
nand U3374 (N_3374,N_3182,N_3207);
and U3375 (N_3375,N_3321,N_3368);
nor U3376 (N_3376,N_3332,N_3256);
xor U3377 (N_3377,N_3365,N_3314);
and U3378 (N_3378,N_3271,N_3305);
xnor U3379 (N_3379,N_3295,N_3262);
and U3380 (N_3380,N_3320,N_3264);
or U3381 (N_3381,N_3267,N_3306);
nand U3382 (N_3382,N_3373,N_3277);
nor U3383 (N_3383,N_3269,N_3315);
nand U3384 (N_3384,N_3349,N_3336);
or U3385 (N_3385,N_3309,N_3301);
nor U3386 (N_3386,N_3308,N_3364);
nand U3387 (N_3387,N_3313,N_3316);
nand U3388 (N_3388,N_3352,N_3251);
nor U3389 (N_3389,N_3353,N_3293);
or U3390 (N_3390,N_3268,N_3322);
or U3391 (N_3391,N_3257,N_3288);
nand U3392 (N_3392,N_3359,N_3286);
nor U3393 (N_3393,N_3260,N_3327);
and U3394 (N_3394,N_3326,N_3371);
nand U3395 (N_3395,N_3278,N_3261);
or U3396 (N_3396,N_3355,N_3276);
nand U3397 (N_3397,N_3362,N_3283);
nand U3398 (N_3398,N_3297,N_3275);
xor U3399 (N_3399,N_3319,N_3338);
and U3400 (N_3400,N_3255,N_3290);
nand U3401 (N_3401,N_3285,N_3259);
nor U3402 (N_3402,N_3281,N_3280);
nor U3403 (N_3403,N_3345,N_3330);
nand U3404 (N_3404,N_3342,N_3284);
xor U3405 (N_3405,N_3361,N_3367);
or U3406 (N_3406,N_3250,N_3354);
xor U3407 (N_3407,N_3298,N_3374);
nor U3408 (N_3408,N_3258,N_3333);
nor U3409 (N_3409,N_3358,N_3337);
nor U3410 (N_3410,N_3254,N_3317);
nand U3411 (N_3411,N_3334,N_3351);
and U3412 (N_3412,N_3299,N_3265);
and U3413 (N_3413,N_3296,N_3294);
nand U3414 (N_3414,N_3335,N_3303);
or U3415 (N_3415,N_3266,N_3287);
nor U3416 (N_3416,N_3328,N_3329);
nor U3417 (N_3417,N_3366,N_3372);
xnor U3418 (N_3418,N_3340,N_3291);
nor U3419 (N_3419,N_3302,N_3331);
or U3420 (N_3420,N_3270,N_3289);
or U3421 (N_3421,N_3300,N_3292);
xnor U3422 (N_3422,N_3312,N_3350);
and U3423 (N_3423,N_3339,N_3274);
nor U3424 (N_3424,N_3363,N_3344);
or U3425 (N_3425,N_3346,N_3307);
xor U3426 (N_3426,N_3341,N_3279);
nand U3427 (N_3427,N_3252,N_3369);
nor U3428 (N_3428,N_3370,N_3318);
nor U3429 (N_3429,N_3348,N_3356);
nor U3430 (N_3430,N_3310,N_3343);
nor U3431 (N_3431,N_3311,N_3272);
or U3432 (N_3432,N_3263,N_3273);
or U3433 (N_3433,N_3304,N_3347);
xnor U3434 (N_3434,N_3357,N_3325);
nand U3435 (N_3435,N_3360,N_3282);
and U3436 (N_3436,N_3253,N_3324);
or U3437 (N_3437,N_3323,N_3340);
xor U3438 (N_3438,N_3310,N_3353);
and U3439 (N_3439,N_3280,N_3285);
nor U3440 (N_3440,N_3270,N_3332);
or U3441 (N_3441,N_3312,N_3265);
or U3442 (N_3442,N_3258,N_3319);
nor U3443 (N_3443,N_3254,N_3295);
or U3444 (N_3444,N_3335,N_3283);
nor U3445 (N_3445,N_3317,N_3279);
and U3446 (N_3446,N_3332,N_3301);
or U3447 (N_3447,N_3324,N_3294);
nor U3448 (N_3448,N_3301,N_3349);
nor U3449 (N_3449,N_3372,N_3306);
xnor U3450 (N_3450,N_3365,N_3293);
nand U3451 (N_3451,N_3277,N_3288);
and U3452 (N_3452,N_3264,N_3290);
nor U3453 (N_3453,N_3356,N_3279);
nand U3454 (N_3454,N_3344,N_3326);
nand U3455 (N_3455,N_3292,N_3359);
xor U3456 (N_3456,N_3316,N_3259);
and U3457 (N_3457,N_3319,N_3347);
and U3458 (N_3458,N_3314,N_3342);
and U3459 (N_3459,N_3344,N_3252);
nand U3460 (N_3460,N_3254,N_3355);
nor U3461 (N_3461,N_3350,N_3290);
nand U3462 (N_3462,N_3354,N_3265);
nand U3463 (N_3463,N_3360,N_3307);
nand U3464 (N_3464,N_3277,N_3271);
xor U3465 (N_3465,N_3353,N_3331);
or U3466 (N_3466,N_3339,N_3297);
or U3467 (N_3467,N_3290,N_3315);
and U3468 (N_3468,N_3299,N_3279);
and U3469 (N_3469,N_3330,N_3268);
nand U3470 (N_3470,N_3291,N_3328);
or U3471 (N_3471,N_3273,N_3252);
or U3472 (N_3472,N_3275,N_3357);
xnor U3473 (N_3473,N_3312,N_3260);
xnor U3474 (N_3474,N_3356,N_3274);
and U3475 (N_3475,N_3281,N_3301);
xnor U3476 (N_3476,N_3276,N_3331);
nand U3477 (N_3477,N_3293,N_3322);
nand U3478 (N_3478,N_3320,N_3318);
nand U3479 (N_3479,N_3373,N_3360);
xor U3480 (N_3480,N_3361,N_3293);
nor U3481 (N_3481,N_3364,N_3344);
and U3482 (N_3482,N_3256,N_3292);
and U3483 (N_3483,N_3264,N_3279);
and U3484 (N_3484,N_3339,N_3330);
nor U3485 (N_3485,N_3321,N_3301);
xnor U3486 (N_3486,N_3278,N_3317);
nand U3487 (N_3487,N_3314,N_3294);
nor U3488 (N_3488,N_3272,N_3282);
nand U3489 (N_3489,N_3313,N_3265);
nor U3490 (N_3490,N_3356,N_3253);
and U3491 (N_3491,N_3281,N_3251);
or U3492 (N_3492,N_3260,N_3315);
xnor U3493 (N_3493,N_3369,N_3314);
nor U3494 (N_3494,N_3258,N_3342);
nor U3495 (N_3495,N_3253,N_3351);
and U3496 (N_3496,N_3280,N_3299);
nor U3497 (N_3497,N_3305,N_3295);
or U3498 (N_3498,N_3373,N_3267);
or U3499 (N_3499,N_3258,N_3357);
nand U3500 (N_3500,N_3498,N_3398);
and U3501 (N_3501,N_3433,N_3487);
nor U3502 (N_3502,N_3394,N_3403);
nand U3503 (N_3503,N_3437,N_3423);
nor U3504 (N_3504,N_3462,N_3376);
nand U3505 (N_3505,N_3420,N_3391);
and U3506 (N_3506,N_3414,N_3427);
nand U3507 (N_3507,N_3445,N_3377);
nand U3508 (N_3508,N_3387,N_3444);
nand U3509 (N_3509,N_3466,N_3496);
and U3510 (N_3510,N_3426,N_3421);
or U3511 (N_3511,N_3383,N_3397);
and U3512 (N_3512,N_3453,N_3492);
nand U3513 (N_3513,N_3405,N_3494);
nor U3514 (N_3514,N_3456,N_3399);
nor U3515 (N_3515,N_3448,N_3484);
or U3516 (N_3516,N_3393,N_3473);
nand U3517 (N_3517,N_3485,N_3458);
and U3518 (N_3518,N_3447,N_3480);
or U3519 (N_3519,N_3375,N_3439);
nor U3520 (N_3520,N_3419,N_3428);
nand U3521 (N_3521,N_3443,N_3401);
or U3522 (N_3522,N_3431,N_3407);
nor U3523 (N_3523,N_3460,N_3475);
xnor U3524 (N_3524,N_3479,N_3379);
nand U3525 (N_3525,N_3470,N_3469);
or U3526 (N_3526,N_3415,N_3438);
nor U3527 (N_3527,N_3392,N_3434);
nand U3528 (N_3528,N_3491,N_3422);
and U3529 (N_3529,N_3408,N_3495);
and U3530 (N_3530,N_3380,N_3389);
xnor U3531 (N_3531,N_3385,N_3432);
nand U3532 (N_3532,N_3384,N_3483);
or U3533 (N_3533,N_3442,N_3395);
nor U3534 (N_3534,N_3450,N_3467);
xor U3535 (N_3535,N_3468,N_3435);
nor U3536 (N_3536,N_3497,N_3457);
xnor U3537 (N_3537,N_3430,N_3441);
or U3538 (N_3538,N_3446,N_3455);
or U3539 (N_3539,N_3477,N_3449);
and U3540 (N_3540,N_3413,N_3481);
or U3541 (N_3541,N_3402,N_3452);
nor U3542 (N_3542,N_3382,N_3486);
nor U3543 (N_3543,N_3478,N_3488);
nor U3544 (N_3544,N_3409,N_3404);
and U3545 (N_3545,N_3400,N_3436);
nor U3546 (N_3546,N_3416,N_3396);
xnor U3547 (N_3547,N_3406,N_3454);
or U3548 (N_3548,N_3381,N_3386);
and U3549 (N_3549,N_3463,N_3412);
nor U3550 (N_3550,N_3390,N_3378);
nor U3551 (N_3551,N_3482,N_3388);
xnor U3552 (N_3552,N_3490,N_3493);
or U3553 (N_3553,N_3499,N_3411);
or U3554 (N_3554,N_3464,N_3489);
or U3555 (N_3555,N_3425,N_3440);
and U3556 (N_3556,N_3459,N_3474);
nand U3557 (N_3557,N_3465,N_3471);
and U3558 (N_3558,N_3472,N_3410);
nor U3559 (N_3559,N_3451,N_3476);
or U3560 (N_3560,N_3418,N_3424);
nor U3561 (N_3561,N_3429,N_3461);
xnor U3562 (N_3562,N_3417,N_3493);
nor U3563 (N_3563,N_3471,N_3418);
or U3564 (N_3564,N_3444,N_3389);
nor U3565 (N_3565,N_3419,N_3466);
nor U3566 (N_3566,N_3397,N_3454);
and U3567 (N_3567,N_3421,N_3380);
nor U3568 (N_3568,N_3495,N_3401);
nand U3569 (N_3569,N_3426,N_3393);
nor U3570 (N_3570,N_3487,N_3388);
xnor U3571 (N_3571,N_3441,N_3419);
and U3572 (N_3572,N_3467,N_3483);
or U3573 (N_3573,N_3403,N_3384);
and U3574 (N_3574,N_3494,N_3480);
and U3575 (N_3575,N_3389,N_3438);
nor U3576 (N_3576,N_3377,N_3466);
nand U3577 (N_3577,N_3471,N_3490);
nand U3578 (N_3578,N_3410,N_3451);
nor U3579 (N_3579,N_3429,N_3497);
xnor U3580 (N_3580,N_3497,N_3470);
and U3581 (N_3581,N_3491,N_3399);
or U3582 (N_3582,N_3392,N_3398);
xor U3583 (N_3583,N_3486,N_3489);
xnor U3584 (N_3584,N_3456,N_3446);
nand U3585 (N_3585,N_3491,N_3414);
nand U3586 (N_3586,N_3443,N_3454);
or U3587 (N_3587,N_3486,N_3495);
or U3588 (N_3588,N_3496,N_3387);
xor U3589 (N_3589,N_3491,N_3430);
nor U3590 (N_3590,N_3380,N_3408);
nand U3591 (N_3591,N_3445,N_3440);
nand U3592 (N_3592,N_3382,N_3457);
xor U3593 (N_3593,N_3402,N_3433);
or U3594 (N_3594,N_3448,N_3381);
xor U3595 (N_3595,N_3418,N_3488);
or U3596 (N_3596,N_3481,N_3476);
nand U3597 (N_3597,N_3404,N_3380);
or U3598 (N_3598,N_3407,N_3439);
xnor U3599 (N_3599,N_3466,N_3400);
and U3600 (N_3600,N_3408,N_3483);
xnor U3601 (N_3601,N_3382,N_3408);
or U3602 (N_3602,N_3483,N_3424);
or U3603 (N_3603,N_3379,N_3405);
nand U3604 (N_3604,N_3450,N_3409);
nor U3605 (N_3605,N_3426,N_3466);
and U3606 (N_3606,N_3388,N_3386);
nand U3607 (N_3607,N_3483,N_3488);
and U3608 (N_3608,N_3392,N_3413);
nand U3609 (N_3609,N_3491,N_3484);
nor U3610 (N_3610,N_3439,N_3423);
or U3611 (N_3611,N_3471,N_3482);
or U3612 (N_3612,N_3401,N_3390);
xnor U3613 (N_3613,N_3382,N_3416);
nor U3614 (N_3614,N_3407,N_3440);
nand U3615 (N_3615,N_3492,N_3481);
and U3616 (N_3616,N_3467,N_3463);
nor U3617 (N_3617,N_3383,N_3451);
nor U3618 (N_3618,N_3482,N_3381);
and U3619 (N_3619,N_3407,N_3454);
nand U3620 (N_3620,N_3382,N_3498);
or U3621 (N_3621,N_3391,N_3398);
or U3622 (N_3622,N_3496,N_3427);
or U3623 (N_3623,N_3401,N_3387);
xnor U3624 (N_3624,N_3416,N_3475);
nor U3625 (N_3625,N_3562,N_3510);
nand U3626 (N_3626,N_3605,N_3569);
nor U3627 (N_3627,N_3536,N_3583);
xnor U3628 (N_3628,N_3596,N_3620);
and U3629 (N_3629,N_3579,N_3544);
and U3630 (N_3630,N_3601,N_3556);
xnor U3631 (N_3631,N_3527,N_3595);
nand U3632 (N_3632,N_3559,N_3554);
and U3633 (N_3633,N_3607,N_3572);
or U3634 (N_3634,N_3535,N_3528);
nand U3635 (N_3635,N_3520,N_3546);
nand U3636 (N_3636,N_3543,N_3622);
and U3637 (N_3637,N_3555,N_3533);
nor U3638 (N_3638,N_3557,N_3578);
or U3639 (N_3639,N_3534,N_3537);
nor U3640 (N_3640,N_3552,N_3621);
nor U3641 (N_3641,N_3500,N_3624);
or U3642 (N_3642,N_3608,N_3511);
or U3643 (N_3643,N_3506,N_3542);
nor U3644 (N_3644,N_3560,N_3539);
and U3645 (N_3645,N_3576,N_3603);
or U3646 (N_3646,N_3521,N_3564);
nand U3647 (N_3647,N_3577,N_3558);
xnor U3648 (N_3648,N_3617,N_3575);
or U3649 (N_3649,N_3594,N_3547);
nor U3650 (N_3650,N_3529,N_3604);
xnor U3651 (N_3651,N_3549,N_3548);
xor U3652 (N_3652,N_3609,N_3573);
nand U3653 (N_3653,N_3522,N_3592);
nor U3654 (N_3654,N_3611,N_3553);
or U3655 (N_3655,N_3570,N_3516);
nor U3656 (N_3656,N_3602,N_3591);
xnor U3657 (N_3657,N_3610,N_3563);
xor U3658 (N_3658,N_3581,N_3585);
nor U3659 (N_3659,N_3530,N_3580);
xor U3660 (N_3660,N_3565,N_3589);
and U3661 (N_3661,N_3523,N_3613);
and U3662 (N_3662,N_3623,N_3606);
xnor U3663 (N_3663,N_3588,N_3504);
nor U3664 (N_3664,N_3540,N_3574);
and U3665 (N_3665,N_3566,N_3512);
xnor U3666 (N_3666,N_3618,N_3503);
nand U3667 (N_3667,N_3598,N_3593);
and U3668 (N_3668,N_3525,N_3524);
nand U3669 (N_3669,N_3519,N_3545);
xnor U3670 (N_3670,N_3505,N_3518);
nand U3671 (N_3671,N_3612,N_3502);
or U3672 (N_3672,N_3597,N_3507);
and U3673 (N_3673,N_3532,N_3550);
xnor U3674 (N_3674,N_3616,N_3541);
or U3675 (N_3675,N_3586,N_3615);
or U3676 (N_3676,N_3587,N_3514);
xor U3677 (N_3677,N_3614,N_3619);
and U3678 (N_3678,N_3551,N_3526);
xor U3679 (N_3679,N_3508,N_3509);
and U3680 (N_3680,N_3513,N_3561);
xnor U3681 (N_3681,N_3584,N_3517);
or U3682 (N_3682,N_3538,N_3600);
xnor U3683 (N_3683,N_3567,N_3568);
nand U3684 (N_3684,N_3571,N_3590);
and U3685 (N_3685,N_3531,N_3515);
xnor U3686 (N_3686,N_3501,N_3599);
nand U3687 (N_3687,N_3582,N_3608);
nor U3688 (N_3688,N_3611,N_3624);
nor U3689 (N_3689,N_3566,N_3605);
xor U3690 (N_3690,N_3536,N_3557);
nor U3691 (N_3691,N_3515,N_3574);
nand U3692 (N_3692,N_3579,N_3612);
or U3693 (N_3693,N_3585,N_3529);
xnor U3694 (N_3694,N_3569,N_3551);
or U3695 (N_3695,N_3569,N_3565);
or U3696 (N_3696,N_3608,N_3567);
and U3697 (N_3697,N_3529,N_3540);
xor U3698 (N_3698,N_3508,N_3548);
xor U3699 (N_3699,N_3568,N_3551);
and U3700 (N_3700,N_3601,N_3503);
and U3701 (N_3701,N_3603,N_3596);
and U3702 (N_3702,N_3581,N_3507);
or U3703 (N_3703,N_3574,N_3557);
xor U3704 (N_3704,N_3526,N_3529);
nor U3705 (N_3705,N_3516,N_3574);
or U3706 (N_3706,N_3581,N_3609);
or U3707 (N_3707,N_3595,N_3577);
nor U3708 (N_3708,N_3582,N_3564);
or U3709 (N_3709,N_3517,N_3502);
nor U3710 (N_3710,N_3608,N_3510);
nand U3711 (N_3711,N_3596,N_3614);
or U3712 (N_3712,N_3544,N_3573);
nand U3713 (N_3713,N_3601,N_3616);
nand U3714 (N_3714,N_3561,N_3609);
and U3715 (N_3715,N_3517,N_3586);
nand U3716 (N_3716,N_3590,N_3599);
and U3717 (N_3717,N_3622,N_3539);
nor U3718 (N_3718,N_3507,N_3573);
nand U3719 (N_3719,N_3573,N_3528);
and U3720 (N_3720,N_3563,N_3557);
and U3721 (N_3721,N_3608,N_3598);
and U3722 (N_3722,N_3519,N_3530);
or U3723 (N_3723,N_3609,N_3543);
and U3724 (N_3724,N_3594,N_3587);
or U3725 (N_3725,N_3532,N_3503);
or U3726 (N_3726,N_3571,N_3624);
xor U3727 (N_3727,N_3509,N_3608);
nand U3728 (N_3728,N_3589,N_3622);
nor U3729 (N_3729,N_3573,N_3542);
nor U3730 (N_3730,N_3614,N_3526);
and U3731 (N_3731,N_3551,N_3607);
or U3732 (N_3732,N_3599,N_3550);
and U3733 (N_3733,N_3591,N_3621);
xor U3734 (N_3734,N_3619,N_3601);
xor U3735 (N_3735,N_3528,N_3514);
nor U3736 (N_3736,N_3513,N_3570);
nand U3737 (N_3737,N_3560,N_3588);
nand U3738 (N_3738,N_3611,N_3550);
nor U3739 (N_3739,N_3574,N_3556);
xnor U3740 (N_3740,N_3620,N_3500);
xnor U3741 (N_3741,N_3549,N_3531);
nand U3742 (N_3742,N_3507,N_3563);
nand U3743 (N_3743,N_3514,N_3548);
and U3744 (N_3744,N_3575,N_3585);
nand U3745 (N_3745,N_3577,N_3579);
nand U3746 (N_3746,N_3546,N_3565);
or U3747 (N_3747,N_3575,N_3601);
nand U3748 (N_3748,N_3526,N_3544);
or U3749 (N_3749,N_3624,N_3516);
nand U3750 (N_3750,N_3667,N_3674);
nor U3751 (N_3751,N_3634,N_3650);
or U3752 (N_3752,N_3643,N_3653);
xor U3753 (N_3753,N_3737,N_3663);
xnor U3754 (N_3754,N_3719,N_3740);
and U3755 (N_3755,N_3641,N_3651);
nand U3756 (N_3756,N_3733,N_3696);
or U3757 (N_3757,N_3654,N_3725);
nand U3758 (N_3758,N_3741,N_3706);
nor U3759 (N_3759,N_3633,N_3664);
and U3760 (N_3760,N_3680,N_3701);
or U3761 (N_3761,N_3632,N_3662);
xor U3762 (N_3762,N_3747,N_3697);
nand U3763 (N_3763,N_3656,N_3657);
or U3764 (N_3764,N_3670,N_3721);
xor U3765 (N_3765,N_3636,N_3715);
xor U3766 (N_3766,N_3673,N_3660);
or U3767 (N_3767,N_3698,N_3744);
or U3768 (N_3768,N_3724,N_3720);
nor U3769 (N_3769,N_3742,N_3732);
xor U3770 (N_3770,N_3718,N_3642);
xor U3771 (N_3771,N_3694,N_3699);
nand U3772 (N_3772,N_3745,N_3709);
and U3773 (N_3773,N_3691,N_3628);
xnor U3774 (N_3774,N_3648,N_3711);
nand U3775 (N_3775,N_3731,N_3700);
nand U3776 (N_3776,N_3710,N_3659);
or U3777 (N_3777,N_3734,N_3644);
nor U3778 (N_3778,N_3682,N_3723);
or U3779 (N_3779,N_3702,N_3743);
or U3780 (N_3780,N_3681,N_3748);
xor U3781 (N_3781,N_3730,N_3666);
or U3782 (N_3782,N_3655,N_3672);
or U3783 (N_3783,N_3729,N_3626);
nand U3784 (N_3784,N_3638,N_3713);
or U3785 (N_3785,N_3695,N_3679);
and U3786 (N_3786,N_3627,N_3692);
xor U3787 (N_3787,N_3736,N_3693);
and U3788 (N_3788,N_3739,N_3738);
xnor U3789 (N_3789,N_3716,N_3625);
xnor U3790 (N_3790,N_3678,N_3722);
or U3791 (N_3791,N_3668,N_3629);
and U3792 (N_3792,N_3688,N_3728);
and U3793 (N_3793,N_3685,N_3683);
nand U3794 (N_3794,N_3669,N_3717);
nor U3795 (N_3795,N_3677,N_3635);
nand U3796 (N_3796,N_3689,N_3684);
and U3797 (N_3797,N_3645,N_3705);
and U3798 (N_3798,N_3727,N_3746);
nor U3799 (N_3799,N_3637,N_3735);
or U3800 (N_3800,N_3703,N_3675);
xnor U3801 (N_3801,N_3665,N_3707);
and U3802 (N_3802,N_3671,N_3631);
xnor U3803 (N_3803,N_3686,N_3639);
nor U3804 (N_3804,N_3690,N_3652);
and U3805 (N_3805,N_3726,N_3646);
xor U3806 (N_3806,N_3630,N_3640);
nor U3807 (N_3807,N_3704,N_3708);
or U3808 (N_3808,N_3714,N_3676);
xnor U3809 (N_3809,N_3658,N_3649);
and U3810 (N_3810,N_3687,N_3647);
xnor U3811 (N_3811,N_3661,N_3712);
nand U3812 (N_3812,N_3749,N_3642);
xnor U3813 (N_3813,N_3650,N_3695);
nor U3814 (N_3814,N_3669,N_3693);
xor U3815 (N_3815,N_3689,N_3664);
xnor U3816 (N_3816,N_3677,N_3722);
nor U3817 (N_3817,N_3743,N_3747);
nand U3818 (N_3818,N_3724,N_3661);
or U3819 (N_3819,N_3713,N_3719);
nand U3820 (N_3820,N_3731,N_3659);
nand U3821 (N_3821,N_3728,N_3740);
nor U3822 (N_3822,N_3736,N_3685);
or U3823 (N_3823,N_3694,N_3674);
xor U3824 (N_3824,N_3733,N_3657);
nor U3825 (N_3825,N_3702,N_3744);
xnor U3826 (N_3826,N_3647,N_3748);
or U3827 (N_3827,N_3668,N_3705);
xor U3828 (N_3828,N_3728,N_3646);
or U3829 (N_3829,N_3662,N_3669);
xnor U3830 (N_3830,N_3660,N_3694);
nand U3831 (N_3831,N_3667,N_3681);
nand U3832 (N_3832,N_3715,N_3733);
nand U3833 (N_3833,N_3705,N_3693);
nand U3834 (N_3834,N_3660,N_3736);
nor U3835 (N_3835,N_3688,N_3723);
nor U3836 (N_3836,N_3685,N_3679);
nand U3837 (N_3837,N_3728,N_3700);
nand U3838 (N_3838,N_3640,N_3724);
or U3839 (N_3839,N_3651,N_3636);
nor U3840 (N_3840,N_3689,N_3749);
xnor U3841 (N_3841,N_3716,N_3693);
xor U3842 (N_3842,N_3637,N_3665);
and U3843 (N_3843,N_3658,N_3736);
and U3844 (N_3844,N_3718,N_3741);
and U3845 (N_3845,N_3730,N_3639);
and U3846 (N_3846,N_3732,N_3708);
or U3847 (N_3847,N_3743,N_3646);
and U3848 (N_3848,N_3647,N_3747);
xor U3849 (N_3849,N_3656,N_3658);
xnor U3850 (N_3850,N_3666,N_3682);
or U3851 (N_3851,N_3731,N_3684);
nor U3852 (N_3852,N_3646,N_3676);
nor U3853 (N_3853,N_3692,N_3666);
or U3854 (N_3854,N_3707,N_3749);
nand U3855 (N_3855,N_3638,N_3639);
xor U3856 (N_3856,N_3656,N_3669);
and U3857 (N_3857,N_3718,N_3654);
and U3858 (N_3858,N_3709,N_3647);
nor U3859 (N_3859,N_3663,N_3735);
and U3860 (N_3860,N_3711,N_3703);
or U3861 (N_3861,N_3696,N_3699);
or U3862 (N_3862,N_3743,N_3636);
nand U3863 (N_3863,N_3735,N_3727);
or U3864 (N_3864,N_3677,N_3724);
nor U3865 (N_3865,N_3719,N_3646);
or U3866 (N_3866,N_3745,N_3733);
nor U3867 (N_3867,N_3690,N_3682);
xor U3868 (N_3868,N_3714,N_3652);
nand U3869 (N_3869,N_3700,N_3695);
nand U3870 (N_3870,N_3661,N_3703);
nor U3871 (N_3871,N_3634,N_3655);
nor U3872 (N_3872,N_3710,N_3745);
nor U3873 (N_3873,N_3701,N_3707);
nand U3874 (N_3874,N_3634,N_3648);
nand U3875 (N_3875,N_3870,N_3778);
nand U3876 (N_3876,N_3835,N_3865);
nand U3877 (N_3877,N_3771,N_3768);
or U3878 (N_3878,N_3813,N_3760);
and U3879 (N_3879,N_3794,N_3860);
or U3880 (N_3880,N_3802,N_3789);
and U3881 (N_3881,N_3750,N_3783);
or U3882 (N_3882,N_3777,N_3753);
and U3883 (N_3883,N_3866,N_3805);
nor U3884 (N_3884,N_3759,N_3772);
nand U3885 (N_3885,N_3827,N_3793);
or U3886 (N_3886,N_3845,N_3814);
or U3887 (N_3887,N_3801,N_3761);
nor U3888 (N_3888,N_3803,N_3785);
and U3889 (N_3889,N_3844,N_3804);
nand U3890 (N_3890,N_3810,N_3829);
xnor U3891 (N_3891,N_3811,N_3766);
or U3892 (N_3892,N_3790,N_3792);
or U3893 (N_3893,N_3779,N_3787);
nand U3894 (N_3894,N_3769,N_3840);
and U3895 (N_3895,N_3826,N_3873);
and U3896 (N_3896,N_3822,N_3854);
and U3897 (N_3897,N_3800,N_3820);
and U3898 (N_3898,N_3856,N_3861);
xor U3899 (N_3899,N_3780,N_3839);
xnor U3900 (N_3900,N_3819,N_3837);
or U3901 (N_3901,N_3770,N_3773);
nor U3902 (N_3902,N_3857,N_3830);
and U3903 (N_3903,N_3797,N_3776);
and U3904 (N_3904,N_3834,N_3815);
xor U3905 (N_3905,N_3752,N_3751);
xor U3906 (N_3906,N_3850,N_3812);
nor U3907 (N_3907,N_3756,N_3808);
and U3908 (N_3908,N_3754,N_3775);
and U3909 (N_3909,N_3849,N_3825);
and U3910 (N_3910,N_3828,N_3824);
nor U3911 (N_3911,N_3758,N_3765);
xnor U3912 (N_3912,N_3791,N_3858);
nand U3913 (N_3913,N_3841,N_3823);
and U3914 (N_3914,N_3862,N_3872);
and U3915 (N_3915,N_3799,N_3871);
xnor U3916 (N_3916,N_3853,N_3782);
xnor U3917 (N_3917,N_3762,N_3874);
or U3918 (N_3918,N_3868,N_3831);
and U3919 (N_3919,N_3842,N_3855);
nor U3920 (N_3920,N_3757,N_3807);
nand U3921 (N_3921,N_3869,N_3816);
nor U3922 (N_3922,N_3848,N_3863);
xnor U3923 (N_3923,N_3763,N_3774);
xor U3924 (N_3924,N_3867,N_3809);
xor U3925 (N_3925,N_3781,N_3818);
and U3926 (N_3926,N_3852,N_3833);
xor U3927 (N_3927,N_3788,N_3764);
or U3928 (N_3928,N_3859,N_3832);
nor U3929 (N_3929,N_3784,N_3806);
or U3930 (N_3930,N_3795,N_3817);
nor U3931 (N_3931,N_3821,N_3843);
and U3932 (N_3932,N_3838,N_3847);
nand U3933 (N_3933,N_3846,N_3786);
nand U3934 (N_3934,N_3755,N_3864);
nor U3935 (N_3935,N_3796,N_3836);
nand U3936 (N_3936,N_3767,N_3798);
and U3937 (N_3937,N_3851,N_3864);
or U3938 (N_3938,N_3777,N_3809);
nor U3939 (N_3939,N_3770,N_3854);
xnor U3940 (N_3940,N_3821,N_3767);
and U3941 (N_3941,N_3776,N_3795);
or U3942 (N_3942,N_3752,N_3851);
nand U3943 (N_3943,N_3817,N_3866);
nand U3944 (N_3944,N_3805,N_3776);
nand U3945 (N_3945,N_3777,N_3769);
xor U3946 (N_3946,N_3833,N_3773);
nand U3947 (N_3947,N_3839,N_3857);
nand U3948 (N_3948,N_3786,N_3785);
nand U3949 (N_3949,N_3855,N_3806);
or U3950 (N_3950,N_3775,N_3788);
and U3951 (N_3951,N_3822,N_3817);
nor U3952 (N_3952,N_3843,N_3781);
nand U3953 (N_3953,N_3795,N_3818);
or U3954 (N_3954,N_3789,N_3837);
nand U3955 (N_3955,N_3845,N_3873);
xnor U3956 (N_3956,N_3782,N_3800);
and U3957 (N_3957,N_3769,N_3816);
xnor U3958 (N_3958,N_3804,N_3761);
nand U3959 (N_3959,N_3854,N_3806);
nand U3960 (N_3960,N_3753,N_3779);
nor U3961 (N_3961,N_3757,N_3845);
xor U3962 (N_3962,N_3757,N_3859);
or U3963 (N_3963,N_3866,N_3811);
nand U3964 (N_3964,N_3871,N_3762);
nand U3965 (N_3965,N_3842,N_3850);
and U3966 (N_3966,N_3843,N_3754);
xnor U3967 (N_3967,N_3821,N_3854);
nor U3968 (N_3968,N_3851,N_3772);
or U3969 (N_3969,N_3813,N_3759);
nand U3970 (N_3970,N_3821,N_3866);
xor U3971 (N_3971,N_3843,N_3820);
nor U3972 (N_3972,N_3849,N_3786);
or U3973 (N_3973,N_3760,N_3826);
xor U3974 (N_3974,N_3818,N_3750);
xnor U3975 (N_3975,N_3751,N_3763);
xor U3976 (N_3976,N_3849,N_3867);
nor U3977 (N_3977,N_3829,N_3858);
or U3978 (N_3978,N_3758,N_3809);
and U3979 (N_3979,N_3832,N_3823);
nor U3980 (N_3980,N_3753,N_3847);
nand U3981 (N_3981,N_3786,N_3826);
nor U3982 (N_3982,N_3852,N_3765);
nand U3983 (N_3983,N_3778,N_3753);
xnor U3984 (N_3984,N_3780,N_3792);
nor U3985 (N_3985,N_3751,N_3867);
or U3986 (N_3986,N_3855,N_3867);
xnor U3987 (N_3987,N_3824,N_3783);
or U3988 (N_3988,N_3777,N_3774);
xor U3989 (N_3989,N_3789,N_3853);
nor U3990 (N_3990,N_3789,N_3819);
or U3991 (N_3991,N_3837,N_3790);
nor U3992 (N_3992,N_3831,N_3829);
or U3993 (N_3993,N_3856,N_3838);
and U3994 (N_3994,N_3773,N_3832);
or U3995 (N_3995,N_3784,N_3779);
or U3996 (N_3996,N_3787,N_3866);
nand U3997 (N_3997,N_3868,N_3852);
and U3998 (N_3998,N_3831,N_3775);
and U3999 (N_3999,N_3829,N_3778);
xnor U4000 (N_4000,N_3928,N_3976);
xor U4001 (N_4001,N_3960,N_3921);
nor U4002 (N_4002,N_3996,N_3899);
nand U4003 (N_4003,N_3970,N_3911);
and U4004 (N_4004,N_3886,N_3997);
or U4005 (N_4005,N_3936,N_3957);
nor U4006 (N_4006,N_3946,N_3944);
xor U4007 (N_4007,N_3918,N_3982);
and U4008 (N_4008,N_3895,N_3902);
or U4009 (N_4009,N_3994,N_3980);
nor U4010 (N_4010,N_3896,N_3907);
xor U4011 (N_4011,N_3954,N_3920);
nor U4012 (N_4012,N_3875,N_3887);
xnor U4013 (N_4013,N_3938,N_3979);
and U4014 (N_4014,N_3922,N_3991);
xor U4015 (N_4015,N_3945,N_3881);
nand U4016 (N_4016,N_3910,N_3962);
nand U4017 (N_4017,N_3914,N_3879);
nor U4018 (N_4018,N_3972,N_3951);
and U4019 (N_4019,N_3880,N_3909);
nand U4020 (N_4020,N_3898,N_3933);
and U4021 (N_4021,N_3998,N_3992);
or U4022 (N_4022,N_3897,N_3961);
nand U4023 (N_4023,N_3892,N_3995);
nor U4024 (N_4024,N_3953,N_3964);
and U4025 (N_4025,N_3915,N_3990);
nand U4026 (N_4026,N_3877,N_3973);
xor U4027 (N_4027,N_3966,N_3988);
xor U4028 (N_4028,N_3893,N_3927);
nor U4029 (N_4029,N_3932,N_3974);
nor U4030 (N_4030,N_3889,N_3985);
xnor U4031 (N_4031,N_3882,N_3941);
and U4032 (N_4032,N_3950,N_3908);
nand U4033 (N_4033,N_3878,N_3948);
and U4034 (N_4034,N_3943,N_3916);
xor U4035 (N_4035,N_3924,N_3987);
nor U4036 (N_4036,N_3891,N_3934);
xor U4037 (N_4037,N_3926,N_3894);
xor U4038 (N_4038,N_3959,N_3903);
nand U4039 (N_4039,N_3975,N_3888);
nand U4040 (N_4040,N_3930,N_3967);
nor U4041 (N_4041,N_3904,N_3986);
and U4042 (N_4042,N_3925,N_3989);
nor U4043 (N_4043,N_3969,N_3929);
and U4044 (N_4044,N_3968,N_3942);
nor U4045 (N_4045,N_3919,N_3981);
or U4046 (N_4046,N_3955,N_3900);
and U4047 (N_4047,N_3949,N_3978);
or U4048 (N_4048,N_3937,N_3984);
nor U4049 (N_4049,N_3931,N_3935);
nand U4050 (N_4050,N_3883,N_3890);
and U4051 (N_4051,N_3993,N_3906);
or U4052 (N_4052,N_3913,N_3923);
nor U4053 (N_4053,N_3884,N_3963);
nor U4054 (N_4054,N_3912,N_3905);
nor U4055 (N_4055,N_3956,N_3958);
and U4056 (N_4056,N_3876,N_3917);
or U4057 (N_4057,N_3965,N_3999);
or U4058 (N_4058,N_3901,N_3939);
nor U4059 (N_4059,N_3977,N_3983);
nand U4060 (N_4060,N_3940,N_3947);
nor U4061 (N_4061,N_3885,N_3971);
and U4062 (N_4062,N_3952,N_3918);
xor U4063 (N_4063,N_3999,N_3915);
nor U4064 (N_4064,N_3989,N_3908);
and U4065 (N_4065,N_3875,N_3948);
and U4066 (N_4066,N_3927,N_3966);
nor U4067 (N_4067,N_3947,N_3975);
nand U4068 (N_4068,N_3988,N_3920);
nand U4069 (N_4069,N_3965,N_3877);
and U4070 (N_4070,N_3964,N_3982);
and U4071 (N_4071,N_3922,N_3975);
nand U4072 (N_4072,N_3935,N_3916);
nand U4073 (N_4073,N_3953,N_3885);
and U4074 (N_4074,N_3933,N_3969);
and U4075 (N_4075,N_3878,N_3880);
nor U4076 (N_4076,N_3922,N_3925);
and U4077 (N_4077,N_3977,N_3932);
or U4078 (N_4078,N_3965,N_3948);
or U4079 (N_4079,N_3924,N_3905);
nor U4080 (N_4080,N_3889,N_3924);
and U4081 (N_4081,N_3938,N_3881);
nor U4082 (N_4082,N_3883,N_3905);
nor U4083 (N_4083,N_3961,N_3955);
or U4084 (N_4084,N_3982,N_3920);
or U4085 (N_4085,N_3932,N_3894);
nand U4086 (N_4086,N_3976,N_3996);
nand U4087 (N_4087,N_3882,N_3888);
xor U4088 (N_4088,N_3958,N_3952);
xnor U4089 (N_4089,N_3984,N_3904);
or U4090 (N_4090,N_3969,N_3898);
nand U4091 (N_4091,N_3897,N_3950);
nand U4092 (N_4092,N_3958,N_3947);
nand U4093 (N_4093,N_3920,N_3975);
nor U4094 (N_4094,N_3978,N_3878);
nand U4095 (N_4095,N_3920,N_3940);
or U4096 (N_4096,N_3925,N_3877);
and U4097 (N_4097,N_3931,N_3875);
nand U4098 (N_4098,N_3902,N_3961);
xnor U4099 (N_4099,N_3910,N_3976);
or U4100 (N_4100,N_3975,N_3973);
xor U4101 (N_4101,N_3985,N_3906);
xor U4102 (N_4102,N_3986,N_3906);
xnor U4103 (N_4103,N_3887,N_3979);
nor U4104 (N_4104,N_3898,N_3942);
or U4105 (N_4105,N_3917,N_3915);
nand U4106 (N_4106,N_3890,N_3968);
or U4107 (N_4107,N_3896,N_3909);
or U4108 (N_4108,N_3945,N_3907);
xnor U4109 (N_4109,N_3957,N_3949);
nand U4110 (N_4110,N_3904,N_3930);
xor U4111 (N_4111,N_3916,N_3888);
nand U4112 (N_4112,N_3986,N_3981);
or U4113 (N_4113,N_3987,N_3938);
nor U4114 (N_4114,N_3960,N_3963);
xnor U4115 (N_4115,N_3964,N_3884);
and U4116 (N_4116,N_3934,N_3932);
xor U4117 (N_4117,N_3993,N_3944);
nand U4118 (N_4118,N_3916,N_3972);
nand U4119 (N_4119,N_3986,N_3971);
nand U4120 (N_4120,N_3982,N_3943);
or U4121 (N_4121,N_3957,N_3997);
and U4122 (N_4122,N_3937,N_3970);
or U4123 (N_4123,N_3997,N_3993);
nand U4124 (N_4124,N_3876,N_3891);
nor U4125 (N_4125,N_4085,N_4113);
nand U4126 (N_4126,N_4046,N_4124);
nand U4127 (N_4127,N_4123,N_4099);
and U4128 (N_4128,N_4116,N_4080);
nand U4129 (N_4129,N_4087,N_4010);
or U4130 (N_4130,N_4047,N_4031);
or U4131 (N_4131,N_4062,N_4039);
and U4132 (N_4132,N_4083,N_4088);
nand U4133 (N_4133,N_4106,N_4096);
or U4134 (N_4134,N_4108,N_4120);
or U4135 (N_4135,N_4001,N_4064);
nand U4136 (N_4136,N_4063,N_4110);
nand U4137 (N_4137,N_4078,N_4050);
and U4138 (N_4138,N_4075,N_4025);
nor U4139 (N_4139,N_4042,N_4024);
xnor U4140 (N_4140,N_4081,N_4054);
xnor U4141 (N_4141,N_4100,N_4015);
xor U4142 (N_4142,N_4014,N_4037);
nor U4143 (N_4143,N_4053,N_4018);
nand U4144 (N_4144,N_4057,N_4027);
nand U4145 (N_4145,N_4105,N_4118);
or U4146 (N_4146,N_4082,N_4104);
and U4147 (N_4147,N_4058,N_4000);
and U4148 (N_4148,N_4077,N_4070);
nand U4149 (N_4149,N_4056,N_4011);
or U4150 (N_4150,N_4065,N_4045);
nor U4151 (N_4151,N_4119,N_4003);
and U4152 (N_4152,N_4028,N_4035);
xnor U4153 (N_4153,N_4049,N_4048);
or U4154 (N_4154,N_4074,N_4115);
xor U4155 (N_4155,N_4095,N_4122);
or U4156 (N_4156,N_4036,N_4098);
nor U4157 (N_4157,N_4006,N_4112);
nand U4158 (N_4158,N_4060,N_4067);
nand U4159 (N_4159,N_4101,N_4068);
or U4160 (N_4160,N_4093,N_4023);
xor U4161 (N_4161,N_4051,N_4090);
or U4162 (N_4162,N_4019,N_4026);
nand U4163 (N_4163,N_4002,N_4071);
or U4164 (N_4164,N_4016,N_4069);
nand U4165 (N_4165,N_4091,N_4079);
or U4166 (N_4166,N_4044,N_4117);
and U4167 (N_4167,N_4041,N_4020);
and U4168 (N_4168,N_4030,N_4114);
and U4169 (N_4169,N_4107,N_4009);
xnor U4170 (N_4170,N_4086,N_4038);
nand U4171 (N_4171,N_4059,N_4032);
and U4172 (N_4172,N_4109,N_4040);
or U4173 (N_4173,N_4111,N_4097);
or U4174 (N_4174,N_4017,N_4034);
xnor U4175 (N_4175,N_4092,N_4052);
xnor U4176 (N_4176,N_4033,N_4007);
nand U4177 (N_4177,N_4089,N_4103);
xor U4178 (N_4178,N_4043,N_4073);
and U4179 (N_4179,N_4021,N_4061);
nand U4180 (N_4180,N_4029,N_4072);
or U4181 (N_4181,N_4102,N_4084);
or U4182 (N_4182,N_4008,N_4066);
or U4183 (N_4183,N_4013,N_4005);
nand U4184 (N_4184,N_4094,N_4012);
and U4185 (N_4185,N_4076,N_4022);
nor U4186 (N_4186,N_4004,N_4121);
nand U4187 (N_4187,N_4055,N_4011);
or U4188 (N_4188,N_4116,N_4083);
or U4189 (N_4189,N_4094,N_4069);
nand U4190 (N_4190,N_4030,N_4111);
and U4191 (N_4191,N_4037,N_4109);
xnor U4192 (N_4192,N_4117,N_4074);
and U4193 (N_4193,N_4003,N_4088);
or U4194 (N_4194,N_4058,N_4014);
xor U4195 (N_4195,N_4013,N_4065);
nand U4196 (N_4196,N_4037,N_4006);
nand U4197 (N_4197,N_4015,N_4088);
or U4198 (N_4198,N_4048,N_4082);
xor U4199 (N_4199,N_4090,N_4076);
and U4200 (N_4200,N_4015,N_4095);
and U4201 (N_4201,N_4114,N_4001);
nand U4202 (N_4202,N_4038,N_4098);
nand U4203 (N_4203,N_4025,N_4087);
nor U4204 (N_4204,N_4092,N_4116);
nand U4205 (N_4205,N_4076,N_4062);
nor U4206 (N_4206,N_4092,N_4023);
or U4207 (N_4207,N_4017,N_4043);
and U4208 (N_4208,N_4044,N_4082);
nand U4209 (N_4209,N_4003,N_4064);
xnor U4210 (N_4210,N_4044,N_4077);
nor U4211 (N_4211,N_4122,N_4002);
nor U4212 (N_4212,N_4078,N_4072);
or U4213 (N_4213,N_4033,N_4035);
or U4214 (N_4214,N_4007,N_4055);
nor U4215 (N_4215,N_4077,N_4042);
or U4216 (N_4216,N_4090,N_4109);
xor U4217 (N_4217,N_4060,N_4076);
and U4218 (N_4218,N_4057,N_4087);
nand U4219 (N_4219,N_4029,N_4057);
xnor U4220 (N_4220,N_4045,N_4060);
and U4221 (N_4221,N_4054,N_4118);
nand U4222 (N_4222,N_4086,N_4082);
or U4223 (N_4223,N_4102,N_4109);
nand U4224 (N_4224,N_4003,N_4104);
nor U4225 (N_4225,N_4065,N_4110);
or U4226 (N_4226,N_4006,N_4109);
nand U4227 (N_4227,N_4074,N_4034);
and U4228 (N_4228,N_4110,N_4028);
and U4229 (N_4229,N_4089,N_4009);
nand U4230 (N_4230,N_4084,N_4077);
and U4231 (N_4231,N_4014,N_4089);
xor U4232 (N_4232,N_4105,N_4052);
or U4233 (N_4233,N_4058,N_4036);
nand U4234 (N_4234,N_4068,N_4067);
nor U4235 (N_4235,N_4073,N_4022);
nor U4236 (N_4236,N_4026,N_4011);
nor U4237 (N_4237,N_4092,N_4053);
nor U4238 (N_4238,N_4067,N_4028);
xor U4239 (N_4239,N_4011,N_4069);
or U4240 (N_4240,N_4051,N_4095);
nand U4241 (N_4241,N_4031,N_4119);
xor U4242 (N_4242,N_4074,N_4061);
nor U4243 (N_4243,N_4026,N_4124);
nand U4244 (N_4244,N_4090,N_4002);
and U4245 (N_4245,N_4018,N_4019);
nand U4246 (N_4246,N_4118,N_4056);
nor U4247 (N_4247,N_4016,N_4120);
nand U4248 (N_4248,N_4052,N_4104);
nor U4249 (N_4249,N_4080,N_4107);
nor U4250 (N_4250,N_4153,N_4172);
and U4251 (N_4251,N_4205,N_4226);
nand U4252 (N_4252,N_4154,N_4136);
nor U4253 (N_4253,N_4176,N_4239);
or U4254 (N_4254,N_4178,N_4249);
nor U4255 (N_4255,N_4131,N_4248);
nor U4256 (N_4256,N_4175,N_4158);
nor U4257 (N_4257,N_4219,N_4189);
nor U4258 (N_4258,N_4214,N_4220);
or U4259 (N_4259,N_4213,N_4245);
nand U4260 (N_4260,N_4177,N_4225);
or U4261 (N_4261,N_4128,N_4144);
and U4262 (N_4262,N_4148,N_4167);
or U4263 (N_4263,N_4199,N_4206);
or U4264 (N_4264,N_4203,N_4138);
or U4265 (N_4265,N_4193,N_4221);
xor U4266 (N_4266,N_4149,N_4146);
and U4267 (N_4267,N_4160,N_4223);
nand U4268 (N_4268,N_4192,N_4209);
or U4269 (N_4269,N_4156,N_4164);
or U4270 (N_4270,N_4182,N_4165);
nor U4271 (N_4271,N_4191,N_4186);
or U4272 (N_4272,N_4162,N_4130);
nor U4273 (N_4273,N_4137,N_4159);
nand U4274 (N_4274,N_4227,N_4125);
or U4275 (N_4275,N_4196,N_4126);
and U4276 (N_4276,N_4210,N_4218);
nor U4277 (N_4277,N_4217,N_4180);
nor U4278 (N_4278,N_4234,N_4173);
xor U4279 (N_4279,N_4151,N_4197);
or U4280 (N_4280,N_4169,N_4238);
nor U4281 (N_4281,N_4201,N_4184);
nor U4282 (N_4282,N_4155,N_4204);
nor U4283 (N_4283,N_4129,N_4194);
and U4284 (N_4284,N_4211,N_4171);
nand U4285 (N_4285,N_4202,N_4187);
or U4286 (N_4286,N_4142,N_4215);
nor U4287 (N_4287,N_4232,N_4229);
nand U4288 (N_4288,N_4163,N_4200);
and U4289 (N_4289,N_4152,N_4216);
nand U4290 (N_4290,N_4185,N_4243);
xor U4291 (N_4291,N_4222,N_4140);
nor U4292 (N_4292,N_4179,N_4127);
nor U4293 (N_4293,N_4190,N_4139);
nor U4294 (N_4294,N_4242,N_4170);
xnor U4295 (N_4295,N_4166,N_4241);
and U4296 (N_4296,N_4198,N_4181);
nand U4297 (N_4297,N_4134,N_4133);
nor U4298 (N_4298,N_4228,N_4208);
and U4299 (N_4299,N_4240,N_4247);
and U4300 (N_4300,N_4145,N_4147);
xor U4301 (N_4301,N_4150,N_4244);
or U4302 (N_4302,N_4183,N_4168);
xor U4303 (N_4303,N_4224,N_4143);
and U4304 (N_4304,N_4246,N_4141);
xor U4305 (N_4305,N_4230,N_4195);
xor U4306 (N_4306,N_4236,N_4157);
xnor U4307 (N_4307,N_4231,N_4132);
xor U4308 (N_4308,N_4207,N_4235);
nand U4309 (N_4309,N_4174,N_4161);
and U4310 (N_4310,N_4237,N_4188);
or U4311 (N_4311,N_4233,N_4135);
nand U4312 (N_4312,N_4212,N_4201);
nor U4313 (N_4313,N_4217,N_4244);
and U4314 (N_4314,N_4217,N_4233);
nand U4315 (N_4315,N_4182,N_4132);
or U4316 (N_4316,N_4161,N_4164);
and U4317 (N_4317,N_4179,N_4183);
nor U4318 (N_4318,N_4235,N_4171);
and U4319 (N_4319,N_4225,N_4148);
and U4320 (N_4320,N_4131,N_4178);
nand U4321 (N_4321,N_4240,N_4150);
xnor U4322 (N_4322,N_4240,N_4213);
xnor U4323 (N_4323,N_4227,N_4204);
or U4324 (N_4324,N_4204,N_4239);
or U4325 (N_4325,N_4127,N_4182);
and U4326 (N_4326,N_4129,N_4177);
and U4327 (N_4327,N_4139,N_4155);
and U4328 (N_4328,N_4169,N_4214);
or U4329 (N_4329,N_4241,N_4239);
or U4330 (N_4330,N_4126,N_4132);
or U4331 (N_4331,N_4190,N_4211);
nand U4332 (N_4332,N_4145,N_4191);
nand U4333 (N_4333,N_4131,N_4168);
xnor U4334 (N_4334,N_4178,N_4165);
nor U4335 (N_4335,N_4189,N_4129);
xnor U4336 (N_4336,N_4186,N_4193);
and U4337 (N_4337,N_4229,N_4212);
or U4338 (N_4338,N_4201,N_4218);
or U4339 (N_4339,N_4216,N_4132);
xor U4340 (N_4340,N_4133,N_4212);
xor U4341 (N_4341,N_4239,N_4135);
nor U4342 (N_4342,N_4241,N_4188);
nand U4343 (N_4343,N_4227,N_4221);
xor U4344 (N_4344,N_4198,N_4137);
and U4345 (N_4345,N_4216,N_4206);
or U4346 (N_4346,N_4130,N_4176);
and U4347 (N_4347,N_4172,N_4218);
and U4348 (N_4348,N_4220,N_4249);
and U4349 (N_4349,N_4158,N_4126);
xor U4350 (N_4350,N_4179,N_4235);
and U4351 (N_4351,N_4145,N_4195);
or U4352 (N_4352,N_4212,N_4164);
nand U4353 (N_4353,N_4203,N_4195);
nor U4354 (N_4354,N_4145,N_4192);
nor U4355 (N_4355,N_4177,N_4220);
nand U4356 (N_4356,N_4232,N_4130);
xor U4357 (N_4357,N_4230,N_4131);
and U4358 (N_4358,N_4188,N_4129);
nand U4359 (N_4359,N_4227,N_4214);
nand U4360 (N_4360,N_4174,N_4152);
xnor U4361 (N_4361,N_4193,N_4200);
xor U4362 (N_4362,N_4202,N_4183);
xnor U4363 (N_4363,N_4192,N_4198);
nand U4364 (N_4364,N_4241,N_4181);
or U4365 (N_4365,N_4191,N_4217);
xor U4366 (N_4366,N_4166,N_4149);
nor U4367 (N_4367,N_4154,N_4162);
and U4368 (N_4368,N_4220,N_4142);
or U4369 (N_4369,N_4241,N_4204);
nand U4370 (N_4370,N_4195,N_4196);
or U4371 (N_4371,N_4183,N_4186);
nor U4372 (N_4372,N_4242,N_4190);
nor U4373 (N_4373,N_4134,N_4207);
xor U4374 (N_4374,N_4151,N_4176);
or U4375 (N_4375,N_4316,N_4299);
nor U4376 (N_4376,N_4341,N_4323);
nor U4377 (N_4377,N_4282,N_4296);
xnor U4378 (N_4378,N_4365,N_4285);
xnor U4379 (N_4379,N_4287,N_4342);
nor U4380 (N_4380,N_4300,N_4340);
nand U4381 (N_4381,N_4356,N_4336);
xor U4382 (N_4382,N_4346,N_4324);
or U4383 (N_4383,N_4368,N_4253);
nand U4384 (N_4384,N_4322,N_4364);
nand U4385 (N_4385,N_4349,N_4267);
and U4386 (N_4386,N_4259,N_4367);
or U4387 (N_4387,N_4284,N_4250);
and U4388 (N_4388,N_4289,N_4317);
and U4389 (N_4389,N_4274,N_4312);
and U4390 (N_4390,N_4278,N_4273);
or U4391 (N_4391,N_4361,N_4291);
nand U4392 (N_4392,N_4372,N_4254);
or U4393 (N_4393,N_4286,N_4281);
and U4394 (N_4394,N_4327,N_4351);
xor U4395 (N_4395,N_4301,N_4307);
nor U4396 (N_4396,N_4309,N_4359);
or U4397 (N_4397,N_4329,N_4318);
nand U4398 (N_4398,N_4306,N_4256);
nor U4399 (N_4399,N_4298,N_4353);
and U4400 (N_4400,N_4295,N_4339);
nand U4401 (N_4401,N_4268,N_4263);
nor U4402 (N_4402,N_4333,N_4314);
or U4403 (N_4403,N_4347,N_4310);
and U4404 (N_4404,N_4370,N_4362);
nand U4405 (N_4405,N_4338,N_4252);
xor U4406 (N_4406,N_4270,N_4311);
xor U4407 (N_4407,N_4315,N_4290);
and U4408 (N_4408,N_4257,N_4343);
nor U4409 (N_4409,N_4305,N_4369);
or U4410 (N_4410,N_4292,N_4345);
nor U4411 (N_4411,N_4261,N_4374);
and U4412 (N_4412,N_4303,N_4355);
or U4413 (N_4413,N_4262,N_4265);
and U4414 (N_4414,N_4266,N_4288);
nand U4415 (N_4415,N_4371,N_4308);
xnor U4416 (N_4416,N_4330,N_4373);
nor U4417 (N_4417,N_4255,N_4337);
and U4418 (N_4418,N_4276,N_4320);
nand U4419 (N_4419,N_4334,N_4304);
or U4420 (N_4420,N_4350,N_4366);
and U4421 (N_4421,N_4272,N_4352);
nand U4422 (N_4422,N_4269,N_4332);
nand U4423 (N_4423,N_4313,N_4360);
or U4424 (N_4424,N_4319,N_4335);
and U4425 (N_4425,N_4251,N_4325);
xnor U4426 (N_4426,N_4321,N_4280);
or U4427 (N_4427,N_4326,N_4294);
xnor U4428 (N_4428,N_4264,N_4275);
or U4429 (N_4429,N_4358,N_4344);
nor U4430 (N_4430,N_4297,N_4357);
and U4431 (N_4431,N_4283,N_4260);
and U4432 (N_4432,N_4363,N_4331);
xnor U4433 (N_4433,N_4354,N_4302);
xnor U4434 (N_4434,N_4293,N_4348);
nand U4435 (N_4435,N_4277,N_4258);
xnor U4436 (N_4436,N_4271,N_4328);
xor U4437 (N_4437,N_4279,N_4360);
nor U4438 (N_4438,N_4317,N_4276);
nor U4439 (N_4439,N_4311,N_4259);
nand U4440 (N_4440,N_4362,N_4306);
nor U4441 (N_4441,N_4349,N_4345);
and U4442 (N_4442,N_4362,N_4295);
xnor U4443 (N_4443,N_4374,N_4275);
nor U4444 (N_4444,N_4323,N_4363);
xnor U4445 (N_4445,N_4305,N_4258);
or U4446 (N_4446,N_4314,N_4341);
or U4447 (N_4447,N_4310,N_4358);
or U4448 (N_4448,N_4299,N_4267);
nor U4449 (N_4449,N_4347,N_4262);
nor U4450 (N_4450,N_4300,N_4324);
xor U4451 (N_4451,N_4353,N_4288);
xor U4452 (N_4452,N_4267,N_4305);
nand U4453 (N_4453,N_4329,N_4312);
nand U4454 (N_4454,N_4271,N_4373);
nand U4455 (N_4455,N_4297,N_4374);
and U4456 (N_4456,N_4357,N_4324);
xnor U4457 (N_4457,N_4343,N_4272);
and U4458 (N_4458,N_4347,N_4323);
and U4459 (N_4459,N_4309,N_4304);
nand U4460 (N_4460,N_4258,N_4367);
and U4461 (N_4461,N_4361,N_4285);
xnor U4462 (N_4462,N_4318,N_4288);
and U4463 (N_4463,N_4276,N_4272);
or U4464 (N_4464,N_4285,N_4316);
nand U4465 (N_4465,N_4351,N_4296);
xor U4466 (N_4466,N_4318,N_4272);
nor U4467 (N_4467,N_4343,N_4317);
xor U4468 (N_4468,N_4364,N_4273);
and U4469 (N_4469,N_4316,N_4261);
or U4470 (N_4470,N_4337,N_4316);
nor U4471 (N_4471,N_4305,N_4279);
nor U4472 (N_4472,N_4283,N_4341);
nand U4473 (N_4473,N_4317,N_4332);
xnor U4474 (N_4474,N_4364,N_4325);
nor U4475 (N_4475,N_4323,N_4300);
and U4476 (N_4476,N_4323,N_4333);
and U4477 (N_4477,N_4271,N_4306);
or U4478 (N_4478,N_4325,N_4254);
xnor U4479 (N_4479,N_4279,N_4264);
xor U4480 (N_4480,N_4260,N_4352);
or U4481 (N_4481,N_4269,N_4279);
nand U4482 (N_4482,N_4318,N_4353);
nand U4483 (N_4483,N_4292,N_4294);
xnor U4484 (N_4484,N_4320,N_4329);
xor U4485 (N_4485,N_4371,N_4251);
nand U4486 (N_4486,N_4258,N_4283);
and U4487 (N_4487,N_4334,N_4343);
nand U4488 (N_4488,N_4289,N_4266);
or U4489 (N_4489,N_4356,N_4291);
nand U4490 (N_4490,N_4301,N_4308);
or U4491 (N_4491,N_4319,N_4311);
nor U4492 (N_4492,N_4319,N_4361);
or U4493 (N_4493,N_4346,N_4334);
nor U4494 (N_4494,N_4351,N_4322);
nor U4495 (N_4495,N_4265,N_4295);
xor U4496 (N_4496,N_4345,N_4290);
xor U4497 (N_4497,N_4371,N_4285);
and U4498 (N_4498,N_4306,N_4373);
and U4499 (N_4499,N_4253,N_4328);
and U4500 (N_4500,N_4424,N_4416);
or U4501 (N_4501,N_4482,N_4375);
or U4502 (N_4502,N_4390,N_4477);
and U4503 (N_4503,N_4441,N_4442);
nor U4504 (N_4504,N_4458,N_4401);
nor U4505 (N_4505,N_4462,N_4413);
nand U4506 (N_4506,N_4376,N_4403);
nand U4507 (N_4507,N_4410,N_4436);
nand U4508 (N_4508,N_4417,N_4430);
or U4509 (N_4509,N_4412,N_4396);
and U4510 (N_4510,N_4421,N_4463);
nor U4511 (N_4511,N_4464,N_4400);
xor U4512 (N_4512,N_4415,N_4404);
or U4513 (N_4513,N_4382,N_4378);
xnor U4514 (N_4514,N_4499,N_4449);
nand U4515 (N_4515,N_4438,N_4440);
xnor U4516 (N_4516,N_4447,N_4484);
or U4517 (N_4517,N_4381,N_4422);
xor U4518 (N_4518,N_4460,N_4418);
and U4519 (N_4519,N_4445,N_4393);
and U4520 (N_4520,N_4471,N_4470);
nand U4521 (N_4521,N_4383,N_4397);
xor U4522 (N_4522,N_4443,N_4489);
xnor U4523 (N_4523,N_4459,N_4455);
nand U4524 (N_4524,N_4461,N_4486);
nand U4525 (N_4525,N_4432,N_4429);
and U4526 (N_4526,N_4474,N_4481);
or U4527 (N_4527,N_4495,N_4392);
xnor U4528 (N_4528,N_4398,N_4423);
or U4529 (N_4529,N_4439,N_4387);
nor U4530 (N_4530,N_4468,N_4479);
nand U4531 (N_4531,N_4420,N_4395);
and U4532 (N_4532,N_4409,N_4427);
nor U4533 (N_4533,N_4466,N_4444);
xnor U4534 (N_4534,N_4496,N_4431);
nand U4535 (N_4535,N_4433,N_4483);
nor U4536 (N_4536,N_4475,N_4467);
xnor U4537 (N_4537,N_4388,N_4485);
and U4538 (N_4538,N_4446,N_4469);
and U4539 (N_4539,N_4428,N_4407);
xor U4540 (N_4540,N_4419,N_4498);
or U4541 (N_4541,N_4384,N_4472);
or U4542 (N_4542,N_4448,N_4389);
nand U4543 (N_4543,N_4478,N_4406);
nand U4544 (N_4544,N_4377,N_4488);
and U4545 (N_4545,N_4476,N_4402);
nor U4546 (N_4546,N_4451,N_4490);
and U4547 (N_4547,N_4452,N_4487);
xnor U4548 (N_4548,N_4497,N_4456);
nand U4549 (N_4549,N_4493,N_4385);
and U4550 (N_4550,N_4454,N_4492);
xor U4551 (N_4551,N_4457,N_4411);
nand U4552 (N_4552,N_4414,N_4426);
or U4553 (N_4553,N_4425,N_4450);
or U4554 (N_4554,N_4408,N_4465);
and U4555 (N_4555,N_4435,N_4473);
and U4556 (N_4556,N_4379,N_4394);
and U4557 (N_4557,N_4494,N_4391);
xnor U4558 (N_4558,N_4405,N_4386);
nor U4559 (N_4559,N_4399,N_4380);
or U4560 (N_4560,N_4434,N_4437);
nor U4561 (N_4561,N_4453,N_4491);
nand U4562 (N_4562,N_4480,N_4449);
or U4563 (N_4563,N_4452,N_4446);
nor U4564 (N_4564,N_4408,N_4457);
and U4565 (N_4565,N_4466,N_4462);
and U4566 (N_4566,N_4405,N_4430);
nand U4567 (N_4567,N_4417,N_4454);
nand U4568 (N_4568,N_4393,N_4387);
xor U4569 (N_4569,N_4481,N_4429);
nor U4570 (N_4570,N_4409,N_4464);
nor U4571 (N_4571,N_4470,N_4382);
and U4572 (N_4572,N_4459,N_4386);
or U4573 (N_4573,N_4464,N_4455);
and U4574 (N_4574,N_4460,N_4405);
and U4575 (N_4575,N_4409,N_4389);
nor U4576 (N_4576,N_4488,N_4404);
nor U4577 (N_4577,N_4420,N_4403);
xor U4578 (N_4578,N_4463,N_4474);
and U4579 (N_4579,N_4462,N_4409);
nor U4580 (N_4580,N_4424,N_4423);
and U4581 (N_4581,N_4455,N_4466);
or U4582 (N_4582,N_4483,N_4497);
nand U4583 (N_4583,N_4475,N_4471);
nor U4584 (N_4584,N_4499,N_4491);
or U4585 (N_4585,N_4411,N_4387);
nor U4586 (N_4586,N_4425,N_4415);
xnor U4587 (N_4587,N_4405,N_4453);
nor U4588 (N_4588,N_4494,N_4422);
or U4589 (N_4589,N_4441,N_4377);
or U4590 (N_4590,N_4420,N_4499);
nand U4591 (N_4591,N_4460,N_4388);
xor U4592 (N_4592,N_4458,N_4441);
or U4593 (N_4593,N_4396,N_4465);
xnor U4594 (N_4594,N_4377,N_4405);
nor U4595 (N_4595,N_4426,N_4421);
nand U4596 (N_4596,N_4395,N_4412);
nor U4597 (N_4597,N_4459,N_4468);
and U4598 (N_4598,N_4444,N_4426);
nor U4599 (N_4599,N_4435,N_4464);
xnor U4600 (N_4600,N_4452,N_4433);
or U4601 (N_4601,N_4459,N_4479);
or U4602 (N_4602,N_4494,N_4386);
or U4603 (N_4603,N_4425,N_4409);
and U4604 (N_4604,N_4379,N_4493);
nor U4605 (N_4605,N_4403,N_4382);
nand U4606 (N_4606,N_4489,N_4415);
nor U4607 (N_4607,N_4377,N_4412);
nor U4608 (N_4608,N_4482,N_4415);
and U4609 (N_4609,N_4471,N_4379);
xor U4610 (N_4610,N_4425,N_4481);
and U4611 (N_4611,N_4426,N_4403);
and U4612 (N_4612,N_4436,N_4433);
xnor U4613 (N_4613,N_4392,N_4405);
xnor U4614 (N_4614,N_4496,N_4447);
or U4615 (N_4615,N_4493,N_4462);
and U4616 (N_4616,N_4408,N_4387);
or U4617 (N_4617,N_4451,N_4387);
or U4618 (N_4618,N_4393,N_4377);
and U4619 (N_4619,N_4415,N_4402);
nand U4620 (N_4620,N_4415,N_4432);
and U4621 (N_4621,N_4451,N_4384);
nand U4622 (N_4622,N_4483,N_4398);
and U4623 (N_4623,N_4384,N_4417);
nand U4624 (N_4624,N_4494,N_4461);
xnor U4625 (N_4625,N_4569,N_4536);
and U4626 (N_4626,N_4600,N_4567);
xnor U4627 (N_4627,N_4509,N_4609);
and U4628 (N_4628,N_4576,N_4563);
or U4629 (N_4629,N_4546,N_4544);
and U4630 (N_4630,N_4606,N_4585);
or U4631 (N_4631,N_4610,N_4568);
xnor U4632 (N_4632,N_4594,N_4511);
xor U4633 (N_4633,N_4512,N_4557);
xor U4634 (N_4634,N_4526,N_4503);
or U4635 (N_4635,N_4501,N_4547);
and U4636 (N_4636,N_4597,N_4518);
nor U4637 (N_4637,N_4564,N_4616);
nand U4638 (N_4638,N_4588,N_4506);
and U4639 (N_4639,N_4566,N_4595);
or U4640 (N_4640,N_4604,N_4577);
nor U4641 (N_4641,N_4525,N_4592);
or U4642 (N_4642,N_4502,N_4580);
or U4643 (N_4643,N_4589,N_4559);
xor U4644 (N_4644,N_4558,N_4510);
and U4645 (N_4645,N_4578,N_4619);
or U4646 (N_4646,N_4534,N_4527);
nor U4647 (N_4647,N_4605,N_4504);
and U4648 (N_4648,N_4602,N_4621);
nor U4649 (N_4649,N_4554,N_4521);
xor U4650 (N_4650,N_4593,N_4551);
nand U4651 (N_4651,N_4607,N_4520);
nand U4652 (N_4652,N_4515,N_4587);
or U4653 (N_4653,N_4516,N_4565);
nor U4654 (N_4654,N_4591,N_4620);
nor U4655 (N_4655,N_4507,N_4601);
or U4656 (N_4656,N_4505,N_4541);
xnor U4657 (N_4657,N_4524,N_4533);
nand U4658 (N_4658,N_4582,N_4537);
and U4659 (N_4659,N_4613,N_4530);
and U4660 (N_4660,N_4519,N_4535);
nor U4661 (N_4661,N_4561,N_4560);
nor U4662 (N_4662,N_4514,N_4548);
and U4663 (N_4663,N_4523,N_4513);
nand U4664 (N_4664,N_4624,N_4603);
xor U4665 (N_4665,N_4539,N_4581);
nand U4666 (N_4666,N_4579,N_4612);
xnor U4667 (N_4667,N_4555,N_4584);
nand U4668 (N_4668,N_4552,N_4583);
and U4669 (N_4669,N_4542,N_4622);
or U4670 (N_4670,N_4528,N_4517);
and U4671 (N_4671,N_4573,N_4545);
nand U4672 (N_4672,N_4615,N_4574);
nand U4673 (N_4673,N_4556,N_4531);
nor U4674 (N_4674,N_4586,N_4572);
or U4675 (N_4675,N_4590,N_4614);
and U4676 (N_4676,N_4623,N_4538);
or U4677 (N_4677,N_4529,N_4618);
xnor U4678 (N_4678,N_4550,N_4540);
and U4679 (N_4679,N_4508,N_4532);
or U4680 (N_4680,N_4553,N_4500);
nand U4681 (N_4681,N_4570,N_4617);
nor U4682 (N_4682,N_4598,N_4562);
nor U4683 (N_4683,N_4608,N_4611);
nand U4684 (N_4684,N_4543,N_4575);
xor U4685 (N_4685,N_4596,N_4571);
nand U4686 (N_4686,N_4549,N_4599);
xor U4687 (N_4687,N_4522,N_4528);
xor U4688 (N_4688,N_4546,N_4537);
or U4689 (N_4689,N_4549,N_4525);
nand U4690 (N_4690,N_4558,N_4542);
and U4691 (N_4691,N_4547,N_4614);
xnor U4692 (N_4692,N_4543,N_4513);
nor U4693 (N_4693,N_4569,N_4599);
xor U4694 (N_4694,N_4537,N_4549);
nor U4695 (N_4695,N_4542,N_4562);
or U4696 (N_4696,N_4621,N_4581);
and U4697 (N_4697,N_4513,N_4615);
xor U4698 (N_4698,N_4611,N_4583);
or U4699 (N_4699,N_4561,N_4501);
nand U4700 (N_4700,N_4539,N_4511);
or U4701 (N_4701,N_4525,N_4580);
or U4702 (N_4702,N_4609,N_4619);
nand U4703 (N_4703,N_4568,N_4591);
nand U4704 (N_4704,N_4526,N_4582);
nor U4705 (N_4705,N_4578,N_4555);
or U4706 (N_4706,N_4547,N_4596);
and U4707 (N_4707,N_4531,N_4553);
nand U4708 (N_4708,N_4576,N_4615);
and U4709 (N_4709,N_4590,N_4528);
and U4710 (N_4710,N_4517,N_4549);
nor U4711 (N_4711,N_4593,N_4582);
nand U4712 (N_4712,N_4509,N_4546);
nand U4713 (N_4713,N_4573,N_4547);
and U4714 (N_4714,N_4543,N_4614);
xor U4715 (N_4715,N_4558,N_4617);
and U4716 (N_4716,N_4527,N_4610);
nor U4717 (N_4717,N_4507,N_4558);
or U4718 (N_4718,N_4579,N_4519);
nor U4719 (N_4719,N_4556,N_4564);
or U4720 (N_4720,N_4503,N_4524);
nor U4721 (N_4721,N_4522,N_4607);
and U4722 (N_4722,N_4500,N_4524);
or U4723 (N_4723,N_4507,N_4570);
nor U4724 (N_4724,N_4555,N_4553);
and U4725 (N_4725,N_4505,N_4549);
and U4726 (N_4726,N_4507,N_4503);
nor U4727 (N_4727,N_4621,N_4503);
or U4728 (N_4728,N_4596,N_4569);
and U4729 (N_4729,N_4577,N_4622);
xnor U4730 (N_4730,N_4578,N_4515);
nand U4731 (N_4731,N_4557,N_4537);
nor U4732 (N_4732,N_4516,N_4572);
nor U4733 (N_4733,N_4575,N_4523);
and U4734 (N_4734,N_4589,N_4597);
xnor U4735 (N_4735,N_4558,N_4578);
and U4736 (N_4736,N_4532,N_4619);
nand U4737 (N_4737,N_4522,N_4592);
or U4738 (N_4738,N_4605,N_4542);
nand U4739 (N_4739,N_4573,N_4567);
or U4740 (N_4740,N_4604,N_4576);
nor U4741 (N_4741,N_4567,N_4596);
nand U4742 (N_4742,N_4535,N_4500);
or U4743 (N_4743,N_4578,N_4540);
or U4744 (N_4744,N_4514,N_4601);
or U4745 (N_4745,N_4514,N_4609);
or U4746 (N_4746,N_4511,N_4503);
or U4747 (N_4747,N_4541,N_4504);
and U4748 (N_4748,N_4527,N_4620);
and U4749 (N_4749,N_4585,N_4560);
nand U4750 (N_4750,N_4745,N_4736);
nand U4751 (N_4751,N_4705,N_4634);
or U4752 (N_4752,N_4711,N_4749);
or U4753 (N_4753,N_4628,N_4656);
xor U4754 (N_4754,N_4658,N_4670);
or U4755 (N_4755,N_4723,N_4715);
nor U4756 (N_4756,N_4709,N_4689);
and U4757 (N_4757,N_4669,N_4686);
and U4758 (N_4758,N_4662,N_4676);
xnor U4759 (N_4759,N_4635,N_4639);
xor U4760 (N_4760,N_4666,N_4701);
and U4761 (N_4761,N_4722,N_4719);
nand U4762 (N_4762,N_4668,N_4743);
and U4763 (N_4763,N_4744,N_4721);
nor U4764 (N_4764,N_4648,N_4657);
and U4765 (N_4765,N_4644,N_4702);
nor U4766 (N_4766,N_4684,N_4699);
and U4767 (N_4767,N_4692,N_4659);
and U4768 (N_4768,N_4626,N_4728);
xnor U4769 (N_4769,N_4643,N_4718);
xnor U4770 (N_4770,N_4695,N_4698);
nor U4771 (N_4771,N_4690,N_4714);
xor U4772 (N_4772,N_4683,N_4737);
and U4773 (N_4773,N_4724,N_4694);
or U4774 (N_4774,N_4627,N_4703);
or U4775 (N_4775,N_4716,N_4679);
nor U4776 (N_4776,N_4733,N_4674);
or U4777 (N_4777,N_4681,N_4673);
and U4778 (N_4778,N_4739,N_4665);
xnor U4779 (N_4779,N_4660,N_4691);
nand U4780 (N_4780,N_4667,N_4636);
nor U4781 (N_4781,N_4740,N_4672);
nand U4782 (N_4782,N_4712,N_4649);
xnor U4783 (N_4783,N_4647,N_4706);
nor U4784 (N_4784,N_4640,N_4677);
nand U4785 (N_4785,N_4687,N_4642);
nand U4786 (N_4786,N_4688,N_4731);
and U4787 (N_4787,N_4654,N_4717);
or U4788 (N_4788,N_4704,N_4638);
xor U4789 (N_4789,N_4713,N_4707);
and U4790 (N_4790,N_4664,N_4645);
or U4791 (N_4791,N_4675,N_4742);
nor U4792 (N_4792,N_4726,N_4631);
or U4793 (N_4793,N_4735,N_4637);
xor U4794 (N_4794,N_4653,N_4732);
nor U4795 (N_4795,N_4748,N_4729);
and U4796 (N_4796,N_4685,N_4746);
and U4797 (N_4797,N_4720,N_4629);
nor U4798 (N_4798,N_4734,N_4747);
xnor U4799 (N_4799,N_4655,N_4652);
xnor U4800 (N_4800,N_4663,N_4680);
nand U4801 (N_4801,N_4625,N_4633);
or U4802 (N_4802,N_4682,N_4741);
nand U4803 (N_4803,N_4700,N_4727);
nand U4804 (N_4804,N_4678,N_4651);
and U4805 (N_4805,N_4632,N_4641);
nor U4806 (N_4806,N_4650,N_4710);
and U4807 (N_4807,N_4738,N_4646);
nand U4808 (N_4808,N_4708,N_4671);
xnor U4809 (N_4809,N_4630,N_4730);
xor U4810 (N_4810,N_4661,N_4693);
and U4811 (N_4811,N_4725,N_4696);
xor U4812 (N_4812,N_4697,N_4711);
nor U4813 (N_4813,N_4714,N_4672);
xor U4814 (N_4814,N_4736,N_4694);
and U4815 (N_4815,N_4715,N_4661);
and U4816 (N_4816,N_4684,N_4670);
or U4817 (N_4817,N_4686,N_4677);
xor U4818 (N_4818,N_4721,N_4748);
xnor U4819 (N_4819,N_4713,N_4704);
and U4820 (N_4820,N_4729,N_4675);
and U4821 (N_4821,N_4656,N_4694);
and U4822 (N_4822,N_4648,N_4672);
xor U4823 (N_4823,N_4698,N_4666);
or U4824 (N_4824,N_4739,N_4740);
nand U4825 (N_4825,N_4640,N_4697);
nor U4826 (N_4826,N_4729,N_4646);
and U4827 (N_4827,N_4709,N_4681);
xor U4828 (N_4828,N_4696,N_4643);
nor U4829 (N_4829,N_4736,N_4692);
xnor U4830 (N_4830,N_4701,N_4721);
nor U4831 (N_4831,N_4707,N_4733);
nand U4832 (N_4832,N_4672,N_4662);
xor U4833 (N_4833,N_4697,N_4736);
and U4834 (N_4834,N_4648,N_4656);
xnor U4835 (N_4835,N_4659,N_4749);
or U4836 (N_4836,N_4726,N_4673);
xor U4837 (N_4837,N_4629,N_4651);
xnor U4838 (N_4838,N_4731,N_4692);
nor U4839 (N_4839,N_4677,N_4641);
or U4840 (N_4840,N_4731,N_4730);
or U4841 (N_4841,N_4686,N_4646);
xnor U4842 (N_4842,N_4697,N_4733);
nor U4843 (N_4843,N_4647,N_4638);
or U4844 (N_4844,N_4651,N_4687);
nor U4845 (N_4845,N_4706,N_4644);
nand U4846 (N_4846,N_4686,N_4651);
and U4847 (N_4847,N_4714,N_4727);
nand U4848 (N_4848,N_4628,N_4703);
or U4849 (N_4849,N_4701,N_4745);
xnor U4850 (N_4850,N_4708,N_4743);
nor U4851 (N_4851,N_4694,N_4667);
nor U4852 (N_4852,N_4642,N_4731);
or U4853 (N_4853,N_4748,N_4627);
nor U4854 (N_4854,N_4718,N_4637);
nand U4855 (N_4855,N_4631,N_4702);
nor U4856 (N_4856,N_4730,N_4715);
and U4857 (N_4857,N_4674,N_4661);
nor U4858 (N_4858,N_4699,N_4648);
nor U4859 (N_4859,N_4677,N_4718);
or U4860 (N_4860,N_4664,N_4699);
nor U4861 (N_4861,N_4682,N_4642);
nor U4862 (N_4862,N_4724,N_4656);
nor U4863 (N_4863,N_4748,N_4717);
nor U4864 (N_4864,N_4695,N_4688);
nand U4865 (N_4865,N_4743,N_4698);
nor U4866 (N_4866,N_4720,N_4679);
and U4867 (N_4867,N_4721,N_4708);
nor U4868 (N_4868,N_4698,N_4748);
nand U4869 (N_4869,N_4742,N_4625);
and U4870 (N_4870,N_4628,N_4707);
and U4871 (N_4871,N_4714,N_4687);
or U4872 (N_4872,N_4702,N_4706);
or U4873 (N_4873,N_4680,N_4668);
xnor U4874 (N_4874,N_4669,N_4659);
or U4875 (N_4875,N_4759,N_4800);
xor U4876 (N_4876,N_4751,N_4765);
nor U4877 (N_4877,N_4867,N_4784);
nand U4878 (N_4878,N_4860,N_4804);
and U4879 (N_4879,N_4874,N_4859);
xor U4880 (N_4880,N_4752,N_4866);
and U4881 (N_4881,N_4862,N_4848);
and U4882 (N_4882,N_4754,N_4826);
nand U4883 (N_4883,N_4810,N_4763);
nor U4884 (N_4884,N_4819,N_4834);
nor U4885 (N_4885,N_4824,N_4841);
nor U4886 (N_4886,N_4785,N_4787);
xnor U4887 (N_4887,N_4846,N_4766);
or U4888 (N_4888,N_4775,N_4870);
xor U4889 (N_4889,N_4780,N_4829);
and U4890 (N_4890,N_4840,N_4770);
nor U4891 (N_4891,N_4791,N_4811);
or U4892 (N_4892,N_4807,N_4816);
nor U4893 (N_4893,N_4798,N_4777);
xor U4894 (N_4894,N_4750,N_4845);
and U4895 (N_4895,N_4852,N_4842);
and U4896 (N_4896,N_4792,N_4851);
or U4897 (N_4897,N_4821,N_4818);
xnor U4898 (N_4898,N_4858,N_4795);
nor U4899 (N_4899,N_4864,N_4797);
xnor U4900 (N_4900,N_4831,N_4776);
or U4901 (N_4901,N_4758,N_4872);
xor U4902 (N_4902,N_4794,N_4806);
or U4903 (N_4903,N_4782,N_4772);
nor U4904 (N_4904,N_4769,N_4833);
and U4905 (N_4905,N_4760,N_4762);
or U4906 (N_4906,N_4786,N_4868);
xor U4907 (N_4907,N_4849,N_4828);
or U4908 (N_4908,N_4843,N_4788);
nor U4909 (N_4909,N_4790,N_4761);
xor U4910 (N_4910,N_4812,N_4757);
nand U4911 (N_4911,N_4844,N_4815);
or U4912 (N_4912,N_4767,N_4771);
nor U4913 (N_4913,N_4768,N_4817);
xor U4914 (N_4914,N_4820,N_4779);
xor U4915 (N_4915,N_4822,N_4789);
nand U4916 (N_4916,N_4753,N_4803);
nand U4917 (N_4917,N_4773,N_4814);
and U4918 (N_4918,N_4850,N_4847);
or U4919 (N_4919,N_4863,N_4796);
and U4920 (N_4920,N_4871,N_4793);
nand U4921 (N_4921,N_4854,N_4799);
xnor U4922 (N_4922,N_4805,N_4869);
nor U4923 (N_4923,N_4838,N_4755);
and U4924 (N_4924,N_4802,N_4778);
xnor U4925 (N_4925,N_4861,N_4801);
and U4926 (N_4926,N_4813,N_4823);
nand U4927 (N_4927,N_4783,N_4756);
nor U4928 (N_4928,N_4825,N_4830);
and U4929 (N_4929,N_4781,N_4835);
nor U4930 (N_4930,N_4808,N_4873);
or U4931 (N_4931,N_4809,N_4836);
and U4932 (N_4932,N_4827,N_4853);
nor U4933 (N_4933,N_4774,N_4837);
or U4934 (N_4934,N_4855,N_4764);
and U4935 (N_4935,N_4839,N_4832);
or U4936 (N_4936,N_4857,N_4856);
xnor U4937 (N_4937,N_4865,N_4752);
and U4938 (N_4938,N_4770,N_4794);
xor U4939 (N_4939,N_4825,N_4756);
nand U4940 (N_4940,N_4762,N_4781);
xnor U4941 (N_4941,N_4868,N_4805);
nor U4942 (N_4942,N_4778,N_4846);
xor U4943 (N_4943,N_4791,N_4873);
and U4944 (N_4944,N_4772,N_4870);
xnor U4945 (N_4945,N_4845,N_4775);
nand U4946 (N_4946,N_4769,N_4872);
or U4947 (N_4947,N_4861,N_4751);
xor U4948 (N_4948,N_4866,N_4783);
xnor U4949 (N_4949,N_4784,N_4768);
nand U4950 (N_4950,N_4785,N_4797);
nor U4951 (N_4951,N_4794,N_4854);
nor U4952 (N_4952,N_4770,N_4774);
or U4953 (N_4953,N_4771,N_4866);
and U4954 (N_4954,N_4824,N_4776);
and U4955 (N_4955,N_4859,N_4873);
xor U4956 (N_4956,N_4850,N_4783);
nand U4957 (N_4957,N_4838,N_4784);
or U4958 (N_4958,N_4873,N_4750);
and U4959 (N_4959,N_4858,N_4841);
nand U4960 (N_4960,N_4803,N_4793);
or U4961 (N_4961,N_4842,N_4804);
nand U4962 (N_4962,N_4767,N_4836);
xnor U4963 (N_4963,N_4826,N_4859);
nand U4964 (N_4964,N_4792,N_4865);
and U4965 (N_4965,N_4774,N_4794);
or U4966 (N_4966,N_4769,N_4819);
nand U4967 (N_4967,N_4874,N_4811);
nand U4968 (N_4968,N_4858,N_4842);
nand U4969 (N_4969,N_4795,N_4857);
and U4970 (N_4970,N_4836,N_4839);
nor U4971 (N_4971,N_4769,N_4796);
nor U4972 (N_4972,N_4757,N_4821);
and U4973 (N_4973,N_4820,N_4864);
nor U4974 (N_4974,N_4839,N_4835);
and U4975 (N_4975,N_4861,N_4776);
or U4976 (N_4976,N_4763,N_4795);
nand U4977 (N_4977,N_4755,N_4792);
and U4978 (N_4978,N_4752,N_4750);
and U4979 (N_4979,N_4768,N_4781);
xor U4980 (N_4980,N_4792,N_4805);
or U4981 (N_4981,N_4818,N_4843);
and U4982 (N_4982,N_4852,N_4870);
xor U4983 (N_4983,N_4818,N_4851);
nor U4984 (N_4984,N_4817,N_4770);
or U4985 (N_4985,N_4755,N_4819);
or U4986 (N_4986,N_4804,N_4809);
or U4987 (N_4987,N_4867,N_4815);
nand U4988 (N_4988,N_4762,N_4871);
xnor U4989 (N_4989,N_4774,N_4782);
nand U4990 (N_4990,N_4807,N_4866);
nand U4991 (N_4991,N_4796,N_4782);
and U4992 (N_4992,N_4766,N_4827);
nor U4993 (N_4993,N_4801,N_4757);
and U4994 (N_4994,N_4838,N_4766);
nor U4995 (N_4995,N_4870,N_4781);
xnor U4996 (N_4996,N_4855,N_4827);
xor U4997 (N_4997,N_4754,N_4796);
xnor U4998 (N_4998,N_4778,N_4766);
or U4999 (N_4999,N_4864,N_4785);
and U5000 (N_5000,N_4899,N_4931);
nand U5001 (N_5001,N_4960,N_4901);
nor U5002 (N_5002,N_4920,N_4894);
or U5003 (N_5003,N_4979,N_4896);
and U5004 (N_5004,N_4980,N_4902);
xnor U5005 (N_5005,N_4996,N_4878);
or U5006 (N_5006,N_4954,N_4966);
xnor U5007 (N_5007,N_4970,N_4905);
and U5008 (N_5008,N_4881,N_4950);
nor U5009 (N_5009,N_4959,N_4976);
nand U5010 (N_5010,N_4986,N_4952);
and U5011 (N_5011,N_4913,N_4941);
xor U5012 (N_5012,N_4898,N_4947);
and U5013 (N_5013,N_4967,N_4989);
nand U5014 (N_5014,N_4912,N_4922);
nor U5015 (N_5015,N_4883,N_4915);
nand U5016 (N_5016,N_4946,N_4963);
and U5017 (N_5017,N_4914,N_4998);
and U5018 (N_5018,N_4984,N_4876);
or U5019 (N_5019,N_4927,N_4943);
nor U5020 (N_5020,N_4990,N_4992);
or U5021 (N_5021,N_4937,N_4956);
or U5022 (N_5022,N_4875,N_4958);
and U5023 (N_5023,N_4907,N_4925);
xor U5024 (N_5024,N_4945,N_4936);
or U5025 (N_5025,N_4991,N_4917);
or U5026 (N_5026,N_4933,N_4918);
and U5027 (N_5027,N_4891,N_4971);
and U5028 (N_5028,N_4968,N_4957);
nand U5029 (N_5029,N_4887,N_4888);
or U5030 (N_5030,N_4951,N_4892);
xor U5031 (N_5031,N_4978,N_4903);
nor U5032 (N_5032,N_4999,N_4889);
or U5033 (N_5033,N_4964,N_4940);
or U5034 (N_5034,N_4911,N_4879);
xor U5035 (N_5035,N_4928,N_4890);
xnor U5036 (N_5036,N_4934,N_4877);
xnor U5037 (N_5037,N_4955,N_4897);
and U5038 (N_5038,N_4932,N_4944);
and U5039 (N_5039,N_4923,N_4929);
or U5040 (N_5040,N_4884,N_4880);
xor U5041 (N_5041,N_4942,N_4994);
nor U5042 (N_5042,N_4965,N_4882);
nor U5043 (N_5043,N_4906,N_4919);
and U5044 (N_5044,N_4900,N_4974);
nor U5045 (N_5045,N_4969,N_4953);
or U5046 (N_5046,N_4995,N_4886);
nor U5047 (N_5047,N_4948,N_4895);
and U5048 (N_5048,N_4885,N_4993);
or U5049 (N_5049,N_4972,N_4988);
xnor U5050 (N_5050,N_4975,N_4997);
xor U5051 (N_5051,N_4904,N_4987);
or U5052 (N_5052,N_4926,N_4921);
xnor U5053 (N_5053,N_4893,N_4962);
nor U5054 (N_5054,N_4939,N_4909);
or U5055 (N_5055,N_4949,N_4924);
nor U5056 (N_5056,N_4985,N_4973);
nand U5057 (N_5057,N_4916,N_4935);
and U5058 (N_5058,N_4930,N_4982);
or U5059 (N_5059,N_4938,N_4981);
nor U5060 (N_5060,N_4983,N_4977);
xnor U5061 (N_5061,N_4961,N_4910);
nor U5062 (N_5062,N_4908,N_4996);
nand U5063 (N_5063,N_4924,N_4976);
nand U5064 (N_5064,N_4881,N_4913);
nand U5065 (N_5065,N_4940,N_4978);
nor U5066 (N_5066,N_4941,N_4926);
and U5067 (N_5067,N_4891,N_4991);
xnor U5068 (N_5068,N_4993,N_4937);
nand U5069 (N_5069,N_4969,N_4988);
or U5070 (N_5070,N_4964,N_4877);
and U5071 (N_5071,N_4952,N_4923);
nand U5072 (N_5072,N_4879,N_4983);
nor U5073 (N_5073,N_4974,N_4993);
or U5074 (N_5074,N_4977,N_4920);
nor U5075 (N_5075,N_4947,N_4995);
and U5076 (N_5076,N_4882,N_4899);
xor U5077 (N_5077,N_4955,N_4993);
and U5078 (N_5078,N_4961,N_4882);
nand U5079 (N_5079,N_4882,N_4947);
or U5080 (N_5080,N_4904,N_4898);
nor U5081 (N_5081,N_4979,N_4911);
and U5082 (N_5082,N_4970,N_4979);
xor U5083 (N_5083,N_4983,N_4883);
or U5084 (N_5084,N_4886,N_4999);
or U5085 (N_5085,N_4893,N_4974);
xnor U5086 (N_5086,N_4968,N_4951);
nand U5087 (N_5087,N_4879,N_4944);
xor U5088 (N_5088,N_4893,N_4990);
nand U5089 (N_5089,N_4957,N_4906);
or U5090 (N_5090,N_4935,N_4875);
and U5091 (N_5091,N_4942,N_4948);
nand U5092 (N_5092,N_4878,N_4899);
nor U5093 (N_5093,N_4997,N_4977);
or U5094 (N_5094,N_4907,N_4979);
or U5095 (N_5095,N_4881,N_4907);
xor U5096 (N_5096,N_4980,N_4998);
and U5097 (N_5097,N_4908,N_4965);
xor U5098 (N_5098,N_4981,N_4892);
or U5099 (N_5099,N_4879,N_4880);
and U5100 (N_5100,N_4981,N_4974);
or U5101 (N_5101,N_4944,N_4972);
nor U5102 (N_5102,N_4935,N_4950);
and U5103 (N_5103,N_4911,N_4910);
xor U5104 (N_5104,N_4996,N_4879);
and U5105 (N_5105,N_4943,N_4935);
nand U5106 (N_5106,N_4934,N_4924);
or U5107 (N_5107,N_4929,N_4957);
xnor U5108 (N_5108,N_4907,N_4883);
and U5109 (N_5109,N_4875,N_4936);
or U5110 (N_5110,N_4992,N_4969);
and U5111 (N_5111,N_4970,N_4896);
xnor U5112 (N_5112,N_4875,N_4954);
nand U5113 (N_5113,N_4978,N_4987);
or U5114 (N_5114,N_4977,N_4948);
or U5115 (N_5115,N_4952,N_4920);
xnor U5116 (N_5116,N_4964,N_4901);
and U5117 (N_5117,N_4943,N_4995);
nor U5118 (N_5118,N_4913,N_4876);
xnor U5119 (N_5119,N_4925,N_4915);
nand U5120 (N_5120,N_4931,N_4903);
or U5121 (N_5121,N_4901,N_4985);
nand U5122 (N_5122,N_4988,N_4881);
nand U5123 (N_5123,N_4953,N_4919);
xor U5124 (N_5124,N_4880,N_4922);
nand U5125 (N_5125,N_5060,N_5075);
and U5126 (N_5126,N_5055,N_5005);
nand U5127 (N_5127,N_5115,N_5116);
and U5128 (N_5128,N_5088,N_5020);
xnor U5129 (N_5129,N_5080,N_5110);
xor U5130 (N_5130,N_5014,N_5033);
and U5131 (N_5131,N_5121,N_5002);
or U5132 (N_5132,N_5095,N_5008);
nand U5133 (N_5133,N_5022,N_5105);
xnor U5134 (N_5134,N_5083,N_5037);
and U5135 (N_5135,N_5059,N_5078);
nor U5136 (N_5136,N_5036,N_5065);
or U5137 (N_5137,N_5032,N_5018);
and U5138 (N_5138,N_5040,N_5103);
nor U5139 (N_5139,N_5118,N_5007);
xnor U5140 (N_5140,N_5091,N_5077);
or U5141 (N_5141,N_5124,N_5101);
nand U5142 (N_5142,N_5086,N_5109);
nor U5143 (N_5143,N_5062,N_5084);
nand U5144 (N_5144,N_5004,N_5122);
xnor U5145 (N_5145,N_5111,N_5120);
nor U5146 (N_5146,N_5013,N_5073);
or U5147 (N_5147,N_5042,N_5079);
nand U5148 (N_5148,N_5098,N_5010);
nand U5149 (N_5149,N_5049,N_5023);
nor U5150 (N_5150,N_5099,N_5053);
xor U5151 (N_5151,N_5009,N_5061);
xor U5152 (N_5152,N_5089,N_5017);
and U5153 (N_5153,N_5001,N_5071);
nor U5154 (N_5154,N_5016,N_5067);
nor U5155 (N_5155,N_5038,N_5076);
xnor U5156 (N_5156,N_5051,N_5069);
and U5157 (N_5157,N_5056,N_5090);
xnor U5158 (N_5158,N_5000,N_5123);
or U5159 (N_5159,N_5112,N_5034);
nand U5160 (N_5160,N_5019,N_5011);
nand U5161 (N_5161,N_5015,N_5104);
or U5162 (N_5162,N_5070,N_5094);
and U5163 (N_5163,N_5052,N_5100);
and U5164 (N_5164,N_5027,N_5041);
xor U5165 (N_5165,N_5046,N_5107);
nand U5166 (N_5166,N_5097,N_5096);
or U5167 (N_5167,N_5093,N_5047);
xnor U5168 (N_5168,N_5048,N_5025);
and U5169 (N_5169,N_5058,N_5039);
xnor U5170 (N_5170,N_5087,N_5074);
and U5171 (N_5171,N_5054,N_5072);
nor U5172 (N_5172,N_5063,N_5031);
nor U5173 (N_5173,N_5085,N_5106);
and U5174 (N_5174,N_5108,N_5117);
and U5175 (N_5175,N_5030,N_5021);
xor U5176 (N_5176,N_5012,N_5064);
and U5177 (N_5177,N_5066,N_5044);
nor U5178 (N_5178,N_5050,N_5024);
or U5179 (N_5179,N_5006,N_5102);
or U5180 (N_5180,N_5119,N_5057);
xor U5181 (N_5181,N_5092,N_5114);
and U5182 (N_5182,N_5045,N_5043);
nor U5183 (N_5183,N_5029,N_5028);
xnor U5184 (N_5184,N_5026,N_5035);
nor U5185 (N_5185,N_5082,N_5003);
xor U5186 (N_5186,N_5113,N_5068);
xor U5187 (N_5187,N_5081,N_5047);
or U5188 (N_5188,N_5051,N_5006);
nand U5189 (N_5189,N_5006,N_5101);
and U5190 (N_5190,N_5042,N_5017);
and U5191 (N_5191,N_5074,N_5001);
nand U5192 (N_5192,N_5028,N_5078);
or U5193 (N_5193,N_5020,N_5026);
nor U5194 (N_5194,N_5069,N_5021);
or U5195 (N_5195,N_5003,N_5018);
xnor U5196 (N_5196,N_5005,N_5033);
nor U5197 (N_5197,N_5054,N_5047);
nand U5198 (N_5198,N_5072,N_5013);
nor U5199 (N_5199,N_5111,N_5022);
or U5200 (N_5200,N_5035,N_5041);
xnor U5201 (N_5201,N_5061,N_5044);
or U5202 (N_5202,N_5079,N_5005);
xor U5203 (N_5203,N_5039,N_5106);
xor U5204 (N_5204,N_5037,N_5110);
and U5205 (N_5205,N_5069,N_5035);
and U5206 (N_5206,N_5026,N_5094);
or U5207 (N_5207,N_5110,N_5040);
nand U5208 (N_5208,N_5017,N_5003);
xnor U5209 (N_5209,N_5005,N_5006);
and U5210 (N_5210,N_5055,N_5010);
and U5211 (N_5211,N_5017,N_5050);
xor U5212 (N_5212,N_5006,N_5082);
nand U5213 (N_5213,N_5013,N_5088);
and U5214 (N_5214,N_5012,N_5115);
or U5215 (N_5215,N_5035,N_5011);
nand U5216 (N_5216,N_5035,N_5058);
and U5217 (N_5217,N_5045,N_5080);
nand U5218 (N_5218,N_5037,N_5071);
and U5219 (N_5219,N_5118,N_5064);
nand U5220 (N_5220,N_5047,N_5120);
nand U5221 (N_5221,N_5060,N_5098);
xnor U5222 (N_5222,N_5014,N_5006);
xor U5223 (N_5223,N_5063,N_5086);
xor U5224 (N_5224,N_5035,N_5008);
xor U5225 (N_5225,N_5120,N_5008);
or U5226 (N_5226,N_5123,N_5042);
nor U5227 (N_5227,N_5033,N_5048);
nand U5228 (N_5228,N_5023,N_5022);
nand U5229 (N_5229,N_5039,N_5041);
or U5230 (N_5230,N_5069,N_5081);
and U5231 (N_5231,N_5055,N_5071);
nand U5232 (N_5232,N_5038,N_5082);
nand U5233 (N_5233,N_5124,N_5037);
nor U5234 (N_5234,N_5054,N_5062);
nor U5235 (N_5235,N_5040,N_5028);
and U5236 (N_5236,N_5116,N_5067);
nor U5237 (N_5237,N_5067,N_5099);
and U5238 (N_5238,N_5078,N_5068);
and U5239 (N_5239,N_5120,N_5081);
or U5240 (N_5240,N_5012,N_5118);
or U5241 (N_5241,N_5003,N_5089);
xnor U5242 (N_5242,N_5090,N_5017);
xnor U5243 (N_5243,N_5001,N_5107);
nand U5244 (N_5244,N_5062,N_5100);
nand U5245 (N_5245,N_5093,N_5108);
nor U5246 (N_5246,N_5111,N_5024);
xnor U5247 (N_5247,N_5046,N_5006);
and U5248 (N_5248,N_5086,N_5007);
or U5249 (N_5249,N_5003,N_5067);
nor U5250 (N_5250,N_5228,N_5155);
or U5251 (N_5251,N_5182,N_5195);
nor U5252 (N_5252,N_5128,N_5233);
nor U5253 (N_5253,N_5234,N_5216);
and U5254 (N_5254,N_5222,N_5173);
and U5255 (N_5255,N_5165,N_5156);
xnor U5256 (N_5256,N_5180,N_5199);
nor U5257 (N_5257,N_5130,N_5248);
xor U5258 (N_5258,N_5168,N_5148);
xor U5259 (N_5259,N_5153,N_5240);
nor U5260 (N_5260,N_5249,N_5206);
nor U5261 (N_5261,N_5198,N_5246);
or U5262 (N_5262,N_5183,N_5169);
nor U5263 (N_5263,N_5170,N_5139);
or U5264 (N_5264,N_5208,N_5140);
or U5265 (N_5265,N_5188,N_5196);
xnor U5266 (N_5266,N_5181,N_5138);
or U5267 (N_5267,N_5166,N_5224);
xnor U5268 (N_5268,N_5221,N_5151);
or U5269 (N_5269,N_5136,N_5214);
nand U5270 (N_5270,N_5152,N_5193);
nor U5271 (N_5271,N_5232,N_5157);
nand U5272 (N_5272,N_5185,N_5176);
xnor U5273 (N_5273,N_5205,N_5229);
nand U5274 (N_5274,N_5213,N_5134);
or U5275 (N_5275,N_5160,N_5177);
or U5276 (N_5276,N_5244,N_5197);
and U5277 (N_5277,N_5203,N_5141);
or U5278 (N_5278,N_5147,N_5187);
or U5279 (N_5279,N_5161,N_5143);
or U5280 (N_5280,N_5145,N_5158);
xnor U5281 (N_5281,N_5209,N_5192);
nor U5282 (N_5282,N_5142,N_5149);
xor U5283 (N_5283,N_5231,N_5204);
and U5284 (N_5284,N_5211,N_5127);
nor U5285 (N_5285,N_5242,N_5144);
and U5286 (N_5286,N_5178,N_5167);
xor U5287 (N_5287,N_5245,N_5227);
or U5288 (N_5288,N_5241,N_5247);
xor U5289 (N_5289,N_5230,N_5238);
or U5290 (N_5290,N_5217,N_5189);
and U5291 (N_5291,N_5179,N_5154);
nor U5292 (N_5292,N_5132,N_5133);
nor U5293 (N_5293,N_5125,N_5210);
or U5294 (N_5294,N_5239,N_5194);
nand U5295 (N_5295,N_5201,N_5223);
or U5296 (N_5296,N_5184,N_5146);
nor U5297 (N_5297,N_5131,N_5226);
or U5298 (N_5298,N_5186,N_5215);
or U5299 (N_5299,N_5219,N_5174);
nor U5300 (N_5300,N_5135,N_5212);
or U5301 (N_5301,N_5126,N_5164);
and U5302 (N_5302,N_5220,N_5159);
or U5303 (N_5303,N_5202,N_5237);
or U5304 (N_5304,N_5225,N_5190);
nand U5305 (N_5305,N_5162,N_5172);
and U5306 (N_5306,N_5218,N_5137);
and U5307 (N_5307,N_5200,N_5191);
nand U5308 (N_5308,N_5171,N_5236);
or U5309 (N_5309,N_5207,N_5235);
nand U5310 (N_5310,N_5163,N_5243);
and U5311 (N_5311,N_5129,N_5175);
or U5312 (N_5312,N_5150,N_5247);
xnor U5313 (N_5313,N_5129,N_5217);
or U5314 (N_5314,N_5193,N_5147);
nand U5315 (N_5315,N_5196,N_5165);
nand U5316 (N_5316,N_5220,N_5233);
nor U5317 (N_5317,N_5175,N_5241);
or U5318 (N_5318,N_5152,N_5141);
nand U5319 (N_5319,N_5245,N_5200);
or U5320 (N_5320,N_5147,N_5186);
nand U5321 (N_5321,N_5189,N_5138);
xnor U5322 (N_5322,N_5142,N_5198);
xor U5323 (N_5323,N_5183,N_5148);
or U5324 (N_5324,N_5163,N_5216);
nand U5325 (N_5325,N_5142,N_5138);
or U5326 (N_5326,N_5191,N_5173);
nor U5327 (N_5327,N_5198,N_5238);
and U5328 (N_5328,N_5186,N_5146);
nand U5329 (N_5329,N_5242,N_5219);
and U5330 (N_5330,N_5199,N_5158);
nor U5331 (N_5331,N_5140,N_5205);
nand U5332 (N_5332,N_5204,N_5170);
xnor U5333 (N_5333,N_5202,N_5173);
and U5334 (N_5334,N_5191,N_5192);
and U5335 (N_5335,N_5144,N_5137);
nor U5336 (N_5336,N_5235,N_5177);
nand U5337 (N_5337,N_5132,N_5195);
and U5338 (N_5338,N_5140,N_5203);
or U5339 (N_5339,N_5197,N_5178);
or U5340 (N_5340,N_5203,N_5135);
nand U5341 (N_5341,N_5171,N_5142);
or U5342 (N_5342,N_5227,N_5224);
nand U5343 (N_5343,N_5139,N_5245);
or U5344 (N_5344,N_5140,N_5164);
or U5345 (N_5345,N_5167,N_5155);
or U5346 (N_5346,N_5158,N_5202);
nand U5347 (N_5347,N_5151,N_5140);
nor U5348 (N_5348,N_5133,N_5177);
nor U5349 (N_5349,N_5229,N_5202);
nor U5350 (N_5350,N_5175,N_5188);
and U5351 (N_5351,N_5196,N_5219);
and U5352 (N_5352,N_5243,N_5204);
nand U5353 (N_5353,N_5133,N_5217);
nand U5354 (N_5354,N_5215,N_5190);
and U5355 (N_5355,N_5217,N_5231);
xor U5356 (N_5356,N_5248,N_5224);
nor U5357 (N_5357,N_5154,N_5233);
xnor U5358 (N_5358,N_5232,N_5143);
or U5359 (N_5359,N_5249,N_5149);
and U5360 (N_5360,N_5130,N_5211);
xor U5361 (N_5361,N_5128,N_5194);
or U5362 (N_5362,N_5188,N_5159);
nand U5363 (N_5363,N_5209,N_5220);
xor U5364 (N_5364,N_5200,N_5150);
or U5365 (N_5365,N_5159,N_5149);
xor U5366 (N_5366,N_5249,N_5159);
nor U5367 (N_5367,N_5238,N_5131);
xnor U5368 (N_5368,N_5189,N_5222);
xor U5369 (N_5369,N_5248,N_5185);
or U5370 (N_5370,N_5204,N_5226);
or U5371 (N_5371,N_5221,N_5248);
nand U5372 (N_5372,N_5148,N_5241);
and U5373 (N_5373,N_5230,N_5229);
nand U5374 (N_5374,N_5211,N_5210);
and U5375 (N_5375,N_5287,N_5322);
xor U5376 (N_5376,N_5333,N_5367);
xor U5377 (N_5377,N_5268,N_5288);
nand U5378 (N_5378,N_5327,N_5301);
or U5379 (N_5379,N_5340,N_5331);
xor U5380 (N_5380,N_5334,N_5260);
xnor U5381 (N_5381,N_5342,N_5341);
xnor U5382 (N_5382,N_5269,N_5358);
nor U5383 (N_5383,N_5256,N_5262);
or U5384 (N_5384,N_5298,N_5300);
and U5385 (N_5385,N_5309,N_5363);
xnor U5386 (N_5386,N_5326,N_5357);
or U5387 (N_5387,N_5360,N_5279);
and U5388 (N_5388,N_5347,N_5275);
xor U5389 (N_5389,N_5337,N_5373);
nand U5390 (N_5390,N_5281,N_5280);
nor U5391 (N_5391,N_5346,N_5368);
nor U5392 (N_5392,N_5251,N_5305);
and U5393 (N_5393,N_5290,N_5315);
or U5394 (N_5394,N_5265,N_5310);
nand U5395 (N_5395,N_5297,N_5338);
and U5396 (N_5396,N_5344,N_5278);
nand U5397 (N_5397,N_5271,N_5354);
nor U5398 (N_5398,N_5293,N_5339);
and U5399 (N_5399,N_5351,N_5255);
nand U5400 (N_5400,N_5359,N_5283);
xnor U5401 (N_5401,N_5345,N_5261);
xor U5402 (N_5402,N_5336,N_5258);
or U5403 (N_5403,N_5252,N_5324);
nand U5404 (N_5404,N_5319,N_5284);
or U5405 (N_5405,N_5307,N_5289);
nor U5406 (N_5406,N_5316,N_5328);
or U5407 (N_5407,N_5325,N_5371);
or U5408 (N_5408,N_5299,N_5291);
and U5409 (N_5409,N_5374,N_5296);
xnor U5410 (N_5410,N_5329,N_5356);
nor U5411 (N_5411,N_5343,N_5292);
nand U5412 (N_5412,N_5308,N_5274);
nand U5413 (N_5413,N_5264,N_5294);
and U5414 (N_5414,N_5321,N_5366);
nor U5415 (N_5415,N_5352,N_5332);
or U5416 (N_5416,N_5323,N_5361);
and U5417 (N_5417,N_5259,N_5266);
nand U5418 (N_5418,N_5270,N_5302);
nor U5419 (N_5419,N_5276,N_5365);
nor U5420 (N_5420,N_5286,N_5314);
and U5421 (N_5421,N_5306,N_5285);
or U5422 (N_5422,N_5257,N_5263);
or U5423 (N_5423,N_5282,N_5312);
or U5424 (N_5424,N_5273,N_5311);
nor U5425 (N_5425,N_5350,N_5370);
xnor U5426 (N_5426,N_5348,N_5349);
nor U5427 (N_5427,N_5254,N_5313);
xnor U5428 (N_5428,N_5253,N_5304);
xnor U5429 (N_5429,N_5320,N_5355);
nor U5430 (N_5430,N_5250,N_5318);
nand U5431 (N_5431,N_5303,N_5364);
nand U5432 (N_5432,N_5330,N_5353);
nor U5433 (N_5433,N_5317,N_5267);
xor U5434 (N_5434,N_5362,N_5277);
nand U5435 (N_5435,N_5372,N_5272);
and U5436 (N_5436,N_5369,N_5335);
nand U5437 (N_5437,N_5295,N_5270);
xor U5438 (N_5438,N_5325,N_5310);
nor U5439 (N_5439,N_5299,N_5254);
nand U5440 (N_5440,N_5297,N_5359);
xnor U5441 (N_5441,N_5251,N_5292);
and U5442 (N_5442,N_5273,N_5281);
or U5443 (N_5443,N_5267,N_5297);
xor U5444 (N_5444,N_5271,N_5251);
nand U5445 (N_5445,N_5296,N_5336);
nor U5446 (N_5446,N_5333,N_5275);
nor U5447 (N_5447,N_5307,N_5314);
and U5448 (N_5448,N_5361,N_5321);
or U5449 (N_5449,N_5362,N_5298);
nor U5450 (N_5450,N_5287,N_5264);
nor U5451 (N_5451,N_5374,N_5288);
xnor U5452 (N_5452,N_5277,N_5283);
or U5453 (N_5453,N_5272,N_5348);
nand U5454 (N_5454,N_5336,N_5317);
nor U5455 (N_5455,N_5319,N_5365);
nor U5456 (N_5456,N_5331,N_5364);
nand U5457 (N_5457,N_5352,N_5254);
xor U5458 (N_5458,N_5258,N_5294);
nor U5459 (N_5459,N_5332,N_5297);
nand U5460 (N_5460,N_5370,N_5250);
or U5461 (N_5461,N_5288,N_5302);
xor U5462 (N_5462,N_5250,N_5366);
xor U5463 (N_5463,N_5298,N_5330);
xnor U5464 (N_5464,N_5310,N_5318);
and U5465 (N_5465,N_5271,N_5310);
nand U5466 (N_5466,N_5352,N_5356);
nand U5467 (N_5467,N_5276,N_5315);
and U5468 (N_5468,N_5343,N_5263);
nand U5469 (N_5469,N_5338,N_5333);
or U5470 (N_5470,N_5305,N_5291);
nor U5471 (N_5471,N_5315,N_5372);
nand U5472 (N_5472,N_5340,N_5252);
xnor U5473 (N_5473,N_5277,N_5332);
xnor U5474 (N_5474,N_5313,N_5330);
nor U5475 (N_5475,N_5365,N_5346);
and U5476 (N_5476,N_5310,N_5314);
or U5477 (N_5477,N_5344,N_5259);
or U5478 (N_5478,N_5268,N_5341);
nand U5479 (N_5479,N_5297,N_5257);
and U5480 (N_5480,N_5368,N_5313);
nand U5481 (N_5481,N_5304,N_5310);
xor U5482 (N_5482,N_5289,N_5253);
or U5483 (N_5483,N_5310,N_5363);
xor U5484 (N_5484,N_5303,N_5290);
or U5485 (N_5485,N_5260,N_5332);
nor U5486 (N_5486,N_5297,N_5299);
and U5487 (N_5487,N_5253,N_5310);
nand U5488 (N_5488,N_5271,N_5365);
xnor U5489 (N_5489,N_5350,N_5265);
or U5490 (N_5490,N_5272,N_5258);
nor U5491 (N_5491,N_5333,N_5313);
nor U5492 (N_5492,N_5264,N_5299);
nand U5493 (N_5493,N_5316,N_5355);
and U5494 (N_5494,N_5318,N_5319);
or U5495 (N_5495,N_5321,N_5342);
or U5496 (N_5496,N_5363,N_5275);
nand U5497 (N_5497,N_5337,N_5311);
nand U5498 (N_5498,N_5265,N_5258);
nand U5499 (N_5499,N_5305,N_5322);
xnor U5500 (N_5500,N_5448,N_5483);
nor U5501 (N_5501,N_5434,N_5451);
xnor U5502 (N_5502,N_5378,N_5486);
nand U5503 (N_5503,N_5485,N_5436);
nor U5504 (N_5504,N_5493,N_5412);
nor U5505 (N_5505,N_5377,N_5489);
or U5506 (N_5506,N_5411,N_5482);
xnor U5507 (N_5507,N_5398,N_5428);
nor U5508 (N_5508,N_5456,N_5397);
or U5509 (N_5509,N_5442,N_5454);
and U5510 (N_5510,N_5409,N_5443);
nor U5511 (N_5511,N_5497,N_5471);
and U5512 (N_5512,N_5479,N_5460);
nor U5513 (N_5513,N_5403,N_5474);
nand U5514 (N_5514,N_5468,N_5376);
and U5515 (N_5515,N_5408,N_5492);
xor U5516 (N_5516,N_5437,N_5457);
nor U5517 (N_5517,N_5496,N_5452);
nand U5518 (N_5518,N_5381,N_5407);
nor U5519 (N_5519,N_5406,N_5495);
nand U5520 (N_5520,N_5379,N_5430);
or U5521 (N_5521,N_5491,N_5490);
xnor U5522 (N_5522,N_5446,N_5385);
xor U5523 (N_5523,N_5414,N_5417);
nor U5524 (N_5524,N_5404,N_5432);
xor U5525 (N_5525,N_5401,N_5396);
or U5526 (N_5526,N_5413,N_5423);
or U5527 (N_5527,N_5440,N_5494);
nand U5528 (N_5528,N_5499,N_5480);
or U5529 (N_5529,N_5400,N_5402);
and U5530 (N_5530,N_5433,N_5449);
nand U5531 (N_5531,N_5386,N_5463);
nand U5532 (N_5532,N_5420,N_5394);
nand U5533 (N_5533,N_5395,N_5444);
nand U5534 (N_5534,N_5447,N_5393);
nand U5535 (N_5535,N_5383,N_5445);
xnor U5536 (N_5536,N_5458,N_5384);
nand U5537 (N_5537,N_5425,N_5487);
xnor U5538 (N_5538,N_5465,N_5459);
nand U5539 (N_5539,N_5426,N_5450);
or U5540 (N_5540,N_5431,N_5481);
nor U5541 (N_5541,N_5410,N_5476);
nand U5542 (N_5542,N_5415,N_5375);
and U5543 (N_5543,N_5382,N_5498);
xor U5544 (N_5544,N_5461,N_5418);
nand U5545 (N_5545,N_5380,N_5469);
or U5546 (N_5546,N_5484,N_5399);
xnor U5547 (N_5547,N_5464,N_5387);
or U5548 (N_5548,N_5391,N_5470);
xor U5549 (N_5549,N_5419,N_5405);
or U5550 (N_5550,N_5472,N_5488);
xnor U5551 (N_5551,N_5389,N_5473);
and U5552 (N_5552,N_5462,N_5427);
and U5553 (N_5553,N_5455,N_5475);
nand U5554 (N_5554,N_5392,N_5438);
and U5555 (N_5555,N_5416,N_5439);
xnor U5556 (N_5556,N_5453,N_5441);
nor U5557 (N_5557,N_5429,N_5421);
nor U5558 (N_5558,N_5435,N_5424);
nor U5559 (N_5559,N_5466,N_5477);
xnor U5560 (N_5560,N_5422,N_5388);
nor U5561 (N_5561,N_5478,N_5390);
or U5562 (N_5562,N_5467,N_5434);
nor U5563 (N_5563,N_5384,N_5424);
or U5564 (N_5564,N_5384,N_5445);
nor U5565 (N_5565,N_5419,N_5453);
or U5566 (N_5566,N_5416,N_5393);
and U5567 (N_5567,N_5422,N_5410);
nor U5568 (N_5568,N_5401,N_5421);
xnor U5569 (N_5569,N_5430,N_5378);
xnor U5570 (N_5570,N_5496,N_5468);
xnor U5571 (N_5571,N_5411,N_5404);
xnor U5572 (N_5572,N_5433,N_5388);
or U5573 (N_5573,N_5476,N_5419);
or U5574 (N_5574,N_5467,N_5478);
and U5575 (N_5575,N_5475,N_5405);
xnor U5576 (N_5576,N_5445,N_5429);
and U5577 (N_5577,N_5485,N_5404);
or U5578 (N_5578,N_5404,N_5486);
or U5579 (N_5579,N_5434,N_5458);
or U5580 (N_5580,N_5415,N_5476);
or U5581 (N_5581,N_5404,N_5494);
nor U5582 (N_5582,N_5440,N_5412);
nor U5583 (N_5583,N_5481,N_5425);
nand U5584 (N_5584,N_5413,N_5452);
xor U5585 (N_5585,N_5382,N_5413);
nand U5586 (N_5586,N_5432,N_5431);
nand U5587 (N_5587,N_5491,N_5377);
and U5588 (N_5588,N_5452,N_5376);
and U5589 (N_5589,N_5486,N_5414);
nor U5590 (N_5590,N_5435,N_5471);
and U5591 (N_5591,N_5494,N_5422);
nand U5592 (N_5592,N_5423,N_5398);
xnor U5593 (N_5593,N_5398,N_5463);
nor U5594 (N_5594,N_5408,N_5394);
nor U5595 (N_5595,N_5461,N_5379);
nor U5596 (N_5596,N_5399,N_5378);
and U5597 (N_5597,N_5491,N_5470);
and U5598 (N_5598,N_5476,N_5466);
and U5599 (N_5599,N_5376,N_5485);
or U5600 (N_5600,N_5446,N_5390);
or U5601 (N_5601,N_5426,N_5407);
and U5602 (N_5602,N_5423,N_5444);
or U5603 (N_5603,N_5495,N_5487);
or U5604 (N_5604,N_5450,N_5493);
xnor U5605 (N_5605,N_5480,N_5400);
xor U5606 (N_5606,N_5406,N_5417);
or U5607 (N_5607,N_5449,N_5480);
and U5608 (N_5608,N_5488,N_5455);
nor U5609 (N_5609,N_5483,N_5388);
nand U5610 (N_5610,N_5376,N_5455);
nand U5611 (N_5611,N_5399,N_5449);
or U5612 (N_5612,N_5402,N_5385);
nand U5613 (N_5613,N_5463,N_5456);
xnor U5614 (N_5614,N_5462,N_5477);
or U5615 (N_5615,N_5419,N_5463);
and U5616 (N_5616,N_5474,N_5483);
or U5617 (N_5617,N_5403,N_5483);
nor U5618 (N_5618,N_5414,N_5468);
or U5619 (N_5619,N_5397,N_5473);
or U5620 (N_5620,N_5439,N_5426);
nor U5621 (N_5621,N_5378,N_5423);
or U5622 (N_5622,N_5441,N_5420);
and U5623 (N_5623,N_5378,N_5478);
nor U5624 (N_5624,N_5412,N_5490);
or U5625 (N_5625,N_5552,N_5619);
nand U5626 (N_5626,N_5525,N_5567);
and U5627 (N_5627,N_5548,N_5527);
xnor U5628 (N_5628,N_5600,N_5609);
xnor U5629 (N_5629,N_5512,N_5588);
xor U5630 (N_5630,N_5515,N_5544);
and U5631 (N_5631,N_5604,N_5558);
xor U5632 (N_5632,N_5549,N_5614);
nand U5633 (N_5633,N_5577,N_5621);
nor U5634 (N_5634,N_5586,N_5618);
and U5635 (N_5635,N_5505,N_5538);
xnor U5636 (N_5636,N_5547,N_5556);
nand U5637 (N_5637,N_5534,N_5601);
nand U5638 (N_5638,N_5579,N_5503);
or U5639 (N_5639,N_5540,N_5570);
or U5640 (N_5640,N_5599,N_5511);
and U5641 (N_5641,N_5546,N_5605);
nand U5642 (N_5642,N_5612,N_5530);
nand U5643 (N_5643,N_5518,N_5531);
or U5644 (N_5644,N_5542,N_5550);
nor U5645 (N_5645,N_5541,N_5574);
nand U5646 (N_5646,N_5539,N_5524);
xnor U5647 (N_5647,N_5572,N_5555);
xor U5648 (N_5648,N_5522,N_5616);
and U5649 (N_5649,N_5598,N_5576);
nand U5650 (N_5650,N_5578,N_5533);
xnor U5651 (N_5651,N_5543,N_5615);
nand U5652 (N_5652,N_5528,N_5562);
nor U5653 (N_5653,N_5551,N_5620);
xnor U5654 (N_5654,N_5559,N_5573);
xor U5655 (N_5655,N_5523,N_5536);
nor U5656 (N_5656,N_5535,N_5501);
nor U5657 (N_5657,N_5596,N_5591);
and U5658 (N_5658,N_5594,N_5580);
nand U5659 (N_5659,N_5593,N_5521);
nand U5660 (N_5660,N_5565,N_5571);
and U5661 (N_5661,N_5500,N_5623);
nand U5662 (N_5662,N_5545,N_5510);
or U5663 (N_5663,N_5583,N_5582);
nand U5664 (N_5664,N_5557,N_5608);
and U5665 (N_5665,N_5507,N_5508);
nand U5666 (N_5666,N_5590,N_5502);
and U5667 (N_5667,N_5592,N_5568);
and U5668 (N_5668,N_5564,N_5506);
or U5669 (N_5669,N_5585,N_5606);
and U5670 (N_5670,N_5509,N_5617);
xor U5671 (N_5671,N_5602,N_5560);
or U5672 (N_5672,N_5613,N_5519);
or U5673 (N_5673,N_5566,N_5569);
nand U5674 (N_5674,N_5589,N_5610);
nor U5675 (N_5675,N_5513,N_5520);
nor U5676 (N_5676,N_5561,N_5554);
or U5677 (N_5677,N_5514,N_5526);
nand U5678 (N_5678,N_5563,N_5532);
nand U5679 (N_5679,N_5575,N_5553);
or U5680 (N_5680,N_5597,N_5537);
nand U5681 (N_5681,N_5603,N_5584);
nand U5682 (N_5682,N_5622,N_5517);
nor U5683 (N_5683,N_5581,N_5611);
and U5684 (N_5684,N_5595,N_5587);
and U5685 (N_5685,N_5516,N_5624);
xnor U5686 (N_5686,N_5504,N_5607);
nor U5687 (N_5687,N_5529,N_5558);
nor U5688 (N_5688,N_5578,N_5582);
and U5689 (N_5689,N_5518,N_5605);
and U5690 (N_5690,N_5612,N_5517);
nand U5691 (N_5691,N_5544,N_5539);
or U5692 (N_5692,N_5588,N_5502);
nand U5693 (N_5693,N_5576,N_5568);
nor U5694 (N_5694,N_5554,N_5556);
nor U5695 (N_5695,N_5557,N_5593);
nand U5696 (N_5696,N_5572,N_5505);
or U5697 (N_5697,N_5614,N_5605);
nand U5698 (N_5698,N_5524,N_5620);
xor U5699 (N_5699,N_5511,N_5611);
nand U5700 (N_5700,N_5543,N_5533);
nand U5701 (N_5701,N_5592,N_5598);
nor U5702 (N_5702,N_5518,N_5556);
or U5703 (N_5703,N_5531,N_5594);
nand U5704 (N_5704,N_5573,N_5579);
nand U5705 (N_5705,N_5611,N_5536);
or U5706 (N_5706,N_5541,N_5526);
or U5707 (N_5707,N_5624,N_5542);
and U5708 (N_5708,N_5613,N_5570);
and U5709 (N_5709,N_5509,N_5586);
nor U5710 (N_5710,N_5525,N_5604);
nor U5711 (N_5711,N_5596,N_5535);
and U5712 (N_5712,N_5502,N_5570);
nand U5713 (N_5713,N_5587,N_5532);
nor U5714 (N_5714,N_5557,N_5530);
nand U5715 (N_5715,N_5516,N_5574);
nor U5716 (N_5716,N_5597,N_5574);
or U5717 (N_5717,N_5585,N_5602);
nor U5718 (N_5718,N_5590,N_5555);
and U5719 (N_5719,N_5582,N_5575);
or U5720 (N_5720,N_5613,N_5562);
nand U5721 (N_5721,N_5543,N_5536);
nor U5722 (N_5722,N_5503,N_5559);
and U5723 (N_5723,N_5589,N_5580);
xnor U5724 (N_5724,N_5584,N_5573);
nor U5725 (N_5725,N_5570,N_5537);
or U5726 (N_5726,N_5565,N_5585);
nand U5727 (N_5727,N_5522,N_5591);
or U5728 (N_5728,N_5502,N_5508);
nand U5729 (N_5729,N_5600,N_5624);
xnor U5730 (N_5730,N_5508,N_5559);
xnor U5731 (N_5731,N_5531,N_5563);
and U5732 (N_5732,N_5624,N_5540);
and U5733 (N_5733,N_5598,N_5568);
xor U5734 (N_5734,N_5505,N_5579);
and U5735 (N_5735,N_5516,N_5592);
and U5736 (N_5736,N_5592,N_5581);
and U5737 (N_5737,N_5615,N_5575);
or U5738 (N_5738,N_5570,N_5529);
nor U5739 (N_5739,N_5542,N_5537);
nand U5740 (N_5740,N_5556,N_5576);
nor U5741 (N_5741,N_5620,N_5582);
nand U5742 (N_5742,N_5550,N_5526);
or U5743 (N_5743,N_5548,N_5525);
xor U5744 (N_5744,N_5542,N_5520);
xor U5745 (N_5745,N_5591,N_5519);
nor U5746 (N_5746,N_5587,N_5580);
or U5747 (N_5747,N_5544,N_5540);
nand U5748 (N_5748,N_5506,N_5590);
or U5749 (N_5749,N_5590,N_5509);
xor U5750 (N_5750,N_5742,N_5683);
or U5751 (N_5751,N_5677,N_5644);
or U5752 (N_5752,N_5670,N_5626);
nand U5753 (N_5753,N_5687,N_5691);
or U5754 (N_5754,N_5725,N_5637);
xnor U5755 (N_5755,N_5635,N_5633);
nand U5756 (N_5756,N_5726,N_5661);
xnor U5757 (N_5757,N_5748,N_5650);
and U5758 (N_5758,N_5735,N_5666);
and U5759 (N_5759,N_5668,N_5709);
or U5760 (N_5760,N_5696,N_5693);
xnor U5761 (N_5761,N_5636,N_5727);
nand U5762 (N_5762,N_5656,N_5699);
nor U5763 (N_5763,N_5627,N_5667);
nand U5764 (N_5764,N_5684,N_5679);
and U5765 (N_5765,N_5680,N_5625);
xnor U5766 (N_5766,N_5739,N_5662);
or U5767 (N_5767,N_5729,N_5640);
or U5768 (N_5768,N_5718,N_5744);
nand U5769 (N_5769,N_5749,N_5686);
nand U5770 (N_5770,N_5653,N_5655);
xor U5771 (N_5771,N_5663,N_5708);
and U5772 (N_5772,N_5738,N_5701);
nand U5773 (N_5773,N_5690,N_5716);
and U5774 (N_5774,N_5659,N_5643);
or U5775 (N_5775,N_5737,N_5664);
nor U5776 (N_5776,N_5741,N_5675);
nor U5777 (N_5777,N_5734,N_5676);
and U5778 (N_5778,N_5747,N_5673);
or U5779 (N_5779,N_5732,N_5736);
nand U5780 (N_5780,N_5722,N_5712);
nor U5781 (N_5781,N_5730,N_5665);
nand U5782 (N_5782,N_5720,N_5698);
xnor U5783 (N_5783,N_5704,N_5697);
xnor U5784 (N_5784,N_5630,N_5634);
and U5785 (N_5785,N_5731,N_5658);
nand U5786 (N_5786,N_5703,N_5628);
and U5787 (N_5787,N_5681,N_5695);
and U5788 (N_5788,N_5692,N_5723);
nor U5789 (N_5789,N_5669,N_5639);
nand U5790 (N_5790,N_5631,N_5678);
nand U5791 (N_5791,N_5728,N_5710);
nand U5792 (N_5792,N_5724,N_5671);
nor U5793 (N_5793,N_5700,N_5646);
nand U5794 (N_5794,N_5652,N_5649);
xnor U5795 (N_5795,N_5711,N_5689);
and U5796 (N_5796,N_5706,N_5688);
xor U5797 (N_5797,N_5642,N_5702);
nor U5798 (N_5798,N_5645,N_5715);
nor U5799 (N_5799,N_5674,N_5629);
nand U5800 (N_5800,N_5719,N_5672);
nand U5801 (N_5801,N_5647,N_5713);
nand U5802 (N_5802,N_5694,N_5746);
and U5803 (N_5803,N_5654,N_5657);
nor U5804 (N_5804,N_5648,N_5660);
nand U5805 (N_5805,N_5641,N_5707);
nor U5806 (N_5806,N_5733,N_5721);
or U5807 (N_5807,N_5740,N_5705);
and U5808 (N_5808,N_5743,N_5745);
or U5809 (N_5809,N_5685,N_5717);
and U5810 (N_5810,N_5682,N_5651);
nand U5811 (N_5811,N_5714,N_5632);
nand U5812 (N_5812,N_5638,N_5740);
xnor U5813 (N_5813,N_5721,N_5654);
xor U5814 (N_5814,N_5659,N_5700);
xnor U5815 (N_5815,N_5730,N_5715);
nand U5816 (N_5816,N_5712,N_5665);
or U5817 (N_5817,N_5657,N_5637);
nor U5818 (N_5818,N_5629,N_5662);
and U5819 (N_5819,N_5671,N_5747);
xnor U5820 (N_5820,N_5693,N_5687);
or U5821 (N_5821,N_5731,N_5726);
and U5822 (N_5822,N_5644,N_5634);
and U5823 (N_5823,N_5695,N_5743);
or U5824 (N_5824,N_5653,N_5728);
or U5825 (N_5825,N_5737,N_5713);
and U5826 (N_5826,N_5685,N_5637);
nand U5827 (N_5827,N_5675,N_5705);
nor U5828 (N_5828,N_5633,N_5649);
and U5829 (N_5829,N_5627,N_5647);
nor U5830 (N_5830,N_5706,N_5696);
and U5831 (N_5831,N_5685,N_5669);
xor U5832 (N_5832,N_5726,N_5708);
xor U5833 (N_5833,N_5628,N_5633);
and U5834 (N_5834,N_5716,N_5704);
and U5835 (N_5835,N_5665,N_5699);
or U5836 (N_5836,N_5709,N_5749);
and U5837 (N_5837,N_5702,N_5648);
nor U5838 (N_5838,N_5672,N_5716);
and U5839 (N_5839,N_5634,N_5686);
nand U5840 (N_5840,N_5713,N_5691);
and U5841 (N_5841,N_5663,N_5658);
nand U5842 (N_5842,N_5630,N_5632);
nand U5843 (N_5843,N_5728,N_5625);
nand U5844 (N_5844,N_5661,N_5746);
xnor U5845 (N_5845,N_5633,N_5728);
and U5846 (N_5846,N_5634,N_5717);
xor U5847 (N_5847,N_5680,N_5649);
nor U5848 (N_5848,N_5650,N_5630);
nor U5849 (N_5849,N_5697,N_5653);
and U5850 (N_5850,N_5643,N_5719);
nand U5851 (N_5851,N_5626,N_5735);
and U5852 (N_5852,N_5678,N_5704);
or U5853 (N_5853,N_5703,N_5625);
and U5854 (N_5854,N_5639,N_5698);
or U5855 (N_5855,N_5632,N_5627);
xor U5856 (N_5856,N_5625,N_5734);
xor U5857 (N_5857,N_5746,N_5634);
and U5858 (N_5858,N_5677,N_5629);
xnor U5859 (N_5859,N_5716,N_5738);
and U5860 (N_5860,N_5659,N_5703);
xnor U5861 (N_5861,N_5718,N_5736);
or U5862 (N_5862,N_5731,N_5637);
and U5863 (N_5863,N_5730,N_5680);
nand U5864 (N_5864,N_5718,N_5695);
or U5865 (N_5865,N_5669,N_5677);
xnor U5866 (N_5866,N_5641,N_5628);
nor U5867 (N_5867,N_5740,N_5631);
or U5868 (N_5868,N_5724,N_5638);
or U5869 (N_5869,N_5702,N_5699);
and U5870 (N_5870,N_5679,N_5633);
xnor U5871 (N_5871,N_5639,N_5628);
and U5872 (N_5872,N_5676,N_5670);
nor U5873 (N_5873,N_5628,N_5710);
nor U5874 (N_5874,N_5705,N_5635);
or U5875 (N_5875,N_5819,N_5847);
nor U5876 (N_5876,N_5775,N_5858);
and U5877 (N_5877,N_5864,N_5784);
nand U5878 (N_5878,N_5792,N_5757);
nand U5879 (N_5879,N_5843,N_5852);
or U5880 (N_5880,N_5836,N_5818);
nor U5881 (N_5881,N_5767,N_5754);
and U5882 (N_5882,N_5865,N_5872);
or U5883 (N_5883,N_5874,N_5823);
nand U5884 (N_5884,N_5768,N_5822);
xnor U5885 (N_5885,N_5815,N_5857);
nand U5886 (N_5886,N_5830,N_5856);
nor U5887 (N_5887,N_5835,N_5766);
or U5888 (N_5888,N_5838,N_5829);
nand U5889 (N_5889,N_5787,N_5855);
xor U5890 (N_5890,N_5846,N_5825);
xnor U5891 (N_5891,N_5803,N_5790);
or U5892 (N_5892,N_5854,N_5793);
nand U5893 (N_5893,N_5770,N_5764);
nor U5894 (N_5894,N_5828,N_5805);
and U5895 (N_5895,N_5850,N_5786);
xnor U5896 (N_5896,N_5867,N_5831);
nor U5897 (N_5897,N_5842,N_5849);
nand U5898 (N_5898,N_5779,N_5789);
nor U5899 (N_5899,N_5776,N_5769);
and U5900 (N_5900,N_5871,N_5860);
and U5901 (N_5901,N_5808,N_5848);
xnor U5902 (N_5902,N_5817,N_5774);
xor U5903 (N_5903,N_5834,N_5863);
and U5904 (N_5904,N_5810,N_5800);
or U5905 (N_5905,N_5785,N_5833);
nor U5906 (N_5906,N_5765,N_5782);
and U5907 (N_5907,N_5801,N_5781);
nand U5908 (N_5908,N_5794,N_5809);
nand U5909 (N_5909,N_5869,N_5840);
xor U5910 (N_5910,N_5851,N_5796);
nand U5911 (N_5911,N_5859,N_5813);
nand U5912 (N_5912,N_5821,N_5750);
nand U5913 (N_5913,N_5844,N_5806);
and U5914 (N_5914,N_5826,N_5762);
and U5915 (N_5915,N_5772,N_5845);
and U5916 (N_5916,N_5799,N_5763);
and U5917 (N_5917,N_5771,N_5756);
nand U5918 (N_5918,N_5777,N_5804);
or U5919 (N_5919,N_5751,N_5778);
xor U5920 (N_5920,N_5791,N_5873);
nor U5921 (N_5921,N_5795,N_5802);
nor U5922 (N_5922,N_5797,N_5832);
nand U5923 (N_5923,N_5811,N_5824);
xnor U5924 (N_5924,N_5759,N_5870);
and U5925 (N_5925,N_5773,N_5866);
nor U5926 (N_5926,N_5760,N_5841);
xor U5927 (N_5927,N_5807,N_5853);
and U5928 (N_5928,N_5761,N_5755);
or U5929 (N_5929,N_5827,N_5780);
or U5930 (N_5930,N_5839,N_5783);
or U5931 (N_5931,N_5820,N_5752);
and U5932 (N_5932,N_5753,N_5816);
nand U5933 (N_5933,N_5862,N_5868);
xnor U5934 (N_5934,N_5861,N_5814);
or U5935 (N_5935,N_5812,N_5788);
or U5936 (N_5936,N_5837,N_5798);
nand U5937 (N_5937,N_5758,N_5793);
xor U5938 (N_5938,N_5835,N_5751);
nor U5939 (N_5939,N_5800,N_5849);
xor U5940 (N_5940,N_5781,N_5828);
and U5941 (N_5941,N_5869,N_5758);
and U5942 (N_5942,N_5842,N_5764);
nor U5943 (N_5943,N_5865,N_5820);
nand U5944 (N_5944,N_5841,N_5796);
and U5945 (N_5945,N_5845,N_5848);
nor U5946 (N_5946,N_5855,N_5791);
and U5947 (N_5947,N_5831,N_5755);
or U5948 (N_5948,N_5846,N_5872);
nand U5949 (N_5949,N_5870,N_5825);
and U5950 (N_5950,N_5858,N_5753);
and U5951 (N_5951,N_5835,N_5861);
or U5952 (N_5952,N_5861,N_5856);
nand U5953 (N_5953,N_5778,N_5855);
and U5954 (N_5954,N_5870,N_5843);
xor U5955 (N_5955,N_5829,N_5756);
and U5956 (N_5956,N_5818,N_5854);
nor U5957 (N_5957,N_5811,N_5872);
or U5958 (N_5958,N_5866,N_5838);
or U5959 (N_5959,N_5751,N_5776);
and U5960 (N_5960,N_5766,N_5842);
xor U5961 (N_5961,N_5873,N_5777);
and U5962 (N_5962,N_5757,N_5806);
and U5963 (N_5963,N_5869,N_5827);
nand U5964 (N_5964,N_5779,N_5838);
xor U5965 (N_5965,N_5756,N_5761);
nor U5966 (N_5966,N_5787,N_5847);
xor U5967 (N_5967,N_5787,N_5863);
xnor U5968 (N_5968,N_5768,N_5846);
nand U5969 (N_5969,N_5870,N_5798);
xor U5970 (N_5970,N_5844,N_5805);
nor U5971 (N_5971,N_5800,N_5751);
nor U5972 (N_5972,N_5788,N_5869);
or U5973 (N_5973,N_5856,N_5806);
and U5974 (N_5974,N_5814,N_5867);
or U5975 (N_5975,N_5776,N_5775);
nor U5976 (N_5976,N_5850,N_5801);
xor U5977 (N_5977,N_5808,N_5813);
nor U5978 (N_5978,N_5796,N_5775);
nand U5979 (N_5979,N_5822,N_5779);
nand U5980 (N_5980,N_5864,N_5870);
nor U5981 (N_5981,N_5769,N_5792);
xnor U5982 (N_5982,N_5773,N_5828);
or U5983 (N_5983,N_5758,N_5799);
xnor U5984 (N_5984,N_5867,N_5780);
nor U5985 (N_5985,N_5764,N_5828);
or U5986 (N_5986,N_5784,N_5756);
xor U5987 (N_5987,N_5812,N_5815);
or U5988 (N_5988,N_5785,N_5830);
and U5989 (N_5989,N_5760,N_5787);
or U5990 (N_5990,N_5826,N_5782);
nand U5991 (N_5991,N_5870,N_5750);
or U5992 (N_5992,N_5804,N_5850);
or U5993 (N_5993,N_5756,N_5772);
nor U5994 (N_5994,N_5827,N_5820);
nand U5995 (N_5995,N_5872,N_5792);
nor U5996 (N_5996,N_5815,N_5835);
nor U5997 (N_5997,N_5780,N_5830);
xor U5998 (N_5998,N_5809,N_5838);
nor U5999 (N_5999,N_5843,N_5761);
nor U6000 (N_6000,N_5991,N_5925);
and U6001 (N_6001,N_5960,N_5972);
nand U6002 (N_6002,N_5902,N_5917);
xor U6003 (N_6003,N_5936,N_5898);
nand U6004 (N_6004,N_5956,N_5982);
and U6005 (N_6005,N_5878,N_5896);
nor U6006 (N_6006,N_5926,N_5879);
nor U6007 (N_6007,N_5911,N_5975);
or U6008 (N_6008,N_5907,N_5881);
nor U6009 (N_6009,N_5952,N_5959);
nor U6010 (N_6010,N_5942,N_5887);
or U6011 (N_6011,N_5889,N_5892);
nand U6012 (N_6012,N_5886,N_5893);
nand U6013 (N_6013,N_5987,N_5932);
xor U6014 (N_6014,N_5998,N_5914);
xnor U6015 (N_6015,N_5993,N_5882);
nor U6016 (N_6016,N_5970,N_5920);
xor U6017 (N_6017,N_5910,N_5919);
or U6018 (N_6018,N_5974,N_5915);
and U6019 (N_6019,N_5999,N_5958);
nor U6020 (N_6020,N_5966,N_5943);
or U6021 (N_6021,N_5890,N_5909);
nand U6022 (N_6022,N_5888,N_5969);
xor U6023 (N_6023,N_5980,N_5885);
xnor U6024 (N_6024,N_5884,N_5876);
and U6025 (N_6025,N_5957,N_5880);
nor U6026 (N_6026,N_5953,N_5976);
or U6027 (N_6027,N_5922,N_5954);
and U6028 (N_6028,N_5931,N_5948);
nand U6029 (N_6029,N_5899,N_5941);
and U6030 (N_6030,N_5895,N_5961);
nor U6031 (N_6031,N_5950,N_5937);
nand U6032 (N_6032,N_5985,N_5904);
or U6033 (N_6033,N_5921,N_5923);
or U6034 (N_6034,N_5981,N_5997);
nand U6035 (N_6035,N_5913,N_5990);
nand U6036 (N_6036,N_5897,N_5992);
nand U6037 (N_6037,N_5938,N_5988);
xnor U6038 (N_6038,N_5996,N_5995);
nor U6039 (N_6039,N_5946,N_5951);
and U6040 (N_6040,N_5978,N_5940);
or U6041 (N_6041,N_5930,N_5983);
nor U6042 (N_6042,N_5905,N_5900);
and U6043 (N_6043,N_5947,N_5903);
or U6044 (N_6044,N_5934,N_5984);
xor U6045 (N_6045,N_5964,N_5994);
or U6046 (N_6046,N_5986,N_5955);
and U6047 (N_6047,N_5924,N_5891);
and U6048 (N_6048,N_5949,N_5906);
and U6049 (N_6049,N_5989,N_5918);
xnor U6050 (N_6050,N_5965,N_5967);
nor U6051 (N_6051,N_5883,N_5935);
and U6052 (N_6052,N_5877,N_5927);
and U6053 (N_6053,N_5968,N_5908);
xnor U6054 (N_6054,N_5973,N_5912);
nand U6055 (N_6055,N_5944,N_5933);
or U6056 (N_6056,N_5875,N_5971);
nor U6057 (N_6057,N_5962,N_5939);
xor U6058 (N_6058,N_5977,N_5945);
nand U6059 (N_6059,N_5916,N_5963);
xor U6060 (N_6060,N_5979,N_5928);
xnor U6061 (N_6061,N_5894,N_5901);
nand U6062 (N_6062,N_5929,N_5941);
nor U6063 (N_6063,N_5975,N_5973);
and U6064 (N_6064,N_5994,N_5934);
and U6065 (N_6065,N_5938,N_5955);
nand U6066 (N_6066,N_5917,N_5960);
or U6067 (N_6067,N_5980,N_5983);
nand U6068 (N_6068,N_5977,N_5970);
xor U6069 (N_6069,N_5963,N_5932);
nand U6070 (N_6070,N_5928,N_5977);
nand U6071 (N_6071,N_5920,N_5987);
or U6072 (N_6072,N_5955,N_5927);
nor U6073 (N_6073,N_5914,N_5979);
xor U6074 (N_6074,N_5901,N_5899);
and U6075 (N_6075,N_5887,N_5893);
xor U6076 (N_6076,N_5875,N_5919);
nand U6077 (N_6077,N_5943,N_5911);
xor U6078 (N_6078,N_5923,N_5895);
xor U6079 (N_6079,N_5896,N_5969);
nor U6080 (N_6080,N_5896,N_5886);
nor U6081 (N_6081,N_5896,N_5953);
or U6082 (N_6082,N_5897,N_5993);
nand U6083 (N_6083,N_5941,N_5901);
nand U6084 (N_6084,N_5965,N_5896);
or U6085 (N_6085,N_5993,N_5994);
nand U6086 (N_6086,N_5972,N_5929);
and U6087 (N_6087,N_5906,N_5930);
nor U6088 (N_6088,N_5916,N_5923);
xnor U6089 (N_6089,N_5982,N_5930);
xor U6090 (N_6090,N_5938,N_5880);
xor U6091 (N_6091,N_5905,N_5947);
xnor U6092 (N_6092,N_5902,N_5944);
and U6093 (N_6093,N_5920,N_5896);
nor U6094 (N_6094,N_5944,N_5955);
and U6095 (N_6095,N_5917,N_5876);
and U6096 (N_6096,N_5953,N_5973);
nand U6097 (N_6097,N_5900,N_5917);
or U6098 (N_6098,N_5997,N_5962);
nand U6099 (N_6099,N_5942,N_5926);
nor U6100 (N_6100,N_5934,N_5995);
nor U6101 (N_6101,N_5900,N_5991);
nand U6102 (N_6102,N_5954,N_5918);
or U6103 (N_6103,N_5933,N_5922);
xnor U6104 (N_6104,N_5896,N_5908);
or U6105 (N_6105,N_5997,N_5946);
and U6106 (N_6106,N_5901,N_5996);
or U6107 (N_6107,N_5939,N_5919);
xnor U6108 (N_6108,N_5994,N_5911);
xnor U6109 (N_6109,N_5927,N_5944);
or U6110 (N_6110,N_5956,N_5945);
xnor U6111 (N_6111,N_5915,N_5934);
nor U6112 (N_6112,N_5973,N_5957);
nand U6113 (N_6113,N_5969,N_5882);
or U6114 (N_6114,N_5895,N_5986);
nor U6115 (N_6115,N_5941,N_5957);
xor U6116 (N_6116,N_5927,N_5959);
and U6117 (N_6117,N_5878,N_5993);
and U6118 (N_6118,N_5969,N_5968);
nand U6119 (N_6119,N_5875,N_5959);
and U6120 (N_6120,N_5897,N_5921);
and U6121 (N_6121,N_5977,N_5888);
xor U6122 (N_6122,N_5949,N_5895);
nor U6123 (N_6123,N_5952,N_5953);
nand U6124 (N_6124,N_5897,N_5959);
and U6125 (N_6125,N_6031,N_6042);
nand U6126 (N_6126,N_6040,N_6107);
and U6127 (N_6127,N_6073,N_6076);
nand U6128 (N_6128,N_6078,N_6043);
xor U6129 (N_6129,N_6032,N_6004);
and U6130 (N_6130,N_6116,N_6092);
or U6131 (N_6131,N_6086,N_6112);
nor U6132 (N_6132,N_6101,N_6052);
nand U6133 (N_6133,N_6023,N_6102);
nand U6134 (N_6134,N_6016,N_6124);
nand U6135 (N_6135,N_6100,N_6071);
and U6136 (N_6136,N_6065,N_6110);
or U6137 (N_6137,N_6051,N_6055);
nor U6138 (N_6138,N_6070,N_6027);
and U6139 (N_6139,N_6087,N_6018);
nor U6140 (N_6140,N_6064,N_6111);
nand U6141 (N_6141,N_6013,N_6057);
and U6142 (N_6142,N_6096,N_6011);
nor U6143 (N_6143,N_6010,N_6119);
xor U6144 (N_6144,N_6089,N_6091);
or U6145 (N_6145,N_6060,N_6117);
or U6146 (N_6146,N_6113,N_6108);
nor U6147 (N_6147,N_6099,N_6053);
nand U6148 (N_6148,N_6050,N_6035);
nor U6149 (N_6149,N_6094,N_6095);
and U6150 (N_6150,N_6029,N_6058);
xnor U6151 (N_6151,N_6088,N_6066);
and U6152 (N_6152,N_6025,N_6005);
xor U6153 (N_6153,N_6046,N_6034);
nor U6154 (N_6154,N_6068,N_6072);
xor U6155 (N_6155,N_6009,N_6056);
nor U6156 (N_6156,N_6014,N_6118);
or U6157 (N_6157,N_6038,N_6084);
nor U6158 (N_6158,N_6001,N_6026);
nor U6159 (N_6159,N_6063,N_6039);
nand U6160 (N_6160,N_6002,N_6083);
nand U6161 (N_6161,N_6098,N_6024);
xor U6162 (N_6162,N_6120,N_6085);
nand U6163 (N_6163,N_6082,N_6041);
nand U6164 (N_6164,N_6059,N_6021);
nand U6165 (N_6165,N_6093,N_6017);
xor U6166 (N_6166,N_6007,N_6074);
nor U6167 (N_6167,N_6062,N_6033);
nor U6168 (N_6168,N_6079,N_6036);
xnor U6169 (N_6169,N_6045,N_6122);
and U6170 (N_6170,N_6048,N_6012);
and U6171 (N_6171,N_6109,N_6067);
nand U6172 (N_6172,N_6047,N_6030);
nor U6173 (N_6173,N_6081,N_6003);
and U6174 (N_6174,N_6022,N_6037);
nor U6175 (N_6175,N_6020,N_6105);
and U6176 (N_6176,N_6015,N_6019);
and U6177 (N_6177,N_6090,N_6104);
or U6178 (N_6178,N_6049,N_6121);
nand U6179 (N_6179,N_6054,N_6077);
and U6180 (N_6180,N_6080,N_6123);
and U6181 (N_6181,N_6000,N_6028);
nand U6182 (N_6182,N_6044,N_6106);
xor U6183 (N_6183,N_6006,N_6061);
or U6184 (N_6184,N_6069,N_6008);
and U6185 (N_6185,N_6114,N_6115);
and U6186 (N_6186,N_6097,N_6075);
and U6187 (N_6187,N_6103,N_6079);
nor U6188 (N_6188,N_6108,N_6116);
and U6189 (N_6189,N_6013,N_6097);
nor U6190 (N_6190,N_6061,N_6089);
and U6191 (N_6191,N_6111,N_6103);
or U6192 (N_6192,N_6107,N_6066);
or U6193 (N_6193,N_6124,N_6075);
nand U6194 (N_6194,N_6008,N_6009);
nor U6195 (N_6195,N_6055,N_6001);
nand U6196 (N_6196,N_6042,N_6079);
or U6197 (N_6197,N_6082,N_6102);
or U6198 (N_6198,N_6005,N_6039);
nand U6199 (N_6199,N_6057,N_6109);
nand U6200 (N_6200,N_6077,N_6055);
xor U6201 (N_6201,N_6098,N_6025);
and U6202 (N_6202,N_6092,N_6007);
or U6203 (N_6203,N_6063,N_6008);
and U6204 (N_6204,N_6097,N_6039);
xor U6205 (N_6205,N_6026,N_6071);
nand U6206 (N_6206,N_6037,N_6035);
nand U6207 (N_6207,N_6028,N_6002);
or U6208 (N_6208,N_6006,N_6073);
or U6209 (N_6209,N_6083,N_6097);
nor U6210 (N_6210,N_6051,N_6040);
nor U6211 (N_6211,N_6076,N_6050);
and U6212 (N_6212,N_6101,N_6039);
and U6213 (N_6213,N_6055,N_6120);
and U6214 (N_6214,N_6054,N_6100);
nor U6215 (N_6215,N_6020,N_6047);
nor U6216 (N_6216,N_6093,N_6094);
or U6217 (N_6217,N_6085,N_6047);
nand U6218 (N_6218,N_6095,N_6034);
xnor U6219 (N_6219,N_6021,N_6015);
nor U6220 (N_6220,N_6013,N_6025);
and U6221 (N_6221,N_6074,N_6058);
and U6222 (N_6222,N_6079,N_6034);
xnor U6223 (N_6223,N_6123,N_6029);
or U6224 (N_6224,N_6124,N_6032);
and U6225 (N_6225,N_6119,N_6022);
or U6226 (N_6226,N_6119,N_6105);
or U6227 (N_6227,N_6010,N_6076);
xor U6228 (N_6228,N_6056,N_6076);
nand U6229 (N_6229,N_6056,N_6084);
nand U6230 (N_6230,N_6114,N_6089);
xnor U6231 (N_6231,N_6086,N_6021);
or U6232 (N_6232,N_6031,N_6007);
or U6233 (N_6233,N_6088,N_6038);
nand U6234 (N_6234,N_6061,N_6053);
nor U6235 (N_6235,N_6090,N_6084);
or U6236 (N_6236,N_6114,N_6049);
xnor U6237 (N_6237,N_6097,N_6005);
or U6238 (N_6238,N_6087,N_6055);
nor U6239 (N_6239,N_6089,N_6006);
nor U6240 (N_6240,N_6057,N_6049);
and U6241 (N_6241,N_6097,N_6070);
and U6242 (N_6242,N_6036,N_6040);
nand U6243 (N_6243,N_6063,N_6102);
xor U6244 (N_6244,N_6017,N_6013);
nand U6245 (N_6245,N_6064,N_6124);
xnor U6246 (N_6246,N_6093,N_6018);
xor U6247 (N_6247,N_6061,N_6004);
xnor U6248 (N_6248,N_6103,N_6120);
nand U6249 (N_6249,N_6066,N_6009);
and U6250 (N_6250,N_6193,N_6169);
and U6251 (N_6251,N_6127,N_6149);
or U6252 (N_6252,N_6196,N_6236);
nand U6253 (N_6253,N_6225,N_6217);
nor U6254 (N_6254,N_6126,N_6135);
xor U6255 (N_6255,N_6164,N_6220);
nand U6256 (N_6256,N_6177,N_6239);
xor U6257 (N_6257,N_6235,N_6152);
nand U6258 (N_6258,N_6183,N_6155);
nand U6259 (N_6259,N_6132,N_6175);
and U6260 (N_6260,N_6187,N_6222);
nand U6261 (N_6261,N_6130,N_6182);
nand U6262 (N_6262,N_6189,N_6208);
nand U6263 (N_6263,N_6234,N_6249);
xor U6264 (N_6264,N_6139,N_6246);
or U6265 (N_6265,N_6214,N_6201);
nand U6266 (N_6266,N_6160,N_6204);
or U6267 (N_6267,N_6188,N_6159);
xnor U6268 (N_6268,N_6148,N_6248);
nor U6269 (N_6269,N_6206,N_6154);
xor U6270 (N_6270,N_6185,N_6218);
and U6271 (N_6271,N_6141,N_6145);
and U6272 (N_6272,N_6229,N_6162);
or U6273 (N_6273,N_6125,N_6194);
xor U6274 (N_6274,N_6163,N_6211);
nor U6275 (N_6275,N_6147,N_6212);
nand U6276 (N_6276,N_6176,N_6156);
nor U6277 (N_6277,N_6143,N_6198);
xor U6278 (N_6278,N_6247,N_6144);
nand U6279 (N_6279,N_6137,N_6179);
xnor U6280 (N_6280,N_6166,N_6219);
nor U6281 (N_6281,N_6178,N_6140);
nor U6282 (N_6282,N_6158,N_6231);
or U6283 (N_6283,N_6221,N_6200);
and U6284 (N_6284,N_6184,N_6207);
and U6285 (N_6285,N_6242,N_6171);
and U6286 (N_6286,N_6167,N_6138);
nor U6287 (N_6287,N_6142,N_6216);
xnor U6288 (N_6288,N_6128,N_6245);
and U6289 (N_6289,N_6136,N_6191);
and U6290 (N_6290,N_6228,N_6180);
and U6291 (N_6291,N_6227,N_6134);
nor U6292 (N_6292,N_6243,N_6150);
or U6293 (N_6293,N_6233,N_6153);
nor U6294 (N_6294,N_6195,N_6202);
nand U6295 (N_6295,N_6157,N_6215);
nor U6296 (N_6296,N_6186,N_6146);
nor U6297 (N_6297,N_6237,N_6238);
and U6298 (N_6298,N_6230,N_6192);
nor U6299 (N_6299,N_6161,N_6205);
nand U6300 (N_6300,N_6203,N_6223);
and U6301 (N_6301,N_6133,N_6197);
nand U6302 (N_6302,N_6209,N_6129);
nor U6303 (N_6303,N_6241,N_6168);
xnor U6304 (N_6304,N_6151,N_6226);
or U6305 (N_6305,N_6232,N_6240);
or U6306 (N_6306,N_6244,N_6131);
and U6307 (N_6307,N_6165,N_6173);
nand U6308 (N_6308,N_6224,N_6181);
xnor U6309 (N_6309,N_6199,N_6174);
and U6310 (N_6310,N_6170,N_6172);
or U6311 (N_6311,N_6210,N_6190);
or U6312 (N_6312,N_6213,N_6169);
and U6313 (N_6313,N_6236,N_6220);
nor U6314 (N_6314,N_6222,N_6211);
nand U6315 (N_6315,N_6126,N_6170);
xor U6316 (N_6316,N_6161,N_6154);
and U6317 (N_6317,N_6171,N_6167);
or U6318 (N_6318,N_6205,N_6136);
and U6319 (N_6319,N_6129,N_6160);
and U6320 (N_6320,N_6173,N_6245);
xnor U6321 (N_6321,N_6235,N_6192);
xor U6322 (N_6322,N_6189,N_6166);
nor U6323 (N_6323,N_6129,N_6125);
nor U6324 (N_6324,N_6188,N_6245);
and U6325 (N_6325,N_6189,N_6231);
and U6326 (N_6326,N_6195,N_6214);
nor U6327 (N_6327,N_6229,N_6137);
or U6328 (N_6328,N_6245,N_6176);
or U6329 (N_6329,N_6177,N_6187);
or U6330 (N_6330,N_6219,N_6210);
and U6331 (N_6331,N_6167,N_6193);
or U6332 (N_6332,N_6220,N_6227);
nor U6333 (N_6333,N_6183,N_6147);
or U6334 (N_6334,N_6202,N_6203);
nand U6335 (N_6335,N_6243,N_6216);
xnor U6336 (N_6336,N_6130,N_6249);
or U6337 (N_6337,N_6205,N_6218);
or U6338 (N_6338,N_6242,N_6232);
nand U6339 (N_6339,N_6196,N_6195);
xnor U6340 (N_6340,N_6236,N_6156);
or U6341 (N_6341,N_6206,N_6152);
or U6342 (N_6342,N_6189,N_6215);
nand U6343 (N_6343,N_6219,N_6127);
nor U6344 (N_6344,N_6165,N_6217);
and U6345 (N_6345,N_6202,N_6248);
nor U6346 (N_6346,N_6134,N_6185);
or U6347 (N_6347,N_6144,N_6163);
nand U6348 (N_6348,N_6180,N_6165);
and U6349 (N_6349,N_6196,N_6201);
nand U6350 (N_6350,N_6151,N_6237);
xnor U6351 (N_6351,N_6181,N_6226);
nand U6352 (N_6352,N_6199,N_6243);
nand U6353 (N_6353,N_6248,N_6178);
nor U6354 (N_6354,N_6163,N_6227);
xor U6355 (N_6355,N_6249,N_6200);
nor U6356 (N_6356,N_6178,N_6133);
nand U6357 (N_6357,N_6139,N_6189);
or U6358 (N_6358,N_6132,N_6218);
nand U6359 (N_6359,N_6148,N_6166);
nor U6360 (N_6360,N_6198,N_6197);
and U6361 (N_6361,N_6201,N_6163);
and U6362 (N_6362,N_6160,N_6126);
and U6363 (N_6363,N_6183,N_6151);
xnor U6364 (N_6364,N_6179,N_6155);
nor U6365 (N_6365,N_6179,N_6190);
nand U6366 (N_6366,N_6137,N_6227);
nand U6367 (N_6367,N_6173,N_6186);
xor U6368 (N_6368,N_6143,N_6141);
or U6369 (N_6369,N_6135,N_6136);
nand U6370 (N_6370,N_6180,N_6139);
and U6371 (N_6371,N_6212,N_6238);
or U6372 (N_6372,N_6173,N_6180);
xnor U6373 (N_6373,N_6242,N_6185);
and U6374 (N_6374,N_6198,N_6226);
and U6375 (N_6375,N_6289,N_6320);
or U6376 (N_6376,N_6268,N_6279);
xor U6377 (N_6377,N_6334,N_6315);
xnor U6378 (N_6378,N_6366,N_6271);
xor U6379 (N_6379,N_6347,N_6277);
or U6380 (N_6380,N_6357,N_6344);
or U6381 (N_6381,N_6371,N_6374);
nor U6382 (N_6382,N_6345,N_6287);
or U6383 (N_6383,N_6251,N_6361);
nand U6384 (N_6384,N_6253,N_6254);
and U6385 (N_6385,N_6343,N_6317);
nand U6386 (N_6386,N_6352,N_6358);
nand U6387 (N_6387,N_6321,N_6294);
nor U6388 (N_6388,N_6328,N_6295);
nor U6389 (N_6389,N_6325,N_6274);
and U6390 (N_6390,N_6342,N_6263);
or U6391 (N_6391,N_6331,N_6359);
nor U6392 (N_6392,N_6350,N_6354);
and U6393 (N_6393,N_6337,N_6270);
or U6394 (N_6394,N_6282,N_6362);
xor U6395 (N_6395,N_6252,N_6355);
nand U6396 (N_6396,N_6258,N_6330);
xnor U6397 (N_6397,N_6286,N_6329);
xnor U6398 (N_6398,N_6340,N_6335);
xnor U6399 (N_6399,N_6281,N_6314);
nand U6400 (N_6400,N_6319,N_6250);
xnor U6401 (N_6401,N_6273,N_6280);
and U6402 (N_6402,N_6256,N_6272);
nand U6403 (N_6403,N_6297,N_6356);
nand U6404 (N_6404,N_6299,N_6283);
and U6405 (N_6405,N_6278,N_6364);
nand U6406 (N_6406,N_6363,N_6276);
nor U6407 (N_6407,N_6296,N_6266);
and U6408 (N_6408,N_6262,N_6261);
nor U6409 (N_6409,N_6372,N_6265);
and U6410 (N_6410,N_6255,N_6327);
and U6411 (N_6411,N_6370,N_6288);
nor U6412 (N_6412,N_6311,N_6339);
nand U6413 (N_6413,N_6353,N_6307);
and U6414 (N_6414,N_6341,N_6309);
nand U6415 (N_6415,N_6312,N_6298);
and U6416 (N_6416,N_6323,N_6284);
nor U6417 (N_6417,N_6308,N_6313);
nand U6418 (N_6418,N_6316,N_6338);
xor U6419 (N_6419,N_6301,N_6292);
or U6420 (N_6420,N_6349,N_6285);
nand U6421 (N_6421,N_6259,N_6300);
and U6422 (N_6422,N_6332,N_6260);
nor U6423 (N_6423,N_6346,N_6369);
nand U6424 (N_6424,N_6318,N_6267);
and U6425 (N_6425,N_6310,N_6293);
xor U6426 (N_6426,N_6322,N_6257);
and U6427 (N_6427,N_6368,N_6306);
and U6428 (N_6428,N_6304,N_6326);
xor U6429 (N_6429,N_6351,N_6269);
nor U6430 (N_6430,N_6303,N_6302);
nor U6431 (N_6431,N_6264,N_6365);
nand U6432 (N_6432,N_6290,N_6348);
or U6433 (N_6433,N_6324,N_6275);
xor U6434 (N_6434,N_6336,N_6305);
and U6435 (N_6435,N_6291,N_6333);
and U6436 (N_6436,N_6373,N_6367);
xnor U6437 (N_6437,N_6360,N_6256);
or U6438 (N_6438,N_6294,N_6296);
and U6439 (N_6439,N_6340,N_6350);
and U6440 (N_6440,N_6263,N_6279);
nor U6441 (N_6441,N_6351,N_6258);
or U6442 (N_6442,N_6290,N_6295);
xor U6443 (N_6443,N_6296,N_6272);
nand U6444 (N_6444,N_6295,N_6324);
or U6445 (N_6445,N_6352,N_6344);
nor U6446 (N_6446,N_6368,N_6252);
or U6447 (N_6447,N_6251,N_6267);
xnor U6448 (N_6448,N_6331,N_6323);
xnor U6449 (N_6449,N_6372,N_6323);
or U6450 (N_6450,N_6366,N_6251);
xnor U6451 (N_6451,N_6363,N_6348);
or U6452 (N_6452,N_6282,N_6363);
nor U6453 (N_6453,N_6297,N_6358);
xnor U6454 (N_6454,N_6371,N_6315);
nor U6455 (N_6455,N_6275,N_6265);
and U6456 (N_6456,N_6269,N_6297);
xor U6457 (N_6457,N_6347,N_6348);
xnor U6458 (N_6458,N_6338,N_6372);
or U6459 (N_6459,N_6276,N_6274);
or U6460 (N_6460,N_6302,N_6362);
or U6461 (N_6461,N_6327,N_6281);
nor U6462 (N_6462,N_6276,N_6292);
nand U6463 (N_6463,N_6349,N_6342);
or U6464 (N_6464,N_6348,N_6351);
nor U6465 (N_6465,N_6316,N_6351);
xnor U6466 (N_6466,N_6328,N_6331);
and U6467 (N_6467,N_6317,N_6267);
and U6468 (N_6468,N_6320,N_6301);
and U6469 (N_6469,N_6299,N_6288);
nor U6470 (N_6470,N_6343,N_6252);
nor U6471 (N_6471,N_6308,N_6272);
or U6472 (N_6472,N_6349,N_6295);
or U6473 (N_6473,N_6353,N_6289);
nor U6474 (N_6474,N_6282,N_6267);
xnor U6475 (N_6475,N_6288,N_6260);
and U6476 (N_6476,N_6365,N_6303);
or U6477 (N_6477,N_6340,N_6363);
nor U6478 (N_6478,N_6257,N_6332);
nor U6479 (N_6479,N_6289,N_6341);
xnor U6480 (N_6480,N_6324,N_6342);
nand U6481 (N_6481,N_6363,N_6368);
xor U6482 (N_6482,N_6299,N_6353);
nor U6483 (N_6483,N_6343,N_6324);
nand U6484 (N_6484,N_6261,N_6270);
xnor U6485 (N_6485,N_6294,N_6334);
nand U6486 (N_6486,N_6344,N_6362);
or U6487 (N_6487,N_6317,N_6312);
and U6488 (N_6488,N_6324,N_6255);
nand U6489 (N_6489,N_6287,N_6348);
nand U6490 (N_6490,N_6291,N_6269);
or U6491 (N_6491,N_6264,N_6299);
and U6492 (N_6492,N_6329,N_6299);
xor U6493 (N_6493,N_6291,N_6368);
nor U6494 (N_6494,N_6252,N_6305);
xnor U6495 (N_6495,N_6310,N_6351);
or U6496 (N_6496,N_6310,N_6338);
or U6497 (N_6497,N_6251,N_6306);
or U6498 (N_6498,N_6370,N_6270);
nor U6499 (N_6499,N_6325,N_6250);
xor U6500 (N_6500,N_6475,N_6441);
or U6501 (N_6501,N_6427,N_6429);
nand U6502 (N_6502,N_6468,N_6444);
xor U6503 (N_6503,N_6467,N_6419);
or U6504 (N_6504,N_6489,N_6400);
or U6505 (N_6505,N_6417,N_6454);
and U6506 (N_6506,N_6438,N_6393);
or U6507 (N_6507,N_6381,N_6447);
nand U6508 (N_6508,N_6412,N_6394);
nor U6509 (N_6509,N_6473,N_6395);
nor U6510 (N_6510,N_6422,N_6469);
nand U6511 (N_6511,N_6464,N_6391);
xnor U6512 (N_6512,N_6420,N_6477);
and U6513 (N_6513,N_6380,N_6471);
nor U6514 (N_6514,N_6396,N_6385);
and U6515 (N_6515,N_6411,N_6431);
or U6516 (N_6516,N_6414,N_6426);
or U6517 (N_6517,N_6432,N_6463);
nor U6518 (N_6518,N_6498,N_6401);
nand U6519 (N_6519,N_6440,N_6458);
nor U6520 (N_6520,N_6390,N_6495);
or U6521 (N_6521,N_6497,N_6491);
xor U6522 (N_6522,N_6375,N_6428);
nand U6523 (N_6523,N_6494,N_6416);
nor U6524 (N_6524,N_6499,N_6485);
nand U6525 (N_6525,N_6442,N_6392);
nor U6526 (N_6526,N_6436,N_6418);
or U6527 (N_6527,N_6453,N_6404);
xor U6528 (N_6528,N_6488,N_6397);
and U6529 (N_6529,N_6483,N_6408);
or U6530 (N_6530,N_6478,N_6433);
nand U6531 (N_6531,N_6465,N_6466);
nor U6532 (N_6532,N_6455,N_6482);
and U6533 (N_6533,N_6387,N_6383);
nor U6534 (N_6534,N_6445,N_6384);
and U6535 (N_6535,N_6446,N_6496);
or U6536 (N_6536,N_6484,N_6410);
or U6537 (N_6537,N_6415,N_6448);
xnor U6538 (N_6538,N_6443,N_6382);
nor U6539 (N_6539,N_6492,N_6490);
xor U6540 (N_6540,N_6377,N_6424);
or U6541 (N_6541,N_6462,N_6421);
nand U6542 (N_6542,N_6452,N_6423);
nand U6543 (N_6543,N_6487,N_6451);
nor U6544 (N_6544,N_6435,N_6430);
or U6545 (N_6545,N_6450,N_6434);
and U6546 (N_6546,N_6470,N_6461);
nor U6547 (N_6547,N_6437,N_6481);
and U6548 (N_6548,N_6376,N_6457);
nand U6549 (N_6549,N_6459,N_6409);
xnor U6550 (N_6550,N_6460,N_6449);
nand U6551 (N_6551,N_6405,N_6403);
or U6552 (N_6552,N_6379,N_6398);
nor U6553 (N_6553,N_6456,N_6439);
and U6554 (N_6554,N_6476,N_6402);
xnor U6555 (N_6555,N_6389,N_6425);
and U6556 (N_6556,N_6388,N_6486);
and U6557 (N_6557,N_6378,N_6480);
and U6558 (N_6558,N_6474,N_6386);
and U6559 (N_6559,N_6407,N_6479);
or U6560 (N_6560,N_6472,N_6406);
or U6561 (N_6561,N_6493,N_6413);
xnor U6562 (N_6562,N_6399,N_6454);
nand U6563 (N_6563,N_6409,N_6414);
xnor U6564 (N_6564,N_6384,N_6450);
nor U6565 (N_6565,N_6469,N_6460);
xnor U6566 (N_6566,N_6389,N_6397);
xnor U6567 (N_6567,N_6406,N_6454);
xor U6568 (N_6568,N_6391,N_6399);
or U6569 (N_6569,N_6395,N_6385);
nor U6570 (N_6570,N_6431,N_6406);
and U6571 (N_6571,N_6449,N_6448);
and U6572 (N_6572,N_6434,N_6461);
nor U6573 (N_6573,N_6439,N_6437);
or U6574 (N_6574,N_6409,N_6448);
xnor U6575 (N_6575,N_6385,N_6456);
nand U6576 (N_6576,N_6431,N_6433);
nand U6577 (N_6577,N_6376,N_6431);
and U6578 (N_6578,N_6404,N_6473);
nor U6579 (N_6579,N_6457,N_6400);
nand U6580 (N_6580,N_6436,N_6489);
nand U6581 (N_6581,N_6487,N_6416);
and U6582 (N_6582,N_6447,N_6433);
nand U6583 (N_6583,N_6452,N_6429);
or U6584 (N_6584,N_6470,N_6466);
or U6585 (N_6585,N_6465,N_6381);
xnor U6586 (N_6586,N_6394,N_6459);
or U6587 (N_6587,N_6421,N_6375);
nor U6588 (N_6588,N_6382,N_6411);
or U6589 (N_6589,N_6417,N_6497);
xor U6590 (N_6590,N_6396,N_6479);
nor U6591 (N_6591,N_6378,N_6424);
xnor U6592 (N_6592,N_6413,N_6495);
xor U6593 (N_6593,N_6460,N_6439);
and U6594 (N_6594,N_6495,N_6457);
xnor U6595 (N_6595,N_6437,N_6466);
or U6596 (N_6596,N_6400,N_6381);
or U6597 (N_6597,N_6451,N_6384);
or U6598 (N_6598,N_6434,N_6437);
or U6599 (N_6599,N_6481,N_6411);
or U6600 (N_6600,N_6468,N_6430);
xnor U6601 (N_6601,N_6479,N_6495);
and U6602 (N_6602,N_6402,N_6493);
and U6603 (N_6603,N_6455,N_6490);
nand U6604 (N_6604,N_6462,N_6423);
or U6605 (N_6605,N_6431,N_6386);
nor U6606 (N_6606,N_6413,N_6425);
nor U6607 (N_6607,N_6412,N_6434);
nor U6608 (N_6608,N_6477,N_6422);
nor U6609 (N_6609,N_6406,N_6440);
nor U6610 (N_6610,N_6411,N_6412);
nand U6611 (N_6611,N_6436,N_6475);
or U6612 (N_6612,N_6410,N_6404);
nor U6613 (N_6613,N_6492,N_6448);
and U6614 (N_6614,N_6450,N_6397);
and U6615 (N_6615,N_6458,N_6470);
nor U6616 (N_6616,N_6430,N_6412);
or U6617 (N_6617,N_6450,N_6407);
and U6618 (N_6618,N_6409,N_6412);
or U6619 (N_6619,N_6447,N_6471);
nand U6620 (N_6620,N_6411,N_6497);
xor U6621 (N_6621,N_6378,N_6496);
xnor U6622 (N_6622,N_6408,N_6430);
nand U6623 (N_6623,N_6495,N_6398);
or U6624 (N_6624,N_6499,N_6412);
nand U6625 (N_6625,N_6589,N_6573);
nand U6626 (N_6626,N_6516,N_6617);
nor U6627 (N_6627,N_6609,N_6588);
and U6628 (N_6628,N_6513,N_6613);
and U6629 (N_6629,N_6556,N_6526);
xnor U6630 (N_6630,N_6577,N_6622);
xor U6631 (N_6631,N_6533,N_6549);
nand U6632 (N_6632,N_6523,N_6603);
and U6633 (N_6633,N_6565,N_6608);
nand U6634 (N_6634,N_6501,N_6606);
xnor U6635 (N_6635,N_6527,N_6576);
and U6636 (N_6636,N_6600,N_6515);
or U6637 (N_6637,N_6596,N_6570);
nand U6638 (N_6638,N_6534,N_6503);
and U6639 (N_6639,N_6605,N_6517);
nor U6640 (N_6640,N_6557,N_6543);
or U6641 (N_6641,N_6539,N_6624);
nand U6642 (N_6642,N_6508,N_6590);
nand U6643 (N_6643,N_6510,N_6528);
and U6644 (N_6644,N_6532,N_6550);
nor U6645 (N_6645,N_6555,N_6502);
nand U6646 (N_6646,N_6521,N_6524);
or U6647 (N_6647,N_6615,N_6580);
nor U6648 (N_6648,N_6530,N_6522);
and U6649 (N_6649,N_6561,N_6614);
nor U6650 (N_6650,N_6619,N_6616);
nor U6651 (N_6651,N_6507,N_6604);
and U6652 (N_6652,N_6531,N_6568);
and U6653 (N_6653,N_6574,N_6538);
nor U6654 (N_6654,N_6567,N_6602);
xnor U6655 (N_6655,N_6601,N_6563);
nor U6656 (N_6656,N_6562,N_6506);
xor U6657 (N_6657,N_6500,N_6511);
xnor U6658 (N_6658,N_6548,N_6542);
and U6659 (N_6659,N_6578,N_6618);
and U6660 (N_6660,N_6553,N_6540);
xnor U6661 (N_6661,N_6593,N_6621);
xor U6662 (N_6662,N_6581,N_6504);
or U6663 (N_6663,N_6587,N_6518);
nor U6664 (N_6664,N_6505,N_6544);
and U6665 (N_6665,N_6607,N_6512);
or U6666 (N_6666,N_6610,N_6620);
nand U6667 (N_6667,N_6551,N_6545);
xnor U6668 (N_6668,N_6558,N_6547);
and U6669 (N_6669,N_6554,N_6572);
nand U6670 (N_6670,N_6594,N_6564);
xor U6671 (N_6671,N_6546,N_6598);
or U6672 (N_6672,N_6612,N_6611);
or U6673 (N_6673,N_6535,N_6592);
nand U6674 (N_6674,N_6599,N_6575);
or U6675 (N_6675,N_6582,N_6591);
nor U6676 (N_6676,N_6579,N_6623);
xor U6677 (N_6677,N_6519,N_6536);
or U6678 (N_6678,N_6509,N_6541);
nor U6679 (N_6679,N_6520,N_6597);
nand U6680 (N_6680,N_6566,N_6571);
nor U6681 (N_6681,N_6560,N_6585);
nand U6682 (N_6682,N_6514,N_6595);
nor U6683 (N_6683,N_6552,N_6584);
xnor U6684 (N_6684,N_6569,N_6583);
nor U6685 (N_6685,N_6529,N_6586);
nand U6686 (N_6686,N_6537,N_6559);
and U6687 (N_6687,N_6525,N_6600);
and U6688 (N_6688,N_6540,N_6550);
and U6689 (N_6689,N_6582,N_6529);
nand U6690 (N_6690,N_6582,N_6608);
or U6691 (N_6691,N_6594,N_6588);
nor U6692 (N_6692,N_6583,N_6551);
xnor U6693 (N_6693,N_6618,N_6586);
nand U6694 (N_6694,N_6564,N_6601);
or U6695 (N_6695,N_6617,N_6564);
and U6696 (N_6696,N_6620,N_6609);
nor U6697 (N_6697,N_6611,N_6535);
and U6698 (N_6698,N_6610,N_6549);
xor U6699 (N_6699,N_6604,N_6505);
xnor U6700 (N_6700,N_6620,N_6579);
and U6701 (N_6701,N_6521,N_6526);
nand U6702 (N_6702,N_6500,N_6593);
or U6703 (N_6703,N_6618,N_6584);
xnor U6704 (N_6704,N_6608,N_6562);
nor U6705 (N_6705,N_6519,N_6558);
or U6706 (N_6706,N_6559,N_6512);
or U6707 (N_6707,N_6621,N_6602);
and U6708 (N_6708,N_6556,N_6534);
or U6709 (N_6709,N_6547,N_6540);
nor U6710 (N_6710,N_6592,N_6534);
or U6711 (N_6711,N_6574,N_6597);
xor U6712 (N_6712,N_6532,N_6582);
xnor U6713 (N_6713,N_6504,N_6574);
nor U6714 (N_6714,N_6611,N_6508);
nand U6715 (N_6715,N_6622,N_6556);
or U6716 (N_6716,N_6614,N_6503);
nand U6717 (N_6717,N_6535,N_6603);
nand U6718 (N_6718,N_6613,N_6556);
or U6719 (N_6719,N_6612,N_6607);
nor U6720 (N_6720,N_6615,N_6581);
nor U6721 (N_6721,N_6523,N_6553);
or U6722 (N_6722,N_6508,N_6592);
or U6723 (N_6723,N_6598,N_6525);
nand U6724 (N_6724,N_6615,N_6529);
nand U6725 (N_6725,N_6528,N_6592);
nand U6726 (N_6726,N_6597,N_6590);
nand U6727 (N_6727,N_6548,N_6523);
nand U6728 (N_6728,N_6541,N_6621);
nand U6729 (N_6729,N_6531,N_6621);
and U6730 (N_6730,N_6549,N_6584);
nor U6731 (N_6731,N_6582,N_6603);
nor U6732 (N_6732,N_6525,N_6583);
and U6733 (N_6733,N_6541,N_6558);
or U6734 (N_6734,N_6556,N_6603);
and U6735 (N_6735,N_6588,N_6616);
and U6736 (N_6736,N_6543,N_6624);
or U6737 (N_6737,N_6511,N_6550);
or U6738 (N_6738,N_6615,N_6541);
or U6739 (N_6739,N_6590,N_6522);
and U6740 (N_6740,N_6524,N_6556);
nand U6741 (N_6741,N_6595,N_6574);
nand U6742 (N_6742,N_6607,N_6541);
nor U6743 (N_6743,N_6562,N_6565);
and U6744 (N_6744,N_6537,N_6529);
and U6745 (N_6745,N_6579,N_6503);
and U6746 (N_6746,N_6550,N_6576);
and U6747 (N_6747,N_6565,N_6571);
nor U6748 (N_6748,N_6539,N_6501);
or U6749 (N_6749,N_6563,N_6562);
nor U6750 (N_6750,N_6683,N_6702);
and U6751 (N_6751,N_6738,N_6639);
xnor U6752 (N_6752,N_6636,N_6642);
nand U6753 (N_6753,N_6696,N_6736);
xnor U6754 (N_6754,N_6716,N_6731);
or U6755 (N_6755,N_6632,N_6704);
nand U6756 (N_6756,N_6643,N_6633);
nand U6757 (N_6757,N_6697,N_6688);
nand U6758 (N_6758,N_6725,N_6705);
nand U6759 (N_6759,N_6637,N_6666);
xor U6760 (N_6760,N_6734,N_6682);
or U6761 (N_6761,N_6733,N_6739);
nand U6762 (N_6762,N_6692,N_6654);
xnor U6763 (N_6763,N_6680,N_6651);
nand U6764 (N_6764,N_6742,N_6628);
nor U6765 (N_6765,N_6719,N_6690);
nand U6766 (N_6766,N_6700,N_6741);
and U6767 (N_6767,N_6701,N_6689);
nand U6768 (N_6768,N_6687,N_6706);
xnor U6769 (N_6769,N_6652,N_6629);
nor U6770 (N_6770,N_6747,N_6743);
nor U6771 (N_6771,N_6723,N_6685);
nor U6772 (N_6772,N_6727,N_6711);
nor U6773 (N_6773,N_6678,N_6679);
or U6774 (N_6774,N_6693,N_6648);
nor U6775 (N_6775,N_6658,N_6667);
nor U6776 (N_6776,N_6634,N_6710);
nand U6777 (N_6777,N_6681,N_6640);
and U6778 (N_6778,N_6674,N_6684);
nand U6779 (N_6779,N_6712,N_6703);
or U6780 (N_6780,N_6669,N_6728);
and U6781 (N_6781,N_6745,N_6670);
nor U6782 (N_6782,N_6677,N_6714);
nor U6783 (N_6783,N_6661,N_6708);
xor U6784 (N_6784,N_6645,N_6732);
nand U6785 (N_6785,N_6656,N_6724);
xor U6786 (N_6786,N_6748,N_6744);
and U6787 (N_6787,N_6746,N_6653);
nand U6788 (N_6788,N_6707,N_6635);
xor U6789 (N_6789,N_6631,N_6627);
or U6790 (N_6790,N_6717,N_6647);
or U6791 (N_6791,N_6676,N_6662);
xor U6792 (N_6792,N_6650,N_6649);
nor U6793 (N_6793,N_6722,N_6665);
nor U6794 (N_6794,N_6668,N_6646);
or U6795 (N_6795,N_6720,N_6673);
and U6796 (N_6796,N_6721,N_6625);
nand U6797 (N_6797,N_6663,N_6672);
nor U6798 (N_6798,N_6675,N_6730);
nor U6799 (N_6799,N_6709,N_6749);
nor U6800 (N_6800,N_6671,N_6715);
nor U6801 (N_6801,N_6664,N_6737);
xor U6802 (N_6802,N_6735,N_6740);
nand U6803 (N_6803,N_6626,N_6694);
xnor U6804 (N_6804,N_6644,N_6713);
nand U6805 (N_6805,N_6698,N_6630);
or U6806 (N_6806,N_6726,N_6641);
nor U6807 (N_6807,N_6655,N_6691);
nand U6808 (N_6808,N_6699,N_6686);
or U6809 (N_6809,N_6657,N_6659);
nor U6810 (N_6810,N_6638,N_6695);
and U6811 (N_6811,N_6718,N_6729);
nand U6812 (N_6812,N_6660,N_6746);
and U6813 (N_6813,N_6688,N_6647);
xnor U6814 (N_6814,N_6749,N_6730);
nor U6815 (N_6815,N_6702,N_6735);
nor U6816 (N_6816,N_6735,N_6749);
xor U6817 (N_6817,N_6628,N_6635);
nand U6818 (N_6818,N_6703,N_6744);
nor U6819 (N_6819,N_6626,N_6684);
or U6820 (N_6820,N_6704,N_6732);
xnor U6821 (N_6821,N_6704,N_6747);
nor U6822 (N_6822,N_6692,N_6684);
or U6823 (N_6823,N_6743,N_6692);
and U6824 (N_6824,N_6668,N_6645);
xor U6825 (N_6825,N_6649,N_6733);
nand U6826 (N_6826,N_6707,N_6696);
nand U6827 (N_6827,N_6709,N_6661);
nor U6828 (N_6828,N_6638,N_6670);
xor U6829 (N_6829,N_6681,N_6725);
nor U6830 (N_6830,N_6724,N_6685);
xnor U6831 (N_6831,N_6729,N_6747);
and U6832 (N_6832,N_6682,N_6748);
nand U6833 (N_6833,N_6743,N_6707);
nand U6834 (N_6834,N_6705,N_6716);
nor U6835 (N_6835,N_6677,N_6642);
nand U6836 (N_6836,N_6641,N_6738);
or U6837 (N_6837,N_6648,N_6711);
nor U6838 (N_6838,N_6717,N_6712);
xor U6839 (N_6839,N_6678,N_6648);
or U6840 (N_6840,N_6712,N_6643);
or U6841 (N_6841,N_6683,N_6628);
xnor U6842 (N_6842,N_6728,N_6747);
nor U6843 (N_6843,N_6691,N_6644);
xnor U6844 (N_6844,N_6696,N_6631);
or U6845 (N_6845,N_6743,N_6640);
or U6846 (N_6846,N_6630,N_6725);
xnor U6847 (N_6847,N_6698,N_6711);
and U6848 (N_6848,N_6682,N_6726);
and U6849 (N_6849,N_6670,N_6662);
and U6850 (N_6850,N_6673,N_6669);
or U6851 (N_6851,N_6684,N_6709);
nor U6852 (N_6852,N_6683,N_6629);
and U6853 (N_6853,N_6728,N_6743);
nor U6854 (N_6854,N_6695,N_6697);
nand U6855 (N_6855,N_6646,N_6717);
nor U6856 (N_6856,N_6662,N_6658);
nand U6857 (N_6857,N_6632,N_6740);
nor U6858 (N_6858,N_6646,N_6725);
and U6859 (N_6859,N_6705,N_6744);
and U6860 (N_6860,N_6683,N_6692);
or U6861 (N_6861,N_6728,N_6644);
nand U6862 (N_6862,N_6676,N_6718);
and U6863 (N_6863,N_6659,N_6717);
or U6864 (N_6864,N_6708,N_6665);
or U6865 (N_6865,N_6718,N_6711);
xnor U6866 (N_6866,N_6712,N_6744);
nand U6867 (N_6867,N_6680,N_6683);
or U6868 (N_6868,N_6681,N_6657);
xnor U6869 (N_6869,N_6671,N_6735);
or U6870 (N_6870,N_6654,N_6704);
nor U6871 (N_6871,N_6743,N_6695);
nand U6872 (N_6872,N_6647,N_6660);
nor U6873 (N_6873,N_6700,N_6746);
and U6874 (N_6874,N_6676,N_6634);
and U6875 (N_6875,N_6850,N_6781);
xor U6876 (N_6876,N_6866,N_6801);
xnor U6877 (N_6877,N_6846,N_6822);
or U6878 (N_6878,N_6864,N_6754);
or U6879 (N_6879,N_6836,N_6751);
nand U6880 (N_6880,N_6793,N_6791);
nand U6881 (N_6881,N_6807,N_6845);
xnor U6882 (N_6882,N_6873,N_6863);
or U6883 (N_6883,N_6831,N_6756);
nand U6884 (N_6884,N_6800,N_6786);
or U6885 (N_6885,N_6853,N_6858);
nor U6886 (N_6886,N_6805,N_6811);
xnor U6887 (N_6887,N_6779,N_6799);
and U6888 (N_6888,N_6851,N_6762);
nand U6889 (N_6889,N_6788,N_6812);
nand U6890 (N_6890,N_6797,N_6780);
and U6891 (N_6891,N_6760,N_6827);
nand U6892 (N_6892,N_6871,N_6803);
and U6893 (N_6893,N_6839,N_6837);
nor U6894 (N_6894,N_6773,N_6813);
and U6895 (N_6895,N_6792,N_6774);
nor U6896 (N_6896,N_6809,N_6874);
nand U6897 (N_6897,N_6778,N_6772);
nand U6898 (N_6898,N_6757,N_6834);
xor U6899 (N_6899,N_6784,N_6828);
nor U6900 (N_6900,N_6767,N_6859);
xor U6901 (N_6901,N_6849,N_6794);
nor U6902 (N_6902,N_6798,N_6854);
and U6903 (N_6903,N_6769,N_6833);
or U6904 (N_6904,N_6872,N_6841);
or U6905 (N_6905,N_6771,N_6868);
xnor U6906 (N_6906,N_6840,N_6847);
and U6907 (N_6907,N_6856,N_6802);
or U6908 (N_6908,N_6870,N_6867);
or U6909 (N_6909,N_6775,N_6816);
nand U6910 (N_6910,N_6832,N_6796);
or U6911 (N_6911,N_6852,N_6843);
or U6912 (N_6912,N_6752,N_6844);
xnor U6913 (N_6913,N_6750,N_6776);
and U6914 (N_6914,N_6819,N_6830);
and U6915 (N_6915,N_6821,N_6765);
nand U6916 (N_6916,N_6804,N_6817);
and U6917 (N_6917,N_6810,N_6825);
nand U6918 (N_6918,N_6787,N_6824);
or U6919 (N_6919,N_6808,N_6758);
and U6920 (N_6920,N_6826,N_6764);
or U6921 (N_6921,N_6835,N_6770);
xnor U6922 (N_6922,N_6818,N_6869);
or U6923 (N_6923,N_6789,N_6838);
or U6924 (N_6924,N_6815,N_6782);
or U6925 (N_6925,N_6755,N_6783);
nand U6926 (N_6926,N_6814,N_6763);
nor U6927 (N_6927,N_6790,N_6857);
nor U6928 (N_6928,N_6768,N_6823);
or U6929 (N_6929,N_6820,N_6777);
nor U6930 (N_6930,N_6865,N_6842);
or U6931 (N_6931,N_6855,N_6862);
and U6932 (N_6932,N_6766,N_6806);
xnor U6933 (N_6933,N_6861,N_6795);
nand U6934 (N_6934,N_6848,N_6860);
or U6935 (N_6935,N_6759,N_6785);
nand U6936 (N_6936,N_6753,N_6761);
or U6937 (N_6937,N_6829,N_6843);
or U6938 (N_6938,N_6822,N_6782);
or U6939 (N_6939,N_6817,N_6860);
nor U6940 (N_6940,N_6792,N_6834);
nor U6941 (N_6941,N_6852,N_6761);
and U6942 (N_6942,N_6762,N_6803);
nand U6943 (N_6943,N_6851,N_6771);
nor U6944 (N_6944,N_6771,N_6857);
xor U6945 (N_6945,N_6776,N_6798);
nand U6946 (N_6946,N_6782,N_6780);
xnor U6947 (N_6947,N_6862,N_6789);
and U6948 (N_6948,N_6818,N_6769);
or U6949 (N_6949,N_6826,N_6830);
xnor U6950 (N_6950,N_6845,N_6775);
and U6951 (N_6951,N_6869,N_6852);
nor U6952 (N_6952,N_6836,N_6754);
xnor U6953 (N_6953,N_6857,N_6775);
nor U6954 (N_6954,N_6803,N_6792);
or U6955 (N_6955,N_6833,N_6834);
or U6956 (N_6956,N_6765,N_6772);
nor U6957 (N_6957,N_6770,N_6795);
xnor U6958 (N_6958,N_6811,N_6866);
nand U6959 (N_6959,N_6788,N_6851);
and U6960 (N_6960,N_6804,N_6816);
or U6961 (N_6961,N_6804,N_6787);
xor U6962 (N_6962,N_6831,N_6788);
nand U6963 (N_6963,N_6854,N_6824);
nand U6964 (N_6964,N_6787,N_6816);
or U6965 (N_6965,N_6859,N_6828);
xor U6966 (N_6966,N_6868,N_6866);
or U6967 (N_6967,N_6871,N_6800);
nand U6968 (N_6968,N_6813,N_6765);
xor U6969 (N_6969,N_6842,N_6861);
nand U6970 (N_6970,N_6789,N_6846);
xnor U6971 (N_6971,N_6811,N_6834);
xor U6972 (N_6972,N_6809,N_6797);
xnor U6973 (N_6973,N_6856,N_6787);
xor U6974 (N_6974,N_6759,N_6757);
nand U6975 (N_6975,N_6813,N_6791);
nor U6976 (N_6976,N_6834,N_6759);
nand U6977 (N_6977,N_6770,N_6768);
and U6978 (N_6978,N_6806,N_6837);
nor U6979 (N_6979,N_6783,N_6844);
or U6980 (N_6980,N_6765,N_6855);
xor U6981 (N_6981,N_6807,N_6861);
or U6982 (N_6982,N_6788,N_6857);
or U6983 (N_6983,N_6793,N_6816);
or U6984 (N_6984,N_6796,N_6868);
nor U6985 (N_6985,N_6844,N_6781);
or U6986 (N_6986,N_6754,N_6802);
and U6987 (N_6987,N_6823,N_6773);
nand U6988 (N_6988,N_6759,N_6825);
xor U6989 (N_6989,N_6816,N_6821);
nor U6990 (N_6990,N_6769,N_6845);
xnor U6991 (N_6991,N_6772,N_6854);
nor U6992 (N_6992,N_6810,N_6802);
nor U6993 (N_6993,N_6825,N_6756);
or U6994 (N_6994,N_6837,N_6855);
nor U6995 (N_6995,N_6854,N_6787);
nand U6996 (N_6996,N_6847,N_6803);
nand U6997 (N_6997,N_6832,N_6754);
nand U6998 (N_6998,N_6785,N_6823);
xnor U6999 (N_6999,N_6860,N_6836);
xnor U7000 (N_7000,N_6967,N_6923);
nor U7001 (N_7001,N_6986,N_6970);
or U7002 (N_7002,N_6945,N_6984);
nand U7003 (N_7003,N_6971,N_6951);
xnor U7004 (N_7004,N_6973,N_6911);
nand U7005 (N_7005,N_6940,N_6918);
or U7006 (N_7006,N_6987,N_6963);
nand U7007 (N_7007,N_6924,N_6976);
or U7008 (N_7008,N_6931,N_6978);
and U7009 (N_7009,N_6896,N_6959);
or U7010 (N_7010,N_6905,N_6889);
xor U7011 (N_7011,N_6972,N_6954);
and U7012 (N_7012,N_6899,N_6941);
xnor U7013 (N_7013,N_6916,N_6919);
and U7014 (N_7014,N_6937,N_6990);
and U7015 (N_7015,N_6944,N_6927);
and U7016 (N_7016,N_6961,N_6891);
and U7017 (N_7017,N_6878,N_6914);
xor U7018 (N_7018,N_6903,N_6932);
nor U7019 (N_7019,N_6991,N_6958);
nor U7020 (N_7020,N_6902,N_6892);
xnor U7021 (N_7021,N_6994,N_6881);
or U7022 (N_7022,N_6876,N_6955);
or U7023 (N_7023,N_6981,N_6894);
nor U7024 (N_7024,N_6960,N_6962);
nand U7025 (N_7025,N_6912,N_6925);
and U7026 (N_7026,N_6992,N_6922);
xor U7027 (N_7027,N_6883,N_6943);
nand U7028 (N_7028,N_6952,N_6920);
nand U7029 (N_7029,N_6977,N_6980);
nand U7030 (N_7030,N_6907,N_6948);
nand U7031 (N_7031,N_6880,N_6969);
or U7032 (N_7032,N_6938,N_6895);
xnor U7033 (N_7033,N_6926,N_6888);
nor U7034 (N_7034,N_6910,N_6930);
nand U7035 (N_7035,N_6996,N_6947);
nor U7036 (N_7036,N_6998,N_6921);
nor U7037 (N_7037,N_6949,N_6886);
nor U7038 (N_7038,N_6956,N_6939);
and U7039 (N_7039,N_6929,N_6928);
nor U7040 (N_7040,N_6898,N_6966);
nor U7041 (N_7041,N_6909,N_6884);
or U7042 (N_7042,N_6975,N_6974);
nand U7043 (N_7043,N_6936,N_6953);
nor U7044 (N_7044,N_6913,N_6900);
xor U7045 (N_7045,N_6950,N_6982);
or U7046 (N_7046,N_6879,N_6965);
nor U7047 (N_7047,N_6882,N_6893);
nor U7048 (N_7048,N_6964,N_6997);
nor U7049 (N_7049,N_6906,N_6890);
or U7050 (N_7050,N_6993,N_6968);
and U7051 (N_7051,N_6915,N_6935);
and U7052 (N_7052,N_6989,N_6877);
xnor U7053 (N_7053,N_6983,N_6901);
xnor U7054 (N_7054,N_6904,N_6957);
nand U7055 (N_7055,N_6933,N_6988);
or U7056 (N_7056,N_6897,N_6999);
xnor U7057 (N_7057,N_6917,N_6887);
xor U7058 (N_7058,N_6908,N_6875);
nor U7059 (N_7059,N_6885,N_6985);
or U7060 (N_7060,N_6942,N_6946);
xnor U7061 (N_7061,N_6979,N_6995);
and U7062 (N_7062,N_6934,N_6982);
or U7063 (N_7063,N_6896,N_6963);
and U7064 (N_7064,N_6903,N_6898);
xnor U7065 (N_7065,N_6959,N_6997);
nand U7066 (N_7066,N_6914,N_6888);
nand U7067 (N_7067,N_6906,N_6915);
and U7068 (N_7068,N_6876,N_6915);
or U7069 (N_7069,N_6979,N_6996);
or U7070 (N_7070,N_6964,N_6983);
nor U7071 (N_7071,N_6886,N_6881);
or U7072 (N_7072,N_6962,N_6997);
and U7073 (N_7073,N_6933,N_6969);
nand U7074 (N_7074,N_6909,N_6893);
or U7075 (N_7075,N_6971,N_6967);
xnor U7076 (N_7076,N_6999,N_6886);
xor U7077 (N_7077,N_6927,N_6875);
xnor U7078 (N_7078,N_6990,N_6881);
or U7079 (N_7079,N_6914,N_6998);
or U7080 (N_7080,N_6981,N_6996);
xnor U7081 (N_7081,N_6918,N_6979);
nand U7082 (N_7082,N_6901,N_6931);
and U7083 (N_7083,N_6972,N_6911);
and U7084 (N_7084,N_6997,N_6981);
nor U7085 (N_7085,N_6887,N_6945);
xor U7086 (N_7086,N_6895,N_6951);
xnor U7087 (N_7087,N_6971,N_6947);
xnor U7088 (N_7088,N_6933,N_6967);
and U7089 (N_7089,N_6957,N_6961);
xor U7090 (N_7090,N_6999,N_6899);
nand U7091 (N_7091,N_6959,N_6939);
nand U7092 (N_7092,N_6932,N_6886);
or U7093 (N_7093,N_6929,N_6912);
and U7094 (N_7094,N_6937,N_6989);
or U7095 (N_7095,N_6886,N_6912);
or U7096 (N_7096,N_6935,N_6980);
nand U7097 (N_7097,N_6907,N_6937);
nand U7098 (N_7098,N_6935,N_6880);
xor U7099 (N_7099,N_6972,N_6884);
and U7100 (N_7100,N_6976,N_6937);
or U7101 (N_7101,N_6886,N_6933);
xnor U7102 (N_7102,N_6960,N_6954);
nand U7103 (N_7103,N_6892,N_6951);
nand U7104 (N_7104,N_6994,N_6924);
or U7105 (N_7105,N_6949,N_6964);
nor U7106 (N_7106,N_6979,N_6900);
nand U7107 (N_7107,N_6906,N_6944);
and U7108 (N_7108,N_6932,N_6910);
xor U7109 (N_7109,N_6935,N_6978);
or U7110 (N_7110,N_6943,N_6980);
or U7111 (N_7111,N_6966,N_6942);
nand U7112 (N_7112,N_6981,N_6974);
nor U7113 (N_7113,N_6903,N_6982);
nor U7114 (N_7114,N_6890,N_6991);
nand U7115 (N_7115,N_6941,N_6901);
nand U7116 (N_7116,N_6880,N_6921);
nor U7117 (N_7117,N_6983,N_6912);
or U7118 (N_7118,N_6927,N_6918);
nand U7119 (N_7119,N_6905,N_6898);
xor U7120 (N_7120,N_6904,N_6986);
or U7121 (N_7121,N_6906,N_6899);
or U7122 (N_7122,N_6928,N_6913);
and U7123 (N_7123,N_6907,N_6920);
nor U7124 (N_7124,N_6934,N_6932);
and U7125 (N_7125,N_7117,N_7030);
nand U7126 (N_7126,N_7102,N_7013);
and U7127 (N_7127,N_7081,N_7111);
and U7128 (N_7128,N_7072,N_7113);
or U7129 (N_7129,N_7063,N_7060);
or U7130 (N_7130,N_7029,N_7124);
nor U7131 (N_7131,N_7059,N_7099);
nor U7132 (N_7132,N_7122,N_7032);
nor U7133 (N_7133,N_7014,N_7007);
nor U7134 (N_7134,N_7026,N_7076);
xor U7135 (N_7135,N_7039,N_7088);
and U7136 (N_7136,N_7078,N_7095);
and U7137 (N_7137,N_7002,N_7101);
xnor U7138 (N_7138,N_7045,N_7022);
and U7139 (N_7139,N_7091,N_7052);
and U7140 (N_7140,N_7004,N_7079);
or U7141 (N_7141,N_7087,N_7105);
and U7142 (N_7142,N_7061,N_7038);
xor U7143 (N_7143,N_7116,N_7018);
xnor U7144 (N_7144,N_7016,N_7056);
xor U7145 (N_7145,N_7068,N_7121);
nand U7146 (N_7146,N_7027,N_7009);
or U7147 (N_7147,N_7046,N_7083);
or U7148 (N_7148,N_7065,N_7057);
nand U7149 (N_7149,N_7067,N_7098);
nand U7150 (N_7150,N_7120,N_7097);
nand U7151 (N_7151,N_7048,N_7089);
nand U7152 (N_7152,N_7073,N_7110);
nor U7153 (N_7153,N_7090,N_7096);
nand U7154 (N_7154,N_7041,N_7010);
and U7155 (N_7155,N_7011,N_7006);
and U7156 (N_7156,N_7070,N_7103);
xnor U7157 (N_7157,N_7054,N_7031);
nand U7158 (N_7158,N_7023,N_7092);
nand U7159 (N_7159,N_7003,N_7008);
nand U7160 (N_7160,N_7084,N_7049);
and U7161 (N_7161,N_7104,N_7112);
or U7162 (N_7162,N_7050,N_7020);
and U7163 (N_7163,N_7034,N_7062);
nand U7164 (N_7164,N_7107,N_7055);
or U7165 (N_7165,N_7019,N_7025);
or U7166 (N_7166,N_7033,N_7035);
nand U7167 (N_7167,N_7024,N_7040);
xnor U7168 (N_7168,N_7047,N_7108);
nor U7169 (N_7169,N_7001,N_7042);
and U7170 (N_7170,N_7074,N_7000);
and U7171 (N_7171,N_7015,N_7100);
and U7172 (N_7172,N_7106,N_7005);
xor U7173 (N_7173,N_7071,N_7021);
xnor U7174 (N_7174,N_7080,N_7064);
nor U7175 (N_7175,N_7037,N_7119);
nand U7176 (N_7176,N_7069,N_7077);
or U7177 (N_7177,N_7053,N_7043);
or U7178 (N_7178,N_7085,N_7028);
or U7179 (N_7179,N_7075,N_7086);
or U7180 (N_7180,N_7066,N_7044);
nand U7181 (N_7181,N_7051,N_7123);
nor U7182 (N_7182,N_7036,N_7093);
xnor U7183 (N_7183,N_7115,N_7012);
nor U7184 (N_7184,N_7109,N_7017);
xor U7185 (N_7185,N_7118,N_7082);
nand U7186 (N_7186,N_7094,N_7058);
or U7187 (N_7187,N_7114,N_7063);
xor U7188 (N_7188,N_7112,N_7122);
or U7189 (N_7189,N_7050,N_7073);
and U7190 (N_7190,N_7010,N_7110);
xnor U7191 (N_7191,N_7034,N_7063);
nor U7192 (N_7192,N_7114,N_7079);
nor U7193 (N_7193,N_7124,N_7123);
nand U7194 (N_7194,N_7016,N_7062);
or U7195 (N_7195,N_7097,N_7072);
or U7196 (N_7196,N_7050,N_7104);
xor U7197 (N_7197,N_7075,N_7056);
and U7198 (N_7198,N_7102,N_7104);
or U7199 (N_7199,N_7022,N_7120);
nand U7200 (N_7200,N_7059,N_7104);
nor U7201 (N_7201,N_7023,N_7042);
xor U7202 (N_7202,N_7086,N_7004);
or U7203 (N_7203,N_7062,N_7071);
nor U7204 (N_7204,N_7007,N_7054);
nor U7205 (N_7205,N_7116,N_7110);
and U7206 (N_7206,N_7121,N_7056);
xor U7207 (N_7207,N_7052,N_7119);
or U7208 (N_7208,N_7062,N_7107);
and U7209 (N_7209,N_7110,N_7074);
and U7210 (N_7210,N_7085,N_7030);
or U7211 (N_7211,N_7038,N_7075);
and U7212 (N_7212,N_7091,N_7080);
xnor U7213 (N_7213,N_7008,N_7030);
nand U7214 (N_7214,N_7034,N_7042);
and U7215 (N_7215,N_7085,N_7078);
and U7216 (N_7216,N_7089,N_7046);
nor U7217 (N_7217,N_7042,N_7084);
or U7218 (N_7218,N_7054,N_7032);
nor U7219 (N_7219,N_7024,N_7044);
nand U7220 (N_7220,N_7102,N_7100);
nor U7221 (N_7221,N_7085,N_7018);
or U7222 (N_7222,N_7077,N_7104);
nand U7223 (N_7223,N_7018,N_7003);
xor U7224 (N_7224,N_7044,N_7005);
nand U7225 (N_7225,N_7034,N_7073);
or U7226 (N_7226,N_7020,N_7091);
nand U7227 (N_7227,N_7059,N_7107);
or U7228 (N_7228,N_7032,N_7022);
nand U7229 (N_7229,N_7124,N_7056);
nand U7230 (N_7230,N_7029,N_7022);
and U7231 (N_7231,N_7035,N_7039);
nand U7232 (N_7232,N_7077,N_7016);
and U7233 (N_7233,N_7090,N_7086);
nand U7234 (N_7234,N_7000,N_7003);
xor U7235 (N_7235,N_7100,N_7028);
and U7236 (N_7236,N_7040,N_7016);
and U7237 (N_7237,N_7008,N_7072);
or U7238 (N_7238,N_7093,N_7072);
nand U7239 (N_7239,N_7010,N_7002);
nor U7240 (N_7240,N_7118,N_7099);
xnor U7241 (N_7241,N_7011,N_7046);
xnor U7242 (N_7242,N_7040,N_7089);
and U7243 (N_7243,N_7045,N_7047);
xnor U7244 (N_7244,N_7013,N_7112);
or U7245 (N_7245,N_7123,N_7004);
nor U7246 (N_7246,N_7058,N_7042);
or U7247 (N_7247,N_7037,N_7026);
xor U7248 (N_7248,N_7090,N_7056);
xor U7249 (N_7249,N_7070,N_7035);
xnor U7250 (N_7250,N_7152,N_7193);
nand U7251 (N_7251,N_7206,N_7203);
or U7252 (N_7252,N_7169,N_7238);
and U7253 (N_7253,N_7146,N_7153);
nand U7254 (N_7254,N_7142,N_7199);
nor U7255 (N_7255,N_7231,N_7191);
nor U7256 (N_7256,N_7167,N_7148);
nand U7257 (N_7257,N_7149,N_7233);
nand U7258 (N_7258,N_7130,N_7134);
nor U7259 (N_7259,N_7219,N_7150);
nor U7260 (N_7260,N_7245,N_7144);
or U7261 (N_7261,N_7241,N_7248);
nand U7262 (N_7262,N_7177,N_7176);
nor U7263 (N_7263,N_7125,N_7202);
nor U7264 (N_7264,N_7154,N_7208);
nand U7265 (N_7265,N_7147,N_7174);
or U7266 (N_7266,N_7159,N_7247);
nor U7267 (N_7267,N_7216,N_7249);
nor U7268 (N_7268,N_7242,N_7166);
nor U7269 (N_7269,N_7151,N_7237);
nor U7270 (N_7270,N_7162,N_7239);
or U7271 (N_7271,N_7225,N_7197);
and U7272 (N_7272,N_7129,N_7164);
nand U7273 (N_7273,N_7223,N_7186);
or U7274 (N_7274,N_7195,N_7133);
xor U7275 (N_7275,N_7183,N_7209);
xor U7276 (N_7276,N_7160,N_7243);
nand U7277 (N_7277,N_7132,N_7220);
nor U7278 (N_7278,N_7218,N_7180);
nand U7279 (N_7279,N_7141,N_7187);
or U7280 (N_7280,N_7131,N_7145);
nor U7281 (N_7281,N_7217,N_7228);
nand U7282 (N_7282,N_7236,N_7221);
xor U7283 (N_7283,N_7158,N_7196);
nand U7284 (N_7284,N_7173,N_7207);
or U7285 (N_7285,N_7212,N_7179);
and U7286 (N_7286,N_7213,N_7165);
nor U7287 (N_7287,N_7240,N_7184);
nor U7288 (N_7288,N_7214,N_7234);
xnor U7289 (N_7289,N_7136,N_7198);
or U7290 (N_7290,N_7188,N_7126);
nor U7291 (N_7291,N_7224,N_7200);
or U7292 (N_7292,N_7227,N_7232);
or U7293 (N_7293,N_7192,N_7222);
nor U7294 (N_7294,N_7171,N_7190);
or U7295 (N_7295,N_7127,N_7175);
xnor U7296 (N_7296,N_7143,N_7229);
xnor U7297 (N_7297,N_7140,N_7181);
nor U7298 (N_7298,N_7178,N_7246);
nand U7299 (N_7299,N_7163,N_7189);
xnor U7300 (N_7300,N_7155,N_7172);
xor U7301 (N_7301,N_7156,N_7157);
nand U7302 (N_7302,N_7205,N_7210);
nor U7303 (N_7303,N_7137,N_7201);
nor U7304 (N_7304,N_7170,N_7204);
or U7305 (N_7305,N_7182,N_7135);
xnor U7306 (N_7306,N_7194,N_7185);
and U7307 (N_7307,N_7211,N_7230);
xor U7308 (N_7308,N_7128,N_7161);
nand U7309 (N_7309,N_7138,N_7235);
nand U7310 (N_7310,N_7215,N_7226);
xnor U7311 (N_7311,N_7139,N_7244);
nor U7312 (N_7312,N_7168,N_7223);
nand U7313 (N_7313,N_7151,N_7185);
xor U7314 (N_7314,N_7233,N_7194);
nor U7315 (N_7315,N_7243,N_7209);
nor U7316 (N_7316,N_7226,N_7143);
nor U7317 (N_7317,N_7201,N_7170);
nand U7318 (N_7318,N_7130,N_7216);
or U7319 (N_7319,N_7182,N_7222);
or U7320 (N_7320,N_7167,N_7241);
xnor U7321 (N_7321,N_7207,N_7179);
nand U7322 (N_7322,N_7188,N_7164);
nand U7323 (N_7323,N_7130,N_7220);
and U7324 (N_7324,N_7220,N_7128);
xor U7325 (N_7325,N_7129,N_7234);
nor U7326 (N_7326,N_7148,N_7153);
or U7327 (N_7327,N_7174,N_7189);
and U7328 (N_7328,N_7182,N_7168);
nor U7329 (N_7329,N_7247,N_7220);
nor U7330 (N_7330,N_7207,N_7229);
and U7331 (N_7331,N_7126,N_7179);
and U7332 (N_7332,N_7153,N_7195);
nor U7333 (N_7333,N_7206,N_7134);
xnor U7334 (N_7334,N_7246,N_7148);
xor U7335 (N_7335,N_7240,N_7149);
nor U7336 (N_7336,N_7169,N_7209);
or U7337 (N_7337,N_7197,N_7178);
and U7338 (N_7338,N_7167,N_7192);
xor U7339 (N_7339,N_7141,N_7181);
nor U7340 (N_7340,N_7180,N_7184);
nand U7341 (N_7341,N_7205,N_7219);
nand U7342 (N_7342,N_7127,N_7242);
nand U7343 (N_7343,N_7213,N_7126);
nand U7344 (N_7344,N_7199,N_7222);
nand U7345 (N_7345,N_7217,N_7166);
or U7346 (N_7346,N_7192,N_7133);
nor U7347 (N_7347,N_7216,N_7212);
and U7348 (N_7348,N_7229,N_7152);
or U7349 (N_7349,N_7226,N_7242);
and U7350 (N_7350,N_7220,N_7186);
or U7351 (N_7351,N_7218,N_7173);
xnor U7352 (N_7352,N_7171,N_7137);
xor U7353 (N_7353,N_7206,N_7211);
xnor U7354 (N_7354,N_7159,N_7237);
or U7355 (N_7355,N_7132,N_7165);
or U7356 (N_7356,N_7232,N_7195);
xnor U7357 (N_7357,N_7228,N_7246);
nor U7358 (N_7358,N_7168,N_7148);
nand U7359 (N_7359,N_7133,N_7223);
and U7360 (N_7360,N_7237,N_7155);
or U7361 (N_7361,N_7187,N_7234);
nor U7362 (N_7362,N_7216,N_7168);
xor U7363 (N_7363,N_7199,N_7143);
or U7364 (N_7364,N_7200,N_7125);
nor U7365 (N_7365,N_7227,N_7243);
or U7366 (N_7366,N_7145,N_7222);
and U7367 (N_7367,N_7163,N_7227);
and U7368 (N_7368,N_7225,N_7181);
nand U7369 (N_7369,N_7155,N_7209);
xnor U7370 (N_7370,N_7248,N_7136);
xnor U7371 (N_7371,N_7153,N_7138);
nand U7372 (N_7372,N_7145,N_7198);
nand U7373 (N_7373,N_7217,N_7153);
nand U7374 (N_7374,N_7197,N_7238);
nand U7375 (N_7375,N_7274,N_7339);
or U7376 (N_7376,N_7336,N_7338);
nand U7377 (N_7377,N_7347,N_7314);
nor U7378 (N_7378,N_7353,N_7273);
and U7379 (N_7379,N_7333,N_7348);
and U7380 (N_7380,N_7346,N_7351);
or U7381 (N_7381,N_7253,N_7308);
xor U7382 (N_7382,N_7312,N_7278);
nand U7383 (N_7383,N_7309,N_7321);
xnor U7384 (N_7384,N_7355,N_7259);
nand U7385 (N_7385,N_7256,N_7254);
or U7386 (N_7386,N_7287,N_7330);
xnor U7387 (N_7387,N_7334,N_7335);
or U7388 (N_7388,N_7266,N_7272);
xor U7389 (N_7389,N_7320,N_7257);
nor U7390 (N_7390,N_7306,N_7297);
or U7391 (N_7391,N_7362,N_7284);
and U7392 (N_7392,N_7275,N_7269);
nand U7393 (N_7393,N_7252,N_7327);
xnor U7394 (N_7394,N_7317,N_7326);
or U7395 (N_7395,N_7277,N_7303);
or U7396 (N_7396,N_7343,N_7307);
nor U7397 (N_7397,N_7315,N_7371);
and U7398 (N_7398,N_7370,N_7352);
and U7399 (N_7399,N_7270,N_7296);
xor U7400 (N_7400,N_7369,N_7301);
xnor U7401 (N_7401,N_7342,N_7285);
nor U7402 (N_7402,N_7286,N_7310);
nor U7403 (N_7403,N_7264,N_7304);
or U7404 (N_7404,N_7322,N_7368);
xnor U7405 (N_7405,N_7324,N_7271);
or U7406 (N_7406,N_7328,N_7276);
nand U7407 (N_7407,N_7354,N_7261);
or U7408 (N_7408,N_7292,N_7279);
or U7409 (N_7409,N_7318,N_7372);
xor U7410 (N_7410,N_7358,N_7356);
nand U7411 (N_7411,N_7265,N_7263);
nand U7412 (N_7412,N_7373,N_7300);
nor U7413 (N_7413,N_7337,N_7299);
xnor U7414 (N_7414,N_7282,N_7302);
nor U7415 (N_7415,N_7260,N_7250);
nor U7416 (N_7416,N_7350,N_7255);
and U7417 (N_7417,N_7367,N_7268);
nor U7418 (N_7418,N_7316,N_7313);
nand U7419 (N_7419,N_7364,N_7319);
or U7420 (N_7420,N_7283,N_7344);
nand U7421 (N_7421,N_7331,N_7349);
or U7422 (N_7422,N_7341,N_7288);
or U7423 (N_7423,N_7360,N_7329);
and U7424 (N_7424,N_7357,N_7345);
nor U7425 (N_7425,N_7363,N_7262);
or U7426 (N_7426,N_7325,N_7290);
nand U7427 (N_7427,N_7374,N_7366);
xnor U7428 (N_7428,N_7365,N_7295);
or U7429 (N_7429,N_7289,N_7305);
and U7430 (N_7430,N_7361,N_7251);
nand U7431 (N_7431,N_7359,N_7294);
nor U7432 (N_7432,N_7281,N_7291);
nand U7433 (N_7433,N_7258,N_7332);
xnor U7434 (N_7434,N_7298,N_7340);
and U7435 (N_7435,N_7323,N_7293);
xor U7436 (N_7436,N_7280,N_7267);
nand U7437 (N_7437,N_7311,N_7254);
xnor U7438 (N_7438,N_7324,N_7266);
and U7439 (N_7439,N_7306,N_7311);
or U7440 (N_7440,N_7252,N_7325);
xor U7441 (N_7441,N_7366,N_7307);
or U7442 (N_7442,N_7296,N_7373);
and U7443 (N_7443,N_7324,N_7286);
xor U7444 (N_7444,N_7307,N_7280);
and U7445 (N_7445,N_7250,N_7326);
or U7446 (N_7446,N_7302,N_7356);
and U7447 (N_7447,N_7254,N_7369);
or U7448 (N_7448,N_7345,N_7374);
nor U7449 (N_7449,N_7360,N_7263);
or U7450 (N_7450,N_7266,N_7295);
or U7451 (N_7451,N_7317,N_7350);
and U7452 (N_7452,N_7368,N_7254);
and U7453 (N_7453,N_7258,N_7294);
nand U7454 (N_7454,N_7263,N_7270);
xor U7455 (N_7455,N_7300,N_7259);
and U7456 (N_7456,N_7300,N_7273);
or U7457 (N_7457,N_7316,N_7284);
and U7458 (N_7458,N_7347,N_7309);
or U7459 (N_7459,N_7356,N_7372);
nand U7460 (N_7460,N_7298,N_7339);
xor U7461 (N_7461,N_7320,N_7270);
xnor U7462 (N_7462,N_7324,N_7366);
and U7463 (N_7463,N_7350,N_7277);
or U7464 (N_7464,N_7278,N_7317);
xor U7465 (N_7465,N_7316,N_7288);
and U7466 (N_7466,N_7356,N_7291);
nor U7467 (N_7467,N_7325,N_7324);
and U7468 (N_7468,N_7256,N_7353);
nand U7469 (N_7469,N_7269,N_7268);
or U7470 (N_7470,N_7305,N_7372);
and U7471 (N_7471,N_7327,N_7329);
xnor U7472 (N_7472,N_7252,N_7330);
or U7473 (N_7473,N_7318,N_7274);
nor U7474 (N_7474,N_7327,N_7299);
xor U7475 (N_7475,N_7346,N_7348);
nor U7476 (N_7476,N_7323,N_7257);
and U7477 (N_7477,N_7261,N_7352);
nor U7478 (N_7478,N_7351,N_7308);
and U7479 (N_7479,N_7326,N_7336);
or U7480 (N_7480,N_7278,N_7293);
nand U7481 (N_7481,N_7308,N_7336);
nor U7482 (N_7482,N_7269,N_7316);
nand U7483 (N_7483,N_7355,N_7289);
and U7484 (N_7484,N_7284,N_7312);
xor U7485 (N_7485,N_7352,N_7292);
nand U7486 (N_7486,N_7374,N_7256);
nor U7487 (N_7487,N_7364,N_7336);
and U7488 (N_7488,N_7328,N_7345);
nor U7489 (N_7489,N_7263,N_7303);
xor U7490 (N_7490,N_7259,N_7312);
nor U7491 (N_7491,N_7280,N_7293);
nor U7492 (N_7492,N_7261,N_7304);
xnor U7493 (N_7493,N_7352,N_7307);
and U7494 (N_7494,N_7280,N_7276);
xor U7495 (N_7495,N_7290,N_7304);
and U7496 (N_7496,N_7349,N_7374);
nor U7497 (N_7497,N_7316,N_7252);
xnor U7498 (N_7498,N_7289,N_7259);
or U7499 (N_7499,N_7325,N_7354);
xor U7500 (N_7500,N_7448,N_7389);
nor U7501 (N_7501,N_7475,N_7405);
nor U7502 (N_7502,N_7481,N_7396);
nor U7503 (N_7503,N_7421,N_7466);
nor U7504 (N_7504,N_7388,N_7473);
nor U7505 (N_7505,N_7441,N_7447);
xor U7506 (N_7506,N_7399,N_7476);
nand U7507 (N_7507,N_7437,N_7387);
or U7508 (N_7508,N_7495,N_7402);
nand U7509 (N_7509,N_7436,N_7425);
nor U7510 (N_7510,N_7455,N_7403);
xnor U7511 (N_7511,N_7468,N_7496);
xnor U7512 (N_7512,N_7412,N_7477);
nand U7513 (N_7513,N_7414,N_7428);
nand U7514 (N_7514,N_7451,N_7452);
and U7515 (N_7515,N_7419,N_7493);
xor U7516 (N_7516,N_7486,N_7462);
xnor U7517 (N_7517,N_7406,N_7482);
and U7518 (N_7518,N_7409,N_7456);
nor U7519 (N_7519,N_7424,N_7478);
and U7520 (N_7520,N_7398,N_7383);
or U7521 (N_7521,N_7483,N_7384);
and U7522 (N_7522,N_7434,N_7465);
xor U7523 (N_7523,N_7407,N_7458);
and U7524 (N_7524,N_7498,N_7435);
and U7525 (N_7525,N_7394,N_7479);
and U7526 (N_7526,N_7440,N_7385);
xor U7527 (N_7527,N_7461,N_7491);
nor U7528 (N_7528,N_7463,N_7490);
nor U7529 (N_7529,N_7431,N_7420);
nand U7530 (N_7530,N_7433,N_7469);
xnor U7531 (N_7531,N_7392,N_7485);
nor U7532 (N_7532,N_7376,N_7472);
xnor U7533 (N_7533,N_7497,N_7422);
or U7534 (N_7534,N_7415,N_7454);
and U7535 (N_7535,N_7400,N_7442);
xor U7536 (N_7536,N_7457,N_7378);
or U7537 (N_7537,N_7423,N_7459);
nor U7538 (N_7538,N_7449,N_7386);
nand U7539 (N_7539,N_7474,N_7411);
nor U7540 (N_7540,N_7489,N_7438);
or U7541 (N_7541,N_7418,N_7480);
or U7542 (N_7542,N_7426,N_7471);
or U7543 (N_7543,N_7395,N_7382);
or U7544 (N_7544,N_7499,N_7375);
nand U7545 (N_7545,N_7381,N_7429);
or U7546 (N_7546,N_7377,N_7380);
xnor U7547 (N_7547,N_7467,N_7416);
nor U7548 (N_7548,N_7444,N_7445);
or U7549 (N_7549,N_7390,N_7401);
and U7550 (N_7550,N_7410,N_7487);
or U7551 (N_7551,N_7470,N_7393);
and U7552 (N_7552,N_7430,N_7391);
xor U7553 (N_7553,N_7488,N_7494);
and U7554 (N_7554,N_7417,N_7413);
nor U7555 (N_7555,N_7379,N_7427);
nand U7556 (N_7556,N_7492,N_7484);
xnor U7557 (N_7557,N_7432,N_7453);
or U7558 (N_7558,N_7464,N_7408);
nor U7559 (N_7559,N_7404,N_7439);
xnor U7560 (N_7560,N_7450,N_7443);
nor U7561 (N_7561,N_7446,N_7460);
nand U7562 (N_7562,N_7397,N_7476);
nand U7563 (N_7563,N_7461,N_7437);
nor U7564 (N_7564,N_7459,N_7413);
nor U7565 (N_7565,N_7444,N_7420);
nor U7566 (N_7566,N_7492,N_7440);
xnor U7567 (N_7567,N_7379,N_7407);
xor U7568 (N_7568,N_7455,N_7453);
and U7569 (N_7569,N_7399,N_7443);
xnor U7570 (N_7570,N_7383,N_7457);
xor U7571 (N_7571,N_7424,N_7474);
and U7572 (N_7572,N_7460,N_7399);
xor U7573 (N_7573,N_7462,N_7481);
xnor U7574 (N_7574,N_7403,N_7460);
nand U7575 (N_7575,N_7489,N_7490);
nor U7576 (N_7576,N_7461,N_7452);
nor U7577 (N_7577,N_7393,N_7394);
and U7578 (N_7578,N_7417,N_7431);
and U7579 (N_7579,N_7471,N_7458);
xnor U7580 (N_7580,N_7376,N_7397);
nor U7581 (N_7581,N_7460,N_7433);
or U7582 (N_7582,N_7493,N_7376);
xor U7583 (N_7583,N_7402,N_7440);
nand U7584 (N_7584,N_7444,N_7440);
xnor U7585 (N_7585,N_7375,N_7393);
nor U7586 (N_7586,N_7452,N_7396);
and U7587 (N_7587,N_7389,N_7440);
or U7588 (N_7588,N_7399,N_7455);
or U7589 (N_7589,N_7496,N_7461);
xnor U7590 (N_7590,N_7450,N_7387);
xnor U7591 (N_7591,N_7435,N_7405);
or U7592 (N_7592,N_7399,N_7432);
xor U7593 (N_7593,N_7404,N_7472);
xor U7594 (N_7594,N_7411,N_7405);
and U7595 (N_7595,N_7477,N_7446);
nor U7596 (N_7596,N_7453,N_7401);
and U7597 (N_7597,N_7402,N_7408);
or U7598 (N_7598,N_7411,N_7480);
and U7599 (N_7599,N_7403,N_7466);
nor U7600 (N_7600,N_7489,N_7386);
xnor U7601 (N_7601,N_7418,N_7388);
or U7602 (N_7602,N_7427,N_7433);
or U7603 (N_7603,N_7442,N_7449);
xor U7604 (N_7604,N_7439,N_7396);
xnor U7605 (N_7605,N_7489,N_7395);
or U7606 (N_7606,N_7431,N_7480);
and U7607 (N_7607,N_7475,N_7398);
and U7608 (N_7608,N_7479,N_7432);
nor U7609 (N_7609,N_7483,N_7462);
and U7610 (N_7610,N_7384,N_7376);
or U7611 (N_7611,N_7392,N_7499);
xnor U7612 (N_7612,N_7450,N_7445);
and U7613 (N_7613,N_7380,N_7455);
nand U7614 (N_7614,N_7479,N_7416);
and U7615 (N_7615,N_7405,N_7399);
nor U7616 (N_7616,N_7407,N_7488);
nand U7617 (N_7617,N_7412,N_7387);
nor U7618 (N_7618,N_7470,N_7380);
or U7619 (N_7619,N_7449,N_7389);
nor U7620 (N_7620,N_7448,N_7497);
and U7621 (N_7621,N_7418,N_7463);
and U7622 (N_7622,N_7494,N_7492);
xnor U7623 (N_7623,N_7418,N_7380);
xor U7624 (N_7624,N_7391,N_7411);
nor U7625 (N_7625,N_7547,N_7602);
nor U7626 (N_7626,N_7616,N_7504);
xnor U7627 (N_7627,N_7595,N_7578);
nor U7628 (N_7628,N_7560,N_7589);
and U7629 (N_7629,N_7550,N_7617);
and U7630 (N_7630,N_7603,N_7549);
nor U7631 (N_7631,N_7524,N_7606);
nor U7632 (N_7632,N_7597,N_7598);
or U7633 (N_7633,N_7613,N_7579);
or U7634 (N_7634,N_7588,N_7591);
nand U7635 (N_7635,N_7546,N_7577);
and U7636 (N_7636,N_7571,N_7565);
nor U7637 (N_7637,N_7516,N_7500);
or U7638 (N_7638,N_7580,N_7506);
and U7639 (N_7639,N_7584,N_7624);
nor U7640 (N_7640,N_7554,N_7545);
nor U7641 (N_7641,N_7505,N_7615);
nor U7642 (N_7642,N_7511,N_7618);
xnor U7643 (N_7643,N_7534,N_7590);
nor U7644 (N_7644,N_7502,N_7561);
and U7645 (N_7645,N_7523,N_7563);
nand U7646 (N_7646,N_7536,N_7576);
or U7647 (N_7647,N_7509,N_7513);
or U7648 (N_7648,N_7611,N_7537);
xnor U7649 (N_7649,N_7592,N_7558);
nand U7650 (N_7650,N_7512,N_7538);
and U7651 (N_7651,N_7553,N_7610);
and U7652 (N_7652,N_7583,N_7604);
nor U7653 (N_7653,N_7568,N_7530);
nor U7654 (N_7654,N_7501,N_7620);
xnor U7655 (N_7655,N_7562,N_7582);
nand U7656 (N_7656,N_7541,N_7612);
nand U7657 (N_7657,N_7569,N_7593);
and U7658 (N_7658,N_7559,N_7526);
nand U7659 (N_7659,N_7574,N_7544);
and U7660 (N_7660,N_7539,N_7529);
nor U7661 (N_7661,N_7535,N_7551);
xor U7662 (N_7662,N_7564,N_7542);
or U7663 (N_7663,N_7521,N_7514);
xnor U7664 (N_7664,N_7622,N_7596);
or U7665 (N_7665,N_7517,N_7581);
nand U7666 (N_7666,N_7525,N_7575);
and U7667 (N_7667,N_7557,N_7573);
or U7668 (N_7668,N_7540,N_7619);
xor U7669 (N_7669,N_7587,N_7572);
xnor U7670 (N_7670,N_7607,N_7510);
nor U7671 (N_7671,N_7543,N_7515);
and U7672 (N_7672,N_7519,N_7508);
nand U7673 (N_7673,N_7533,N_7520);
and U7674 (N_7674,N_7503,N_7522);
or U7675 (N_7675,N_7594,N_7555);
xnor U7676 (N_7676,N_7528,N_7601);
nor U7677 (N_7677,N_7566,N_7600);
nand U7678 (N_7678,N_7586,N_7531);
nor U7679 (N_7679,N_7556,N_7609);
nor U7680 (N_7680,N_7518,N_7552);
nand U7681 (N_7681,N_7527,N_7532);
nor U7682 (N_7682,N_7605,N_7623);
or U7683 (N_7683,N_7548,N_7621);
and U7684 (N_7684,N_7507,N_7567);
nand U7685 (N_7685,N_7608,N_7599);
nand U7686 (N_7686,N_7614,N_7585);
nand U7687 (N_7687,N_7570,N_7567);
xnor U7688 (N_7688,N_7503,N_7530);
nor U7689 (N_7689,N_7586,N_7553);
and U7690 (N_7690,N_7607,N_7579);
nor U7691 (N_7691,N_7544,N_7610);
or U7692 (N_7692,N_7550,N_7594);
xnor U7693 (N_7693,N_7606,N_7557);
and U7694 (N_7694,N_7563,N_7508);
and U7695 (N_7695,N_7578,N_7621);
or U7696 (N_7696,N_7601,N_7549);
nand U7697 (N_7697,N_7504,N_7615);
or U7698 (N_7698,N_7548,N_7603);
xor U7699 (N_7699,N_7527,N_7545);
xor U7700 (N_7700,N_7614,N_7623);
xnor U7701 (N_7701,N_7605,N_7580);
and U7702 (N_7702,N_7532,N_7549);
nor U7703 (N_7703,N_7554,N_7571);
nand U7704 (N_7704,N_7548,N_7570);
nor U7705 (N_7705,N_7593,N_7515);
xnor U7706 (N_7706,N_7598,N_7546);
nand U7707 (N_7707,N_7545,N_7579);
nand U7708 (N_7708,N_7591,N_7615);
nand U7709 (N_7709,N_7532,N_7541);
xor U7710 (N_7710,N_7607,N_7615);
xnor U7711 (N_7711,N_7568,N_7553);
or U7712 (N_7712,N_7538,N_7620);
nor U7713 (N_7713,N_7569,N_7532);
or U7714 (N_7714,N_7566,N_7583);
nand U7715 (N_7715,N_7613,N_7612);
nand U7716 (N_7716,N_7570,N_7547);
nor U7717 (N_7717,N_7585,N_7505);
nand U7718 (N_7718,N_7624,N_7591);
nand U7719 (N_7719,N_7603,N_7573);
and U7720 (N_7720,N_7545,N_7584);
and U7721 (N_7721,N_7530,N_7620);
nor U7722 (N_7722,N_7623,N_7508);
or U7723 (N_7723,N_7570,N_7541);
nor U7724 (N_7724,N_7502,N_7572);
nand U7725 (N_7725,N_7590,N_7567);
or U7726 (N_7726,N_7582,N_7623);
and U7727 (N_7727,N_7610,N_7515);
nand U7728 (N_7728,N_7569,N_7576);
nor U7729 (N_7729,N_7582,N_7616);
or U7730 (N_7730,N_7512,N_7603);
nand U7731 (N_7731,N_7563,N_7594);
xnor U7732 (N_7732,N_7555,N_7621);
nand U7733 (N_7733,N_7574,N_7612);
nand U7734 (N_7734,N_7605,N_7599);
nor U7735 (N_7735,N_7617,N_7547);
nor U7736 (N_7736,N_7606,N_7614);
and U7737 (N_7737,N_7623,N_7514);
and U7738 (N_7738,N_7555,N_7597);
and U7739 (N_7739,N_7537,N_7578);
and U7740 (N_7740,N_7525,N_7528);
or U7741 (N_7741,N_7508,N_7548);
nand U7742 (N_7742,N_7500,N_7542);
nand U7743 (N_7743,N_7547,N_7594);
nor U7744 (N_7744,N_7501,N_7609);
and U7745 (N_7745,N_7604,N_7592);
nor U7746 (N_7746,N_7575,N_7574);
nand U7747 (N_7747,N_7510,N_7606);
nor U7748 (N_7748,N_7585,N_7582);
and U7749 (N_7749,N_7587,N_7553);
or U7750 (N_7750,N_7668,N_7745);
nand U7751 (N_7751,N_7715,N_7641);
xnor U7752 (N_7752,N_7749,N_7684);
nand U7753 (N_7753,N_7645,N_7670);
nand U7754 (N_7754,N_7739,N_7646);
nand U7755 (N_7755,N_7706,N_7724);
nand U7756 (N_7756,N_7735,N_7673);
nor U7757 (N_7757,N_7644,N_7740);
and U7758 (N_7758,N_7719,N_7705);
nand U7759 (N_7759,N_7671,N_7675);
nor U7760 (N_7760,N_7703,N_7674);
xnor U7761 (N_7761,N_7662,N_7730);
nand U7762 (N_7762,N_7630,N_7710);
nand U7763 (N_7763,N_7738,N_7713);
or U7764 (N_7764,N_7744,N_7725);
nor U7765 (N_7765,N_7704,N_7702);
and U7766 (N_7766,N_7691,N_7690);
xor U7767 (N_7767,N_7692,N_7728);
nand U7768 (N_7768,N_7661,N_7732);
xor U7769 (N_7769,N_7741,N_7666);
nand U7770 (N_7770,N_7634,N_7748);
or U7771 (N_7771,N_7747,N_7627);
nor U7772 (N_7772,N_7685,N_7643);
nor U7773 (N_7773,N_7716,N_7676);
xor U7774 (N_7774,N_7625,N_7717);
xor U7775 (N_7775,N_7731,N_7681);
and U7776 (N_7776,N_7683,N_7648);
or U7777 (N_7777,N_7727,N_7726);
nand U7778 (N_7778,N_7631,N_7640);
xnor U7779 (N_7779,N_7654,N_7743);
xor U7780 (N_7780,N_7651,N_7711);
nand U7781 (N_7781,N_7687,N_7734);
nand U7782 (N_7782,N_7677,N_7686);
or U7783 (N_7783,N_7698,N_7678);
xnor U7784 (N_7784,N_7656,N_7655);
nor U7785 (N_7785,N_7720,N_7672);
nor U7786 (N_7786,N_7657,N_7707);
or U7787 (N_7787,N_7693,N_7628);
xor U7788 (N_7788,N_7697,N_7700);
and U7789 (N_7789,N_7701,N_7632);
xor U7790 (N_7790,N_7746,N_7729);
and U7791 (N_7791,N_7667,N_7708);
nand U7792 (N_7792,N_7647,N_7733);
or U7793 (N_7793,N_7723,N_7721);
nor U7794 (N_7794,N_7635,N_7742);
xnor U7795 (N_7795,N_7689,N_7688);
nor U7796 (N_7796,N_7638,N_7736);
xor U7797 (N_7797,N_7718,N_7649);
nand U7798 (N_7798,N_7737,N_7663);
nand U7799 (N_7799,N_7722,N_7650);
or U7800 (N_7800,N_7699,N_7665);
xor U7801 (N_7801,N_7682,N_7696);
nor U7802 (N_7802,N_7658,N_7639);
or U7803 (N_7803,N_7680,N_7712);
nor U7804 (N_7804,N_7660,N_7694);
or U7805 (N_7805,N_7642,N_7669);
or U7806 (N_7806,N_7653,N_7714);
xnor U7807 (N_7807,N_7637,N_7679);
nand U7808 (N_7808,N_7664,N_7636);
nand U7809 (N_7809,N_7709,N_7695);
xnor U7810 (N_7810,N_7652,N_7626);
or U7811 (N_7811,N_7629,N_7633);
and U7812 (N_7812,N_7659,N_7703);
and U7813 (N_7813,N_7701,N_7631);
and U7814 (N_7814,N_7734,N_7647);
and U7815 (N_7815,N_7628,N_7709);
or U7816 (N_7816,N_7635,N_7746);
nor U7817 (N_7817,N_7725,N_7661);
nand U7818 (N_7818,N_7651,N_7650);
nand U7819 (N_7819,N_7683,N_7635);
xnor U7820 (N_7820,N_7716,N_7691);
and U7821 (N_7821,N_7657,N_7626);
nand U7822 (N_7822,N_7643,N_7710);
xnor U7823 (N_7823,N_7626,N_7632);
xnor U7824 (N_7824,N_7671,N_7730);
nor U7825 (N_7825,N_7701,N_7671);
nand U7826 (N_7826,N_7713,N_7730);
xor U7827 (N_7827,N_7723,N_7703);
and U7828 (N_7828,N_7704,N_7743);
and U7829 (N_7829,N_7665,N_7688);
or U7830 (N_7830,N_7642,N_7738);
xnor U7831 (N_7831,N_7638,N_7640);
xor U7832 (N_7832,N_7648,N_7682);
nand U7833 (N_7833,N_7649,N_7727);
nor U7834 (N_7834,N_7683,N_7703);
nor U7835 (N_7835,N_7631,N_7638);
xnor U7836 (N_7836,N_7643,N_7627);
nor U7837 (N_7837,N_7640,N_7634);
and U7838 (N_7838,N_7741,N_7684);
nor U7839 (N_7839,N_7706,N_7679);
or U7840 (N_7840,N_7697,N_7632);
xor U7841 (N_7841,N_7690,N_7671);
and U7842 (N_7842,N_7632,N_7625);
and U7843 (N_7843,N_7738,N_7649);
and U7844 (N_7844,N_7728,N_7669);
or U7845 (N_7845,N_7713,N_7714);
nor U7846 (N_7846,N_7705,N_7714);
nor U7847 (N_7847,N_7713,N_7625);
nand U7848 (N_7848,N_7644,N_7718);
nor U7849 (N_7849,N_7727,N_7697);
or U7850 (N_7850,N_7656,N_7694);
xnor U7851 (N_7851,N_7636,N_7720);
and U7852 (N_7852,N_7636,N_7725);
or U7853 (N_7853,N_7662,N_7651);
nor U7854 (N_7854,N_7699,N_7660);
and U7855 (N_7855,N_7653,N_7701);
xor U7856 (N_7856,N_7639,N_7654);
or U7857 (N_7857,N_7733,N_7661);
nor U7858 (N_7858,N_7704,N_7656);
and U7859 (N_7859,N_7738,N_7690);
nor U7860 (N_7860,N_7697,N_7665);
and U7861 (N_7861,N_7729,N_7631);
nor U7862 (N_7862,N_7699,N_7729);
and U7863 (N_7863,N_7645,N_7693);
and U7864 (N_7864,N_7749,N_7727);
xor U7865 (N_7865,N_7649,N_7627);
xnor U7866 (N_7866,N_7646,N_7717);
or U7867 (N_7867,N_7673,N_7645);
xnor U7868 (N_7868,N_7740,N_7707);
nand U7869 (N_7869,N_7684,N_7743);
nor U7870 (N_7870,N_7673,N_7680);
and U7871 (N_7871,N_7655,N_7635);
and U7872 (N_7872,N_7659,N_7747);
or U7873 (N_7873,N_7721,N_7738);
nand U7874 (N_7874,N_7680,N_7674);
xnor U7875 (N_7875,N_7775,N_7800);
or U7876 (N_7876,N_7823,N_7752);
or U7877 (N_7877,N_7860,N_7785);
nor U7878 (N_7878,N_7806,N_7787);
nand U7879 (N_7879,N_7767,N_7788);
and U7880 (N_7880,N_7762,N_7814);
nand U7881 (N_7881,N_7850,N_7754);
nor U7882 (N_7882,N_7818,N_7851);
xnor U7883 (N_7883,N_7779,N_7786);
nand U7884 (N_7884,N_7870,N_7840);
nor U7885 (N_7885,N_7825,N_7854);
and U7886 (N_7886,N_7872,N_7821);
xnor U7887 (N_7887,N_7819,N_7764);
nor U7888 (N_7888,N_7833,N_7830);
and U7889 (N_7889,N_7862,N_7824);
nand U7890 (N_7890,N_7837,N_7780);
and U7891 (N_7891,N_7809,N_7865);
nand U7892 (N_7892,N_7797,N_7783);
nor U7893 (N_7893,N_7790,N_7864);
xor U7894 (N_7894,N_7772,N_7807);
nand U7895 (N_7895,N_7831,N_7753);
nand U7896 (N_7896,N_7855,N_7760);
and U7897 (N_7897,N_7750,N_7838);
or U7898 (N_7898,N_7852,N_7849);
and U7899 (N_7899,N_7756,N_7773);
xnor U7900 (N_7900,N_7816,N_7817);
xor U7901 (N_7901,N_7805,N_7808);
or U7902 (N_7902,N_7836,N_7869);
nand U7903 (N_7903,N_7846,N_7798);
nand U7904 (N_7904,N_7751,N_7863);
and U7905 (N_7905,N_7822,N_7845);
xnor U7906 (N_7906,N_7835,N_7802);
and U7907 (N_7907,N_7867,N_7874);
or U7908 (N_7908,N_7777,N_7792);
nand U7909 (N_7909,N_7858,N_7853);
xor U7910 (N_7910,N_7801,N_7843);
or U7911 (N_7911,N_7781,N_7861);
or U7912 (N_7912,N_7841,N_7866);
xnor U7913 (N_7913,N_7868,N_7782);
nand U7914 (N_7914,N_7810,N_7847);
xor U7915 (N_7915,N_7776,N_7848);
nor U7916 (N_7916,N_7761,N_7771);
xor U7917 (N_7917,N_7804,N_7795);
xor U7918 (N_7918,N_7844,N_7758);
nor U7919 (N_7919,N_7755,N_7856);
nand U7920 (N_7920,N_7796,N_7793);
xor U7921 (N_7921,N_7871,N_7832);
and U7922 (N_7922,N_7820,N_7759);
and U7923 (N_7923,N_7778,N_7811);
nor U7924 (N_7924,N_7769,N_7842);
xnor U7925 (N_7925,N_7763,N_7873);
and U7926 (N_7926,N_7789,N_7757);
or U7927 (N_7927,N_7794,N_7857);
xnor U7928 (N_7928,N_7815,N_7839);
or U7929 (N_7929,N_7784,N_7766);
nor U7930 (N_7930,N_7791,N_7828);
and U7931 (N_7931,N_7829,N_7834);
or U7932 (N_7932,N_7859,N_7770);
xor U7933 (N_7933,N_7765,N_7768);
nor U7934 (N_7934,N_7827,N_7799);
nor U7935 (N_7935,N_7813,N_7812);
nor U7936 (N_7936,N_7774,N_7826);
nand U7937 (N_7937,N_7803,N_7806);
xnor U7938 (N_7938,N_7762,N_7857);
xor U7939 (N_7939,N_7762,N_7828);
nand U7940 (N_7940,N_7790,N_7768);
xor U7941 (N_7941,N_7802,N_7856);
xnor U7942 (N_7942,N_7872,N_7837);
xor U7943 (N_7943,N_7773,N_7867);
nand U7944 (N_7944,N_7863,N_7782);
or U7945 (N_7945,N_7777,N_7822);
and U7946 (N_7946,N_7874,N_7856);
and U7947 (N_7947,N_7785,N_7827);
or U7948 (N_7948,N_7842,N_7756);
nor U7949 (N_7949,N_7824,N_7857);
and U7950 (N_7950,N_7786,N_7854);
nand U7951 (N_7951,N_7785,N_7850);
or U7952 (N_7952,N_7786,N_7845);
and U7953 (N_7953,N_7823,N_7757);
nor U7954 (N_7954,N_7815,N_7832);
or U7955 (N_7955,N_7816,N_7776);
nand U7956 (N_7956,N_7788,N_7783);
and U7957 (N_7957,N_7752,N_7779);
nand U7958 (N_7958,N_7789,N_7846);
nand U7959 (N_7959,N_7864,N_7834);
nor U7960 (N_7960,N_7834,N_7789);
nand U7961 (N_7961,N_7814,N_7842);
nand U7962 (N_7962,N_7851,N_7789);
nand U7963 (N_7963,N_7839,N_7832);
nand U7964 (N_7964,N_7757,N_7873);
xnor U7965 (N_7965,N_7801,N_7775);
nor U7966 (N_7966,N_7846,N_7775);
and U7967 (N_7967,N_7854,N_7819);
xnor U7968 (N_7968,N_7835,N_7849);
and U7969 (N_7969,N_7813,N_7872);
and U7970 (N_7970,N_7759,N_7756);
xor U7971 (N_7971,N_7852,N_7874);
and U7972 (N_7972,N_7861,N_7841);
and U7973 (N_7973,N_7816,N_7788);
and U7974 (N_7974,N_7794,N_7752);
xnor U7975 (N_7975,N_7764,N_7853);
or U7976 (N_7976,N_7770,N_7791);
xnor U7977 (N_7977,N_7851,N_7844);
or U7978 (N_7978,N_7781,N_7808);
nor U7979 (N_7979,N_7752,N_7843);
xor U7980 (N_7980,N_7833,N_7806);
nor U7981 (N_7981,N_7794,N_7866);
and U7982 (N_7982,N_7871,N_7830);
nor U7983 (N_7983,N_7820,N_7818);
and U7984 (N_7984,N_7806,N_7768);
xnor U7985 (N_7985,N_7797,N_7819);
xnor U7986 (N_7986,N_7835,N_7790);
xor U7987 (N_7987,N_7786,N_7823);
nor U7988 (N_7988,N_7853,N_7840);
nor U7989 (N_7989,N_7755,N_7873);
xor U7990 (N_7990,N_7784,N_7871);
and U7991 (N_7991,N_7751,N_7782);
and U7992 (N_7992,N_7820,N_7822);
and U7993 (N_7993,N_7826,N_7874);
nor U7994 (N_7994,N_7840,N_7790);
nand U7995 (N_7995,N_7800,N_7824);
and U7996 (N_7996,N_7792,N_7809);
or U7997 (N_7997,N_7822,N_7783);
nor U7998 (N_7998,N_7791,N_7845);
or U7999 (N_7999,N_7873,N_7855);
xnor U8000 (N_8000,N_7941,N_7894);
nand U8001 (N_8001,N_7918,N_7949);
nand U8002 (N_8002,N_7942,N_7904);
and U8003 (N_8003,N_7977,N_7952);
xor U8004 (N_8004,N_7939,N_7979);
nor U8005 (N_8005,N_7888,N_7994);
xnor U8006 (N_8006,N_7990,N_7876);
xnor U8007 (N_8007,N_7999,N_7922);
nor U8008 (N_8008,N_7954,N_7878);
or U8009 (N_8009,N_7946,N_7983);
or U8010 (N_8010,N_7956,N_7934);
or U8011 (N_8011,N_7961,N_7992);
nand U8012 (N_8012,N_7997,N_7884);
or U8013 (N_8013,N_7955,N_7899);
or U8014 (N_8014,N_7885,N_7987);
and U8015 (N_8015,N_7936,N_7959);
or U8016 (N_8016,N_7933,N_7938);
nand U8017 (N_8017,N_7917,N_7927);
nor U8018 (N_8018,N_7996,N_7879);
and U8019 (N_8019,N_7882,N_7893);
xnor U8020 (N_8020,N_7985,N_7912);
or U8021 (N_8021,N_7930,N_7953);
nand U8022 (N_8022,N_7906,N_7883);
and U8023 (N_8023,N_7892,N_7978);
or U8024 (N_8024,N_7980,N_7908);
and U8025 (N_8025,N_7982,N_7890);
xnor U8026 (N_8026,N_7937,N_7995);
nand U8027 (N_8027,N_7896,N_7931);
xor U8028 (N_8028,N_7969,N_7919);
or U8029 (N_8029,N_7898,N_7963);
xnor U8030 (N_8030,N_7993,N_7971);
nand U8031 (N_8031,N_7958,N_7901);
xor U8032 (N_8032,N_7966,N_7947);
or U8033 (N_8033,N_7932,N_7920);
nand U8034 (N_8034,N_7967,N_7875);
xnor U8035 (N_8035,N_7964,N_7921);
or U8036 (N_8036,N_7909,N_7903);
or U8037 (N_8037,N_7925,N_7905);
xor U8038 (N_8038,N_7910,N_7944);
nor U8039 (N_8039,N_7986,N_7897);
or U8040 (N_8040,N_7886,N_7887);
and U8041 (N_8041,N_7928,N_7972);
or U8042 (N_8042,N_7877,N_7965);
or U8043 (N_8043,N_7948,N_7924);
nor U8044 (N_8044,N_7907,N_7911);
xnor U8045 (N_8045,N_7957,N_7943);
xor U8046 (N_8046,N_7900,N_7988);
nand U8047 (N_8047,N_7926,N_7950);
or U8048 (N_8048,N_7975,N_7915);
and U8049 (N_8049,N_7935,N_7940);
nand U8050 (N_8050,N_7880,N_7984);
or U8051 (N_8051,N_7968,N_7914);
or U8052 (N_8052,N_7976,N_7991);
xor U8053 (N_8053,N_7913,N_7916);
xnor U8054 (N_8054,N_7881,N_7929);
nand U8055 (N_8055,N_7923,N_7998);
nand U8056 (N_8056,N_7970,N_7889);
nor U8057 (N_8057,N_7960,N_7973);
or U8058 (N_8058,N_7945,N_7951);
nand U8059 (N_8059,N_7989,N_7962);
xor U8060 (N_8060,N_7891,N_7902);
or U8061 (N_8061,N_7895,N_7974);
or U8062 (N_8062,N_7981,N_7956);
nand U8063 (N_8063,N_7917,N_7897);
or U8064 (N_8064,N_7993,N_7942);
nor U8065 (N_8065,N_7961,N_7902);
xor U8066 (N_8066,N_7945,N_7954);
or U8067 (N_8067,N_7879,N_7975);
nor U8068 (N_8068,N_7936,N_7894);
nor U8069 (N_8069,N_7920,N_7892);
nor U8070 (N_8070,N_7953,N_7996);
and U8071 (N_8071,N_7935,N_7981);
nand U8072 (N_8072,N_7923,N_7939);
nand U8073 (N_8073,N_7906,N_7994);
nor U8074 (N_8074,N_7953,N_7973);
nand U8075 (N_8075,N_7943,N_7893);
nand U8076 (N_8076,N_7905,N_7920);
nor U8077 (N_8077,N_7911,N_7942);
xnor U8078 (N_8078,N_7915,N_7997);
nor U8079 (N_8079,N_7935,N_7905);
nand U8080 (N_8080,N_7935,N_7919);
xor U8081 (N_8081,N_7926,N_7993);
nand U8082 (N_8082,N_7965,N_7959);
xnor U8083 (N_8083,N_7974,N_7883);
nand U8084 (N_8084,N_7912,N_7953);
nor U8085 (N_8085,N_7965,N_7941);
or U8086 (N_8086,N_7922,N_7961);
and U8087 (N_8087,N_7876,N_7894);
xor U8088 (N_8088,N_7946,N_7920);
nor U8089 (N_8089,N_7938,N_7971);
xnor U8090 (N_8090,N_7953,N_7944);
nor U8091 (N_8091,N_7969,N_7974);
nor U8092 (N_8092,N_7891,N_7887);
or U8093 (N_8093,N_7925,N_7994);
nor U8094 (N_8094,N_7919,N_7878);
nor U8095 (N_8095,N_7909,N_7961);
or U8096 (N_8096,N_7931,N_7921);
nor U8097 (N_8097,N_7898,N_7917);
nor U8098 (N_8098,N_7931,N_7962);
or U8099 (N_8099,N_7895,N_7969);
nor U8100 (N_8100,N_7913,N_7968);
or U8101 (N_8101,N_7958,N_7903);
nor U8102 (N_8102,N_7958,N_7924);
xor U8103 (N_8103,N_7980,N_7960);
nor U8104 (N_8104,N_7912,N_7904);
nor U8105 (N_8105,N_7993,N_7946);
or U8106 (N_8106,N_7879,N_7991);
nor U8107 (N_8107,N_7939,N_7889);
nor U8108 (N_8108,N_7890,N_7914);
nor U8109 (N_8109,N_7957,N_7992);
nor U8110 (N_8110,N_7987,N_7939);
or U8111 (N_8111,N_7903,N_7975);
and U8112 (N_8112,N_7939,N_7959);
xnor U8113 (N_8113,N_7915,N_7960);
or U8114 (N_8114,N_7995,N_7992);
nand U8115 (N_8115,N_7925,N_7897);
xor U8116 (N_8116,N_7882,N_7983);
xnor U8117 (N_8117,N_7989,N_7876);
or U8118 (N_8118,N_7895,N_7965);
or U8119 (N_8119,N_7960,N_7965);
or U8120 (N_8120,N_7918,N_7905);
xor U8121 (N_8121,N_7907,N_7881);
or U8122 (N_8122,N_7974,N_7938);
and U8123 (N_8123,N_7969,N_7910);
nor U8124 (N_8124,N_7927,N_7990);
and U8125 (N_8125,N_8083,N_8032);
or U8126 (N_8126,N_8036,N_8047);
nor U8127 (N_8127,N_8010,N_8035);
xor U8128 (N_8128,N_8018,N_8075);
xor U8129 (N_8129,N_8105,N_8085);
xor U8130 (N_8130,N_8012,N_8071);
nand U8131 (N_8131,N_8096,N_8052);
or U8132 (N_8132,N_8008,N_8122);
or U8133 (N_8133,N_8060,N_8123);
nor U8134 (N_8134,N_8033,N_8077);
xnor U8135 (N_8135,N_8084,N_8079);
xor U8136 (N_8136,N_8034,N_8061);
and U8137 (N_8137,N_8054,N_8062);
nand U8138 (N_8138,N_8022,N_8064);
xnor U8139 (N_8139,N_8037,N_8014);
or U8140 (N_8140,N_8049,N_8087);
or U8141 (N_8141,N_8103,N_8042);
nand U8142 (N_8142,N_8043,N_8058);
xnor U8143 (N_8143,N_8055,N_8073);
or U8144 (N_8144,N_8070,N_8082);
and U8145 (N_8145,N_8067,N_8039);
and U8146 (N_8146,N_8007,N_8050);
nand U8147 (N_8147,N_8066,N_8112);
nor U8148 (N_8148,N_8081,N_8013);
nand U8149 (N_8149,N_8053,N_8063);
nand U8150 (N_8150,N_8069,N_8000);
nor U8151 (N_8151,N_8030,N_8005);
or U8152 (N_8152,N_8102,N_8076);
nor U8153 (N_8153,N_8006,N_8046);
and U8154 (N_8154,N_8003,N_8045);
nand U8155 (N_8155,N_8119,N_8089);
nor U8156 (N_8156,N_8109,N_8038);
nor U8157 (N_8157,N_8057,N_8028);
nor U8158 (N_8158,N_8080,N_8100);
or U8159 (N_8159,N_8059,N_8111);
and U8160 (N_8160,N_8099,N_8091);
or U8161 (N_8161,N_8124,N_8023);
or U8162 (N_8162,N_8088,N_8011);
xnor U8163 (N_8163,N_8004,N_8015);
nand U8164 (N_8164,N_8020,N_8002);
and U8165 (N_8165,N_8041,N_8110);
xor U8166 (N_8166,N_8101,N_8092);
nor U8167 (N_8167,N_8009,N_8107);
or U8168 (N_8168,N_8106,N_8040);
and U8169 (N_8169,N_8001,N_8090);
nor U8170 (N_8170,N_8051,N_8120);
and U8171 (N_8171,N_8065,N_8044);
nand U8172 (N_8172,N_8114,N_8016);
xnor U8173 (N_8173,N_8121,N_8025);
nor U8174 (N_8174,N_8029,N_8104);
xor U8175 (N_8175,N_8019,N_8048);
and U8176 (N_8176,N_8116,N_8056);
nor U8177 (N_8177,N_8097,N_8074);
xnor U8178 (N_8178,N_8093,N_8027);
and U8179 (N_8179,N_8021,N_8094);
and U8180 (N_8180,N_8078,N_8115);
xnor U8181 (N_8181,N_8117,N_8095);
or U8182 (N_8182,N_8086,N_8026);
and U8183 (N_8183,N_8118,N_8072);
or U8184 (N_8184,N_8108,N_8098);
or U8185 (N_8185,N_8024,N_8113);
xor U8186 (N_8186,N_8068,N_8031);
or U8187 (N_8187,N_8017,N_8035);
and U8188 (N_8188,N_8010,N_8096);
nor U8189 (N_8189,N_8061,N_8095);
or U8190 (N_8190,N_8084,N_8058);
nand U8191 (N_8191,N_8071,N_8081);
or U8192 (N_8192,N_8111,N_8035);
nor U8193 (N_8193,N_8043,N_8118);
nand U8194 (N_8194,N_8071,N_8015);
nor U8195 (N_8195,N_8081,N_8113);
nand U8196 (N_8196,N_8059,N_8040);
nor U8197 (N_8197,N_8026,N_8011);
and U8198 (N_8198,N_8017,N_8074);
xnor U8199 (N_8199,N_8065,N_8037);
xnor U8200 (N_8200,N_8007,N_8006);
xor U8201 (N_8201,N_8044,N_8064);
nand U8202 (N_8202,N_8086,N_8096);
or U8203 (N_8203,N_8079,N_8032);
or U8204 (N_8204,N_8043,N_8002);
and U8205 (N_8205,N_8018,N_8106);
and U8206 (N_8206,N_8064,N_8120);
nand U8207 (N_8207,N_8113,N_8115);
xnor U8208 (N_8208,N_8075,N_8115);
and U8209 (N_8209,N_8043,N_8033);
and U8210 (N_8210,N_8001,N_8040);
nand U8211 (N_8211,N_8102,N_8082);
xor U8212 (N_8212,N_8080,N_8018);
nand U8213 (N_8213,N_8067,N_8004);
nand U8214 (N_8214,N_8084,N_8099);
nor U8215 (N_8215,N_8105,N_8049);
xor U8216 (N_8216,N_8107,N_8064);
nor U8217 (N_8217,N_8090,N_8015);
nand U8218 (N_8218,N_8000,N_8028);
and U8219 (N_8219,N_8089,N_8067);
nor U8220 (N_8220,N_8004,N_8039);
and U8221 (N_8221,N_8107,N_8014);
and U8222 (N_8222,N_8095,N_8100);
or U8223 (N_8223,N_8110,N_8084);
or U8224 (N_8224,N_8010,N_8093);
nor U8225 (N_8225,N_8045,N_8116);
nor U8226 (N_8226,N_8063,N_8016);
xnor U8227 (N_8227,N_8112,N_8069);
or U8228 (N_8228,N_8021,N_8082);
xor U8229 (N_8229,N_8041,N_8108);
or U8230 (N_8230,N_8016,N_8044);
or U8231 (N_8231,N_8044,N_8120);
or U8232 (N_8232,N_8122,N_8027);
and U8233 (N_8233,N_8120,N_8066);
nor U8234 (N_8234,N_8078,N_8057);
nand U8235 (N_8235,N_8053,N_8011);
nor U8236 (N_8236,N_8048,N_8013);
or U8237 (N_8237,N_8085,N_8084);
xor U8238 (N_8238,N_8081,N_8062);
nand U8239 (N_8239,N_8044,N_8077);
xor U8240 (N_8240,N_8016,N_8052);
nor U8241 (N_8241,N_8113,N_8058);
xor U8242 (N_8242,N_8041,N_8005);
nor U8243 (N_8243,N_8057,N_8041);
and U8244 (N_8244,N_8099,N_8117);
nand U8245 (N_8245,N_8029,N_8033);
or U8246 (N_8246,N_8109,N_8093);
and U8247 (N_8247,N_8080,N_8015);
and U8248 (N_8248,N_8070,N_8029);
nand U8249 (N_8249,N_8116,N_8013);
xor U8250 (N_8250,N_8241,N_8164);
or U8251 (N_8251,N_8180,N_8209);
nor U8252 (N_8252,N_8165,N_8247);
xor U8253 (N_8253,N_8240,N_8244);
nand U8254 (N_8254,N_8188,N_8202);
nor U8255 (N_8255,N_8184,N_8157);
nand U8256 (N_8256,N_8192,N_8217);
nor U8257 (N_8257,N_8204,N_8171);
and U8258 (N_8258,N_8168,N_8178);
and U8259 (N_8259,N_8215,N_8141);
or U8260 (N_8260,N_8183,N_8221);
or U8261 (N_8261,N_8142,N_8144);
and U8262 (N_8262,N_8199,N_8214);
or U8263 (N_8263,N_8216,N_8198);
and U8264 (N_8264,N_8200,N_8159);
or U8265 (N_8265,N_8151,N_8243);
nor U8266 (N_8266,N_8166,N_8155);
nand U8267 (N_8267,N_8158,N_8173);
nor U8268 (N_8268,N_8237,N_8163);
and U8269 (N_8269,N_8189,N_8233);
xnor U8270 (N_8270,N_8125,N_8154);
xor U8271 (N_8271,N_8203,N_8211);
xnor U8272 (N_8272,N_8145,N_8149);
or U8273 (N_8273,N_8210,N_8179);
nor U8274 (N_8274,N_8150,N_8174);
or U8275 (N_8275,N_8246,N_8167);
nor U8276 (N_8276,N_8242,N_8205);
and U8277 (N_8277,N_8162,N_8186);
and U8278 (N_8278,N_8170,N_8130);
or U8279 (N_8279,N_8207,N_8126);
nor U8280 (N_8280,N_8222,N_8236);
nand U8281 (N_8281,N_8187,N_8148);
nor U8282 (N_8282,N_8139,N_8245);
and U8283 (N_8283,N_8127,N_8146);
and U8284 (N_8284,N_8208,N_8143);
nand U8285 (N_8285,N_8128,N_8135);
xor U8286 (N_8286,N_8248,N_8197);
or U8287 (N_8287,N_8206,N_8177);
xnor U8288 (N_8288,N_8239,N_8193);
nand U8289 (N_8289,N_8138,N_8228);
nor U8290 (N_8290,N_8220,N_8156);
xor U8291 (N_8291,N_8194,N_8218);
nor U8292 (N_8292,N_8224,N_8136);
nand U8293 (N_8293,N_8238,N_8196);
or U8294 (N_8294,N_8137,N_8223);
or U8295 (N_8295,N_8235,N_8147);
nand U8296 (N_8296,N_8225,N_8234);
nand U8297 (N_8297,N_8249,N_8229);
or U8298 (N_8298,N_8129,N_8132);
nand U8299 (N_8299,N_8169,N_8175);
nor U8300 (N_8300,N_8140,N_8190);
nand U8301 (N_8301,N_8172,N_8133);
xnor U8302 (N_8302,N_8176,N_8191);
nor U8303 (N_8303,N_8213,N_8182);
nor U8304 (N_8304,N_8152,N_8212);
nand U8305 (N_8305,N_8231,N_8232);
nor U8306 (N_8306,N_8195,N_8227);
nor U8307 (N_8307,N_8185,N_8131);
nor U8308 (N_8308,N_8219,N_8153);
or U8309 (N_8309,N_8181,N_8201);
or U8310 (N_8310,N_8134,N_8230);
and U8311 (N_8311,N_8161,N_8226);
xor U8312 (N_8312,N_8160,N_8138);
xor U8313 (N_8313,N_8144,N_8186);
and U8314 (N_8314,N_8155,N_8152);
nand U8315 (N_8315,N_8230,N_8153);
or U8316 (N_8316,N_8207,N_8183);
and U8317 (N_8317,N_8148,N_8214);
nor U8318 (N_8318,N_8127,N_8226);
nand U8319 (N_8319,N_8171,N_8174);
nor U8320 (N_8320,N_8245,N_8180);
or U8321 (N_8321,N_8146,N_8190);
and U8322 (N_8322,N_8218,N_8142);
xor U8323 (N_8323,N_8147,N_8227);
xnor U8324 (N_8324,N_8133,N_8235);
and U8325 (N_8325,N_8125,N_8163);
or U8326 (N_8326,N_8245,N_8154);
or U8327 (N_8327,N_8133,N_8152);
and U8328 (N_8328,N_8215,N_8222);
xnor U8329 (N_8329,N_8192,N_8173);
xor U8330 (N_8330,N_8224,N_8242);
nor U8331 (N_8331,N_8201,N_8220);
and U8332 (N_8332,N_8226,N_8178);
nand U8333 (N_8333,N_8204,N_8126);
nand U8334 (N_8334,N_8234,N_8242);
xnor U8335 (N_8335,N_8247,N_8167);
and U8336 (N_8336,N_8159,N_8244);
or U8337 (N_8337,N_8234,N_8230);
or U8338 (N_8338,N_8243,N_8155);
nor U8339 (N_8339,N_8193,N_8174);
nand U8340 (N_8340,N_8194,N_8192);
and U8341 (N_8341,N_8171,N_8185);
xor U8342 (N_8342,N_8199,N_8151);
and U8343 (N_8343,N_8129,N_8140);
or U8344 (N_8344,N_8207,N_8129);
and U8345 (N_8345,N_8143,N_8244);
nor U8346 (N_8346,N_8156,N_8172);
and U8347 (N_8347,N_8175,N_8224);
and U8348 (N_8348,N_8186,N_8248);
xor U8349 (N_8349,N_8207,N_8172);
nor U8350 (N_8350,N_8227,N_8205);
nand U8351 (N_8351,N_8166,N_8165);
or U8352 (N_8352,N_8164,N_8196);
xnor U8353 (N_8353,N_8239,N_8204);
nor U8354 (N_8354,N_8248,N_8249);
or U8355 (N_8355,N_8191,N_8164);
nand U8356 (N_8356,N_8146,N_8172);
nand U8357 (N_8357,N_8158,N_8152);
and U8358 (N_8358,N_8218,N_8150);
and U8359 (N_8359,N_8195,N_8196);
or U8360 (N_8360,N_8244,N_8203);
nand U8361 (N_8361,N_8179,N_8154);
nor U8362 (N_8362,N_8148,N_8198);
xnor U8363 (N_8363,N_8218,N_8179);
xnor U8364 (N_8364,N_8126,N_8182);
and U8365 (N_8365,N_8186,N_8154);
nand U8366 (N_8366,N_8189,N_8241);
xor U8367 (N_8367,N_8205,N_8186);
nand U8368 (N_8368,N_8162,N_8164);
and U8369 (N_8369,N_8135,N_8144);
xnor U8370 (N_8370,N_8190,N_8196);
nand U8371 (N_8371,N_8223,N_8236);
nand U8372 (N_8372,N_8187,N_8167);
xor U8373 (N_8373,N_8163,N_8158);
xor U8374 (N_8374,N_8210,N_8191);
and U8375 (N_8375,N_8303,N_8368);
and U8376 (N_8376,N_8262,N_8253);
nand U8377 (N_8377,N_8308,N_8366);
or U8378 (N_8378,N_8250,N_8321);
nand U8379 (N_8379,N_8325,N_8364);
and U8380 (N_8380,N_8302,N_8260);
and U8381 (N_8381,N_8310,N_8272);
xnor U8382 (N_8382,N_8338,N_8255);
nor U8383 (N_8383,N_8354,N_8293);
nand U8384 (N_8384,N_8358,N_8335);
nand U8385 (N_8385,N_8267,N_8345);
xor U8386 (N_8386,N_8276,N_8355);
xor U8387 (N_8387,N_8340,N_8307);
nor U8388 (N_8388,N_8283,N_8264);
xor U8389 (N_8389,N_8373,N_8269);
and U8390 (N_8390,N_8298,N_8339);
xor U8391 (N_8391,N_8282,N_8320);
and U8392 (N_8392,N_8331,N_8311);
nor U8393 (N_8393,N_8319,N_8263);
or U8394 (N_8394,N_8297,N_8299);
nor U8395 (N_8395,N_8281,N_8256);
nand U8396 (N_8396,N_8268,N_8360);
nor U8397 (N_8397,N_8343,N_8369);
xor U8398 (N_8398,N_8254,N_8341);
xnor U8399 (N_8399,N_8295,N_8324);
or U8400 (N_8400,N_8286,N_8344);
xnor U8401 (N_8401,N_8314,N_8291);
xnor U8402 (N_8402,N_8329,N_8367);
xor U8403 (N_8403,N_8348,N_8353);
xor U8404 (N_8404,N_8334,N_8359);
nand U8405 (N_8405,N_8350,N_8328);
or U8406 (N_8406,N_8316,N_8288);
nand U8407 (N_8407,N_8357,N_8361);
nand U8408 (N_8408,N_8278,N_8347);
xnor U8409 (N_8409,N_8300,N_8371);
nor U8410 (N_8410,N_8374,N_8259);
or U8411 (N_8411,N_8289,N_8323);
nand U8412 (N_8412,N_8306,N_8290);
and U8413 (N_8413,N_8279,N_8285);
nand U8414 (N_8414,N_8312,N_8349);
or U8415 (N_8415,N_8273,N_8317);
and U8416 (N_8416,N_8322,N_8275);
and U8417 (N_8417,N_8342,N_8326);
and U8418 (N_8418,N_8270,N_8352);
nor U8419 (N_8419,N_8261,N_8266);
or U8420 (N_8420,N_8287,N_8363);
xor U8421 (N_8421,N_8271,N_8332);
or U8422 (N_8422,N_8274,N_8337);
and U8423 (N_8423,N_8327,N_8258);
and U8424 (N_8424,N_8277,N_8333);
or U8425 (N_8425,N_8304,N_8346);
and U8426 (N_8426,N_8301,N_8309);
and U8427 (N_8427,N_8356,N_8257);
nor U8428 (N_8428,N_8252,N_8296);
and U8429 (N_8429,N_8336,N_8284);
xnor U8430 (N_8430,N_8251,N_8351);
nand U8431 (N_8431,N_8365,N_8294);
and U8432 (N_8432,N_8330,N_8292);
xnor U8433 (N_8433,N_8313,N_8265);
nand U8434 (N_8434,N_8370,N_8305);
nor U8435 (N_8435,N_8318,N_8280);
and U8436 (N_8436,N_8372,N_8362);
or U8437 (N_8437,N_8315,N_8277);
or U8438 (N_8438,N_8267,N_8332);
xnor U8439 (N_8439,N_8268,N_8350);
nand U8440 (N_8440,N_8289,N_8271);
nand U8441 (N_8441,N_8368,N_8345);
nor U8442 (N_8442,N_8327,N_8269);
nand U8443 (N_8443,N_8348,N_8285);
and U8444 (N_8444,N_8259,N_8276);
nand U8445 (N_8445,N_8252,N_8371);
nor U8446 (N_8446,N_8253,N_8374);
nand U8447 (N_8447,N_8332,N_8365);
nor U8448 (N_8448,N_8308,N_8266);
nand U8449 (N_8449,N_8257,N_8310);
and U8450 (N_8450,N_8353,N_8304);
or U8451 (N_8451,N_8324,N_8371);
nor U8452 (N_8452,N_8320,N_8286);
and U8453 (N_8453,N_8296,N_8326);
and U8454 (N_8454,N_8344,N_8367);
xnor U8455 (N_8455,N_8361,N_8262);
and U8456 (N_8456,N_8253,N_8285);
nand U8457 (N_8457,N_8367,N_8270);
xnor U8458 (N_8458,N_8339,N_8356);
nor U8459 (N_8459,N_8340,N_8309);
or U8460 (N_8460,N_8334,N_8362);
or U8461 (N_8461,N_8304,N_8271);
nand U8462 (N_8462,N_8350,N_8262);
xnor U8463 (N_8463,N_8354,N_8256);
xor U8464 (N_8464,N_8282,N_8311);
xnor U8465 (N_8465,N_8286,N_8271);
nor U8466 (N_8466,N_8309,N_8367);
nor U8467 (N_8467,N_8312,N_8290);
nand U8468 (N_8468,N_8355,N_8348);
nor U8469 (N_8469,N_8261,N_8335);
xnor U8470 (N_8470,N_8266,N_8362);
nand U8471 (N_8471,N_8350,N_8332);
and U8472 (N_8472,N_8330,N_8258);
nor U8473 (N_8473,N_8370,N_8252);
nor U8474 (N_8474,N_8298,N_8371);
or U8475 (N_8475,N_8298,N_8350);
xor U8476 (N_8476,N_8252,N_8271);
xnor U8477 (N_8477,N_8345,N_8275);
and U8478 (N_8478,N_8251,N_8305);
and U8479 (N_8479,N_8374,N_8356);
and U8480 (N_8480,N_8373,N_8360);
nand U8481 (N_8481,N_8307,N_8278);
and U8482 (N_8482,N_8253,N_8290);
nor U8483 (N_8483,N_8329,N_8283);
nor U8484 (N_8484,N_8355,N_8320);
nand U8485 (N_8485,N_8304,N_8328);
and U8486 (N_8486,N_8302,N_8308);
and U8487 (N_8487,N_8327,N_8337);
nand U8488 (N_8488,N_8283,N_8364);
xnor U8489 (N_8489,N_8366,N_8328);
and U8490 (N_8490,N_8323,N_8310);
nor U8491 (N_8491,N_8330,N_8338);
and U8492 (N_8492,N_8282,N_8278);
nand U8493 (N_8493,N_8287,N_8353);
or U8494 (N_8494,N_8371,N_8288);
nor U8495 (N_8495,N_8334,N_8253);
xnor U8496 (N_8496,N_8256,N_8263);
or U8497 (N_8497,N_8353,N_8272);
or U8498 (N_8498,N_8303,N_8373);
or U8499 (N_8499,N_8259,N_8318);
xor U8500 (N_8500,N_8491,N_8423);
nor U8501 (N_8501,N_8488,N_8448);
and U8502 (N_8502,N_8389,N_8427);
or U8503 (N_8503,N_8384,N_8402);
nor U8504 (N_8504,N_8405,N_8493);
xor U8505 (N_8505,N_8428,N_8429);
nor U8506 (N_8506,N_8446,N_8407);
xnor U8507 (N_8507,N_8475,N_8441);
or U8508 (N_8508,N_8454,N_8489);
xor U8509 (N_8509,N_8456,N_8485);
nand U8510 (N_8510,N_8430,N_8455);
or U8511 (N_8511,N_8409,N_8464);
nand U8512 (N_8512,N_8497,N_8385);
or U8513 (N_8513,N_8462,N_8473);
nor U8514 (N_8514,N_8471,N_8482);
or U8515 (N_8515,N_8378,N_8387);
nand U8516 (N_8516,N_8474,N_8496);
or U8517 (N_8517,N_8465,N_8444);
and U8518 (N_8518,N_8377,N_8443);
xor U8519 (N_8519,N_8393,N_8418);
nor U8520 (N_8520,N_8492,N_8420);
and U8521 (N_8521,N_8438,N_8381);
xnor U8522 (N_8522,N_8422,N_8419);
or U8523 (N_8523,N_8408,N_8480);
xor U8524 (N_8524,N_8457,N_8458);
nand U8525 (N_8525,N_8451,N_8450);
and U8526 (N_8526,N_8416,N_8404);
nor U8527 (N_8527,N_8417,N_8477);
or U8528 (N_8528,N_8498,N_8388);
nand U8529 (N_8529,N_8452,N_8403);
nor U8530 (N_8530,N_8442,N_8466);
and U8531 (N_8531,N_8432,N_8413);
and U8532 (N_8532,N_8433,N_8470);
and U8533 (N_8533,N_8376,N_8449);
nand U8534 (N_8534,N_8494,N_8399);
nor U8535 (N_8535,N_8412,N_8490);
nand U8536 (N_8536,N_8447,N_8394);
or U8537 (N_8537,N_8406,N_8467);
xnor U8538 (N_8538,N_8440,N_8380);
nand U8539 (N_8539,N_8460,N_8437);
xor U8540 (N_8540,N_8453,N_8375);
xnor U8541 (N_8541,N_8436,N_8495);
nor U8542 (N_8542,N_8469,N_8390);
and U8543 (N_8543,N_8425,N_8411);
and U8544 (N_8544,N_8414,N_8401);
and U8545 (N_8545,N_8479,N_8499);
nor U8546 (N_8546,N_8383,N_8478);
and U8547 (N_8547,N_8382,N_8476);
nor U8548 (N_8548,N_8431,N_8396);
or U8549 (N_8549,N_8410,N_8487);
nand U8550 (N_8550,N_8435,N_8434);
nor U8551 (N_8551,N_8468,N_8424);
xnor U8552 (N_8552,N_8481,N_8439);
nand U8553 (N_8553,N_8459,N_8379);
xnor U8554 (N_8554,N_8415,N_8445);
and U8555 (N_8555,N_8391,N_8461);
nand U8556 (N_8556,N_8392,N_8395);
and U8557 (N_8557,N_8483,N_8426);
nor U8558 (N_8558,N_8398,N_8397);
nor U8559 (N_8559,N_8484,N_8386);
or U8560 (N_8560,N_8472,N_8463);
nand U8561 (N_8561,N_8421,N_8486);
xor U8562 (N_8562,N_8400,N_8380);
nor U8563 (N_8563,N_8491,N_8445);
and U8564 (N_8564,N_8391,N_8469);
xor U8565 (N_8565,N_8399,N_8481);
nand U8566 (N_8566,N_8394,N_8439);
and U8567 (N_8567,N_8487,N_8425);
nor U8568 (N_8568,N_8489,N_8380);
nor U8569 (N_8569,N_8408,N_8464);
or U8570 (N_8570,N_8421,N_8381);
and U8571 (N_8571,N_8499,N_8417);
nor U8572 (N_8572,N_8455,N_8421);
or U8573 (N_8573,N_8482,N_8461);
nor U8574 (N_8574,N_8446,N_8488);
nand U8575 (N_8575,N_8383,N_8434);
and U8576 (N_8576,N_8447,N_8438);
nor U8577 (N_8577,N_8389,N_8480);
nor U8578 (N_8578,N_8404,N_8491);
and U8579 (N_8579,N_8436,N_8399);
xnor U8580 (N_8580,N_8468,N_8432);
and U8581 (N_8581,N_8443,N_8461);
nand U8582 (N_8582,N_8486,N_8380);
xor U8583 (N_8583,N_8487,N_8432);
xor U8584 (N_8584,N_8477,N_8461);
or U8585 (N_8585,N_8404,N_8493);
nand U8586 (N_8586,N_8379,N_8498);
nand U8587 (N_8587,N_8423,N_8380);
or U8588 (N_8588,N_8376,N_8442);
xor U8589 (N_8589,N_8389,N_8474);
nor U8590 (N_8590,N_8455,N_8486);
nor U8591 (N_8591,N_8497,N_8395);
xnor U8592 (N_8592,N_8499,N_8465);
xnor U8593 (N_8593,N_8445,N_8447);
nor U8594 (N_8594,N_8414,N_8423);
xor U8595 (N_8595,N_8433,N_8375);
nand U8596 (N_8596,N_8383,N_8469);
or U8597 (N_8597,N_8408,N_8469);
nor U8598 (N_8598,N_8427,N_8444);
or U8599 (N_8599,N_8428,N_8437);
or U8600 (N_8600,N_8380,N_8448);
or U8601 (N_8601,N_8415,N_8431);
xnor U8602 (N_8602,N_8377,N_8388);
nor U8603 (N_8603,N_8412,N_8485);
xnor U8604 (N_8604,N_8440,N_8461);
xnor U8605 (N_8605,N_8405,N_8447);
nand U8606 (N_8606,N_8478,N_8467);
nor U8607 (N_8607,N_8477,N_8377);
nand U8608 (N_8608,N_8456,N_8467);
nor U8609 (N_8609,N_8408,N_8454);
nor U8610 (N_8610,N_8462,N_8469);
and U8611 (N_8611,N_8384,N_8439);
nor U8612 (N_8612,N_8385,N_8484);
and U8613 (N_8613,N_8375,N_8440);
nand U8614 (N_8614,N_8402,N_8466);
or U8615 (N_8615,N_8375,N_8481);
xnor U8616 (N_8616,N_8465,N_8459);
nor U8617 (N_8617,N_8430,N_8487);
or U8618 (N_8618,N_8399,N_8477);
or U8619 (N_8619,N_8433,N_8493);
xor U8620 (N_8620,N_8440,N_8474);
nand U8621 (N_8621,N_8399,N_8471);
nand U8622 (N_8622,N_8462,N_8400);
and U8623 (N_8623,N_8433,N_8476);
or U8624 (N_8624,N_8401,N_8420);
and U8625 (N_8625,N_8556,N_8604);
nor U8626 (N_8626,N_8512,N_8609);
nor U8627 (N_8627,N_8583,N_8564);
and U8628 (N_8628,N_8503,N_8562);
and U8629 (N_8629,N_8593,N_8552);
or U8630 (N_8630,N_8601,N_8605);
or U8631 (N_8631,N_8585,N_8561);
nand U8632 (N_8632,N_8570,N_8567);
nor U8633 (N_8633,N_8619,N_8530);
nand U8634 (N_8634,N_8571,N_8534);
and U8635 (N_8635,N_8525,N_8578);
nor U8636 (N_8636,N_8584,N_8524);
or U8637 (N_8637,N_8518,N_8513);
nor U8638 (N_8638,N_8608,N_8523);
xnor U8639 (N_8639,N_8577,N_8529);
or U8640 (N_8640,N_8536,N_8526);
xnor U8641 (N_8641,N_8540,N_8614);
or U8642 (N_8642,N_8545,N_8528);
xnor U8643 (N_8643,N_8595,N_8527);
or U8644 (N_8644,N_8617,N_8542);
or U8645 (N_8645,N_8533,N_8610);
nand U8646 (N_8646,N_8566,N_8511);
nand U8647 (N_8647,N_8517,N_8613);
or U8648 (N_8648,N_8618,N_8569);
and U8649 (N_8649,N_8506,N_8600);
and U8650 (N_8650,N_8621,N_8507);
and U8651 (N_8651,N_8549,N_8514);
nor U8652 (N_8652,N_8521,N_8568);
and U8653 (N_8653,N_8612,N_8502);
nor U8654 (N_8654,N_8535,N_8504);
xor U8655 (N_8655,N_8501,N_8592);
nand U8656 (N_8656,N_8599,N_8563);
and U8657 (N_8657,N_8576,N_8510);
or U8658 (N_8658,N_8532,N_8550);
nand U8659 (N_8659,N_8546,N_8622);
nor U8660 (N_8660,N_8505,N_8522);
nor U8661 (N_8661,N_8580,N_8581);
or U8662 (N_8662,N_8586,N_8603);
xnor U8663 (N_8663,N_8565,N_8531);
or U8664 (N_8664,N_8520,N_8596);
or U8665 (N_8665,N_8559,N_8615);
nand U8666 (N_8666,N_8572,N_8539);
and U8667 (N_8667,N_8537,N_8590);
nor U8668 (N_8668,N_8547,N_8508);
or U8669 (N_8669,N_8611,N_8544);
or U8670 (N_8670,N_8554,N_8519);
xor U8671 (N_8671,N_8548,N_8543);
xnor U8672 (N_8672,N_8555,N_8516);
nor U8673 (N_8673,N_8573,N_8538);
nor U8674 (N_8674,N_8551,N_8598);
nor U8675 (N_8675,N_8594,N_8623);
nand U8676 (N_8676,N_8541,N_8553);
and U8677 (N_8677,N_8616,N_8560);
xor U8678 (N_8678,N_8620,N_8557);
nor U8679 (N_8679,N_8624,N_8602);
nor U8680 (N_8680,N_8589,N_8587);
or U8681 (N_8681,N_8582,N_8515);
and U8682 (N_8682,N_8575,N_8597);
nand U8683 (N_8683,N_8558,N_8606);
xor U8684 (N_8684,N_8579,N_8574);
or U8685 (N_8685,N_8500,N_8607);
nor U8686 (N_8686,N_8588,N_8509);
nor U8687 (N_8687,N_8591,N_8578);
nand U8688 (N_8688,N_8501,N_8566);
nor U8689 (N_8689,N_8500,N_8531);
or U8690 (N_8690,N_8538,N_8598);
and U8691 (N_8691,N_8562,N_8500);
nand U8692 (N_8692,N_8580,N_8623);
nor U8693 (N_8693,N_8562,N_8521);
or U8694 (N_8694,N_8568,N_8611);
nor U8695 (N_8695,N_8614,N_8537);
nor U8696 (N_8696,N_8590,N_8572);
nand U8697 (N_8697,N_8614,N_8577);
and U8698 (N_8698,N_8517,N_8530);
nand U8699 (N_8699,N_8500,N_8555);
nand U8700 (N_8700,N_8616,N_8601);
nor U8701 (N_8701,N_8514,N_8609);
nor U8702 (N_8702,N_8536,N_8586);
and U8703 (N_8703,N_8552,N_8577);
or U8704 (N_8704,N_8507,N_8550);
or U8705 (N_8705,N_8505,N_8588);
nand U8706 (N_8706,N_8526,N_8621);
nor U8707 (N_8707,N_8606,N_8514);
nor U8708 (N_8708,N_8527,N_8553);
xnor U8709 (N_8709,N_8506,N_8605);
xor U8710 (N_8710,N_8575,N_8525);
nand U8711 (N_8711,N_8504,N_8546);
and U8712 (N_8712,N_8568,N_8572);
xnor U8713 (N_8713,N_8566,N_8528);
nor U8714 (N_8714,N_8615,N_8566);
or U8715 (N_8715,N_8507,N_8542);
nand U8716 (N_8716,N_8546,N_8500);
or U8717 (N_8717,N_8606,N_8620);
xnor U8718 (N_8718,N_8517,N_8574);
nor U8719 (N_8719,N_8532,N_8577);
nor U8720 (N_8720,N_8606,N_8607);
nand U8721 (N_8721,N_8554,N_8579);
and U8722 (N_8722,N_8591,N_8501);
nand U8723 (N_8723,N_8554,N_8592);
xor U8724 (N_8724,N_8600,N_8540);
nand U8725 (N_8725,N_8605,N_8519);
and U8726 (N_8726,N_8591,N_8547);
or U8727 (N_8727,N_8621,N_8584);
nand U8728 (N_8728,N_8539,N_8569);
xor U8729 (N_8729,N_8538,N_8531);
nand U8730 (N_8730,N_8619,N_8584);
nand U8731 (N_8731,N_8589,N_8582);
or U8732 (N_8732,N_8501,N_8542);
or U8733 (N_8733,N_8504,N_8548);
xor U8734 (N_8734,N_8554,N_8606);
and U8735 (N_8735,N_8532,N_8538);
and U8736 (N_8736,N_8574,N_8605);
xnor U8737 (N_8737,N_8579,N_8565);
or U8738 (N_8738,N_8508,N_8560);
nand U8739 (N_8739,N_8520,N_8576);
nor U8740 (N_8740,N_8595,N_8563);
nor U8741 (N_8741,N_8518,N_8622);
nand U8742 (N_8742,N_8595,N_8558);
or U8743 (N_8743,N_8600,N_8580);
xor U8744 (N_8744,N_8591,N_8521);
nor U8745 (N_8745,N_8594,N_8559);
nand U8746 (N_8746,N_8505,N_8575);
nor U8747 (N_8747,N_8570,N_8500);
or U8748 (N_8748,N_8582,N_8592);
and U8749 (N_8749,N_8589,N_8584);
nand U8750 (N_8750,N_8684,N_8648);
or U8751 (N_8751,N_8719,N_8663);
xnor U8752 (N_8752,N_8729,N_8697);
and U8753 (N_8753,N_8634,N_8686);
or U8754 (N_8754,N_8734,N_8642);
xnor U8755 (N_8755,N_8645,N_8651);
and U8756 (N_8756,N_8725,N_8733);
nand U8757 (N_8757,N_8741,N_8673);
nand U8758 (N_8758,N_8636,N_8660);
and U8759 (N_8759,N_8744,N_8694);
or U8760 (N_8760,N_8666,N_8655);
nand U8761 (N_8761,N_8637,N_8742);
nor U8762 (N_8762,N_8676,N_8625);
nor U8763 (N_8763,N_8709,N_8708);
nor U8764 (N_8764,N_8702,N_8714);
and U8765 (N_8765,N_8720,N_8746);
nor U8766 (N_8766,N_8704,N_8703);
nor U8767 (N_8767,N_8639,N_8681);
nor U8768 (N_8768,N_8728,N_8679);
nand U8769 (N_8769,N_8653,N_8726);
nor U8770 (N_8770,N_8747,N_8727);
xnor U8771 (N_8771,N_8627,N_8721);
or U8772 (N_8772,N_8659,N_8696);
or U8773 (N_8773,N_8672,N_8692);
nor U8774 (N_8774,N_8730,N_8633);
nor U8775 (N_8775,N_8713,N_8695);
or U8776 (N_8776,N_8678,N_8712);
or U8777 (N_8777,N_8738,N_8656);
nand U8778 (N_8778,N_8683,N_8724);
nand U8779 (N_8779,N_8677,N_8665);
xor U8780 (N_8780,N_8739,N_8675);
nand U8781 (N_8781,N_8687,N_8740);
or U8782 (N_8782,N_8630,N_8710);
nand U8783 (N_8783,N_8640,N_8646);
or U8784 (N_8784,N_8638,N_8669);
or U8785 (N_8785,N_8718,N_8705);
nand U8786 (N_8786,N_8690,N_8715);
nand U8787 (N_8787,N_8654,N_8682);
and U8788 (N_8788,N_8658,N_8731);
nor U8789 (N_8789,N_8628,N_8700);
or U8790 (N_8790,N_8674,N_8661);
or U8791 (N_8791,N_8650,N_8717);
nand U8792 (N_8792,N_8711,N_8699);
nand U8793 (N_8793,N_8641,N_8671);
nand U8794 (N_8794,N_8668,N_8743);
or U8795 (N_8795,N_8647,N_8749);
nand U8796 (N_8796,N_8685,N_8664);
nand U8797 (N_8797,N_8632,N_8631);
nand U8798 (N_8798,N_8670,N_8667);
xnor U8799 (N_8799,N_8688,N_8644);
and U8800 (N_8800,N_8635,N_8689);
or U8801 (N_8801,N_8662,N_8716);
xnor U8802 (N_8802,N_8745,N_8706);
or U8803 (N_8803,N_8701,N_8698);
nor U8804 (N_8804,N_8629,N_8657);
nand U8805 (N_8805,N_8652,N_8722);
nor U8806 (N_8806,N_8748,N_8732);
nand U8807 (N_8807,N_8649,N_8736);
or U8808 (N_8808,N_8707,N_8680);
nor U8809 (N_8809,N_8737,N_8626);
or U8810 (N_8810,N_8643,N_8723);
and U8811 (N_8811,N_8693,N_8735);
nand U8812 (N_8812,N_8691,N_8707);
or U8813 (N_8813,N_8749,N_8687);
and U8814 (N_8814,N_8692,N_8669);
or U8815 (N_8815,N_8676,N_8672);
and U8816 (N_8816,N_8677,N_8682);
xnor U8817 (N_8817,N_8740,N_8656);
or U8818 (N_8818,N_8667,N_8738);
nor U8819 (N_8819,N_8733,N_8650);
nor U8820 (N_8820,N_8648,N_8724);
nand U8821 (N_8821,N_8694,N_8714);
xor U8822 (N_8822,N_8626,N_8724);
nand U8823 (N_8823,N_8716,N_8727);
or U8824 (N_8824,N_8681,N_8645);
and U8825 (N_8825,N_8745,N_8648);
or U8826 (N_8826,N_8723,N_8674);
nand U8827 (N_8827,N_8684,N_8732);
nand U8828 (N_8828,N_8721,N_8671);
or U8829 (N_8829,N_8693,N_8642);
nor U8830 (N_8830,N_8742,N_8625);
xor U8831 (N_8831,N_8687,N_8685);
and U8832 (N_8832,N_8745,N_8723);
xnor U8833 (N_8833,N_8734,N_8683);
or U8834 (N_8834,N_8680,N_8648);
or U8835 (N_8835,N_8709,N_8691);
and U8836 (N_8836,N_8700,N_8629);
nor U8837 (N_8837,N_8703,N_8732);
xnor U8838 (N_8838,N_8659,N_8677);
and U8839 (N_8839,N_8671,N_8729);
xor U8840 (N_8840,N_8646,N_8729);
nand U8841 (N_8841,N_8714,N_8718);
or U8842 (N_8842,N_8636,N_8686);
and U8843 (N_8843,N_8732,N_8723);
nand U8844 (N_8844,N_8662,N_8651);
or U8845 (N_8845,N_8710,N_8691);
xnor U8846 (N_8846,N_8639,N_8748);
nand U8847 (N_8847,N_8704,N_8694);
nor U8848 (N_8848,N_8658,N_8661);
and U8849 (N_8849,N_8747,N_8655);
or U8850 (N_8850,N_8720,N_8654);
and U8851 (N_8851,N_8641,N_8698);
xor U8852 (N_8852,N_8667,N_8737);
nor U8853 (N_8853,N_8720,N_8679);
nor U8854 (N_8854,N_8706,N_8657);
or U8855 (N_8855,N_8725,N_8729);
and U8856 (N_8856,N_8723,N_8630);
xnor U8857 (N_8857,N_8744,N_8678);
or U8858 (N_8858,N_8694,N_8728);
nor U8859 (N_8859,N_8734,N_8633);
or U8860 (N_8860,N_8741,N_8747);
and U8861 (N_8861,N_8744,N_8723);
or U8862 (N_8862,N_8725,N_8678);
xnor U8863 (N_8863,N_8690,N_8705);
nor U8864 (N_8864,N_8682,N_8717);
and U8865 (N_8865,N_8705,N_8749);
or U8866 (N_8866,N_8661,N_8709);
nand U8867 (N_8867,N_8701,N_8674);
xor U8868 (N_8868,N_8678,N_8733);
nor U8869 (N_8869,N_8642,N_8727);
nor U8870 (N_8870,N_8694,N_8718);
xor U8871 (N_8871,N_8738,N_8728);
and U8872 (N_8872,N_8631,N_8670);
nand U8873 (N_8873,N_8683,N_8670);
or U8874 (N_8874,N_8678,N_8641);
and U8875 (N_8875,N_8867,N_8794);
nor U8876 (N_8876,N_8774,N_8815);
or U8877 (N_8877,N_8809,N_8769);
xor U8878 (N_8878,N_8776,N_8833);
nand U8879 (N_8879,N_8840,N_8831);
xor U8880 (N_8880,N_8786,N_8810);
nand U8881 (N_8881,N_8872,N_8773);
nor U8882 (N_8882,N_8799,N_8797);
or U8883 (N_8883,N_8821,N_8830);
or U8884 (N_8884,N_8814,N_8808);
nand U8885 (N_8885,N_8853,N_8858);
nand U8886 (N_8886,N_8762,N_8804);
and U8887 (N_8887,N_8826,N_8857);
and U8888 (N_8888,N_8846,N_8855);
nor U8889 (N_8889,N_8870,N_8750);
nand U8890 (N_8890,N_8819,N_8865);
or U8891 (N_8891,N_8861,N_8752);
nor U8892 (N_8892,N_8869,N_8784);
nand U8893 (N_8893,N_8841,N_8850);
nor U8894 (N_8894,N_8780,N_8759);
nand U8895 (N_8895,N_8866,N_8798);
nor U8896 (N_8896,N_8766,N_8771);
xnor U8897 (N_8897,N_8832,N_8851);
and U8898 (N_8898,N_8756,N_8755);
or U8899 (N_8899,N_8765,N_8806);
xnor U8900 (N_8900,N_8775,N_8795);
or U8901 (N_8901,N_8767,N_8778);
nand U8902 (N_8902,N_8849,N_8801);
and U8903 (N_8903,N_8844,N_8847);
nor U8904 (N_8904,N_8789,N_8817);
or U8905 (N_8905,N_8864,N_8845);
xor U8906 (N_8906,N_8757,N_8816);
xnor U8907 (N_8907,N_8790,N_8803);
nor U8908 (N_8908,N_8785,N_8793);
or U8909 (N_8909,N_8760,N_8852);
nor U8910 (N_8910,N_8779,N_8818);
nor U8911 (N_8911,N_8802,N_8812);
and U8912 (N_8912,N_8859,N_8813);
or U8913 (N_8913,N_8764,N_8863);
nor U8914 (N_8914,N_8837,N_8824);
and U8915 (N_8915,N_8770,N_8782);
or U8916 (N_8916,N_8868,N_8874);
nand U8917 (N_8917,N_8828,N_8761);
and U8918 (N_8918,N_8796,N_8842);
and U8919 (N_8919,N_8783,N_8777);
or U8920 (N_8920,N_8836,N_8811);
nor U8921 (N_8921,N_8805,N_8827);
nand U8922 (N_8922,N_8751,N_8820);
nand U8923 (N_8923,N_8838,N_8854);
xnor U8924 (N_8924,N_8825,N_8848);
or U8925 (N_8925,N_8871,N_8791);
and U8926 (N_8926,N_8788,N_8763);
xnor U8927 (N_8927,N_8839,N_8792);
nor U8928 (N_8928,N_8843,N_8787);
nand U8929 (N_8929,N_8753,N_8829);
and U8930 (N_8930,N_8823,N_8860);
xnor U8931 (N_8931,N_8856,N_8768);
or U8932 (N_8932,N_8835,N_8800);
or U8933 (N_8933,N_8834,N_8758);
and U8934 (N_8934,N_8807,N_8772);
or U8935 (N_8935,N_8862,N_8781);
and U8936 (N_8936,N_8822,N_8873);
or U8937 (N_8937,N_8754,N_8765);
and U8938 (N_8938,N_8871,N_8835);
and U8939 (N_8939,N_8806,N_8762);
or U8940 (N_8940,N_8813,N_8764);
xnor U8941 (N_8941,N_8804,N_8842);
nand U8942 (N_8942,N_8866,N_8836);
and U8943 (N_8943,N_8811,N_8833);
nand U8944 (N_8944,N_8759,N_8812);
or U8945 (N_8945,N_8811,N_8860);
or U8946 (N_8946,N_8835,N_8750);
or U8947 (N_8947,N_8847,N_8865);
nand U8948 (N_8948,N_8850,N_8845);
nor U8949 (N_8949,N_8764,N_8770);
and U8950 (N_8950,N_8828,N_8835);
nand U8951 (N_8951,N_8766,N_8824);
or U8952 (N_8952,N_8855,N_8807);
nor U8953 (N_8953,N_8873,N_8797);
xnor U8954 (N_8954,N_8773,N_8751);
nand U8955 (N_8955,N_8772,N_8760);
or U8956 (N_8956,N_8866,N_8761);
or U8957 (N_8957,N_8754,N_8864);
and U8958 (N_8958,N_8830,N_8862);
or U8959 (N_8959,N_8798,N_8870);
xnor U8960 (N_8960,N_8826,N_8801);
and U8961 (N_8961,N_8782,N_8864);
xor U8962 (N_8962,N_8768,N_8824);
nor U8963 (N_8963,N_8854,N_8815);
xor U8964 (N_8964,N_8803,N_8807);
and U8965 (N_8965,N_8870,N_8857);
and U8966 (N_8966,N_8794,N_8828);
xnor U8967 (N_8967,N_8784,N_8834);
or U8968 (N_8968,N_8818,N_8777);
and U8969 (N_8969,N_8820,N_8809);
nor U8970 (N_8970,N_8791,N_8849);
xnor U8971 (N_8971,N_8764,N_8838);
nand U8972 (N_8972,N_8824,N_8786);
xnor U8973 (N_8973,N_8834,N_8768);
xnor U8974 (N_8974,N_8806,N_8816);
nand U8975 (N_8975,N_8829,N_8785);
or U8976 (N_8976,N_8782,N_8819);
and U8977 (N_8977,N_8785,N_8774);
or U8978 (N_8978,N_8766,N_8813);
nand U8979 (N_8979,N_8772,N_8770);
and U8980 (N_8980,N_8838,N_8835);
and U8981 (N_8981,N_8755,N_8763);
xnor U8982 (N_8982,N_8820,N_8867);
nor U8983 (N_8983,N_8828,N_8861);
and U8984 (N_8984,N_8818,N_8833);
nand U8985 (N_8985,N_8788,N_8757);
xnor U8986 (N_8986,N_8781,N_8825);
nand U8987 (N_8987,N_8829,N_8861);
xor U8988 (N_8988,N_8784,N_8871);
xor U8989 (N_8989,N_8811,N_8855);
and U8990 (N_8990,N_8866,N_8769);
nand U8991 (N_8991,N_8843,N_8837);
nor U8992 (N_8992,N_8794,N_8793);
xnor U8993 (N_8993,N_8832,N_8775);
nand U8994 (N_8994,N_8850,N_8873);
nand U8995 (N_8995,N_8824,N_8753);
and U8996 (N_8996,N_8798,N_8839);
or U8997 (N_8997,N_8754,N_8796);
or U8998 (N_8998,N_8767,N_8771);
or U8999 (N_8999,N_8779,N_8820);
nor U9000 (N_9000,N_8927,N_8979);
nor U9001 (N_9001,N_8904,N_8992);
nor U9002 (N_9002,N_8994,N_8991);
nand U9003 (N_9003,N_8993,N_8950);
nand U9004 (N_9004,N_8980,N_8989);
or U9005 (N_9005,N_8940,N_8912);
or U9006 (N_9006,N_8899,N_8881);
nand U9007 (N_9007,N_8971,N_8883);
xor U9008 (N_9008,N_8944,N_8970);
and U9009 (N_9009,N_8875,N_8923);
or U9010 (N_9010,N_8907,N_8965);
and U9011 (N_9011,N_8901,N_8924);
or U9012 (N_9012,N_8946,N_8922);
and U9013 (N_9013,N_8954,N_8930);
nor U9014 (N_9014,N_8948,N_8910);
or U9015 (N_9015,N_8882,N_8937);
and U9016 (N_9016,N_8920,N_8945);
and U9017 (N_9017,N_8889,N_8938);
nor U9018 (N_9018,N_8895,N_8933);
xor U9019 (N_9019,N_8961,N_8952);
nand U9020 (N_9020,N_8995,N_8963);
nand U9021 (N_9021,N_8880,N_8984);
or U9022 (N_9022,N_8981,N_8960);
or U9023 (N_9023,N_8934,N_8947);
nand U9024 (N_9024,N_8997,N_8884);
nand U9025 (N_9025,N_8915,N_8998);
or U9026 (N_9026,N_8982,N_8879);
nand U9027 (N_9027,N_8898,N_8969);
nand U9028 (N_9028,N_8962,N_8917);
xor U9029 (N_9029,N_8908,N_8986);
nand U9030 (N_9030,N_8976,N_8918);
and U9031 (N_9031,N_8876,N_8941);
and U9032 (N_9032,N_8968,N_8888);
and U9033 (N_9033,N_8921,N_8951);
xor U9034 (N_9034,N_8975,N_8974);
nand U9035 (N_9035,N_8914,N_8977);
nand U9036 (N_9036,N_8978,N_8972);
nor U9037 (N_9037,N_8990,N_8919);
nand U9038 (N_9038,N_8949,N_8905);
xor U9039 (N_9039,N_8999,N_8939);
nand U9040 (N_9040,N_8892,N_8886);
xor U9041 (N_9041,N_8957,N_8877);
and U9042 (N_9042,N_8973,N_8959);
nand U9043 (N_9043,N_8903,N_8878);
xnor U9044 (N_9044,N_8983,N_8958);
nor U9045 (N_9045,N_8955,N_8891);
nor U9046 (N_9046,N_8928,N_8967);
and U9047 (N_9047,N_8896,N_8931);
or U9048 (N_9048,N_8911,N_8929);
nor U9049 (N_9049,N_8887,N_8964);
or U9050 (N_9050,N_8909,N_8890);
nor U9051 (N_9051,N_8996,N_8897);
and U9052 (N_9052,N_8902,N_8985);
xor U9053 (N_9053,N_8943,N_8966);
and U9054 (N_9054,N_8935,N_8893);
or U9055 (N_9055,N_8906,N_8953);
and U9056 (N_9056,N_8885,N_8900);
or U9057 (N_9057,N_8987,N_8926);
nor U9058 (N_9058,N_8894,N_8936);
nor U9059 (N_9059,N_8916,N_8956);
and U9060 (N_9060,N_8932,N_8913);
nor U9061 (N_9061,N_8942,N_8925);
and U9062 (N_9062,N_8988,N_8914);
and U9063 (N_9063,N_8916,N_8954);
xnor U9064 (N_9064,N_8917,N_8978);
and U9065 (N_9065,N_8987,N_8901);
and U9066 (N_9066,N_8989,N_8885);
or U9067 (N_9067,N_8913,N_8918);
xnor U9068 (N_9068,N_8995,N_8974);
nand U9069 (N_9069,N_8951,N_8911);
and U9070 (N_9070,N_8997,N_8948);
nor U9071 (N_9071,N_8985,N_8998);
and U9072 (N_9072,N_8892,N_8958);
nor U9073 (N_9073,N_8950,N_8933);
and U9074 (N_9074,N_8914,N_8932);
or U9075 (N_9075,N_8979,N_8924);
nor U9076 (N_9076,N_8936,N_8988);
and U9077 (N_9077,N_8928,N_8917);
nor U9078 (N_9078,N_8987,N_8978);
nand U9079 (N_9079,N_8939,N_8974);
nor U9080 (N_9080,N_8890,N_8938);
or U9081 (N_9081,N_8997,N_8931);
nand U9082 (N_9082,N_8890,N_8931);
nand U9083 (N_9083,N_8925,N_8999);
or U9084 (N_9084,N_8991,N_8928);
nor U9085 (N_9085,N_8984,N_8977);
or U9086 (N_9086,N_8943,N_8985);
xor U9087 (N_9087,N_8986,N_8996);
and U9088 (N_9088,N_8977,N_8974);
nor U9089 (N_9089,N_8885,N_8955);
or U9090 (N_9090,N_8926,N_8946);
nor U9091 (N_9091,N_8959,N_8943);
nor U9092 (N_9092,N_8966,N_8922);
or U9093 (N_9093,N_8912,N_8896);
xnor U9094 (N_9094,N_8955,N_8903);
and U9095 (N_9095,N_8938,N_8998);
nor U9096 (N_9096,N_8889,N_8964);
and U9097 (N_9097,N_8891,N_8900);
or U9098 (N_9098,N_8958,N_8969);
nand U9099 (N_9099,N_8996,N_8904);
and U9100 (N_9100,N_8911,N_8918);
or U9101 (N_9101,N_8922,N_8937);
nand U9102 (N_9102,N_8948,N_8968);
nand U9103 (N_9103,N_8973,N_8902);
xor U9104 (N_9104,N_8962,N_8880);
nand U9105 (N_9105,N_8995,N_8897);
xor U9106 (N_9106,N_8993,N_8990);
nand U9107 (N_9107,N_8904,N_8910);
or U9108 (N_9108,N_8917,N_8911);
xor U9109 (N_9109,N_8946,N_8962);
or U9110 (N_9110,N_8897,N_8896);
and U9111 (N_9111,N_8878,N_8994);
xor U9112 (N_9112,N_8908,N_8937);
or U9113 (N_9113,N_8977,N_8994);
nand U9114 (N_9114,N_8993,N_8983);
xor U9115 (N_9115,N_8950,N_8940);
or U9116 (N_9116,N_8908,N_8901);
nand U9117 (N_9117,N_8885,N_8912);
xor U9118 (N_9118,N_8886,N_8924);
nor U9119 (N_9119,N_8999,N_8901);
nor U9120 (N_9120,N_8918,N_8892);
nand U9121 (N_9121,N_8963,N_8931);
nand U9122 (N_9122,N_8951,N_8903);
and U9123 (N_9123,N_8980,N_8978);
nor U9124 (N_9124,N_8963,N_8891);
or U9125 (N_9125,N_9011,N_9100);
or U9126 (N_9126,N_9005,N_9081);
nor U9127 (N_9127,N_9123,N_9001);
and U9128 (N_9128,N_9003,N_9104);
and U9129 (N_9129,N_9042,N_9102);
or U9130 (N_9130,N_9087,N_9085);
and U9131 (N_9131,N_9002,N_9113);
nor U9132 (N_9132,N_9067,N_9022);
nor U9133 (N_9133,N_9059,N_9040);
and U9134 (N_9134,N_9064,N_9082);
xnor U9135 (N_9135,N_9009,N_9036);
or U9136 (N_9136,N_9027,N_9025);
and U9137 (N_9137,N_9074,N_9073);
and U9138 (N_9138,N_9086,N_9026);
nand U9139 (N_9139,N_9077,N_9056);
and U9140 (N_9140,N_9109,N_9076);
nor U9141 (N_9141,N_9120,N_9045);
or U9142 (N_9142,N_9084,N_9112);
and U9143 (N_9143,N_9016,N_9018);
xnor U9144 (N_9144,N_9024,N_9008);
xor U9145 (N_9145,N_9110,N_9108);
nor U9146 (N_9146,N_9058,N_9019);
and U9147 (N_9147,N_9121,N_9078);
or U9148 (N_9148,N_9052,N_9043);
xnor U9149 (N_9149,N_9017,N_9096);
and U9150 (N_9150,N_9049,N_9031);
xor U9151 (N_9151,N_9035,N_9046);
and U9152 (N_9152,N_9028,N_9079);
xnor U9153 (N_9153,N_9010,N_9083);
nor U9154 (N_9154,N_9041,N_9101);
and U9155 (N_9155,N_9038,N_9103);
nand U9156 (N_9156,N_9091,N_9111);
xnor U9157 (N_9157,N_9007,N_9044);
or U9158 (N_9158,N_9090,N_9061);
xnor U9159 (N_9159,N_9054,N_9032);
or U9160 (N_9160,N_9106,N_9047);
nand U9161 (N_9161,N_9115,N_9029);
nor U9162 (N_9162,N_9000,N_9066);
nand U9163 (N_9163,N_9039,N_9097);
and U9164 (N_9164,N_9094,N_9053);
or U9165 (N_9165,N_9030,N_9093);
or U9166 (N_9166,N_9013,N_9034);
xor U9167 (N_9167,N_9080,N_9089);
xor U9168 (N_9168,N_9057,N_9105);
nor U9169 (N_9169,N_9055,N_9069);
nor U9170 (N_9170,N_9060,N_9114);
nor U9171 (N_9171,N_9122,N_9098);
and U9172 (N_9172,N_9065,N_9014);
nand U9173 (N_9173,N_9068,N_9050);
nor U9174 (N_9174,N_9088,N_9118);
or U9175 (N_9175,N_9124,N_9006);
nand U9176 (N_9176,N_9051,N_9092);
or U9177 (N_9177,N_9037,N_9020);
or U9178 (N_9178,N_9071,N_9004);
or U9179 (N_9179,N_9072,N_9116);
and U9180 (N_9180,N_9099,N_9119);
or U9181 (N_9181,N_9107,N_9062);
nand U9182 (N_9182,N_9117,N_9023);
xnor U9183 (N_9183,N_9012,N_9063);
xor U9184 (N_9184,N_9015,N_9048);
and U9185 (N_9185,N_9095,N_9033);
nand U9186 (N_9186,N_9021,N_9075);
and U9187 (N_9187,N_9070,N_9039);
xnor U9188 (N_9188,N_9040,N_9005);
xnor U9189 (N_9189,N_9121,N_9116);
nand U9190 (N_9190,N_9114,N_9002);
nand U9191 (N_9191,N_9025,N_9113);
xor U9192 (N_9192,N_9004,N_9085);
or U9193 (N_9193,N_9084,N_9074);
nor U9194 (N_9194,N_9053,N_9122);
xnor U9195 (N_9195,N_9114,N_9067);
and U9196 (N_9196,N_9035,N_9097);
xor U9197 (N_9197,N_9032,N_9068);
or U9198 (N_9198,N_9090,N_9079);
xnor U9199 (N_9199,N_9067,N_9110);
nand U9200 (N_9200,N_9103,N_9088);
or U9201 (N_9201,N_9006,N_9024);
nand U9202 (N_9202,N_9045,N_9098);
xor U9203 (N_9203,N_9087,N_9003);
xor U9204 (N_9204,N_9007,N_9101);
nand U9205 (N_9205,N_9063,N_9002);
and U9206 (N_9206,N_9048,N_9032);
nand U9207 (N_9207,N_9000,N_9057);
or U9208 (N_9208,N_9011,N_9091);
nand U9209 (N_9209,N_9038,N_9069);
nand U9210 (N_9210,N_9066,N_9092);
xor U9211 (N_9211,N_9011,N_9029);
nand U9212 (N_9212,N_9030,N_9091);
and U9213 (N_9213,N_9025,N_9057);
or U9214 (N_9214,N_9115,N_9043);
or U9215 (N_9215,N_9105,N_9117);
nor U9216 (N_9216,N_9036,N_9011);
xor U9217 (N_9217,N_9000,N_9109);
xor U9218 (N_9218,N_9107,N_9106);
xnor U9219 (N_9219,N_9044,N_9103);
and U9220 (N_9220,N_9012,N_9079);
nand U9221 (N_9221,N_9089,N_9026);
xnor U9222 (N_9222,N_9008,N_9048);
xor U9223 (N_9223,N_9006,N_9086);
and U9224 (N_9224,N_9059,N_9046);
nor U9225 (N_9225,N_9092,N_9107);
and U9226 (N_9226,N_9080,N_9027);
nor U9227 (N_9227,N_9074,N_9029);
nand U9228 (N_9228,N_9119,N_9100);
nand U9229 (N_9229,N_9075,N_9011);
and U9230 (N_9230,N_9108,N_9112);
xnor U9231 (N_9231,N_9006,N_9065);
and U9232 (N_9232,N_9033,N_9002);
xor U9233 (N_9233,N_9031,N_9065);
nand U9234 (N_9234,N_9040,N_9119);
nand U9235 (N_9235,N_9051,N_9097);
nand U9236 (N_9236,N_9030,N_9029);
and U9237 (N_9237,N_9005,N_9065);
and U9238 (N_9238,N_9030,N_9106);
and U9239 (N_9239,N_9035,N_9033);
xor U9240 (N_9240,N_9104,N_9047);
nand U9241 (N_9241,N_9109,N_9108);
or U9242 (N_9242,N_9098,N_9002);
xnor U9243 (N_9243,N_9115,N_9099);
and U9244 (N_9244,N_9064,N_9094);
or U9245 (N_9245,N_9072,N_9098);
nand U9246 (N_9246,N_9003,N_9123);
and U9247 (N_9247,N_9009,N_9054);
xnor U9248 (N_9248,N_9107,N_9045);
nand U9249 (N_9249,N_9022,N_9102);
xnor U9250 (N_9250,N_9167,N_9125);
nor U9251 (N_9251,N_9249,N_9210);
or U9252 (N_9252,N_9215,N_9159);
and U9253 (N_9253,N_9133,N_9162);
nand U9254 (N_9254,N_9234,N_9220);
nor U9255 (N_9255,N_9142,N_9233);
and U9256 (N_9256,N_9160,N_9176);
and U9257 (N_9257,N_9187,N_9186);
or U9258 (N_9258,N_9140,N_9164);
nor U9259 (N_9259,N_9175,N_9132);
xnor U9260 (N_9260,N_9169,N_9185);
nand U9261 (N_9261,N_9136,N_9214);
nor U9262 (N_9262,N_9194,N_9157);
nor U9263 (N_9263,N_9203,N_9221);
nor U9264 (N_9264,N_9199,N_9246);
xnor U9265 (N_9265,N_9178,N_9173);
nor U9266 (N_9266,N_9216,N_9148);
xnor U9267 (N_9267,N_9206,N_9138);
nor U9268 (N_9268,N_9201,N_9241);
and U9269 (N_9269,N_9129,N_9128);
or U9270 (N_9270,N_9189,N_9161);
nor U9271 (N_9271,N_9180,N_9247);
nor U9272 (N_9272,N_9155,N_9166);
nand U9273 (N_9273,N_9228,N_9196);
nor U9274 (N_9274,N_9127,N_9143);
or U9275 (N_9275,N_9239,N_9126);
xnor U9276 (N_9276,N_9245,N_9181);
and U9277 (N_9277,N_9222,N_9182);
nor U9278 (N_9278,N_9146,N_9135);
and U9279 (N_9279,N_9218,N_9150);
or U9280 (N_9280,N_9158,N_9179);
or U9281 (N_9281,N_9154,N_9151);
xor U9282 (N_9282,N_9197,N_9248);
nor U9283 (N_9283,N_9144,N_9193);
xor U9284 (N_9284,N_9141,N_9137);
xnor U9285 (N_9285,N_9171,N_9198);
nand U9286 (N_9286,N_9225,N_9145);
or U9287 (N_9287,N_9204,N_9205);
nor U9288 (N_9288,N_9149,N_9231);
and U9289 (N_9289,N_9226,N_9223);
and U9290 (N_9290,N_9207,N_9163);
xor U9291 (N_9291,N_9243,N_9152);
or U9292 (N_9292,N_9217,N_9170);
nor U9293 (N_9293,N_9202,N_9213);
xor U9294 (N_9294,N_9235,N_9188);
and U9295 (N_9295,N_9236,N_9208);
nor U9296 (N_9296,N_9184,N_9227);
nand U9297 (N_9297,N_9195,N_9172);
nand U9298 (N_9298,N_9153,N_9139);
nand U9299 (N_9299,N_9219,N_9183);
xor U9300 (N_9300,N_9147,N_9244);
and U9301 (N_9301,N_9211,N_9224);
nand U9302 (N_9302,N_9209,N_9131);
nor U9303 (N_9303,N_9232,N_9177);
nor U9304 (N_9304,N_9192,N_9229);
or U9305 (N_9305,N_9242,N_9134);
xor U9306 (N_9306,N_9237,N_9191);
nand U9307 (N_9307,N_9174,N_9212);
nand U9308 (N_9308,N_9165,N_9240);
nor U9309 (N_9309,N_9168,N_9200);
or U9310 (N_9310,N_9130,N_9238);
and U9311 (N_9311,N_9156,N_9190);
and U9312 (N_9312,N_9230,N_9126);
nor U9313 (N_9313,N_9158,N_9132);
xor U9314 (N_9314,N_9246,N_9212);
nor U9315 (N_9315,N_9173,N_9129);
or U9316 (N_9316,N_9142,N_9147);
xor U9317 (N_9317,N_9211,N_9201);
or U9318 (N_9318,N_9213,N_9163);
nor U9319 (N_9319,N_9247,N_9235);
nor U9320 (N_9320,N_9176,N_9198);
and U9321 (N_9321,N_9210,N_9221);
and U9322 (N_9322,N_9234,N_9224);
and U9323 (N_9323,N_9201,N_9248);
nand U9324 (N_9324,N_9165,N_9223);
and U9325 (N_9325,N_9159,N_9220);
and U9326 (N_9326,N_9233,N_9148);
xor U9327 (N_9327,N_9190,N_9171);
or U9328 (N_9328,N_9204,N_9213);
xor U9329 (N_9329,N_9230,N_9224);
nor U9330 (N_9330,N_9194,N_9244);
or U9331 (N_9331,N_9172,N_9240);
nor U9332 (N_9332,N_9238,N_9184);
and U9333 (N_9333,N_9240,N_9236);
nor U9334 (N_9334,N_9163,N_9210);
xor U9335 (N_9335,N_9226,N_9137);
nand U9336 (N_9336,N_9221,N_9229);
nand U9337 (N_9337,N_9241,N_9235);
nor U9338 (N_9338,N_9194,N_9208);
nor U9339 (N_9339,N_9187,N_9199);
and U9340 (N_9340,N_9223,N_9201);
nor U9341 (N_9341,N_9237,N_9155);
or U9342 (N_9342,N_9201,N_9149);
nor U9343 (N_9343,N_9169,N_9132);
or U9344 (N_9344,N_9200,N_9226);
or U9345 (N_9345,N_9132,N_9139);
nor U9346 (N_9346,N_9191,N_9238);
nor U9347 (N_9347,N_9181,N_9172);
nor U9348 (N_9348,N_9241,N_9203);
nand U9349 (N_9349,N_9199,N_9226);
or U9350 (N_9350,N_9187,N_9180);
or U9351 (N_9351,N_9170,N_9147);
and U9352 (N_9352,N_9237,N_9199);
and U9353 (N_9353,N_9227,N_9159);
and U9354 (N_9354,N_9190,N_9181);
or U9355 (N_9355,N_9153,N_9148);
nor U9356 (N_9356,N_9164,N_9219);
nand U9357 (N_9357,N_9165,N_9162);
nand U9358 (N_9358,N_9222,N_9158);
nor U9359 (N_9359,N_9195,N_9187);
nand U9360 (N_9360,N_9143,N_9223);
or U9361 (N_9361,N_9167,N_9178);
xor U9362 (N_9362,N_9172,N_9140);
nor U9363 (N_9363,N_9150,N_9213);
xnor U9364 (N_9364,N_9145,N_9220);
nand U9365 (N_9365,N_9234,N_9174);
nand U9366 (N_9366,N_9181,N_9187);
or U9367 (N_9367,N_9171,N_9199);
nand U9368 (N_9368,N_9183,N_9203);
xnor U9369 (N_9369,N_9178,N_9247);
xor U9370 (N_9370,N_9205,N_9220);
or U9371 (N_9371,N_9155,N_9242);
nor U9372 (N_9372,N_9158,N_9211);
nand U9373 (N_9373,N_9180,N_9238);
or U9374 (N_9374,N_9191,N_9222);
xnor U9375 (N_9375,N_9309,N_9367);
or U9376 (N_9376,N_9291,N_9319);
xor U9377 (N_9377,N_9312,N_9303);
xor U9378 (N_9378,N_9329,N_9261);
and U9379 (N_9379,N_9264,N_9252);
nand U9380 (N_9380,N_9359,N_9307);
nor U9381 (N_9381,N_9292,N_9284);
or U9382 (N_9382,N_9374,N_9278);
xnor U9383 (N_9383,N_9330,N_9350);
and U9384 (N_9384,N_9320,N_9280);
nand U9385 (N_9385,N_9301,N_9373);
and U9386 (N_9386,N_9354,N_9362);
and U9387 (N_9387,N_9251,N_9257);
or U9388 (N_9388,N_9275,N_9315);
xor U9389 (N_9389,N_9349,N_9352);
nand U9390 (N_9390,N_9317,N_9255);
nor U9391 (N_9391,N_9364,N_9360);
and U9392 (N_9392,N_9297,N_9365);
and U9393 (N_9393,N_9316,N_9254);
or U9394 (N_9394,N_9273,N_9328);
or U9395 (N_9395,N_9263,N_9325);
or U9396 (N_9396,N_9260,N_9267);
nand U9397 (N_9397,N_9296,N_9340);
and U9398 (N_9398,N_9274,N_9361);
or U9399 (N_9399,N_9277,N_9289);
nor U9400 (N_9400,N_9294,N_9338);
and U9401 (N_9401,N_9356,N_9295);
nand U9402 (N_9402,N_9304,N_9293);
nor U9403 (N_9403,N_9347,N_9314);
xnor U9404 (N_9404,N_9271,N_9345);
and U9405 (N_9405,N_9268,N_9287);
nand U9406 (N_9406,N_9371,N_9348);
nor U9407 (N_9407,N_9336,N_9272);
xnor U9408 (N_9408,N_9334,N_9300);
nand U9409 (N_9409,N_9318,N_9372);
nand U9410 (N_9410,N_9265,N_9305);
or U9411 (N_9411,N_9333,N_9306);
or U9412 (N_9412,N_9331,N_9342);
or U9413 (N_9413,N_9308,N_9250);
nand U9414 (N_9414,N_9299,N_9262);
nand U9415 (N_9415,N_9324,N_9335);
or U9416 (N_9416,N_9253,N_9285);
or U9417 (N_9417,N_9366,N_9343);
or U9418 (N_9418,N_9286,N_9341);
nand U9419 (N_9419,N_9327,N_9281);
nor U9420 (N_9420,N_9310,N_9311);
or U9421 (N_9421,N_9344,N_9256);
xor U9422 (N_9422,N_9276,N_9258);
and U9423 (N_9423,N_9358,N_9321);
nand U9424 (N_9424,N_9283,N_9302);
xor U9425 (N_9425,N_9326,N_9298);
or U9426 (N_9426,N_9357,N_9323);
xor U9427 (N_9427,N_9269,N_9282);
nor U9428 (N_9428,N_9279,N_9322);
and U9429 (N_9429,N_9363,N_9313);
or U9430 (N_9430,N_9368,N_9346);
nor U9431 (N_9431,N_9259,N_9332);
or U9432 (N_9432,N_9339,N_9266);
nor U9433 (N_9433,N_9353,N_9369);
xnor U9434 (N_9434,N_9290,N_9337);
and U9435 (N_9435,N_9351,N_9355);
nand U9436 (N_9436,N_9270,N_9288);
or U9437 (N_9437,N_9370,N_9349);
nor U9438 (N_9438,N_9340,N_9301);
xnor U9439 (N_9439,N_9316,N_9280);
nand U9440 (N_9440,N_9345,N_9360);
xor U9441 (N_9441,N_9317,N_9263);
xnor U9442 (N_9442,N_9345,N_9374);
or U9443 (N_9443,N_9325,N_9271);
or U9444 (N_9444,N_9288,N_9314);
or U9445 (N_9445,N_9337,N_9278);
or U9446 (N_9446,N_9301,N_9362);
and U9447 (N_9447,N_9323,N_9267);
nand U9448 (N_9448,N_9267,N_9306);
or U9449 (N_9449,N_9363,N_9331);
nor U9450 (N_9450,N_9291,N_9328);
nand U9451 (N_9451,N_9362,N_9353);
or U9452 (N_9452,N_9254,N_9309);
and U9453 (N_9453,N_9299,N_9308);
and U9454 (N_9454,N_9317,N_9252);
or U9455 (N_9455,N_9372,N_9265);
nor U9456 (N_9456,N_9332,N_9364);
nand U9457 (N_9457,N_9335,N_9253);
nor U9458 (N_9458,N_9320,N_9265);
nand U9459 (N_9459,N_9363,N_9295);
or U9460 (N_9460,N_9327,N_9307);
nor U9461 (N_9461,N_9319,N_9279);
or U9462 (N_9462,N_9322,N_9356);
and U9463 (N_9463,N_9254,N_9360);
nor U9464 (N_9464,N_9335,N_9341);
nand U9465 (N_9465,N_9334,N_9372);
or U9466 (N_9466,N_9334,N_9282);
or U9467 (N_9467,N_9294,N_9286);
xor U9468 (N_9468,N_9344,N_9346);
nand U9469 (N_9469,N_9254,N_9354);
nand U9470 (N_9470,N_9353,N_9330);
nand U9471 (N_9471,N_9324,N_9336);
or U9472 (N_9472,N_9262,N_9270);
or U9473 (N_9473,N_9308,N_9271);
xor U9474 (N_9474,N_9329,N_9250);
nor U9475 (N_9475,N_9269,N_9325);
and U9476 (N_9476,N_9301,N_9279);
nor U9477 (N_9477,N_9333,N_9297);
nand U9478 (N_9478,N_9327,N_9316);
or U9479 (N_9479,N_9351,N_9297);
xor U9480 (N_9480,N_9283,N_9361);
or U9481 (N_9481,N_9283,N_9374);
nor U9482 (N_9482,N_9273,N_9290);
xor U9483 (N_9483,N_9352,N_9300);
nor U9484 (N_9484,N_9366,N_9350);
and U9485 (N_9485,N_9262,N_9274);
and U9486 (N_9486,N_9322,N_9321);
or U9487 (N_9487,N_9363,N_9266);
or U9488 (N_9488,N_9305,N_9341);
xor U9489 (N_9489,N_9262,N_9346);
xnor U9490 (N_9490,N_9278,N_9366);
or U9491 (N_9491,N_9322,N_9313);
xor U9492 (N_9492,N_9315,N_9291);
xor U9493 (N_9493,N_9324,N_9366);
nor U9494 (N_9494,N_9356,N_9292);
or U9495 (N_9495,N_9298,N_9333);
and U9496 (N_9496,N_9253,N_9353);
xnor U9497 (N_9497,N_9270,N_9254);
and U9498 (N_9498,N_9308,N_9350);
and U9499 (N_9499,N_9333,N_9259);
and U9500 (N_9500,N_9464,N_9496);
nand U9501 (N_9501,N_9414,N_9457);
xnor U9502 (N_9502,N_9475,N_9455);
nand U9503 (N_9503,N_9389,N_9398);
nor U9504 (N_9504,N_9468,N_9420);
nor U9505 (N_9505,N_9441,N_9425);
or U9506 (N_9506,N_9413,N_9432);
or U9507 (N_9507,N_9439,N_9395);
nor U9508 (N_9508,N_9481,N_9426);
or U9509 (N_9509,N_9458,N_9416);
nor U9510 (N_9510,N_9377,N_9436);
xnor U9511 (N_9511,N_9391,N_9386);
nand U9512 (N_9512,N_9411,N_9392);
xor U9513 (N_9513,N_9471,N_9460);
nand U9514 (N_9514,N_9415,N_9483);
and U9515 (N_9515,N_9440,N_9494);
and U9516 (N_9516,N_9423,N_9448);
xnor U9517 (N_9517,N_9401,N_9394);
and U9518 (N_9518,N_9491,N_9497);
and U9519 (N_9519,N_9495,N_9384);
and U9520 (N_9520,N_9378,N_9428);
nor U9521 (N_9521,N_9469,N_9467);
xnor U9522 (N_9522,N_9447,N_9486);
and U9523 (N_9523,N_9445,N_9476);
xnor U9524 (N_9524,N_9435,N_9480);
or U9525 (N_9525,N_9470,N_9383);
xnor U9526 (N_9526,N_9487,N_9408);
nor U9527 (N_9527,N_9402,N_9465);
or U9528 (N_9528,N_9430,N_9409);
xnor U9529 (N_9529,N_9442,N_9431);
xnor U9530 (N_9530,N_9388,N_9482);
and U9531 (N_9531,N_9412,N_9397);
or U9532 (N_9532,N_9419,N_9490);
nor U9533 (N_9533,N_9449,N_9407);
nor U9534 (N_9534,N_9399,N_9472);
nand U9535 (N_9535,N_9421,N_9387);
xnor U9536 (N_9536,N_9380,N_9463);
xor U9537 (N_9537,N_9479,N_9462);
or U9538 (N_9538,N_9452,N_9489);
xor U9539 (N_9539,N_9450,N_9473);
xor U9540 (N_9540,N_9459,N_9454);
or U9541 (N_9541,N_9406,N_9379);
xor U9542 (N_9542,N_9461,N_9418);
and U9543 (N_9543,N_9453,N_9444);
xnor U9544 (N_9544,N_9385,N_9484);
nand U9545 (N_9545,N_9403,N_9422);
and U9546 (N_9546,N_9417,N_9410);
nand U9547 (N_9547,N_9438,N_9493);
and U9548 (N_9548,N_9393,N_9466);
xnor U9549 (N_9549,N_9446,N_9382);
nor U9550 (N_9550,N_9478,N_9437);
nor U9551 (N_9551,N_9433,N_9405);
xnor U9552 (N_9552,N_9451,N_9499);
xor U9553 (N_9553,N_9390,N_9376);
nor U9554 (N_9554,N_9427,N_9474);
nand U9555 (N_9555,N_9492,N_9400);
nand U9556 (N_9556,N_9404,N_9381);
or U9557 (N_9557,N_9485,N_9456);
nor U9558 (N_9558,N_9488,N_9396);
xor U9559 (N_9559,N_9498,N_9424);
or U9560 (N_9560,N_9375,N_9477);
nand U9561 (N_9561,N_9443,N_9434);
nand U9562 (N_9562,N_9429,N_9455);
or U9563 (N_9563,N_9426,N_9472);
or U9564 (N_9564,N_9459,N_9424);
and U9565 (N_9565,N_9396,N_9413);
or U9566 (N_9566,N_9463,N_9461);
nor U9567 (N_9567,N_9427,N_9426);
and U9568 (N_9568,N_9385,N_9456);
nand U9569 (N_9569,N_9422,N_9458);
and U9570 (N_9570,N_9447,N_9483);
nor U9571 (N_9571,N_9457,N_9402);
nor U9572 (N_9572,N_9414,N_9408);
or U9573 (N_9573,N_9479,N_9447);
nor U9574 (N_9574,N_9422,N_9445);
and U9575 (N_9575,N_9481,N_9427);
xnor U9576 (N_9576,N_9495,N_9431);
or U9577 (N_9577,N_9433,N_9377);
xnor U9578 (N_9578,N_9382,N_9484);
xnor U9579 (N_9579,N_9438,N_9466);
and U9580 (N_9580,N_9451,N_9426);
or U9581 (N_9581,N_9465,N_9408);
nand U9582 (N_9582,N_9416,N_9491);
xor U9583 (N_9583,N_9447,N_9453);
xor U9584 (N_9584,N_9488,N_9456);
xnor U9585 (N_9585,N_9493,N_9394);
and U9586 (N_9586,N_9447,N_9435);
or U9587 (N_9587,N_9455,N_9413);
xnor U9588 (N_9588,N_9392,N_9450);
nor U9589 (N_9589,N_9393,N_9399);
nor U9590 (N_9590,N_9420,N_9415);
nor U9591 (N_9591,N_9470,N_9454);
or U9592 (N_9592,N_9380,N_9456);
nand U9593 (N_9593,N_9393,N_9422);
or U9594 (N_9594,N_9408,N_9498);
or U9595 (N_9595,N_9392,N_9479);
and U9596 (N_9596,N_9404,N_9441);
or U9597 (N_9597,N_9456,N_9442);
nor U9598 (N_9598,N_9484,N_9497);
or U9599 (N_9599,N_9408,N_9394);
or U9600 (N_9600,N_9455,N_9433);
xnor U9601 (N_9601,N_9425,N_9466);
xnor U9602 (N_9602,N_9435,N_9499);
or U9603 (N_9603,N_9479,N_9404);
nand U9604 (N_9604,N_9427,N_9387);
nor U9605 (N_9605,N_9389,N_9405);
nand U9606 (N_9606,N_9489,N_9406);
xor U9607 (N_9607,N_9465,N_9496);
nor U9608 (N_9608,N_9412,N_9442);
or U9609 (N_9609,N_9430,N_9426);
or U9610 (N_9610,N_9476,N_9452);
nor U9611 (N_9611,N_9490,N_9432);
nor U9612 (N_9612,N_9401,N_9490);
or U9613 (N_9613,N_9405,N_9462);
or U9614 (N_9614,N_9477,N_9389);
and U9615 (N_9615,N_9406,N_9465);
nand U9616 (N_9616,N_9410,N_9421);
or U9617 (N_9617,N_9482,N_9442);
and U9618 (N_9618,N_9488,N_9494);
and U9619 (N_9619,N_9427,N_9382);
and U9620 (N_9620,N_9393,N_9423);
nand U9621 (N_9621,N_9439,N_9418);
xnor U9622 (N_9622,N_9387,N_9485);
nor U9623 (N_9623,N_9428,N_9487);
xor U9624 (N_9624,N_9410,N_9408);
nor U9625 (N_9625,N_9545,N_9584);
nand U9626 (N_9626,N_9561,N_9560);
xor U9627 (N_9627,N_9619,N_9587);
nor U9628 (N_9628,N_9623,N_9592);
and U9629 (N_9629,N_9564,N_9500);
nor U9630 (N_9630,N_9549,N_9603);
and U9631 (N_9631,N_9503,N_9527);
nand U9632 (N_9632,N_9568,N_9604);
nor U9633 (N_9633,N_9530,N_9502);
nor U9634 (N_9634,N_9546,N_9501);
xnor U9635 (N_9635,N_9517,N_9504);
or U9636 (N_9636,N_9582,N_9511);
xor U9637 (N_9637,N_9507,N_9565);
nor U9638 (N_9638,N_9533,N_9512);
and U9639 (N_9639,N_9585,N_9596);
or U9640 (N_9640,N_9569,N_9621);
and U9641 (N_9641,N_9553,N_9528);
xor U9642 (N_9642,N_9577,N_9572);
nand U9643 (N_9643,N_9620,N_9522);
and U9644 (N_9644,N_9612,N_9594);
and U9645 (N_9645,N_9506,N_9570);
nor U9646 (N_9646,N_9566,N_9509);
or U9647 (N_9647,N_9543,N_9590);
xnor U9648 (N_9648,N_9550,N_9597);
and U9649 (N_9649,N_9591,N_9540);
nand U9650 (N_9650,N_9554,N_9515);
xor U9651 (N_9651,N_9529,N_9520);
and U9652 (N_9652,N_9562,N_9608);
and U9653 (N_9653,N_9513,N_9593);
nand U9654 (N_9654,N_9556,N_9536);
and U9655 (N_9655,N_9538,N_9600);
or U9656 (N_9656,N_9537,N_9524);
xor U9657 (N_9657,N_9516,N_9548);
nand U9658 (N_9658,N_9624,N_9578);
nand U9659 (N_9659,N_9575,N_9541);
nand U9660 (N_9660,N_9519,N_9544);
xnor U9661 (N_9661,N_9567,N_9579);
nand U9662 (N_9662,N_9605,N_9588);
nand U9663 (N_9663,N_9589,N_9558);
xnor U9664 (N_9664,N_9573,N_9615);
or U9665 (N_9665,N_9602,N_9622);
and U9666 (N_9666,N_9514,N_9598);
nand U9667 (N_9667,N_9532,N_9542);
or U9668 (N_9668,N_9557,N_9611);
and U9669 (N_9669,N_9555,N_9559);
nand U9670 (N_9670,N_9508,N_9599);
or U9671 (N_9671,N_9539,N_9574);
nor U9672 (N_9672,N_9616,N_9581);
and U9673 (N_9673,N_9614,N_9505);
nor U9674 (N_9674,N_9551,N_9595);
xor U9675 (N_9675,N_9535,N_9531);
nand U9676 (N_9676,N_9510,N_9552);
nor U9677 (N_9677,N_9617,N_9618);
or U9678 (N_9678,N_9610,N_9526);
nand U9679 (N_9679,N_9606,N_9613);
or U9680 (N_9680,N_9586,N_9583);
xnor U9681 (N_9681,N_9571,N_9607);
xnor U9682 (N_9682,N_9523,N_9525);
nor U9683 (N_9683,N_9518,N_9521);
or U9684 (N_9684,N_9601,N_9563);
or U9685 (N_9685,N_9576,N_9547);
or U9686 (N_9686,N_9609,N_9534);
nand U9687 (N_9687,N_9580,N_9535);
xnor U9688 (N_9688,N_9624,N_9502);
and U9689 (N_9689,N_9563,N_9500);
nand U9690 (N_9690,N_9555,N_9505);
nand U9691 (N_9691,N_9587,N_9602);
xor U9692 (N_9692,N_9520,N_9618);
or U9693 (N_9693,N_9565,N_9518);
nor U9694 (N_9694,N_9522,N_9502);
or U9695 (N_9695,N_9590,N_9520);
and U9696 (N_9696,N_9555,N_9564);
nand U9697 (N_9697,N_9531,N_9554);
or U9698 (N_9698,N_9514,N_9595);
nor U9699 (N_9699,N_9580,N_9585);
xor U9700 (N_9700,N_9516,N_9513);
xnor U9701 (N_9701,N_9536,N_9546);
nand U9702 (N_9702,N_9615,N_9554);
nor U9703 (N_9703,N_9520,N_9579);
or U9704 (N_9704,N_9543,N_9619);
xnor U9705 (N_9705,N_9602,N_9521);
nor U9706 (N_9706,N_9609,N_9517);
xnor U9707 (N_9707,N_9538,N_9620);
nand U9708 (N_9708,N_9595,N_9545);
nor U9709 (N_9709,N_9552,N_9530);
or U9710 (N_9710,N_9586,N_9548);
nor U9711 (N_9711,N_9576,N_9569);
nor U9712 (N_9712,N_9621,N_9597);
nand U9713 (N_9713,N_9566,N_9607);
or U9714 (N_9714,N_9609,N_9537);
and U9715 (N_9715,N_9529,N_9510);
nand U9716 (N_9716,N_9581,N_9597);
xor U9717 (N_9717,N_9500,N_9581);
nor U9718 (N_9718,N_9551,N_9582);
or U9719 (N_9719,N_9501,N_9527);
nor U9720 (N_9720,N_9523,N_9551);
nor U9721 (N_9721,N_9541,N_9525);
nor U9722 (N_9722,N_9542,N_9510);
or U9723 (N_9723,N_9616,N_9607);
or U9724 (N_9724,N_9604,N_9552);
and U9725 (N_9725,N_9544,N_9562);
xnor U9726 (N_9726,N_9620,N_9507);
or U9727 (N_9727,N_9508,N_9567);
xnor U9728 (N_9728,N_9544,N_9612);
nor U9729 (N_9729,N_9614,N_9553);
nor U9730 (N_9730,N_9508,N_9500);
or U9731 (N_9731,N_9568,N_9575);
nand U9732 (N_9732,N_9521,N_9536);
or U9733 (N_9733,N_9522,N_9596);
and U9734 (N_9734,N_9546,N_9572);
xor U9735 (N_9735,N_9543,N_9604);
and U9736 (N_9736,N_9589,N_9520);
or U9737 (N_9737,N_9616,N_9537);
xnor U9738 (N_9738,N_9588,N_9520);
nand U9739 (N_9739,N_9594,N_9548);
nand U9740 (N_9740,N_9552,N_9623);
xnor U9741 (N_9741,N_9536,N_9616);
or U9742 (N_9742,N_9599,N_9572);
or U9743 (N_9743,N_9602,N_9590);
nor U9744 (N_9744,N_9558,N_9599);
xnor U9745 (N_9745,N_9565,N_9574);
and U9746 (N_9746,N_9513,N_9621);
xnor U9747 (N_9747,N_9538,N_9522);
xnor U9748 (N_9748,N_9556,N_9610);
nor U9749 (N_9749,N_9586,N_9518);
xnor U9750 (N_9750,N_9688,N_9689);
and U9751 (N_9751,N_9659,N_9634);
xor U9752 (N_9752,N_9675,N_9698);
and U9753 (N_9753,N_9732,N_9717);
xnor U9754 (N_9754,N_9644,N_9645);
xor U9755 (N_9755,N_9735,N_9636);
nor U9756 (N_9756,N_9683,N_9707);
and U9757 (N_9757,N_9697,N_9640);
or U9758 (N_9758,N_9670,N_9712);
or U9759 (N_9759,N_9638,N_9684);
or U9760 (N_9760,N_9694,N_9674);
or U9761 (N_9761,N_9678,N_9700);
and U9762 (N_9762,N_9741,N_9711);
xnor U9763 (N_9763,N_9666,N_9733);
nor U9764 (N_9764,N_9661,N_9643);
or U9765 (N_9765,N_9647,N_9627);
and U9766 (N_9766,N_9710,N_9696);
and U9767 (N_9767,N_9651,N_9704);
nor U9768 (N_9768,N_9718,N_9703);
or U9769 (N_9769,N_9695,N_9691);
xor U9770 (N_9770,N_9748,N_9692);
or U9771 (N_9771,N_9629,N_9726);
xor U9772 (N_9772,N_9723,N_9637);
xor U9773 (N_9773,N_9719,N_9722);
and U9774 (N_9774,N_9709,N_9731);
xnor U9775 (N_9775,N_9693,N_9746);
or U9776 (N_9776,N_9669,N_9699);
xor U9777 (N_9777,N_9631,N_9662);
nor U9778 (N_9778,N_9736,N_9702);
nand U9779 (N_9779,N_9749,N_9652);
nor U9780 (N_9780,N_9668,N_9641);
xor U9781 (N_9781,N_9677,N_9715);
nor U9782 (N_9782,N_9655,N_9639);
nor U9783 (N_9783,N_9743,N_9682);
nor U9784 (N_9784,N_9633,N_9660);
nor U9785 (N_9785,N_9686,N_9642);
nor U9786 (N_9786,N_9744,N_9657);
nor U9787 (N_9787,N_9650,N_9747);
or U9788 (N_9788,N_9664,N_9671);
or U9789 (N_9789,N_9721,N_9673);
nor U9790 (N_9790,N_9658,N_9656);
xnor U9791 (N_9791,N_9730,N_9740);
nor U9792 (N_9792,N_9680,N_9690);
xor U9793 (N_9793,N_9729,N_9714);
xor U9794 (N_9794,N_9734,N_9628);
and U9795 (N_9795,N_9716,N_9679);
and U9796 (N_9796,N_9708,N_9648);
nand U9797 (N_9797,N_9672,N_9654);
nand U9798 (N_9798,N_9701,N_9667);
xor U9799 (N_9799,N_9738,N_9724);
nor U9800 (N_9800,N_9739,N_9737);
and U9801 (N_9801,N_9635,N_9649);
xor U9802 (N_9802,N_9706,N_9713);
xnor U9803 (N_9803,N_9720,N_9676);
nand U9804 (N_9804,N_9630,N_9687);
nand U9805 (N_9805,N_9685,N_9725);
xor U9806 (N_9806,N_9742,N_9632);
nand U9807 (N_9807,N_9625,N_9745);
and U9808 (N_9808,N_9626,N_9665);
and U9809 (N_9809,N_9663,N_9728);
xnor U9810 (N_9810,N_9646,N_9705);
xnor U9811 (N_9811,N_9681,N_9653);
nand U9812 (N_9812,N_9727,N_9698);
nand U9813 (N_9813,N_9639,N_9746);
and U9814 (N_9814,N_9643,N_9664);
nor U9815 (N_9815,N_9706,N_9720);
nand U9816 (N_9816,N_9667,N_9689);
or U9817 (N_9817,N_9663,N_9708);
xnor U9818 (N_9818,N_9633,N_9676);
nor U9819 (N_9819,N_9710,N_9694);
xor U9820 (N_9820,N_9667,N_9681);
nor U9821 (N_9821,N_9747,N_9691);
and U9822 (N_9822,N_9723,N_9693);
and U9823 (N_9823,N_9732,N_9735);
xnor U9824 (N_9824,N_9725,N_9686);
nand U9825 (N_9825,N_9736,N_9662);
xor U9826 (N_9826,N_9658,N_9675);
nand U9827 (N_9827,N_9701,N_9666);
and U9828 (N_9828,N_9709,N_9677);
xnor U9829 (N_9829,N_9718,N_9709);
nor U9830 (N_9830,N_9703,N_9740);
nand U9831 (N_9831,N_9653,N_9643);
nor U9832 (N_9832,N_9694,N_9729);
nand U9833 (N_9833,N_9691,N_9745);
or U9834 (N_9834,N_9658,N_9737);
and U9835 (N_9835,N_9628,N_9643);
xor U9836 (N_9836,N_9704,N_9695);
and U9837 (N_9837,N_9703,N_9631);
or U9838 (N_9838,N_9651,N_9691);
nand U9839 (N_9839,N_9673,N_9694);
nor U9840 (N_9840,N_9695,N_9690);
xnor U9841 (N_9841,N_9626,N_9712);
and U9842 (N_9842,N_9643,N_9696);
xnor U9843 (N_9843,N_9686,N_9723);
nand U9844 (N_9844,N_9718,N_9683);
nor U9845 (N_9845,N_9721,N_9668);
or U9846 (N_9846,N_9691,N_9650);
nand U9847 (N_9847,N_9724,N_9740);
or U9848 (N_9848,N_9686,N_9730);
and U9849 (N_9849,N_9632,N_9699);
and U9850 (N_9850,N_9719,N_9736);
nand U9851 (N_9851,N_9675,N_9679);
nor U9852 (N_9852,N_9715,N_9730);
nand U9853 (N_9853,N_9680,N_9639);
or U9854 (N_9854,N_9671,N_9713);
or U9855 (N_9855,N_9677,N_9650);
and U9856 (N_9856,N_9708,N_9720);
or U9857 (N_9857,N_9667,N_9637);
xor U9858 (N_9858,N_9712,N_9729);
xor U9859 (N_9859,N_9664,N_9729);
and U9860 (N_9860,N_9730,N_9732);
xor U9861 (N_9861,N_9727,N_9650);
nand U9862 (N_9862,N_9674,N_9638);
xnor U9863 (N_9863,N_9641,N_9702);
or U9864 (N_9864,N_9737,N_9626);
or U9865 (N_9865,N_9692,N_9661);
nor U9866 (N_9866,N_9702,N_9730);
nor U9867 (N_9867,N_9671,N_9705);
or U9868 (N_9868,N_9668,N_9725);
and U9869 (N_9869,N_9715,N_9645);
nor U9870 (N_9870,N_9746,N_9711);
or U9871 (N_9871,N_9669,N_9651);
nor U9872 (N_9872,N_9669,N_9637);
xor U9873 (N_9873,N_9655,N_9659);
and U9874 (N_9874,N_9664,N_9678);
nor U9875 (N_9875,N_9802,N_9841);
and U9876 (N_9876,N_9793,N_9781);
or U9877 (N_9877,N_9816,N_9837);
xor U9878 (N_9878,N_9768,N_9824);
nand U9879 (N_9879,N_9845,N_9815);
xor U9880 (N_9880,N_9866,N_9753);
or U9881 (N_9881,N_9804,N_9822);
nor U9882 (N_9882,N_9758,N_9828);
xnor U9883 (N_9883,N_9850,N_9806);
nand U9884 (N_9884,N_9790,N_9829);
xor U9885 (N_9885,N_9860,N_9859);
and U9886 (N_9886,N_9799,N_9826);
nand U9887 (N_9887,N_9807,N_9780);
nand U9888 (N_9888,N_9760,N_9801);
or U9889 (N_9889,N_9840,N_9764);
nor U9890 (N_9890,N_9791,N_9770);
or U9891 (N_9891,N_9797,N_9812);
xor U9892 (N_9892,N_9755,N_9846);
nand U9893 (N_9893,N_9789,N_9847);
xnor U9894 (N_9894,N_9874,N_9833);
nand U9895 (N_9895,N_9834,N_9838);
or U9896 (N_9896,N_9783,N_9861);
xor U9897 (N_9897,N_9794,N_9792);
xnor U9898 (N_9898,N_9856,N_9765);
nand U9899 (N_9899,N_9777,N_9870);
and U9900 (N_9900,N_9769,N_9821);
xor U9901 (N_9901,N_9773,N_9803);
and U9902 (N_9902,N_9843,N_9762);
or U9903 (N_9903,N_9863,N_9819);
and U9904 (N_9904,N_9867,N_9752);
xnor U9905 (N_9905,N_9786,N_9756);
and U9906 (N_9906,N_9825,N_9779);
or U9907 (N_9907,N_9817,N_9858);
or U9908 (N_9908,N_9811,N_9788);
and U9909 (N_9909,N_9831,N_9872);
xor U9910 (N_9910,N_9862,N_9808);
nor U9911 (N_9911,N_9772,N_9853);
and U9912 (N_9912,N_9771,N_9763);
xor U9913 (N_9913,N_9782,N_9849);
nor U9914 (N_9914,N_9864,N_9842);
nand U9915 (N_9915,N_9836,N_9823);
and U9916 (N_9916,N_9754,N_9775);
and U9917 (N_9917,N_9751,N_9839);
nor U9918 (N_9918,N_9827,N_9851);
nand U9919 (N_9919,N_9865,N_9761);
xor U9920 (N_9920,N_9787,N_9813);
or U9921 (N_9921,N_9798,N_9795);
nand U9922 (N_9922,N_9848,N_9810);
nor U9923 (N_9923,N_9776,N_9857);
nor U9924 (N_9924,N_9805,N_9855);
or U9925 (N_9925,N_9818,N_9873);
or U9926 (N_9926,N_9785,N_9809);
nand U9927 (N_9927,N_9869,N_9820);
xor U9928 (N_9928,N_9757,N_9832);
or U9929 (N_9929,N_9796,N_9759);
xor U9930 (N_9930,N_9814,N_9844);
xnor U9931 (N_9931,N_9800,N_9835);
nand U9932 (N_9932,N_9750,N_9868);
nand U9933 (N_9933,N_9774,N_9778);
and U9934 (N_9934,N_9766,N_9852);
or U9935 (N_9935,N_9871,N_9830);
nand U9936 (N_9936,N_9767,N_9784);
xor U9937 (N_9937,N_9854,N_9756);
xnor U9938 (N_9938,N_9841,N_9809);
or U9939 (N_9939,N_9791,N_9858);
nand U9940 (N_9940,N_9812,N_9835);
nand U9941 (N_9941,N_9796,N_9828);
and U9942 (N_9942,N_9777,N_9757);
or U9943 (N_9943,N_9781,N_9839);
or U9944 (N_9944,N_9760,N_9805);
and U9945 (N_9945,N_9861,N_9807);
and U9946 (N_9946,N_9828,N_9831);
or U9947 (N_9947,N_9840,N_9864);
nand U9948 (N_9948,N_9753,N_9807);
nand U9949 (N_9949,N_9774,N_9828);
or U9950 (N_9950,N_9837,N_9824);
nand U9951 (N_9951,N_9858,N_9847);
or U9952 (N_9952,N_9779,N_9869);
and U9953 (N_9953,N_9811,N_9789);
xor U9954 (N_9954,N_9833,N_9816);
and U9955 (N_9955,N_9847,N_9872);
or U9956 (N_9956,N_9750,N_9839);
or U9957 (N_9957,N_9804,N_9803);
and U9958 (N_9958,N_9829,N_9836);
or U9959 (N_9959,N_9824,N_9836);
nand U9960 (N_9960,N_9793,N_9803);
xor U9961 (N_9961,N_9822,N_9814);
or U9962 (N_9962,N_9825,N_9805);
nand U9963 (N_9963,N_9814,N_9871);
and U9964 (N_9964,N_9761,N_9856);
and U9965 (N_9965,N_9802,N_9800);
or U9966 (N_9966,N_9797,N_9776);
and U9967 (N_9967,N_9806,N_9837);
and U9968 (N_9968,N_9861,N_9774);
xnor U9969 (N_9969,N_9862,N_9840);
xnor U9970 (N_9970,N_9852,N_9758);
nor U9971 (N_9971,N_9834,N_9792);
and U9972 (N_9972,N_9854,N_9861);
xor U9973 (N_9973,N_9840,N_9753);
nor U9974 (N_9974,N_9803,N_9805);
nand U9975 (N_9975,N_9844,N_9751);
or U9976 (N_9976,N_9862,N_9794);
and U9977 (N_9977,N_9821,N_9776);
nand U9978 (N_9978,N_9838,N_9866);
xor U9979 (N_9979,N_9806,N_9785);
or U9980 (N_9980,N_9862,N_9778);
xor U9981 (N_9981,N_9750,N_9775);
nand U9982 (N_9982,N_9863,N_9811);
or U9983 (N_9983,N_9783,N_9806);
xnor U9984 (N_9984,N_9819,N_9832);
and U9985 (N_9985,N_9772,N_9817);
nand U9986 (N_9986,N_9752,N_9794);
nor U9987 (N_9987,N_9845,N_9798);
nand U9988 (N_9988,N_9811,N_9799);
nand U9989 (N_9989,N_9867,N_9837);
nand U9990 (N_9990,N_9868,N_9858);
nand U9991 (N_9991,N_9848,N_9830);
xor U9992 (N_9992,N_9781,N_9790);
or U9993 (N_9993,N_9771,N_9871);
xor U9994 (N_9994,N_9848,N_9803);
and U9995 (N_9995,N_9811,N_9797);
nor U9996 (N_9996,N_9817,N_9849);
and U9997 (N_9997,N_9754,N_9788);
or U9998 (N_9998,N_9756,N_9873);
nand U9999 (N_9999,N_9808,N_9828);
xnor U10000 (N_10000,N_9923,N_9969);
or U10001 (N_10001,N_9958,N_9935);
nand U10002 (N_10002,N_9903,N_9936);
xnor U10003 (N_10003,N_9999,N_9994);
or U10004 (N_10004,N_9891,N_9884);
and U10005 (N_10005,N_9879,N_9991);
and U10006 (N_10006,N_9886,N_9909);
nor U10007 (N_10007,N_9918,N_9967);
or U10008 (N_10008,N_9897,N_9914);
nand U10009 (N_10009,N_9993,N_9934);
nor U10010 (N_10010,N_9910,N_9920);
xor U10011 (N_10011,N_9921,N_9953);
xnor U10012 (N_10012,N_9950,N_9929);
nand U10013 (N_10013,N_9945,N_9948);
and U10014 (N_10014,N_9988,N_9942);
nand U10015 (N_10015,N_9959,N_9882);
and U10016 (N_10016,N_9980,N_9960);
xnor U10017 (N_10017,N_9916,N_9962);
xnor U10018 (N_10018,N_9976,N_9965);
or U10019 (N_10019,N_9981,N_9968);
nor U10020 (N_10020,N_9892,N_9915);
xor U10021 (N_10021,N_9971,N_9997);
and U10022 (N_10022,N_9901,N_9913);
or U10023 (N_10023,N_9899,N_9970);
or U10024 (N_10024,N_9931,N_9990);
nor U10025 (N_10025,N_9954,N_9937);
and U10026 (N_10026,N_9930,N_9894);
and U10027 (N_10027,N_9964,N_9900);
and U10028 (N_10028,N_9978,N_9917);
nor U10029 (N_10029,N_9922,N_9941);
or U10030 (N_10030,N_9992,N_9911);
nand U10031 (N_10031,N_9946,N_9949);
and U10032 (N_10032,N_9926,N_9956);
or U10033 (N_10033,N_9876,N_9888);
nor U10034 (N_10034,N_9982,N_9986);
nand U10035 (N_10035,N_9933,N_9974);
nand U10036 (N_10036,N_9893,N_9972);
xor U10037 (N_10037,N_9989,N_9905);
nor U10038 (N_10038,N_9938,N_9961);
or U10039 (N_10039,N_9895,N_9907);
nor U10040 (N_10040,N_9995,N_9875);
and U10041 (N_10041,N_9889,N_9966);
xnor U10042 (N_10042,N_9955,N_9943);
nor U10043 (N_10043,N_9890,N_9883);
xor U10044 (N_10044,N_9885,N_9979);
nand U10045 (N_10045,N_9940,N_9996);
nor U10046 (N_10046,N_9977,N_9904);
and U10047 (N_10047,N_9912,N_9881);
xor U10048 (N_10048,N_9928,N_9963);
or U10049 (N_10049,N_9906,N_9925);
and U10050 (N_10050,N_9898,N_9983);
nor U10051 (N_10051,N_9932,N_9987);
and U10052 (N_10052,N_9975,N_9973);
or U10053 (N_10053,N_9877,N_9919);
nor U10054 (N_10054,N_9985,N_9944);
nand U10055 (N_10055,N_9927,N_9908);
and U10056 (N_10056,N_9952,N_9896);
xnor U10057 (N_10057,N_9951,N_9947);
and U10058 (N_10058,N_9878,N_9998);
or U10059 (N_10059,N_9887,N_9939);
xor U10060 (N_10060,N_9984,N_9902);
and U10061 (N_10061,N_9924,N_9880);
nor U10062 (N_10062,N_9957,N_9887);
nand U10063 (N_10063,N_9890,N_9907);
and U10064 (N_10064,N_9967,N_9911);
and U10065 (N_10065,N_9901,N_9894);
nor U10066 (N_10066,N_9949,N_9968);
and U10067 (N_10067,N_9947,N_9882);
xor U10068 (N_10068,N_9961,N_9935);
and U10069 (N_10069,N_9944,N_9932);
or U10070 (N_10070,N_9875,N_9950);
or U10071 (N_10071,N_9973,N_9892);
xor U10072 (N_10072,N_9976,N_9962);
or U10073 (N_10073,N_9994,N_9961);
nor U10074 (N_10074,N_9985,N_9965);
and U10075 (N_10075,N_9996,N_9882);
and U10076 (N_10076,N_9988,N_9886);
nand U10077 (N_10077,N_9984,N_9919);
nand U10078 (N_10078,N_9906,N_9956);
nor U10079 (N_10079,N_9899,N_9998);
or U10080 (N_10080,N_9969,N_9968);
and U10081 (N_10081,N_9940,N_9891);
nand U10082 (N_10082,N_9979,N_9981);
or U10083 (N_10083,N_9944,N_9951);
xnor U10084 (N_10084,N_9937,N_9923);
xor U10085 (N_10085,N_9892,N_9901);
or U10086 (N_10086,N_9999,N_9883);
xor U10087 (N_10087,N_9906,N_9890);
nor U10088 (N_10088,N_9892,N_9912);
xor U10089 (N_10089,N_9916,N_9934);
nand U10090 (N_10090,N_9976,N_9914);
xnor U10091 (N_10091,N_9917,N_9948);
and U10092 (N_10092,N_9939,N_9915);
xor U10093 (N_10093,N_9900,N_9918);
and U10094 (N_10094,N_9969,N_9937);
nor U10095 (N_10095,N_9944,N_9885);
nor U10096 (N_10096,N_9935,N_9968);
xnor U10097 (N_10097,N_9881,N_9895);
xnor U10098 (N_10098,N_9995,N_9892);
xor U10099 (N_10099,N_9897,N_9921);
or U10100 (N_10100,N_9922,N_9913);
and U10101 (N_10101,N_9945,N_9976);
or U10102 (N_10102,N_9970,N_9911);
nand U10103 (N_10103,N_9958,N_9928);
or U10104 (N_10104,N_9980,N_9897);
xor U10105 (N_10105,N_9968,N_9987);
nor U10106 (N_10106,N_9939,N_9968);
or U10107 (N_10107,N_9942,N_9998);
nand U10108 (N_10108,N_9884,N_9944);
xnor U10109 (N_10109,N_9965,N_9937);
nand U10110 (N_10110,N_9895,N_9878);
nand U10111 (N_10111,N_9927,N_9902);
and U10112 (N_10112,N_9953,N_9881);
and U10113 (N_10113,N_9922,N_9880);
or U10114 (N_10114,N_9891,N_9952);
nor U10115 (N_10115,N_9961,N_9962);
nand U10116 (N_10116,N_9990,N_9884);
and U10117 (N_10117,N_9966,N_9897);
or U10118 (N_10118,N_9974,N_9972);
nand U10119 (N_10119,N_9966,N_9941);
and U10120 (N_10120,N_9916,N_9982);
nor U10121 (N_10121,N_9893,N_9890);
nand U10122 (N_10122,N_9904,N_9965);
nor U10123 (N_10123,N_9883,N_9955);
nand U10124 (N_10124,N_9902,N_9876);
and U10125 (N_10125,N_10057,N_10043);
or U10126 (N_10126,N_10067,N_10054);
nor U10127 (N_10127,N_10066,N_10016);
xnor U10128 (N_10128,N_10072,N_10090);
and U10129 (N_10129,N_10011,N_10058);
and U10130 (N_10130,N_10048,N_10038);
nor U10131 (N_10131,N_10076,N_10022);
nand U10132 (N_10132,N_10093,N_10085);
xor U10133 (N_10133,N_10020,N_10112);
xnor U10134 (N_10134,N_10094,N_10092);
nor U10135 (N_10135,N_10102,N_10089);
and U10136 (N_10136,N_10026,N_10025);
nand U10137 (N_10137,N_10095,N_10006);
or U10138 (N_10138,N_10070,N_10003);
xnor U10139 (N_10139,N_10047,N_10036);
xnor U10140 (N_10140,N_10059,N_10060);
or U10141 (N_10141,N_10064,N_10077);
and U10142 (N_10142,N_10039,N_10024);
xor U10143 (N_10143,N_10082,N_10027);
nand U10144 (N_10144,N_10046,N_10033);
and U10145 (N_10145,N_10028,N_10091);
and U10146 (N_10146,N_10008,N_10081);
nor U10147 (N_10147,N_10042,N_10015);
nand U10148 (N_10148,N_10034,N_10084);
nor U10149 (N_10149,N_10100,N_10103);
and U10150 (N_10150,N_10080,N_10114);
xor U10151 (N_10151,N_10001,N_10083);
xor U10152 (N_10152,N_10010,N_10041);
or U10153 (N_10153,N_10104,N_10118);
nor U10154 (N_10154,N_10052,N_10055);
xor U10155 (N_10155,N_10049,N_10107);
and U10156 (N_10156,N_10037,N_10044);
or U10157 (N_10157,N_10021,N_10074);
nand U10158 (N_10158,N_10014,N_10073);
nor U10159 (N_10159,N_10009,N_10029);
nor U10160 (N_10160,N_10079,N_10062);
nand U10161 (N_10161,N_10086,N_10035);
and U10162 (N_10162,N_10099,N_10121);
nor U10163 (N_10163,N_10123,N_10111);
nand U10164 (N_10164,N_10105,N_10088);
and U10165 (N_10165,N_10017,N_10071);
xnor U10166 (N_10166,N_10023,N_10106);
or U10167 (N_10167,N_10019,N_10098);
xnor U10168 (N_10168,N_10063,N_10117);
or U10169 (N_10169,N_10051,N_10065);
xor U10170 (N_10170,N_10110,N_10087);
xor U10171 (N_10171,N_10120,N_10056);
nand U10172 (N_10172,N_10113,N_10030);
or U10173 (N_10173,N_10078,N_10002);
xor U10174 (N_10174,N_10096,N_10013);
nand U10175 (N_10175,N_10032,N_10122);
xnor U10176 (N_10176,N_10115,N_10050);
nand U10177 (N_10177,N_10119,N_10069);
xor U10178 (N_10178,N_10000,N_10061);
or U10179 (N_10179,N_10097,N_10124);
or U10180 (N_10180,N_10005,N_10108);
nand U10181 (N_10181,N_10101,N_10045);
nand U10182 (N_10182,N_10004,N_10040);
xnor U10183 (N_10183,N_10018,N_10109);
and U10184 (N_10184,N_10116,N_10012);
or U10185 (N_10185,N_10075,N_10068);
nor U10186 (N_10186,N_10007,N_10031);
and U10187 (N_10187,N_10053,N_10050);
and U10188 (N_10188,N_10090,N_10114);
nand U10189 (N_10189,N_10109,N_10099);
xnor U10190 (N_10190,N_10114,N_10031);
xor U10191 (N_10191,N_10090,N_10004);
and U10192 (N_10192,N_10093,N_10053);
or U10193 (N_10193,N_10057,N_10086);
nand U10194 (N_10194,N_10091,N_10103);
nand U10195 (N_10195,N_10005,N_10034);
and U10196 (N_10196,N_10046,N_10082);
or U10197 (N_10197,N_10105,N_10121);
and U10198 (N_10198,N_10065,N_10102);
or U10199 (N_10199,N_10010,N_10075);
nor U10200 (N_10200,N_10054,N_10045);
nand U10201 (N_10201,N_10086,N_10089);
xnor U10202 (N_10202,N_10124,N_10002);
nor U10203 (N_10203,N_10100,N_10102);
and U10204 (N_10204,N_10022,N_10106);
or U10205 (N_10205,N_10046,N_10068);
and U10206 (N_10206,N_10054,N_10107);
or U10207 (N_10207,N_10073,N_10097);
and U10208 (N_10208,N_10105,N_10090);
or U10209 (N_10209,N_10096,N_10118);
nor U10210 (N_10210,N_10033,N_10108);
and U10211 (N_10211,N_10081,N_10043);
or U10212 (N_10212,N_10018,N_10000);
and U10213 (N_10213,N_10071,N_10101);
or U10214 (N_10214,N_10007,N_10086);
nand U10215 (N_10215,N_10107,N_10003);
or U10216 (N_10216,N_10097,N_10043);
or U10217 (N_10217,N_10020,N_10117);
xnor U10218 (N_10218,N_10044,N_10094);
xor U10219 (N_10219,N_10043,N_10068);
xor U10220 (N_10220,N_10049,N_10043);
xor U10221 (N_10221,N_10030,N_10088);
and U10222 (N_10222,N_10054,N_10027);
xor U10223 (N_10223,N_10031,N_10083);
or U10224 (N_10224,N_10022,N_10085);
xnor U10225 (N_10225,N_10045,N_10069);
nor U10226 (N_10226,N_10024,N_10117);
nand U10227 (N_10227,N_10023,N_10016);
and U10228 (N_10228,N_10114,N_10016);
nor U10229 (N_10229,N_10095,N_10009);
xor U10230 (N_10230,N_10006,N_10077);
or U10231 (N_10231,N_10041,N_10081);
nand U10232 (N_10232,N_10050,N_10101);
xor U10233 (N_10233,N_10074,N_10055);
xnor U10234 (N_10234,N_10110,N_10016);
nand U10235 (N_10235,N_10073,N_10121);
nand U10236 (N_10236,N_10087,N_10006);
xnor U10237 (N_10237,N_10108,N_10120);
nor U10238 (N_10238,N_10024,N_10014);
and U10239 (N_10239,N_10059,N_10024);
nor U10240 (N_10240,N_10078,N_10103);
xnor U10241 (N_10241,N_10078,N_10052);
or U10242 (N_10242,N_10018,N_10110);
and U10243 (N_10243,N_10081,N_10068);
or U10244 (N_10244,N_10041,N_10062);
nand U10245 (N_10245,N_10112,N_10017);
xor U10246 (N_10246,N_10027,N_10085);
or U10247 (N_10247,N_10098,N_10086);
xnor U10248 (N_10248,N_10038,N_10115);
nor U10249 (N_10249,N_10102,N_10024);
or U10250 (N_10250,N_10191,N_10216);
nor U10251 (N_10251,N_10181,N_10160);
nor U10252 (N_10252,N_10147,N_10174);
nor U10253 (N_10253,N_10221,N_10145);
xor U10254 (N_10254,N_10141,N_10143);
and U10255 (N_10255,N_10235,N_10157);
nor U10256 (N_10256,N_10247,N_10173);
and U10257 (N_10257,N_10214,N_10146);
and U10258 (N_10258,N_10177,N_10217);
and U10259 (N_10259,N_10195,N_10197);
and U10260 (N_10260,N_10189,N_10152);
nor U10261 (N_10261,N_10194,N_10150);
and U10262 (N_10262,N_10224,N_10219);
nor U10263 (N_10263,N_10155,N_10223);
and U10264 (N_10264,N_10153,N_10161);
and U10265 (N_10265,N_10137,N_10234);
nand U10266 (N_10266,N_10245,N_10156);
or U10267 (N_10267,N_10188,N_10164);
or U10268 (N_10268,N_10151,N_10227);
xor U10269 (N_10269,N_10233,N_10139);
nand U10270 (N_10270,N_10163,N_10236);
and U10271 (N_10271,N_10184,N_10138);
nor U10272 (N_10272,N_10212,N_10179);
nor U10273 (N_10273,N_10185,N_10244);
and U10274 (N_10274,N_10211,N_10169);
and U10275 (N_10275,N_10207,N_10192);
nor U10276 (N_10276,N_10232,N_10220);
nand U10277 (N_10277,N_10222,N_10162);
xnor U10278 (N_10278,N_10142,N_10196);
nand U10279 (N_10279,N_10215,N_10186);
xor U10280 (N_10280,N_10131,N_10190);
nor U10281 (N_10281,N_10134,N_10127);
xor U10282 (N_10282,N_10136,N_10210);
xor U10283 (N_10283,N_10135,N_10241);
xor U10284 (N_10284,N_10159,N_10182);
xor U10285 (N_10285,N_10218,N_10239);
or U10286 (N_10286,N_10133,N_10199);
nand U10287 (N_10287,N_10237,N_10132);
xnor U10288 (N_10288,N_10148,N_10230);
nand U10289 (N_10289,N_10165,N_10140);
xor U10290 (N_10290,N_10213,N_10125);
or U10291 (N_10291,N_10238,N_10240);
and U10292 (N_10292,N_10248,N_10209);
and U10293 (N_10293,N_10193,N_10168);
or U10294 (N_10294,N_10229,N_10130);
or U10295 (N_10295,N_10144,N_10154);
xnor U10296 (N_10296,N_10166,N_10225);
xnor U10297 (N_10297,N_10249,N_10201);
nand U10298 (N_10298,N_10242,N_10171);
xnor U10299 (N_10299,N_10178,N_10205);
xnor U10300 (N_10300,N_10129,N_10204);
xnor U10301 (N_10301,N_10180,N_10246);
nand U10302 (N_10302,N_10208,N_10128);
xor U10303 (N_10303,N_10172,N_10167);
and U10304 (N_10304,N_10183,N_10243);
or U10305 (N_10305,N_10206,N_10149);
or U10306 (N_10306,N_10176,N_10198);
xor U10307 (N_10307,N_10202,N_10126);
and U10308 (N_10308,N_10228,N_10231);
xor U10309 (N_10309,N_10158,N_10226);
xor U10310 (N_10310,N_10175,N_10203);
or U10311 (N_10311,N_10187,N_10200);
and U10312 (N_10312,N_10170,N_10193);
nor U10313 (N_10313,N_10162,N_10139);
and U10314 (N_10314,N_10226,N_10151);
and U10315 (N_10315,N_10192,N_10162);
xor U10316 (N_10316,N_10249,N_10161);
or U10317 (N_10317,N_10130,N_10153);
and U10318 (N_10318,N_10180,N_10147);
and U10319 (N_10319,N_10189,N_10139);
xor U10320 (N_10320,N_10248,N_10215);
and U10321 (N_10321,N_10131,N_10166);
and U10322 (N_10322,N_10183,N_10161);
nand U10323 (N_10323,N_10138,N_10152);
xnor U10324 (N_10324,N_10219,N_10197);
xor U10325 (N_10325,N_10141,N_10148);
and U10326 (N_10326,N_10201,N_10143);
xnor U10327 (N_10327,N_10205,N_10176);
or U10328 (N_10328,N_10169,N_10208);
nand U10329 (N_10329,N_10138,N_10141);
nand U10330 (N_10330,N_10186,N_10192);
nand U10331 (N_10331,N_10153,N_10129);
or U10332 (N_10332,N_10200,N_10125);
nand U10333 (N_10333,N_10142,N_10184);
and U10334 (N_10334,N_10206,N_10170);
and U10335 (N_10335,N_10215,N_10237);
nand U10336 (N_10336,N_10136,N_10139);
nor U10337 (N_10337,N_10232,N_10192);
nand U10338 (N_10338,N_10188,N_10126);
nor U10339 (N_10339,N_10134,N_10230);
nand U10340 (N_10340,N_10146,N_10235);
nand U10341 (N_10341,N_10189,N_10232);
nor U10342 (N_10342,N_10235,N_10187);
xnor U10343 (N_10343,N_10163,N_10189);
and U10344 (N_10344,N_10137,N_10183);
nor U10345 (N_10345,N_10185,N_10243);
and U10346 (N_10346,N_10179,N_10152);
nand U10347 (N_10347,N_10247,N_10185);
nor U10348 (N_10348,N_10209,N_10169);
or U10349 (N_10349,N_10141,N_10242);
and U10350 (N_10350,N_10193,N_10206);
or U10351 (N_10351,N_10202,N_10221);
xnor U10352 (N_10352,N_10126,N_10144);
or U10353 (N_10353,N_10182,N_10210);
xnor U10354 (N_10354,N_10164,N_10208);
nor U10355 (N_10355,N_10132,N_10206);
and U10356 (N_10356,N_10168,N_10216);
nor U10357 (N_10357,N_10204,N_10131);
nand U10358 (N_10358,N_10224,N_10169);
and U10359 (N_10359,N_10185,N_10144);
and U10360 (N_10360,N_10138,N_10234);
nor U10361 (N_10361,N_10238,N_10126);
and U10362 (N_10362,N_10201,N_10135);
xor U10363 (N_10363,N_10130,N_10210);
and U10364 (N_10364,N_10229,N_10174);
or U10365 (N_10365,N_10172,N_10142);
xnor U10366 (N_10366,N_10219,N_10189);
or U10367 (N_10367,N_10235,N_10246);
nand U10368 (N_10368,N_10248,N_10198);
or U10369 (N_10369,N_10218,N_10199);
or U10370 (N_10370,N_10203,N_10197);
nand U10371 (N_10371,N_10227,N_10198);
nor U10372 (N_10372,N_10182,N_10192);
or U10373 (N_10373,N_10137,N_10136);
xor U10374 (N_10374,N_10162,N_10146);
or U10375 (N_10375,N_10308,N_10341);
and U10376 (N_10376,N_10344,N_10329);
or U10377 (N_10377,N_10260,N_10300);
and U10378 (N_10378,N_10320,N_10343);
and U10379 (N_10379,N_10254,N_10351);
and U10380 (N_10380,N_10301,N_10258);
xnor U10381 (N_10381,N_10285,N_10257);
and U10382 (N_10382,N_10337,N_10290);
xnor U10383 (N_10383,N_10342,N_10347);
or U10384 (N_10384,N_10269,N_10263);
or U10385 (N_10385,N_10360,N_10339);
xor U10386 (N_10386,N_10302,N_10270);
or U10387 (N_10387,N_10370,N_10322);
nand U10388 (N_10388,N_10371,N_10330);
nor U10389 (N_10389,N_10373,N_10304);
nor U10390 (N_10390,N_10352,N_10282);
nand U10391 (N_10391,N_10357,N_10296);
nor U10392 (N_10392,N_10338,N_10303);
and U10393 (N_10393,N_10275,N_10350);
xnor U10394 (N_10394,N_10334,N_10250);
nand U10395 (N_10395,N_10312,N_10264);
xnor U10396 (N_10396,N_10331,N_10255);
or U10397 (N_10397,N_10278,N_10326);
and U10398 (N_10398,N_10368,N_10372);
xor U10399 (N_10399,N_10292,N_10333);
xnor U10400 (N_10400,N_10356,N_10365);
or U10401 (N_10401,N_10299,N_10253);
nor U10402 (N_10402,N_10354,N_10362);
and U10403 (N_10403,N_10319,N_10324);
xnor U10404 (N_10404,N_10318,N_10369);
nor U10405 (N_10405,N_10294,N_10361);
nand U10406 (N_10406,N_10374,N_10297);
nand U10407 (N_10407,N_10267,N_10272);
nand U10408 (N_10408,N_10295,N_10281);
nor U10409 (N_10409,N_10277,N_10313);
and U10410 (N_10410,N_10358,N_10328);
nor U10411 (N_10411,N_10307,N_10321);
xnor U10412 (N_10412,N_10314,N_10348);
or U10413 (N_10413,N_10327,N_10349);
nor U10414 (N_10414,N_10364,N_10274);
xnor U10415 (N_10415,N_10305,N_10265);
and U10416 (N_10416,N_10268,N_10309);
nor U10417 (N_10417,N_10359,N_10283);
nor U10418 (N_10418,N_10286,N_10261);
xor U10419 (N_10419,N_10353,N_10355);
xor U10420 (N_10420,N_10266,N_10311);
and U10421 (N_10421,N_10288,N_10315);
xor U10422 (N_10422,N_10289,N_10332);
nand U10423 (N_10423,N_10256,N_10345);
nor U10424 (N_10424,N_10335,N_10340);
nand U10425 (N_10425,N_10310,N_10323);
nor U10426 (N_10426,N_10252,N_10276);
nand U10427 (N_10427,N_10306,N_10325);
nor U10428 (N_10428,N_10363,N_10316);
and U10429 (N_10429,N_10284,N_10367);
and U10430 (N_10430,N_10336,N_10366);
and U10431 (N_10431,N_10273,N_10262);
nand U10432 (N_10432,N_10346,N_10280);
nand U10433 (N_10433,N_10251,N_10259);
and U10434 (N_10434,N_10298,N_10317);
or U10435 (N_10435,N_10287,N_10293);
xnor U10436 (N_10436,N_10291,N_10271);
nand U10437 (N_10437,N_10279,N_10296);
and U10438 (N_10438,N_10358,N_10332);
and U10439 (N_10439,N_10296,N_10359);
xor U10440 (N_10440,N_10372,N_10340);
or U10441 (N_10441,N_10286,N_10346);
xnor U10442 (N_10442,N_10338,N_10366);
or U10443 (N_10443,N_10314,N_10253);
and U10444 (N_10444,N_10310,N_10251);
xnor U10445 (N_10445,N_10372,N_10285);
and U10446 (N_10446,N_10266,N_10351);
nor U10447 (N_10447,N_10272,N_10260);
and U10448 (N_10448,N_10312,N_10325);
and U10449 (N_10449,N_10287,N_10252);
nor U10450 (N_10450,N_10311,N_10341);
or U10451 (N_10451,N_10371,N_10333);
nor U10452 (N_10452,N_10286,N_10308);
nand U10453 (N_10453,N_10270,N_10288);
xor U10454 (N_10454,N_10261,N_10328);
or U10455 (N_10455,N_10280,N_10301);
or U10456 (N_10456,N_10296,N_10346);
nand U10457 (N_10457,N_10310,N_10294);
xor U10458 (N_10458,N_10371,N_10343);
nand U10459 (N_10459,N_10336,N_10296);
xnor U10460 (N_10460,N_10296,N_10307);
nor U10461 (N_10461,N_10370,N_10277);
xnor U10462 (N_10462,N_10251,N_10372);
xnor U10463 (N_10463,N_10324,N_10368);
and U10464 (N_10464,N_10337,N_10315);
nor U10465 (N_10465,N_10257,N_10289);
nor U10466 (N_10466,N_10350,N_10264);
xor U10467 (N_10467,N_10343,N_10369);
xnor U10468 (N_10468,N_10316,N_10276);
and U10469 (N_10469,N_10275,N_10320);
and U10470 (N_10470,N_10323,N_10345);
and U10471 (N_10471,N_10324,N_10254);
xor U10472 (N_10472,N_10256,N_10281);
and U10473 (N_10473,N_10274,N_10356);
or U10474 (N_10474,N_10347,N_10293);
or U10475 (N_10475,N_10281,N_10282);
nor U10476 (N_10476,N_10276,N_10317);
xor U10477 (N_10477,N_10285,N_10291);
and U10478 (N_10478,N_10260,N_10355);
and U10479 (N_10479,N_10371,N_10315);
and U10480 (N_10480,N_10284,N_10317);
xor U10481 (N_10481,N_10338,N_10319);
nor U10482 (N_10482,N_10285,N_10269);
and U10483 (N_10483,N_10256,N_10323);
and U10484 (N_10484,N_10308,N_10326);
or U10485 (N_10485,N_10254,N_10300);
nand U10486 (N_10486,N_10301,N_10286);
and U10487 (N_10487,N_10352,N_10283);
xnor U10488 (N_10488,N_10325,N_10343);
xor U10489 (N_10489,N_10285,N_10276);
and U10490 (N_10490,N_10362,N_10324);
xor U10491 (N_10491,N_10251,N_10334);
and U10492 (N_10492,N_10291,N_10342);
or U10493 (N_10493,N_10262,N_10370);
xnor U10494 (N_10494,N_10250,N_10291);
or U10495 (N_10495,N_10312,N_10348);
or U10496 (N_10496,N_10370,N_10260);
or U10497 (N_10497,N_10349,N_10264);
xor U10498 (N_10498,N_10345,N_10348);
nor U10499 (N_10499,N_10293,N_10256);
xor U10500 (N_10500,N_10422,N_10487);
or U10501 (N_10501,N_10489,N_10468);
and U10502 (N_10502,N_10389,N_10483);
or U10503 (N_10503,N_10382,N_10467);
nand U10504 (N_10504,N_10490,N_10499);
nand U10505 (N_10505,N_10396,N_10376);
nand U10506 (N_10506,N_10415,N_10469);
nand U10507 (N_10507,N_10416,N_10493);
and U10508 (N_10508,N_10436,N_10413);
xor U10509 (N_10509,N_10399,N_10401);
or U10510 (N_10510,N_10461,N_10404);
and U10511 (N_10511,N_10482,N_10494);
xnor U10512 (N_10512,N_10395,N_10486);
nand U10513 (N_10513,N_10429,N_10443);
or U10514 (N_10514,N_10492,N_10440);
or U10515 (N_10515,N_10423,N_10479);
nor U10516 (N_10516,N_10427,N_10420);
nor U10517 (N_10517,N_10466,N_10442);
nor U10518 (N_10518,N_10475,N_10459);
nand U10519 (N_10519,N_10383,N_10380);
and U10520 (N_10520,N_10477,N_10497);
nand U10521 (N_10521,N_10484,N_10438);
and U10522 (N_10522,N_10447,N_10428);
nor U10523 (N_10523,N_10397,N_10394);
nor U10524 (N_10524,N_10454,N_10470);
nor U10525 (N_10525,N_10400,N_10412);
or U10526 (N_10526,N_10462,N_10439);
nor U10527 (N_10527,N_10455,N_10456);
or U10528 (N_10528,N_10418,N_10476);
nand U10529 (N_10529,N_10391,N_10451);
nor U10530 (N_10530,N_10426,N_10402);
nand U10531 (N_10531,N_10444,N_10452);
or U10532 (N_10532,N_10481,N_10417);
nor U10533 (N_10533,N_10387,N_10424);
or U10534 (N_10534,N_10425,N_10464);
nor U10535 (N_10535,N_10495,N_10448);
nor U10536 (N_10536,N_10421,N_10378);
or U10537 (N_10537,N_10431,N_10449);
nand U10538 (N_10538,N_10407,N_10433);
nand U10539 (N_10539,N_10460,N_10390);
xnor U10540 (N_10540,N_10480,N_10435);
and U10541 (N_10541,N_10450,N_10472);
xnor U10542 (N_10542,N_10408,N_10379);
and U10543 (N_10543,N_10414,N_10441);
or U10544 (N_10544,N_10485,N_10381);
and U10545 (N_10545,N_10406,N_10445);
nand U10546 (N_10546,N_10405,N_10388);
and U10547 (N_10547,N_10385,N_10419);
nor U10548 (N_10548,N_10403,N_10446);
xnor U10549 (N_10549,N_10457,N_10465);
or U10550 (N_10550,N_10434,N_10411);
nor U10551 (N_10551,N_10432,N_10409);
xnor U10552 (N_10552,N_10398,N_10471);
xor U10553 (N_10553,N_10473,N_10393);
xor U10554 (N_10554,N_10496,N_10488);
or U10555 (N_10555,N_10384,N_10386);
xor U10556 (N_10556,N_10498,N_10478);
nor U10557 (N_10557,N_10430,N_10463);
xnor U10558 (N_10558,N_10474,N_10375);
nor U10559 (N_10559,N_10377,N_10410);
or U10560 (N_10560,N_10458,N_10491);
or U10561 (N_10561,N_10453,N_10437);
xor U10562 (N_10562,N_10392,N_10464);
nor U10563 (N_10563,N_10434,N_10461);
or U10564 (N_10564,N_10468,N_10477);
or U10565 (N_10565,N_10426,N_10463);
or U10566 (N_10566,N_10444,N_10461);
nand U10567 (N_10567,N_10479,N_10409);
or U10568 (N_10568,N_10413,N_10405);
or U10569 (N_10569,N_10396,N_10438);
and U10570 (N_10570,N_10399,N_10485);
nor U10571 (N_10571,N_10408,N_10407);
nand U10572 (N_10572,N_10391,N_10377);
xor U10573 (N_10573,N_10393,N_10440);
and U10574 (N_10574,N_10448,N_10480);
or U10575 (N_10575,N_10414,N_10406);
xor U10576 (N_10576,N_10472,N_10493);
xor U10577 (N_10577,N_10398,N_10385);
and U10578 (N_10578,N_10461,N_10483);
nor U10579 (N_10579,N_10473,N_10489);
nor U10580 (N_10580,N_10456,N_10398);
or U10581 (N_10581,N_10438,N_10436);
xnor U10582 (N_10582,N_10384,N_10434);
xor U10583 (N_10583,N_10470,N_10445);
or U10584 (N_10584,N_10440,N_10381);
nor U10585 (N_10585,N_10470,N_10438);
and U10586 (N_10586,N_10412,N_10462);
nor U10587 (N_10587,N_10490,N_10482);
nor U10588 (N_10588,N_10450,N_10393);
and U10589 (N_10589,N_10483,N_10445);
and U10590 (N_10590,N_10384,N_10395);
nor U10591 (N_10591,N_10385,N_10486);
or U10592 (N_10592,N_10476,N_10481);
or U10593 (N_10593,N_10493,N_10382);
or U10594 (N_10594,N_10401,N_10443);
and U10595 (N_10595,N_10398,N_10451);
nor U10596 (N_10596,N_10450,N_10391);
or U10597 (N_10597,N_10488,N_10417);
and U10598 (N_10598,N_10437,N_10445);
nand U10599 (N_10599,N_10424,N_10427);
and U10600 (N_10600,N_10391,N_10462);
nand U10601 (N_10601,N_10434,N_10499);
nand U10602 (N_10602,N_10396,N_10385);
or U10603 (N_10603,N_10475,N_10430);
nand U10604 (N_10604,N_10401,N_10490);
xnor U10605 (N_10605,N_10451,N_10408);
nand U10606 (N_10606,N_10482,N_10441);
or U10607 (N_10607,N_10464,N_10375);
nor U10608 (N_10608,N_10492,N_10444);
xnor U10609 (N_10609,N_10469,N_10375);
or U10610 (N_10610,N_10394,N_10491);
and U10611 (N_10611,N_10437,N_10432);
or U10612 (N_10612,N_10451,N_10449);
or U10613 (N_10613,N_10445,N_10458);
nand U10614 (N_10614,N_10483,N_10479);
and U10615 (N_10615,N_10380,N_10423);
nand U10616 (N_10616,N_10403,N_10483);
and U10617 (N_10617,N_10469,N_10402);
nand U10618 (N_10618,N_10451,N_10413);
nor U10619 (N_10619,N_10379,N_10490);
xor U10620 (N_10620,N_10401,N_10457);
xnor U10621 (N_10621,N_10468,N_10469);
or U10622 (N_10622,N_10491,N_10418);
xor U10623 (N_10623,N_10456,N_10402);
nand U10624 (N_10624,N_10496,N_10381);
nor U10625 (N_10625,N_10605,N_10586);
nor U10626 (N_10626,N_10523,N_10579);
nor U10627 (N_10627,N_10584,N_10509);
nand U10628 (N_10628,N_10610,N_10532);
xor U10629 (N_10629,N_10594,N_10531);
or U10630 (N_10630,N_10576,N_10524);
nor U10631 (N_10631,N_10540,N_10609);
xor U10632 (N_10632,N_10599,N_10504);
nand U10633 (N_10633,N_10511,N_10596);
nor U10634 (N_10634,N_10590,N_10530);
nor U10635 (N_10635,N_10578,N_10541);
nand U10636 (N_10636,N_10622,N_10613);
nand U10637 (N_10637,N_10595,N_10607);
nor U10638 (N_10638,N_10542,N_10544);
nor U10639 (N_10639,N_10569,N_10601);
nand U10640 (N_10640,N_10589,N_10620);
and U10641 (N_10641,N_10554,N_10562);
nand U10642 (N_10642,N_10552,N_10551);
or U10643 (N_10643,N_10533,N_10571);
xor U10644 (N_10644,N_10518,N_10557);
nand U10645 (N_10645,N_10508,N_10565);
xnor U10646 (N_10646,N_10560,N_10500);
nor U10647 (N_10647,N_10514,N_10520);
or U10648 (N_10648,N_10612,N_10618);
or U10649 (N_10649,N_10570,N_10505);
and U10650 (N_10650,N_10507,N_10623);
nand U10651 (N_10651,N_10563,N_10545);
nand U10652 (N_10652,N_10585,N_10591);
xnor U10653 (N_10653,N_10539,N_10602);
nor U10654 (N_10654,N_10502,N_10575);
nor U10655 (N_10655,N_10501,N_10567);
nand U10656 (N_10656,N_10566,N_10503);
nor U10657 (N_10657,N_10573,N_10598);
and U10658 (N_10658,N_10521,N_10546);
or U10659 (N_10659,N_10534,N_10538);
nand U10660 (N_10660,N_10522,N_10572);
and U10661 (N_10661,N_10614,N_10597);
nand U10662 (N_10662,N_10537,N_10543);
nor U10663 (N_10663,N_10624,N_10561);
nor U10664 (N_10664,N_10529,N_10515);
and U10665 (N_10665,N_10582,N_10600);
xor U10666 (N_10666,N_10587,N_10525);
nand U10667 (N_10667,N_10621,N_10608);
nor U10668 (N_10668,N_10512,N_10588);
or U10669 (N_10669,N_10580,N_10535);
or U10670 (N_10670,N_10611,N_10593);
xnor U10671 (N_10671,N_10516,N_10559);
or U10672 (N_10672,N_10581,N_10619);
and U10673 (N_10673,N_10549,N_10506);
nor U10674 (N_10674,N_10517,N_10577);
xor U10675 (N_10675,N_10616,N_10564);
xnor U10676 (N_10676,N_10513,N_10615);
nor U10677 (N_10677,N_10527,N_10604);
nor U10678 (N_10678,N_10553,N_10526);
nand U10679 (N_10679,N_10550,N_10583);
xnor U10680 (N_10680,N_10592,N_10558);
nor U10681 (N_10681,N_10528,N_10510);
and U10682 (N_10682,N_10574,N_10547);
nor U10683 (N_10683,N_10536,N_10603);
nand U10684 (N_10684,N_10519,N_10617);
or U10685 (N_10685,N_10556,N_10606);
xor U10686 (N_10686,N_10548,N_10555);
nand U10687 (N_10687,N_10568,N_10591);
nand U10688 (N_10688,N_10620,N_10504);
nor U10689 (N_10689,N_10526,N_10587);
nor U10690 (N_10690,N_10614,N_10610);
or U10691 (N_10691,N_10578,N_10616);
and U10692 (N_10692,N_10622,N_10579);
nand U10693 (N_10693,N_10621,N_10524);
and U10694 (N_10694,N_10590,N_10578);
or U10695 (N_10695,N_10599,N_10524);
and U10696 (N_10696,N_10554,N_10587);
or U10697 (N_10697,N_10538,N_10589);
and U10698 (N_10698,N_10596,N_10577);
nor U10699 (N_10699,N_10532,N_10618);
and U10700 (N_10700,N_10549,N_10551);
or U10701 (N_10701,N_10606,N_10620);
and U10702 (N_10702,N_10619,N_10587);
xnor U10703 (N_10703,N_10538,N_10605);
or U10704 (N_10704,N_10500,N_10553);
or U10705 (N_10705,N_10557,N_10602);
or U10706 (N_10706,N_10591,N_10556);
and U10707 (N_10707,N_10586,N_10516);
xor U10708 (N_10708,N_10523,N_10534);
nor U10709 (N_10709,N_10585,N_10547);
and U10710 (N_10710,N_10543,N_10511);
nand U10711 (N_10711,N_10506,N_10520);
xnor U10712 (N_10712,N_10526,N_10606);
nand U10713 (N_10713,N_10612,N_10518);
xnor U10714 (N_10714,N_10608,N_10502);
nor U10715 (N_10715,N_10516,N_10533);
and U10716 (N_10716,N_10509,N_10617);
or U10717 (N_10717,N_10589,N_10614);
nor U10718 (N_10718,N_10571,N_10623);
nor U10719 (N_10719,N_10591,N_10617);
nand U10720 (N_10720,N_10574,N_10617);
and U10721 (N_10721,N_10607,N_10500);
nand U10722 (N_10722,N_10508,N_10578);
and U10723 (N_10723,N_10621,N_10559);
nor U10724 (N_10724,N_10503,N_10516);
nor U10725 (N_10725,N_10558,N_10595);
nand U10726 (N_10726,N_10607,N_10549);
nand U10727 (N_10727,N_10510,N_10558);
nor U10728 (N_10728,N_10568,N_10575);
xor U10729 (N_10729,N_10554,N_10611);
or U10730 (N_10730,N_10615,N_10621);
and U10731 (N_10731,N_10568,N_10540);
and U10732 (N_10732,N_10532,N_10543);
and U10733 (N_10733,N_10523,N_10535);
xor U10734 (N_10734,N_10518,N_10601);
and U10735 (N_10735,N_10513,N_10523);
or U10736 (N_10736,N_10529,N_10623);
nand U10737 (N_10737,N_10621,N_10587);
nand U10738 (N_10738,N_10507,N_10593);
or U10739 (N_10739,N_10521,N_10543);
nor U10740 (N_10740,N_10565,N_10546);
and U10741 (N_10741,N_10524,N_10587);
nor U10742 (N_10742,N_10623,N_10611);
and U10743 (N_10743,N_10623,N_10533);
and U10744 (N_10744,N_10549,N_10555);
nand U10745 (N_10745,N_10514,N_10623);
nor U10746 (N_10746,N_10509,N_10585);
nand U10747 (N_10747,N_10529,N_10555);
or U10748 (N_10748,N_10608,N_10542);
nor U10749 (N_10749,N_10599,N_10567);
nand U10750 (N_10750,N_10738,N_10657);
xor U10751 (N_10751,N_10641,N_10704);
nand U10752 (N_10752,N_10683,N_10733);
nand U10753 (N_10753,N_10659,N_10690);
xor U10754 (N_10754,N_10697,N_10742);
nor U10755 (N_10755,N_10743,N_10667);
xnor U10756 (N_10756,N_10652,N_10675);
and U10757 (N_10757,N_10746,N_10722);
or U10758 (N_10758,N_10707,N_10650);
or U10759 (N_10759,N_10672,N_10747);
xor U10760 (N_10760,N_10735,N_10721);
xor U10761 (N_10761,N_10705,N_10674);
nor U10762 (N_10762,N_10635,N_10646);
and U10763 (N_10763,N_10693,N_10682);
nand U10764 (N_10764,N_10698,N_10744);
or U10765 (N_10765,N_10627,N_10739);
nand U10766 (N_10766,N_10655,N_10666);
nor U10767 (N_10767,N_10661,N_10632);
xor U10768 (N_10768,N_10636,N_10731);
xor U10769 (N_10769,N_10685,N_10718);
nor U10770 (N_10770,N_10708,N_10729);
xor U10771 (N_10771,N_10649,N_10668);
or U10772 (N_10772,N_10681,N_10732);
or U10773 (N_10773,N_10687,N_10651);
xnor U10774 (N_10774,N_10692,N_10737);
or U10775 (N_10775,N_10660,N_10699);
xor U10776 (N_10776,N_10656,N_10630);
nor U10777 (N_10777,N_10740,N_10691);
and U10778 (N_10778,N_10736,N_10724);
and U10779 (N_10779,N_10702,N_10639);
nand U10780 (N_10780,N_10679,N_10665);
nand U10781 (N_10781,N_10727,N_10748);
and U10782 (N_10782,N_10716,N_10714);
or U10783 (N_10783,N_10648,N_10701);
and U10784 (N_10784,N_10680,N_10642);
nor U10785 (N_10785,N_10717,N_10684);
nor U10786 (N_10786,N_10676,N_10663);
or U10787 (N_10787,N_10723,N_10671);
nor U10788 (N_10788,N_10749,N_10670);
and U10789 (N_10789,N_10700,N_10695);
nor U10790 (N_10790,N_10734,N_10633);
xnor U10791 (N_10791,N_10706,N_10625);
xnor U10792 (N_10792,N_10730,N_10741);
nor U10793 (N_10793,N_10710,N_10728);
and U10794 (N_10794,N_10653,N_10678);
and U10795 (N_10795,N_10725,N_10694);
or U10796 (N_10796,N_10688,N_10673);
xnor U10797 (N_10797,N_10689,N_10654);
nor U10798 (N_10798,N_10720,N_10719);
or U10799 (N_10799,N_10712,N_10696);
xor U10800 (N_10800,N_10647,N_10726);
nor U10801 (N_10801,N_10640,N_10643);
nor U10802 (N_10802,N_10629,N_10664);
nor U10803 (N_10803,N_10631,N_10658);
nand U10804 (N_10804,N_10709,N_10715);
nand U10805 (N_10805,N_10669,N_10713);
xnor U10806 (N_10806,N_10626,N_10703);
nor U10807 (N_10807,N_10677,N_10638);
nor U10808 (N_10808,N_10645,N_10711);
nor U10809 (N_10809,N_10628,N_10686);
nor U10810 (N_10810,N_10662,N_10637);
nand U10811 (N_10811,N_10644,N_10745);
nor U10812 (N_10812,N_10634,N_10654);
xnor U10813 (N_10813,N_10701,N_10627);
or U10814 (N_10814,N_10687,N_10675);
nor U10815 (N_10815,N_10631,N_10743);
or U10816 (N_10816,N_10704,N_10660);
and U10817 (N_10817,N_10691,N_10631);
or U10818 (N_10818,N_10745,N_10713);
and U10819 (N_10819,N_10699,N_10659);
or U10820 (N_10820,N_10648,N_10649);
nor U10821 (N_10821,N_10667,N_10725);
nand U10822 (N_10822,N_10653,N_10676);
nand U10823 (N_10823,N_10736,N_10633);
nand U10824 (N_10824,N_10654,N_10747);
and U10825 (N_10825,N_10710,N_10694);
xnor U10826 (N_10826,N_10709,N_10731);
nor U10827 (N_10827,N_10679,N_10712);
nor U10828 (N_10828,N_10648,N_10708);
xnor U10829 (N_10829,N_10732,N_10740);
or U10830 (N_10830,N_10680,N_10659);
nor U10831 (N_10831,N_10638,N_10668);
xor U10832 (N_10832,N_10655,N_10693);
or U10833 (N_10833,N_10682,N_10706);
nor U10834 (N_10834,N_10661,N_10738);
xor U10835 (N_10835,N_10658,N_10718);
nand U10836 (N_10836,N_10659,N_10716);
and U10837 (N_10837,N_10658,N_10724);
xnor U10838 (N_10838,N_10634,N_10637);
or U10839 (N_10839,N_10676,N_10660);
xor U10840 (N_10840,N_10674,N_10688);
and U10841 (N_10841,N_10740,N_10661);
xnor U10842 (N_10842,N_10737,N_10641);
and U10843 (N_10843,N_10728,N_10640);
or U10844 (N_10844,N_10737,N_10721);
xnor U10845 (N_10845,N_10675,N_10685);
xor U10846 (N_10846,N_10638,N_10713);
nor U10847 (N_10847,N_10660,N_10657);
nor U10848 (N_10848,N_10704,N_10642);
nand U10849 (N_10849,N_10647,N_10701);
and U10850 (N_10850,N_10686,N_10627);
nand U10851 (N_10851,N_10686,N_10669);
or U10852 (N_10852,N_10716,N_10637);
and U10853 (N_10853,N_10735,N_10647);
and U10854 (N_10854,N_10668,N_10726);
and U10855 (N_10855,N_10638,N_10669);
nor U10856 (N_10856,N_10730,N_10721);
and U10857 (N_10857,N_10730,N_10678);
or U10858 (N_10858,N_10689,N_10671);
or U10859 (N_10859,N_10639,N_10714);
or U10860 (N_10860,N_10729,N_10715);
nor U10861 (N_10861,N_10714,N_10738);
nand U10862 (N_10862,N_10676,N_10703);
xor U10863 (N_10863,N_10693,N_10672);
xnor U10864 (N_10864,N_10738,N_10727);
nand U10865 (N_10865,N_10703,N_10672);
or U10866 (N_10866,N_10627,N_10704);
xor U10867 (N_10867,N_10638,N_10699);
nor U10868 (N_10868,N_10677,N_10647);
xor U10869 (N_10869,N_10717,N_10676);
nand U10870 (N_10870,N_10653,N_10662);
xor U10871 (N_10871,N_10655,N_10653);
or U10872 (N_10872,N_10625,N_10714);
xnor U10873 (N_10873,N_10652,N_10644);
nor U10874 (N_10874,N_10749,N_10715);
or U10875 (N_10875,N_10801,N_10872);
nor U10876 (N_10876,N_10820,N_10813);
nor U10877 (N_10877,N_10808,N_10812);
nand U10878 (N_10878,N_10818,N_10874);
xor U10879 (N_10879,N_10853,N_10854);
or U10880 (N_10880,N_10759,N_10857);
nor U10881 (N_10881,N_10868,N_10772);
or U10882 (N_10882,N_10774,N_10842);
and U10883 (N_10883,N_10758,N_10779);
nand U10884 (N_10884,N_10841,N_10787);
xnor U10885 (N_10885,N_10834,N_10753);
or U10886 (N_10886,N_10786,N_10762);
nand U10887 (N_10887,N_10836,N_10838);
nand U10888 (N_10888,N_10837,N_10798);
xnor U10889 (N_10889,N_10821,N_10784);
and U10890 (N_10890,N_10816,N_10822);
or U10891 (N_10891,N_10800,N_10832);
nor U10892 (N_10892,N_10783,N_10797);
and U10893 (N_10893,N_10756,N_10809);
nor U10894 (N_10894,N_10827,N_10869);
and U10895 (N_10895,N_10811,N_10829);
nand U10896 (N_10896,N_10755,N_10850);
nor U10897 (N_10897,N_10764,N_10830);
and U10898 (N_10898,N_10839,N_10771);
xnor U10899 (N_10899,N_10776,N_10871);
or U10900 (N_10900,N_10828,N_10794);
or U10901 (N_10901,N_10819,N_10824);
and U10902 (N_10902,N_10856,N_10752);
and U10903 (N_10903,N_10826,N_10806);
xor U10904 (N_10904,N_10840,N_10845);
xnor U10905 (N_10905,N_10867,N_10788);
nor U10906 (N_10906,N_10817,N_10852);
or U10907 (N_10907,N_10763,N_10803);
nand U10908 (N_10908,N_10792,N_10810);
nor U10909 (N_10909,N_10780,N_10751);
nor U10910 (N_10910,N_10860,N_10793);
nand U10911 (N_10911,N_10757,N_10844);
or U10912 (N_10912,N_10777,N_10862);
nor U10913 (N_10913,N_10835,N_10859);
xor U10914 (N_10914,N_10768,N_10781);
and U10915 (N_10915,N_10760,N_10831);
and U10916 (N_10916,N_10790,N_10823);
xnor U10917 (N_10917,N_10848,N_10769);
and U10918 (N_10918,N_10846,N_10866);
and U10919 (N_10919,N_10847,N_10778);
nor U10920 (N_10920,N_10864,N_10796);
or U10921 (N_10921,N_10773,N_10785);
nand U10922 (N_10922,N_10807,N_10770);
xor U10923 (N_10923,N_10766,N_10802);
or U10924 (N_10924,N_10814,N_10870);
or U10925 (N_10925,N_10849,N_10865);
or U10926 (N_10926,N_10782,N_10833);
nor U10927 (N_10927,N_10795,N_10804);
xor U10928 (N_10928,N_10815,N_10789);
xnor U10929 (N_10929,N_10799,N_10825);
and U10930 (N_10930,N_10858,N_10843);
or U10931 (N_10931,N_10754,N_10765);
and U10932 (N_10932,N_10775,N_10863);
nand U10933 (N_10933,N_10767,N_10855);
xor U10934 (N_10934,N_10805,N_10873);
nor U10935 (N_10935,N_10761,N_10750);
and U10936 (N_10936,N_10861,N_10791);
xor U10937 (N_10937,N_10851,N_10846);
and U10938 (N_10938,N_10778,N_10773);
nor U10939 (N_10939,N_10802,N_10863);
and U10940 (N_10940,N_10856,N_10751);
xnor U10941 (N_10941,N_10847,N_10850);
nor U10942 (N_10942,N_10767,N_10795);
nor U10943 (N_10943,N_10826,N_10797);
or U10944 (N_10944,N_10750,N_10837);
nand U10945 (N_10945,N_10830,N_10783);
or U10946 (N_10946,N_10858,N_10769);
xor U10947 (N_10947,N_10827,N_10757);
nand U10948 (N_10948,N_10757,N_10862);
xor U10949 (N_10949,N_10863,N_10856);
or U10950 (N_10950,N_10801,N_10856);
nor U10951 (N_10951,N_10756,N_10823);
nand U10952 (N_10952,N_10872,N_10823);
or U10953 (N_10953,N_10820,N_10840);
nor U10954 (N_10954,N_10798,N_10785);
and U10955 (N_10955,N_10839,N_10856);
nor U10956 (N_10956,N_10822,N_10859);
or U10957 (N_10957,N_10841,N_10828);
nor U10958 (N_10958,N_10779,N_10756);
and U10959 (N_10959,N_10801,N_10765);
and U10960 (N_10960,N_10784,N_10847);
and U10961 (N_10961,N_10844,N_10851);
or U10962 (N_10962,N_10865,N_10835);
nor U10963 (N_10963,N_10860,N_10753);
nand U10964 (N_10964,N_10779,N_10761);
or U10965 (N_10965,N_10871,N_10805);
and U10966 (N_10966,N_10808,N_10769);
xnor U10967 (N_10967,N_10755,N_10861);
nand U10968 (N_10968,N_10775,N_10868);
nand U10969 (N_10969,N_10757,N_10871);
nand U10970 (N_10970,N_10829,N_10775);
or U10971 (N_10971,N_10802,N_10874);
nor U10972 (N_10972,N_10765,N_10874);
xnor U10973 (N_10973,N_10799,N_10807);
xor U10974 (N_10974,N_10864,N_10840);
nand U10975 (N_10975,N_10810,N_10839);
and U10976 (N_10976,N_10752,N_10842);
or U10977 (N_10977,N_10769,N_10822);
and U10978 (N_10978,N_10766,N_10799);
and U10979 (N_10979,N_10768,N_10804);
nand U10980 (N_10980,N_10842,N_10785);
nor U10981 (N_10981,N_10829,N_10796);
xor U10982 (N_10982,N_10798,N_10787);
nand U10983 (N_10983,N_10824,N_10809);
or U10984 (N_10984,N_10815,N_10760);
nand U10985 (N_10985,N_10812,N_10782);
or U10986 (N_10986,N_10781,N_10842);
nor U10987 (N_10987,N_10769,N_10821);
xor U10988 (N_10988,N_10874,N_10799);
or U10989 (N_10989,N_10870,N_10864);
and U10990 (N_10990,N_10778,N_10856);
nor U10991 (N_10991,N_10864,N_10861);
or U10992 (N_10992,N_10779,N_10817);
xnor U10993 (N_10993,N_10815,N_10761);
xnor U10994 (N_10994,N_10776,N_10765);
nand U10995 (N_10995,N_10866,N_10785);
and U10996 (N_10996,N_10852,N_10803);
nor U10997 (N_10997,N_10871,N_10771);
and U10998 (N_10998,N_10873,N_10788);
and U10999 (N_10999,N_10864,N_10818);
xnor U11000 (N_11000,N_10954,N_10950);
nor U11001 (N_11001,N_10889,N_10922);
xnor U11002 (N_11002,N_10919,N_10916);
and U11003 (N_11003,N_10939,N_10938);
xnor U11004 (N_11004,N_10957,N_10942);
nor U11005 (N_11005,N_10990,N_10935);
and U11006 (N_11006,N_10996,N_10960);
and U11007 (N_11007,N_10876,N_10886);
nand U11008 (N_11008,N_10902,N_10893);
and U11009 (N_11009,N_10884,N_10968);
nor U11010 (N_11010,N_10965,N_10944);
xor U11011 (N_11011,N_10878,N_10976);
and U11012 (N_11012,N_10953,N_10991);
and U11013 (N_11013,N_10897,N_10914);
or U11014 (N_11014,N_10988,N_10956);
and U11015 (N_11015,N_10894,N_10891);
and U11016 (N_11016,N_10959,N_10929);
xnor U11017 (N_11017,N_10906,N_10995);
xnor U11018 (N_11018,N_10971,N_10955);
nor U11019 (N_11019,N_10994,N_10920);
nor U11020 (N_11020,N_10973,N_10948);
nand U11021 (N_11021,N_10963,N_10877);
or U11022 (N_11022,N_10977,N_10993);
and U11023 (N_11023,N_10961,N_10909);
and U11024 (N_11024,N_10964,N_10951);
or U11025 (N_11025,N_10901,N_10937);
nor U11026 (N_11026,N_10905,N_10892);
and U11027 (N_11027,N_10925,N_10875);
and U11028 (N_11028,N_10984,N_10883);
nor U11029 (N_11029,N_10927,N_10900);
xnor U11030 (N_11030,N_10898,N_10992);
xnor U11031 (N_11031,N_10928,N_10969);
nor U11032 (N_11032,N_10903,N_10911);
xnor U11033 (N_11033,N_10941,N_10931);
xor U11034 (N_11034,N_10908,N_10936);
xnor U11035 (N_11035,N_10983,N_10943);
and U11036 (N_11036,N_10932,N_10921);
or U11037 (N_11037,N_10989,N_10924);
xor U11038 (N_11038,N_10958,N_10879);
nor U11039 (N_11039,N_10888,N_10975);
nor U11040 (N_11040,N_10952,N_10885);
or U11041 (N_11041,N_10918,N_10910);
nor U11042 (N_11042,N_10946,N_10895);
or U11043 (N_11043,N_10947,N_10896);
nand U11044 (N_11044,N_10912,N_10987);
xnor U11045 (N_11045,N_10999,N_10967);
and U11046 (N_11046,N_10979,N_10982);
or U11047 (N_11047,N_10899,N_10945);
or U11048 (N_11048,N_10981,N_10907);
and U11049 (N_11049,N_10986,N_10940);
nor U11050 (N_11050,N_10887,N_10985);
nor U11051 (N_11051,N_10890,N_10998);
xor U11052 (N_11052,N_10933,N_10997);
nor U11053 (N_11053,N_10881,N_10882);
nor U11054 (N_11054,N_10923,N_10962);
xnor U11055 (N_11055,N_10930,N_10974);
and U11056 (N_11056,N_10966,N_10917);
or U11057 (N_11057,N_10972,N_10980);
nand U11058 (N_11058,N_10880,N_10913);
nor U11059 (N_11059,N_10978,N_10934);
nor U11060 (N_11060,N_10915,N_10970);
nor U11061 (N_11061,N_10926,N_10904);
nand U11062 (N_11062,N_10949,N_10987);
nand U11063 (N_11063,N_10939,N_10875);
nand U11064 (N_11064,N_10910,N_10933);
or U11065 (N_11065,N_10879,N_10877);
nand U11066 (N_11066,N_10935,N_10988);
xnor U11067 (N_11067,N_10975,N_10987);
nor U11068 (N_11068,N_10961,N_10944);
nand U11069 (N_11069,N_10971,N_10984);
nor U11070 (N_11070,N_10892,N_10891);
nor U11071 (N_11071,N_10895,N_10876);
xnor U11072 (N_11072,N_10928,N_10960);
and U11073 (N_11073,N_10876,N_10981);
or U11074 (N_11074,N_10949,N_10969);
or U11075 (N_11075,N_10915,N_10986);
and U11076 (N_11076,N_10900,N_10986);
xnor U11077 (N_11077,N_10930,N_10969);
nor U11078 (N_11078,N_10892,N_10951);
nor U11079 (N_11079,N_10964,N_10950);
nor U11080 (N_11080,N_10937,N_10910);
and U11081 (N_11081,N_10941,N_10881);
nand U11082 (N_11082,N_10941,N_10961);
nand U11083 (N_11083,N_10925,N_10989);
nand U11084 (N_11084,N_10947,N_10930);
nand U11085 (N_11085,N_10932,N_10929);
nor U11086 (N_11086,N_10941,N_10944);
nor U11087 (N_11087,N_10879,N_10914);
and U11088 (N_11088,N_10901,N_10994);
xor U11089 (N_11089,N_10985,N_10948);
or U11090 (N_11090,N_10893,N_10979);
and U11091 (N_11091,N_10893,N_10958);
or U11092 (N_11092,N_10875,N_10994);
xnor U11093 (N_11093,N_10927,N_10996);
or U11094 (N_11094,N_10976,N_10979);
xnor U11095 (N_11095,N_10973,N_10969);
nand U11096 (N_11096,N_10925,N_10893);
and U11097 (N_11097,N_10896,N_10985);
or U11098 (N_11098,N_10893,N_10940);
nand U11099 (N_11099,N_10970,N_10945);
xnor U11100 (N_11100,N_10916,N_10955);
xor U11101 (N_11101,N_10942,N_10904);
or U11102 (N_11102,N_10944,N_10897);
nor U11103 (N_11103,N_10943,N_10881);
xor U11104 (N_11104,N_10901,N_10987);
nor U11105 (N_11105,N_10925,N_10930);
nand U11106 (N_11106,N_10946,N_10875);
nand U11107 (N_11107,N_10946,N_10905);
nor U11108 (N_11108,N_10951,N_10927);
nand U11109 (N_11109,N_10882,N_10896);
nor U11110 (N_11110,N_10880,N_10937);
nand U11111 (N_11111,N_10936,N_10941);
or U11112 (N_11112,N_10926,N_10942);
xor U11113 (N_11113,N_10993,N_10955);
nor U11114 (N_11114,N_10892,N_10965);
xnor U11115 (N_11115,N_10928,N_10981);
and U11116 (N_11116,N_10933,N_10941);
and U11117 (N_11117,N_10963,N_10959);
nand U11118 (N_11118,N_10930,N_10909);
and U11119 (N_11119,N_10977,N_10916);
xnor U11120 (N_11120,N_10951,N_10985);
or U11121 (N_11121,N_10976,N_10897);
xnor U11122 (N_11122,N_10962,N_10963);
xnor U11123 (N_11123,N_10995,N_10936);
nor U11124 (N_11124,N_10888,N_10996);
and U11125 (N_11125,N_11026,N_11092);
and U11126 (N_11126,N_11043,N_11114);
nor U11127 (N_11127,N_11074,N_11040);
and U11128 (N_11128,N_11022,N_11101);
or U11129 (N_11129,N_11124,N_11091);
nand U11130 (N_11130,N_11003,N_11057);
nand U11131 (N_11131,N_11024,N_11123);
nor U11132 (N_11132,N_11104,N_11117);
xnor U11133 (N_11133,N_11048,N_11113);
nor U11134 (N_11134,N_11058,N_11005);
nor U11135 (N_11135,N_11106,N_11122);
nand U11136 (N_11136,N_11054,N_11021);
xnor U11137 (N_11137,N_11009,N_11050);
and U11138 (N_11138,N_11019,N_11053);
xor U11139 (N_11139,N_11087,N_11051);
nor U11140 (N_11140,N_11018,N_11121);
xnor U11141 (N_11141,N_11011,N_11036);
nor U11142 (N_11142,N_11049,N_11033);
nor U11143 (N_11143,N_11004,N_11072);
or U11144 (N_11144,N_11060,N_11082);
or U11145 (N_11145,N_11037,N_11035);
or U11146 (N_11146,N_11093,N_11067);
and U11147 (N_11147,N_11069,N_11120);
xnor U11148 (N_11148,N_11013,N_11112);
and U11149 (N_11149,N_11062,N_11007);
or U11150 (N_11150,N_11078,N_11002);
xnor U11151 (N_11151,N_11115,N_11025);
xor U11152 (N_11152,N_11094,N_11028);
or U11153 (N_11153,N_11000,N_11032);
and U11154 (N_11154,N_11052,N_11097);
and U11155 (N_11155,N_11096,N_11006);
or U11156 (N_11156,N_11086,N_11073);
nor U11157 (N_11157,N_11055,N_11020);
nand U11158 (N_11158,N_11029,N_11088);
nor U11159 (N_11159,N_11030,N_11061);
xnor U11160 (N_11160,N_11016,N_11059);
xnor U11161 (N_11161,N_11105,N_11014);
nor U11162 (N_11162,N_11118,N_11064);
xnor U11163 (N_11163,N_11023,N_11068);
nand U11164 (N_11164,N_11095,N_11034);
or U11165 (N_11165,N_11100,N_11119);
xnor U11166 (N_11166,N_11010,N_11017);
nor U11167 (N_11167,N_11102,N_11116);
and U11168 (N_11168,N_11045,N_11015);
xor U11169 (N_11169,N_11081,N_11080);
or U11170 (N_11170,N_11012,N_11090);
nand U11171 (N_11171,N_11027,N_11079);
or U11172 (N_11172,N_11108,N_11039);
nand U11173 (N_11173,N_11098,N_11083);
nor U11174 (N_11174,N_11075,N_11056);
xnor U11175 (N_11175,N_11008,N_11046);
xor U11176 (N_11176,N_11110,N_11076);
nor U11177 (N_11177,N_11038,N_11065);
and U11178 (N_11178,N_11109,N_11031);
nor U11179 (N_11179,N_11047,N_11084);
or U11180 (N_11180,N_11085,N_11089);
nand U11181 (N_11181,N_11044,N_11063);
nor U11182 (N_11182,N_11111,N_11099);
nor U11183 (N_11183,N_11103,N_11107);
and U11184 (N_11184,N_11042,N_11071);
and U11185 (N_11185,N_11070,N_11066);
nand U11186 (N_11186,N_11001,N_11041);
xor U11187 (N_11187,N_11077,N_11099);
and U11188 (N_11188,N_11108,N_11093);
or U11189 (N_11189,N_11009,N_11079);
or U11190 (N_11190,N_11059,N_11093);
or U11191 (N_11191,N_11099,N_11119);
nand U11192 (N_11192,N_11109,N_11077);
and U11193 (N_11193,N_11117,N_11026);
or U11194 (N_11194,N_11091,N_11033);
xnor U11195 (N_11195,N_11112,N_11119);
xor U11196 (N_11196,N_11021,N_11016);
xnor U11197 (N_11197,N_11039,N_11109);
nand U11198 (N_11198,N_11095,N_11028);
or U11199 (N_11199,N_11012,N_11061);
nand U11200 (N_11200,N_11002,N_11088);
nand U11201 (N_11201,N_11049,N_11088);
and U11202 (N_11202,N_11097,N_11064);
nand U11203 (N_11203,N_11084,N_11079);
nand U11204 (N_11204,N_11026,N_11024);
and U11205 (N_11205,N_11043,N_11070);
nor U11206 (N_11206,N_11041,N_11030);
nor U11207 (N_11207,N_11088,N_11097);
or U11208 (N_11208,N_11066,N_11033);
nand U11209 (N_11209,N_11049,N_11061);
nand U11210 (N_11210,N_11071,N_11044);
nor U11211 (N_11211,N_11063,N_11111);
xor U11212 (N_11212,N_11011,N_11070);
or U11213 (N_11213,N_11038,N_11006);
nor U11214 (N_11214,N_11026,N_11102);
or U11215 (N_11215,N_11045,N_11009);
nor U11216 (N_11216,N_11119,N_11062);
nand U11217 (N_11217,N_11045,N_11004);
nand U11218 (N_11218,N_11107,N_11047);
nor U11219 (N_11219,N_11059,N_11080);
xor U11220 (N_11220,N_11062,N_11001);
nand U11221 (N_11221,N_11115,N_11060);
nand U11222 (N_11222,N_11057,N_11005);
nor U11223 (N_11223,N_11073,N_11011);
and U11224 (N_11224,N_11068,N_11008);
nor U11225 (N_11225,N_11107,N_11009);
and U11226 (N_11226,N_11058,N_11051);
xnor U11227 (N_11227,N_11107,N_11073);
nand U11228 (N_11228,N_11018,N_11071);
nor U11229 (N_11229,N_11046,N_11082);
nand U11230 (N_11230,N_11097,N_11023);
nor U11231 (N_11231,N_11036,N_11056);
nor U11232 (N_11232,N_11004,N_11009);
nand U11233 (N_11233,N_11047,N_11009);
nor U11234 (N_11234,N_11081,N_11013);
nand U11235 (N_11235,N_11093,N_11116);
and U11236 (N_11236,N_11109,N_11052);
xor U11237 (N_11237,N_11011,N_11124);
nand U11238 (N_11238,N_11017,N_11075);
and U11239 (N_11239,N_11052,N_11078);
and U11240 (N_11240,N_11039,N_11107);
or U11241 (N_11241,N_11094,N_11074);
xnor U11242 (N_11242,N_11032,N_11087);
nand U11243 (N_11243,N_11079,N_11102);
nand U11244 (N_11244,N_11015,N_11050);
or U11245 (N_11245,N_11023,N_11060);
nand U11246 (N_11246,N_11092,N_11080);
nor U11247 (N_11247,N_11096,N_11045);
or U11248 (N_11248,N_11032,N_11080);
xnor U11249 (N_11249,N_11005,N_11028);
and U11250 (N_11250,N_11164,N_11185);
and U11251 (N_11251,N_11240,N_11175);
xor U11252 (N_11252,N_11230,N_11207);
xor U11253 (N_11253,N_11160,N_11193);
nand U11254 (N_11254,N_11199,N_11203);
and U11255 (N_11255,N_11197,N_11153);
nand U11256 (N_11256,N_11239,N_11179);
and U11257 (N_11257,N_11138,N_11129);
and U11258 (N_11258,N_11169,N_11150);
or U11259 (N_11259,N_11167,N_11177);
nor U11260 (N_11260,N_11245,N_11187);
or U11261 (N_11261,N_11142,N_11152);
nand U11262 (N_11262,N_11228,N_11236);
and U11263 (N_11263,N_11154,N_11243);
and U11264 (N_11264,N_11180,N_11238);
xor U11265 (N_11265,N_11144,N_11229);
nand U11266 (N_11266,N_11231,N_11163);
nor U11267 (N_11267,N_11232,N_11168);
nor U11268 (N_11268,N_11139,N_11141);
or U11269 (N_11269,N_11202,N_11247);
and U11270 (N_11270,N_11221,N_11224);
xnor U11271 (N_11271,N_11217,N_11131);
nor U11272 (N_11272,N_11186,N_11216);
nand U11273 (N_11273,N_11205,N_11136);
and U11274 (N_11274,N_11151,N_11145);
nor U11275 (N_11275,N_11132,N_11206);
nand U11276 (N_11276,N_11227,N_11220);
and U11277 (N_11277,N_11219,N_11246);
xor U11278 (N_11278,N_11134,N_11210);
xor U11279 (N_11279,N_11182,N_11172);
xor U11280 (N_11280,N_11171,N_11198);
and U11281 (N_11281,N_11127,N_11148);
nor U11282 (N_11282,N_11176,N_11249);
or U11283 (N_11283,N_11194,N_11226);
nand U11284 (N_11284,N_11242,N_11183);
nand U11285 (N_11285,N_11174,N_11140);
nand U11286 (N_11286,N_11223,N_11222);
and U11287 (N_11287,N_11196,N_11162);
xnor U11288 (N_11288,N_11170,N_11125);
nand U11289 (N_11289,N_11211,N_11191);
or U11290 (N_11290,N_11133,N_11130);
and U11291 (N_11291,N_11200,N_11189);
xor U11292 (N_11292,N_11147,N_11178);
nand U11293 (N_11293,N_11173,N_11201);
and U11294 (N_11294,N_11248,N_11234);
xor U11295 (N_11295,N_11159,N_11225);
xor U11296 (N_11296,N_11188,N_11215);
or U11297 (N_11297,N_11208,N_11244);
and U11298 (N_11298,N_11213,N_11156);
nand U11299 (N_11299,N_11143,N_11158);
nand U11300 (N_11300,N_11204,N_11195);
nor U11301 (N_11301,N_11181,N_11149);
xnor U11302 (N_11302,N_11237,N_11184);
nor U11303 (N_11303,N_11126,N_11212);
nand U11304 (N_11304,N_11218,N_11146);
or U11305 (N_11305,N_11241,N_11161);
nand U11306 (N_11306,N_11192,N_11233);
nor U11307 (N_11307,N_11128,N_11155);
nor U11308 (N_11308,N_11235,N_11157);
nand U11309 (N_11309,N_11137,N_11166);
and U11310 (N_11310,N_11214,N_11135);
nand U11311 (N_11311,N_11209,N_11190);
nor U11312 (N_11312,N_11165,N_11164);
or U11313 (N_11313,N_11147,N_11222);
xor U11314 (N_11314,N_11162,N_11208);
and U11315 (N_11315,N_11153,N_11178);
nor U11316 (N_11316,N_11163,N_11156);
or U11317 (N_11317,N_11130,N_11189);
xnor U11318 (N_11318,N_11126,N_11159);
nor U11319 (N_11319,N_11241,N_11176);
nor U11320 (N_11320,N_11140,N_11175);
xnor U11321 (N_11321,N_11155,N_11150);
or U11322 (N_11322,N_11187,N_11212);
or U11323 (N_11323,N_11145,N_11159);
or U11324 (N_11324,N_11218,N_11132);
nand U11325 (N_11325,N_11207,N_11160);
nand U11326 (N_11326,N_11239,N_11193);
xor U11327 (N_11327,N_11182,N_11189);
nor U11328 (N_11328,N_11224,N_11192);
or U11329 (N_11329,N_11155,N_11178);
and U11330 (N_11330,N_11170,N_11129);
and U11331 (N_11331,N_11196,N_11210);
or U11332 (N_11332,N_11201,N_11168);
xor U11333 (N_11333,N_11232,N_11142);
xnor U11334 (N_11334,N_11151,N_11131);
or U11335 (N_11335,N_11153,N_11239);
or U11336 (N_11336,N_11162,N_11159);
and U11337 (N_11337,N_11145,N_11233);
xor U11338 (N_11338,N_11144,N_11227);
nand U11339 (N_11339,N_11238,N_11162);
nand U11340 (N_11340,N_11135,N_11233);
nor U11341 (N_11341,N_11190,N_11194);
nand U11342 (N_11342,N_11240,N_11209);
nand U11343 (N_11343,N_11208,N_11138);
xnor U11344 (N_11344,N_11181,N_11155);
or U11345 (N_11345,N_11200,N_11240);
and U11346 (N_11346,N_11245,N_11173);
nand U11347 (N_11347,N_11222,N_11220);
xor U11348 (N_11348,N_11188,N_11201);
nand U11349 (N_11349,N_11211,N_11142);
xnor U11350 (N_11350,N_11199,N_11142);
nor U11351 (N_11351,N_11147,N_11238);
nor U11352 (N_11352,N_11187,N_11227);
xor U11353 (N_11353,N_11143,N_11163);
and U11354 (N_11354,N_11243,N_11200);
nand U11355 (N_11355,N_11194,N_11160);
xor U11356 (N_11356,N_11223,N_11244);
nor U11357 (N_11357,N_11212,N_11221);
or U11358 (N_11358,N_11203,N_11204);
nor U11359 (N_11359,N_11143,N_11135);
xor U11360 (N_11360,N_11228,N_11234);
nor U11361 (N_11361,N_11127,N_11153);
nand U11362 (N_11362,N_11184,N_11206);
or U11363 (N_11363,N_11193,N_11155);
or U11364 (N_11364,N_11244,N_11189);
or U11365 (N_11365,N_11139,N_11237);
nor U11366 (N_11366,N_11133,N_11188);
nor U11367 (N_11367,N_11241,N_11240);
xnor U11368 (N_11368,N_11185,N_11127);
nor U11369 (N_11369,N_11153,N_11217);
and U11370 (N_11370,N_11203,N_11214);
nor U11371 (N_11371,N_11130,N_11165);
or U11372 (N_11372,N_11152,N_11219);
and U11373 (N_11373,N_11135,N_11205);
nand U11374 (N_11374,N_11239,N_11245);
nor U11375 (N_11375,N_11327,N_11320);
nand U11376 (N_11376,N_11281,N_11353);
xor U11377 (N_11377,N_11255,N_11299);
nor U11378 (N_11378,N_11371,N_11372);
and U11379 (N_11379,N_11274,N_11329);
xnor U11380 (N_11380,N_11270,N_11340);
or U11381 (N_11381,N_11286,N_11357);
or U11382 (N_11382,N_11288,N_11290);
xor U11383 (N_11383,N_11284,N_11355);
and U11384 (N_11384,N_11295,N_11252);
and U11385 (N_11385,N_11253,N_11336);
or U11386 (N_11386,N_11300,N_11254);
and U11387 (N_11387,N_11278,N_11356);
and U11388 (N_11388,N_11264,N_11360);
and U11389 (N_11389,N_11337,N_11368);
or U11390 (N_11390,N_11263,N_11346);
or U11391 (N_11391,N_11314,N_11351);
or U11392 (N_11392,N_11297,N_11266);
xor U11393 (N_11393,N_11362,N_11305);
nand U11394 (N_11394,N_11302,N_11365);
nand U11395 (N_11395,N_11341,N_11366);
nand U11396 (N_11396,N_11324,N_11352);
nand U11397 (N_11397,N_11277,N_11269);
and U11398 (N_11398,N_11309,N_11322);
nand U11399 (N_11399,N_11370,N_11313);
nand U11400 (N_11400,N_11294,N_11369);
or U11401 (N_11401,N_11258,N_11359);
xor U11402 (N_11402,N_11280,N_11328);
xnor U11403 (N_11403,N_11271,N_11317);
or U11404 (N_11404,N_11303,N_11316);
xor U11405 (N_11405,N_11310,N_11374);
or U11406 (N_11406,N_11259,N_11334);
and U11407 (N_11407,N_11331,N_11326);
nand U11408 (N_11408,N_11307,N_11339);
and U11409 (N_11409,N_11279,N_11256);
nand U11410 (N_11410,N_11338,N_11296);
xnor U11411 (N_11411,N_11349,N_11260);
nor U11412 (N_11412,N_11321,N_11291);
or U11413 (N_11413,N_11275,N_11282);
nor U11414 (N_11414,N_11268,N_11289);
nand U11415 (N_11415,N_11358,N_11267);
nor U11416 (N_11416,N_11287,N_11304);
xnor U11417 (N_11417,N_11318,N_11283);
nand U11418 (N_11418,N_11342,N_11308);
nor U11419 (N_11419,N_11276,N_11361);
nand U11420 (N_11420,N_11319,N_11311);
nor U11421 (N_11421,N_11257,N_11315);
xnor U11422 (N_11422,N_11343,N_11323);
and U11423 (N_11423,N_11265,N_11306);
or U11424 (N_11424,N_11262,N_11273);
or U11425 (N_11425,N_11373,N_11367);
nand U11426 (N_11426,N_11272,N_11335);
nand U11427 (N_11427,N_11292,N_11354);
nand U11428 (N_11428,N_11325,N_11330);
or U11429 (N_11429,N_11333,N_11348);
nand U11430 (N_11430,N_11332,N_11363);
or U11431 (N_11431,N_11364,N_11301);
and U11432 (N_11432,N_11298,N_11344);
nand U11433 (N_11433,N_11293,N_11261);
nor U11434 (N_11434,N_11250,N_11251);
xor U11435 (N_11435,N_11285,N_11312);
or U11436 (N_11436,N_11345,N_11347);
or U11437 (N_11437,N_11350,N_11250);
nand U11438 (N_11438,N_11372,N_11316);
nand U11439 (N_11439,N_11289,N_11309);
and U11440 (N_11440,N_11277,N_11301);
xnor U11441 (N_11441,N_11298,N_11254);
and U11442 (N_11442,N_11360,N_11349);
nand U11443 (N_11443,N_11338,N_11263);
or U11444 (N_11444,N_11252,N_11321);
nor U11445 (N_11445,N_11366,N_11373);
or U11446 (N_11446,N_11301,N_11355);
nor U11447 (N_11447,N_11343,N_11335);
xor U11448 (N_11448,N_11316,N_11288);
and U11449 (N_11449,N_11360,N_11333);
nand U11450 (N_11450,N_11321,N_11264);
or U11451 (N_11451,N_11261,N_11345);
or U11452 (N_11452,N_11373,N_11269);
nor U11453 (N_11453,N_11261,N_11339);
xnor U11454 (N_11454,N_11366,N_11359);
or U11455 (N_11455,N_11285,N_11317);
or U11456 (N_11456,N_11283,N_11338);
xnor U11457 (N_11457,N_11350,N_11279);
nor U11458 (N_11458,N_11369,N_11312);
and U11459 (N_11459,N_11272,N_11302);
and U11460 (N_11460,N_11259,N_11357);
xnor U11461 (N_11461,N_11292,N_11348);
nand U11462 (N_11462,N_11342,N_11338);
and U11463 (N_11463,N_11254,N_11282);
and U11464 (N_11464,N_11315,N_11274);
nand U11465 (N_11465,N_11351,N_11256);
nand U11466 (N_11466,N_11274,N_11283);
or U11467 (N_11467,N_11256,N_11338);
and U11468 (N_11468,N_11266,N_11366);
or U11469 (N_11469,N_11308,N_11346);
and U11470 (N_11470,N_11373,N_11340);
or U11471 (N_11471,N_11297,N_11280);
xnor U11472 (N_11472,N_11338,N_11367);
xnor U11473 (N_11473,N_11342,N_11339);
nor U11474 (N_11474,N_11280,N_11281);
nand U11475 (N_11475,N_11333,N_11317);
xor U11476 (N_11476,N_11364,N_11263);
and U11477 (N_11477,N_11308,N_11350);
and U11478 (N_11478,N_11342,N_11303);
or U11479 (N_11479,N_11374,N_11365);
nand U11480 (N_11480,N_11370,N_11328);
or U11481 (N_11481,N_11368,N_11287);
or U11482 (N_11482,N_11353,N_11340);
nor U11483 (N_11483,N_11336,N_11281);
nor U11484 (N_11484,N_11359,N_11334);
or U11485 (N_11485,N_11291,N_11304);
nand U11486 (N_11486,N_11292,N_11276);
nor U11487 (N_11487,N_11329,N_11343);
nand U11488 (N_11488,N_11260,N_11344);
nor U11489 (N_11489,N_11368,N_11316);
xnor U11490 (N_11490,N_11294,N_11273);
xor U11491 (N_11491,N_11339,N_11258);
nand U11492 (N_11492,N_11356,N_11354);
nand U11493 (N_11493,N_11360,N_11295);
nor U11494 (N_11494,N_11366,N_11365);
or U11495 (N_11495,N_11283,N_11290);
nor U11496 (N_11496,N_11269,N_11329);
or U11497 (N_11497,N_11366,N_11311);
xor U11498 (N_11498,N_11310,N_11270);
or U11499 (N_11499,N_11304,N_11286);
nand U11500 (N_11500,N_11391,N_11410);
or U11501 (N_11501,N_11458,N_11386);
nand U11502 (N_11502,N_11387,N_11456);
and U11503 (N_11503,N_11419,N_11470);
or U11504 (N_11504,N_11380,N_11482);
and U11505 (N_11505,N_11465,N_11473);
nor U11506 (N_11506,N_11427,N_11494);
nor U11507 (N_11507,N_11488,N_11397);
xnor U11508 (N_11508,N_11406,N_11411);
nand U11509 (N_11509,N_11455,N_11394);
or U11510 (N_11510,N_11404,N_11375);
or U11511 (N_11511,N_11441,N_11491);
nor U11512 (N_11512,N_11412,N_11384);
or U11513 (N_11513,N_11442,N_11415);
and U11514 (N_11514,N_11477,N_11451);
and U11515 (N_11515,N_11424,N_11408);
xnor U11516 (N_11516,N_11421,N_11498);
and U11517 (N_11517,N_11385,N_11377);
or U11518 (N_11518,N_11446,N_11471);
nand U11519 (N_11519,N_11459,N_11378);
nand U11520 (N_11520,N_11463,N_11420);
nand U11521 (N_11521,N_11390,N_11487);
nand U11522 (N_11522,N_11423,N_11413);
xor U11523 (N_11523,N_11399,N_11433);
nand U11524 (N_11524,N_11483,N_11416);
nand U11525 (N_11525,N_11418,N_11492);
xor U11526 (N_11526,N_11382,N_11388);
xor U11527 (N_11527,N_11429,N_11381);
nand U11528 (N_11528,N_11435,N_11403);
and U11529 (N_11529,N_11448,N_11430);
xnor U11530 (N_11530,N_11445,N_11496);
and U11531 (N_11531,N_11490,N_11431);
or U11532 (N_11532,N_11467,N_11393);
or U11533 (N_11533,N_11398,N_11480);
and U11534 (N_11534,N_11439,N_11379);
or U11535 (N_11535,N_11401,N_11464);
nand U11536 (N_11536,N_11395,N_11414);
xor U11537 (N_11537,N_11447,N_11383);
and U11538 (N_11538,N_11438,N_11462);
nand U11539 (N_11539,N_11432,N_11417);
nand U11540 (N_11540,N_11453,N_11485);
and U11541 (N_11541,N_11426,N_11497);
nor U11542 (N_11542,N_11457,N_11472);
or U11543 (N_11543,N_11461,N_11376);
nor U11544 (N_11544,N_11479,N_11454);
or U11545 (N_11545,N_11481,N_11434);
and U11546 (N_11546,N_11409,N_11475);
nand U11547 (N_11547,N_11422,N_11476);
xnor U11548 (N_11548,N_11474,N_11468);
and U11549 (N_11549,N_11436,N_11452);
and U11550 (N_11550,N_11449,N_11407);
or U11551 (N_11551,N_11392,N_11405);
nand U11552 (N_11552,N_11450,N_11460);
nor U11553 (N_11553,N_11466,N_11440);
and U11554 (N_11554,N_11428,N_11489);
or U11555 (N_11555,N_11484,N_11469);
nor U11556 (N_11556,N_11389,N_11478);
and U11557 (N_11557,N_11443,N_11396);
and U11558 (N_11558,N_11493,N_11425);
nor U11559 (N_11559,N_11486,N_11499);
nor U11560 (N_11560,N_11402,N_11444);
or U11561 (N_11561,N_11437,N_11495);
xnor U11562 (N_11562,N_11400,N_11392);
or U11563 (N_11563,N_11465,N_11464);
nor U11564 (N_11564,N_11476,N_11414);
or U11565 (N_11565,N_11479,N_11418);
nor U11566 (N_11566,N_11381,N_11481);
xnor U11567 (N_11567,N_11487,N_11383);
xnor U11568 (N_11568,N_11430,N_11481);
and U11569 (N_11569,N_11398,N_11462);
nand U11570 (N_11570,N_11482,N_11403);
xnor U11571 (N_11571,N_11418,N_11488);
or U11572 (N_11572,N_11410,N_11405);
or U11573 (N_11573,N_11384,N_11439);
nor U11574 (N_11574,N_11394,N_11482);
and U11575 (N_11575,N_11412,N_11407);
and U11576 (N_11576,N_11432,N_11474);
xnor U11577 (N_11577,N_11401,N_11378);
and U11578 (N_11578,N_11455,N_11415);
or U11579 (N_11579,N_11443,N_11464);
and U11580 (N_11580,N_11472,N_11483);
nand U11581 (N_11581,N_11452,N_11466);
and U11582 (N_11582,N_11447,N_11460);
nor U11583 (N_11583,N_11390,N_11489);
nor U11584 (N_11584,N_11456,N_11440);
nor U11585 (N_11585,N_11454,N_11490);
xnor U11586 (N_11586,N_11390,N_11420);
or U11587 (N_11587,N_11453,N_11401);
or U11588 (N_11588,N_11387,N_11465);
xnor U11589 (N_11589,N_11454,N_11493);
nor U11590 (N_11590,N_11398,N_11493);
xor U11591 (N_11591,N_11444,N_11494);
and U11592 (N_11592,N_11404,N_11491);
and U11593 (N_11593,N_11382,N_11415);
xnor U11594 (N_11594,N_11417,N_11460);
and U11595 (N_11595,N_11490,N_11439);
or U11596 (N_11596,N_11413,N_11419);
and U11597 (N_11597,N_11413,N_11386);
and U11598 (N_11598,N_11396,N_11388);
xnor U11599 (N_11599,N_11377,N_11424);
nor U11600 (N_11600,N_11438,N_11433);
and U11601 (N_11601,N_11442,N_11412);
nand U11602 (N_11602,N_11450,N_11399);
and U11603 (N_11603,N_11447,N_11424);
nor U11604 (N_11604,N_11426,N_11377);
nand U11605 (N_11605,N_11391,N_11490);
nor U11606 (N_11606,N_11474,N_11392);
nor U11607 (N_11607,N_11390,N_11494);
nand U11608 (N_11608,N_11494,N_11421);
and U11609 (N_11609,N_11491,N_11396);
and U11610 (N_11610,N_11444,N_11455);
nor U11611 (N_11611,N_11384,N_11432);
and U11612 (N_11612,N_11445,N_11414);
and U11613 (N_11613,N_11406,N_11403);
or U11614 (N_11614,N_11409,N_11466);
xnor U11615 (N_11615,N_11412,N_11448);
and U11616 (N_11616,N_11440,N_11447);
xor U11617 (N_11617,N_11397,N_11427);
and U11618 (N_11618,N_11463,N_11384);
or U11619 (N_11619,N_11432,N_11455);
xor U11620 (N_11620,N_11471,N_11412);
and U11621 (N_11621,N_11377,N_11442);
nor U11622 (N_11622,N_11437,N_11473);
nor U11623 (N_11623,N_11393,N_11459);
nand U11624 (N_11624,N_11469,N_11400);
xnor U11625 (N_11625,N_11609,N_11531);
xnor U11626 (N_11626,N_11595,N_11619);
nor U11627 (N_11627,N_11538,N_11580);
xor U11628 (N_11628,N_11577,N_11551);
xnor U11629 (N_11629,N_11616,N_11511);
nand U11630 (N_11630,N_11588,N_11516);
nand U11631 (N_11631,N_11565,N_11547);
xnor U11632 (N_11632,N_11546,N_11549);
xor U11633 (N_11633,N_11552,N_11584);
nor U11634 (N_11634,N_11581,N_11526);
and U11635 (N_11635,N_11600,N_11621);
or U11636 (N_11636,N_11512,N_11611);
or U11637 (N_11637,N_11521,N_11576);
nand U11638 (N_11638,N_11540,N_11561);
or U11639 (N_11639,N_11541,N_11567);
or U11640 (N_11640,N_11523,N_11542);
or U11641 (N_11641,N_11519,N_11624);
or U11642 (N_11642,N_11504,N_11507);
nor U11643 (N_11643,N_11501,N_11613);
nand U11644 (N_11644,N_11596,N_11590);
xor U11645 (N_11645,N_11559,N_11524);
nor U11646 (N_11646,N_11614,N_11607);
or U11647 (N_11647,N_11599,N_11608);
nor U11648 (N_11648,N_11536,N_11601);
nor U11649 (N_11649,N_11537,N_11593);
nor U11650 (N_11650,N_11605,N_11570);
nor U11651 (N_11651,N_11583,N_11517);
nor U11652 (N_11652,N_11503,N_11587);
nor U11653 (N_11653,N_11500,N_11532);
and U11654 (N_11654,N_11569,N_11555);
xor U11655 (N_11655,N_11586,N_11527);
nor U11656 (N_11656,N_11513,N_11618);
nand U11657 (N_11657,N_11502,N_11564);
xnor U11658 (N_11658,N_11566,N_11622);
xor U11659 (N_11659,N_11592,N_11515);
nor U11660 (N_11660,N_11545,N_11548);
nand U11661 (N_11661,N_11602,N_11603);
xnor U11662 (N_11662,N_11525,N_11579);
or U11663 (N_11663,N_11589,N_11558);
xor U11664 (N_11664,N_11560,N_11571);
nor U11665 (N_11665,N_11506,N_11594);
nor U11666 (N_11666,N_11617,N_11568);
nand U11667 (N_11667,N_11505,N_11591);
nor U11668 (N_11668,N_11509,N_11574);
or U11669 (N_11669,N_11562,N_11508);
and U11670 (N_11670,N_11620,N_11578);
and U11671 (N_11671,N_11556,N_11539);
xnor U11672 (N_11672,N_11572,N_11615);
nor U11673 (N_11673,N_11612,N_11598);
xnor U11674 (N_11674,N_11530,N_11533);
nor U11675 (N_11675,N_11575,N_11534);
nand U11676 (N_11676,N_11557,N_11623);
xnor U11677 (N_11677,N_11522,N_11582);
nor U11678 (N_11678,N_11573,N_11543);
and U11679 (N_11679,N_11528,N_11563);
nor U11680 (N_11680,N_11544,N_11529);
or U11681 (N_11681,N_11597,N_11553);
nand U11682 (N_11682,N_11554,N_11585);
nor U11683 (N_11683,N_11520,N_11535);
xnor U11684 (N_11684,N_11550,N_11604);
xor U11685 (N_11685,N_11510,N_11514);
and U11686 (N_11686,N_11606,N_11518);
xnor U11687 (N_11687,N_11610,N_11609);
or U11688 (N_11688,N_11595,N_11548);
or U11689 (N_11689,N_11521,N_11506);
nand U11690 (N_11690,N_11559,N_11503);
nand U11691 (N_11691,N_11611,N_11575);
nor U11692 (N_11692,N_11503,N_11611);
xor U11693 (N_11693,N_11505,N_11603);
xor U11694 (N_11694,N_11605,N_11616);
nor U11695 (N_11695,N_11590,N_11618);
and U11696 (N_11696,N_11504,N_11574);
xor U11697 (N_11697,N_11621,N_11540);
xnor U11698 (N_11698,N_11621,N_11578);
nor U11699 (N_11699,N_11538,N_11527);
and U11700 (N_11700,N_11620,N_11555);
xor U11701 (N_11701,N_11501,N_11579);
or U11702 (N_11702,N_11565,N_11520);
nand U11703 (N_11703,N_11525,N_11564);
xor U11704 (N_11704,N_11504,N_11544);
xnor U11705 (N_11705,N_11521,N_11513);
nand U11706 (N_11706,N_11570,N_11547);
nand U11707 (N_11707,N_11601,N_11552);
or U11708 (N_11708,N_11529,N_11520);
nor U11709 (N_11709,N_11534,N_11545);
nor U11710 (N_11710,N_11588,N_11566);
and U11711 (N_11711,N_11577,N_11518);
or U11712 (N_11712,N_11580,N_11583);
or U11713 (N_11713,N_11552,N_11510);
or U11714 (N_11714,N_11530,N_11604);
nand U11715 (N_11715,N_11591,N_11568);
xor U11716 (N_11716,N_11569,N_11556);
xnor U11717 (N_11717,N_11590,N_11511);
nor U11718 (N_11718,N_11551,N_11615);
xnor U11719 (N_11719,N_11599,N_11620);
or U11720 (N_11720,N_11608,N_11614);
and U11721 (N_11721,N_11601,N_11532);
nand U11722 (N_11722,N_11502,N_11537);
xnor U11723 (N_11723,N_11603,N_11586);
and U11724 (N_11724,N_11624,N_11527);
and U11725 (N_11725,N_11584,N_11596);
nand U11726 (N_11726,N_11604,N_11545);
and U11727 (N_11727,N_11597,N_11608);
or U11728 (N_11728,N_11549,N_11598);
nor U11729 (N_11729,N_11567,N_11534);
nor U11730 (N_11730,N_11504,N_11529);
and U11731 (N_11731,N_11501,N_11548);
xor U11732 (N_11732,N_11599,N_11594);
xnor U11733 (N_11733,N_11556,N_11510);
or U11734 (N_11734,N_11609,N_11571);
xor U11735 (N_11735,N_11533,N_11531);
xnor U11736 (N_11736,N_11586,N_11564);
nor U11737 (N_11737,N_11515,N_11543);
nor U11738 (N_11738,N_11502,N_11544);
and U11739 (N_11739,N_11617,N_11540);
nand U11740 (N_11740,N_11546,N_11522);
xor U11741 (N_11741,N_11540,N_11570);
nor U11742 (N_11742,N_11572,N_11534);
nor U11743 (N_11743,N_11556,N_11542);
nand U11744 (N_11744,N_11538,N_11502);
or U11745 (N_11745,N_11593,N_11542);
or U11746 (N_11746,N_11583,N_11620);
or U11747 (N_11747,N_11518,N_11504);
xor U11748 (N_11748,N_11624,N_11535);
nand U11749 (N_11749,N_11535,N_11603);
and U11750 (N_11750,N_11734,N_11689);
xnor U11751 (N_11751,N_11677,N_11720);
or U11752 (N_11752,N_11703,N_11675);
and U11753 (N_11753,N_11690,N_11641);
and U11754 (N_11754,N_11652,N_11711);
xor U11755 (N_11755,N_11634,N_11732);
or U11756 (N_11756,N_11716,N_11638);
xor U11757 (N_11757,N_11661,N_11743);
nor U11758 (N_11758,N_11678,N_11653);
or U11759 (N_11759,N_11747,N_11713);
or U11760 (N_11760,N_11680,N_11635);
nand U11761 (N_11761,N_11651,N_11649);
and U11762 (N_11762,N_11637,N_11633);
nor U11763 (N_11763,N_11659,N_11715);
or U11764 (N_11764,N_11710,N_11670);
and U11765 (N_11765,N_11654,N_11636);
or U11766 (N_11766,N_11669,N_11682);
nand U11767 (N_11767,N_11665,N_11681);
or U11768 (N_11768,N_11664,N_11658);
nor U11769 (N_11769,N_11740,N_11714);
and U11770 (N_11770,N_11679,N_11643);
or U11771 (N_11771,N_11663,N_11712);
xor U11772 (N_11772,N_11697,N_11729);
nand U11773 (N_11773,N_11724,N_11736);
nor U11774 (N_11774,N_11684,N_11674);
or U11775 (N_11775,N_11647,N_11671);
xnor U11776 (N_11776,N_11625,N_11629);
nor U11777 (N_11777,N_11672,N_11630);
xnor U11778 (N_11778,N_11639,N_11662);
and U11779 (N_11779,N_11640,N_11696);
and U11780 (N_11780,N_11685,N_11704);
or U11781 (N_11781,N_11718,N_11688);
nand U11782 (N_11782,N_11737,N_11748);
xor U11783 (N_11783,N_11701,N_11699);
or U11784 (N_11784,N_11723,N_11705);
xor U11785 (N_11785,N_11683,N_11744);
xnor U11786 (N_11786,N_11698,N_11668);
xnor U11787 (N_11787,N_11627,N_11650);
and U11788 (N_11788,N_11739,N_11692);
or U11789 (N_11789,N_11632,N_11695);
or U11790 (N_11790,N_11673,N_11721);
xnor U11791 (N_11791,N_11719,N_11656);
nor U11792 (N_11792,N_11733,N_11655);
xor U11793 (N_11793,N_11666,N_11738);
nor U11794 (N_11794,N_11645,N_11687);
xor U11795 (N_11795,N_11706,N_11707);
or U11796 (N_11796,N_11646,N_11626);
nor U11797 (N_11797,N_11694,N_11691);
xnor U11798 (N_11798,N_11749,N_11709);
nor U11799 (N_11799,N_11660,N_11725);
or U11800 (N_11800,N_11731,N_11631);
or U11801 (N_11801,N_11657,N_11727);
xor U11802 (N_11802,N_11717,N_11667);
or U11803 (N_11803,N_11642,N_11628);
xor U11804 (N_11804,N_11700,N_11644);
or U11805 (N_11805,N_11730,N_11676);
xor U11806 (N_11806,N_11708,N_11741);
nand U11807 (N_11807,N_11726,N_11686);
and U11808 (N_11808,N_11648,N_11745);
and U11809 (N_11809,N_11746,N_11722);
nand U11810 (N_11810,N_11742,N_11735);
or U11811 (N_11811,N_11693,N_11702);
xor U11812 (N_11812,N_11728,N_11681);
nand U11813 (N_11813,N_11648,N_11738);
nor U11814 (N_11814,N_11672,N_11734);
nand U11815 (N_11815,N_11627,N_11697);
nor U11816 (N_11816,N_11662,N_11744);
nor U11817 (N_11817,N_11661,N_11652);
and U11818 (N_11818,N_11631,N_11713);
nor U11819 (N_11819,N_11638,N_11702);
nand U11820 (N_11820,N_11723,N_11740);
or U11821 (N_11821,N_11730,N_11679);
xor U11822 (N_11822,N_11643,N_11707);
nand U11823 (N_11823,N_11687,N_11651);
and U11824 (N_11824,N_11732,N_11631);
or U11825 (N_11825,N_11690,N_11632);
nand U11826 (N_11826,N_11723,N_11635);
xor U11827 (N_11827,N_11706,N_11712);
nand U11828 (N_11828,N_11695,N_11726);
xor U11829 (N_11829,N_11728,N_11689);
and U11830 (N_11830,N_11664,N_11715);
and U11831 (N_11831,N_11645,N_11691);
or U11832 (N_11832,N_11696,N_11639);
nand U11833 (N_11833,N_11679,N_11629);
nand U11834 (N_11834,N_11727,N_11717);
xor U11835 (N_11835,N_11654,N_11730);
nor U11836 (N_11836,N_11641,N_11717);
or U11837 (N_11837,N_11666,N_11636);
or U11838 (N_11838,N_11725,N_11657);
or U11839 (N_11839,N_11644,N_11688);
nand U11840 (N_11840,N_11649,N_11694);
xor U11841 (N_11841,N_11716,N_11667);
nor U11842 (N_11842,N_11713,N_11731);
xnor U11843 (N_11843,N_11629,N_11686);
or U11844 (N_11844,N_11655,N_11689);
or U11845 (N_11845,N_11684,N_11689);
and U11846 (N_11846,N_11662,N_11716);
or U11847 (N_11847,N_11666,N_11745);
nand U11848 (N_11848,N_11677,N_11663);
nor U11849 (N_11849,N_11636,N_11679);
nand U11850 (N_11850,N_11662,N_11682);
and U11851 (N_11851,N_11702,N_11660);
or U11852 (N_11852,N_11660,N_11737);
xnor U11853 (N_11853,N_11725,N_11726);
nand U11854 (N_11854,N_11635,N_11720);
xnor U11855 (N_11855,N_11639,N_11626);
nor U11856 (N_11856,N_11729,N_11683);
nand U11857 (N_11857,N_11631,N_11682);
nor U11858 (N_11858,N_11629,N_11741);
nand U11859 (N_11859,N_11707,N_11645);
nor U11860 (N_11860,N_11675,N_11664);
xnor U11861 (N_11861,N_11639,N_11723);
nor U11862 (N_11862,N_11687,N_11642);
nor U11863 (N_11863,N_11688,N_11645);
and U11864 (N_11864,N_11696,N_11729);
nand U11865 (N_11865,N_11724,N_11657);
and U11866 (N_11866,N_11748,N_11636);
and U11867 (N_11867,N_11718,N_11744);
or U11868 (N_11868,N_11719,N_11710);
xor U11869 (N_11869,N_11719,N_11725);
or U11870 (N_11870,N_11738,N_11711);
xnor U11871 (N_11871,N_11644,N_11714);
nand U11872 (N_11872,N_11719,N_11658);
and U11873 (N_11873,N_11737,N_11679);
nor U11874 (N_11874,N_11733,N_11656);
xor U11875 (N_11875,N_11820,N_11852);
and U11876 (N_11876,N_11765,N_11850);
nor U11877 (N_11877,N_11816,N_11770);
xnor U11878 (N_11878,N_11763,N_11803);
nand U11879 (N_11879,N_11817,N_11869);
and U11880 (N_11880,N_11789,N_11751);
nor U11881 (N_11881,N_11785,N_11856);
xnor U11882 (N_11882,N_11872,N_11835);
xnor U11883 (N_11883,N_11792,N_11854);
or U11884 (N_11884,N_11855,N_11857);
or U11885 (N_11885,N_11756,N_11810);
xor U11886 (N_11886,N_11818,N_11762);
nand U11887 (N_11887,N_11863,N_11750);
or U11888 (N_11888,N_11831,N_11809);
and U11889 (N_11889,N_11859,N_11757);
xor U11890 (N_11890,N_11851,N_11798);
or U11891 (N_11891,N_11844,N_11759);
or U11892 (N_11892,N_11777,N_11769);
or U11893 (N_11893,N_11853,N_11841);
xor U11894 (N_11894,N_11767,N_11823);
and U11895 (N_11895,N_11801,N_11834);
or U11896 (N_11896,N_11788,N_11752);
xor U11897 (N_11897,N_11813,N_11866);
nand U11898 (N_11898,N_11864,N_11774);
or U11899 (N_11899,N_11827,N_11848);
nor U11900 (N_11900,N_11807,N_11782);
and U11901 (N_11901,N_11815,N_11806);
or U11902 (N_11902,N_11768,N_11867);
or U11903 (N_11903,N_11843,N_11758);
and U11904 (N_11904,N_11830,N_11786);
and U11905 (N_11905,N_11861,N_11865);
nor U11906 (N_11906,N_11760,N_11793);
nor U11907 (N_11907,N_11804,N_11838);
nor U11908 (N_11908,N_11772,N_11870);
and U11909 (N_11909,N_11833,N_11828);
or U11910 (N_11910,N_11784,N_11874);
and U11911 (N_11911,N_11825,N_11790);
xnor U11912 (N_11912,N_11754,N_11871);
or U11913 (N_11913,N_11814,N_11766);
or U11914 (N_11914,N_11780,N_11824);
nand U11915 (N_11915,N_11821,N_11862);
and U11916 (N_11916,N_11808,N_11773);
nand U11917 (N_11917,N_11832,N_11842);
nand U11918 (N_11918,N_11778,N_11771);
and U11919 (N_11919,N_11873,N_11755);
nand U11920 (N_11920,N_11840,N_11812);
or U11921 (N_11921,N_11860,N_11829);
nor U11922 (N_11922,N_11753,N_11846);
and U11923 (N_11923,N_11849,N_11775);
nand U11924 (N_11924,N_11847,N_11795);
nand U11925 (N_11925,N_11802,N_11783);
nand U11926 (N_11926,N_11791,N_11822);
nand U11927 (N_11927,N_11800,N_11794);
nand U11928 (N_11928,N_11805,N_11796);
nor U11929 (N_11929,N_11845,N_11787);
or U11930 (N_11930,N_11797,N_11764);
nand U11931 (N_11931,N_11836,N_11858);
or U11932 (N_11932,N_11811,N_11799);
and U11933 (N_11933,N_11781,N_11868);
nand U11934 (N_11934,N_11826,N_11839);
nor U11935 (N_11935,N_11776,N_11779);
and U11936 (N_11936,N_11837,N_11761);
xor U11937 (N_11937,N_11819,N_11857);
and U11938 (N_11938,N_11779,N_11794);
nor U11939 (N_11939,N_11825,N_11760);
and U11940 (N_11940,N_11872,N_11760);
nand U11941 (N_11941,N_11827,N_11870);
xnor U11942 (N_11942,N_11754,N_11833);
and U11943 (N_11943,N_11810,N_11799);
nand U11944 (N_11944,N_11829,N_11863);
or U11945 (N_11945,N_11825,N_11777);
nand U11946 (N_11946,N_11759,N_11862);
nand U11947 (N_11947,N_11811,N_11866);
nor U11948 (N_11948,N_11813,N_11845);
xor U11949 (N_11949,N_11799,N_11838);
nand U11950 (N_11950,N_11761,N_11847);
nor U11951 (N_11951,N_11813,N_11779);
or U11952 (N_11952,N_11832,N_11807);
nor U11953 (N_11953,N_11829,N_11793);
and U11954 (N_11954,N_11845,N_11764);
nand U11955 (N_11955,N_11765,N_11792);
xnor U11956 (N_11956,N_11819,N_11813);
xnor U11957 (N_11957,N_11772,N_11818);
nand U11958 (N_11958,N_11806,N_11788);
nor U11959 (N_11959,N_11780,N_11857);
nand U11960 (N_11960,N_11772,N_11764);
and U11961 (N_11961,N_11811,N_11812);
xor U11962 (N_11962,N_11797,N_11851);
nor U11963 (N_11963,N_11795,N_11840);
xnor U11964 (N_11964,N_11783,N_11867);
or U11965 (N_11965,N_11769,N_11752);
nor U11966 (N_11966,N_11872,N_11763);
or U11967 (N_11967,N_11870,N_11787);
nor U11968 (N_11968,N_11844,N_11799);
nor U11969 (N_11969,N_11789,N_11773);
or U11970 (N_11970,N_11760,N_11774);
or U11971 (N_11971,N_11789,N_11753);
or U11972 (N_11972,N_11757,N_11811);
or U11973 (N_11973,N_11805,N_11774);
or U11974 (N_11974,N_11845,N_11778);
or U11975 (N_11975,N_11834,N_11814);
xnor U11976 (N_11976,N_11760,N_11811);
nor U11977 (N_11977,N_11833,N_11832);
xor U11978 (N_11978,N_11812,N_11847);
nand U11979 (N_11979,N_11866,N_11773);
xor U11980 (N_11980,N_11760,N_11803);
nor U11981 (N_11981,N_11863,N_11799);
xor U11982 (N_11982,N_11753,N_11780);
nor U11983 (N_11983,N_11830,N_11792);
or U11984 (N_11984,N_11794,N_11826);
and U11985 (N_11985,N_11788,N_11808);
nor U11986 (N_11986,N_11828,N_11787);
or U11987 (N_11987,N_11857,N_11862);
or U11988 (N_11988,N_11766,N_11794);
or U11989 (N_11989,N_11767,N_11824);
or U11990 (N_11990,N_11836,N_11833);
or U11991 (N_11991,N_11871,N_11850);
nor U11992 (N_11992,N_11775,N_11754);
xor U11993 (N_11993,N_11831,N_11865);
xor U11994 (N_11994,N_11816,N_11823);
or U11995 (N_11995,N_11867,N_11863);
nor U11996 (N_11996,N_11867,N_11839);
or U11997 (N_11997,N_11773,N_11778);
nand U11998 (N_11998,N_11756,N_11809);
nor U11999 (N_11999,N_11799,N_11864);
or U12000 (N_12000,N_11911,N_11945);
nand U12001 (N_12001,N_11988,N_11899);
or U12002 (N_12002,N_11953,N_11881);
nor U12003 (N_12003,N_11955,N_11992);
xnor U12004 (N_12004,N_11980,N_11925);
nor U12005 (N_12005,N_11879,N_11969);
nand U12006 (N_12006,N_11904,N_11933);
nor U12007 (N_12007,N_11885,N_11944);
xor U12008 (N_12008,N_11948,N_11954);
xor U12009 (N_12009,N_11993,N_11985);
nand U12010 (N_12010,N_11887,N_11943);
xor U12011 (N_12011,N_11908,N_11981);
nor U12012 (N_12012,N_11877,N_11882);
xnor U12013 (N_12013,N_11990,N_11976);
and U12014 (N_12014,N_11940,N_11906);
or U12015 (N_12015,N_11889,N_11966);
or U12016 (N_12016,N_11936,N_11901);
nor U12017 (N_12017,N_11995,N_11912);
or U12018 (N_12018,N_11907,N_11975);
and U12019 (N_12019,N_11997,N_11909);
or U12020 (N_12020,N_11958,N_11898);
xnor U12021 (N_12021,N_11935,N_11914);
and U12022 (N_12022,N_11890,N_11983);
nand U12023 (N_12023,N_11959,N_11949);
xnor U12024 (N_12024,N_11961,N_11915);
nand U12025 (N_12025,N_11896,N_11970);
nand U12026 (N_12026,N_11893,N_11886);
or U12027 (N_12027,N_11876,N_11986);
nor U12028 (N_12028,N_11878,N_11957);
nor U12029 (N_12029,N_11977,N_11875);
or U12030 (N_12030,N_11964,N_11987);
and U12031 (N_12031,N_11938,N_11895);
or U12032 (N_12032,N_11952,N_11973);
and U12033 (N_12033,N_11978,N_11941);
and U12034 (N_12034,N_11965,N_11891);
nor U12035 (N_12035,N_11918,N_11921);
nor U12036 (N_12036,N_11897,N_11930);
or U12037 (N_12037,N_11994,N_11971);
nor U12038 (N_12038,N_11942,N_11905);
nand U12039 (N_12039,N_11910,N_11946);
nor U12040 (N_12040,N_11989,N_11968);
and U12041 (N_12041,N_11888,N_11928);
and U12042 (N_12042,N_11916,N_11972);
nand U12043 (N_12043,N_11926,N_11924);
nor U12044 (N_12044,N_11894,N_11892);
or U12045 (N_12045,N_11947,N_11996);
and U12046 (N_12046,N_11967,N_11927);
and U12047 (N_12047,N_11931,N_11951);
and U12048 (N_12048,N_11974,N_11982);
nand U12049 (N_12049,N_11950,N_11883);
xnor U12050 (N_12050,N_11903,N_11929);
nor U12051 (N_12051,N_11991,N_11984);
and U12052 (N_12052,N_11923,N_11919);
and U12053 (N_12053,N_11963,N_11937);
and U12054 (N_12054,N_11956,N_11900);
and U12055 (N_12055,N_11934,N_11902);
xor U12056 (N_12056,N_11922,N_11932);
nor U12057 (N_12057,N_11880,N_11913);
xor U12058 (N_12058,N_11917,N_11999);
nand U12059 (N_12059,N_11920,N_11962);
or U12060 (N_12060,N_11939,N_11884);
and U12061 (N_12061,N_11979,N_11998);
and U12062 (N_12062,N_11960,N_11904);
or U12063 (N_12063,N_11968,N_11960);
xor U12064 (N_12064,N_11919,N_11921);
nor U12065 (N_12065,N_11894,N_11923);
and U12066 (N_12066,N_11892,N_11897);
xor U12067 (N_12067,N_11941,N_11875);
or U12068 (N_12068,N_11989,N_11882);
nor U12069 (N_12069,N_11941,N_11961);
nand U12070 (N_12070,N_11879,N_11927);
xor U12071 (N_12071,N_11975,N_11885);
and U12072 (N_12072,N_11912,N_11900);
xnor U12073 (N_12073,N_11886,N_11954);
and U12074 (N_12074,N_11987,N_11996);
nor U12075 (N_12075,N_11925,N_11916);
xnor U12076 (N_12076,N_11950,N_11899);
nand U12077 (N_12077,N_11923,N_11901);
xnor U12078 (N_12078,N_11966,N_11898);
and U12079 (N_12079,N_11947,N_11932);
xor U12080 (N_12080,N_11931,N_11934);
nand U12081 (N_12081,N_11913,N_11899);
nor U12082 (N_12082,N_11969,N_11935);
and U12083 (N_12083,N_11988,N_11927);
and U12084 (N_12084,N_11974,N_11961);
xnor U12085 (N_12085,N_11882,N_11958);
nand U12086 (N_12086,N_11928,N_11894);
nor U12087 (N_12087,N_11950,N_11982);
or U12088 (N_12088,N_11939,N_11878);
and U12089 (N_12089,N_11969,N_11885);
or U12090 (N_12090,N_11917,N_11925);
nand U12091 (N_12091,N_11949,N_11902);
nor U12092 (N_12092,N_11979,N_11958);
xor U12093 (N_12093,N_11947,N_11904);
nand U12094 (N_12094,N_11909,N_11953);
nand U12095 (N_12095,N_11914,N_11974);
nor U12096 (N_12096,N_11931,N_11891);
nand U12097 (N_12097,N_11967,N_11930);
and U12098 (N_12098,N_11977,N_11903);
xnor U12099 (N_12099,N_11992,N_11946);
and U12100 (N_12100,N_11981,N_11892);
or U12101 (N_12101,N_11882,N_11875);
xnor U12102 (N_12102,N_11943,N_11888);
and U12103 (N_12103,N_11991,N_11892);
nand U12104 (N_12104,N_11929,N_11922);
nor U12105 (N_12105,N_11897,N_11919);
xor U12106 (N_12106,N_11947,N_11878);
or U12107 (N_12107,N_11947,N_11939);
and U12108 (N_12108,N_11933,N_11964);
nor U12109 (N_12109,N_11912,N_11957);
or U12110 (N_12110,N_11905,N_11931);
nor U12111 (N_12111,N_11895,N_11972);
xor U12112 (N_12112,N_11962,N_11932);
and U12113 (N_12113,N_11972,N_11995);
xor U12114 (N_12114,N_11932,N_11890);
and U12115 (N_12115,N_11976,N_11887);
and U12116 (N_12116,N_11937,N_11882);
xnor U12117 (N_12117,N_11884,N_11901);
nor U12118 (N_12118,N_11933,N_11945);
nor U12119 (N_12119,N_11981,N_11927);
or U12120 (N_12120,N_11958,N_11893);
and U12121 (N_12121,N_11943,N_11902);
nand U12122 (N_12122,N_11921,N_11993);
nand U12123 (N_12123,N_11970,N_11922);
and U12124 (N_12124,N_11975,N_11956);
xor U12125 (N_12125,N_12042,N_12049);
nor U12126 (N_12126,N_12111,N_12097);
and U12127 (N_12127,N_12030,N_12032);
nand U12128 (N_12128,N_12122,N_12092);
nor U12129 (N_12129,N_12113,N_12057);
xor U12130 (N_12130,N_12034,N_12017);
nor U12131 (N_12131,N_12119,N_12053);
or U12132 (N_12132,N_12020,N_12101);
xor U12133 (N_12133,N_12073,N_12090);
nand U12134 (N_12134,N_12060,N_12071);
nand U12135 (N_12135,N_12118,N_12027);
or U12136 (N_12136,N_12108,N_12091);
nand U12137 (N_12137,N_12123,N_12079);
xnor U12138 (N_12138,N_12100,N_12089);
or U12139 (N_12139,N_12063,N_12067);
or U12140 (N_12140,N_12099,N_12096);
xor U12141 (N_12141,N_12052,N_12103);
nand U12142 (N_12142,N_12094,N_12045);
nand U12143 (N_12143,N_12084,N_12033);
nand U12144 (N_12144,N_12044,N_12066);
nand U12145 (N_12145,N_12115,N_12098);
xor U12146 (N_12146,N_12062,N_12016);
and U12147 (N_12147,N_12048,N_12005);
nor U12148 (N_12148,N_12117,N_12024);
xor U12149 (N_12149,N_12028,N_12035);
nor U12150 (N_12150,N_12031,N_12061);
or U12151 (N_12151,N_12075,N_12043);
xor U12152 (N_12152,N_12077,N_12010);
or U12153 (N_12153,N_12065,N_12055);
and U12154 (N_12154,N_12102,N_12085);
or U12155 (N_12155,N_12106,N_12041);
xor U12156 (N_12156,N_12081,N_12022);
and U12157 (N_12157,N_12012,N_12021);
nand U12158 (N_12158,N_12023,N_12105);
nor U12159 (N_12159,N_12088,N_12013);
and U12160 (N_12160,N_12083,N_12107);
or U12161 (N_12161,N_12009,N_12070);
and U12162 (N_12162,N_12121,N_12093);
nor U12163 (N_12163,N_12038,N_12087);
xnor U12164 (N_12164,N_12058,N_12046);
xnor U12165 (N_12165,N_12056,N_12114);
nand U12166 (N_12166,N_12047,N_12050);
xor U12167 (N_12167,N_12109,N_12116);
nand U12168 (N_12168,N_12037,N_12002);
nor U12169 (N_12169,N_12054,N_12059);
or U12170 (N_12170,N_12026,N_12112);
and U12171 (N_12171,N_12036,N_12015);
nor U12172 (N_12172,N_12014,N_12080);
or U12173 (N_12173,N_12006,N_12011);
xnor U12174 (N_12174,N_12040,N_12029);
or U12175 (N_12175,N_12110,N_12095);
or U12176 (N_12176,N_12051,N_12082);
and U12177 (N_12177,N_12000,N_12008);
or U12178 (N_12178,N_12025,N_12018);
nor U12179 (N_12179,N_12019,N_12001);
nand U12180 (N_12180,N_12039,N_12072);
nor U12181 (N_12181,N_12004,N_12104);
or U12182 (N_12182,N_12069,N_12007);
nor U12183 (N_12183,N_12068,N_12078);
or U12184 (N_12184,N_12074,N_12064);
xnor U12185 (N_12185,N_12076,N_12086);
nor U12186 (N_12186,N_12003,N_12120);
nand U12187 (N_12187,N_12124,N_12072);
nand U12188 (N_12188,N_12005,N_12051);
nand U12189 (N_12189,N_12089,N_12039);
xor U12190 (N_12190,N_12002,N_12110);
or U12191 (N_12191,N_12118,N_12037);
nand U12192 (N_12192,N_12097,N_12056);
nand U12193 (N_12193,N_12077,N_12045);
nor U12194 (N_12194,N_12070,N_12115);
nand U12195 (N_12195,N_12010,N_12005);
or U12196 (N_12196,N_12094,N_12028);
nand U12197 (N_12197,N_12059,N_12074);
or U12198 (N_12198,N_12014,N_12021);
xor U12199 (N_12199,N_12048,N_12004);
nand U12200 (N_12200,N_12076,N_12118);
and U12201 (N_12201,N_12103,N_12108);
nor U12202 (N_12202,N_12013,N_12033);
nand U12203 (N_12203,N_12122,N_12020);
xor U12204 (N_12204,N_12057,N_12021);
or U12205 (N_12205,N_12113,N_12014);
xor U12206 (N_12206,N_12068,N_12009);
or U12207 (N_12207,N_12075,N_12057);
nand U12208 (N_12208,N_12045,N_12070);
or U12209 (N_12209,N_12099,N_12076);
nor U12210 (N_12210,N_12064,N_12076);
or U12211 (N_12211,N_12040,N_12120);
or U12212 (N_12212,N_12055,N_12032);
and U12213 (N_12213,N_12070,N_12007);
nand U12214 (N_12214,N_12116,N_12009);
or U12215 (N_12215,N_12124,N_12046);
and U12216 (N_12216,N_12062,N_12086);
or U12217 (N_12217,N_12051,N_12069);
and U12218 (N_12218,N_12054,N_12093);
nor U12219 (N_12219,N_12046,N_12004);
or U12220 (N_12220,N_12028,N_12064);
xnor U12221 (N_12221,N_12006,N_12098);
or U12222 (N_12222,N_12093,N_12090);
or U12223 (N_12223,N_12002,N_12061);
nand U12224 (N_12224,N_12097,N_12030);
and U12225 (N_12225,N_12057,N_12080);
nor U12226 (N_12226,N_12052,N_12111);
and U12227 (N_12227,N_12025,N_12114);
nor U12228 (N_12228,N_12094,N_12026);
xnor U12229 (N_12229,N_12037,N_12040);
xor U12230 (N_12230,N_12059,N_12068);
or U12231 (N_12231,N_12059,N_12062);
nand U12232 (N_12232,N_12054,N_12024);
or U12233 (N_12233,N_12026,N_12058);
nand U12234 (N_12234,N_12038,N_12014);
nor U12235 (N_12235,N_12075,N_12055);
or U12236 (N_12236,N_12062,N_12013);
xor U12237 (N_12237,N_12063,N_12083);
nand U12238 (N_12238,N_12101,N_12111);
nor U12239 (N_12239,N_12043,N_12082);
or U12240 (N_12240,N_12063,N_12114);
or U12241 (N_12241,N_12048,N_12053);
nor U12242 (N_12242,N_12050,N_12090);
nand U12243 (N_12243,N_12009,N_12109);
or U12244 (N_12244,N_12029,N_12032);
xnor U12245 (N_12245,N_12068,N_12037);
xor U12246 (N_12246,N_12012,N_12121);
xnor U12247 (N_12247,N_12036,N_12070);
nand U12248 (N_12248,N_12061,N_12120);
and U12249 (N_12249,N_12032,N_12085);
and U12250 (N_12250,N_12206,N_12209);
xnor U12251 (N_12251,N_12174,N_12200);
nor U12252 (N_12252,N_12208,N_12203);
nand U12253 (N_12253,N_12218,N_12156);
and U12254 (N_12254,N_12213,N_12157);
and U12255 (N_12255,N_12211,N_12133);
xor U12256 (N_12256,N_12129,N_12226);
or U12257 (N_12257,N_12172,N_12222);
and U12258 (N_12258,N_12236,N_12233);
xor U12259 (N_12259,N_12215,N_12131);
and U12260 (N_12260,N_12194,N_12248);
or U12261 (N_12261,N_12212,N_12201);
nor U12262 (N_12262,N_12238,N_12242);
xor U12263 (N_12263,N_12240,N_12184);
nor U12264 (N_12264,N_12165,N_12160);
and U12265 (N_12265,N_12237,N_12126);
xor U12266 (N_12266,N_12158,N_12192);
nand U12267 (N_12267,N_12151,N_12163);
nor U12268 (N_12268,N_12169,N_12197);
or U12269 (N_12269,N_12199,N_12152);
nand U12270 (N_12270,N_12180,N_12159);
nand U12271 (N_12271,N_12128,N_12176);
xnor U12272 (N_12272,N_12140,N_12146);
nand U12273 (N_12273,N_12150,N_12216);
and U12274 (N_12274,N_12139,N_12135);
xnor U12275 (N_12275,N_12195,N_12182);
nor U12276 (N_12276,N_12220,N_12247);
or U12277 (N_12277,N_12223,N_12177);
and U12278 (N_12278,N_12205,N_12190);
nand U12279 (N_12279,N_12153,N_12170);
or U12280 (N_12280,N_12224,N_12125);
and U12281 (N_12281,N_12141,N_12186);
nand U12282 (N_12282,N_12245,N_12149);
nor U12283 (N_12283,N_12132,N_12171);
and U12284 (N_12284,N_12181,N_12228);
or U12285 (N_12285,N_12229,N_12243);
nand U12286 (N_12286,N_12227,N_12185);
xnor U12287 (N_12287,N_12217,N_12137);
and U12288 (N_12288,N_12127,N_12225);
xnor U12289 (N_12289,N_12178,N_12239);
nor U12290 (N_12290,N_12173,N_12134);
or U12291 (N_12291,N_12207,N_12179);
or U12292 (N_12292,N_12189,N_12167);
nor U12293 (N_12293,N_12161,N_12143);
or U12294 (N_12294,N_12144,N_12235);
or U12295 (N_12295,N_12234,N_12230);
xor U12296 (N_12296,N_12249,N_12241);
xnor U12297 (N_12297,N_12155,N_12130);
xor U12298 (N_12298,N_12142,N_12187);
xnor U12299 (N_12299,N_12221,N_12193);
or U12300 (N_12300,N_12198,N_12202);
xor U12301 (N_12301,N_12162,N_12188);
xor U12302 (N_12302,N_12214,N_12244);
nor U12303 (N_12303,N_12168,N_12166);
nor U12304 (N_12304,N_12196,N_12191);
and U12305 (N_12305,N_12175,N_12164);
nand U12306 (N_12306,N_12148,N_12219);
nor U12307 (N_12307,N_12136,N_12204);
nor U12308 (N_12308,N_12183,N_12145);
xor U12309 (N_12309,N_12231,N_12154);
and U12310 (N_12310,N_12210,N_12232);
or U12311 (N_12311,N_12246,N_12147);
xnor U12312 (N_12312,N_12138,N_12143);
or U12313 (N_12313,N_12218,N_12243);
nor U12314 (N_12314,N_12221,N_12177);
xnor U12315 (N_12315,N_12199,N_12177);
nor U12316 (N_12316,N_12232,N_12226);
nand U12317 (N_12317,N_12155,N_12205);
nor U12318 (N_12318,N_12155,N_12158);
or U12319 (N_12319,N_12190,N_12228);
and U12320 (N_12320,N_12230,N_12144);
xnor U12321 (N_12321,N_12209,N_12199);
xor U12322 (N_12322,N_12222,N_12139);
or U12323 (N_12323,N_12242,N_12216);
nand U12324 (N_12324,N_12197,N_12134);
nand U12325 (N_12325,N_12197,N_12244);
or U12326 (N_12326,N_12233,N_12179);
and U12327 (N_12327,N_12203,N_12210);
xor U12328 (N_12328,N_12187,N_12158);
and U12329 (N_12329,N_12167,N_12239);
and U12330 (N_12330,N_12140,N_12241);
nand U12331 (N_12331,N_12168,N_12228);
nand U12332 (N_12332,N_12155,N_12190);
or U12333 (N_12333,N_12243,N_12176);
nor U12334 (N_12334,N_12227,N_12147);
nor U12335 (N_12335,N_12182,N_12203);
and U12336 (N_12336,N_12142,N_12139);
and U12337 (N_12337,N_12177,N_12228);
or U12338 (N_12338,N_12165,N_12137);
xnor U12339 (N_12339,N_12209,N_12246);
xor U12340 (N_12340,N_12161,N_12165);
nor U12341 (N_12341,N_12130,N_12236);
xnor U12342 (N_12342,N_12134,N_12186);
xnor U12343 (N_12343,N_12132,N_12182);
nor U12344 (N_12344,N_12150,N_12144);
and U12345 (N_12345,N_12139,N_12244);
and U12346 (N_12346,N_12170,N_12234);
nand U12347 (N_12347,N_12246,N_12154);
xor U12348 (N_12348,N_12188,N_12143);
or U12349 (N_12349,N_12201,N_12141);
or U12350 (N_12350,N_12157,N_12163);
nand U12351 (N_12351,N_12140,N_12170);
and U12352 (N_12352,N_12177,N_12178);
and U12353 (N_12353,N_12125,N_12245);
xnor U12354 (N_12354,N_12182,N_12202);
nand U12355 (N_12355,N_12162,N_12217);
or U12356 (N_12356,N_12128,N_12192);
nor U12357 (N_12357,N_12229,N_12246);
nor U12358 (N_12358,N_12210,N_12188);
nand U12359 (N_12359,N_12207,N_12243);
xor U12360 (N_12360,N_12215,N_12246);
and U12361 (N_12361,N_12184,N_12145);
nand U12362 (N_12362,N_12208,N_12211);
nand U12363 (N_12363,N_12203,N_12205);
nand U12364 (N_12364,N_12170,N_12214);
or U12365 (N_12365,N_12134,N_12167);
and U12366 (N_12366,N_12167,N_12200);
nand U12367 (N_12367,N_12246,N_12165);
xnor U12368 (N_12368,N_12213,N_12214);
or U12369 (N_12369,N_12180,N_12170);
xor U12370 (N_12370,N_12188,N_12198);
nor U12371 (N_12371,N_12191,N_12134);
nand U12372 (N_12372,N_12201,N_12214);
or U12373 (N_12373,N_12214,N_12132);
and U12374 (N_12374,N_12156,N_12249);
nor U12375 (N_12375,N_12347,N_12334);
nand U12376 (N_12376,N_12348,N_12311);
or U12377 (N_12377,N_12291,N_12270);
or U12378 (N_12378,N_12276,N_12321);
or U12379 (N_12379,N_12329,N_12349);
and U12380 (N_12380,N_12343,N_12350);
or U12381 (N_12381,N_12274,N_12259);
nor U12382 (N_12382,N_12360,N_12286);
xnor U12383 (N_12383,N_12332,N_12325);
or U12384 (N_12384,N_12331,N_12372);
xor U12385 (N_12385,N_12359,N_12313);
nand U12386 (N_12386,N_12341,N_12269);
xor U12387 (N_12387,N_12322,N_12361);
nand U12388 (N_12388,N_12336,N_12305);
nor U12389 (N_12389,N_12346,N_12292);
or U12390 (N_12390,N_12275,N_12309);
xor U12391 (N_12391,N_12271,N_12354);
or U12392 (N_12392,N_12287,N_12339);
and U12393 (N_12393,N_12253,N_12315);
or U12394 (N_12394,N_12307,N_12316);
nand U12395 (N_12395,N_12318,N_12333);
and U12396 (N_12396,N_12280,N_12289);
nand U12397 (N_12397,N_12299,N_12371);
nor U12398 (N_12398,N_12262,N_12258);
or U12399 (N_12399,N_12277,N_12370);
and U12400 (N_12400,N_12282,N_12351);
and U12401 (N_12401,N_12319,N_12368);
and U12402 (N_12402,N_12327,N_12310);
and U12403 (N_12403,N_12363,N_12297);
nor U12404 (N_12404,N_12254,N_12304);
nor U12405 (N_12405,N_12364,N_12251);
nand U12406 (N_12406,N_12358,N_12278);
nand U12407 (N_12407,N_12308,N_12296);
xnor U12408 (N_12408,N_12335,N_12314);
xnor U12409 (N_12409,N_12303,N_12353);
xnor U12410 (N_12410,N_12365,N_12300);
xor U12411 (N_12411,N_12272,N_12281);
nor U12412 (N_12412,N_12317,N_12298);
nor U12413 (N_12413,N_12340,N_12279);
nand U12414 (N_12414,N_12356,N_12273);
and U12415 (N_12415,N_12284,N_12302);
or U12416 (N_12416,N_12366,N_12344);
or U12417 (N_12417,N_12267,N_12330);
or U12418 (N_12418,N_12369,N_12295);
and U12419 (N_12419,N_12337,N_12345);
nor U12420 (N_12420,N_12268,N_12362);
xnor U12421 (N_12421,N_12288,N_12257);
nand U12422 (N_12422,N_12261,N_12252);
nand U12423 (N_12423,N_12293,N_12264);
or U12424 (N_12424,N_12357,N_12290);
or U12425 (N_12425,N_12367,N_12328);
nor U12426 (N_12426,N_12373,N_12320);
and U12427 (N_12427,N_12260,N_12324);
nor U12428 (N_12428,N_12285,N_12326);
nor U12429 (N_12429,N_12342,N_12250);
nor U12430 (N_12430,N_12294,N_12323);
or U12431 (N_12431,N_12256,N_12283);
nand U12432 (N_12432,N_12265,N_12355);
nor U12433 (N_12433,N_12312,N_12266);
nor U12434 (N_12434,N_12352,N_12338);
or U12435 (N_12435,N_12263,N_12306);
and U12436 (N_12436,N_12301,N_12374);
or U12437 (N_12437,N_12255,N_12337);
nand U12438 (N_12438,N_12298,N_12274);
nand U12439 (N_12439,N_12261,N_12255);
nand U12440 (N_12440,N_12295,N_12309);
nand U12441 (N_12441,N_12321,N_12275);
nand U12442 (N_12442,N_12287,N_12281);
nand U12443 (N_12443,N_12310,N_12305);
or U12444 (N_12444,N_12278,N_12365);
or U12445 (N_12445,N_12294,N_12264);
or U12446 (N_12446,N_12330,N_12349);
nor U12447 (N_12447,N_12315,N_12325);
and U12448 (N_12448,N_12253,N_12297);
nor U12449 (N_12449,N_12342,N_12307);
and U12450 (N_12450,N_12285,N_12329);
xnor U12451 (N_12451,N_12338,N_12370);
and U12452 (N_12452,N_12269,N_12288);
and U12453 (N_12453,N_12285,N_12258);
and U12454 (N_12454,N_12337,N_12350);
xor U12455 (N_12455,N_12356,N_12261);
nor U12456 (N_12456,N_12364,N_12278);
and U12457 (N_12457,N_12304,N_12333);
or U12458 (N_12458,N_12312,N_12320);
nand U12459 (N_12459,N_12337,N_12368);
xnor U12460 (N_12460,N_12254,N_12269);
nand U12461 (N_12461,N_12350,N_12267);
and U12462 (N_12462,N_12345,N_12374);
xor U12463 (N_12463,N_12344,N_12319);
nor U12464 (N_12464,N_12323,N_12366);
or U12465 (N_12465,N_12250,N_12341);
or U12466 (N_12466,N_12300,N_12316);
nand U12467 (N_12467,N_12276,N_12338);
or U12468 (N_12468,N_12252,N_12373);
nor U12469 (N_12469,N_12360,N_12269);
nand U12470 (N_12470,N_12346,N_12294);
nor U12471 (N_12471,N_12363,N_12373);
nand U12472 (N_12472,N_12330,N_12366);
or U12473 (N_12473,N_12302,N_12251);
nand U12474 (N_12474,N_12259,N_12340);
xnor U12475 (N_12475,N_12281,N_12340);
xnor U12476 (N_12476,N_12269,N_12259);
nor U12477 (N_12477,N_12347,N_12285);
nor U12478 (N_12478,N_12324,N_12261);
or U12479 (N_12479,N_12319,N_12279);
or U12480 (N_12480,N_12278,N_12263);
xnor U12481 (N_12481,N_12282,N_12256);
or U12482 (N_12482,N_12277,N_12253);
xnor U12483 (N_12483,N_12264,N_12265);
nor U12484 (N_12484,N_12287,N_12343);
or U12485 (N_12485,N_12271,N_12311);
or U12486 (N_12486,N_12290,N_12358);
or U12487 (N_12487,N_12355,N_12262);
nor U12488 (N_12488,N_12311,N_12365);
nor U12489 (N_12489,N_12315,N_12357);
or U12490 (N_12490,N_12372,N_12351);
and U12491 (N_12491,N_12290,N_12263);
and U12492 (N_12492,N_12370,N_12324);
nor U12493 (N_12493,N_12318,N_12326);
xnor U12494 (N_12494,N_12285,N_12283);
and U12495 (N_12495,N_12313,N_12335);
nor U12496 (N_12496,N_12286,N_12344);
and U12497 (N_12497,N_12270,N_12293);
nor U12498 (N_12498,N_12305,N_12328);
xnor U12499 (N_12499,N_12329,N_12338);
xnor U12500 (N_12500,N_12444,N_12378);
nand U12501 (N_12501,N_12416,N_12470);
nor U12502 (N_12502,N_12490,N_12462);
nor U12503 (N_12503,N_12398,N_12382);
xor U12504 (N_12504,N_12432,N_12385);
nor U12505 (N_12505,N_12376,N_12492);
xnor U12506 (N_12506,N_12498,N_12406);
nand U12507 (N_12507,N_12387,N_12471);
or U12508 (N_12508,N_12409,N_12390);
xor U12509 (N_12509,N_12399,N_12453);
nand U12510 (N_12510,N_12389,N_12461);
xnor U12511 (N_12511,N_12386,N_12473);
and U12512 (N_12512,N_12428,N_12481);
or U12513 (N_12513,N_12417,N_12475);
nand U12514 (N_12514,N_12383,N_12419);
and U12515 (N_12515,N_12426,N_12442);
and U12516 (N_12516,N_12430,N_12452);
xor U12517 (N_12517,N_12435,N_12379);
or U12518 (N_12518,N_12451,N_12381);
xor U12519 (N_12519,N_12384,N_12445);
xor U12520 (N_12520,N_12469,N_12413);
xor U12521 (N_12521,N_12395,N_12410);
nand U12522 (N_12522,N_12496,N_12418);
xor U12523 (N_12523,N_12429,N_12438);
and U12524 (N_12524,N_12495,N_12479);
and U12525 (N_12525,N_12474,N_12472);
or U12526 (N_12526,N_12491,N_12478);
and U12527 (N_12527,N_12392,N_12436);
nand U12528 (N_12528,N_12402,N_12441);
xnor U12529 (N_12529,N_12465,N_12454);
or U12530 (N_12530,N_12412,N_12487);
nand U12531 (N_12531,N_12424,N_12422);
and U12532 (N_12532,N_12476,N_12407);
or U12533 (N_12533,N_12403,N_12457);
xnor U12534 (N_12534,N_12391,N_12466);
or U12535 (N_12535,N_12425,N_12464);
xnor U12536 (N_12536,N_12468,N_12421);
nand U12537 (N_12537,N_12408,N_12477);
and U12538 (N_12538,N_12482,N_12443);
nand U12539 (N_12539,N_12448,N_12447);
and U12540 (N_12540,N_12460,N_12439);
or U12541 (N_12541,N_12420,N_12393);
or U12542 (N_12542,N_12411,N_12437);
nand U12543 (N_12543,N_12450,N_12404);
nor U12544 (N_12544,N_12488,N_12449);
xnor U12545 (N_12545,N_12458,N_12377);
nor U12546 (N_12546,N_12380,N_12415);
nor U12547 (N_12547,N_12401,N_12483);
nor U12548 (N_12548,N_12427,N_12486);
or U12549 (N_12549,N_12485,N_12440);
nor U12550 (N_12550,N_12463,N_12394);
nor U12551 (N_12551,N_12497,N_12388);
nor U12552 (N_12552,N_12499,N_12489);
and U12553 (N_12553,N_12493,N_12480);
xor U12554 (N_12554,N_12467,N_12456);
and U12555 (N_12555,N_12423,N_12414);
or U12556 (N_12556,N_12396,N_12494);
xnor U12557 (N_12557,N_12375,N_12433);
and U12558 (N_12558,N_12405,N_12431);
nor U12559 (N_12559,N_12455,N_12446);
and U12560 (N_12560,N_12397,N_12400);
nand U12561 (N_12561,N_12484,N_12459);
xnor U12562 (N_12562,N_12434,N_12413);
and U12563 (N_12563,N_12426,N_12412);
xor U12564 (N_12564,N_12467,N_12465);
xor U12565 (N_12565,N_12404,N_12474);
nand U12566 (N_12566,N_12495,N_12395);
and U12567 (N_12567,N_12420,N_12471);
nand U12568 (N_12568,N_12418,N_12450);
or U12569 (N_12569,N_12484,N_12489);
and U12570 (N_12570,N_12381,N_12467);
xor U12571 (N_12571,N_12375,N_12450);
or U12572 (N_12572,N_12440,N_12457);
nand U12573 (N_12573,N_12397,N_12410);
xor U12574 (N_12574,N_12443,N_12428);
or U12575 (N_12575,N_12476,N_12383);
xor U12576 (N_12576,N_12390,N_12422);
xor U12577 (N_12577,N_12470,N_12435);
xor U12578 (N_12578,N_12455,N_12424);
nor U12579 (N_12579,N_12413,N_12435);
nor U12580 (N_12580,N_12411,N_12480);
and U12581 (N_12581,N_12453,N_12459);
and U12582 (N_12582,N_12397,N_12491);
xor U12583 (N_12583,N_12410,N_12459);
or U12584 (N_12584,N_12437,N_12488);
or U12585 (N_12585,N_12456,N_12441);
or U12586 (N_12586,N_12420,N_12466);
nor U12587 (N_12587,N_12480,N_12479);
xnor U12588 (N_12588,N_12411,N_12430);
nand U12589 (N_12589,N_12418,N_12386);
and U12590 (N_12590,N_12412,N_12429);
nor U12591 (N_12591,N_12473,N_12474);
nand U12592 (N_12592,N_12496,N_12381);
xnor U12593 (N_12593,N_12440,N_12479);
or U12594 (N_12594,N_12432,N_12384);
or U12595 (N_12595,N_12440,N_12445);
nand U12596 (N_12596,N_12496,N_12455);
and U12597 (N_12597,N_12426,N_12468);
nor U12598 (N_12598,N_12467,N_12426);
or U12599 (N_12599,N_12467,N_12413);
nand U12600 (N_12600,N_12396,N_12425);
xor U12601 (N_12601,N_12444,N_12387);
or U12602 (N_12602,N_12444,N_12476);
or U12603 (N_12603,N_12447,N_12382);
nand U12604 (N_12604,N_12485,N_12477);
or U12605 (N_12605,N_12413,N_12394);
and U12606 (N_12606,N_12457,N_12377);
or U12607 (N_12607,N_12425,N_12424);
nor U12608 (N_12608,N_12418,N_12456);
and U12609 (N_12609,N_12415,N_12462);
nand U12610 (N_12610,N_12404,N_12380);
and U12611 (N_12611,N_12413,N_12401);
nand U12612 (N_12612,N_12403,N_12392);
xnor U12613 (N_12613,N_12407,N_12381);
or U12614 (N_12614,N_12478,N_12390);
xnor U12615 (N_12615,N_12386,N_12495);
nor U12616 (N_12616,N_12458,N_12493);
nor U12617 (N_12617,N_12453,N_12492);
and U12618 (N_12618,N_12421,N_12392);
nand U12619 (N_12619,N_12491,N_12408);
nor U12620 (N_12620,N_12401,N_12391);
or U12621 (N_12621,N_12485,N_12428);
and U12622 (N_12622,N_12418,N_12381);
nand U12623 (N_12623,N_12454,N_12410);
or U12624 (N_12624,N_12451,N_12446);
or U12625 (N_12625,N_12579,N_12601);
nand U12626 (N_12626,N_12507,N_12534);
nor U12627 (N_12627,N_12506,N_12580);
nor U12628 (N_12628,N_12541,N_12508);
or U12629 (N_12629,N_12581,N_12538);
nor U12630 (N_12630,N_12607,N_12609);
and U12631 (N_12631,N_12519,N_12553);
xnor U12632 (N_12632,N_12582,N_12585);
or U12633 (N_12633,N_12610,N_12563);
or U12634 (N_12634,N_12559,N_12592);
nand U12635 (N_12635,N_12540,N_12603);
xnor U12636 (N_12636,N_12526,N_12532);
nor U12637 (N_12637,N_12522,N_12557);
xnor U12638 (N_12638,N_12588,N_12567);
or U12639 (N_12639,N_12566,N_12548);
and U12640 (N_12640,N_12578,N_12516);
xor U12641 (N_12641,N_12536,N_12593);
nor U12642 (N_12642,N_12562,N_12568);
nand U12643 (N_12643,N_12544,N_12509);
xor U12644 (N_12644,N_12621,N_12556);
xor U12645 (N_12645,N_12546,N_12620);
and U12646 (N_12646,N_12596,N_12503);
and U12647 (N_12647,N_12612,N_12615);
or U12648 (N_12648,N_12515,N_12616);
and U12649 (N_12649,N_12552,N_12576);
nand U12650 (N_12650,N_12511,N_12598);
or U12651 (N_12651,N_12569,N_12602);
nor U12652 (N_12652,N_12575,N_12524);
and U12653 (N_12653,N_12586,N_12547);
nor U12654 (N_12654,N_12600,N_12517);
nor U12655 (N_12655,N_12611,N_12565);
and U12656 (N_12656,N_12590,N_12520);
nand U12657 (N_12657,N_12500,N_12624);
and U12658 (N_12658,N_12613,N_12525);
nand U12659 (N_12659,N_12549,N_12622);
and U12660 (N_12660,N_12571,N_12554);
xor U12661 (N_12661,N_12597,N_12619);
and U12662 (N_12662,N_12574,N_12539);
xnor U12663 (N_12663,N_12533,N_12583);
and U12664 (N_12664,N_12617,N_12555);
or U12665 (N_12665,N_12564,N_12573);
and U12666 (N_12666,N_12606,N_12595);
and U12667 (N_12667,N_12528,N_12543);
xnor U12668 (N_12668,N_12584,N_12504);
and U12669 (N_12669,N_12542,N_12608);
xor U12670 (N_12670,N_12513,N_12614);
nor U12671 (N_12671,N_12550,N_12587);
nand U12672 (N_12672,N_12545,N_12604);
nor U12673 (N_12673,N_12502,N_12510);
xor U12674 (N_12674,N_12514,N_12589);
or U12675 (N_12675,N_12623,N_12530);
or U12676 (N_12676,N_12605,N_12505);
and U12677 (N_12677,N_12523,N_12561);
or U12678 (N_12678,N_12572,N_12560);
nor U12679 (N_12679,N_12512,N_12529);
and U12680 (N_12680,N_12521,N_12531);
nand U12681 (N_12681,N_12518,N_12551);
xnor U12682 (N_12682,N_12570,N_12501);
and U12683 (N_12683,N_12527,N_12591);
nor U12684 (N_12684,N_12535,N_12594);
and U12685 (N_12685,N_12558,N_12618);
nand U12686 (N_12686,N_12599,N_12577);
xor U12687 (N_12687,N_12537,N_12524);
nand U12688 (N_12688,N_12535,N_12561);
nor U12689 (N_12689,N_12521,N_12502);
xor U12690 (N_12690,N_12555,N_12522);
or U12691 (N_12691,N_12500,N_12583);
and U12692 (N_12692,N_12552,N_12594);
nor U12693 (N_12693,N_12614,N_12512);
nor U12694 (N_12694,N_12573,N_12620);
xor U12695 (N_12695,N_12521,N_12533);
nor U12696 (N_12696,N_12606,N_12553);
or U12697 (N_12697,N_12562,N_12559);
nor U12698 (N_12698,N_12574,N_12514);
and U12699 (N_12699,N_12531,N_12539);
or U12700 (N_12700,N_12588,N_12592);
nor U12701 (N_12701,N_12542,N_12598);
or U12702 (N_12702,N_12591,N_12511);
nor U12703 (N_12703,N_12562,N_12598);
and U12704 (N_12704,N_12530,N_12598);
xnor U12705 (N_12705,N_12595,N_12592);
nand U12706 (N_12706,N_12500,N_12600);
nand U12707 (N_12707,N_12559,N_12595);
nand U12708 (N_12708,N_12556,N_12540);
nor U12709 (N_12709,N_12560,N_12518);
xor U12710 (N_12710,N_12525,N_12606);
and U12711 (N_12711,N_12509,N_12604);
or U12712 (N_12712,N_12595,N_12545);
nand U12713 (N_12713,N_12566,N_12510);
nand U12714 (N_12714,N_12595,N_12512);
nand U12715 (N_12715,N_12503,N_12509);
or U12716 (N_12716,N_12612,N_12537);
or U12717 (N_12717,N_12577,N_12613);
or U12718 (N_12718,N_12540,N_12529);
and U12719 (N_12719,N_12526,N_12611);
or U12720 (N_12720,N_12597,N_12560);
and U12721 (N_12721,N_12591,N_12620);
and U12722 (N_12722,N_12560,N_12603);
and U12723 (N_12723,N_12621,N_12528);
xnor U12724 (N_12724,N_12618,N_12514);
and U12725 (N_12725,N_12561,N_12585);
xnor U12726 (N_12726,N_12619,N_12574);
and U12727 (N_12727,N_12504,N_12503);
and U12728 (N_12728,N_12607,N_12611);
xnor U12729 (N_12729,N_12620,N_12503);
and U12730 (N_12730,N_12521,N_12596);
nor U12731 (N_12731,N_12589,N_12608);
nand U12732 (N_12732,N_12577,N_12513);
xor U12733 (N_12733,N_12612,N_12502);
or U12734 (N_12734,N_12515,N_12564);
and U12735 (N_12735,N_12521,N_12585);
and U12736 (N_12736,N_12601,N_12573);
nand U12737 (N_12737,N_12538,N_12610);
xor U12738 (N_12738,N_12612,N_12594);
and U12739 (N_12739,N_12568,N_12583);
nor U12740 (N_12740,N_12618,N_12521);
nand U12741 (N_12741,N_12591,N_12622);
nor U12742 (N_12742,N_12620,N_12537);
xnor U12743 (N_12743,N_12566,N_12553);
xnor U12744 (N_12744,N_12512,N_12514);
nand U12745 (N_12745,N_12506,N_12592);
and U12746 (N_12746,N_12560,N_12623);
nand U12747 (N_12747,N_12524,N_12590);
and U12748 (N_12748,N_12508,N_12515);
nor U12749 (N_12749,N_12501,N_12507);
nand U12750 (N_12750,N_12717,N_12728);
or U12751 (N_12751,N_12678,N_12643);
and U12752 (N_12752,N_12733,N_12682);
nand U12753 (N_12753,N_12710,N_12732);
xor U12754 (N_12754,N_12741,N_12671);
and U12755 (N_12755,N_12680,N_12684);
nand U12756 (N_12756,N_12725,N_12743);
nand U12757 (N_12757,N_12652,N_12727);
and U12758 (N_12758,N_12746,N_12683);
or U12759 (N_12759,N_12676,N_12674);
nor U12760 (N_12760,N_12657,N_12706);
nor U12761 (N_12761,N_12644,N_12631);
and U12762 (N_12762,N_12735,N_12662);
nand U12763 (N_12763,N_12688,N_12632);
or U12764 (N_12764,N_12726,N_12707);
nand U12765 (N_12765,N_12656,N_12705);
xnor U12766 (N_12766,N_12627,N_12698);
xor U12767 (N_12767,N_12679,N_12700);
or U12768 (N_12768,N_12711,N_12668);
and U12769 (N_12769,N_12691,N_12740);
nand U12770 (N_12770,N_12670,N_12712);
and U12771 (N_12771,N_12692,N_12695);
xnor U12772 (N_12772,N_12709,N_12738);
nor U12773 (N_12773,N_12666,N_12690);
xor U12774 (N_12774,N_12655,N_12730);
xnor U12775 (N_12775,N_12630,N_12633);
or U12776 (N_12776,N_12659,N_12653);
and U12777 (N_12777,N_12639,N_12689);
nor U12778 (N_12778,N_12686,N_12637);
nor U12779 (N_12779,N_12703,N_12723);
xnor U12780 (N_12780,N_12747,N_12714);
nand U12781 (N_12781,N_12685,N_12636);
xor U12782 (N_12782,N_12693,N_12696);
nand U12783 (N_12783,N_12677,N_12658);
or U12784 (N_12784,N_12716,N_12654);
or U12785 (N_12785,N_12661,N_12675);
and U12786 (N_12786,N_12708,N_12737);
or U12787 (N_12787,N_12651,N_12642);
nor U12788 (N_12788,N_12646,N_12650);
nand U12789 (N_12789,N_12699,N_12739);
nand U12790 (N_12790,N_12672,N_12720);
and U12791 (N_12791,N_12629,N_12634);
or U12792 (N_12792,N_12640,N_12664);
nor U12793 (N_12793,N_12649,N_12702);
xnor U12794 (N_12794,N_12718,N_12744);
or U12795 (N_12795,N_12748,N_12715);
nor U12796 (N_12796,N_12729,N_12638);
xnor U12797 (N_12797,N_12694,N_12734);
or U12798 (N_12798,N_12669,N_12681);
nor U12799 (N_12799,N_12687,N_12635);
or U12800 (N_12800,N_12673,N_12724);
or U12801 (N_12801,N_12660,N_12665);
or U12802 (N_12802,N_12749,N_12628);
nor U12803 (N_12803,N_12736,N_12645);
nor U12804 (N_12804,N_12713,N_12745);
nand U12805 (N_12805,N_12625,N_12721);
xor U12806 (N_12806,N_12641,N_12719);
or U12807 (N_12807,N_12701,N_12626);
nand U12808 (N_12808,N_12704,N_12663);
nand U12809 (N_12809,N_12667,N_12697);
and U12810 (N_12810,N_12648,N_12722);
and U12811 (N_12811,N_12742,N_12731);
and U12812 (N_12812,N_12647,N_12718);
xnor U12813 (N_12813,N_12695,N_12641);
nor U12814 (N_12814,N_12634,N_12660);
and U12815 (N_12815,N_12702,N_12642);
or U12816 (N_12816,N_12674,N_12747);
or U12817 (N_12817,N_12636,N_12724);
nand U12818 (N_12818,N_12727,N_12648);
and U12819 (N_12819,N_12665,N_12672);
nand U12820 (N_12820,N_12732,N_12632);
xor U12821 (N_12821,N_12734,N_12741);
nand U12822 (N_12822,N_12739,N_12697);
or U12823 (N_12823,N_12626,N_12727);
nor U12824 (N_12824,N_12635,N_12677);
xor U12825 (N_12825,N_12629,N_12648);
nand U12826 (N_12826,N_12657,N_12729);
nor U12827 (N_12827,N_12625,N_12726);
and U12828 (N_12828,N_12747,N_12658);
xor U12829 (N_12829,N_12639,N_12633);
nor U12830 (N_12830,N_12706,N_12745);
xor U12831 (N_12831,N_12675,N_12709);
and U12832 (N_12832,N_12727,N_12662);
or U12833 (N_12833,N_12744,N_12675);
or U12834 (N_12834,N_12652,N_12670);
xnor U12835 (N_12835,N_12724,N_12653);
and U12836 (N_12836,N_12692,N_12687);
and U12837 (N_12837,N_12633,N_12677);
nand U12838 (N_12838,N_12687,N_12703);
or U12839 (N_12839,N_12634,N_12648);
xnor U12840 (N_12840,N_12718,N_12726);
and U12841 (N_12841,N_12736,N_12749);
and U12842 (N_12842,N_12714,N_12701);
nor U12843 (N_12843,N_12723,N_12632);
nand U12844 (N_12844,N_12654,N_12692);
nor U12845 (N_12845,N_12647,N_12662);
or U12846 (N_12846,N_12708,N_12633);
or U12847 (N_12847,N_12646,N_12748);
and U12848 (N_12848,N_12680,N_12695);
nor U12849 (N_12849,N_12721,N_12676);
nor U12850 (N_12850,N_12745,N_12655);
nand U12851 (N_12851,N_12688,N_12650);
nand U12852 (N_12852,N_12714,N_12654);
nand U12853 (N_12853,N_12712,N_12659);
or U12854 (N_12854,N_12732,N_12678);
nand U12855 (N_12855,N_12713,N_12642);
nor U12856 (N_12856,N_12705,N_12716);
xnor U12857 (N_12857,N_12715,N_12717);
nand U12858 (N_12858,N_12674,N_12660);
xor U12859 (N_12859,N_12713,N_12653);
nor U12860 (N_12860,N_12660,N_12652);
xnor U12861 (N_12861,N_12716,N_12739);
nand U12862 (N_12862,N_12645,N_12698);
or U12863 (N_12863,N_12683,N_12679);
xor U12864 (N_12864,N_12705,N_12647);
nand U12865 (N_12865,N_12687,N_12735);
nor U12866 (N_12866,N_12728,N_12637);
nor U12867 (N_12867,N_12726,N_12641);
xnor U12868 (N_12868,N_12710,N_12650);
xnor U12869 (N_12869,N_12654,N_12696);
or U12870 (N_12870,N_12655,N_12679);
xnor U12871 (N_12871,N_12640,N_12625);
or U12872 (N_12872,N_12647,N_12691);
nand U12873 (N_12873,N_12669,N_12683);
xnor U12874 (N_12874,N_12661,N_12635);
or U12875 (N_12875,N_12778,N_12768);
nand U12876 (N_12876,N_12751,N_12769);
and U12877 (N_12877,N_12805,N_12854);
nand U12878 (N_12878,N_12796,N_12818);
and U12879 (N_12879,N_12771,N_12766);
nor U12880 (N_12880,N_12853,N_12832);
nor U12881 (N_12881,N_12824,N_12781);
nor U12882 (N_12882,N_12812,N_12865);
nand U12883 (N_12883,N_12844,N_12803);
and U12884 (N_12884,N_12850,N_12775);
xnor U12885 (N_12885,N_12780,N_12794);
nand U12886 (N_12886,N_12787,N_12756);
nand U12887 (N_12887,N_12856,N_12867);
or U12888 (N_12888,N_12862,N_12785);
and U12889 (N_12889,N_12870,N_12762);
nand U12890 (N_12890,N_12842,N_12814);
nor U12891 (N_12891,N_12852,N_12791);
nand U12892 (N_12892,N_12855,N_12829);
and U12893 (N_12893,N_12828,N_12871);
nand U12894 (N_12894,N_12831,N_12765);
xnor U12895 (N_12895,N_12807,N_12767);
and U12896 (N_12896,N_12763,N_12868);
nor U12897 (N_12897,N_12806,N_12817);
and U12898 (N_12898,N_12863,N_12802);
nand U12899 (N_12899,N_12754,N_12822);
nand U12900 (N_12900,N_12782,N_12873);
and U12901 (N_12901,N_12793,N_12825);
xor U12902 (N_12902,N_12797,N_12869);
or U12903 (N_12903,N_12760,N_12774);
and U12904 (N_12904,N_12815,N_12821);
nor U12905 (N_12905,N_12776,N_12819);
or U12906 (N_12906,N_12859,N_12837);
xnor U12907 (N_12907,N_12777,N_12752);
and U12908 (N_12908,N_12835,N_12798);
and U12909 (N_12909,N_12833,N_12788);
and U12910 (N_12910,N_12857,N_12847);
or U12911 (N_12911,N_12841,N_12866);
nor U12912 (N_12912,N_12840,N_12753);
nor U12913 (N_12913,N_12848,N_12826);
and U12914 (N_12914,N_12845,N_12830);
nor U12915 (N_12915,N_12864,N_12811);
nor U12916 (N_12916,N_12799,N_12757);
nand U12917 (N_12917,N_12820,N_12851);
nor U12918 (N_12918,N_12772,N_12810);
nand U12919 (N_12919,N_12801,N_12784);
nor U12920 (N_12920,N_12761,N_12846);
nand U12921 (N_12921,N_12860,N_12816);
nor U12922 (N_12922,N_12790,N_12843);
nand U12923 (N_12923,N_12795,N_12786);
nand U12924 (N_12924,N_12792,N_12849);
or U12925 (N_12925,N_12823,N_12759);
nand U12926 (N_12926,N_12874,N_12808);
or U12927 (N_12927,N_12755,N_12804);
and U12928 (N_12928,N_12827,N_12872);
xor U12929 (N_12929,N_12783,N_12764);
xnor U12930 (N_12930,N_12858,N_12813);
nand U12931 (N_12931,N_12758,N_12789);
nor U12932 (N_12932,N_12861,N_12770);
nor U12933 (N_12933,N_12839,N_12779);
nor U12934 (N_12934,N_12836,N_12750);
nor U12935 (N_12935,N_12773,N_12809);
and U12936 (N_12936,N_12834,N_12800);
nand U12937 (N_12937,N_12838,N_12757);
nor U12938 (N_12938,N_12870,N_12824);
nor U12939 (N_12939,N_12859,N_12758);
nand U12940 (N_12940,N_12776,N_12865);
nor U12941 (N_12941,N_12816,N_12762);
and U12942 (N_12942,N_12802,N_12852);
nor U12943 (N_12943,N_12850,N_12782);
xor U12944 (N_12944,N_12817,N_12767);
and U12945 (N_12945,N_12786,N_12861);
nand U12946 (N_12946,N_12815,N_12811);
xor U12947 (N_12947,N_12798,N_12847);
nor U12948 (N_12948,N_12777,N_12780);
nand U12949 (N_12949,N_12769,N_12801);
or U12950 (N_12950,N_12865,N_12869);
xor U12951 (N_12951,N_12793,N_12781);
nor U12952 (N_12952,N_12830,N_12866);
xor U12953 (N_12953,N_12842,N_12771);
xor U12954 (N_12954,N_12781,N_12791);
nor U12955 (N_12955,N_12776,N_12784);
nand U12956 (N_12956,N_12769,N_12773);
nor U12957 (N_12957,N_12776,N_12832);
or U12958 (N_12958,N_12806,N_12764);
xor U12959 (N_12959,N_12785,N_12861);
nor U12960 (N_12960,N_12752,N_12764);
xnor U12961 (N_12961,N_12794,N_12856);
nor U12962 (N_12962,N_12768,N_12780);
nor U12963 (N_12963,N_12822,N_12855);
or U12964 (N_12964,N_12845,N_12823);
or U12965 (N_12965,N_12868,N_12825);
nor U12966 (N_12966,N_12760,N_12812);
xnor U12967 (N_12967,N_12872,N_12769);
and U12968 (N_12968,N_12821,N_12798);
and U12969 (N_12969,N_12798,N_12819);
and U12970 (N_12970,N_12784,N_12866);
or U12971 (N_12971,N_12857,N_12819);
or U12972 (N_12972,N_12820,N_12872);
and U12973 (N_12973,N_12871,N_12777);
xnor U12974 (N_12974,N_12840,N_12854);
and U12975 (N_12975,N_12841,N_12853);
or U12976 (N_12976,N_12763,N_12760);
nor U12977 (N_12977,N_12770,N_12808);
nor U12978 (N_12978,N_12814,N_12849);
and U12979 (N_12979,N_12861,N_12766);
nand U12980 (N_12980,N_12780,N_12751);
nand U12981 (N_12981,N_12851,N_12807);
nor U12982 (N_12982,N_12753,N_12812);
xnor U12983 (N_12983,N_12820,N_12817);
and U12984 (N_12984,N_12817,N_12799);
and U12985 (N_12985,N_12753,N_12788);
and U12986 (N_12986,N_12777,N_12755);
and U12987 (N_12987,N_12788,N_12782);
xor U12988 (N_12988,N_12836,N_12856);
xnor U12989 (N_12989,N_12752,N_12823);
nand U12990 (N_12990,N_12751,N_12850);
or U12991 (N_12991,N_12792,N_12798);
xor U12992 (N_12992,N_12833,N_12821);
nor U12993 (N_12993,N_12823,N_12866);
xnor U12994 (N_12994,N_12819,N_12859);
nand U12995 (N_12995,N_12824,N_12853);
or U12996 (N_12996,N_12796,N_12757);
xnor U12997 (N_12997,N_12857,N_12785);
nand U12998 (N_12998,N_12800,N_12868);
or U12999 (N_12999,N_12839,N_12804);
nor U13000 (N_13000,N_12950,N_12887);
or U13001 (N_13001,N_12962,N_12933);
or U13002 (N_13002,N_12941,N_12969);
or U13003 (N_13003,N_12964,N_12900);
xor U13004 (N_13004,N_12926,N_12890);
nor U13005 (N_13005,N_12908,N_12907);
nor U13006 (N_13006,N_12963,N_12966);
xor U13007 (N_13007,N_12883,N_12975);
nand U13008 (N_13008,N_12879,N_12994);
xnor U13009 (N_13009,N_12917,N_12939);
nand U13010 (N_13010,N_12953,N_12955);
xnor U13011 (N_13011,N_12995,N_12997);
nand U13012 (N_13012,N_12911,N_12896);
nor U13013 (N_13013,N_12988,N_12936);
and U13014 (N_13014,N_12987,N_12924);
nor U13015 (N_13015,N_12948,N_12930);
or U13016 (N_13016,N_12932,N_12970);
xnor U13017 (N_13017,N_12905,N_12897);
nand U13018 (N_13018,N_12946,N_12980);
xor U13019 (N_13019,N_12959,N_12923);
nand U13020 (N_13020,N_12938,N_12876);
nor U13021 (N_13021,N_12903,N_12881);
nand U13022 (N_13022,N_12989,N_12934);
xor U13023 (N_13023,N_12940,N_12882);
and U13024 (N_13024,N_12958,N_12921);
xor U13025 (N_13025,N_12954,N_12929);
or U13026 (N_13026,N_12947,N_12945);
nand U13027 (N_13027,N_12993,N_12880);
nand U13028 (N_13028,N_12922,N_12898);
nand U13029 (N_13029,N_12951,N_12979);
and U13030 (N_13030,N_12944,N_12877);
xor U13031 (N_13031,N_12996,N_12893);
nor U13032 (N_13032,N_12937,N_12992);
nor U13033 (N_13033,N_12985,N_12971);
xnor U13034 (N_13034,N_12931,N_12986);
or U13035 (N_13035,N_12957,N_12998);
xnor U13036 (N_13036,N_12984,N_12981);
or U13037 (N_13037,N_12888,N_12973);
nor U13038 (N_13038,N_12915,N_12904);
nor U13039 (N_13039,N_12967,N_12978);
and U13040 (N_13040,N_12906,N_12999);
xnor U13041 (N_13041,N_12909,N_12914);
xnor U13042 (N_13042,N_12935,N_12878);
xnor U13043 (N_13043,N_12885,N_12956);
or U13044 (N_13044,N_12974,N_12972);
xor U13045 (N_13045,N_12990,N_12961);
nand U13046 (N_13046,N_12919,N_12912);
nor U13047 (N_13047,N_12920,N_12892);
xor U13048 (N_13048,N_12983,N_12925);
nor U13049 (N_13049,N_12928,N_12918);
and U13050 (N_13050,N_12884,N_12889);
nand U13051 (N_13051,N_12977,N_12991);
nor U13052 (N_13052,N_12902,N_12894);
or U13053 (N_13053,N_12960,N_12976);
nand U13054 (N_13054,N_12942,N_12927);
or U13055 (N_13055,N_12910,N_12875);
xor U13056 (N_13056,N_12901,N_12886);
xnor U13057 (N_13057,N_12913,N_12982);
nand U13058 (N_13058,N_12891,N_12968);
or U13059 (N_13059,N_12949,N_12952);
and U13060 (N_13060,N_12943,N_12916);
xor U13061 (N_13061,N_12895,N_12899);
and U13062 (N_13062,N_12965,N_12943);
or U13063 (N_13063,N_12965,N_12986);
or U13064 (N_13064,N_12992,N_12959);
xor U13065 (N_13065,N_12947,N_12885);
or U13066 (N_13066,N_12930,N_12919);
and U13067 (N_13067,N_12960,N_12924);
and U13068 (N_13068,N_12935,N_12916);
nor U13069 (N_13069,N_12940,N_12996);
nand U13070 (N_13070,N_12904,N_12884);
and U13071 (N_13071,N_12934,N_12959);
or U13072 (N_13072,N_12979,N_12989);
and U13073 (N_13073,N_12918,N_12917);
xnor U13074 (N_13074,N_12917,N_12904);
nand U13075 (N_13075,N_12926,N_12956);
xnor U13076 (N_13076,N_12912,N_12977);
or U13077 (N_13077,N_12949,N_12907);
and U13078 (N_13078,N_12877,N_12936);
xnor U13079 (N_13079,N_12948,N_12908);
and U13080 (N_13080,N_12950,N_12930);
nand U13081 (N_13081,N_12973,N_12962);
and U13082 (N_13082,N_12917,N_12911);
nand U13083 (N_13083,N_12890,N_12880);
nand U13084 (N_13084,N_12937,N_12902);
nor U13085 (N_13085,N_12966,N_12918);
nand U13086 (N_13086,N_12943,N_12878);
xor U13087 (N_13087,N_12905,N_12986);
nor U13088 (N_13088,N_12974,N_12992);
and U13089 (N_13089,N_12964,N_12999);
xor U13090 (N_13090,N_12879,N_12890);
xnor U13091 (N_13091,N_12983,N_12912);
and U13092 (N_13092,N_12983,N_12990);
nand U13093 (N_13093,N_12900,N_12911);
nor U13094 (N_13094,N_12942,N_12911);
xnor U13095 (N_13095,N_12920,N_12960);
xor U13096 (N_13096,N_12946,N_12973);
nand U13097 (N_13097,N_12919,N_12924);
or U13098 (N_13098,N_12934,N_12914);
xor U13099 (N_13099,N_12936,N_12957);
or U13100 (N_13100,N_12989,N_12997);
xor U13101 (N_13101,N_12917,N_12875);
or U13102 (N_13102,N_12887,N_12888);
and U13103 (N_13103,N_12876,N_12890);
nor U13104 (N_13104,N_12892,N_12905);
xnor U13105 (N_13105,N_12908,N_12936);
and U13106 (N_13106,N_12896,N_12955);
nand U13107 (N_13107,N_12911,N_12949);
nand U13108 (N_13108,N_12912,N_12910);
nand U13109 (N_13109,N_12904,N_12886);
and U13110 (N_13110,N_12875,N_12898);
xnor U13111 (N_13111,N_12891,N_12989);
nand U13112 (N_13112,N_12989,N_12971);
or U13113 (N_13113,N_12912,N_12992);
or U13114 (N_13114,N_12880,N_12911);
nand U13115 (N_13115,N_12905,N_12943);
xor U13116 (N_13116,N_12899,N_12932);
or U13117 (N_13117,N_12953,N_12979);
or U13118 (N_13118,N_12924,N_12888);
nand U13119 (N_13119,N_12995,N_12974);
xnor U13120 (N_13120,N_12910,N_12887);
nand U13121 (N_13121,N_12945,N_12896);
and U13122 (N_13122,N_12892,N_12917);
nor U13123 (N_13123,N_12879,N_12998);
or U13124 (N_13124,N_12891,N_12897);
nor U13125 (N_13125,N_13077,N_13119);
and U13126 (N_13126,N_13010,N_13023);
and U13127 (N_13127,N_13056,N_13004);
and U13128 (N_13128,N_13079,N_13039);
nand U13129 (N_13129,N_13046,N_13052);
xor U13130 (N_13130,N_13008,N_13053);
xor U13131 (N_13131,N_13091,N_13019);
xnor U13132 (N_13132,N_13067,N_13120);
or U13133 (N_13133,N_13109,N_13071);
and U13134 (N_13134,N_13058,N_13003);
nor U13135 (N_13135,N_13098,N_13107);
xor U13136 (N_13136,N_13082,N_13122);
or U13137 (N_13137,N_13049,N_13088);
xnor U13138 (N_13138,N_13114,N_13016);
xnor U13139 (N_13139,N_13047,N_13095);
or U13140 (N_13140,N_13017,N_13036);
xnor U13141 (N_13141,N_13033,N_13031);
xor U13142 (N_13142,N_13045,N_13061);
xor U13143 (N_13143,N_13013,N_13044);
and U13144 (N_13144,N_13117,N_13086);
and U13145 (N_13145,N_13078,N_13057);
nand U13146 (N_13146,N_13099,N_13068);
xor U13147 (N_13147,N_13034,N_13014);
nand U13148 (N_13148,N_13076,N_13073);
or U13149 (N_13149,N_13038,N_13000);
or U13150 (N_13150,N_13085,N_13035);
xor U13151 (N_13151,N_13075,N_13104);
or U13152 (N_13152,N_13106,N_13024);
and U13153 (N_13153,N_13103,N_13066);
and U13154 (N_13154,N_13025,N_13060);
nor U13155 (N_13155,N_13027,N_13041);
nor U13156 (N_13156,N_13054,N_13090);
or U13157 (N_13157,N_13018,N_13009);
nor U13158 (N_13158,N_13080,N_13084);
nand U13159 (N_13159,N_13020,N_13118);
nand U13160 (N_13160,N_13102,N_13113);
or U13161 (N_13161,N_13065,N_13002);
nand U13162 (N_13162,N_13040,N_13121);
nor U13163 (N_13163,N_13097,N_13062);
nor U13164 (N_13164,N_13042,N_13123);
xnor U13165 (N_13165,N_13096,N_13081);
nand U13166 (N_13166,N_13105,N_13072);
and U13167 (N_13167,N_13116,N_13007);
xnor U13168 (N_13168,N_13055,N_13059);
nand U13169 (N_13169,N_13087,N_13030);
nand U13170 (N_13170,N_13011,N_13037);
and U13171 (N_13171,N_13022,N_13012);
nor U13172 (N_13172,N_13032,N_13110);
and U13173 (N_13173,N_13026,N_13100);
nand U13174 (N_13174,N_13089,N_13092);
and U13175 (N_13175,N_13115,N_13005);
or U13176 (N_13176,N_13051,N_13070);
and U13177 (N_13177,N_13050,N_13093);
and U13178 (N_13178,N_13043,N_13112);
nor U13179 (N_13179,N_13111,N_13064);
nand U13180 (N_13180,N_13006,N_13094);
or U13181 (N_13181,N_13048,N_13074);
nand U13182 (N_13182,N_13015,N_13069);
and U13183 (N_13183,N_13063,N_13108);
xor U13184 (N_13184,N_13083,N_13101);
or U13185 (N_13185,N_13028,N_13001);
xor U13186 (N_13186,N_13029,N_13124);
or U13187 (N_13187,N_13021,N_13042);
nor U13188 (N_13188,N_13050,N_13085);
nand U13189 (N_13189,N_13007,N_13080);
nand U13190 (N_13190,N_13046,N_13028);
nand U13191 (N_13191,N_13039,N_13056);
nand U13192 (N_13192,N_13059,N_13113);
nand U13193 (N_13193,N_13043,N_13070);
nand U13194 (N_13194,N_13034,N_13035);
and U13195 (N_13195,N_13103,N_13030);
and U13196 (N_13196,N_13124,N_13010);
xnor U13197 (N_13197,N_13058,N_13078);
nand U13198 (N_13198,N_13005,N_13045);
or U13199 (N_13199,N_13064,N_13077);
xnor U13200 (N_13200,N_13022,N_13088);
and U13201 (N_13201,N_13033,N_13025);
or U13202 (N_13202,N_13066,N_13111);
xor U13203 (N_13203,N_13068,N_13103);
or U13204 (N_13204,N_13053,N_13077);
xor U13205 (N_13205,N_13103,N_13005);
or U13206 (N_13206,N_13013,N_13085);
nand U13207 (N_13207,N_13025,N_13110);
and U13208 (N_13208,N_13048,N_13065);
nand U13209 (N_13209,N_13004,N_13001);
nor U13210 (N_13210,N_13065,N_13121);
nor U13211 (N_13211,N_13093,N_13063);
or U13212 (N_13212,N_13050,N_13072);
or U13213 (N_13213,N_13075,N_13106);
or U13214 (N_13214,N_13056,N_13110);
xor U13215 (N_13215,N_13034,N_13056);
and U13216 (N_13216,N_13095,N_13080);
nor U13217 (N_13217,N_13044,N_13045);
nor U13218 (N_13218,N_13069,N_13030);
xnor U13219 (N_13219,N_13030,N_13014);
and U13220 (N_13220,N_13069,N_13054);
nor U13221 (N_13221,N_13070,N_13100);
xnor U13222 (N_13222,N_13104,N_13033);
nand U13223 (N_13223,N_13044,N_13025);
nand U13224 (N_13224,N_13119,N_13121);
or U13225 (N_13225,N_13081,N_13030);
or U13226 (N_13226,N_13048,N_13050);
or U13227 (N_13227,N_13042,N_13101);
or U13228 (N_13228,N_13095,N_13058);
or U13229 (N_13229,N_13095,N_13092);
and U13230 (N_13230,N_13077,N_13005);
and U13231 (N_13231,N_13036,N_13101);
and U13232 (N_13232,N_13021,N_13076);
and U13233 (N_13233,N_13015,N_13025);
and U13234 (N_13234,N_13112,N_13103);
xnor U13235 (N_13235,N_13093,N_13095);
and U13236 (N_13236,N_13009,N_13041);
nand U13237 (N_13237,N_13057,N_13107);
nand U13238 (N_13238,N_13051,N_13000);
and U13239 (N_13239,N_13002,N_13110);
xor U13240 (N_13240,N_13098,N_13005);
xor U13241 (N_13241,N_13057,N_13023);
or U13242 (N_13242,N_13082,N_13065);
and U13243 (N_13243,N_13119,N_13034);
or U13244 (N_13244,N_13032,N_13114);
and U13245 (N_13245,N_13076,N_13063);
or U13246 (N_13246,N_13078,N_13021);
or U13247 (N_13247,N_13049,N_13083);
xor U13248 (N_13248,N_13047,N_13036);
xor U13249 (N_13249,N_13049,N_13042);
xnor U13250 (N_13250,N_13127,N_13202);
and U13251 (N_13251,N_13219,N_13147);
and U13252 (N_13252,N_13198,N_13224);
or U13253 (N_13253,N_13248,N_13146);
or U13254 (N_13254,N_13243,N_13209);
nor U13255 (N_13255,N_13132,N_13196);
xor U13256 (N_13256,N_13215,N_13189);
and U13257 (N_13257,N_13130,N_13195);
or U13258 (N_13258,N_13235,N_13186);
xnor U13259 (N_13259,N_13182,N_13199);
or U13260 (N_13260,N_13156,N_13126);
and U13261 (N_13261,N_13154,N_13184);
or U13262 (N_13262,N_13159,N_13249);
xnor U13263 (N_13263,N_13133,N_13246);
nor U13264 (N_13264,N_13229,N_13232);
nor U13265 (N_13265,N_13225,N_13178);
nand U13266 (N_13266,N_13173,N_13171);
xnor U13267 (N_13267,N_13192,N_13221);
or U13268 (N_13268,N_13181,N_13172);
nor U13269 (N_13269,N_13213,N_13241);
nor U13270 (N_13270,N_13148,N_13128);
xor U13271 (N_13271,N_13206,N_13138);
and U13272 (N_13272,N_13245,N_13185);
xnor U13273 (N_13273,N_13234,N_13169);
or U13274 (N_13274,N_13160,N_13145);
nor U13275 (N_13275,N_13239,N_13180);
nor U13276 (N_13276,N_13141,N_13136);
and U13277 (N_13277,N_13157,N_13142);
xnor U13278 (N_13278,N_13131,N_13150);
xnor U13279 (N_13279,N_13220,N_13161);
nor U13280 (N_13280,N_13176,N_13167);
nor U13281 (N_13281,N_13238,N_13194);
xor U13282 (N_13282,N_13214,N_13125);
or U13283 (N_13283,N_13140,N_13197);
nand U13284 (N_13284,N_13151,N_13193);
and U13285 (N_13285,N_13208,N_13152);
xnor U13286 (N_13286,N_13166,N_13240);
or U13287 (N_13287,N_13179,N_13230);
and U13288 (N_13288,N_13139,N_13218);
or U13289 (N_13289,N_13174,N_13217);
nor U13290 (N_13290,N_13134,N_13203);
or U13291 (N_13291,N_13143,N_13222);
xor U13292 (N_13292,N_13135,N_13223);
nand U13293 (N_13293,N_13153,N_13226);
and U13294 (N_13294,N_13175,N_13210);
xor U13295 (N_13295,N_13236,N_13168);
nand U13296 (N_13296,N_13216,N_13155);
or U13297 (N_13297,N_13231,N_13163);
or U13298 (N_13298,N_13227,N_13137);
and U13299 (N_13299,N_13212,N_13233);
or U13300 (N_13300,N_13200,N_13188);
xnor U13301 (N_13301,N_13187,N_13237);
or U13302 (N_13302,N_13190,N_13228);
and U13303 (N_13303,N_13211,N_13164);
and U13304 (N_13304,N_13170,N_13191);
nand U13305 (N_13305,N_13242,N_13204);
nor U13306 (N_13306,N_13158,N_13244);
nand U13307 (N_13307,N_13205,N_13177);
xor U13308 (N_13308,N_13162,N_13129);
or U13309 (N_13309,N_13144,N_13149);
xor U13310 (N_13310,N_13207,N_13201);
or U13311 (N_13311,N_13247,N_13183);
nor U13312 (N_13312,N_13165,N_13176);
nand U13313 (N_13313,N_13130,N_13216);
xnor U13314 (N_13314,N_13195,N_13249);
xor U13315 (N_13315,N_13130,N_13219);
nor U13316 (N_13316,N_13145,N_13228);
or U13317 (N_13317,N_13219,N_13243);
nor U13318 (N_13318,N_13136,N_13178);
nor U13319 (N_13319,N_13235,N_13233);
or U13320 (N_13320,N_13228,N_13194);
nor U13321 (N_13321,N_13209,N_13165);
and U13322 (N_13322,N_13198,N_13143);
or U13323 (N_13323,N_13186,N_13195);
nor U13324 (N_13324,N_13148,N_13147);
and U13325 (N_13325,N_13169,N_13244);
or U13326 (N_13326,N_13204,N_13224);
nand U13327 (N_13327,N_13226,N_13216);
or U13328 (N_13328,N_13238,N_13170);
and U13329 (N_13329,N_13150,N_13175);
and U13330 (N_13330,N_13215,N_13246);
nand U13331 (N_13331,N_13180,N_13188);
xnor U13332 (N_13332,N_13183,N_13180);
or U13333 (N_13333,N_13218,N_13131);
and U13334 (N_13334,N_13149,N_13172);
nor U13335 (N_13335,N_13171,N_13164);
or U13336 (N_13336,N_13161,N_13242);
nor U13337 (N_13337,N_13225,N_13180);
xnor U13338 (N_13338,N_13183,N_13178);
or U13339 (N_13339,N_13147,N_13236);
and U13340 (N_13340,N_13203,N_13247);
or U13341 (N_13341,N_13130,N_13210);
nand U13342 (N_13342,N_13197,N_13190);
nand U13343 (N_13343,N_13168,N_13187);
nand U13344 (N_13344,N_13154,N_13231);
nand U13345 (N_13345,N_13151,N_13169);
or U13346 (N_13346,N_13219,N_13171);
or U13347 (N_13347,N_13133,N_13165);
nor U13348 (N_13348,N_13147,N_13132);
or U13349 (N_13349,N_13193,N_13128);
nor U13350 (N_13350,N_13145,N_13171);
nand U13351 (N_13351,N_13209,N_13239);
and U13352 (N_13352,N_13198,N_13196);
or U13353 (N_13353,N_13241,N_13235);
and U13354 (N_13354,N_13192,N_13190);
and U13355 (N_13355,N_13139,N_13222);
or U13356 (N_13356,N_13221,N_13243);
nor U13357 (N_13357,N_13211,N_13174);
nand U13358 (N_13358,N_13126,N_13148);
and U13359 (N_13359,N_13212,N_13230);
nand U13360 (N_13360,N_13130,N_13161);
nand U13361 (N_13361,N_13218,N_13162);
or U13362 (N_13362,N_13138,N_13133);
or U13363 (N_13363,N_13208,N_13225);
or U13364 (N_13364,N_13156,N_13207);
xor U13365 (N_13365,N_13177,N_13170);
nor U13366 (N_13366,N_13127,N_13221);
or U13367 (N_13367,N_13200,N_13177);
or U13368 (N_13368,N_13237,N_13222);
nor U13369 (N_13369,N_13238,N_13173);
xnor U13370 (N_13370,N_13242,N_13159);
nor U13371 (N_13371,N_13184,N_13131);
and U13372 (N_13372,N_13136,N_13227);
nand U13373 (N_13373,N_13158,N_13140);
xor U13374 (N_13374,N_13151,N_13186);
or U13375 (N_13375,N_13287,N_13262);
nor U13376 (N_13376,N_13363,N_13372);
or U13377 (N_13377,N_13252,N_13281);
or U13378 (N_13378,N_13373,N_13294);
nand U13379 (N_13379,N_13368,N_13370);
nand U13380 (N_13380,N_13296,N_13317);
nor U13381 (N_13381,N_13335,N_13282);
nand U13382 (N_13382,N_13293,N_13319);
xnor U13383 (N_13383,N_13374,N_13286);
xor U13384 (N_13384,N_13332,N_13269);
xnor U13385 (N_13385,N_13289,N_13348);
nor U13386 (N_13386,N_13360,N_13353);
and U13387 (N_13387,N_13284,N_13329);
nor U13388 (N_13388,N_13295,N_13250);
nand U13389 (N_13389,N_13251,N_13318);
nand U13390 (N_13390,N_13265,N_13283);
and U13391 (N_13391,N_13371,N_13345);
nor U13392 (N_13392,N_13280,N_13343);
and U13393 (N_13393,N_13341,N_13357);
or U13394 (N_13394,N_13321,N_13333);
or U13395 (N_13395,N_13346,N_13266);
nand U13396 (N_13396,N_13256,N_13362);
or U13397 (N_13397,N_13304,N_13347);
or U13398 (N_13398,N_13331,N_13285);
or U13399 (N_13399,N_13261,N_13358);
or U13400 (N_13400,N_13338,N_13271);
xnor U13401 (N_13401,N_13327,N_13350);
or U13402 (N_13402,N_13355,N_13258);
nor U13403 (N_13403,N_13308,N_13259);
or U13404 (N_13404,N_13326,N_13255);
or U13405 (N_13405,N_13276,N_13320);
nand U13406 (N_13406,N_13334,N_13356);
or U13407 (N_13407,N_13300,N_13328);
or U13408 (N_13408,N_13344,N_13324);
nand U13409 (N_13409,N_13288,N_13322);
and U13410 (N_13410,N_13325,N_13301);
xnor U13411 (N_13411,N_13254,N_13279);
nand U13412 (N_13412,N_13369,N_13342);
and U13413 (N_13413,N_13291,N_13268);
nand U13414 (N_13414,N_13310,N_13270);
nand U13415 (N_13415,N_13303,N_13354);
nand U13416 (N_13416,N_13306,N_13315);
nor U13417 (N_13417,N_13330,N_13264);
nand U13418 (N_13418,N_13352,N_13292);
or U13419 (N_13419,N_13302,N_13311);
xnor U13420 (N_13420,N_13349,N_13313);
xnor U13421 (N_13421,N_13307,N_13367);
nor U13422 (N_13422,N_13260,N_13253);
nor U13423 (N_13423,N_13365,N_13359);
nor U13424 (N_13424,N_13263,N_13277);
xnor U13425 (N_13425,N_13298,N_13361);
nand U13426 (N_13426,N_13273,N_13267);
nor U13427 (N_13427,N_13309,N_13305);
xnor U13428 (N_13428,N_13274,N_13299);
nand U13429 (N_13429,N_13366,N_13337);
nor U13430 (N_13430,N_13272,N_13278);
nor U13431 (N_13431,N_13340,N_13275);
or U13432 (N_13432,N_13323,N_13351);
or U13433 (N_13433,N_13257,N_13339);
nor U13434 (N_13434,N_13336,N_13316);
and U13435 (N_13435,N_13312,N_13314);
and U13436 (N_13436,N_13290,N_13364);
nand U13437 (N_13437,N_13297,N_13313);
or U13438 (N_13438,N_13309,N_13289);
xor U13439 (N_13439,N_13296,N_13274);
or U13440 (N_13440,N_13332,N_13311);
nand U13441 (N_13441,N_13311,N_13327);
nand U13442 (N_13442,N_13345,N_13360);
xnor U13443 (N_13443,N_13302,N_13256);
nor U13444 (N_13444,N_13253,N_13316);
nor U13445 (N_13445,N_13262,N_13354);
or U13446 (N_13446,N_13251,N_13337);
and U13447 (N_13447,N_13254,N_13358);
and U13448 (N_13448,N_13291,N_13332);
nor U13449 (N_13449,N_13364,N_13269);
nand U13450 (N_13450,N_13374,N_13250);
nand U13451 (N_13451,N_13297,N_13341);
nand U13452 (N_13452,N_13319,N_13281);
xor U13453 (N_13453,N_13334,N_13351);
nand U13454 (N_13454,N_13343,N_13313);
or U13455 (N_13455,N_13287,N_13301);
nor U13456 (N_13456,N_13257,N_13357);
and U13457 (N_13457,N_13345,N_13254);
nand U13458 (N_13458,N_13311,N_13283);
nand U13459 (N_13459,N_13339,N_13310);
and U13460 (N_13460,N_13274,N_13345);
nor U13461 (N_13461,N_13304,N_13322);
nand U13462 (N_13462,N_13266,N_13322);
nor U13463 (N_13463,N_13357,N_13270);
nand U13464 (N_13464,N_13337,N_13257);
nor U13465 (N_13465,N_13306,N_13257);
nor U13466 (N_13466,N_13315,N_13361);
nor U13467 (N_13467,N_13302,N_13361);
xnor U13468 (N_13468,N_13266,N_13269);
xnor U13469 (N_13469,N_13316,N_13346);
and U13470 (N_13470,N_13357,N_13280);
nand U13471 (N_13471,N_13264,N_13368);
nor U13472 (N_13472,N_13291,N_13371);
nor U13473 (N_13473,N_13265,N_13281);
nor U13474 (N_13474,N_13356,N_13260);
nand U13475 (N_13475,N_13349,N_13282);
xor U13476 (N_13476,N_13259,N_13349);
nor U13477 (N_13477,N_13357,N_13330);
nand U13478 (N_13478,N_13347,N_13251);
nand U13479 (N_13479,N_13296,N_13307);
xor U13480 (N_13480,N_13266,N_13313);
xor U13481 (N_13481,N_13370,N_13365);
or U13482 (N_13482,N_13365,N_13345);
nor U13483 (N_13483,N_13261,N_13304);
or U13484 (N_13484,N_13270,N_13359);
nand U13485 (N_13485,N_13370,N_13330);
nand U13486 (N_13486,N_13269,N_13290);
nand U13487 (N_13487,N_13281,N_13328);
nor U13488 (N_13488,N_13363,N_13295);
nor U13489 (N_13489,N_13276,N_13257);
and U13490 (N_13490,N_13347,N_13267);
nor U13491 (N_13491,N_13348,N_13320);
and U13492 (N_13492,N_13318,N_13333);
nor U13493 (N_13493,N_13322,N_13373);
or U13494 (N_13494,N_13335,N_13308);
nand U13495 (N_13495,N_13366,N_13325);
nor U13496 (N_13496,N_13350,N_13368);
nor U13497 (N_13497,N_13286,N_13264);
or U13498 (N_13498,N_13346,N_13329);
and U13499 (N_13499,N_13294,N_13305);
xnor U13500 (N_13500,N_13490,N_13475);
xnor U13501 (N_13501,N_13417,N_13424);
nor U13502 (N_13502,N_13408,N_13375);
nor U13503 (N_13503,N_13430,N_13399);
or U13504 (N_13504,N_13426,N_13387);
or U13505 (N_13505,N_13459,N_13420);
nand U13506 (N_13506,N_13394,N_13380);
nand U13507 (N_13507,N_13434,N_13383);
and U13508 (N_13508,N_13427,N_13378);
xor U13509 (N_13509,N_13382,N_13429);
or U13510 (N_13510,N_13440,N_13488);
nor U13511 (N_13511,N_13403,N_13481);
nand U13512 (N_13512,N_13428,N_13467);
and U13513 (N_13513,N_13453,N_13478);
nand U13514 (N_13514,N_13423,N_13419);
xnor U13515 (N_13515,N_13442,N_13445);
and U13516 (N_13516,N_13471,N_13395);
and U13517 (N_13517,N_13496,N_13379);
and U13518 (N_13518,N_13413,N_13452);
nand U13519 (N_13519,N_13454,N_13415);
nand U13520 (N_13520,N_13389,N_13492);
and U13521 (N_13521,N_13414,N_13497);
nor U13522 (N_13522,N_13499,N_13435);
xor U13523 (N_13523,N_13450,N_13432);
nand U13524 (N_13524,N_13460,N_13495);
nor U13525 (N_13525,N_13451,N_13464);
nand U13526 (N_13526,N_13480,N_13470);
nor U13527 (N_13527,N_13412,N_13418);
xor U13528 (N_13528,N_13461,N_13487);
or U13529 (N_13529,N_13409,N_13463);
nor U13530 (N_13530,N_13407,N_13391);
xnor U13531 (N_13531,N_13491,N_13458);
xnor U13532 (N_13532,N_13479,N_13474);
xnor U13533 (N_13533,N_13468,N_13441);
or U13534 (N_13534,N_13436,N_13411);
or U13535 (N_13535,N_13425,N_13438);
nand U13536 (N_13536,N_13498,N_13483);
nor U13537 (N_13537,N_13485,N_13386);
nor U13538 (N_13538,N_13473,N_13455);
and U13539 (N_13539,N_13489,N_13465);
and U13540 (N_13540,N_13437,N_13393);
xor U13541 (N_13541,N_13482,N_13444);
and U13542 (N_13542,N_13416,N_13446);
or U13543 (N_13543,N_13439,N_13397);
or U13544 (N_13544,N_13381,N_13404);
xnor U13545 (N_13545,N_13422,N_13447);
or U13546 (N_13546,N_13472,N_13398);
nand U13547 (N_13547,N_13384,N_13456);
xnor U13548 (N_13548,N_13466,N_13477);
xnor U13549 (N_13549,N_13388,N_13443);
nor U13550 (N_13550,N_13396,N_13449);
or U13551 (N_13551,N_13401,N_13457);
nor U13552 (N_13552,N_13376,N_13433);
nand U13553 (N_13553,N_13392,N_13469);
nand U13554 (N_13554,N_13410,N_13400);
nor U13555 (N_13555,N_13448,N_13390);
xnor U13556 (N_13556,N_13476,N_13484);
or U13557 (N_13557,N_13402,N_13377);
nor U13558 (N_13558,N_13493,N_13421);
xor U13559 (N_13559,N_13405,N_13486);
nand U13560 (N_13560,N_13494,N_13385);
xor U13561 (N_13561,N_13406,N_13431);
or U13562 (N_13562,N_13462,N_13406);
nor U13563 (N_13563,N_13462,N_13436);
xnor U13564 (N_13564,N_13417,N_13490);
nand U13565 (N_13565,N_13477,N_13423);
nor U13566 (N_13566,N_13437,N_13381);
nor U13567 (N_13567,N_13413,N_13400);
nand U13568 (N_13568,N_13398,N_13473);
or U13569 (N_13569,N_13403,N_13475);
or U13570 (N_13570,N_13460,N_13488);
and U13571 (N_13571,N_13439,N_13463);
nand U13572 (N_13572,N_13380,N_13414);
and U13573 (N_13573,N_13382,N_13477);
or U13574 (N_13574,N_13433,N_13405);
xnor U13575 (N_13575,N_13380,N_13388);
nor U13576 (N_13576,N_13440,N_13421);
nand U13577 (N_13577,N_13497,N_13471);
xor U13578 (N_13578,N_13461,N_13492);
and U13579 (N_13579,N_13422,N_13464);
nor U13580 (N_13580,N_13395,N_13496);
and U13581 (N_13581,N_13468,N_13482);
and U13582 (N_13582,N_13407,N_13451);
or U13583 (N_13583,N_13451,N_13490);
and U13584 (N_13584,N_13421,N_13494);
and U13585 (N_13585,N_13458,N_13381);
nand U13586 (N_13586,N_13493,N_13397);
nor U13587 (N_13587,N_13477,N_13496);
nand U13588 (N_13588,N_13408,N_13442);
xnor U13589 (N_13589,N_13492,N_13469);
xor U13590 (N_13590,N_13401,N_13431);
xnor U13591 (N_13591,N_13413,N_13481);
nor U13592 (N_13592,N_13480,N_13490);
xor U13593 (N_13593,N_13402,N_13470);
and U13594 (N_13594,N_13437,N_13471);
or U13595 (N_13595,N_13375,N_13457);
nor U13596 (N_13596,N_13451,N_13377);
xor U13597 (N_13597,N_13396,N_13400);
and U13598 (N_13598,N_13472,N_13495);
and U13599 (N_13599,N_13389,N_13426);
nor U13600 (N_13600,N_13426,N_13481);
nor U13601 (N_13601,N_13438,N_13406);
xor U13602 (N_13602,N_13378,N_13420);
nor U13603 (N_13603,N_13378,N_13488);
xnor U13604 (N_13604,N_13440,N_13420);
and U13605 (N_13605,N_13401,N_13418);
or U13606 (N_13606,N_13486,N_13434);
nand U13607 (N_13607,N_13429,N_13477);
xnor U13608 (N_13608,N_13431,N_13437);
nor U13609 (N_13609,N_13471,N_13415);
nand U13610 (N_13610,N_13483,N_13428);
and U13611 (N_13611,N_13495,N_13386);
or U13612 (N_13612,N_13377,N_13468);
and U13613 (N_13613,N_13410,N_13412);
nor U13614 (N_13614,N_13409,N_13413);
and U13615 (N_13615,N_13431,N_13467);
and U13616 (N_13616,N_13392,N_13471);
and U13617 (N_13617,N_13433,N_13438);
and U13618 (N_13618,N_13409,N_13454);
nor U13619 (N_13619,N_13432,N_13407);
nor U13620 (N_13620,N_13379,N_13392);
or U13621 (N_13621,N_13466,N_13455);
and U13622 (N_13622,N_13438,N_13412);
nor U13623 (N_13623,N_13486,N_13487);
and U13624 (N_13624,N_13471,N_13377);
or U13625 (N_13625,N_13622,N_13585);
xnor U13626 (N_13626,N_13504,N_13533);
nand U13627 (N_13627,N_13577,N_13520);
nor U13628 (N_13628,N_13613,N_13525);
or U13629 (N_13629,N_13605,N_13584);
and U13630 (N_13630,N_13586,N_13553);
nor U13631 (N_13631,N_13593,N_13540);
nand U13632 (N_13632,N_13576,N_13524);
or U13633 (N_13633,N_13548,N_13606);
xnor U13634 (N_13634,N_13621,N_13550);
and U13635 (N_13635,N_13568,N_13541);
xnor U13636 (N_13636,N_13545,N_13614);
nor U13637 (N_13637,N_13523,N_13611);
xor U13638 (N_13638,N_13512,N_13594);
and U13639 (N_13639,N_13566,N_13589);
or U13640 (N_13640,N_13517,N_13515);
and U13641 (N_13641,N_13527,N_13560);
or U13642 (N_13642,N_13575,N_13501);
nand U13643 (N_13643,N_13569,N_13508);
xor U13644 (N_13644,N_13509,N_13506);
and U13645 (N_13645,N_13581,N_13574);
xnor U13646 (N_13646,N_13624,N_13552);
nand U13647 (N_13647,N_13591,N_13546);
and U13648 (N_13648,N_13538,N_13513);
and U13649 (N_13649,N_13556,N_13616);
nand U13650 (N_13650,N_13604,N_13602);
and U13651 (N_13651,N_13592,N_13519);
xnor U13652 (N_13652,N_13583,N_13514);
and U13653 (N_13653,N_13539,N_13572);
nor U13654 (N_13654,N_13564,N_13597);
nor U13655 (N_13655,N_13559,N_13543);
or U13656 (N_13656,N_13607,N_13547);
nor U13657 (N_13657,N_13578,N_13599);
nor U13658 (N_13658,N_13510,N_13557);
nand U13659 (N_13659,N_13535,N_13518);
nand U13660 (N_13660,N_13582,N_13600);
xnor U13661 (N_13661,N_13521,N_13596);
xor U13662 (N_13662,N_13571,N_13563);
nand U13663 (N_13663,N_13558,N_13526);
nor U13664 (N_13664,N_13598,N_13502);
and U13665 (N_13665,N_13610,N_13561);
nand U13666 (N_13666,N_13542,N_13507);
or U13667 (N_13667,N_13549,N_13528);
nand U13668 (N_13668,N_13565,N_13511);
and U13669 (N_13669,N_13617,N_13619);
or U13670 (N_13670,N_13573,N_13608);
xor U13671 (N_13671,N_13609,N_13536);
nand U13672 (N_13672,N_13532,N_13601);
or U13673 (N_13673,N_13522,N_13505);
or U13674 (N_13674,N_13554,N_13603);
or U13675 (N_13675,N_13537,N_13516);
and U13676 (N_13676,N_13615,N_13587);
xor U13677 (N_13677,N_13500,N_13530);
or U13678 (N_13678,N_13534,N_13623);
xnor U13679 (N_13679,N_13579,N_13567);
nor U13680 (N_13680,N_13580,N_13612);
and U13681 (N_13681,N_13544,N_13529);
and U13682 (N_13682,N_13503,N_13588);
nand U13683 (N_13683,N_13531,N_13570);
and U13684 (N_13684,N_13595,N_13555);
nand U13685 (N_13685,N_13618,N_13562);
nor U13686 (N_13686,N_13551,N_13590);
nand U13687 (N_13687,N_13620,N_13618);
or U13688 (N_13688,N_13588,N_13579);
nand U13689 (N_13689,N_13500,N_13619);
and U13690 (N_13690,N_13560,N_13618);
nand U13691 (N_13691,N_13501,N_13567);
xnor U13692 (N_13692,N_13559,N_13511);
nor U13693 (N_13693,N_13612,N_13524);
and U13694 (N_13694,N_13520,N_13564);
nor U13695 (N_13695,N_13619,N_13577);
nor U13696 (N_13696,N_13612,N_13562);
and U13697 (N_13697,N_13574,N_13542);
xor U13698 (N_13698,N_13536,N_13575);
and U13699 (N_13699,N_13622,N_13506);
xor U13700 (N_13700,N_13576,N_13510);
and U13701 (N_13701,N_13595,N_13618);
and U13702 (N_13702,N_13599,N_13507);
nor U13703 (N_13703,N_13623,N_13556);
or U13704 (N_13704,N_13504,N_13608);
and U13705 (N_13705,N_13552,N_13543);
nand U13706 (N_13706,N_13574,N_13532);
nor U13707 (N_13707,N_13587,N_13525);
or U13708 (N_13708,N_13588,N_13544);
or U13709 (N_13709,N_13560,N_13537);
nor U13710 (N_13710,N_13559,N_13539);
nor U13711 (N_13711,N_13622,N_13575);
nor U13712 (N_13712,N_13526,N_13582);
or U13713 (N_13713,N_13580,N_13557);
nand U13714 (N_13714,N_13529,N_13556);
xnor U13715 (N_13715,N_13601,N_13509);
nand U13716 (N_13716,N_13611,N_13573);
or U13717 (N_13717,N_13506,N_13545);
and U13718 (N_13718,N_13501,N_13516);
or U13719 (N_13719,N_13500,N_13575);
or U13720 (N_13720,N_13507,N_13526);
nor U13721 (N_13721,N_13540,N_13557);
and U13722 (N_13722,N_13500,N_13541);
nor U13723 (N_13723,N_13553,N_13593);
nand U13724 (N_13724,N_13501,N_13510);
and U13725 (N_13725,N_13558,N_13565);
or U13726 (N_13726,N_13532,N_13598);
nand U13727 (N_13727,N_13549,N_13550);
and U13728 (N_13728,N_13513,N_13501);
and U13729 (N_13729,N_13569,N_13612);
and U13730 (N_13730,N_13568,N_13587);
xnor U13731 (N_13731,N_13536,N_13503);
or U13732 (N_13732,N_13614,N_13548);
and U13733 (N_13733,N_13570,N_13555);
and U13734 (N_13734,N_13577,N_13601);
and U13735 (N_13735,N_13602,N_13573);
and U13736 (N_13736,N_13541,N_13537);
xnor U13737 (N_13737,N_13603,N_13522);
or U13738 (N_13738,N_13616,N_13579);
or U13739 (N_13739,N_13603,N_13568);
nand U13740 (N_13740,N_13575,N_13623);
and U13741 (N_13741,N_13585,N_13544);
nand U13742 (N_13742,N_13561,N_13504);
nor U13743 (N_13743,N_13617,N_13543);
and U13744 (N_13744,N_13604,N_13600);
nand U13745 (N_13745,N_13541,N_13607);
nor U13746 (N_13746,N_13615,N_13520);
nand U13747 (N_13747,N_13608,N_13617);
xnor U13748 (N_13748,N_13512,N_13600);
and U13749 (N_13749,N_13604,N_13549);
xor U13750 (N_13750,N_13742,N_13694);
xor U13751 (N_13751,N_13713,N_13741);
nor U13752 (N_13752,N_13682,N_13651);
and U13753 (N_13753,N_13730,N_13735);
nor U13754 (N_13754,N_13748,N_13710);
and U13755 (N_13755,N_13648,N_13629);
xor U13756 (N_13756,N_13683,N_13643);
nor U13757 (N_13757,N_13696,N_13702);
xnor U13758 (N_13758,N_13650,N_13640);
or U13759 (N_13759,N_13666,N_13734);
xor U13760 (N_13760,N_13711,N_13699);
nor U13761 (N_13761,N_13680,N_13658);
xnor U13762 (N_13762,N_13698,N_13642);
xor U13763 (N_13763,N_13728,N_13632);
nor U13764 (N_13764,N_13663,N_13655);
nor U13765 (N_13765,N_13636,N_13724);
or U13766 (N_13766,N_13675,N_13657);
and U13767 (N_13767,N_13739,N_13747);
and U13768 (N_13768,N_13644,N_13635);
nand U13769 (N_13769,N_13630,N_13708);
or U13770 (N_13770,N_13652,N_13720);
xor U13771 (N_13771,N_13678,N_13726);
nand U13772 (N_13772,N_13638,N_13725);
xor U13773 (N_13773,N_13661,N_13656);
nor U13774 (N_13774,N_13681,N_13674);
nor U13775 (N_13775,N_13628,N_13721);
xnor U13776 (N_13776,N_13715,N_13718);
and U13777 (N_13777,N_13740,N_13701);
nand U13778 (N_13778,N_13737,N_13660);
or U13779 (N_13779,N_13684,N_13695);
and U13780 (N_13780,N_13662,N_13687);
or U13781 (N_13781,N_13685,N_13727);
xnor U13782 (N_13782,N_13693,N_13679);
xor U13783 (N_13783,N_13639,N_13697);
nor U13784 (N_13784,N_13700,N_13631);
or U13785 (N_13785,N_13716,N_13634);
nor U13786 (N_13786,N_13641,N_13677);
nand U13787 (N_13787,N_13625,N_13729);
nand U13788 (N_13788,N_13744,N_13670);
nand U13789 (N_13789,N_13690,N_13627);
nor U13790 (N_13790,N_13707,N_13705);
and U13791 (N_13791,N_13659,N_13732);
xnor U13792 (N_13792,N_13709,N_13686);
nand U13793 (N_13793,N_13717,N_13647);
and U13794 (N_13794,N_13626,N_13749);
and U13795 (N_13795,N_13665,N_13714);
or U13796 (N_13796,N_13692,N_13671);
nand U13797 (N_13797,N_13645,N_13722);
and U13798 (N_13798,N_13746,N_13654);
xor U13799 (N_13799,N_13676,N_13731);
xnor U13800 (N_13800,N_13689,N_13637);
nand U13801 (N_13801,N_13673,N_13649);
or U13802 (N_13802,N_13691,N_13723);
and U13803 (N_13803,N_13633,N_13719);
nand U13804 (N_13804,N_13706,N_13646);
or U13805 (N_13805,N_13688,N_13736);
nor U13806 (N_13806,N_13738,N_13672);
nand U13807 (N_13807,N_13669,N_13667);
nor U13808 (N_13808,N_13733,N_13745);
or U13809 (N_13809,N_13653,N_13704);
nand U13810 (N_13810,N_13743,N_13703);
xor U13811 (N_13811,N_13664,N_13712);
or U13812 (N_13812,N_13668,N_13680);
nand U13813 (N_13813,N_13626,N_13719);
xor U13814 (N_13814,N_13684,N_13637);
and U13815 (N_13815,N_13693,N_13709);
nor U13816 (N_13816,N_13702,N_13724);
and U13817 (N_13817,N_13679,N_13688);
nand U13818 (N_13818,N_13657,N_13684);
xnor U13819 (N_13819,N_13723,N_13699);
xnor U13820 (N_13820,N_13683,N_13711);
xor U13821 (N_13821,N_13640,N_13710);
nor U13822 (N_13822,N_13724,N_13645);
and U13823 (N_13823,N_13644,N_13656);
and U13824 (N_13824,N_13651,N_13697);
or U13825 (N_13825,N_13631,N_13713);
and U13826 (N_13826,N_13635,N_13741);
or U13827 (N_13827,N_13688,N_13677);
nand U13828 (N_13828,N_13715,N_13741);
nor U13829 (N_13829,N_13738,N_13659);
nor U13830 (N_13830,N_13627,N_13719);
nor U13831 (N_13831,N_13649,N_13690);
nor U13832 (N_13832,N_13657,N_13710);
nand U13833 (N_13833,N_13654,N_13707);
nand U13834 (N_13834,N_13650,N_13676);
nand U13835 (N_13835,N_13707,N_13729);
nand U13836 (N_13836,N_13689,N_13725);
nand U13837 (N_13837,N_13739,N_13682);
nor U13838 (N_13838,N_13659,N_13700);
nor U13839 (N_13839,N_13646,N_13641);
and U13840 (N_13840,N_13639,N_13636);
and U13841 (N_13841,N_13625,N_13741);
nand U13842 (N_13842,N_13678,N_13693);
nand U13843 (N_13843,N_13661,N_13631);
nor U13844 (N_13844,N_13682,N_13629);
nor U13845 (N_13845,N_13658,N_13718);
or U13846 (N_13846,N_13705,N_13678);
nand U13847 (N_13847,N_13686,N_13742);
xnor U13848 (N_13848,N_13723,N_13634);
or U13849 (N_13849,N_13641,N_13721);
xnor U13850 (N_13850,N_13652,N_13717);
nor U13851 (N_13851,N_13630,N_13716);
and U13852 (N_13852,N_13676,N_13665);
or U13853 (N_13853,N_13682,N_13636);
or U13854 (N_13854,N_13739,N_13680);
nand U13855 (N_13855,N_13626,N_13656);
and U13856 (N_13856,N_13725,N_13680);
nand U13857 (N_13857,N_13674,N_13662);
nor U13858 (N_13858,N_13685,N_13651);
and U13859 (N_13859,N_13665,N_13718);
or U13860 (N_13860,N_13734,N_13654);
and U13861 (N_13861,N_13738,N_13683);
and U13862 (N_13862,N_13731,N_13744);
nand U13863 (N_13863,N_13672,N_13681);
nor U13864 (N_13864,N_13701,N_13660);
nand U13865 (N_13865,N_13673,N_13672);
nor U13866 (N_13866,N_13690,N_13670);
xnor U13867 (N_13867,N_13696,N_13719);
nand U13868 (N_13868,N_13657,N_13736);
xnor U13869 (N_13869,N_13647,N_13680);
nor U13870 (N_13870,N_13641,N_13672);
or U13871 (N_13871,N_13692,N_13673);
nand U13872 (N_13872,N_13663,N_13680);
or U13873 (N_13873,N_13723,N_13698);
nor U13874 (N_13874,N_13741,N_13673);
nor U13875 (N_13875,N_13818,N_13842);
xnor U13876 (N_13876,N_13817,N_13853);
or U13877 (N_13877,N_13750,N_13811);
and U13878 (N_13878,N_13819,N_13862);
nor U13879 (N_13879,N_13784,N_13755);
nand U13880 (N_13880,N_13833,N_13855);
nand U13881 (N_13881,N_13843,N_13756);
nand U13882 (N_13882,N_13788,N_13795);
nor U13883 (N_13883,N_13868,N_13780);
xnor U13884 (N_13884,N_13774,N_13797);
or U13885 (N_13885,N_13807,N_13849);
xor U13886 (N_13886,N_13814,N_13804);
nand U13887 (N_13887,N_13856,N_13844);
and U13888 (N_13888,N_13777,N_13823);
and U13889 (N_13889,N_13753,N_13866);
and U13890 (N_13890,N_13826,N_13752);
nand U13891 (N_13891,N_13813,N_13799);
or U13892 (N_13892,N_13761,N_13779);
xnor U13893 (N_13893,N_13794,N_13763);
nor U13894 (N_13894,N_13791,N_13835);
xor U13895 (N_13895,N_13839,N_13810);
nor U13896 (N_13896,N_13783,N_13751);
nor U13897 (N_13897,N_13836,N_13758);
and U13898 (N_13898,N_13834,N_13861);
and U13899 (N_13899,N_13765,N_13789);
xnor U13900 (N_13900,N_13785,N_13767);
and U13901 (N_13901,N_13820,N_13858);
nor U13902 (N_13902,N_13828,N_13792);
and U13903 (N_13903,N_13840,N_13852);
nor U13904 (N_13904,N_13821,N_13860);
xor U13905 (N_13905,N_13841,N_13865);
nand U13906 (N_13906,N_13806,N_13859);
and U13907 (N_13907,N_13854,N_13845);
nand U13908 (N_13908,N_13848,N_13822);
and U13909 (N_13909,N_13801,N_13798);
nand U13910 (N_13910,N_13796,N_13776);
xnor U13911 (N_13911,N_13769,N_13815);
xnor U13912 (N_13912,N_13764,N_13770);
xnor U13913 (N_13913,N_13782,N_13805);
nor U13914 (N_13914,N_13803,N_13873);
and U13915 (N_13915,N_13832,N_13831);
nor U13916 (N_13916,N_13864,N_13816);
xnor U13917 (N_13917,N_13771,N_13863);
xor U13918 (N_13918,N_13802,N_13870);
nand U13919 (N_13919,N_13790,N_13847);
or U13920 (N_13920,N_13872,N_13768);
nor U13921 (N_13921,N_13837,N_13827);
nand U13922 (N_13922,N_13809,N_13830);
nand U13923 (N_13923,N_13781,N_13760);
nand U13924 (N_13924,N_13869,N_13812);
nor U13925 (N_13925,N_13754,N_13867);
and U13926 (N_13926,N_13772,N_13778);
nor U13927 (N_13927,N_13775,N_13851);
nor U13928 (N_13928,N_13824,N_13846);
nand U13929 (N_13929,N_13829,N_13786);
nor U13930 (N_13930,N_13825,N_13874);
or U13931 (N_13931,N_13808,N_13766);
and U13932 (N_13932,N_13773,N_13850);
and U13933 (N_13933,N_13800,N_13857);
xor U13934 (N_13934,N_13787,N_13762);
xor U13935 (N_13935,N_13871,N_13793);
and U13936 (N_13936,N_13757,N_13759);
xor U13937 (N_13937,N_13838,N_13797);
or U13938 (N_13938,N_13799,N_13780);
or U13939 (N_13939,N_13800,N_13850);
and U13940 (N_13940,N_13759,N_13847);
or U13941 (N_13941,N_13847,N_13762);
and U13942 (N_13942,N_13759,N_13796);
or U13943 (N_13943,N_13828,N_13764);
and U13944 (N_13944,N_13813,N_13840);
xor U13945 (N_13945,N_13785,N_13848);
and U13946 (N_13946,N_13765,N_13759);
nand U13947 (N_13947,N_13811,N_13782);
and U13948 (N_13948,N_13853,N_13823);
and U13949 (N_13949,N_13856,N_13802);
xnor U13950 (N_13950,N_13770,N_13857);
nor U13951 (N_13951,N_13799,N_13859);
nand U13952 (N_13952,N_13754,N_13807);
and U13953 (N_13953,N_13773,N_13858);
or U13954 (N_13954,N_13786,N_13833);
nand U13955 (N_13955,N_13779,N_13764);
nand U13956 (N_13956,N_13853,N_13751);
nor U13957 (N_13957,N_13866,N_13847);
nor U13958 (N_13958,N_13820,N_13789);
nor U13959 (N_13959,N_13758,N_13815);
or U13960 (N_13960,N_13766,N_13859);
and U13961 (N_13961,N_13809,N_13818);
nand U13962 (N_13962,N_13865,N_13766);
and U13963 (N_13963,N_13802,N_13857);
nand U13964 (N_13964,N_13795,N_13832);
xnor U13965 (N_13965,N_13814,N_13794);
nor U13966 (N_13966,N_13858,N_13798);
xor U13967 (N_13967,N_13774,N_13789);
and U13968 (N_13968,N_13866,N_13873);
xnor U13969 (N_13969,N_13874,N_13777);
xnor U13970 (N_13970,N_13868,N_13763);
and U13971 (N_13971,N_13862,N_13799);
and U13972 (N_13972,N_13768,N_13769);
and U13973 (N_13973,N_13851,N_13861);
or U13974 (N_13974,N_13832,N_13750);
and U13975 (N_13975,N_13827,N_13835);
xor U13976 (N_13976,N_13831,N_13830);
or U13977 (N_13977,N_13799,N_13856);
nand U13978 (N_13978,N_13820,N_13782);
xor U13979 (N_13979,N_13824,N_13865);
and U13980 (N_13980,N_13768,N_13826);
nor U13981 (N_13981,N_13794,N_13784);
and U13982 (N_13982,N_13847,N_13776);
or U13983 (N_13983,N_13811,N_13772);
nor U13984 (N_13984,N_13872,N_13811);
xnor U13985 (N_13985,N_13823,N_13821);
nor U13986 (N_13986,N_13832,N_13784);
nand U13987 (N_13987,N_13760,N_13858);
or U13988 (N_13988,N_13813,N_13860);
nor U13989 (N_13989,N_13807,N_13818);
nand U13990 (N_13990,N_13778,N_13792);
nor U13991 (N_13991,N_13758,N_13753);
and U13992 (N_13992,N_13871,N_13825);
nor U13993 (N_13993,N_13781,N_13821);
or U13994 (N_13994,N_13803,N_13784);
nand U13995 (N_13995,N_13757,N_13798);
or U13996 (N_13996,N_13810,N_13751);
nand U13997 (N_13997,N_13759,N_13834);
xor U13998 (N_13998,N_13760,N_13792);
and U13999 (N_13999,N_13842,N_13756);
xor U14000 (N_14000,N_13956,N_13916);
and U14001 (N_14001,N_13888,N_13989);
and U14002 (N_14002,N_13886,N_13927);
nor U14003 (N_14003,N_13966,N_13995);
nor U14004 (N_14004,N_13951,N_13944);
nor U14005 (N_14005,N_13953,N_13997);
or U14006 (N_14006,N_13938,N_13941);
nand U14007 (N_14007,N_13923,N_13892);
nor U14008 (N_14008,N_13894,N_13972);
xnor U14009 (N_14009,N_13887,N_13949);
nand U14010 (N_14010,N_13942,N_13919);
and U14011 (N_14011,N_13975,N_13904);
xnor U14012 (N_14012,N_13906,N_13876);
xor U14013 (N_14013,N_13912,N_13915);
nor U14014 (N_14014,N_13910,N_13963);
and U14015 (N_14015,N_13982,N_13914);
xor U14016 (N_14016,N_13943,N_13969);
nand U14017 (N_14017,N_13946,N_13962);
nand U14018 (N_14018,N_13999,N_13958);
or U14019 (N_14019,N_13885,N_13952);
nor U14020 (N_14020,N_13984,N_13925);
nor U14021 (N_14021,N_13882,N_13889);
nor U14022 (N_14022,N_13974,N_13961);
nor U14023 (N_14023,N_13968,N_13891);
or U14024 (N_14024,N_13896,N_13909);
or U14025 (N_14025,N_13900,N_13911);
nand U14026 (N_14026,N_13990,N_13893);
nor U14027 (N_14027,N_13981,N_13898);
and U14028 (N_14028,N_13988,N_13932);
nand U14029 (N_14029,N_13971,N_13931);
nand U14030 (N_14030,N_13955,N_13905);
and U14031 (N_14031,N_13970,N_13985);
nand U14032 (N_14032,N_13879,N_13940);
xor U14033 (N_14033,N_13991,N_13908);
or U14034 (N_14034,N_13878,N_13895);
nor U14035 (N_14035,N_13987,N_13959);
xor U14036 (N_14036,N_13980,N_13921);
nor U14037 (N_14037,N_13992,N_13947);
xor U14038 (N_14038,N_13950,N_13986);
xnor U14039 (N_14039,N_13899,N_13933);
or U14040 (N_14040,N_13875,N_13937);
nor U14041 (N_14041,N_13945,N_13983);
nand U14042 (N_14042,N_13998,N_13973);
or U14043 (N_14043,N_13897,N_13924);
nor U14044 (N_14044,N_13996,N_13926);
xnor U14045 (N_14045,N_13993,N_13907);
xnor U14046 (N_14046,N_13979,N_13967);
nand U14047 (N_14047,N_13960,N_13901);
xnor U14048 (N_14048,N_13934,N_13976);
xnor U14049 (N_14049,N_13930,N_13994);
xnor U14050 (N_14050,N_13978,N_13913);
xor U14051 (N_14051,N_13936,N_13920);
and U14052 (N_14052,N_13935,N_13948);
xor U14053 (N_14053,N_13881,N_13918);
nand U14054 (N_14054,N_13954,N_13880);
or U14055 (N_14055,N_13890,N_13902);
and U14056 (N_14056,N_13957,N_13928);
xor U14057 (N_14057,N_13964,N_13965);
or U14058 (N_14058,N_13922,N_13883);
or U14059 (N_14059,N_13903,N_13877);
xor U14060 (N_14060,N_13917,N_13929);
or U14061 (N_14061,N_13939,N_13884);
nand U14062 (N_14062,N_13977,N_13909);
and U14063 (N_14063,N_13885,N_13932);
nor U14064 (N_14064,N_13901,N_13990);
or U14065 (N_14065,N_13970,N_13984);
and U14066 (N_14066,N_13932,N_13914);
nor U14067 (N_14067,N_13974,N_13895);
or U14068 (N_14068,N_13933,N_13954);
or U14069 (N_14069,N_13960,N_13976);
nor U14070 (N_14070,N_13964,N_13989);
nand U14071 (N_14071,N_13999,N_13895);
nand U14072 (N_14072,N_13886,N_13925);
nand U14073 (N_14073,N_13910,N_13885);
nand U14074 (N_14074,N_13954,N_13920);
nand U14075 (N_14075,N_13946,N_13969);
or U14076 (N_14076,N_13927,N_13963);
and U14077 (N_14077,N_13886,N_13940);
xnor U14078 (N_14078,N_13900,N_13952);
and U14079 (N_14079,N_13941,N_13883);
nand U14080 (N_14080,N_13995,N_13959);
or U14081 (N_14081,N_13970,N_13968);
nand U14082 (N_14082,N_13941,N_13997);
and U14083 (N_14083,N_13934,N_13936);
or U14084 (N_14084,N_13915,N_13963);
or U14085 (N_14085,N_13895,N_13931);
and U14086 (N_14086,N_13995,N_13926);
or U14087 (N_14087,N_13944,N_13888);
and U14088 (N_14088,N_13946,N_13948);
nor U14089 (N_14089,N_13885,N_13987);
nor U14090 (N_14090,N_13881,N_13926);
or U14091 (N_14091,N_13937,N_13978);
nor U14092 (N_14092,N_13995,N_13971);
nand U14093 (N_14093,N_13909,N_13972);
and U14094 (N_14094,N_13997,N_13883);
nor U14095 (N_14095,N_13908,N_13965);
nor U14096 (N_14096,N_13908,N_13930);
and U14097 (N_14097,N_13881,N_13939);
xor U14098 (N_14098,N_13913,N_13990);
and U14099 (N_14099,N_13875,N_13887);
and U14100 (N_14100,N_13938,N_13922);
xnor U14101 (N_14101,N_13987,N_13958);
xnor U14102 (N_14102,N_13967,N_13901);
nor U14103 (N_14103,N_13930,N_13955);
nor U14104 (N_14104,N_13997,N_13973);
or U14105 (N_14105,N_13943,N_13920);
nand U14106 (N_14106,N_13879,N_13878);
and U14107 (N_14107,N_13982,N_13972);
nor U14108 (N_14108,N_13954,N_13983);
or U14109 (N_14109,N_13922,N_13886);
and U14110 (N_14110,N_13948,N_13953);
or U14111 (N_14111,N_13890,N_13953);
nor U14112 (N_14112,N_13995,N_13920);
and U14113 (N_14113,N_13995,N_13912);
and U14114 (N_14114,N_13970,N_13959);
nand U14115 (N_14115,N_13993,N_13961);
and U14116 (N_14116,N_13914,N_13879);
or U14117 (N_14117,N_13947,N_13919);
nand U14118 (N_14118,N_13951,N_13950);
or U14119 (N_14119,N_13985,N_13913);
nand U14120 (N_14120,N_13940,N_13990);
xor U14121 (N_14121,N_13983,N_13918);
and U14122 (N_14122,N_13882,N_13902);
nand U14123 (N_14123,N_13957,N_13925);
or U14124 (N_14124,N_13998,N_13919);
xnor U14125 (N_14125,N_14081,N_14005);
nand U14126 (N_14126,N_14065,N_14009);
nor U14127 (N_14127,N_14045,N_14072);
nand U14128 (N_14128,N_14074,N_14117);
or U14129 (N_14129,N_14069,N_14122);
nor U14130 (N_14130,N_14036,N_14120);
nor U14131 (N_14131,N_14050,N_14107);
nor U14132 (N_14132,N_14032,N_14093);
or U14133 (N_14133,N_14018,N_14082);
and U14134 (N_14134,N_14111,N_14087);
xnor U14135 (N_14135,N_14085,N_14004);
nor U14136 (N_14136,N_14083,N_14024);
nand U14137 (N_14137,N_14030,N_14080);
nand U14138 (N_14138,N_14096,N_14100);
nor U14139 (N_14139,N_14091,N_14046);
and U14140 (N_14140,N_14031,N_14121);
nand U14141 (N_14141,N_14020,N_14021);
or U14142 (N_14142,N_14025,N_14040);
nor U14143 (N_14143,N_14098,N_14101);
nor U14144 (N_14144,N_14104,N_14061);
nor U14145 (N_14145,N_14079,N_14037);
or U14146 (N_14146,N_14113,N_14053);
nand U14147 (N_14147,N_14067,N_14095);
and U14148 (N_14148,N_14042,N_14013);
or U14149 (N_14149,N_14092,N_14114);
or U14150 (N_14150,N_14084,N_14068);
or U14151 (N_14151,N_14029,N_14066);
nand U14152 (N_14152,N_14016,N_14119);
and U14153 (N_14153,N_14123,N_14023);
nand U14154 (N_14154,N_14112,N_14051);
xnor U14155 (N_14155,N_14044,N_14110);
and U14156 (N_14156,N_14124,N_14102);
nand U14157 (N_14157,N_14010,N_14070);
xnor U14158 (N_14158,N_14106,N_14109);
nand U14159 (N_14159,N_14094,N_14056);
nor U14160 (N_14160,N_14011,N_14108);
or U14161 (N_14161,N_14003,N_14019);
xnor U14162 (N_14162,N_14052,N_14035);
and U14163 (N_14163,N_14001,N_14103);
and U14164 (N_14164,N_14014,N_14057);
nand U14165 (N_14165,N_14060,N_14041);
xor U14166 (N_14166,N_14077,N_14055);
nor U14167 (N_14167,N_14017,N_14076);
and U14168 (N_14168,N_14034,N_14038);
xnor U14169 (N_14169,N_14062,N_14033);
and U14170 (N_14170,N_14054,N_14105);
nand U14171 (N_14171,N_14058,N_14006);
or U14172 (N_14172,N_14022,N_14039);
or U14173 (N_14173,N_14115,N_14048);
and U14174 (N_14174,N_14078,N_14097);
xor U14175 (N_14175,N_14064,N_14043);
nor U14176 (N_14176,N_14073,N_14086);
and U14177 (N_14177,N_14026,N_14015);
nor U14178 (N_14178,N_14063,N_14116);
nand U14179 (N_14179,N_14049,N_14002);
or U14180 (N_14180,N_14075,N_14099);
nand U14181 (N_14181,N_14007,N_14089);
nand U14182 (N_14182,N_14027,N_14059);
or U14183 (N_14183,N_14090,N_14008);
xor U14184 (N_14184,N_14118,N_14088);
and U14185 (N_14185,N_14028,N_14000);
nand U14186 (N_14186,N_14012,N_14071);
or U14187 (N_14187,N_14047,N_14039);
or U14188 (N_14188,N_14112,N_14052);
nor U14189 (N_14189,N_14095,N_14038);
xor U14190 (N_14190,N_14046,N_14045);
or U14191 (N_14191,N_14095,N_14052);
and U14192 (N_14192,N_14066,N_14024);
and U14193 (N_14193,N_14093,N_14061);
nand U14194 (N_14194,N_14042,N_14106);
nor U14195 (N_14195,N_14001,N_14023);
nand U14196 (N_14196,N_14044,N_14033);
nor U14197 (N_14197,N_14053,N_14016);
or U14198 (N_14198,N_14083,N_14110);
nand U14199 (N_14199,N_14087,N_14098);
and U14200 (N_14200,N_14111,N_14077);
and U14201 (N_14201,N_14037,N_14035);
xnor U14202 (N_14202,N_14003,N_14087);
or U14203 (N_14203,N_14049,N_14023);
and U14204 (N_14204,N_14056,N_14074);
xor U14205 (N_14205,N_14104,N_14003);
nor U14206 (N_14206,N_14013,N_14044);
nand U14207 (N_14207,N_14090,N_14118);
nor U14208 (N_14208,N_14098,N_14007);
nand U14209 (N_14209,N_14065,N_14047);
or U14210 (N_14210,N_14085,N_14012);
or U14211 (N_14211,N_14072,N_14022);
nor U14212 (N_14212,N_14003,N_14027);
and U14213 (N_14213,N_14093,N_14094);
or U14214 (N_14214,N_14047,N_14095);
xnor U14215 (N_14215,N_14046,N_14116);
nand U14216 (N_14216,N_14008,N_14039);
nor U14217 (N_14217,N_14043,N_14042);
nand U14218 (N_14218,N_14056,N_14024);
xnor U14219 (N_14219,N_14041,N_14091);
or U14220 (N_14220,N_14064,N_14030);
nor U14221 (N_14221,N_14122,N_14096);
xnor U14222 (N_14222,N_14104,N_14035);
nor U14223 (N_14223,N_14083,N_14048);
xnor U14224 (N_14224,N_14097,N_14000);
xor U14225 (N_14225,N_14006,N_14025);
nand U14226 (N_14226,N_14078,N_14063);
xor U14227 (N_14227,N_14067,N_14071);
nor U14228 (N_14228,N_14072,N_14104);
and U14229 (N_14229,N_14093,N_14000);
nor U14230 (N_14230,N_14064,N_14091);
or U14231 (N_14231,N_14094,N_14048);
and U14232 (N_14232,N_14042,N_14022);
or U14233 (N_14233,N_14076,N_14035);
xor U14234 (N_14234,N_14011,N_14124);
nor U14235 (N_14235,N_14121,N_14106);
xnor U14236 (N_14236,N_14058,N_14069);
and U14237 (N_14237,N_14023,N_14075);
nor U14238 (N_14238,N_14122,N_14013);
or U14239 (N_14239,N_14120,N_14053);
xor U14240 (N_14240,N_14099,N_14092);
and U14241 (N_14241,N_14010,N_14045);
nand U14242 (N_14242,N_14037,N_14030);
xor U14243 (N_14243,N_14077,N_14027);
nor U14244 (N_14244,N_14079,N_14061);
nor U14245 (N_14245,N_14077,N_14013);
and U14246 (N_14246,N_14060,N_14103);
xnor U14247 (N_14247,N_14043,N_14013);
or U14248 (N_14248,N_14111,N_14056);
nand U14249 (N_14249,N_14081,N_14025);
and U14250 (N_14250,N_14233,N_14238);
nand U14251 (N_14251,N_14159,N_14231);
nor U14252 (N_14252,N_14209,N_14167);
or U14253 (N_14253,N_14165,N_14208);
nand U14254 (N_14254,N_14178,N_14179);
and U14255 (N_14255,N_14211,N_14152);
xor U14256 (N_14256,N_14151,N_14142);
nand U14257 (N_14257,N_14205,N_14184);
or U14258 (N_14258,N_14187,N_14170);
and U14259 (N_14259,N_14140,N_14162);
nor U14260 (N_14260,N_14168,N_14207);
nor U14261 (N_14261,N_14240,N_14197);
and U14262 (N_14262,N_14171,N_14200);
xor U14263 (N_14263,N_14246,N_14169);
nor U14264 (N_14264,N_14173,N_14134);
nor U14265 (N_14265,N_14181,N_14243);
xor U14266 (N_14266,N_14130,N_14236);
or U14267 (N_14267,N_14232,N_14235);
nand U14268 (N_14268,N_14180,N_14198);
and U14269 (N_14269,N_14199,N_14161);
or U14270 (N_14270,N_14242,N_14237);
or U14271 (N_14271,N_14150,N_14212);
xnor U14272 (N_14272,N_14218,N_14172);
nor U14273 (N_14273,N_14213,N_14129);
or U14274 (N_14274,N_14222,N_14202);
and U14275 (N_14275,N_14190,N_14158);
or U14276 (N_14276,N_14196,N_14177);
nor U14277 (N_14277,N_14192,N_14226);
and U14278 (N_14278,N_14146,N_14230);
and U14279 (N_14279,N_14217,N_14133);
xor U14280 (N_14280,N_14225,N_14139);
nand U14281 (N_14281,N_14160,N_14229);
xnor U14282 (N_14282,N_14174,N_14248);
nand U14283 (N_14283,N_14155,N_14201);
xor U14284 (N_14284,N_14149,N_14185);
nor U14285 (N_14285,N_14147,N_14194);
xor U14286 (N_14286,N_14215,N_14143);
or U14287 (N_14287,N_14220,N_14204);
nand U14288 (N_14288,N_14188,N_14182);
nand U14289 (N_14289,N_14137,N_14249);
nor U14290 (N_14290,N_14228,N_14244);
or U14291 (N_14291,N_14239,N_14191);
xor U14292 (N_14292,N_14221,N_14241);
xnor U14293 (N_14293,N_14163,N_14136);
or U14294 (N_14294,N_14223,N_14144);
nor U14295 (N_14295,N_14183,N_14138);
nor U14296 (N_14296,N_14216,N_14125);
and U14297 (N_14297,N_14214,N_14141);
nor U14298 (N_14298,N_14126,N_14219);
nor U14299 (N_14299,N_14164,N_14153);
xnor U14300 (N_14300,N_14206,N_14227);
or U14301 (N_14301,N_14166,N_14247);
xnor U14302 (N_14302,N_14154,N_14245);
or U14303 (N_14303,N_14186,N_14127);
xnor U14304 (N_14304,N_14176,N_14195);
nand U14305 (N_14305,N_14157,N_14128);
xnor U14306 (N_14306,N_14145,N_14135);
nand U14307 (N_14307,N_14175,N_14148);
nand U14308 (N_14308,N_14132,N_14234);
xnor U14309 (N_14309,N_14131,N_14193);
xor U14310 (N_14310,N_14224,N_14156);
or U14311 (N_14311,N_14210,N_14189);
nor U14312 (N_14312,N_14203,N_14190);
and U14313 (N_14313,N_14178,N_14175);
or U14314 (N_14314,N_14239,N_14175);
or U14315 (N_14315,N_14192,N_14222);
nor U14316 (N_14316,N_14223,N_14228);
nand U14317 (N_14317,N_14136,N_14203);
nand U14318 (N_14318,N_14161,N_14217);
nor U14319 (N_14319,N_14230,N_14136);
nand U14320 (N_14320,N_14186,N_14152);
or U14321 (N_14321,N_14247,N_14189);
xor U14322 (N_14322,N_14246,N_14166);
xor U14323 (N_14323,N_14212,N_14143);
nor U14324 (N_14324,N_14159,N_14125);
or U14325 (N_14325,N_14168,N_14244);
nand U14326 (N_14326,N_14141,N_14149);
or U14327 (N_14327,N_14206,N_14229);
nor U14328 (N_14328,N_14144,N_14199);
and U14329 (N_14329,N_14144,N_14184);
and U14330 (N_14330,N_14130,N_14191);
or U14331 (N_14331,N_14161,N_14235);
xor U14332 (N_14332,N_14238,N_14243);
and U14333 (N_14333,N_14238,N_14141);
xnor U14334 (N_14334,N_14239,N_14211);
xnor U14335 (N_14335,N_14172,N_14197);
nand U14336 (N_14336,N_14158,N_14199);
and U14337 (N_14337,N_14172,N_14211);
nand U14338 (N_14338,N_14177,N_14214);
nor U14339 (N_14339,N_14225,N_14165);
and U14340 (N_14340,N_14150,N_14181);
or U14341 (N_14341,N_14177,N_14211);
or U14342 (N_14342,N_14141,N_14240);
and U14343 (N_14343,N_14188,N_14173);
and U14344 (N_14344,N_14146,N_14139);
and U14345 (N_14345,N_14127,N_14148);
nand U14346 (N_14346,N_14219,N_14181);
and U14347 (N_14347,N_14213,N_14137);
nor U14348 (N_14348,N_14239,N_14147);
nor U14349 (N_14349,N_14185,N_14211);
and U14350 (N_14350,N_14249,N_14193);
nor U14351 (N_14351,N_14246,N_14182);
xor U14352 (N_14352,N_14127,N_14239);
nand U14353 (N_14353,N_14156,N_14143);
or U14354 (N_14354,N_14145,N_14246);
and U14355 (N_14355,N_14232,N_14162);
nor U14356 (N_14356,N_14222,N_14141);
nand U14357 (N_14357,N_14194,N_14154);
xor U14358 (N_14358,N_14140,N_14183);
nand U14359 (N_14359,N_14239,N_14173);
xnor U14360 (N_14360,N_14237,N_14154);
xor U14361 (N_14361,N_14174,N_14141);
nand U14362 (N_14362,N_14210,N_14237);
and U14363 (N_14363,N_14237,N_14151);
nor U14364 (N_14364,N_14136,N_14202);
xnor U14365 (N_14365,N_14168,N_14205);
xnor U14366 (N_14366,N_14211,N_14223);
xnor U14367 (N_14367,N_14200,N_14233);
nor U14368 (N_14368,N_14201,N_14136);
and U14369 (N_14369,N_14177,N_14169);
and U14370 (N_14370,N_14168,N_14173);
or U14371 (N_14371,N_14158,N_14135);
and U14372 (N_14372,N_14222,N_14139);
nor U14373 (N_14373,N_14186,N_14221);
xnor U14374 (N_14374,N_14211,N_14159);
xor U14375 (N_14375,N_14365,N_14313);
nand U14376 (N_14376,N_14270,N_14334);
or U14377 (N_14377,N_14358,N_14287);
or U14378 (N_14378,N_14343,N_14342);
or U14379 (N_14379,N_14308,N_14302);
nor U14380 (N_14380,N_14257,N_14332);
or U14381 (N_14381,N_14292,N_14323);
and U14382 (N_14382,N_14262,N_14279);
nor U14383 (N_14383,N_14321,N_14288);
and U14384 (N_14384,N_14344,N_14260);
or U14385 (N_14385,N_14254,N_14290);
xnor U14386 (N_14386,N_14364,N_14312);
nand U14387 (N_14387,N_14337,N_14299);
nor U14388 (N_14388,N_14267,N_14335);
xor U14389 (N_14389,N_14275,N_14258);
nor U14390 (N_14390,N_14280,N_14369);
and U14391 (N_14391,N_14372,N_14278);
or U14392 (N_14392,N_14320,N_14360);
nor U14393 (N_14393,N_14368,N_14304);
xor U14394 (N_14394,N_14329,N_14317);
or U14395 (N_14395,N_14307,N_14252);
xor U14396 (N_14396,N_14284,N_14301);
and U14397 (N_14397,N_14361,N_14354);
and U14398 (N_14398,N_14370,N_14327);
nor U14399 (N_14399,N_14314,N_14311);
nand U14400 (N_14400,N_14363,N_14300);
or U14401 (N_14401,N_14352,N_14367);
nor U14402 (N_14402,N_14346,N_14285);
or U14403 (N_14403,N_14255,N_14340);
and U14404 (N_14404,N_14263,N_14281);
nor U14405 (N_14405,N_14324,N_14336);
xnor U14406 (N_14406,N_14305,N_14298);
nor U14407 (N_14407,N_14373,N_14356);
xnor U14408 (N_14408,N_14333,N_14297);
and U14409 (N_14409,N_14250,N_14269);
xor U14410 (N_14410,N_14318,N_14341);
xor U14411 (N_14411,N_14371,N_14309);
nand U14412 (N_14412,N_14253,N_14274);
xnor U14413 (N_14413,N_14289,N_14347);
xnor U14414 (N_14414,N_14310,N_14315);
nand U14415 (N_14415,N_14350,N_14362);
or U14416 (N_14416,N_14348,N_14330);
nand U14417 (N_14417,N_14349,N_14277);
xor U14418 (N_14418,N_14296,N_14339);
or U14419 (N_14419,N_14303,N_14268);
nand U14420 (N_14420,N_14319,N_14294);
nor U14421 (N_14421,N_14306,N_14286);
nor U14422 (N_14422,N_14295,N_14345);
xor U14423 (N_14423,N_14283,N_14272);
or U14424 (N_14424,N_14326,N_14351);
or U14425 (N_14425,N_14359,N_14357);
nor U14426 (N_14426,N_14338,N_14256);
and U14427 (N_14427,N_14266,N_14273);
or U14428 (N_14428,N_14325,N_14264);
or U14429 (N_14429,N_14291,N_14282);
nand U14430 (N_14430,N_14374,N_14322);
nor U14431 (N_14431,N_14331,N_14353);
or U14432 (N_14432,N_14261,N_14259);
nand U14433 (N_14433,N_14316,N_14355);
nor U14434 (N_14434,N_14366,N_14265);
nor U14435 (N_14435,N_14251,N_14276);
xnor U14436 (N_14436,N_14328,N_14271);
and U14437 (N_14437,N_14293,N_14285);
or U14438 (N_14438,N_14309,N_14300);
or U14439 (N_14439,N_14327,N_14331);
xor U14440 (N_14440,N_14289,N_14276);
and U14441 (N_14441,N_14312,N_14276);
and U14442 (N_14442,N_14277,N_14369);
or U14443 (N_14443,N_14277,N_14321);
nand U14444 (N_14444,N_14370,N_14313);
nand U14445 (N_14445,N_14315,N_14335);
or U14446 (N_14446,N_14353,N_14356);
and U14447 (N_14447,N_14351,N_14288);
xnor U14448 (N_14448,N_14350,N_14263);
nor U14449 (N_14449,N_14284,N_14266);
and U14450 (N_14450,N_14314,N_14315);
nor U14451 (N_14451,N_14306,N_14342);
and U14452 (N_14452,N_14331,N_14267);
xnor U14453 (N_14453,N_14296,N_14307);
and U14454 (N_14454,N_14291,N_14257);
nand U14455 (N_14455,N_14363,N_14359);
and U14456 (N_14456,N_14258,N_14351);
nor U14457 (N_14457,N_14276,N_14341);
xnor U14458 (N_14458,N_14332,N_14281);
xor U14459 (N_14459,N_14278,N_14281);
and U14460 (N_14460,N_14292,N_14306);
and U14461 (N_14461,N_14357,N_14367);
xnor U14462 (N_14462,N_14312,N_14370);
and U14463 (N_14463,N_14333,N_14326);
nand U14464 (N_14464,N_14317,N_14270);
nand U14465 (N_14465,N_14325,N_14279);
nor U14466 (N_14466,N_14340,N_14327);
and U14467 (N_14467,N_14267,N_14253);
nand U14468 (N_14468,N_14357,N_14266);
xnor U14469 (N_14469,N_14275,N_14260);
nor U14470 (N_14470,N_14370,N_14254);
nor U14471 (N_14471,N_14301,N_14279);
or U14472 (N_14472,N_14295,N_14289);
nor U14473 (N_14473,N_14269,N_14284);
xnor U14474 (N_14474,N_14264,N_14313);
xor U14475 (N_14475,N_14308,N_14307);
nor U14476 (N_14476,N_14363,N_14301);
nor U14477 (N_14477,N_14331,N_14282);
xnor U14478 (N_14478,N_14345,N_14347);
nor U14479 (N_14479,N_14329,N_14307);
xor U14480 (N_14480,N_14320,N_14299);
xor U14481 (N_14481,N_14334,N_14271);
and U14482 (N_14482,N_14323,N_14260);
or U14483 (N_14483,N_14264,N_14251);
nand U14484 (N_14484,N_14313,N_14293);
xnor U14485 (N_14485,N_14278,N_14353);
xor U14486 (N_14486,N_14258,N_14343);
and U14487 (N_14487,N_14294,N_14270);
nand U14488 (N_14488,N_14355,N_14354);
and U14489 (N_14489,N_14351,N_14334);
nand U14490 (N_14490,N_14359,N_14340);
and U14491 (N_14491,N_14250,N_14347);
or U14492 (N_14492,N_14335,N_14273);
and U14493 (N_14493,N_14361,N_14281);
and U14494 (N_14494,N_14352,N_14327);
xnor U14495 (N_14495,N_14338,N_14361);
or U14496 (N_14496,N_14294,N_14348);
xor U14497 (N_14497,N_14351,N_14337);
or U14498 (N_14498,N_14336,N_14335);
and U14499 (N_14499,N_14358,N_14326);
xnor U14500 (N_14500,N_14380,N_14462);
and U14501 (N_14501,N_14392,N_14457);
nand U14502 (N_14502,N_14461,N_14493);
nor U14503 (N_14503,N_14417,N_14481);
nand U14504 (N_14504,N_14408,N_14424);
or U14505 (N_14505,N_14496,N_14459);
nor U14506 (N_14506,N_14485,N_14396);
nor U14507 (N_14507,N_14386,N_14470);
xnor U14508 (N_14508,N_14456,N_14479);
nand U14509 (N_14509,N_14406,N_14378);
xnor U14510 (N_14510,N_14497,N_14420);
or U14511 (N_14511,N_14393,N_14438);
nor U14512 (N_14512,N_14494,N_14413);
xor U14513 (N_14513,N_14458,N_14441);
xnor U14514 (N_14514,N_14465,N_14452);
and U14515 (N_14515,N_14435,N_14401);
nand U14516 (N_14516,N_14433,N_14426);
xor U14517 (N_14517,N_14454,N_14397);
xor U14518 (N_14518,N_14383,N_14476);
xnor U14519 (N_14519,N_14495,N_14416);
or U14520 (N_14520,N_14398,N_14473);
nor U14521 (N_14521,N_14487,N_14409);
nor U14522 (N_14522,N_14444,N_14423);
nor U14523 (N_14523,N_14414,N_14407);
nor U14524 (N_14524,N_14483,N_14474);
or U14525 (N_14525,N_14455,N_14419);
nor U14526 (N_14526,N_14477,N_14432);
or U14527 (N_14527,N_14490,N_14384);
or U14528 (N_14528,N_14448,N_14449);
nor U14529 (N_14529,N_14377,N_14412);
and U14530 (N_14530,N_14463,N_14427);
nand U14531 (N_14531,N_14428,N_14404);
xor U14532 (N_14532,N_14402,N_14499);
nand U14533 (N_14533,N_14415,N_14443);
xor U14534 (N_14534,N_14447,N_14430);
nor U14535 (N_14535,N_14381,N_14388);
or U14536 (N_14536,N_14421,N_14375);
and U14537 (N_14537,N_14403,N_14486);
nand U14538 (N_14538,N_14482,N_14442);
or U14539 (N_14539,N_14385,N_14446);
nor U14540 (N_14540,N_14382,N_14489);
or U14541 (N_14541,N_14471,N_14434);
xor U14542 (N_14542,N_14418,N_14467);
nor U14543 (N_14543,N_14399,N_14492);
xor U14544 (N_14544,N_14498,N_14391);
nor U14545 (N_14545,N_14439,N_14460);
or U14546 (N_14546,N_14376,N_14464);
or U14547 (N_14547,N_14379,N_14480);
xnor U14548 (N_14548,N_14491,N_14395);
and U14549 (N_14549,N_14468,N_14469);
xor U14550 (N_14550,N_14389,N_14390);
and U14551 (N_14551,N_14400,N_14440);
xor U14552 (N_14552,N_14436,N_14453);
or U14553 (N_14553,N_14445,N_14451);
and U14554 (N_14554,N_14488,N_14425);
nor U14555 (N_14555,N_14394,N_14484);
or U14556 (N_14556,N_14478,N_14450);
and U14557 (N_14557,N_14422,N_14429);
nor U14558 (N_14558,N_14472,N_14437);
nand U14559 (N_14559,N_14466,N_14405);
and U14560 (N_14560,N_14411,N_14475);
and U14561 (N_14561,N_14387,N_14431);
nor U14562 (N_14562,N_14410,N_14400);
or U14563 (N_14563,N_14390,N_14436);
nor U14564 (N_14564,N_14397,N_14496);
xnor U14565 (N_14565,N_14390,N_14403);
nand U14566 (N_14566,N_14477,N_14419);
xor U14567 (N_14567,N_14467,N_14424);
nor U14568 (N_14568,N_14457,N_14425);
xor U14569 (N_14569,N_14474,N_14465);
xor U14570 (N_14570,N_14440,N_14491);
nor U14571 (N_14571,N_14445,N_14484);
nand U14572 (N_14572,N_14407,N_14380);
nor U14573 (N_14573,N_14408,N_14445);
nor U14574 (N_14574,N_14476,N_14438);
and U14575 (N_14575,N_14461,N_14415);
nand U14576 (N_14576,N_14380,N_14392);
and U14577 (N_14577,N_14474,N_14398);
nand U14578 (N_14578,N_14375,N_14422);
xor U14579 (N_14579,N_14423,N_14419);
or U14580 (N_14580,N_14414,N_14478);
xnor U14581 (N_14581,N_14467,N_14412);
or U14582 (N_14582,N_14466,N_14454);
xnor U14583 (N_14583,N_14452,N_14473);
nor U14584 (N_14584,N_14395,N_14383);
nand U14585 (N_14585,N_14444,N_14412);
or U14586 (N_14586,N_14423,N_14403);
xor U14587 (N_14587,N_14424,N_14476);
xnor U14588 (N_14588,N_14384,N_14424);
or U14589 (N_14589,N_14444,N_14486);
and U14590 (N_14590,N_14378,N_14400);
and U14591 (N_14591,N_14447,N_14388);
or U14592 (N_14592,N_14472,N_14482);
xor U14593 (N_14593,N_14432,N_14389);
or U14594 (N_14594,N_14401,N_14404);
or U14595 (N_14595,N_14436,N_14468);
xnor U14596 (N_14596,N_14403,N_14437);
nand U14597 (N_14597,N_14410,N_14461);
or U14598 (N_14598,N_14432,N_14447);
and U14599 (N_14599,N_14431,N_14435);
xnor U14600 (N_14600,N_14467,N_14446);
and U14601 (N_14601,N_14458,N_14451);
nor U14602 (N_14602,N_14477,N_14450);
nor U14603 (N_14603,N_14404,N_14422);
xor U14604 (N_14604,N_14415,N_14397);
or U14605 (N_14605,N_14445,N_14450);
and U14606 (N_14606,N_14380,N_14485);
nor U14607 (N_14607,N_14395,N_14435);
nor U14608 (N_14608,N_14393,N_14479);
nand U14609 (N_14609,N_14420,N_14430);
xor U14610 (N_14610,N_14499,N_14493);
or U14611 (N_14611,N_14453,N_14411);
and U14612 (N_14612,N_14473,N_14390);
xnor U14613 (N_14613,N_14418,N_14442);
xnor U14614 (N_14614,N_14389,N_14439);
nand U14615 (N_14615,N_14481,N_14427);
and U14616 (N_14616,N_14448,N_14459);
xnor U14617 (N_14617,N_14458,N_14423);
nand U14618 (N_14618,N_14384,N_14449);
or U14619 (N_14619,N_14375,N_14416);
nand U14620 (N_14620,N_14429,N_14406);
xnor U14621 (N_14621,N_14482,N_14382);
xnor U14622 (N_14622,N_14394,N_14417);
or U14623 (N_14623,N_14377,N_14495);
nor U14624 (N_14624,N_14478,N_14456);
nand U14625 (N_14625,N_14536,N_14568);
or U14626 (N_14626,N_14501,N_14591);
nor U14627 (N_14627,N_14590,N_14537);
or U14628 (N_14628,N_14508,N_14592);
nor U14629 (N_14629,N_14517,N_14524);
or U14630 (N_14630,N_14594,N_14566);
and U14631 (N_14631,N_14526,N_14525);
or U14632 (N_14632,N_14576,N_14613);
xnor U14633 (N_14633,N_14543,N_14552);
nand U14634 (N_14634,N_14504,N_14582);
and U14635 (N_14635,N_14606,N_14500);
and U14636 (N_14636,N_14503,N_14528);
nor U14637 (N_14637,N_14527,N_14575);
and U14638 (N_14638,N_14541,N_14614);
nand U14639 (N_14639,N_14580,N_14587);
xnor U14640 (N_14640,N_14619,N_14588);
and U14641 (N_14641,N_14565,N_14596);
xnor U14642 (N_14642,N_14540,N_14547);
or U14643 (N_14643,N_14549,N_14512);
xnor U14644 (N_14644,N_14583,N_14520);
nand U14645 (N_14645,N_14581,N_14554);
or U14646 (N_14646,N_14607,N_14521);
xnor U14647 (N_14647,N_14509,N_14544);
and U14648 (N_14648,N_14564,N_14553);
xnor U14649 (N_14649,N_14622,N_14593);
nor U14650 (N_14650,N_14522,N_14585);
or U14651 (N_14651,N_14542,N_14609);
nor U14652 (N_14652,N_14618,N_14621);
or U14653 (N_14653,N_14538,N_14567);
or U14654 (N_14654,N_14558,N_14595);
nand U14655 (N_14655,N_14506,N_14573);
nor U14656 (N_14656,N_14608,N_14620);
and U14657 (N_14657,N_14577,N_14570);
and U14658 (N_14658,N_14556,N_14589);
nand U14659 (N_14659,N_14605,N_14515);
nand U14660 (N_14660,N_14615,N_14530);
nor U14661 (N_14661,N_14616,N_14604);
nor U14662 (N_14662,N_14557,N_14599);
and U14663 (N_14663,N_14563,N_14561);
xor U14664 (N_14664,N_14529,N_14555);
nor U14665 (N_14665,N_14578,N_14533);
nand U14666 (N_14666,N_14569,N_14603);
and U14667 (N_14667,N_14612,N_14531);
or U14668 (N_14668,N_14546,N_14548);
nand U14669 (N_14669,N_14562,N_14617);
nor U14670 (N_14670,N_14518,N_14602);
and U14671 (N_14671,N_14534,N_14502);
xor U14672 (N_14672,N_14598,N_14601);
and U14673 (N_14673,N_14532,N_14545);
or U14674 (N_14674,N_14584,N_14571);
or U14675 (N_14675,N_14611,N_14574);
nor U14676 (N_14676,N_14579,N_14510);
nand U14677 (N_14677,N_14505,N_14539);
nor U14678 (N_14678,N_14623,N_14586);
and U14679 (N_14679,N_14516,N_14519);
and U14680 (N_14680,N_14507,N_14535);
or U14681 (N_14681,N_14551,N_14610);
nor U14682 (N_14682,N_14511,N_14550);
nand U14683 (N_14683,N_14597,N_14600);
nand U14684 (N_14684,N_14523,N_14559);
xnor U14685 (N_14685,N_14514,N_14572);
nand U14686 (N_14686,N_14624,N_14560);
nand U14687 (N_14687,N_14513,N_14558);
nand U14688 (N_14688,N_14541,N_14556);
or U14689 (N_14689,N_14574,N_14607);
or U14690 (N_14690,N_14615,N_14533);
or U14691 (N_14691,N_14527,N_14505);
nor U14692 (N_14692,N_14556,N_14581);
xnor U14693 (N_14693,N_14526,N_14582);
nand U14694 (N_14694,N_14603,N_14533);
and U14695 (N_14695,N_14503,N_14516);
and U14696 (N_14696,N_14602,N_14615);
and U14697 (N_14697,N_14541,N_14521);
and U14698 (N_14698,N_14599,N_14549);
nor U14699 (N_14699,N_14596,N_14603);
or U14700 (N_14700,N_14603,N_14536);
xnor U14701 (N_14701,N_14520,N_14542);
nor U14702 (N_14702,N_14609,N_14530);
and U14703 (N_14703,N_14540,N_14526);
nor U14704 (N_14704,N_14524,N_14603);
xor U14705 (N_14705,N_14540,N_14579);
nor U14706 (N_14706,N_14582,N_14593);
xnor U14707 (N_14707,N_14546,N_14519);
nand U14708 (N_14708,N_14598,N_14589);
or U14709 (N_14709,N_14583,N_14534);
or U14710 (N_14710,N_14570,N_14579);
xnor U14711 (N_14711,N_14604,N_14513);
nand U14712 (N_14712,N_14514,N_14590);
nand U14713 (N_14713,N_14528,N_14569);
xnor U14714 (N_14714,N_14549,N_14580);
nand U14715 (N_14715,N_14597,N_14555);
or U14716 (N_14716,N_14541,N_14603);
nor U14717 (N_14717,N_14582,N_14520);
nor U14718 (N_14718,N_14529,N_14585);
nor U14719 (N_14719,N_14500,N_14595);
nand U14720 (N_14720,N_14516,N_14548);
nand U14721 (N_14721,N_14588,N_14560);
or U14722 (N_14722,N_14546,N_14557);
or U14723 (N_14723,N_14596,N_14504);
xnor U14724 (N_14724,N_14598,N_14587);
and U14725 (N_14725,N_14617,N_14613);
xnor U14726 (N_14726,N_14506,N_14503);
nand U14727 (N_14727,N_14501,N_14553);
nand U14728 (N_14728,N_14505,N_14574);
nor U14729 (N_14729,N_14508,N_14624);
xnor U14730 (N_14730,N_14548,N_14510);
and U14731 (N_14731,N_14510,N_14581);
nand U14732 (N_14732,N_14537,N_14536);
nand U14733 (N_14733,N_14515,N_14617);
xnor U14734 (N_14734,N_14506,N_14587);
xor U14735 (N_14735,N_14522,N_14511);
nor U14736 (N_14736,N_14510,N_14557);
nand U14737 (N_14737,N_14540,N_14550);
or U14738 (N_14738,N_14589,N_14516);
xor U14739 (N_14739,N_14558,N_14573);
nand U14740 (N_14740,N_14588,N_14572);
xor U14741 (N_14741,N_14517,N_14589);
nor U14742 (N_14742,N_14584,N_14505);
nand U14743 (N_14743,N_14603,N_14546);
and U14744 (N_14744,N_14530,N_14571);
nand U14745 (N_14745,N_14594,N_14552);
and U14746 (N_14746,N_14509,N_14569);
and U14747 (N_14747,N_14534,N_14539);
nand U14748 (N_14748,N_14533,N_14502);
nand U14749 (N_14749,N_14541,N_14624);
and U14750 (N_14750,N_14706,N_14713);
nor U14751 (N_14751,N_14698,N_14679);
xor U14752 (N_14752,N_14634,N_14662);
and U14753 (N_14753,N_14716,N_14673);
nand U14754 (N_14754,N_14636,N_14687);
xor U14755 (N_14755,N_14633,N_14709);
nand U14756 (N_14756,N_14629,N_14663);
nor U14757 (N_14757,N_14643,N_14727);
nand U14758 (N_14758,N_14671,N_14735);
nor U14759 (N_14759,N_14748,N_14726);
nand U14760 (N_14760,N_14642,N_14667);
xnor U14761 (N_14761,N_14690,N_14696);
or U14762 (N_14762,N_14734,N_14637);
nand U14763 (N_14763,N_14725,N_14689);
nand U14764 (N_14764,N_14675,N_14659);
nand U14765 (N_14765,N_14658,N_14740);
and U14766 (N_14766,N_14627,N_14743);
and U14767 (N_14767,N_14656,N_14638);
or U14768 (N_14768,N_14641,N_14652);
xor U14769 (N_14769,N_14632,N_14670);
xor U14770 (N_14770,N_14708,N_14686);
nand U14771 (N_14771,N_14721,N_14651);
nand U14772 (N_14772,N_14718,N_14684);
nor U14773 (N_14773,N_14742,N_14647);
or U14774 (N_14774,N_14700,N_14682);
and U14775 (N_14775,N_14715,N_14646);
nor U14776 (N_14776,N_14699,N_14674);
xor U14777 (N_14777,N_14732,N_14668);
or U14778 (N_14778,N_14719,N_14714);
nand U14779 (N_14779,N_14695,N_14640);
nor U14780 (N_14780,N_14683,N_14648);
or U14781 (N_14781,N_14717,N_14661);
nand U14782 (N_14782,N_14707,N_14676);
nor U14783 (N_14783,N_14681,N_14693);
xor U14784 (N_14784,N_14657,N_14720);
nor U14785 (N_14785,N_14664,N_14625);
nand U14786 (N_14786,N_14702,N_14738);
xnor U14787 (N_14787,N_14731,N_14630);
nor U14788 (N_14788,N_14712,N_14728);
and U14789 (N_14789,N_14691,N_14736);
xor U14790 (N_14790,N_14697,N_14654);
and U14791 (N_14791,N_14649,N_14729);
nand U14792 (N_14792,N_14703,N_14628);
and U14793 (N_14793,N_14705,N_14730);
xnor U14794 (N_14794,N_14677,N_14665);
nor U14795 (N_14795,N_14672,N_14680);
xnor U14796 (N_14796,N_14722,N_14678);
or U14797 (N_14797,N_14711,N_14688);
nand U14798 (N_14798,N_14666,N_14724);
nor U14799 (N_14799,N_14746,N_14626);
xor U14800 (N_14800,N_14660,N_14741);
xor U14801 (N_14801,N_14739,N_14631);
xor U14802 (N_14802,N_14653,N_14747);
or U14803 (N_14803,N_14669,N_14723);
xor U14804 (N_14804,N_14639,N_14635);
xor U14805 (N_14805,N_14685,N_14704);
xor U14806 (N_14806,N_14645,N_14745);
xnor U14807 (N_14807,N_14710,N_14744);
or U14808 (N_14808,N_14737,N_14749);
and U14809 (N_14809,N_14650,N_14694);
and U14810 (N_14810,N_14692,N_14655);
and U14811 (N_14811,N_14701,N_14733);
nand U14812 (N_14812,N_14644,N_14748);
and U14813 (N_14813,N_14680,N_14626);
or U14814 (N_14814,N_14658,N_14691);
nand U14815 (N_14815,N_14674,N_14680);
or U14816 (N_14816,N_14716,N_14683);
xor U14817 (N_14817,N_14728,N_14708);
or U14818 (N_14818,N_14721,N_14747);
or U14819 (N_14819,N_14629,N_14738);
nor U14820 (N_14820,N_14741,N_14661);
xor U14821 (N_14821,N_14679,N_14658);
xor U14822 (N_14822,N_14744,N_14724);
nand U14823 (N_14823,N_14668,N_14737);
nand U14824 (N_14824,N_14655,N_14733);
nor U14825 (N_14825,N_14667,N_14655);
nor U14826 (N_14826,N_14744,N_14640);
or U14827 (N_14827,N_14686,N_14646);
nor U14828 (N_14828,N_14713,N_14627);
and U14829 (N_14829,N_14672,N_14625);
xnor U14830 (N_14830,N_14642,N_14668);
nand U14831 (N_14831,N_14703,N_14657);
and U14832 (N_14832,N_14668,N_14702);
nor U14833 (N_14833,N_14705,N_14701);
nand U14834 (N_14834,N_14718,N_14663);
or U14835 (N_14835,N_14663,N_14700);
nand U14836 (N_14836,N_14693,N_14677);
nor U14837 (N_14837,N_14644,N_14652);
or U14838 (N_14838,N_14713,N_14746);
and U14839 (N_14839,N_14695,N_14639);
nand U14840 (N_14840,N_14648,N_14655);
or U14841 (N_14841,N_14709,N_14646);
xnor U14842 (N_14842,N_14744,N_14743);
nand U14843 (N_14843,N_14665,N_14731);
and U14844 (N_14844,N_14746,N_14659);
or U14845 (N_14845,N_14667,N_14676);
nor U14846 (N_14846,N_14719,N_14725);
nor U14847 (N_14847,N_14697,N_14678);
nor U14848 (N_14848,N_14683,N_14700);
or U14849 (N_14849,N_14733,N_14693);
nor U14850 (N_14850,N_14729,N_14715);
xnor U14851 (N_14851,N_14714,N_14648);
nand U14852 (N_14852,N_14649,N_14720);
or U14853 (N_14853,N_14711,N_14662);
nand U14854 (N_14854,N_14648,N_14637);
or U14855 (N_14855,N_14727,N_14682);
and U14856 (N_14856,N_14723,N_14711);
and U14857 (N_14857,N_14634,N_14658);
and U14858 (N_14858,N_14651,N_14676);
or U14859 (N_14859,N_14672,N_14740);
and U14860 (N_14860,N_14688,N_14736);
or U14861 (N_14861,N_14648,N_14652);
and U14862 (N_14862,N_14718,N_14692);
nor U14863 (N_14863,N_14680,N_14731);
or U14864 (N_14864,N_14735,N_14706);
xor U14865 (N_14865,N_14733,N_14662);
or U14866 (N_14866,N_14696,N_14733);
and U14867 (N_14867,N_14648,N_14693);
xnor U14868 (N_14868,N_14682,N_14712);
xnor U14869 (N_14869,N_14625,N_14710);
and U14870 (N_14870,N_14726,N_14708);
or U14871 (N_14871,N_14722,N_14724);
xor U14872 (N_14872,N_14659,N_14736);
or U14873 (N_14873,N_14716,N_14742);
xor U14874 (N_14874,N_14706,N_14652);
xor U14875 (N_14875,N_14788,N_14754);
or U14876 (N_14876,N_14751,N_14752);
nor U14877 (N_14877,N_14761,N_14807);
xnor U14878 (N_14878,N_14873,N_14764);
nand U14879 (N_14879,N_14773,N_14818);
xnor U14880 (N_14880,N_14862,N_14750);
nor U14881 (N_14881,N_14860,N_14838);
nand U14882 (N_14882,N_14869,N_14817);
and U14883 (N_14883,N_14847,N_14796);
xnor U14884 (N_14884,N_14806,N_14768);
or U14885 (N_14885,N_14782,N_14874);
nand U14886 (N_14886,N_14845,N_14783);
xnor U14887 (N_14887,N_14852,N_14819);
and U14888 (N_14888,N_14836,N_14767);
nor U14889 (N_14889,N_14861,N_14822);
nor U14890 (N_14890,N_14795,N_14849);
nor U14891 (N_14891,N_14853,N_14824);
or U14892 (N_14892,N_14835,N_14801);
xor U14893 (N_14893,N_14780,N_14839);
nand U14894 (N_14894,N_14864,N_14759);
nand U14895 (N_14895,N_14774,N_14805);
and U14896 (N_14896,N_14810,N_14809);
and U14897 (N_14897,N_14855,N_14800);
and U14898 (N_14898,N_14770,N_14785);
and U14899 (N_14899,N_14794,N_14816);
xnor U14900 (N_14900,N_14828,N_14763);
and U14901 (N_14901,N_14840,N_14856);
nand U14902 (N_14902,N_14863,N_14789);
nor U14903 (N_14903,N_14846,N_14766);
and U14904 (N_14904,N_14867,N_14753);
xor U14905 (N_14905,N_14790,N_14833);
nand U14906 (N_14906,N_14808,N_14776);
nor U14907 (N_14907,N_14812,N_14786);
xor U14908 (N_14908,N_14813,N_14866);
xnor U14909 (N_14909,N_14850,N_14755);
nand U14910 (N_14910,N_14827,N_14823);
nand U14911 (N_14911,N_14811,N_14857);
nand U14912 (N_14912,N_14865,N_14843);
xnor U14913 (N_14913,N_14769,N_14792);
or U14914 (N_14914,N_14804,N_14765);
xnor U14915 (N_14915,N_14851,N_14837);
nor U14916 (N_14916,N_14771,N_14781);
or U14917 (N_14917,N_14830,N_14772);
nand U14918 (N_14918,N_14775,N_14784);
and U14919 (N_14919,N_14799,N_14815);
xor U14920 (N_14920,N_14757,N_14777);
and U14921 (N_14921,N_14821,N_14842);
nor U14922 (N_14922,N_14798,N_14756);
or U14923 (N_14923,N_14820,N_14778);
and U14924 (N_14924,N_14814,N_14762);
nor U14925 (N_14925,N_14868,N_14802);
nand U14926 (N_14926,N_14841,N_14803);
and U14927 (N_14927,N_14844,N_14832);
xor U14928 (N_14928,N_14779,N_14826);
nor U14929 (N_14929,N_14859,N_14854);
nand U14930 (N_14930,N_14871,N_14793);
and U14931 (N_14931,N_14858,N_14834);
nand U14932 (N_14932,N_14831,N_14758);
and U14933 (N_14933,N_14760,N_14829);
and U14934 (N_14934,N_14791,N_14787);
or U14935 (N_14935,N_14797,N_14825);
xnor U14936 (N_14936,N_14848,N_14870);
nor U14937 (N_14937,N_14872,N_14816);
or U14938 (N_14938,N_14802,N_14797);
or U14939 (N_14939,N_14781,N_14805);
nand U14940 (N_14940,N_14816,N_14786);
nand U14941 (N_14941,N_14874,N_14829);
or U14942 (N_14942,N_14844,N_14817);
and U14943 (N_14943,N_14783,N_14778);
and U14944 (N_14944,N_14754,N_14805);
and U14945 (N_14945,N_14787,N_14851);
xor U14946 (N_14946,N_14838,N_14863);
xor U14947 (N_14947,N_14852,N_14872);
xor U14948 (N_14948,N_14848,N_14829);
nand U14949 (N_14949,N_14755,N_14833);
nor U14950 (N_14950,N_14755,N_14769);
or U14951 (N_14951,N_14823,N_14795);
xnor U14952 (N_14952,N_14756,N_14870);
nor U14953 (N_14953,N_14790,N_14846);
or U14954 (N_14954,N_14769,N_14778);
nor U14955 (N_14955,N_14852,N_14800);
nand U14956 (N_14956,N_14769,N_14816);
and U14957 (N_14957,N_14796,N_14810);
xor U14958 (N_14958,N_14751,N_14814);
xnor U14959 (N_14959,N_14861,N_14856);
nor U14960 (N_14960,N_14782,N_14798);
and U14961 (N_14961,N_14839,N_14850);
xnor U14962 (N_14962,N_14806,N_14820);
nand U14963 (N_14963,N_14773,N_14762);
nand U14964 (N_14964,N_14781,N_14863);
nor U14965 (N_14965,N_14772,N_14853);
nor U14966 (N_14966,N_14865,N_14791);
and U14967 (N_14967,N_14783,N_14802);
nand U14968 (N_14968,N_14855,N_14756);
and U14969 (N_14969,N_14838,N_14803);
xor U14970 (N_14970,N_14851,N_14814);
or U14971 (N_14971,N_14781,N_14761);
nand U14972 (N_14972,N_14751,N_14860);
and U14973 (N_14973,N_14811,N_14845);
nand U14974 (N_14974,N_14756,N_14818);
nor U14975 (N_14975,N_14872,N_14855);
or U14976 (N_14976,N_14779,N_14750);
or U14977 (N_14977,N_14806,N_14838);
or U14978 (N_14978,N_14844,N_14770);
xor U14979 (N_14979,N_14829,N_14838);
and U14980 (N_14980,N_14835,N_14854);
nand U14981 (N_14981,N_14779,N_14798);
and U14982 (N_14982,N_14768,N_14766);
nand U14983 (N_14983,N_14841,N_14786);
nor U14984 (N_14984,N_14806,N_14756);
nand U14985 (N_14985,N_14861,N_14809);
or U14986 (N_14986,N_14819,N_14806);
and U14987 (N_14987,N_14857,N_14833);
or U14988 (N_14988,N_14844,N_14837);
nor U14989 (N_14989,N_14755,N_14799);
and U14990 (N_14990,N_14756,N_14824);
nor U14991 (N_14991,N_14874,N_14822);
xnor U14992 (N_14992,N_14859,N_14772);
nor U14993 (N_14993,N_14840,N_14862);
and U14994 (N_14994,N_14859,N_14840);
and U14995 (N_14995,N_14781,N_14840);
nor U14996 (N_14996,N_14804,N_14860);
nor U14997 (N_14997,N_14767,N_14756);
nand U14998 (N_14998,N_14828,N_14855);
nand U14999 (N_14999,N_14871,N_14850);
or UO_0 (O_0,N_14916,N_14986);
nand UO_1 (O_1,N_14891,N_14960);
and UO_2 (O_2,N_14983,N_14918);
nand UO_3 (O_3,N_14887,N_14928);
and UO_4 (O_4,N_14990,N_14926);
nand UO_5 (O_5,N_14875,N_14957);
nor UO_6 (O_6,N_14884,N_14956);
xor UO_7 (O_7,N_14921,N_14915);
or UO_8 (O_8,N_14896,N_14944);
xnor UO_9 (O_9,N_14964,N_14978);
nor UO_10 (O_10,N_14922,N_14999);
xor UO_11 (O_11,N_14967,N_14985);
and UO_12 (O_12,N_14908,N_14946);
nand UO_13 (O_13,N_14933,N_14973);
nand UO_14 (O_14,N_14894,N_14919);
nand UO_15 (O_15,N_14996,N_14976);
nor UO_16 (O_16,N_14880,N_14959);
xor UO_17 (O_17,N_14877,N_14937);
xnor UO_18 (O_18,N_14900,N_14989);
nand UO_19 (O_19,N_14958,N_14906);
nand UO_20 (O_20,N_14923,N_14950);
nand UO_21 (O_21,N_14941,N_14987);
nand UO_22 (O_22,N_14925,N_14905);
xor UO_23 (O_23,N_14998,N_14947);
nor UO_24 (O_24,N_14924,N_14943);
nand UO_25 (O_25,N_14901,N_14980);
xor UO_26 (O_26,N_14904,N_14979);
nor UO_27 (O_27,N_14914,N_14886);
nor UO_28 (O_28,N_14907,N_14942);
and UO_29 (O_29,N_14997,N_14951);
nor UO_30 (O_30,N_14954,N_14889);
nand UO_31 (O_31,N_14882,N_14932);
xor UO_32 (O_32,N_14949,N_14961);
xor UO_33 (O_33,N_14984,N_14963);
xor UO_34 (O_34,N_14988,N_14948);
nor UO_35 (O_35,N_14927,N_14940);
and UO_36 (O_36,N_14892,N_14883);
and UO_37 (O_37,N_14992,N_14991);
or UO_38 (O_38,N_14930,N_14935);
nand UO_39 (O_39,N_14929,N_14934);
xor UO_40 (O_40,N_14917,N_14945);
and UO_41 (O_41,N_14962,N_14970);
xnor UO_42 (O_42,N_14920,N_14895);
xor UO_43 (O_43,N_14893,N_14912);
and UO_44 (O_44,N_14938,N_14890);
or UO_45 (O_45,N_14936,N_14981);
nor UO_46 (O_46,N_14910,N_14965);
xnor UO_47 (O_47,N_14977,N_14931);
xnor UO_48 (O_48,N_14953,N_14971);
xor UO_49 (O_49,N_14902,N_14881);
nor UO_50 (O_50,N_14903,N_14911);
xor UO_51 (O_51,N_14972,N_14982);
xor UO_52 (O_52,N_14879,N_14994);
and UO_53 (O_53,N_14885,N_14968);
and UO_54 (O_54,N_14952,N_14888);
or UO_55 (O_55,N_14897,N_14898);
xor UO_56 (O_56,N_14995,N_14955);
nand UO_57 (O_57,N_14909,N_14939);
xnor UO_58 (O_58,N_14899,N_14878);
xnor UO_59 (O_59,N_14975,N_14913);
or UO_60 (O_60,N_14876,N_14993);
xnor UO_61 (O_61,N_14969,N_14974);
and UO_62 (O_62,N_14966,N_14994);
xor UO_63 (O_63,N_14985,N_14978);
or UO_64 (O_64,N_14931,N_14998);
nor UO_65 (O_65,N_14946,N_14941);
and UO_66 (O_66,N_14963,N_14972);
xnor UO_67 (O_67,N_14979,N_14921);
or UO_68 (O_68,N_14919,N_14979);
nor UO_69 (O_69,N_14884,N_14913);
and UO_70 (O_70,N_14941,N_14970);
and UO_71 (O_71,N_14931,N_14902);
or UO_72 (O_72,N_14935,N_14980);
and UO_73 (O_73,N_14900,N_14883);
xnor UO_74 (O_74,N_14986,N_14949);
xor UO_75 (O_75,N_14994,N_14891);
or UO_76 (O_76,N_14988,N_14897);
and UO_77 (O_77,N_14963,N_14911);
xnor UO_78 (O_78,N_14963,N_14945);
or UO_79 (O_79,N_14958,N_14983);
nand UO_80 (O_80,N_14971,N_14889);
and UO_81 (O_81,N_14915,N_14953);
nor UO_82 (O_82,N_14952,N_14985);
nand UO_83 (O_83,N_14891,N_14898);
nor UO_84 (O_84,N_14876,N_14878);
xor UO_85 (O_85,N_14964,N_14891);
xor UO_86 (O_86,N_14954,N_14904);
and UO_87 (O_87,N_14917,N_14925);
nor UO_88 (O_88,N_14976,N_14887);
and UO_89 (O_89,N_14923,N_14934);
xor UO_90 (O_90,N_14952,N_14917);
xnor UO_91 (O_91,N_14947,N_14892);
xor UO_92 (O_92,N_14896,N_14960);
nor UO_93 (O_93,N_14975,N_14962);
xnor UO_94 (O_94,N_14950,N_14936);
nor UO_95 (O_95,N_14947,N_14954);
nor UO_96 (O_96,N_14950,N_14879);
and UO_97 (O_97,N_14879,N_14962);
and UO_98 (O_98,N_14879,N_14977);
nor UO_99 (O_99,N_14916,N_14984);
xnor UO_100 (O_100,N_14918,N_14962);
xnor UO_101 (O_101,N_14915,N_14891);
nand UO_102 (O_102,N_14887,N_14948);
nor UO_103 (O_103,N_14883,N_14920);
xnor UO_104 (O_104,N_14982,N_14923);
and UO_105 (O_105,N_14924,N_14933);
nor UO_106 (O_106,N_14931,N_14973);
nand UO_107 (O_107,N_14998,N_14943);
and UO_108 (O_108,N_14972,N_14936);
nand UO_109 (O_109,N_14908,N_14983);
xnor UO_110 (O_110,N_14927,N_14943);
nand UO_111 (O_111,N_14877,N_14892);
and UO_112 (O_112,N_14912,N_14990);
xnor UO_113 (O_113,N_14934,N_14921);
nand UO_114 (O_114,N_14912,N_14949);
and UO_115 (O_115,N_14933,N_14962);
and UO_116 (O_116,N_14917,N_14983);
nor UO_117 (O_117,N_14892,N_14893);
xor UO_118 (O_118,N_14976,N_14880);
xnor UO_119 (O_119,N_14943,N_14966);
or UO_120 (O_120,N_14968,N_14974);
xor UO_121 (O_121,N_14936,N_14905);
xor UO_122 (O_122,N_14927,N_14892);
and UO_123 (O_123,N_14947,N_14976);
xor UO_124 (O_124,N_14980,N_14970);
xor UO_125 (O_125,N_14885,N_14936);
and UO_126 (O_126,N_14909,N_14990);
or UO_127 (O_127,N_14981,N_14995);
or UO_128 (O_128,N_14891,N_14939);
nor UO_129 (O_129,N_14988,N_14878);
nor UO_130 (O_130,N_14900,N_14887);
and UO_131 (O_131,N_14880,N_14904);
nor UO_132 (O_132,N_14985,N_14933);
nor UO_133 (O_133,N_14995,N_14960);
or UO_134 (O_134,N_14958,N_14949);
nand UO_135 (O_135,N_14954,N_14942);
nor UO_136 (O_136,N_14919,N_14935);
nand UO_137 (O_137,N_14971,N_14897);
and UO_138 (O_138,N_14981,N_14917);
and UO_139 (O_139,N_14904,N_14902);
nor UO_140 (O_140,N_14958,N_14934);
or UO_141 (O_141,N_14983,N_14912);
xnor UO_142 (O_142,N_14877,N_14994);
and UO_143 (O_143,N_14917,N_14919);
nor UO_144 (O_144,N_14988,N_14980);
and UO_145 (O_145,N_14895,N_14907);
nand UO_146 (O_146,N_14919,N_14931);
xnor UO_147 (O_147,N_14903,N_14972);
xor UO_148 (O_148,N_14925,N_14927);
or UO_149 (O_149,N_14886,N_14922);
xor UO_150 (O_150,N_14904,N_14924);
and UO_151 (O_151,N_14953,N_14928);
nor UO_152 (O_152,N_14962,N_14988);
xnor UO_153 (O_153,N_14885,N_14950);
nor UO_154 (O_154,N_14897,N_14939);
and UO_155 (O_155,N_14882,N_14914);
or UO_156 (O_156,N_14901,N_14935);
and UO_157 (O_157,N_14905,N_14904);
nor UO_158 (O_158,N_14989,N_14901);
or UO_159 (O_159,N_14900,N_14923);
nor UO_160 (O_160,N_14981,N_14950);
and UO_161 (O_161,N_14952,N_14962);
xor UO_162 (O_162,N_14982,N_14910);
nor UO_163 (O_163,N_14984,N_14947);
xnor UO_164 (O_164,N_14970,N_14935);
or UO_165 (O_165,N_14887,N_14984);
nor UO_166 (O_166,N_14932,N_14947);
nor UO_167 (O_167,N_14995,N_14877);
and UO_168 (O_168,N_14925,N_14964);
or UO_169 (O_169,N_14910,N_14887);
nand UO_170 (O_170,N_14972,N_14921);
or UO_171 (O_171,N_14999,N_14987);
xor UO_172 (O_172,N_14991,N_14890);
nand UO_173 (O_173,N_14926,N_14998);
nor UO_174 (O_174,N_14961,N_14947);
or UO_175 (O_175,N_14969,N_14948);
and UO_176 (O_176,N_14982,N_14983);
nor UO_177 (O_177,N_14951,N_14906);
and UO_178 (O_178,N_14877,N_14963);
and UO_179 (O_179,N_14879,N_14918);
or UO_180 (O_180,N_14952,N_14970);
and UO_181 (O_181,N_14965,N_14977);
nor UO_182 (O_182,N_14977,N_14985);
and UO_183 (O_183,N_14980,N_14950);
and UO_184 (O_184,N_14967,N_14892);
or UO_185 (O_185,N_14969,N_14888);
or UO_186 (O_186,N_14881,N_14983);
and UO_187 (O_187,N_14915,N_14946);
nand UO_188 (O_188,N_14877,N_14912);
nand UO_189 (O_189,N_14926,N_14922);
xor UO_190 (O_190,N_14891,N_14886);
and UO_191 (O_191,N_14886,N_14898);
nand UO_192 (O_192,N_14883,N_14888);
or UO_193 (O_193,N_14957,N_14878);
and UO_194 (O_194,N_14899,N_14949);
xor UO_195 (O_195,N_14936,N_14903);
and UO_196 (O_196,N_14981,N_14972);
and UO_197 (O_197,N_14886,N_14944);
or UO_198 (O_198,N_14996,N_14985);
or UO_199 (O_199,N_14887,N_14905);
nand UO_200 (O_200,N_14928,N_14918);
or UO_201 (O_201,N_14966,N_14919);
xnor UO_202 (O_202,N_14997,N_14966);
nor UO_203 (O_203,N_14933,N_14944);
xnor UO_204 (O_204,N_14920,N_14876);
xor UO_205 (O_205,N_14999,N_14893);
nor UO_206 (O_206,N_14906,N_14961);
and UO_207 (O_207,N_14981,N_14973);
nor UO_208 (O_208,N_14977,N_14967);
nor UO_209 (O_209,N_14977,N_14976);
or UO_210 (O_210,N_14962,N_14969);
nor UO_211 (O_211,N_14946,N_14878);
xor UO_212 (O_212,N_14901,N_14893);
and UO_213 (O_213,N_14886,N_14980);
or UO_214 (O_214,N_14890,N_14996);
nor UO_215 (O_215,N_14963,N_14983);
nand UO_216 (O_216,N_14972,N_14968);
xor UO_217 (O_217,N_14997,N_14897);
or UO_218 (O_218,N_14934,N_14905);
nand UO_219 (O_219,N_14967,N_14996);
and UO_220 (O_220,N_14877,N_14920);
nand UO_221 (O_221,N_14951,N_14964);
nand UO_222 (O_222,N_14963,N_14888);
and UO_223 (O_223,N_14925,N_14947);
or UO_224 (O_224,N_14941,N_14913);
nand UO_225 (O_225,N_14941,N_14909);
and UO_226 (O_226,N_14933,N_14893);
nor UO_227 (O_227,N_14972,N_14939);
and UO_228 (O_228,N_14981,N_14878);
nor UO_229 (O_229,N_14987,N_14910);
nor UO_230 (O_230,N_14927,N_14976);
xor UO_231 (O_231,N_14989,N_14986);
nor UO_232 (O_232,N_14957,N_14892);
nand UO_233 (O_233,N_14980,N_14972);
or UO_234 (O_234,N_14960,N_14913);
nand UO_235 (O_235,N_14928,N_14890);
and UO_236 (O_236,N_14886,N_14921);
nand UO_237 (O_237,N_14979,N_14984);
xor UO_238 (O_238,N_14912,N_14956);
nor UO_239 (O_239,N_14902,N_14966);
and UO_240 (O_240,N_14916,N_14997);
and UO_241 (O_241,N_14999,N_14995);
nand UO_242 (O_242,N_14969,N_14881);
nand UO_243 (O_243,N_14944,N_14921);
nand UO_244 (O_244,N_14877,N_14944);
and UO_245 (O_245,N_14974,N_14926);
xnor UO_246 (O_246,N_14900,N_14981);
xor UO_247 (O_247,N_14964,N_14914);
nor UO_248 (O_248,N_14911,N_14973);
nor UO_249 (O_249,N_14875,N_14988);
nor UO_250 (O_250,N_14918,N_14942);
xor UO_251 (O_251,N_14918,N_14904);
nor UO_252 (O_252,N_14902,N_14941);
or UO_253 (O_253,N_14943,N_14956);
and UO_254 (O_254,N_14902,N_14879);
nand UO_255 (O_255,N_14923,N_14973);
and UO_256 (O_256,N_14974,N_14988);
and UO_257 (O_257,N_14907,N_14903);
and UO_258 (O_258,N_14997,N_14947);
nand UO_259 (O_259,N_14939,N_14959);
nor UO_260 (O_260,N_14890,N_14930);
xor UO_261 (O_261,N_14885,N_14907);
nor UO_262 (O_262,N_14958,N_14969);
xnor UO_263 (O_263,N_14881,N_14876);
nor UO_264 (O_264,N_14926,N_14920);
nand UO_265 (O_265,N_14942,N_14945);
and UO_266 (O_266,N_14975,N_14879);
and UO_267 (O_267,N_14898,N_14996);
and UO_268 (O_268,N_14883,N_14932);
nand UO_269 (O_269,N_14965,N_14913);
or UO_270 (O_270,N_14881,N_14920);
xnor UO_271 (O_271,N_14976,N_14975);
and UO_272 (O_272,N_14884,N_14958);
nor UO_273 (O_273,N_14889,N_14997);
nand UO_274 (O_274,N_14993,N_14963);
and UO_275 (O_275,N_14999,N_14978);
or UO_276 (O_276,N_14892,N_14902);
or UO_277 (O_277,N_14977,N_14951);
nand UO_278 (O_278,N_14893,N_14983);
or UO_279 (O_279,N_14965,N_14912);
xnor UO_280 (O_280,N_14964,N_14903);
nor UO_281 (O_281,N_14953,N_14882);
nor UO_282 (O_282,N_14884,N_14977);
and UO_283 (O_283,N_14969,N_14973);
nand UO_284 (O_284,N_14910,N_14985);
or UO_285 (O_285,N_14975,N_14986);
or UO_286 (O_286,N_14919,N_14891);
nand UO_287 (O_287,N_14997,N_14930);
and UO_288 (O_288,N_14970,N_14984);
xnor UO_289 (O_289,N_14919,N_14895);
and UO_290 (O_290,N_14985,N_14947);
or UO_291 (O_291,N_14929,N_14901);
and UO_292 (O_292,N_14883,N_14927);
xor UO_293 (O_293,N_14980,N_14975);
nand UO_294 (O_294,N_14969,N_14894);
and UO_295 (O_295,N_14933,N_14886);
and UO_296 (O_296,N_14958,N_14989);
nor UO_297 (O_297,N_14917,N_14894);
xnor UO_298 (O_298,N_14993,N_14989);
or UO_299 (O_299,N_14911,N_14916);
xor UO_300 (O_300,N_14882,N_14889);
nand UO_301 (O_301,N_14888,N_14975);
nor UO_302 (O_302,N_14878,N_14980);
nor UO_303 (O_303,N_14920,N_14931);
nor UO_304 (O_304,N_14952,N_14980);
xnor UO_305 (O_305,N_14964,N_14882);
and UO_306 (O_306,N_14882,N_14946);
and UO_307 (O_307,N_14906,N_14944);
xor UO_308 (O_308,N_14978,N_14927);
and UO_309 (O_309,N_14960,N_14949);
xnor UO_310 (O_310,N_14897,N_14903);
nor UO_311 (O_311,N_14956,N_14951);
xor UO_312 (O_312,N_14880,N_14971);
xor UO_313 (O_313,N_14982,N_14959);
or UO_314 (O_314,N_14958,N_14887);
nor UO_315 (O_315,N_14927,N_14987);
xor UO_316 (O_316,N_14958,N_14988);
xnor UO_317 (O_317,N_14919,N_14972);
nor UO_318 (O_318,N_14996,N_14958);
nor UO_319 (O_319,N_14925,N_14988);
xor UO_320 (O_320,N_14888,N_14903);
xnor UO_321 (O_321,N_14918,N_14926);
xor UO_322 (O_322,N_14904,N_14993);
and UO_323 (O_323,N_14968,N_14969);
or UO_324 (O_324,N_14962,N_14876);
nand UO_325 (O_325,N_14881,N_14895);
nand UO_326 (O_326,N_14875,N_14903);
or UO_327 (O_327,N_14973,N_14993);
nor UO_328 (O_328,N_14974,N_14922);
xor UO_329 (O_329,N_14957,N_14907);
nor UO_330 (O_330,N_14953,N_14955);
and UO_331 (O_331,N_14961,N_14901);
and UO_332 (O_332,N_14993,N_14977);
and UO_333 (O_333,N_14939,N_14978);
xor UO_334 (O_334,N_14988,N_14882);
or UO_335 (O_335,N_14944,N_14875);
and UO_336 (O_336,N_14990,N_14984);
nand UO_337 (O_337,N_14921,N_14985);
xnor UO_338 (O_338,N_14997,N_14984);
xor UO_339 (O_339,N_14889,N_14887);
or UO_340 (O_340,N_14997,N_14956);
nor UO_341 (O_341,N_14896,N_14984);
and UO_342 (O_342,N_14908,N_14939);
nand UO_343 (O_343,N_14952,N_14907);
and UO_344 (O_344,N_14917,N_14915);
nand UO_345 (O_345,N_14991,N_14953);
nor UO_346 (O_346,N_14922,N_14956);
or UO_347 (O_347,N_14992,N_14905);
nor UO_348 (O_348,N_14942,N_14903);
nor UO_349 (O_349,N_14962,N_14947);
nand UO_350 (O_350,N_14907,N_14981);
xor UO_351 (O_351,N_14994,N_14993);
and UO_352 (O_352,N_14885,N_14934);
xnor UO_353 (O_353,N_14884,N_14902);
or UO_354 (O_354,N_14944,N_14925);
or UO_355 (O_355,N_14908,N_14976);
nand UO_356 (O_356,N_14905,N_14946);
nor UO_357 (O_357,N_14994,N_14895);
nor UO_358 (O_358,N_14971,N_14933);
xnor UO_359 (O_359,N_14933,N_14901);
nand UO_360 (O_360,N_14941,N_14917);
and UO_361 (O_361,N_14951,N_14884);
or UO_362 (O_362,N_14905,N_14996);
nor UO_363 (O_363,N_14949,N_14941);
nor UO_364 (O_364,N_14950,N_14987);
nand UO_365 (O_365,N_14921,N_14890);
and UO_366 (O_366,N_14960,N_14992);
or UO_367 (O_367,N_14985,N_14997);
nand UO_368 (O_368,N_14912,N_14982);
and UO_369 (O_369,N_14971,N_14881);
xor UO_370 (O_370,N_14997,N_14893);
and UO_371 (O_371,N_14958,N_14985);
nor UO_372 (O_372,N_14920,N_14994);
nor UO_373 (O_373,N_14944,N_14968);
xnor UO_374 (O_374,N_14974,N_14956);
xnor UO_375 (O_375,N_14933,N_14940);
nor UO_376 (O_376,N_14929,N_14883);
nand UO_377 (O_377,N_14948,N_14960);
nor UO_378 (O_378,N_14899,N_14974);
nor UO_379 (O_379,N_14879,N_14976);
nand UO_380 (O_380,N_14925,N_14882);
nor UO_381 (O_381,N_14960,N_14954);
or UO_382 (O_382,N_14919,N_14914);
and UO_383 (O_383,N_14886,N_14900);
or UO_384 (O_384,N_14946,N_14969);
nand UO_385 (O_385,N_14951,N_14998);
xor UO_386 (O_386,N_14907,N_14995);
xnor UO_387 (O_387,N_14895,N_14986);
nand UO_388 (O_388,N_14998,N_14886);
xor UO_389 (O_389,N_14997,N_14978);
nand UO_390 (O_390,N_14950,N_14914);
and UO_391 (O_391,N_14895,N_14950);
and UO_392 (O_392,N_14932,N_14940);
and UO_393 (O_393,N_14951,N_14976);
and UO_394 (O_394,N_14984,N_14941);
xnor UO_395 (O_395,N_14948,N_14905);
or UO_396 (O_396,N_14911,N_14907);
xnor UO_397 (O_397,N_14943,N_14974);
or UO_398 (O_398,N_14950,N_14916);
nand UO_399 (O_399,N_14887,N_14899);
xnor UO_400 (O_400,N_14882,N_14993);
nand UO_401 (O_401,N_14904,N_14978);
or UO_402 (O_402,N_14952,N_14979);
nand UO_403 (O_403,N_14878,N_14961);
and UO_404 (O_404,N_14909,N_14971);
and UO_405 (O_405,N_14987,N_14912);
xor UO_406 (O_406,N_14950,N_14938);
nand UO_407 (O_407,N_14918,N_14958);
nor UO_408 (O_408,N_14951,N_14927);
nand UO_409 (O_409,N_14891,N_14884);
nand UO_410 (O_410,N_14994,N_14880);
and UO_411 (O_411,N_14934,N_14916);
and UO_412 (O_412,N_14950,N_14992);
nor UO_413 (O_413,N_14961,N_14920);
nor UO_414 (O_414,N_14907,N_14960);
or UO_415 (O_415,N_14910,N_14906);
and UO_416 (O_416,N_14997,N_14901);
nand UO_417 (O_417,N_14991,N_14904);
nand UO_418 (O_418,N_14980,N_14897);
or UO_419 (O_419,N_14988,N_14963);
nand UO_420 (O_420,N_14951,N_14918);
nor UO_421 (O_421,N_14894,N_14935);
nor UO_422 (O_422,N_14959,N_14990);
and UO_423 (O_423,N_14879,N_14955);
or UO_424 (O_424,N_14915,N_14986);
nor UO_425 (O_425,N_14951,N_14996);
nand UO_426 (O_426,N_14988,N_14896);
nor UO_427 (O_427,N_14962,N_14928);
nand UO_428 (O_428,N_14925,N_14970);
and UO_429 (O_429,N_14983,N_14930);
xnor UO_430 (O_430,N_14908,N_14961);
nor UO_431 (O_431,N_14935,N_14914);
and UO_432 (O_432,N_14897,N_14984);
or UO_433 (O_433,N_14964,N_14941);
nand UO_434 (O_434,N_14885,N_14943);
or UO_435 (O_435,N_14916,N_14956);
and UO_436 (O_436,N_14877,N_14898);
nand UO_437 (O_437,N_14961,N_14939);
or UO_438 (O_438,N_14960,N_14917);
nor UO_439 (O_439,N_14924,N_14975);
nand UO_440 (O_440,N_14975,N_14984);
xnor UO_441 (O_441,N_14875,N_14904);
nor UO_442 (O_442,N_14884,N_14967);
nor UO_443 (O_443,N_14946,N_14890);
or UO_444 (O_444,N_14965,N_14894);
xnor UO_445 (O_445,N_14990,N_14918);
or UO_446 (O_446,N_14942,N_14994);
nor UO_447 (O_447,N_14952,N_14931);
and UO_448 (O_448,N_14901,N_14903);
and UO_449 (O_449,N_14888,N_14938);
or UO_450 (O_450,N_14926,N_14907);
and UO_451 (O_451,N_14916,N_14949);
xor UO_452 (O_452,N_14937,N_14941);
nand UO_453 (O_453,N_14912,N_14924);
or UO_454 (O_454,N_14941,N_14919);
or UO_455 (O_455,N_14885,N_14894);
xnor UO_456 (O_456,N_14921,N_14948);
xor UO_457 (O_457,N_14995,N_14935);
and UO_458 (O_458,N_14988,N_14876);
nand UO_459 (O_459,N_14885,N_14927);
and UO_460 (O_460,N_14948,N_14878);
nor UO_461 (O_461,N_14943,N_14904);
nand UO_462 (O_462,N_14957,N_14968);
xor UO_463 (O_463,N_14899,N_14969);
or UO_464 (O_464,N_14933,N_14968);
and UO_465 (O_465,N_14962,N_14989);
nor UO_466 (O_466,N_14928,N_14931);
xor UO_467 (O_467,N_14933,N_14932);
and UO_468 (O_468,N_14919,N_14910);
nor UO_469 (O_469,N_14899,N_14884);
or UO_470 (O_470,N_14879,N_14917);
and UO_471 (O_471,N_14999,N_14942);
nand UO_472 (O_472,N_14923,N_14903);
or UO_473 (O_473,N_14945,N_14877);
nor UO_474 (O_474,N_14894,N_14994);
nor UO_475 (O_475,N_14958,N_14977);
and UO_476 (O_476,N_14956,N_14936);
nor UO_477 (O_477,N_14959,N_14914);
xor UO_478 (O_478,N_14985,N_14979);
nor UO_479 (O_479,N_14970,N_14948);
xor UO_480 (O_480,N_14879,N_14901);
or UO_481 (O_481,N_14914,N_14990);
or UO_482 (O_482,N_14899,N_14973);
and UO_483 (O_483,N_14970,N_14892);
nand UO_484 (O_484,N_14916,N_14906);
and UO_485 (O_485,N_14963,N_14948);
or UO_486 (O_486,N_14914,N_14937);
nand UO_487 (O_487,N_14990,N_14968);
nor UO_488 (O_488,N_14895,N_14898);
and UO_489 (O_489,N_14890,N_14973);
xor UO_490 (O_490,N_14884,N_14973);
or UO_491 (O_491,N_14922,N_14957);
xor UO_492 (O_492,N_14974,N_14980);
nor UO_493 (O_493,N_14981,N_14932);
nor UO_494 (O_494,N_14980,N_14934);
or UO_495 (O_495,N_14931,N_14980);
xor UO_496 (O_496,N_14892,N_14931);
xnor UO_497 (O_497,N_14914,N_14917);
and UO_498 (O_498,N_14958,N_14910);
nand UO_499 (O_499,N_14999,N_14894);
nand UO_500 (O_500,N_14968,N_14895);
nor UO_501 (O_501,N_14940,N_14962);
or UO_502 (O_502,N_14926,N_14949);
nand UO_503 (O_503,N_14997,N_14902);
and UO_504 (O_504,N_14915,N_14990);
nor UO_505 (O_505,N_14993,N_14975);
xnor UO_506 (O_506,N_14998,N_14995);
and UO_507 (O_507,N_14915,N_14905);
xor UO_508 (O_508,N_14987,N_14949);
nand UO_509 (O_509,N_14913,N_14882);
and UO_510 (O_510,N_14926,N_14910);
nor UO_511 (O_511,N_14954,N_14885);
nand UO_512 (O_512,N_14918,N_14936);
or UO_513 (O_513,N_14973,N_14913);
or UO_514 (O_514,N_14949,N_14927);
nand UO_515 (O_515,N_14926,N_14883);
and UO_516 (O_516,N_14973,N_14960);
xor UO_517 (O_517,N_14994,N_14948);
xor UO_518 (O_518,N_14926,N_14934);
nand UO_519 (O_519,N_14895,N_14960);
and UO_520 (O_520,N_14936,N_14875);
nor UO_521 (O_521,N_14923,N_14883);
nand UO_522 (O_522,N_14970,N_14895);
and UO_523 (O_523,N_14986,N_14875);
nand UO_524 (O_524,N_14999,N_14909);
xor UO_525 (O_525,N_14953,N_14921);
and UO_526 (O_526,N_14997,N_14995);
xor UO_527 (O_527,N_14909,N_14968);
and UO_528 (O_528,N_14961,N_14931);
nor UO_529 (O_529,N_14919,N_14924);
or UO_530 (O_530,N_14989,N_14959);
xnor UO_531 (O_531,N_14877,N_14981);
and UO_532 (O_532,N_14890,N_14947);
and UO_533 (O_533,N_14976,N_14995);
nand UO_534 (O_534,N_14996,N_14931);
and UO_535 (O_535,N_14968,N_14946);
xor UO_536 (O_536,N_14924,N_14949);
or UO_537 (O_537,N_14899,N_14880);
xnor UO_538 (O_538,N_14895,N_14897);
xnor UO_539 (O_539,N_14881,N_14965);
and UO_540 (O_540,N_14991,N_14911);
nor UO_541 (O_541,N_14876,N_14982);
nand UO_542 (O_542,N_14899,N_14926);
or UO_543 (O_543,N_14970,N_14983);
xor UO_544 (O_544,N_14936,N_14883);
or UO_545 (O_545,N_14982,N_14997);
nand UO_546 (O_546,N_14933,N_14909);
nor UO_547 (O_547,N_14915,N_14892);
nand UO_548 (O_548,N_14967,N_14944);
or UO_549 (O_549,N_14958,N_14953);
or UO_550 (O_550,N_14975,N_14897);
or UO_551 (O_551,N_14943,N_14949);
nand UO_552 (O_552,N_14966,N_14944);
nand UO_553 (O_553,N_14947,N_14921);
and UO_554 (O_554,N_14974,N_14912);
nand UO_555 (O_555,N_14964,N_14997);
nor UO_556 (O_556,N_14931,N_14890);
or UO_557 (O_557,N_14928,N_14963);
xor UO_558 (O_558,N_14944,N_14987);
nor UO_559 (O_559,N_14952,N_14989);
nor UO_560 (O_560,N_14935,N_14879);
and UO_561 (O_561,N_14986,N_14877);
or UO_562 (O_562,N_14990,N_14898);
nand UO_563 (O_563,N_14906,N_14904);
and UO_564 (O_564,N_14929,N_14902);
or UO_565 (O_565,N_14876,N_14961);
nand UO_566 (O_566,N_14997,N_14943);
or UO_567 (O_567,N_14931,N_14945);
and UO_568 (O_568,N_14977,N_14896);
nand UO_569 (O_569,N_14919,N_14945);
and UO_570 (O_570,N_14990,N_14936);
nor UO_571 (O_571,N_14988,N_14916);
nand UO_572 (O_572,N_14892,N_14995);
nor UO_573 (O_573,N_14889,N_14968);
or UO_574 (O_574,N_14960,N_14894);
or UO_575 (O_575,N_14982,N_14943);
nand UO_576 (O_576,N_14956,N_14957);
nor UO_577 (O_577,N_14928,N_14989);
nor UO_578 (O_578,N_14998,N_14929);
nor UO_579 (O_579,N_14902,N_14985);
or UO_580 (O_580,N_14897,N_14928);
nand UO_581 (O_581,N_14992,N_14944);
xnor UO_582 (O_582,N_14954,N_14978);
nand UO_583 (O_583,N_14890,N_14903);
or UO_584 (O_584,N_14892,N_14918);
nor UO_585 (O_585,N_14945,N_14930);
nand UO_586 (O_586,N_14915,N_14933);
nor UO_587 (O_587,N_14928,N_14978);
and UO_588 (O_588,N_14959,N_14943);
nand UO_589 (O_589,N_14916,N_14913);
and UO_590 (O_590,N_14925,N_14996);
nand UO_591 (O_591,N_14961,N_14956);
nand UO_592 (O_592,N_14928,N_14955);
and UO_593 (O_593,N_14893,N_14976);
nand UO_594 (O_594,N_14959,N_14919);
nand UO_595 (O_595,N_14878,N_14987);
or UO_596 (O_596,N_14993,N_14902);
xnor UO_597 (O_597,N_14909,N_14891);
xnor UO_598 (O_598,N_14917,N_14947);
nand UO_599 (O_599,N_14981,N_14987);
nand UO_600 (O_600,N_14981,N_14894);
nor UO_601 (O_601,N_14992,N_14974);
or UO_602 (O_602,N_14969,N_14883);
or UO_603 (O_603,N_14997,N_14973);
and UO_604 (O_604,N_14885,N_14898);
nor UO_605 (O_605,N_14986,N_14951);
or UO_606 (O_606,N_14952,N_14879);
nand UO_607 (O_607,N_14983,N_14905);
or UO_608 (O_608,N_14878,N_14986);
xor UO_609 (O_609,N_14916,N_14995);
or UO_610 (O_610,N_14965,N_14961);
or UO_611 (O_611,N_14976,N_14971);
nand UO_612 (O_612,N_14911,N_14924);
nand UO_613 (O_613,N_14912,N_14994);
nand UO_614 (O_614,N_14953,N_14906);
nand UO_615 (O_615,N_14886,N_14959);
or UO_616 (O_616,N_14937,N_14923);
nand UO_617 (O_617,N_14970,N_14932);
xor UO_618 (O_618,N_14880,N_14942);
xor UO_619 (O_619,N_14952,N_14894);
nor UO_620 (O_620,N_14907,N_14961);
nor UO_621 (O_621,N_14941,N_14894);
nor UO_622 (O_622,N_14999,N_14974);
nor UO_623 (O_623,N_14971,N_14884);
nor UO_624 (O_624,N_14925,N_14911);
and UO_625 (O_625,N_14977,N_14953);
and UO_626 (O_626,N_14902,N_14942);
nand UO_627 (O_627,N_14898,N_14902);
or UO_628 (O_628,N_14976,N_14953);
and UO_629 (O_629,N_14993,N_14986);
nand UO_630 (O_630,N_14985,N_14880);
nor UO_631 (O_631,N_14880,N_14979);
nand UO_632 (O_632,N_14979,N_14930);
or UO_633 (O_633,N_14897,N_14962);
or UO_634 (O_634,N_14894,N_14921);
xnor UO_635 (O_635,N_14952,N_14881);
and UO_636 (O_636,N_14887,N_14996);
or UO_637 (O_637,N_14956,N_14940);
and UO_638 (O_638,N_14990,N_14947);
and UO_639 (O_639,N_14978,N_14908);
nor UO_640 (O_640,N_14966,N_14876);
and UO_641 (O_641,N_14896,N_14978);
or UO_642 (O_642,N_14979,N_14992);
or UO_643 (O_643,N_14907,N_14979);
or UO_644 (O_644,N_14955,N_14878);
or UO_645 (O_645,N_14881,N_14891);
and UO_646 (O_646,N_14910,N_14914);
and UO_647 (O_647,N_14891,N_14982);
xnor UO_648 (O_648,N_14976,N_14941);
nor UO_649 (O_649,N_14934,N_14928);
nor UO_650 (O_650,N_14996,N_14993);
xor UO_651 (O_651,N_14982,N_14909);
and UO_652 (O_652,N_14982,N_14888);
nand UO_653 (O_653,N_14935,N_14886);
nand UO_654 (O_654,N_14890,N_14958);
or UO_655 (O_655,N_14932,N_14916);
xor UO_656 (O_656,N_14941,N_14990);
or UO_657 (O_657,N_14952,N_14986);
xor UO_658 (O_658,N_14934,N_14987);
and UO_659 (O_659,N_14937,N_14961);
nand UO_660 (O_660,N_14892,N_14891);
or UO_661 (O_661,N_14920,N_14899);
nand UO_662 (O_662,N_14977,N_14901);
nand UO_663 (O_663,N_14918,N_14995);
and UO_664 (O_664,N_14948,N_14947);
xor UO_665 (O_665,N_14949,N_14975);
xor UO_666 (O_666,N_14902,N_14974);
and UO_667 (O_667,N_14942,N_14914);
xor UO_668 (O_668,N_14974,N_14958);
or UO_669 (O_669,N_14980,N_14971);
or UO_670 (O_670,N_14955,N_14989);
nor UO_671 (O_671,N_14931,N_14957);
xnor UO_672 (O_672,N_14980,N_14948);
nand UO_673 (O_673,N_14921,N_14916);
and UO_674 (O_674,N_14967,N_14984);
nand UO_675 (O_675,N_14882,N_14928);
xnor UO_676 (O_676,N_14900,N_14914);
and UO_677 (O_677,N_14955,N_14943);
xor UO_678 (O_678,N_14875,N_14911);
nor UO_679 (O_679,N_14954,N_14998);
xor UO_680 (O_680,N_14928,N_14945);
xor UO_681 (O_681,N_14962,N_14949);
nor UO_682 (O_682,N_14909,N_14922);
nand UO_683 (O_683,N_14896,N_14897);
or UO_684 (O_684,N_14915,N_14987);
or UO_685 (O_685,N_14901,N_14968);
nand UO_686 (O_686,N_14933,N_14911);
nand UO_687 (O_687,N_14944,N_14898);
nor UO_688 (O_688,N_14915,N_14887);
or UO_689 (O_689,N_14974,N_14935);
nand UO_690 (O_690,N_14930,N_14987);
xnor UO_691 (O_691,N_14957,N_14974);
nor UO_692 (O_692,N_14926,N_14992);
and UO_693 (O_693,N_14914,N_14930);
and UO_694 (O_694,N_14936,N_14985);
or UO_695 (O_695,N_14891,N_14999);
and UO_696 (O_696,N_14954,N_14900);
or UO_697 (O_697,N_14946,N_14932);
nor UO_698 (O_698,N_14988,N_14907);
nand UO_699 (O_699,N_14932,N_14895);
xnor UO_700 (O_700,N_14987,N_14947);
and UO_701 (O_701,N_14929,N_14921);
and UO_702 (O_702,N_14980,N_14882);
xor UO_703 (O_703,N_14959,N_14965);
or UO_704 (O_704,N_14926,N_14957);
or UO_705 (O_705,N_14915,N_14989);
nand UO_706 (O_706,N_14920,N_14945);
or UO_707 (O_707,N_14982,N_14906);
and UO_708 (O_708,N_14893,N_14929);
nand UO_709 (O_709,N_14959,N_14988);
or UO_710 (O_710,N_14931,N_14940);
nand UO_711 (O_711,N_14937,N_14893);
and UO_712 (O_712,N_14948,N_14971);
or UO_713 (O_713,N_14999,N_14915);
nand UO_714 (O_714,N_14890,N_14892);
nor UO_715 (O_715,N_14903,N_14955);
nor UO_716 (O_716,N_14973,N_14999);
nand UO_717 (O_717,N_14999,N_14878);
and UO_718 (O_718,N_14919,N_14923);
or UO_719 (O_719,N_14925,N_14904);
or UO_720 (O_720,N_14909,N_14989);
and UO_721 (O_721,N_14878,N_14954);
or UO_722 (O_722,N_14908,N_14947);
and UO_723 (O_723,N_14940,N_14968);
xnor UO_724 (O_724,N_14979,N_14980);
nand UO_725 (O_725,N_14995,N_14915);
or UO_726 (O_726,N_14951,N_14952);
nand UO_727 (O_727,N_14940,N_14948);
and UO_728 (O_728,N_14968,N_14985);
or UO_729 (O_729,N_14954,N_14988);
or UO_730 (O_730,N_14994,N_14875);
xor UO_731 (O_731,N_14926,N_14928);
and UO_732 (O_732,N_14920,N_14975);
or UO_733 (O_733,N_14925,N_14921);
or UO_734 (O_734,N_14954,N_14964);
or UO_735 (O_735,N_14990,N_14891);
or UO_736 (O_736,N_14913,N_14952);
or UO_737 (O_737,N_14928,N_14949);
and UO_738 (O_738,N_14925,N_14936);
and UO_739 (O_739,N_14910,N_14891);
nand UO_740 (O_740,N_14966,N_14911);
xnor UO_741 (O_741,N_14970,N_14889);
xor UO_742 (O_742,N_14929,N_14945);
or UO_743 (O_743,N_14965,N_14954);
or UO_744 (O_744,N_14984,N_14937);
or UO_745 (O_745,N_14994,N_14914);
nand UO_746 (O_746,N_14940,N_14937);
or UO_747 (O_747,N_14902,N_14944);
or UO_748 (O_748,N_14983,N_14949);
nand UO_749 (O_749,N_14981,N_14994);
and UO_750 (O_750,N_14966,N_14912);
xor UO_751 (O_751,N_14925,N_14913);
xor UO_752 (O_752,N_14980,N_14933);
nor UO_753 (O_753,N_14900,N_14988);
xor UO_754 (O_754,N_14875,N_14910);
nor UO_755 (O_755,N_14982,N_14928);
xor UO_756 (O_756,N_14959,N_14951);
or UO_757 (O_757,N_14982,N_14895);
and UO_758 (O_758,N_14922,N_14893);
nor UO_759 (O_759,N_14900,N_14941);
or UO_760 (O_760,N_14965,N_14942);
xnor UO_761 (O_761,N_14921,N_14961);
or UO_762 (O_762,N_14950,N_14979);
and UO_763 (O_763,N_14889,N_14958);
xor UO_764 (O_764,N_14991,N_14881);
xnor UO_765 (O_765,N_14878,N_14912);
xnor UO_766 (O_766,N_14921,N_14991);
xor UO_767 (O_767,N_14973,N_14928);
nand UO_768 (O_768,N_14993,N_14925);
or UO_769 (O_769,N_14928,N_14879);
nor UO_770 (O_770,N_14948,N_14987);
nor UO_771 (O_771,N_14974,N_14933);
or UO_772 (O_772,N_14941,N_14920);
or UO_773 (O_773,N_14981,N_14895);
and UO_774 (O_774,N_14956,N_14969);
and UO_775 (O_775,N_14924,N_14959);
nand UO_776 (O_776,N_14954,N_14995);
nand UO_777 (O_777,N_14907,N_14884);
or UO_778 (O_778,N_14886,N_14907);
nor UO_779 (O_779,N_14900,N_14925);
and UO_780 (O_780,N_14912,N_14915);
xor UO_781 (O_781,N_14901,N_14991);
nor UO_782 (O_782,N_14884,N_14911);
or UO_783 (O_783,N_14961,N_14887);
xnor UO_784 (O_784,N_14974,N_14915);
xor UO_785 (O_785,N_14988,N_14965);
and UO_786 (O_786,N_14880,N_14945);
or UO_787 (O_787,N_14971,N_14890);
nor UO_788 (O_788,N_14932,N_14962);
xnor UO_789 (O_789,N_14896,N_14961);
xor UO_790 (O_790,N_14935,N_14926);
xnor UO_791 (O_791,N_14968,N_14893);
or UO_792 (O_792,N_14965,N_14935);
or UO_793 (O_793,N_14895,N_14966);
or UO_794 (O_794,N_14937,N_14906);
xnor UO_795 (O_795,N_14929,N_14891);
xnor UO_796 (O_796,N_14929,N_14981);
and UO_797 (O_797,N_14889,N_14930);
xnor UO_798 (O_798,N_14875,N_14974);
and UO_799 (O_799,N_14946,N_14943);
nor UO_800 (O_800,N_14961,N_14950);
nand UO_801 (O_801,N_14943,N_14919);
nand UO_802 (O_802,N_14928,N_14985);
nor UO_803 (O_803,N_14971,N_14968);
nor UO_804 (O_804,N_14875,N_14915);
nor UO_805 (O_805,N_14892,N_14975);
xnor UO_806 (O_806,N_14982,N_14949);
or UO_807 (O_807,N_14961,N_14897);
or UO_808 (O_808,N_14949,N_14930);
nand UO_809 (O_809,N_14965,N_14885);
nand UO_810 (O_810,N_14944,N_14905);
xor UO_811 (O_811,N_14982,N_14993);
xor UO_812 (O_812,N_14956,N_14907);
nand UO_813 (O_813,N_14978,N_14918);
and UO_814 (O_814,N_14963,N_14892);
or UO_815 (O_815,N_14965,N_14904);
or UO_816 (O_816,N_14925,N_14933);
nor UO_817 (O_817,N_14916,N_14912);
and UO_818 (O_818,N_14924,N_14908);
or UO_819 (O_819,N_14905,N_14906);
nor UO_820 (O_820,N_14892,N_14981);
and UO_821 (O_821,N_14918,N_14998);
or UO_822 (O_822,N_14882,N_14982);
and UO_823 (O_823,N_14980,N_14907);
xor UO_824 (O_824,N_14990,N_14884);
or UO_825 (O_825,N_14970,N_14942);
xnor UO_826 (O_826,N_14902,N_14916);
nand UO_827 (O_827,N_14994,N_14934);
and UO_828 (O_828,N_14911,N_14921);
or UO_829 (O_829,N_14890,N_14966);
or UO_830 (O_830,N_14996,N_14980);
or UO_831 (O_831,N_14976,N_14884);
and UO_832 (O_832,N_14923,N_14892);
and UO_833 (O_833,N_14903,N_14983);
nor UO_834 (O_834,N_14975,N_14884);
xnor UO_835 (O_835,N_14902,N_14908);
xor UO_836 (O_836,N_14936,N_14994);
nand UO_837 (O_837,N_14981,N_14992);
or UO_838 (O_838,N_14880,N_14913);
xor UO_839 (O_839,N_14921,N_14969);
xor UO_840 (O_840,N_14903,N_14931);
xnor UO_841 (O_841,N_14987,N_14908);
and UO_842 (O_842,N_14933,N_14907);
xnor UO_843 (O_843,N_14907,N_14935);
nor UO_844 (O_844,N_14893,N_14883);
and UO_845 (O_845,N_14976,N_14986);
xnor UO_846 (O_846,N_14959,N_14933);
and UO_847 (O_847,N_14953,N_14897);
nor UO_848 (O_848,N_14997,N_14961);
or UO_849 (O_849,N_14887,N_14935);
or UO_850 (O_850,N_14942,N_14940);
xnor UO_851 (O_851,N_14914,N_14970);
nand UO_852 (O_852,N_14915,N_14919);
and UO_853 (O_853,N_14993,N_14909);
or UO_854 (O_854,N_14895,N_14889);
and UO_855 (O_855,N_14998,N_14904);
nor UO_856 (O_856,N_14890,N_14882);
nor UO_857 (O_857,N_14890,N_14944);
xnor UO_858 (O_858,N_14901,N_14878);
xor UO_859 (O_859,N_14926,N_14892);
or UO_860 (O_860,N_14971,N_14907);
nor UO_861 (O_861,N_14946,N_14972);
or UO_862 (O_862,N_14911,N_14975);
xnor UO_863 (O_863,N_14902,N_14948);
and UO_864 (O_864,N_14996,N_14919);
nand UO_865 (O_865,N_14922,N_14945);
and UO_866 (O_866,N_14940,N_14952);
xnor UO_867 (O_867,N_14885,N_14964);
and UO_868 (O_868,N_14958,N_14999);
nand UO_869 (O_869,N_14926,N_14970);
and UO_870 (O_870,N_14954,N_14972);
or UO_871 (O_871,N_14939,N_14950);
or UO_872 (O_872,N_14935,N_14884);
nand UO_873 (O_873,N_14934,N_14939);
xnor UO_874 (O_874,N_14899,N_14943);
xor UO_875 (O_875,N_14954,N_14943);
or UO_876 (O_876,N_14906,N_14896);
or UO_877 (O_877,N_14889,N_14880);
xnor UO_878 (O_878,N_14992,N_14923);
xnor UO_879 (O_879,N_14922,N_14993);
xor UO_880 (O_880,N_14956,N_14899);
or UO_881 (O_881,N_14879,N_14970);
and UO_882 (O_882,N_14957,N_14997);
or UO_883 (O_883,N_14928,N_14942);
or UO_884 (O_884,N_14876,N_14999);
and UO_885 (O_885,N_14886,N_14875);
nand UO_886 (O_886,N_14938,N_14909);
and UO_887 (O_887,N_14996,N_14962);
nor UO_888 (O_888,N_14935,N_14936);
or UO_889 (O_889,N_14883,N_14941);
and UO_890 (O_890,N_14941,N_14912);
and UO_891 (O_891,N_14968,N_14924);
nor UO_892 (O_892,N_14973,N_14982);
nand UO_893 (O_893,N_14909,N_14978);
and UO_894 (O_894,N_14998,N_14983);
or UO_895 (O_895,N_14967,N_14983);
xnor UO_896 (O_896,N_14966,N_14987);
nand UO_897 (O_897,N_14927,N_14989);
nand UO_898 (O_898,N_14982,N_14878);
nand UO_899 (O_899,N_14914,N_14995);
xnor UO_900 (O_900,N_14876,N_14965);
or UO_901 (O_901,N_14884,N_14926);
nand UO_902 (O_902,N_14878,N_14910);
nor UO_903 (O_903,N_14970,N_14964);
or UO_904 (O_904,N_14898,N_14932);
nand UO_905 (O_905,N_14995,N_14991);
and UO_906 (O_906,N_14939,N_14974);
nor UO_907 (O_907,N_14968,N_14878);
and UO_908 (O_908,N_14925,N_14998);
nand UO_909 (O_909,N_14916,N_14964);
nand UO_910 (O_910,N_14963,N_14886);
xnor UO_911 (O_911,N_14936,N_14924);
xor UO_912 (O_912,N_14881,N_14879);
or UO_913 (O_913,N_14983,N_14990);
xnor UO_914 (O_914,N_14961,N_14954);
nand UO_915 (O_915,N_14889,N_14932);
nand UO_916 (O_916,N_14927,N_14984);
xor UO_917 (O_917,N_14905,N_14982);
and UO_918 (O_918,N_14951,N_14983);
xnor UO_919 (O_919,N_14921,N_14938);
xnor UO_920 (O_920,N_14933,N_14949);
nand UO_921 (O_921,N_14894,N_14925);
and UO_922 (O_922,N_14978,N_14923);
nand UO_923 (O_923,N_14983,N_14925);
nor UO_924 (O_924,N_14946,N_14924);
nor UO_925 (O_925,N_14909,N_14878);
nor UO_926 (O_926,N_14982,N_14987);
or UO_927 (O_927,N_14951,N_14989);
and UO_928 (O_928,N_14880,N_14995);
and UO_929 (O_929,N_14888,N_14934);
nand UO_930 (O_930,N_14875,N_14971);
nand UO_931 (O_931,N_14901,N_14881);
nand UO_932 (O_932,N_14938,N_14919);
or UO_933 (O_933,N_14943,N_14928);
nor UO_934 (O_934,N_14919,N_14920);
or UO_935 (O_935,N_14917,N_14987);
nor UO_936 (O_936,N_14889,N_14918);
nand UO_937 (O_937,N_14877,N_14884);
and UO_938 (O_938,N_14931,N_14895);
xor UO_939 (O_939,N_14937,N_14898);
or UO_940 (O_940,N_14906,N_14875);
and UO_941 (O_941,N_14931,N_14997);
and UO_942 (O_942,N_14931,N_14924);
or UO_943 (O_943,N_14985,N_14892);
xnor UO_944 (O_944,N_14968,N_14879);
and UO_945 (O_945,N_14998,N_14909);
or UO_946 (O_946,N_14961,N_14875);
or UO_947 (O_947,N_14897,N_14933);
xor UO_948 (O_948,N_14985,N_14914);
nand UO_949 (O_949,N_14927,N_14913);
and UO_950 (O_950,N_14959,N_14903);
nand UO_951 (O_951,N_14906,N_14993);
and UO_952 (O_952,N_14903,N_14949);
xnor UO_953 (O_953,N_14956,N_14975);
and UO_954 (O_954,N_14900,N_14984);
and UO_955 (O_955,N_14997,N_14921);
and UO_956 (O_956,N_14955,N_14946);
xor UO_957 (O_957,N_14942,N_14905);
and UO_958 (O_958,N_14964,N_14883);
or UO_959 (O_959,N_14885,N_14930);
or UO_960 (O_960,N_14959,N_14887);
xor UO_961 (O_961,N_14957,N_14880);
and UO_962 (O_962,N_14963,N_14957);
or UO_963 (O_963,N_14973,N_14950);
or UO_964 (O_964,N_14948,N_14986);
and UO_965 (O_965,N_14907,N_14929);
nor UO_966 (O_966,N_14921,N_14902);
xor UO_967 (O_967,N_14929,N_14991);
xnor UO_968 (O_968,N_14958,N_14941);
and UO_969 (O_969,N_14902,N_14910);
and UO_970 (O_970,N_14985,N_14957);
or UO_971 (O_971,N_14992,N_14888);
xor UO_972 (O_972,N_14957,N_14906);
nor UO_973 (O_973,N_14901,N_14979);
nand UO_974 (O_974,N_14990,N_14893);
and UO_975 (O_975,N_14931,N_14933);
and UO_976 (O_976,N_14956,N_14901);
xor UO_977 (O_977,N_14969,N_14947);
nor UO_978 (O_978,N_14921,N_14912);
xor UO_979 (O_979,N_14979,N_14963);
or UO_980 (O_980,N_14919,N_14930);
nor UO_981 (O_981,N_14921,N_14990);
or UO_982 (O_982,N_14920,N_14990);
nand UO_983 (O_983,N_14963,N_14997);
and UO_984 (O_984,N_14998,N_14887);
and UO_985 (O_985,N_14993,N_14930);
xor UO_986 (O_986,N_14980,N_14967);
nor UO_987 (O_987,N_14954,N_14880);
xor UO_988 (O_988,N_14960,N_14887);
or UO_989 (O_989,N_14976,N_14952);
or UO_990 (O_990,N_14899,N_14979);
xnor UO_991 (O_991,N_14967,N_14941);
nor UO_992 (O_992,N_14884,N_14930);
xor UO_993 (O_993,N_14955,N_14980);
or UO_994 (O_994,N_14993,N_14916);
or UO_995 (O_995,N_14990,N_14953);
nor UO_996 (O_996,N_14967,N_14927);
nor UO_997 (O_997,N_14949,N_14890);
nand UO_998 (O_998,N_14988,N_14921);
xor UO_999 (O_999,N_14945,N_14933);
nand UO_1000 (O_1000,N_14933,N_14965);
nand UO_1001 (O_1001,N_14936,N_14879);
nand UO_1002 (O_1002,N_14899,N_14945);
and UO_1003 (O_1003,N_14977,N_14952);
nand UO_1004 (O_1004,N_14933,N_14876);
nor UO_1005 (O_1005,N_14959,N_14958);
xor UO_1006 (O_1006,N_14943,N_14971);
xor UO_1007 (O_1007,N_14962,N_14980);
nor UO_1008 (O_1008,N_14876,N_14888);
nand UO_1009 (O_1009,N_14978,N_14940);
or UO_1010 (O_1010,N_14982,N_14985);
or UO_1011 (O_1011,N_14882,N_14900);
or UO_1012 (O_1012,N_14878,N_14897);
and UO_1013 (O_1013,N_14978,N_14960);
xnor UO_1014 (O_1014,N_14938,N_14990);
nand UO_1015 (O_1015,N_14911,N_14950);
nor UO_1016 (O_1016,N_14929,N_14900);
xnor UO_1017 (O_1017,N_14901,N_14877);
nand UO_1018 (O_1018,N_14940,N_14923);
and UO_1019 (O_1019,N_14947,N_14943);
and UO_1020 (O_1020,N_14927,N_14904);
nand UO_1021 (O_1021,N_14920,N_14938);
or UO_1022 (O_1022,N_14932,N_14976);
xor UO_1023 (O_1023,N_14877,N_14946);
nand UO_1024 (O_1024,N_14976,N_14911);
or UO_1025 (O_1025,N_14987,N_14968);
and UO_1026 (O_1026,N_14958,N_14926);
xor UO_1027 (O_1027,N_14943,N_14908);
and UO_1028 (O_1028,N_14939,N_14935);
nor UO_1029 (O_1029,N_14986,N_14984);
or UO_1030 (O_1030,N_14946,N_14913);
and UO_1031 (O_1031,N_14939,N_14878);
nand UO_1032 (O_1032,N_14937,N_14911);
nor UO_1033 (O_1033,N_14893,N_14894);
or UO_1034 (O_1034,N_14991,N_14950);
or UO_1035 (O_1035,N_14962,N_14974);
nor UO_1036 (O_1036,N_14895,N_14890);
nor UO_1037 (O_1037,N_14981,N_14906);
nand UO_1038 (O_1038,N_14910,N_14983);
or UO_1039 (O_1039,N_14934,N_14992);
nand UO_1040 (O_1040,N_14966,N_14883);
nand UO_1041 (O_1041,N_14896,N_14902);
xor UO_1042 (O_1042,N_14893,N_14995);
and UO_1043 (O_1043,N_14938,N_14989);
and UO_1044 (O_1044,N_14955,N_14930);
xnor UO_1045 (O_1045,N_14937,N_14909);
and UO_1046 (O_1046,N_14940,N_14950);
xnor UO_1047 (O_1047,N_14916,N_14960);
and UO_1048 (O_1048,N_14993,N_14913);
nand UO_1049 (O_1049,N_14935,N_14896);
nand UO_1050 (O_1050,N_14905,N_14920);
nand UO_1051 (O_1051,N_14895,N_14922);
nor UO_1052 (O_1052,N_14987,N_14879);
nand UO_1053 (O_1053,N_14935,N_14910);
xnor UO_1054 (O_1054,N_14960,N_14901);
nand UO_1055 (O_1055,N_14949,N_14875);
nor UO_1056 (O_1056,N_14989,N_14935);
nand UO_1057 (O_1057,N_14883,N_14919);
or UO_1058 (O_1058,N_14920,N_14933);
nor UO_1059 (O_1059,N_14891,N_14902);
nor UO_1060 (O_1060,N_14904,N_14939);
xnor UO_1061 (O_1061,N_14902,N_14979);
xnor UO_1062 (O_1062,N_14883,N_14881);
xnor UO_1063 (O_1063,N_14907,N_14888);
xor UO_1064 (O_1064,N_14921,N_14960);
xor UO_1065 (O_1065,N_14927,N_14953);
and UO_1066 (O_1066,N_14900,N_14986);
and UO_1067 (O_1067,N_14955,N_14987);
and UO_1068 (O_1068,N_14988,N_14919);
nand UO_1069 (O_1069,N_14928,N_14912);
and UO_1070 (O_1070,N_14983,N_14915);
and UO_1071 (O_1071,N_14884,N_14896);
xor UO_1072 (O_1072,N_14999,N_14955);
nor UO_1073 (O_1073,N_14940,N_14972);
and UO_1074 (O_1074,N_14934,N_14924);
and UO_1075 (O_1075,N_14975,N_14921);
nand UO_1076 (O_1076,N_14975,N_14990);
nand UO_1077 (O_1077,N_14963,N_14935);
or UO_1078 (O_1078,N_14908,N_14901);
xnor UO_1079 (O_1079,N_14985,N_14895);
or UO_1080 (O_1080,N_14940,N_14913);
xor UO_1081 (O_1081,N_14951,N_14913);
nand UO_1082 (O_1082,N_14968,N_14964);
nor UO_1083 (O_1083,N_14896,N_14964);
xnor UO_1084 (O_1084,N_14941,N_14956);
xor UO_1085 (O_1085,N_14934,N_14954);
nor UO_1086 (O_1086,N_14911,N_14960);
nand UO_1087 (O_1087,N_14937,N_14883);
nand UO_1088 (O_1088,N_14937,N_14958);
or UO_1089 (O_1089,N_14937,N_14997);
nor UO_1090 (O_1090,N_14993,N_14954);
nand UO_1091 (O_1091,N_14947,N_14936);
xor UO_1092 (O_1092,N_14949,N_14913);
and UO_1093 (O_1093,N_14939,N_14995);
xor UO_1094 (O_1094,N_14969,N_14930);
or UO_1095 (O_1095,N_14895,N_14877);
or UO_1096 (O_1096,N_14967,N_14938);
xor UO_1097 (O_1097,N_14942,N_14882);
or UO_1098 (O_1098,N_14916,N_14905);
or UO_1099 (O_1099,N_14979,N_14896);
or UO_1100 (O_1100,N_14878,N_14875);
nor UO_1101 (O_1101,N_14977,N_14996);
and UO_1102 (O_1102,N_14939,N_14890);
xor UO_1103 (O_1103,N_14898,N_14941);
and UO_1104 (O_1104,N_14911,N_14929);
nor UO_1105 (O_1105,N_14985,N_14964);
nand UO_1106 (O_1106,N_14945,N_14996);
or UO_1107 (O_1107,N_14922,N_14981);
xor UO_1108 (O_1108,N_14936,N_14887);
nor UO_1109 (O_1109,N_14880,N_14912);
nand UO_1110 (O_1110,N_14895,N_14912);
or UO_1111 (O_1111,N_14962,N_14906);
nand UO_1112 (O_1112,N_14938,N_14916);
xor UO_1113 (O_1113,N_14974,N_14897);
xnor UO_1114 (O_1114,N_14938,N_14960);
nor UO_1115 (O_1115,N_14991,N_14941);
xor UO_1116 (O_1116,N_14883,N_14877);
nand UO_1117 (O_1117,N_14880,N_14938);
nand UO_1118 (O_1118,N_14876,N_14898);
or UO_1119 (O_1119,N_14963,N_14880);
and UO_1120 (O_1120,N_14932,N_14999);
nand UO_1121 (O_1121,N_14945,N_14954);
xnor UO_1122 (O_1122,N_14875,N_14909);
and UO_1123 (O_1123,N_14986,N_14929);
and UO_1124 (O_1124,N_14928,N_14889);
nand UO_1125 (O_1125,N_14890,N_14913);
xor UO_1126 (O_1126,N_14906,N_14878);
nor UO_1127 (O_1127,N_14918,N_14916);
xnor UO_1128 (O_1128,N_14952,N_14909);
xor UO_1129 (O_1129,N_14905,N_14875);
nor UO_1130 (O_1130,N_14975,N_14973);
nand UO_1131 (O_1131,N_14952,N_14890);
nor UO_1132 (O_1132,N_14887,N_14916);
nor UO_1133 (O_1133,N_14914,N_14938);
nor UO_1134 (O_1134,N_14992,N_14953);
and UO_1135 (O_1135,N_14914,N_14927);
nor UO_1136 (O_1136,N_14950,N_14886);
xnor UO_1137 (O_1137,N_14962,N_14979);
nor UO_1138 (O_1138,N_14904,N_14948);
nor UO_1139 (O_1139,N_14961,N_14919);
nand UO_1140 (O_1140,N_14915,N_14878);
nand UO_1141 (O_1141,N_14906,N_14999);
xnor UO_1142 (O_1142,N_14965,N_14936);
nand UO_1143 (O_1143,N_14885,N_14900);
and UO_1144 (O_1144,N_14962,N_14951);
or UO_1145 (O_1145,N_14981,N_14909);
nand UO_1146 (O_1146,N_14935,N_14888);
nand UO_1147 (O_1147,N_14888,N_14891);
and UO_1148 (O_1148,N_14903,N_14878);
or UO_1149 (O_1149,N_14910,N_14927);
or UO_1150 (O_1150,N_14889,N_14938);
xnor UO_1151 (O_1151,N_14992,N_14968);
xnor UO_1152 (O_1152,N_14972,N_14902);
nor UO_1153 (O_1153,N_14926,N_14980);
or UO_1154 (O_1154,N_14914,N_14916);
or UO_1155 (O_1155,N_14943,N_14951);
nand UO_1156 (O_1156,N_14969,N_14984);
and UO_1157 (O_1157,N_14911,N_14993);
xnor UO_1158 (O_1158,N_14963,N_14929);
nand UO_1159 (O_1159,N_14896,N_14901);
nand UO_1160 (O_1160,N_14917,N_14995);
and UO_1161 (O_1161,N_14983,N_14965);
and UO_1162 (O_1162,N_14877,N_14951);
xor UO_1163 (O_1163,N_14972,N_14971);
nand UO_1164 (O_1164,N_14921,N_14987);
nand UO_1165 (O_1165,N_14887,N_14881);
and UO_1166 (O_1166,N_14944,N_14964);
nor UO_1167 (O_1167,N_14916,N_14879);
xor UO_1168 (O_1168,N_14964,N_14965);
and UO_1169 (O_1169,N_14972,N_14987);
or UO_1170 (O_1170,N_14905,N_14933);
nor UO_1171 (O_1171,N_14946,N_14910);
and UO_1172 (O_1172,N_14878,N_14919);
nor UO_1173 (O_1173,N_14981,N_14938);
nand UO_1174 (O_1174,N_14910,N_14898);
and UO_1175 (O_1175,N_14891,N_14925);
nor UO_1176 (O_1176,N_14954,N_14884);
xor UO_1177 (O_1177,N_14979,N_14957);
nand UO_1178 (O_1178,N_14981,N_14940);
xnor UO_1179 (O_1179,N_14955,N_14918);
nand UO_1180 (O_1180,N_14988,N_14985);
nand UO_1181 (O_1181,N_14992,N_14880);
nor UO_1182 (O_1182,N_14961,N_14915);
nor UO_1183 (O_1183,N_14999,N_14931);
nand UO_1184 (O_1184,N_14937,N_14894);
nand UO_1185 (O_1185,N_14927,N_14930);
xor UO_1186 (O_1186,N_14939,N_14971);
xor UO_1187 (O_1187,N_14996,N_14911);
and UO_1188 (O_1188,N_14972,N_14947);
xnor UO_1189 (O_1189,N_14916,N_14977);
or UO_1190 (O_1190,N_14907,N_14899);
and UO_1191 (O_1191,N_14979,N_14996);
nand UO_1192 (O_1192,N_14983,N_14972);
and UO_1193 (O_1193,N_14941,N_14945);
nand UO_1194 (O_1194,N_14887,N_14907);
or UO_1195 (O_1195,N_14894,N_14892);
or UO_1196 (O_1196,N_14993,N_14953);
xor UO_1197 (O_1197,N_14927,N_14884);
and UO_1198 (O_1198,N_14961,N_14922);
xor UO_1199 (O_1199,N_14920,N_14943);
nor UO_1200 (O_1200,N_14918,N_14914);
xnor UO_1201 (O_1201,N_14990,N_14877);
and UO_1202 (O_1202,N_14917,N_14880);
xor UO_1203 (O_1203,N_14981,N_14876);
nand UO_1204 (O_1204,N_14936,N_14992);
or UO_1205 (O_1205,N_14898,N_14921);
nand UO_1206 (O_1206,N_14974,N_14934);
and UO_1207 (O_1207,N_14919,N_14877);
nand UO_1208 (O_1208,N_14927,N_14982);
or UO_1209 (O_1209,N_14935,N_14877);
and UO_1210 (O_1210,N_14961,N_14909);
xor UO_1211 (O_1211,N_14895,N_14991);
nand UO_1212 (O_1212,N_14976,N_14957);
nor UO_1213 (O_1213,N_14886,N_14987);
nand UO_1214 (O_1214,N_14902,N_14980);
and UO_1215 (O_1215,N_14922,N_14985);
and UO_1216 (O_1216,N_14966,N_14980);
and UO_1217 (O_1217,N_14958,N_14986);
xor UO_1218 (O_1218,N_14901,N_14936);
or UO_1219 (O_1219,N_14949,N_14934);
nor UO_1220 (O_1220,N_14941,N_14953);
nor UO_1221 (O_1221,N_14983,N_14899);
and UO_1222 (O_1222,N_14996,N_14989);
nor UO_1223 (O_1223,N_14895,N_14956);
or UO_1224 (O_1224,N_14977,N_14929);
and UO_1225 (O_1225,N_14996,N_14917);
xnor UO_1226 (O_1226,N_14996,N_14875);
nor UO_1227 (O_1227,N_14982,N_14976);
and UO_1228 (O_1228,N_14881,N_14924);
nand UO_1229 (O_1229,N_14962,N_14888);
or UO_1230 (O_1230,N_14890,N_14990);
nand UO_1231 (O_1231,N_14999,N_14981);
xnor UO_1232 (O_1232,N_14948,N_14894);
or UO_1233 (O_1233,N_14884,N_14912);
and UO_1234 (O_1234,N_14920,N_14928);
nor UO_1235 (O_1235,N_14974,N_14965);
xor UO_1236 (O_1236,N_14937,N_14948);
nand UO_1237 (O_1237,N_14941,N_14972);
nand UO_1238 (O_1238,N_14882,N_14963);
or UO_1239 (O_1239,N_14967,N_14970);
nand UO_1240 (O_1240,N_14915,N_14906);
or UO_1241 (O_1241,N_14926,N_14954);
or UO_1242 (O_1242,N_14920,N_14988);
and UO_1243 (O_1243,N_14923,N_14908);
and UO_1244 (O_1244,N_14929,N_14912);
or UO_1245 (O_1245,N_14949,N_14918);
xor UO_1246 (O_1246,N_14990,N_14879);
nand UO_1247 (O_1247,N_14988,N_14877);
nor UO_1248 (O_1248,N_14935,N_14958);
nor UO_1249 (O_1249,N_14982,N_14935);
xor UO_1250 (O_1250,N_14904,N_14987);
nand UO_1251 (O_1251,N_14997,N_14924);
xor UO_1252 (O_1252,N_14920,N_14916);
and UO_1253 (O_1253,N_14878,N_14893);
and UO_1254 (O_1254,N_14952,N_14971);
nand UO_1255 (O_1255,N_14981,N_14996);
nor UO_1256 (O_1256,N_14965,N_14971);
or UO_1257 (O_1257,N_14923,N_14941);
nor UO_1258 (O_1258,N_14936,N_14940);
nor UO_1259 (O_1259,N_14922,N_14955);
or UO_1260 (O_1260,N_14945,N_14905);
and UO_1261 (O_1261,N_14893,N_14966);
nor UO_1262 (O_1262,N_14877,N_14974);
and UO_1263 (O_1263,N_14903,N_14989);
nor UO_1264 (O_1264,N_14920,N_14970);
nand UO_1265 (O_1265,N_14909,N_14987);
nor UO_1266 (O_1266,N_14987,N_14952);
nor UO_1267 (O_1267,N_14904,N_14899);
nor UO_1268 (O_1268,N_14997,N_14945);
or UO_1269 (O_1269,N_14990,N_14995);
or UO_1270 (O_1270,N_14972,N_14906);
and UO_1271 (O_1271,N_14951,N_14971);
or UO_1272 (O_1272,N_14875,N_14938);
nor UO_1273 (O_1273,N_14975,N_14967);
xnor UO_1274 (O_1274,N_14985,N_14999);
or UO_1275 (O_1275,N_14934,N_14935);
nand UO_1276 (O_1276,N_14949,N_14999);
nand UO_1277 (O_1277,N_14925,N_14931);
nor UO_1278 (O_1278,N_14995,N_14948);
nand UO_1279 (O_1279,N_14931,N_14876);
xnor UO_1280 (O_1280,N_14878,N_14944);
nor UO_1281 (O_1281,N_14939,N_14983);
or UO_1282 (O_1282,N_14951,N_14879);
nor UO_1283 (O_1283,N_14982,N_14992);
xnor UO_1284 (O_1284,N_14903,N_14958);
and UO_1285 (O_1285,N_14919,N_14989);
or UO_1286 (O_1286,N_14999,N_14979);
and UO_1287 (O_1287,N_14947,N_14994);
nand UO_1288 (O_1288,N_14970,N_14917);
and UO_1289 (O_1289,N_14946,N_14965);
xor UO_1290 (O_1290,N_14917,N_14992);
nand UO_1291 (O_1291,N_14952,N_14892);
nand UO_1292 (O_1292,N_14879,N_14966);
xnor UO_1293 (O_1293,N_14928,N_14900);
nor UO_1294 (O_1294,N_14936,N_14894);
nand UO_1295 (O_1295,N_14907,N_14985);
and UO_1296 (O_1296,N_14912,N_14944);
and UO_1297 (O_1297,N_14919,N_14903);
nand UO_1298 (O_1298,N_14999,N_14996);
or UO_1299 (O_1299,N_14930,N_14940);
or UO_1300 (O_1300,N_14999,N_14991);
or UO_1301 (O_1301,N_14976,N_14876);
nor UO_1302 (O_1302,N_14930,N_14897);
or UO_1303 (O_1303,N_14913,N_14976);
nor UO_1304 (O_1304,N_14876,N_14968);
xor UO_1305 (O_1305,N_14910,N_14894);
or UO_1306 (O_1306,N_14911,N_14920);
nand UO_1307 (O_1307,N_14955,N_14984);
and UO_1308 (O_1308,N_14910,N_14913);
nand UO_1309 (O_1309,N_14912,N_14917);
nand UO_1310 (O_1310,N_14901,N_14950);
nand UO_1311 (O_1311,N_14948,N_14901);
and UO_1312 (O_1312,N_14921,N_14917);
nand UO_1313 (O_1313,N_14944,N_14952);
xnor UO_1314 (O_1314,N_14897,N_14978);
nand UO_1315 (O_1315,N_14914,N_14969);
xnor UO_1316 (O_1316,N_14969,N_14913);
nand UO_1317 (O_1317,N_14986,N_14911);
or UO_1318 (O_1318,N_14962,N_14916);
xnor UO_1319 (O_1319,N_14953,N_14973);
nand UO_1320 (O_1320,N_14885,N_14991);
nand UO_1321 (O_1321,N_14892,N_14887);
nor UO_1322 (O_1322,N_14963,N_14923);
xnor UO_1323 (O_1323,N_14991,N_14898);
and UO_1324 (O_1324,N_14907,N_14937);
xor UO_1325 (O_1325,N_14905,N_14889);
and UO_1326 (O_1326,N_14936,N_14989);
nand UO_1327 (O_1327,N_14935,N_14996);
and UO_1328 (O_1328,N_14959,N_14967);
or UO_1329 (O_1329,N_14908,N_14963);
and UO_1330 (O_1330,N_14932,N_14959);
xnor UO_1331 (O_1331,N_14981,N_14930);
nand UO_1332 (O_1332,N_14949,N_14985);
or UO_1333 (O_1333,N_14904,N_14962);
and UO_1334 (O_1334,N_14881,N_14921);
nor UO_1335 (O_1335,N_14888,N_14892);
xnor UO_1336 (O_1336,N_14908,N_14944);
and UO_1337 (O_1337,N_14897,N_14993);
nor UO_1338 (O_1338,N_14971,N_14940);
and UO_1339 (O_1339,N_14939,N_14929);
and UO_1340 (O_1340,N_14915,N_14971);
nand UO_1341 (O_1341,N_14989,N_14973);
nor UO_1342 (O_1342,N_14913,N_14886);
and UO_1343 (O_1343,N_14934,N_14919);
xnor UO_1344 (O_1344,N_14954,N_14992);
or UO_1345 (O_1345,N_14923,N_14957);
and UO_1346 (O_1346,N_14886,N_14918);
nor UO_1347 (O_1347,N_14946,N_14904);
or UO_1348 (O_1348,N_14933,N_14977);
and UO_1349 (O_1349,N_14971,N_14921);
nor UO_1350 (O_1350,N_14943,N_14891);
nand UO_1351 (O_1351,N_14928,N_14937);
nor UO_1352 (O_1352,N_14885,N_14902);
xnor UO_1353 (O_1353,N_14947,N_14938);
and UO_1354 (O_1354,N_14908,N_14918);
or UO_1355 (O_1355,N_14925,N_14949);
nor UO_1356 (O_1356,N_14952,N_14935);
or UO_1357 (O_1357,N_14980,N_14892);
xnor UO_1358 (O_1358,N_14983,N_14898);
nand UO_1359 (O_1359,N_14879,N_14984);
xor UO_1360 (O_1360,N_14990,N_14903);
nor UO_1361 (O_1361,N_14952,N_14891);
and UO_1362 (O_1362,N_14925,N_14965);
nand UO_1363 (O_1363,N_14875,N_14924);
nand UO_1364 (O_1364,N_14950,N_14909);
or UO_1365 (O_1365,N_14918,N_14891);
xnor UO_1366 (O_1366,N_14968,N_14977);
or UO_1367 (O_1367,N_14940,N_14912);
xnor UO_1368 (O_1368,N_14921,N_14905);
nor UO_1369 (O_1369,N_14948,N_14911);
or UO_1370 (O_1370,N_14905,N_14932);
nand UO_1371 (O_1371,N_14987,N_14926);
nand UO_1372 (O_1372,N_14956,N_14976);
nor UO_1373 (O_1373,N_14985,N_14941);
nand UO_1374 (O_1374,N_14923,N_14991);
nand UO_1375 (O_1375,N_14981,N_14942);
nand UO_1376 (O_1376,N_14923,N_14989);
and UO_1377 (O_1377,N_14916,N_14959);
and UO_1378 (O_1378,N_14967,N_14900);
nand UO_1379 (O_1379,N_14923,N_14897);
nor UO_1380 (O_1380,N_14955,N_14972);
xor UO_1381 (O_1381,N_14956,N_14938);
nand UO_1382 (O_1382,N_14938,N_14897);
or UO_1383 (O_1383,N_14893,N_14980);
xor UO_1384 (O_1384,N_14981,N_14974);
and UO_1385 (O_1385,N_14953,N_14997);
or UO_1386 (O_1386,N_14878,N_14937);
and UO_1387 (O_1387,N_14913,N_14905);
nor UO_1388 (O_1388,N_14924,N_14930);
or UO_1389 (O_1389,N_14994,N_14980);
or UO_1390 (O_1390,N_14960,N_14990);
xnor UO_1391 (O_1391,N_14989,N_14914);
nand UO_1392 (O_1392,N_14882,N_14875);
nand UO_1393 (O_1393,N_14986,N_14997);
or UO_1394 (O_1394,N_14949,N_14882);
nand UO_1395 (O_1395,N_14943,N_14999);
or UO_1396 (O_1396,N_14981,N_14927);
xor UO_1397 (O_1397,N_14999,N_14896);
nor UO_1398 (O_1398,N_14892,N_14878);
or UO_1399 (O_1399,N_14965,N_14945);
xnor UO_1400 (O_1400,N_14936,N_14974);
xnor UO_1401 (O_1401,N_14948,N_14952);
xnor UO_1402 (O_1402,N_14942,N_14893);
xor UO_1403 (O_1403,N_14937,N_14967);
nor UO_1404 (O_1404,N_14973,N_14970);
and UO_1405 (O_1405,N_14967,N_14880);
and UO_1406 (O_1406,N_14892,N_14939);
or UO_1407 (O_1407,N_14954,N_14879);
xnor UO_1408 (O_1408,N_14882,N_14994);
nor UO_1409 (O_1409,N_14899,N_14892);
xnor UO_1410 (O_1410,N_14982,N_14880);
nand UO_1411 (O_1411,N_14961,N_14972);
xnor UO_1412 (O_1412,N_14921,N_14984);
nor UO_1413 (O_1413,N_14952,N_14900);
nand UO_1414 (O_1414,N_14909,N_14876);
and UO_1415 (O_1415,N_14936,N_14915);
nand UO_1416 (O_1416,N_14883,N_14934);
nor UO_1417 (O_1417,N_14925,N_14985);
nor UO_1418 (O_1418,N_14911,N_14997);
nor UO_1419 (O_1419,N_14878,N_14888);
xor UO_1420 (O_1420,N_14943,N_14942);
nor UO_1421 (O_1421,N_14995,N_14987);
nand UO_1422 (O_1422,N_14961,N_14948);
nor UO_1423 (O_1423,N_14983,N_14896);
and UO_1424 (O_1424,N_14907,N_14947);
nor UO_1425 (O_1425,N_14906,N_14879);
xnor UO_1426 (O_1426,N_14914,N_14876);
or UO_1427 (O_1427,N_14924,N_14890);
and UO_1428 (O_1428,N_14950,N_14887);
xor UO_1429 (O_1429,N_14942,N_14930);
and UO_1430 (O_1430,N_14996,N_14957);
xnor UO_1431 (O_1431,N_14922,N_14963);
and UO_1432 (O_1432,N_14927,N_14929);
xnor UO_1433 (O_1433,N_14918,N_14929);
nor UO_1434 (O_1434,N_14954,N_14932);
nor UO_1435 (O_1435,N_14981,N_14899);
nand UO_1436 (O_1436,N_14889,N_14906);
nand UO_1437 (O_1437,N_14941,N_14978);
or UO_1438 (O_1438,N_14879,N_14967);
or UO_1439 (O_1439,N_14941,N_14992);
xor UO_1440 (O_1440,N_14937,N_14930);
xnor UO_1441 (O_1441,N_14986,N_14919);
or UO_1442 (O_1442,N_14883,N_14916);
or UO_1443 (O_1443,N_14928,N_14880);
xor UO_1444 (O_1444,N_14939,N_14976);
nand UO_1445 (O_1445,N_14899,N_14932);
and UO_1446 (O_1446,N_14882,N_14897);
or UO_1447 (O_1447,N_14980,N_14925);
or UO_1448 (O_1448,N_14998,N_14972);
xnor UO_1449 (O_1449,N_14999,N_14892);
nand UO_1450 (O_1450,N_14920,N_14980);
xor UO_1451 (O_1451,N_14984,N_14892);
and UO_1452 (O_1452,N_14890,N_14917);
and UO_1453 (O_1453,N_14929,N_14906);
nand UO_1454 (O_1454,N_14938,N_14886);
nor UO_1455 (O_1455,N_14893,N_14919);
or UO_1456 (O_1456,N_14960,N_14933);
nand UO_1457 (O_1457,N_14957,N_14935);
or UO_1458 (O_1458,N_14965,N_14996);
and UO_1459 (O_1459,N_14999,N_14983);
or UO_1460 (O_1460,N_14955,N_14970);
or UO_1461 (O_1461,N_14882,N_14948);
xnor UO_1462 (O_1462,N_14956,N_14878);
and UO_1463 (O_1463,N_14997,N_14971);
xor UO_1464 (O_1464,N_14885,N_14914);
xnor UO_1465 (O_1465,N_14894,N_14929);
nor UO_1466 (O_1466,N_14917,N_14962);
nand UO_1467 (O_1467,N_14987,N_14939);
xnor UO_1468 (O_1468,N_14976,N_14898);
or UO_1469 (O_1469,N_14926,N_14890);
nand UO_1470 (O_1470,N_14913,N_14991);
or UO_1471 (O_1471,N_14928,N_14913);
or UO_1472 (O_1472,N_14985,N_14912);
nor UO_1473 (O_1473,N_14990,N_14886);
and UO_1474 (O_1474,N_14918,N_14957);
xnor UO_1475 (O_1475,N_14917,N_14940);
and UO_1476 (O_1476,N_14926,N_14936);
xor UO_1477 (O_1477,N_14984,N_14928);
and UO_1478 (O_1478,N_14901,N_14907);
nand UO_1479 (O_1479,N_14972,N_14913);
and UO_1480 (O_1480,N_14985,N_14976);
and UO_1481 (O_1481,N_14935,N_14954);
and UO_1482 (O_1482,N_14976,N_14933);
nand UO_1483 (O_1483,N_14997,N_14925);
nand UO_1484 (O_1484,N_14897,N_14877);
xor UO_1485 (O_1485,N_14908,N_14998);
nand UO_1486 (O_1486,N_14993,N_14988);
or UO_1487 (O_1487,N_14900,N_14946);
nand UO_1488 (O_1488,N_14934,N_14898);
nand UO_1489 (O_1489,N_14987,N_14992);
nand UO_1490 (O_1490,N_14998,N_14941);
or UO_1491 (O_1491,N_14953,N_14961);
nor UO_1492 (O_1492,N_14984,N_14936);
xnor UO_1493 (O_1493,N_14945,N_14886);
xnor UO_1494 (O_1494,N_14929,N_14879);
nand UO_1495 (O_1495,N_14942,N_14892);
xor UO_1496 (O_1496,N_14961,N_14967);
xnor UO_1497 (O_1497,N_14962,N_14942);
xnor UO_1498 (O_1498,N_14906,N_14887);
nand UO_1499 (O_1499,N_14968,N_14925);
or UO_1500 (O_1500,N_14932,N_14949);
xnor UO_1501 (O_1501,N_14949,N_14922);
nand UO_1502 (O_1502,N_14966,N_14889);
nor UO_1503 (O_1503,N_14940,N_14979);
and UO_1504 (O_1504,N_14922,N_14996);
nor UO_1505 (O_1505,N_14923,N_14889);
nand UO_1506 (O_1506,N_14914,N_14908);
or UO_1507 (O_1507,N_14999,N_14933);
xor UO_1508 (O_1508,N_14984,N_14974);
or UO_1509 (O_1509,N_14885,N_14895);
nor UO_1510 (O_1510,N_14969,N_14983);
nor UO_1511 (O_1511,N_14984,N_14876);
and UO_1512 (O_1512,N_14893,N_14974);
and UO_1513 (O_1513,N_14913,N_14986);
and UO_1514 (O_1514,N_14975,N_14964);
or UO_1515 (O_1515,N_14876,N_14887);
nor UO_1516 (O_1516,N_14997,N_14999);
xor UO_1517 (O_1517,N_14920,N_14908);
nand UO_1518 (O_1518,N_14997,N_14910);
nor UO_1519 (O_1519,N_14939,N_14911);
and UO_1520 (O_1520,N_14932,N_14879);
nor UO_1521 (O_1521,N_14933,N_14956);
and UO_1522 (O_1522,N_14923,N_14895);
nand UO_1523 (O_1523,N_14954,N_14905);
and UO_1524 (O_1524,N_14895,N_14977);
xor UO_1525 (O_1525,N_14879,N_14964);
or UO_1526 (O_1526,N_14899,N_14903);
xor UO_1527 (O_1527,N_14879,N_14891);
and UO_1528 (O_1528,N_14945,N_14985);
and UO_1529 (O_1529,N_14964,N_14988);
xnor UO_1530 (O_1530,N_14894,N_14891);
and UO_1531 (O_1531,N_14940,N_14954);
and UO_1532 (O_1532,N_14954,N_14913);
and UO_1533 (O_1533,N_14984,N_14958);
nand UO_1534 (O_1534,N_14997,N_14938);
nor UO_1535 (O_1535,N_14976,N_14943);
or UO_1536 (O_1536,N_14961,N_14996);
or UO_1537 (O_1537,N_14981,N_14975);
xor UO_1538 (O_1538,N_14924,N_14947);
xor UO_1539 (O_1539,N_14998,N_14937);
nor UO_1540 (O_1540,N_14965,N_14994);
nand UO_1541 (O_1541,N_14921,N_14904);
nand UO_1542 (O_1542,N_14921,N_14952);
nand UO_1543 (O_1543,N_14970,N_14959);
or UO_1544 (O_1544,N_14985,N_14959);
xnor UO_1545 (O_1545,N_14893,N_14920);
or UO_1546 (O_1546,N_14895,N_14995);
or UO_1547 (O_1547,N_14899,N_14913);
xor UO_1548 (O_1548,N_14958,N_14900);
nand UO_1549 (O_1549,N_14913,N_14979);
nor UO_1550 (O_1550,N_14968,N_14996);
nand UO_1551 (O_1551,N_14882,N_14911);
xor UO_1552 (O_1552,N_14900,N_14893);
xor UO_1553 (O_1553,N_14891,N_14945);
nand UO_1554 (O_1554,N_14908,N_14883);
nand UO_1555 (O_1555,N_14926,N_14938);
nor UO_1556 (O_1556,N_14892,N_14889);
xor UO_1557 (O_1557,N_14973,N_14907);
nand UO_1558 (O_1558,N_14930,N_14968);
nand UO_1559 (O_1559,N_14899,N_14879);
and UO_1560 (O_1560,N_14914,N_14881);
or UO_1561 (O_1561,N_14931,N_14915);
or UO_1562 (O_1562,N_14908,N_14997);
or UO_1563 (O_1563,N_14978,N_14976);
or UO_1564 (O_1564,N_14919,N_14909);
nor UO_1565 (O_1565,N_14882,N_14895);
or UO_1566 (O_1566,N_14919,N_14922);
nor UO_1567 (O_1567,N_14937,N_14980);
nor UO_1568 (O_1568,N_14980,N_14983);
or UO_1569 (O_1569,N_14919,N_14940);
xnor UO_1570 (O_1570,N_14981,N_14983);
xor UO_1571 (O_1571,N_14925,N_14906);
nor UO_1572 (O_1572,N_14929,N_14892);
or UO_1573 (O_1573,N_14884,N_14932);
nor UO_1574 (O_1574,N_14969,N_14918);
or UO_1575 (O_1575,N_14981,N_14920);
or UO_1576 (O_1576,N_14890,N_14963);
or UO_1577 (O_1577,N_14935,N_14893);
nor UO_1578 (O_1578,N_14950,N_14986);
nor UO_1579 (O_1579,N_14882,N_14891);
nor UO_1580 (O_1580,N_14923,N_14968);
nand UO_1581 (O_1581,N_14923,N_14916);
xnor UO_1582 (O_1582,N_14886,N_14977);
nand UO_1583 (O_1583,N_14980,N_14883);
or UO_1584 (O_1584,N_14956,N_14935);
and UO_1585 (O_1585,N_14941,N_14969);
nand UO_1586 (O_1586,N_14887,N_14973);
or UO_1587 (O_1587,N_14999,N_14971);
or UO_1588 (O_1588,N_14924,N_14937);
or UO_1589 (O_1589,N_14952,N_14910);
nand UO_1590 (O_1590,N_14966,N_14957);
nor UO_1591 (O_1591,N_14942,N_14952);
or UO_1592 (O_1592,N_14957,N_14904);
nor UO_1593 (O_1593,N_14876,N_14958);
and UO_1594 (O_1594,N_14900,N_14963);
and UO_1595 (O_1595,N_14897,N_14893);
nor UO_1596 (O_1596,N_14883,N_14982);
or UO_1597 (O_1597,N_14945,N_14950);
nor UO_1598 (O_1598,N_14969,N_14937);
and UO_1599 (O_1599,N_14913,N_14878);
nand UO_1600 (O_1600,N_14930,N_14967);
xnor UO_1601 (O_1601,N_14882,N_14966);
and UO_1602 (O_1602,N_14972,N_14892);
nor UO_1603 (O_1603,N_14884,N_14942);
nand UO_1604 (O_1604,N_14993,N_14894);
xor UO_1605 (O_1605,N_14924,N_14894);
or UO_1606 (O_1606,N_14936,N_14962);
nand UO_1607 (O_1607,N_14926,N_14976);
xor UO_1608 (O_1608,N_14920,N_14891);
and UO_1609 (O_1609,N_14973,N_14966);
nor UO_1610 (O_1610,N_14989,N_14948);
xor UO_1611 (O_1611,N_14945,N_14986);
xnor UO_1612 (O_1612,N_14958,N_14951);
and UO_1613 (O_1613,N_14943,N_14876);
nor UO_1614 (O_1614,N_14892,N_14959);
or UO_1615 (O_1615,N_14966,N_14920);
and UO_1616 (O_1616,N_14942,N_14967);
xnor UO_1617 (O_1617,N_14897,N_14965);
or UO_1618 (O_1618,N_14977,N_14883);
and UO_1619 (O_1619,N_14995,N_14886);
and UO_1620 (O_1620,N_14934,N_14981);
nand UO_1621 (O_1621,N_14928,N_14903);
or UO_1622 (O_1622,N_14976,N_14890);
nand UO_1623 (O_1623,N_14974,N_14963);
and UO_1624 (O_1624,N_14919,N_14978);
nor UO_1625 (O_1625,N_14940,N_14970);
or UO_1626 (O_1626,N_14898,N_14956);
nor UO_1627 (O_1627,N_14944,N_14989);
or UO_1628 (O_1628,N_14881,N_14929);
or UO_1629 (O_1629,N_14920,N_14875);
or UO_1630 (O_1630,N_14897,N_14902);
nor UO_1631 (O_1631,N_14906,N_14930);
or UO_1632 (O_1632,N_14995,N_14920);
and UO_1633 (O_1633,N_14876,N_14932);
nor UO_1634 (O_1634,N_14891,N_14962);
or UO_1635 (O_1635,N_14916,N_14936);
or UO_1636 (O_1636,N_14933,N_14984);
and UO_1637 (O_1637,N_14894,N_14991);
nand UO_1638 (O_1638,N_14921,N_14935);
and UO_1639 (O_1639,N_14939,N_14928);
and UO_1640 (O_1640,N_14968,N_14938);
xor UO_1641 (O_1641,N_14981,N_14990);
nand UO_1642 (O_1642,N_14978,N_14946);
nand UO_1643 (O_1643,N_14889,N_14977);
or UO_1644 (O_1644,N_14888,N_14898);
xnor UO_1645 (O_1645,N_14905,N_14987);
xor UO_1646 (O_1646,N_14968,N_14943);
nor UO_1647 (O_1647,N_14897,N_14995);
xor UO_1648 (O_1648,N_14886,N_14985);
xor UO_1649 (O_1649,N_14976,N_14960);
xnor UO_1650 (O_1650,N_14986,N_14925);
xor UO_1651 (O_1651,N_14905,N_14937);
xnor UO_1652 (O_1652,N_14966,N_14975);
nor UO_1653 (O_1653,N_14883,N_14904);
nor UO_1654 (O_1654,N_14962,N_14892);
nor UO_1655 (O_1655,N_14982,N_14903);
nand UO_1656 (O_1656,N_14970,N_14974);
nor UO_1657 (O_1657,N_14970,N_14924);
nor UO_1658 (O_1658,N_14963,N_14966);
xor UO_1659 (O_1659,N_14877,N_14972);
or UO_1660 (O_1660,N_14895,N_14951);
nand UO_1661 (O_1661,N_14994,N_14991);
nor UO_1662 (O_1662,N_14956,N_14983);
xnor UO_1663 (O_1663,N_14971,N_14975);
and UO_1664 (O_1664,N_14950,N_14875);
xnor UO_1665 (O_1665,N_14903,N_14908);
or UO_1666 (O_1666,N_14944,N_14919);
and UO_1667 (O_1667,N_14940,N_14988);
and UO_1668 (O_1668,N_14889,N_14992);
xnor UO_1669 (O_1669,N_14916,N_14990);
xnor UO_1670 (O_1670,N_14978,N_14975);
and UO_1671 (O_1671,N_14906,N_14918);
nor UO_1672 (O_1672,N_14940,N_14882);
or UO_1673 (O_1673,N_14885,N_14945);
xor UO_1674 (O_1674,N_14951,N_14910);
and UO_1675 (O_1675,N_14932,N_14990);
nor UO_1676 (O_1676,N_14962,N_14955);
nand UO_1677 (O_1677,N_14903,N_14927);
and UO_1678 (O_1678,N_14924,N_14938);
xor UO_1679 (O_1679,N_14960,N_14889);
nor UO_1680 (O_1680,N_14936,N_14902);
and UO_1681 (O_1681,N_14915,N_14902);
nor UO_1682 (O_1682,N_14881,N_14967);
or UO_1683 (O_1683,N_14944,N_14998);
xor UO_1684 (O_1684,N_14878,N_14880);
or UO_1685 (O_1685,N_14920,N_14903);
nand UO_1686 (O_1686,N_14891,N_14908);
nor UO_1687 (O_1687,N_14896,N_14886);
and UO_1688 (O_1688,N_14883,N_14970);
or UO_1689 (O_1689,N_14982,N_14932);
xnor UO_1690 (O_1690,N_14932,N_14927);
and UO_1691 (O_1691,N_14962,N_14948);
and UO_1692 (O_1692,N_14875,N_14889);
or UO_1693 (O_1693,N_14887,N_14979);
or UO_1694 (O_1694,N_14943,N_14988);
or UO_1695 (O_1695,N_14979,N_14946);
xnor UO_1696 (O_1696,N_14971,N_14879);
nand UO_1697 (O_1697,N_14900,N_14948);
and UO_1698 (O_1698,N_14958,N_14914);
nand UO_1699 (O_1699,N_14934,N_14964);
nor UO_1700 (O_1700,N_14949,N_14894);
xor UO_1701 (O_1701,N_14975,N_14989);
nor UO_1702 (O_1702,N_14939,N_14966);
and UO_1703 (O_1703,N_14894,N_14979);
xnor UO_1704 (O_1704,N_14920,N_14958);
xnor UO_1705 (O_1705,N_14991,N_14917);
nand UO_1706 (O_1706,N_14899,N_14998);
nor UO_1707 (O_1707,N_14911,N_14895);
nor UO_1708 (O_1708,N_14876,N_14994);
and UO_1709 (O_1709,N_14986,N_14905);
xnor UO_1710 (O_1710,N_14897,N_14989);
xor UO_1711 (O_1711,N_14940,N_14995);
nand UO_1712 (O_1712,N_14901,N_14902);
or UO_1713 (O_1713,N_14878,N_14936);
and UO_1714 (O_1714,N_14967,N_14913);
and UO_1715 (O_1715,N_14887,N_14999);
xor UO_1716 (O_1716,N_14909,N_14906);
and UO_1717 (O_1717,N_14899,N_14928);
nor UO_1718 (O_1718,N_14932,N_14986);
or UO_1719 (O_1719,N_14949,N_14883);
nand UO_1720 (O_1720,N_14901,N_14982);
or UO_1721 (O_1721,N_14906,N_14931);
nor UO_1722 (O_1722,N_14973,N_14998);
and UO_1723 (O_1723,N_14888,N_14984);
nand UO_1724 (O_1724,N_14937,N_14886);
or UO_1725 (O_1725,N_14991,N_14915);
xnor UO_1726 (O_1726,N_14934,N_14976);
nand UO_1727 (O_1727,N_14951,N_14932);
nand UO_1728 (O_1728,N_14958,N_14899);
nand UO_1729 (O_1729,N_14981,N_14903);
xnor UO_1730 (O_1730,N_14939,N_14893);
and UO_1731 (O_1731,N_14923,N_14993);
xnor UO_1732 (O_1732,N_14936,N_14970);
and UO_1733 (O_1733,N_14971,N_14994);
nand UO_1734 (O_1734,N_14929,N_14992);
or UO_1735 (O_1735,N_14905,N_14961);
xnor UO_1736 (O_1736,N_14919,N_14956);
or UO_1737 (O_1737,N_14899,N_14946);
and UO_1738 (O_1738,N_14930,N_14948);
nand UO_1739 (O_1739,N_14887,N_14924);
nor UO_1740 (O_1740,N_14880,N_14900);
or UO_1741 (O_1741,N_14910,N_14934);
nand UO_1742 (O_1742,N_14938,N_14879);
nand UO_1743 (O_1743,N_14930,N_14878);
xnor UO_1744 (O_1744,N_14956,N_14914);
nor UO_1745 (O_1745,N_14961,N_14892);
or UO_1746 (O_1746,N_14885,N_14958);
xnor UO_1747 (O_1747,N_14957,N_14980);
nor UO_1748 (O_1748,N_14902,N_14986);
and UO_1749 (O_1749,N_14937,N_14880);
or UO_1750 (O_1750,N_14888,N_14928);
or UO_1751 (O_1751,N_14957,N_14933);
xnor UO_1752 (O_1752,N_14977,N_14892);
nor UO_1753 (O_1753,N_14927,N_14980);
and UO_1754 (O_1754,N_14914,N_14931);
nor UO_1755 (O_1755,N_14914,N_14976);
xor UO_1756 (O_1756,N_14897,N_14889);
xor UO_1757 (O_1757,N_14981,N_14918);
nand UO_1758 (O_1758,N_14939,N_14948);
nor UO_1759 (O_1759,N_14902,N_14990);
and UO_1760 (O_1760,N_14949,N_14951);
or UO_1761 (O_1761,N_14931,N_14943);
xor UO_1762 (O_1762,N_14934,N_14938);
nand UO_1763 (O_1763,N_14942,N_14960);
or UO_1764 (O_1764,N_14948,N_14888);
xnor UO_1765 (O_1765,N_14995,N_14961);
nand UO_1766 (O_1766,N_14898,N_14986);
xnor UO_1767 (O_1767,N_14916,N_14979);
or UO_1768 (O_1768,N_14901,N_14894);
and UO_1769 (O_1769,N_14994,N_14911);
nand UO_1770 (O_1770,N_14892,N_14875);
nor UO_1771 (O_1771,N_14972,N_14937);
nand UO_1772 (O_1772,N_14949,N_14976);
or UO_1773 (O_1773,N_14881,N_14987);
xor UO_1774 (O_1774,N_14895,N_14987);
nor UO_1775 (O_1775,N_14876,N_14901);
nor UO_1776 (O_1776,N_14980,N_14876);
xnor UO_1777 (O_1777,N_14906,N_14883);
xnor UO_1778 (O_1778,N_14932,N_14973);
nand UO_1779 (O_1779,N_14951,N_14968);
nor UO_1780 (O_1780,N_14930,N_14977);
nand UO_1781 (O_1781,N_14927,N_14923);
xnor UO_1782 (O_1782,N_14977,N_14907);
or UO_1783 (O_1783,N_14930,N_14876);
nand UO_1784 (O_1784,N_14983,N_14985);
nor UO_1785 (O_1785,N_14948,N_14985);
or UO_1786 (O_1786,N_14941,N_14966);
nor UO_1787 (O_1787,N_14885,N_14949);
nand UO_1788 (O_1788,N_14999,N_14988);
nor UO_1789 (O_1789,N_14953,N_14933);
and UO_1790 (O_1790,N_14929,N_14920);
nor UO_1791 (O_1791,N_14970,N_14909);
nor UO_1792 (O_1792,N_14987,N_14978);
nand UO_1793 (O_1793,N_14931,N_14989);
nand UO_1794 (O_1794,N_14935,N_14898);
nor UO_1795 (O_1795,N_14937,N_14889);
and UO_1796 (O_1796,N_14974,N_14916);
or UO_1797 (O_1797,N_14896,N_14924);
nand UO_1798 (O_1798,N_14900,N_14964);
xnor UO_1799 (O_1799,N_14895,N_14886);
nor UO_1800 (O_1800,N_14880,N_14892);
xor UO_1801 (O_1801,N_14920,N_14892);
and UO_1802 (O_1802,N_14891,N_14885);
nand UO_1803 (O_1803,N_14954,N_14931);
and UO_1804 (O_1804,N_14954,N_14877);
nor UO_1805 (O_1805,N_14971,N_14896);
nor UO_1806 (O_1806,N_14925,N_14920);
or UO_1807 (O_1807,N_14984,N_14994);
nor UO_1808 (O_1808,N_14876,N_14925);
nand UO_1809 (O_1809,N_14959,N_14904);
or UO_1810 (O_1810,N_14885,N_14904);
or UO_1811 (O_1811,N_14980,N_14939);
or UO_1812 (O_1812,N_14931,N_14886);
and UO_1813 (O_1813,N_14894,N_14899);
nor UO_1814 (O_1814,N_14922,N_14940);
or UO_1815 (O_1815,N_14988,N_14991);
nand UO_1816 (O_1816,N_14912,N_14957);
nor UO_1817 (O_1817,N_14975,N_14910);
nor UO_1818 (O_1818,N_14944,N_14990);
nand UO_1819 (O_1819,N_14908,N_14886);
and UO_1820 (O_1820,N_14973,N_14904);
nand UO_1821 (O_1821,N_14896,N_14917);
nor UO_1822 (O_1822,N_14933,N_14970);
nor UO_1823 (O_1823,N_14963,N_14916);
and UO_1824 (O_1824,N_14899,N_14900);
nand UO_1825 (O_1825,N_14953,N_14966);
nor UO_1826 (O_1826,N_14894,N_14904);
or UO_1827 (O_1827,N_14926,N_14952);
nor UO_1828 (O_1828,N_14886,N_14883);
nor UO_1829 (O_1829,N_14989,N_14878);
xor UO_1830 (O_1830,N_14949,N_14900);
or UO_1831 (O_1831,N_14907,N_14904);
or UO_1832 (O_1832,N_14920,N_14886);
nor UO_1833 (O_1833,N_14940,N_14987);
nand UO_1834 (O_1834,N_14898,N_14926);
nor UO_1835 (O_1835,N_14926,N_14877);
nand UO_1836 (O_1836,N_14906,N_14997);
nand UO_1837 (O_1837,N_14978,N_14981);
nor UO_1838 (O_1838,N_14893,N_14886);
nor UO_1839 (O_1839,N_14966,N_14960);
nand UO_1840 (O_1840,N_14933,N_14992);
or UO_1841 (O_1841,N_14958,N_14946);
nor UO_1842 (O_1842,N_14906,N_14901);
and UO_1843 (O_1843,N_14985,N_14992);
nand UO_1844 (O_1844,N_14982,N_14907);
nand UO_1845 (O_1845,N_14983,N_14940);
and UO_1846 (O_1846,N_14999,N_14946);
or UO_1847 (O_1847,N_14875,N_14885);
and UO_1848 (O_1848,N_14900,N_14974);
nor UO_1849 (O_1849,N_14942,N_14950);
or UO_1850 (O_1850,N_14999,N_14966);
nor UO_1851 (O_1851,N_14916,N_14943);
and UO_1852 (O_1852,N_14997,N_14914);
and UO_1853 (O_1853,N_14954,N_14949);
nand UO_1854 (O_1854,N_14928,N_14990);
nand UO_1855 (O_1855,N_14944,N_14999);
nor UO_1856 (O_1856,N_14993,N_14952);
and UO_1857 (O_1857,N_14926,N_14969);
nand UO_1858 (O_1858,N_14931,N_14930);
or UO_1859 (O_1859,N_14977,N_14878);
or UO_1860 (O_1860,N_14961,N_14924);
and UO_1861 (O_1861,N_14936,N_14949);
nor UO_1862 (O_1862,N_14944,N_14926);
xnor UO_1863 (O_1863,N_14982,N_14979);
nor UO_1864 (O_1864,N_14906,N_14892);
and UO_1865 (O_1865,N_14901,N_14974);
nor UO_1866 (O_1866,N_14894,N_14953);
xnor UO_1867 (O_1867,N_14894,N_14913);
and UO_1868 (O_1868,N_14926,N_14931);
or UO_1869 (O_1869,N_14952,N_14897);
and UO_1870 (O_1870,N_14987,N_14900);
or UO_1871 (O_1871,N_14903,N_14997);
or UO_1872 (O_1872,N_14980,N_14998);
nand UO_1873 (O_1873,N_14934,N_14884);
and UO_1874 (O_1874,N_14900,N_14935);
or UO_1875 (O_1875,N_14886,N_14949);
nor UO_1876 (O_1876,N_14959,N_14994);
nor UO_1877 (O_1877,N_14933,N_14895);
and UO_1878 (O_1878,N_14935,N_14971);
nand UO_1879 (O_1879,N_14953,N_14875);
nor UO_1880 (O_1880,N_14954,N_14895);
or UO_1881 (O_1881,N_14958,N_14997);
and UO_1882 (O_1882,N_14930,N_14883);
nor UO_1883 (O_1883,N_14916,N_14937);
nand UO_1884 (O_1884,N_14933,N_14954);
nor UO_1885 (O_1885,N_14977,N_14898);
or UO_1886 (O_1886,N_14923,N_14880);
xor UO_1887 (O_1887,N_14972,N_14966);
or UO_1888 (O_1888,N_14987,N_14875);
xnor UO_1889 (O_1889,N_14881,N_14925);
xor UO_1890 (O_1890,N_14913,N_14929);
nand UO_1891 (O_1891,N_14977,N_14990);
nand UO_1892 (O_1892,N_14891,N_14900);
xnor UO_1893 (O_1893,N_14909,N_14984);
nand UO_1894 (O_1894,N_14883,N_14895);
or UO_1895 (O_1895,N_14979,N_14923);
or UO_1896 (O_1896,N_14918,N_14895);
and UO_1897 (O_1897,N_14928,N_14944);
nor UO_1898 (O_1898,N_14926,N_14975);
and UO_1899 (O_1899,N_14995,N_14959);
and UO_1900 (O_1900,N_14988,N_14966);
xor UO_1901 (O_1901,N_14949,N_14988);
nor UO_1902 (O_1902,N_14951,N_14995);
nor UO_1903 (O_1903,N_14884,N_14915);
or UO_1904 (O_1904,N_14967,N_14988);
xor UO_1905 (O_1905,N_14963,N_14978);
or UO_1906 (O_1906,N_14897,N_14949);
and UO_1907 (O_1907,N_14953,N_14939);
and UO_1908 (O_1908,N_14983,N_14882);
xor UO_1909 (O_1909,N_14944,N_14943);
xnor UO_1910 (O_1910,N_14891,N_14922);
nor UO_1911 (O_1911,N_14918,N_14913);
xor UO_1912 (O_1912,N_14990,N_14999);
xnor UO_1913 (O_1913,N_14878,N_14908);
xnor UO_1914 (O_1914,N_14971,N_14987);
nand UO_1915 (O_1915,N_14897,N_14934);
and UO_1916 (O_1916,N_14901,N_14885);
xor UO_1917 (O_1917,N_14890,N_14988);
nor UO_1918 (O_1918,N_14986,N_14981);
or UO_1919 (O_1919,N_14955,N_14939);
nor UO_1920 (O_1920,N_14968,N_14881);
xnor UO_1921 (O_1921,N_14907,N_14964);
and UO_1922 (O_1922,N_14929,N_14970);
or UO_1923 (O_1923,N_14875,N_14976);
nand UO_1924 (O_1924,N_14977,N_14986);
or UO_1925 (O_1925,N_14901,N_14945);
nand UO_1926 (O_1926,N_14910,N_14995);
xor UO_1927 (O_1927,N_14898,N_14952);
nor UO_1928 (O_1928,N_14918,N_14943);
and UO_1929 (O_1929,N_14974,N_14908);
xor UO_1930 (O_1930,N_14885,N_14937);
and UO_1931 (O_1931,N_14984,N_14932);
nand UO_1932 (O_1932,N_14916,N_14878);
or UO_1933 (O_1933,N_14924,N_14972);
and UO_1934 (O_1934,N_14930,N_14956);
nor UO_1935 (O_1935,N_14962,N_14976);
nor UO_1936 (O_1936,N_14930,N_14984);
nand UO_1937 (O_1937,N_14926,N_14966);
and UO_1938 (O_1938,N_14970,N_14949);
nor UO_1939 (O_1939,N_14939,N_14875);
nor UO_1940 (O_1940,N_14911,N_14969);
nor UO_1941 (O_1941,N_14972,N_14930);
and UO_1942 (O_1942,N_14974,N_14998);
or UO_1943 (O_1943,N_14982,N_14953);
or UO_1944 (O_1944,N_14907,N_14932);
nand UO_1945 (O_1945,N_14964,N_14928);
nor UO_1946 (O_1946,N_14957,N_14954);
nor UO_1947 (O_1947,N_14894,N_14975);
nand UO_1948 (O_1948,N_14989,N_14887);
and UO_1949 (O_1949,N_14884,N_14929);
nor UO_1950 (O_1950,N_14954,N_14888);
or UO_1951 (O_1951,N_14993,N_14997);
xnor UO_1952 (O_1952,N_14946,N_14916);
nand UO_1953 (O_1953,N_14980,N_14947);
nor UO_1954 (O_1954,N_14959,N_14895);
xnor UO_1955 (O_1955,N_14992,N_14919);
or UO_1956 (O_1956,N_14907,N_14990);
and UO_1957 (O_1957,N_14879,N_14908);
nand UO_1958 (O_1958,N_14959,N_14894);
and UO_1959 (O_1959,N_14946,N_14954);
nor UO_1960 (O_1960,N_14986,N_14974);
xor UO_1961 (O_1961,N_14926,N_14882);
or UO_1962 (O_1962,N_14875,N_14908);
and UO_1963 (O_1963,N_14890,N_14972);
or UO_1964 (O_1964,N_14933,N_14972);
and UO_1965 (O_1965,N_14887,N_14875);
and UO_1966 (O_1966,N_14965,N_14919);
nor UO_1967 (O_1967,N_14960,N_14967);
nor UO_1968 (O_1968,N_14881,N_14913);
or UO_1969 (O_1969,N_14964,N_14961);
nor UO_1970 (O_1970,N_14971,N_14929);
and UO_1971 (O_1971,N_14972,N_14897);
and UO_1972 (O_1972,N_14927,N_14983);
and UO_1973 (O_1973,N_14891,N_14876);
nand UO_1974 (O_1974,N_14959,N_14953);
xnor UO_1975 (O_1975,N_14993,N_14933);
nor UO_1976 (O_1976,N_14985,N_14897);
nor UO_1977 (O_1977,N_14928,N_14915);
nand UO_1978 (O_1978,N_14922,N_14967);
nand UO_1979 (O_1979,N_14921,N_14993);
xor UO_1980 (O_1980,N_14923,N_14997);
and UO_1981 (O_1981,N_14987,N_14993);
or UO_1982 (O_1982,N_14884,N_14879);
xnor UO_1983 (O_1983,N_14920,N_14904);
or UO_1984 (O_1984,N_14907,N_14989);
or UO_1985 (O_1985,N_14906,N_14967);
nand UO_1986 (O_1986,N_14940,N_14953);
nor UO_1987 (O_1987,N_14991,N_14882);
and UO_1988 (O_1988,N_14895,N_14894);
or UO_1989 (O_1989,N_14935,N_14903);
nand UO_1990 (O_1990,N_14990,N_14908);
and UO_1991 (O_1991,N_14977,N_14991);
nor UO_1992 (O_1992,N_14886,N_14899);
nor UO_1993 (O_1993,N_14967,N_14890);
or UO_1994 (O_1994,N_14921,N_14939);
or UO_1995 (O_1995,N_14949,N_14884);
or UO_1996 (O_1996,N_14969,N_14978);
or UO_1997 (O_1997,N_14937,N_14892);
nand UO_1998 (O_1998,N_14893,N_14993);
nand UO_1999 (O_1999,N_14937,N_14917);
endmodule