module basic_1500_15000_2000_75_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_497,In_97);
or U1 (N_1,In_1112,In_1435);
or U2 (N_2,In_676,In_1145);
and U3 (N_3,In_1342,In_208);
and U4 (N_4,In_574,In_866);
xor U5 (N_5,In_1488,In_1461);
nor U6 (N_6,In_737,In_1275);
xor U7 (N_7,In_1257,In_20);
xnor U8 (N_8,In_453,In_539);
or U9 (N_9,In_1496,In_157);
xnor U10 (N_10,In_1068,In_1181);
nor U11 (N_11,In_486,In_1439);
xnor U12 (N_12,In_15,In_1369);
xor U13 (N_13,In_10,In_594);
and U14 (N_14,In_1360,In_333);
xor U15 (N_15,In_1373,In_348);
or U16 (N_16,In_1027,In_52);
and U17 (N_17,In_409,In_634);
or U18 (N_18,In_789,In_797);
xnor U19 (N_19,In_806,In_767);
or U20 (N_20,In_440,In_163);
nand U21 (N_21,In_1440,In_295);
xnor U22 (N_22,In_959,In_721);
and U23 (N_23,In_808,In_729);
and U24 (N_24,In_1491,In_1278);
and U25 (N_25,In_108,In_711);
nand U26 (N_26,In_469,In_1333);
nor U27 (N_27,In_533,In_75);
or U28 (N_28,In_11,In_1290);
and U29 (N_29,In_1253,In_1127);
and U30 (N_30,In_918,In_404);
or U31 (N_31,In_1398,In_937);
nand U32 (N_32,In_981,In_759);
nor U33 (N_33,In_383,In_1131);
nand U34 (N_34,In_1429,In_719);
nor U35 (N_35,In_1051,In_1362);
and U36 (N_36,In_1041,In_917);
nor U37 (N_37,In_1144,In_600);
and U38 (N_38,In_876,In_332);
xnor U39 (N_39,In_1138,In_1229);
nor U40 (N_40,In_251,In_940);
and U41 (N_41,In_335,In_458);
or U42 (N_42,In_1326,In_1416);
or U43 (N_43,In_254,In_1106);
xor U44 (N_44,In_1281,In_1391);
and U45 (N_45,In_955,In_727);
xor U46 (N_46,In_285,In_774);
and U47 (N_47,In_1166,In_951);
nor U48 (N_48,In_1334,In_339);
nor U49 (N_49,In_479,In_896);
or U50 (N_50,In_1011,In_869);
and U51 (N_51,In_323,In_669);
or U52 (N_52,In_752,In_903);
xnor U53 (N_53,In_985,In_381);
nor U54 (N_54,In_452,In_1339);
or U55 (N_55,In_631,In_893);
nor U56 (N_56,In_228,In_670);
and U57 (N_57,In_167,In_59);
xor U58 (N_58,In_1483,In_121);
xnor U59 (N_59,In_1350,In_186);
xor U60 (N_60,In_654,In_60);
and U61 (N_61,In_831,In_1366);
nor U62 (N_62,In_708,In_596);
nor U63 (N_63,In_1256,In_1252);
nand U64 (N_64,In_93,In_357);
nand U65 (N_65,In_256,In_1421);
nor U66 (N_66,In_141,In_1409);
and U67 (N_67,In_907,In_1235);
and U68 (N_68,In_441,In_130);
or U69 (N_69,In_198,In_1161);
and U70 (N_70,In_552,In_832);
nor U71 (N_71,In_1262,In_1167);
nor U72 (N_72,In_1220,In_1207);
nand U73 (N_73,In_517,In_143);
nand U74 (N_74,In_480,In_1282);
nor U75 (N_75,In_360,In_783);
nor U76 (N_76,In_21,In_712);
nand U77 (N_77,In_347,In_742);
nor U78 (N_78,In_992,In_550);
nor U79 (N_79,In_1427,In_385);
xnor U80 (N_80,In_697,In_769);
xnor U81 (N_81,In_883,In_505);
nor U82 (N_82,In_28,In_1447);
xor U83 (N_83,In_144,In_1469);
xnor U84 (N_84,In_662,In_575);
xnor U85 (N_85,In_126,In_111);
or U86 (N_86,In_588,In_867);
nand U87 (N_87,In_665,In_1395);
xnor U88 (N_88,In_1316,In_34);
nor U89 (N_89,In_1089,In_1283);
or U90 (N_90,In_77,In_1266);
xor U91 (N_91,In_656,In_399);
xnor U92 (N_92,In_33,In_1345);
and U93 (N_93,In_630,In_948);
or U94 (N_94,In_43,In_154);
or U95 (N_95,In_1265,In_403);
nor U96 (N_96,In_201,In_1441);
nand U97 (N_97,In_64,In_688);
xor U98 (N_98,In_565,In_734);
nand U99 (N_99,In_246,In_1237);
and U100 (N_100,In_725,In_865);
or U101 (N_101,In_42,In_790);
xnor U102 (N_102,In_1132,In_2);
nand U103 (N_103,In_1038,In_816);
nor U104 (N_104,In_267,In_459);
xnor U105 (N_105,In_1155,In_1087);
and U106 (N_106,In_997,In_1174);
and U107 (N_107,In_1411,In_788);
xor U108 (N_108,In_760,In_221);
nand U109 (N_109,In_417,In_1343);
or U110 (N_110,In_1444,In_1486);
xnor U111 (N_111,In_975,In_672);
and U112 (N_112,In_1116,In_1086);
and U113 (N_113,In_4,In_873);
and U114 (N_114,In_1241,In_26);
and U115 (N_115,In_643,In_193);
or U116 (N_116,In_214,In_794);
or U117 (N_117,In_1341,In_1016);
nand U118 (N_118,In_1471,In_442);
xnor U119 (N_119,In_1250,In_1296);
nand U120 (N_120,In_1284,In_107);
nand U121 (N_121,In_912,In_570);
nand U122 (N_122,In_1219,In_319);
and U123 (N_123,In_636,In_835);
xnor U124 (N_124,In_197,In_755);
nor U125 (N_125,In_217,In_1104);
xor U126 (N_126,In_1045,In_142);
and U127 (N_127,In_365,In_1289);
nand U128 (N_128,In_950,In_444);
xnor U129 (N_129,In_36,In_1414);
nor U130 (N_130,In_651,In_1269);
nor U131 (N_131,In_65,In_870);
nor U132 (N_132,In_996,In_1165);
nor U133 (N_133,In_1193,In_0);
nand U134 (N_134,In_1053,In_1497);
xnor U135 (N_135,In_1020,In_922);
xor U136 (N_136,In_1249,In_689);
or U137 (N_137,In_1128,In_560);
or U138 (N_138,In_296,In_987);
nor U139 (N_139,In_164,In_663);
nand U140 (N_140,In_352,In_84);
nor U141 (N_141,In_1094,In_109);
or U142 (N_142,In_943,In_946);
xnor U143 (N_143,In_844,In_438);
or U144 (N_144,In_477,In_1005);
xor U145 (N_145,In_1147,In_465);
and U146 (N_146,In_340,In_523);
or U147 (N_147,In_915,In_1099);
nor U148 (N_148,In_529,In_801);
nor U149 (N_149,In_1494,In_1493);
xor U150 (N_150,In_590,In_681);
xnor U151 (N_151,In_50,In_1291);
and U152 (N_152,In_633,In_956);
nor U153 (N_153,In_294,In_841);
and U154 (N_154,In_674,In_1470);
and U155 (N_155,In_1247,In_259);
and U156 (N_156,In_724,In_472);
and U157 (N_157,In_14,In_484);
nand U158 (N_158,In_990,In_668);
nand U159 (N_159,In_1003,In_436);
or U160 (N_160,In_1372,In_1019);
xnor U161 (N_161,In_435,In_610);
xnor U162 (N_162,In_1209,In_117);
xor U163 (N_163,In_976,In_572);
and U164 (N_164,In_382,In_970);
or U165 (N_165,In_258,In_232);
nor U166 (N_166,In_543,In_351);
or U167 (N_167,In_276,In_977);
xor U168 (N_168,In_1312,In_1190);
and U169 (N_169,In_1160,In_936);
or U170 (N_170,In_1029,In_847);
xnor U171 (N_171,In_836,In_1036);
nand U172 (N_172,In_413,In_326);
nand U173 (N_173,In_1443,In_1319);
nand U174 (N_174,In_1150,In_751);
or U175 (N_175,In_764,In_1212);
xnor U176 (N_176,In_377,In_1404);
nand U177 (N_177,In_671,In_799);
and U178 (N_178,In_1069,In_1472);
and U179 (N_179,In_1495,In_40);
or U180 (N_180,In_1168,In_342);
xnor U181 (N_181,In_1210,In_564);
nor U182 (N_182,In_1157,In_625);
xnor U183 (N_183,In_642,In_705);
or U184 (N_184,In_1308,In_886);
nor U185 (N_185,In_297,In_245);
or U186 (N_186,In_334,In_1426);
nand U187 (N_187,In_1438,In_880);
or U188 (N_188,In_255,In_57);
and U189 (N_189,In_603,In_447);
and U190 (N_190,In_1322,In_279);
nand U191 (N_191,In_895,In_1000);
and U192 (N_192,In_1349,In_1385);
xor U193 (N_193,In_1139,In_1037);
nor U194 (N_194,In_924,In_73);
and U195 (N_195,In_1254,In_1022);
or U196 (N_196,In_96,In_1180);
xnor U197 (N_197,In_115,In_1240);
xnor U198 (N_198,In_1057,In_118);
xnor U199 (N_199,In_703,In_78);
nor U200 (N_200,In_29,In_207);
and U201 (N_201,In_168,N_188);
or U202 (N_202,N_169,In_584);
nand U203 (N_203,In_45,In_682);
nand U204 (N_204,In_778,In_1182);
and U205 (N_205,In_1121,N_55);
nand U206 (N_206,In_1081,N_97);
nor U207 (N_207,In_1232,In_849);
nand U208 (N_208,In_1058,In_1042);
or U209 (N_209,In_723,In_104);
nand U210 (N_210,In_470,In_1039);
nand U211 (N_211,In_765,In_1332);
xnor U212 (N_212,In_1090,N_0);
nor U213 (N_213,N_58,In_942);
nor U214 (N_214,In_820,In_1474);
xnor U215 (N_215,In_317,In_780);
nand U216 (N_216,In_1422,N_133);
nand U217 (N_217,N_161,In_514);
and U218 (N_218,In_1375,In_113);
or U219 (N_219,In_137,In_1134);
and U220 (N_220,In_1030,In_1006);
nand U221 (N_221,In_1007,In_967);
nand U222 (N_222,In_1453,In_763);
nor U223 (N_223,In_49,N_157);
nand U224 (N_224,In_938,In_1076);
nand U225 (N_225,In_978,In_945);
xor U226 (N_226,In_415,In_349);
nand U227 (N_227,N_23,In_81);
xor U228 (N_228,In_645,N_33);
and U229 (N_229,In_746,In_451);
or U230 (N_230,In_1091,N_147);
nand U231 (N_231,In_1335,N_87);
and U232 (N_232,In_839,In_1218);
nand U233 (N_233,In_919,In_772);
and U234 (N_234,N_65,N_152);
or U235 (N_235,In_798,In_134);
nand U236 (N_236,In_973,In_58);
nor U237 (N_237,In_388,In_927);
nand U238 (N_238,In_785,In_454);
nor U239 (N_239,In_1133,In_678);
nand U240 (N_240,N_69,In_1468);
or U241 (N_241,N_187,In_786);
nor U242 (N_242,In_181,In_200);
xor U243 (N_243,In_717,In_1013);
xnor U244 (N_244,In_1305,In_661);
xnor U245 (N_245,N_112,In_307);
or U246 (N_246,In_138,In_851);
nand U247 (N_247,In_226,In_488);
xnor U248 (N_248,In_1476,In_445);
nand U249 (N_249,In_1407,N_123);
or U250 (N_250,In_509,In_1463);
nand U251 (N_251,In_283,In_1226);
nor U252 (N_252,In_61,In_1344);
or U253 (N_253,In_902,In_179);
xnor U254 (N_254,In_414,In_1324);
nor U255 (N_255,N_19,In_99);
xor U256 (N_256,N_21,In_288);
xnor U257 (N_257,In_1143,In_1205);
nor U258 (N_258,In_519,In_105);
nor U259 (N_259,In_683,In_515);
nor U260 (N_260,N_111,In_398);
xor U261 (N_261,In_239,N_13);
xor U262 (N_262,In_632,N_101);
nand U263 (N_263,N_113,N_132);
or U264 (N_264,In_664,In_337);
nor U265 (N_265,In_863,In_127);
and U266 (N_266,In_209,In_1397);
nor U267 (N_267,In_368,In_527);
nand U268 (N_268,N_110,In_722);
or U269 (N_269,In_249,In_1418);
xnor U270 (N_270,In_954,In_1348);
nor U271 (N_271,In_406,In_1055);
and U272 (N_272,In_426,In_732);
nor U273 (N_273,N_8,In_498);
or U274 (N_274,In_202,In_754);
or U275 (N_275,In_1153,In_1263);
xor U276 (N_276,In_1288,In_482);
or U277 (N_277,In_512,In_253);
nor U278 (N_278,In_599,In_1396);
nor U279 (N_279,In_500,In_312);
xnor U280 (N_280,In_268,In_675);
or U281 (N_281,In_944,In_795);
xnor U282 (N_282,In_792,In_252);
nand U283 (N_283,In_748,In_47);
or U284 (N_284,In_995,N_20);
nor U285 (N_285,In_32,In_793);
nand U286 (N_286,In_162,In_1208);
xor U287 (N_287,In_953,In_341);
xnor U288 (N_288,In_434,In_240);
and U289 (N_289,In_932,In_1405);
and U290 (N_290,In_476,In_693);
and U291 (N_291,In_546,In_39);
xor U292 (N_292,In_491,In_1095);
or U293 (N_293,In_1238,N_40);
nor U294 (N_294,N_92,In_913);
xor U295 (N_295,In_1223,N_93);
nor U296 (N_296,In_1123,In_971);
nor U297 (N_297,In_1499,In_233);
nor U298 (N_298,In_604,In_1436);
xor U299 (N_299,In_694,In_1390);
and U300 (N_300,In_1024,In_501);
nor U301 (N_301,In_420,In_1340);
and U302 (N_302,In_1477,In_538);
nand U303 (N_303,In_1410,In_1217);
nor U304 (N_304,In_726,N_3);
nor U305 (N_305,In_1450,In_1080);
or U306 (N_306,In_401,In_1378);
and U307 (N_307,In_416,N_183);
nor U308 (N_308,In_88,In_1118);
nor U309 (N_309,In_684,In_165);
and U310 (N_310,In_1458,In_83);
nor U311 (N_311,In_1259,In_641);
or U312 (N_312,In_686,N_148);
or U313 (N_313,In_287,In_1072);
and U314 (N_314,In_522,N_138);
or U315 (N_315,In_1258,In_577);
nor U316 (N_316,In_679,In_1183);
and U317 (N_317,In_824,In_298);
xnor U318 (N_318,In_293,In_1310);
and U319 (N_319,In_868,In_1023);
or U320 (N_320,N_177,N_41);
or U321 (N_321,In_1432,In_53);
xnor U322 (N_322,In_437,In_150);
and U323 (N_323,In_281,In_964);
nand U324 (N_324,In_627,In_1066);
or U325 (N_325,In_1065,N_186);
xnor U326 (N_326,In_41,In_609);
or U327 (N_327,In_753,In_1047);
nor U328 (N_328,In_1231,In_1424);
xnor U329 (N_329,In_140,In_934);
xnor U330 (N_330,N_24,In_180);
xor U331 (N_331,In_1465,In_356);
xor U332 (N_332,N_77,In_1272);
xor U333 (N_333,In_1277,In_450);
xor U334 (N_334,In_1009,In_153);
nor U335 (N_335,In_156,In_974);
nand U336 (N_336,In_98,In_1480);
and U337 (N_337,N_80,N_6);
or U338 (N_338,In_1475,In_328);
xor U339 (N_339,In_56,In_1164);
xor U340 (N_340,In_872,In_1402);
nor U341 (N_341,In_215,In_407);
nand U342 (N_342,In_1268,In_1412);
nand U343 (N_343,In_386,In_1457);
nand U344 (N_344,In_728,In_390);
xnor U345 (N_345,In_802,In_739);
and U346 (N_346,N_67,In_648);
and U347 (N_347,In_859,In_782);
or U348 (N_348,In_455,N_184);
or U349 (N_349,In_1376,In_291);
xnor U350 (N_350,In_1014,In_898);
and U351 (N_351,N_32,N_71);
nor U352 (N_352,In_1021,In_730);
xnor U353 (N_353,In_813,In_384);
or U354 (N_354,In_6,In_914);
and U355 (N_355,In_687,In_1388);
and U356 (N_356,In_796,In_431);
xnor U357 (N_357,In_850,In_1146);
xnor U358 (N_358,In_908,N_11);
or U359 (N_359,In_1052,In_433);
xnor U360 (N_360,In_79,In_309);
or U361 (N_361,In_861,In_1355);
xnor U362 (N_362,N_10,In_315);
and U363 (N_363,In_696,In_1206);
nand U364 (N_364,In_428,In_1028);
and U365 (N_365,N_134,N_141);
xor U366 (N_366,In_887,In_843);
nor U367 (N_367,In_110,In_526);
xnor U368 (N_368,N_59,In_1415);
xnor U369 (N_369,In_1379,In_875);
nand U370 (N_370,In_1162,In_92);
and U371 (N_371,In_894,In_418);
nor U372 (N_372,In_89,In_834);
xnor U373 (N_373,In_216,In_94);
xor U374 (N_374,N_39,In_524);
xnor U375 (N_375,In_1297,In_508);
nor U376 (N_376,In_1478,In_353);
or U377 (N_377,In_1303,In_206);
or U378 (N_378,In_637,N_192);
xor U379 (N_379,In_483,In_1070);
and U380 (N_380,In_120,N_64);
nor U381 (N_381,In_210,In_531);
nor U382 (N_382,In_1062,N_74);
or U383 (N_383,In_176,In_1245);
and U384 (N_384,In_74,N_73);
or U385 (N_385,N_190,In_1035);
nor U386 (N_386,In_556,In_1498);
nor U387 (N_387,In_1451,In_1420);
nand U388 (N_388,In_1113,In_650);
xnor U389 (N_389,In_779,In_222);
or U390 (N_390,N_14,In_1172);
xor U391 (N_391,In_986,N_78);
xor U392 (N_392,In_346,In_716);
or U393 (N_393,In_102,In_63);
and U394 (N_394,In_1399,In_1054);
nor U395 (N_395,In_1122,In_24);
or U396 (N_396,In_244,In_1321);
or U397 (N_397,In_1169,N_90);
xor U398 (N_398,In_568,In_1100);
nor U399 (N_399,N_76,In_1114);
and U400 (N_400,In_161,In_439);
nor U401 (N_401,N_263,In_741);
and U402 (N_402,In_673,In_147);
nor U403 (N_403,In_1393,In_1489);
nand U404 (N_404,In_635,In_957);
nand U405 (N_405,In_826,N_230);
and U406 (N_406,In_1301,In_1490);
nor U407 (N_407,In_1459,N_384);
or U408 (N_408,N_309,N_43);
nand U409 (N_409,In_991,In_602);
and U410 (N_410,In_231,In_1227);
or U411 (N_411,In_410,In_266);
or U412 (N_412,In_129,In_815);
nor U413 (N_413,In_1187,In_982);
and U414 (N_414,In_554,N_346);
and U415 (N_415,In_460,In_928);
and U416 (N_416,N_338,In_1347);
nand U417 (N_417,In_931,In_833);
nor U418 (N_418,N_288,In_318);
nand U419 (N_419,In_555,In_1425);
nor U420 (N_420,In_62,In_905);
and U421 (N_421,In_536,In_1267);
xnor U422 (N_422,N_205,In_1352);
xnor U423 (N_423,N_70,N_355);
xor U424 (N_424,N_107,In_1050);
or U425 (N_425,In_837,N_109);
or U426 (N_426,N_234,N_335);
and U427 (N_427,In_35,N_203);
nand U428 (N_428,N_293,In_904);
xnor U429 (N_429,In_879,In_446);
or U430 (N_430,N_307,N_389);
and U431 (N_431,In_1374,In_892);
nor U432 (N_432,In_171,In_248);
or U433 (N_433,In_124,In_677);
nor U434 (N_434,In_1192,N_308);
nand U435 (N_435,In_114,In_471);
nand U436 (N_436,In_343,In_182);
nand U437 (N_437,In_1142,N_167);
and U438 (N_438,In_878,In_620);
nor U439 (N_439,In_740,In_989);
nor U440 (N_440,In_457,N_218);
nand U441 (N_441,In_962,In_709);
xnor U442 (N_442,In_361,In_1260);
nand U443 (N_443,N_296,In_1158);
or U444 (N_444,In_618,In_237);
and U445 (N_445,In_311,In_1049);
nor U446 (N_446,N_391,N_398);
and U447 (N_447,N_95,In_475);
nor U448 (N_448,N_314,In_1015);
or U449 (N_449,N_284,In_1179);
nor U450 (N_450,In_583,In_542);
nand U451 (N_451,N_259,In_784);
xnor U452 (N_452,In_375,N_392);
or U453 (N_453,N_311,In_1215);
nor U454 (N_454,In_685,In_374);
xor U455 (N_455,In_422,In_366);
and U456 (N_456,In_3,In_613);
nor U457 (N_457,In_380,N_342);
and U458 (N_458,In_302,In_225);
nor U459 (N_459,N_25,In_284);
nand U460 (N_460,In_757,In_659);
or U461 (N_461,In_1008,N_352);
or U462 (N_462,N_351,In_773);
and U463 (N_463,N_233,In_1124);
nand U464 (N_464,In_322,In_37);
nand U465 (N_465,In_320,In_301);
nand U466 (N_466,N_387,In_653);
nor U467 (N_467,In_1060,In_933);
and U468 (N_468,N_393,In_499);
nor U469 (N_469,In_984,N_162);
and U470 (N_470,In_8,In_1149);
nand U471 (N_471,In_290,In_90);
or U472 (N_472,N_375,In_640);
xnor U473 (N_473,In_647,In_372);
nor U474 (N_474,In_516,In_1276);
nand U475 (N_475,N_165,In_1136);
xor U476 (N_476,In_1228,In_819);
or U477 (N_477,In_1309,N_212);
xnor U478 (N_478,In_525,N_31);
or U479 (N_479,In_185,N_125);
nor U480 (N_480,N_119,N_163);
nand U481 (N_481,N_361,In_227);
or U482 (N_482,In_17,In_1125);
xor U483 (N_483,N_363,In_1200);
nor U484 (N_484,In_1148,In_520);
and U485 (N_485,N_281,In_1431);
and U486 (N_486,In_370,In_735);
xnor U487 (N_487,In_1202,In_489);
xor U488 (N_488,In_900,N_331);
nand U489 (N_489,N_156,In_261);
xnor U490 (N_490,In_949,In_194);
or U491 (N_491,In_1386,In_614);
xor U492 (N_492,N_332,N_173);
nor U493 (N_493,In_1381,In_1389);
nor U494 (N_494,In_1330,N_258);
or U495 (N_495,N_56,N_54);
xnor U496 (N_496,In_5,N_99);
and U497 (N_497,In_1302,In_132);
or U498 (N_498,In_1448,In_1261);
and U499 (N_499,In_321,In_923);
nor U500 (N_500,In_158,N_271);
nand U501 (N_501,In_1364,In_218);
nor U502 (N_502,In_313,In_547);
nor U503 (N_503,N_195,In_173);
nor U504 (N_504,In_7,In_576);
or U505 (N_505,In_1017,In_1285);
xor U506 (N_506,N_143,N_15);
or U507 (N_507,In_1354,In_882);
nor U508 (N_508,In_502,In_421);
and U509 (N_509,N_86,In_119);
or U510 (N_510,N_26,In_324);
or U511 (N_511,N_66,N_390);
nand U512 (N_512,In_1464,N_282);
nor U513 (N_513,In_1129,In_273);
and U514 (N_514,In_775,In_804);
nand U515 (N_515,N_211,In_1025);
xnor U516 (N_516,N_245,N_237);
nor U517 (N_517,N_82,N_137);
and U518 (N_518,N_35,In_534);
and U519 (N_519,In_598,In_1101);
nand U520 (N_520,In_128,In_238);
nand U521 (N_521,In_649,N_179);
and U522 (N_522,In_1199,In_597);
and U523 (N_523,N_320,In_855);
and U524 (N_524,In_544,N_53);
nand U525 (N_525,N_268,In_146);
nand U526 (N_526,In_1093,In_1337);
nand U527 (N_527,In_655,In_354);
nor U528 (N_528,In_190,N_229);
nor U529 (N_529,In_1430,In_269);
xnor U530 (N_530,In_1109,N_322);
or U531 (N_531,N_388,In_941);
and U532 (N_532,N_222,N_27);
xnor U533 (N_533,In_1434,In_811);
nor U534 (N_534,In_692,In_123);
and U535 (N_535,N_96,In_149);
or U536 (N_536,In_1178,In_400);
and U537 (N_537,In_1467,In_807);
xnor U538 (N_538,In_224,N_298);
xor U539 (N_539,In_1111,N_209);
and U540 (N_540,N_171,In_921);
and U541 (N_541,In_282,In_367);
xnor U542 (N_542,N_244,N_185);
nor U543 (N_543,In_690,In_1473);
or U544 (N_544,In_262,In_166);
nor U545 (N_545,N_359,N_373);
xnor U546 (N_546,In_492,In_606);
xor U547 (N_547,In_569,N_232);
nand U548 (N_548,In_1071,N_344);
nor U549 (N_549,N_193,N_240);
xor U550 (N_550,In_814,In_1242);
nand U551 (N_551,In_1239,In_535);
and U552 (N_552,In_749,In_191);
and U553 (N_553,In_885,In_877);
and U554 (N_554,In_23,In_646);
nor U555 (N_555,In_571,In_1034);
nand U556 (N_556,In_1046,In_593);
or U557 (N_557,In_55,In_1204);
and U558 (N_558,N_4,In_762);
and U559 (N_559,N_168,N_150);
and U560 (N_560,In_845,In_1273);
and U561 (N_561,In_76,In_809);
nand U562 (N_562,N_394,In_1064);
or U563 (N_563,In_559,In_330);
or U564 (N_564,In_175,In_485);
nand U565 (N_565,N_358,In_369);
nor U566 (N_566,In_495,In_920);
nor U567 (N_567,N_153,In_736);
or U568 (N_568,N_321,In_125);
xnor U569 (N_569,In_731,In_999);
and U570 (N_570,In_1191,In_1221);
nand U571 (N_571,In_1446,In_155);
nor U572 (N_572,In_698,In_490);
and U573 (N_573,In_1043,In_1189);
nor U574 (N_574,In_223,In_419);
xor U575 (N_575,In_1079,N_362);
xnor U576 (N_576,N_136,In_289);
nor U577 (N_577,N_243,In_994);
or U578 (N_578,In_250,N_140);
nand U579 (N_579,N_155,In_916);
nor U580 (N_580,In_626,In_1286);
nand U581 (N_581,In_980,In_429);
or U582 (N_582,In_387,N_246);
nand U583 (N_583,In_1092,In_172);
xnor U584 (N_584,In_275,In_706);
nand U585 (N_585,N_360,In_397);
and U586 (N_586,In_195,In_12);
or U587 (N_587,In_1120,In_638);
xnor U588 (N_588,In_1359,N_176);
nor U589 (N_589,In_1456,In_211);
nor U590 (N_590,In_183,In_1492);
nor U591 (N_591,In_1482,In_394);
and U592 (N_592,In_1433,N_206);
xor U593 (N_593,N_345,In_18);
or U594 (N_594,In_1119,In_1294);
or U595 (N_595,In_443,N_91);
nand U596 (N_596,N_378,In_1299);
nand U597 (N_597,In_424,In_553);
xor U598 (N_598,In_1403,In_1078);
nor U599 (N_599,In_272,In_344);
xor U600 (N_600,N_439,N_577);
nor U601 (N_601,N_158,N_260);
or U602 (N_602,In_1061,N_459);
nand U603 (N_603,N_563,In_1274);
and U604 (N_604,N_257,N_219);
xnor U605 (N_605,N_175,N_430);
nor U606 (N_606,N_597,N_515);
xnor U607 (N_607,N_562,N_414);
or U608 (N_608,N_483,In_958);
and U609 (N_609,N_417,In_586);
xnor U610 (N_610,In_761,N_540);
nor U611 (N_611,In_1317,In_1195);
nand U612 (N_612,In_1233,N_495);
xnor U613 (N_613,In_644,In_38);
and U614 (N_614,N_371,In_1270);
nand U615 (N_615,N_525,In_1452);
xnor U616 (N_616,N_510,In_363);
xor U617 (N_617,In_329,N_216);
nor U618 (N_618,N_108,N_353);
or U619 (N_619,N_569,N_241);
nor U620 (N_620,N_337,N_255);
and U621 (N_621,N_302,In_1485);
and U622 (N_622,N_469,In_1279);
xnor U623 (N_623,In_304,N_89);
or U624 (N_624,N_274,N_75);
and U625 (N_625,In_1462,In_1222);
and U626 (N_626,N_441,In_1188);
and U627 (N_627,In_818,In_1248);
nand U628 (N_628,In_1361,In_1449);
xor U629 (N_629,N_425,In_617);
and U630 (N_630,In_587,In_1018);
or U631 (N_631,N_450,In_1031);
or U632 (N_632,N_370,N_280);
nor U633 (N_633,In_925,In_376);
or U634 (N_634,In_612,In_456);
nand U635 (N_635,N_572,N_49);
or U636 (N_636,N_406,N_197);
xnor U637 (N_637,In_466,In_1130);
nor U638 (N_638,In_624,N_289);
and U639 (N_639,N_48,In_22);
and U640 (N_640,In_557,N_324);
and U641 (N_641,In_464,In_702);
or U642 (N_642,In_350,N_105);
xnor U643 (N_643,In_1295,In_1298);
and U644 (N_644,N_501,N_316);
nand U645 (N_645,N_253,In_1287);
and U646 (N_646,In_1338,In_1107);
nand U647 (N_647,In_540,In_48);
nand U648 (N_648,N_564,In_1185);
nor U649 (N_649,In_591,In_787);
xnor U650 (N_650,In_336,In_1306);
nor U651 (N_651,In_220,In_30);
nor U652 (N_652,In_715,In_412);
and U653 (N_653,In_67,In_1346);
nor U654 (N_654,In_408,N_416);
nand U655 (N_655,In_1356,N_104);
nor U656 (N_656,N_528,In_871);
and U657 (N_657,N_267,N_506);
and U658 (N_658,N_103,In_510);
and U659 (N_659,In_1323,In_54);
and U660 (N_660,N_382,N_553);
or U661 (N_661,In_212,N_407);
and U662 (N_662,N_539,N_63);
nor U663 (N_663,N_522,N_142);
or U664 (N_664,N_523,In_449);
nor U665 (N_665,In_521,In_1002);
nor U666 (N_666,N_582,N_250);
and U667 (N_667,N_304,In_494);
xor U668 (N_668,N_408,N_536);
xnor U669 (N_669,In_1314,In_899);
nand U670 (N_670,In_280,N_139);
or U671 (N_671,In_791,N_225);
nand U672 (N_672,In_325,In_87);
or U673 (N_673,N_598,N_297);
nand U674 (N_674,In_1225,N_356);
and U675 (N_675,In_13,N_327);
nor U676 (N_676,In_1096,N_559);
nand U677 (N_677,N_117,N_100);
and U678 (N_678,In_947,In_391);
and U679 (N_679,N_499,In_930);
xnor U680 (N_680,N_124,N_299);
xor U681 (N_681,In_639,N_481);
and U682 (N_682,In_1243,In_1455);
nor U683 (N_683,N_535,In_405);
or U684 (N_684,In_897,N_571);
nand U685 (N_685,N_286,In_993);
xor U686 (N_686,N_462,N_383);
nand U687 (N_687,N_575,In_771);
xor U688 (N_688,In_1056,In_968);
nor U689 (N_689,In_481,In_823);
and U690 (N_690,N_468,In_1059);
and U691 (N_691,N_178,In_1357);
or U692 (N_692,In_1216,In_1012);
nor U693 (N_693,In_884,N_512);
and U694 (N_694,N_145,N_482);
xor U695 (N_695,In_1484,In_595);
xor U696 (N_696,In_558,In_247);
nand U697 (N_697,N_130,N_369);
nand U698 (N_698,In_345,N_340);
xor U699 (N_699,In_139,N_42);
or U700 (N_700,N_588,N_410);
or U701 (N_701,In_573,N_488);
nand U702 (N_702,In_184,In_658);
nor U703 (N_703,In_230,N_574);
nand U704 (N_704,In_911,In_578);
nor U705 (N_705,In_1423,In_562);
xnor U706 (N_706,N_88,N_2);
xnor U707 (N_707,In_1173,N_555);
nor U708 (N_708,N_12,In_1413);
xor U709 (N_709,N_433,In_1117);
nor U710 (N_710,In_733,N_599);
nor U711 (N_711,N_264,N_530);
and U712 (N_712,In_777,In_504);
nand U713 (N_713,In_338,N_365);
nand U714 (N_714,In_286,N_194);
nand U715 (N_715,In_204,In_829);
nand U716 (N_716,N_269,N_385);
nor U717 (N_717,In_548,N_266);
nand U718 (N_718,N_305,In_532);
xor U719 (N_719,In_1211,In_660);
or U720 (N_720,N_328,In_1126);
xor U721 (N_721,In_122,N_423);
nand U722 (N_722,N_434,N_326);
xnor U723 (N_723,In_800,N_341);
and U724 (N_724,N_498,N_585);
and U725 (N_725,N_238,In_151);
and U726 (N_726,In_1082,In_952);
xnor U727 (N_727,N_379,N_180);
and U728 (N_728,N_449,N_458);
or U729 (N_729,In_1102,N_457);
or U730 (N_730,In_549,In_178);
xor U731 (N_731,In_699,In_1479);
nand U732 (N_732,N_213,N_83);
xor U733 (N_733,In_1230,In_203);
and U734 (N_734,N_460,N_85);
xor U735 (N_735,In_243,N_586);
and U736 (N_736,In_1201,N_454);
nor U737 (N_737,In_392,In_1246);
nand U738 (N_738,N_166,In_744);
nor U739 (N_739,N_377,N_318);
xor U740 (N_740,N_566,N_347);
nor U741 (N_741,N_448,N_492);
and U742 (N_742,N_144,N_278);
xnor U743 (N_743,N_120,N_30);
nand U744 (N_744,N_405,N_313);
or U745 (N_745,N_556,N_277);
nand U746 (N_746,In_714,In_278);
or U747 (N_747,N_401,N_435);
nor U748 (N_748,N_532,In_890);
xnor U749 (N_749,N_214,N_426);
and U750 (N_750,N_580,In_611);
nand U751 (N_751,In_848,In_1083);
and U752 (N_752,In_1363,N_485);
xor U753 (N_753,In_152,N_518);
and U754 (N_754,In_1110,In_1271);
nor U755 (N_755,N_576,In_373);
and U756 (N_756,N_554,N_228);
xnor U757 (N_757,In_493,In_423);
and U758 (N_758,N_542,N_538);
and U759 (N_759,In_983,In_106);
nor U760 (N_760,In_1445,In_31);
and U761 (N_761,In_513,In_862);
nand U762 (N_762,N_477,In_1026);
nand U763 (N_763,In_1214,N_579);
xor U764 (N_764,In_1358,In_1067);
xnor U765 (N_765,In_358,N_476);
and U766 (N_766,N_224,In_667);
nor U767 (N_767,N_348,In_189);
or U768 (N_768,N_210,N_204);
nor U769 (N_769,N_521,N_7);
or U770 (N_770,In_1224,In_718);
or U771 (N_771,N_1,In_427);
nand U772 (N_772,In_605,N_402);
nor U773 (N_773,N_502,In_135);
nand U774 (N_774,In_1186,In_192);
nand U775 (N_775,N_461,In_308);
and U776 (N_776,N_474,In_1328);
or U777 (N_777,In_1264,In_530);
and U778 (N_778,N_334,In_91);
xor U779 (N_779,In_781,In_628);
nand U780 (N_780,N_189,In_1048);
xnor U781 (N_781,N_79,N_248);
or U782 (N_782,In_1073,In_825);
xnor U783 (N_783,N_46,In_1428);
nor U784 (N_784,N_437,In_838);
or U785 (N_785,In_720,In_1487);
or U786 (N_786,In_411,In_314);
nor U787 (N_787,N_121,N_570);
and U788 (N_788,N_291,N_146);
nor U789 (N_789,N_507,In_966);
nor U790 (N_790,In_25,N_455);
nand U791 (N_791,In_842,N_47);
nor U792 (N_792,In_468,N_596);
xor U793 (N_793,N_590,In_1175);
or U794 (N_794,N_517,N_325);
nand U795 (N_795,N_505,N_61);
and U796 (N_796,In_1141,N_182);
or U797 (N_797,In_1417,In_1105);
or U798 (N_798,In_1077,In_998);
or U799 (N_799,In_1394,In_299);
xnor U800 (N_800,N_673,In_432);
xor U801 (N_801,N_511,N_668);
nand U802 (N_802,N_34,N_789);
xor U803 (N_803,In_566,N_546);
and U804 (N_804,N_428,N_465);
nor U805 (N_805,In_1320,N_122);
or U806 (N_806,N_265,In_821);
or U807 (N_807,In_1442,N_106);
nor U808 (N_808,In_478,In_496);
xor U809 (N_809,In_1380,N_534);
nand U810 (N_810,N_200,N_665);
and U811 (N_811,N_84,N_227);
xor U812 (N_812,N_651,In_463);
nand U813 (N_813,In_1311,N_367);
nor U814 (N_814,N_154,In_112);
or U815 (N_815,N_581,In_1085);
and U816 (N_816,In_131,In_487);
nand U817 (N_817,N_114,N_735);
nand U818 (N_818,N_404,N_589);
nor U819 (N_819,In_159,In_1392);
nor U820 (N_820,In_1098,In_51);
and U821 (N_821,N_223,In_1329);
nor U822 (N_822,N_660,In_1197);
xor U823 (N_823,N_504,In_263);
xnor U824 (N_824,N_757,N_753);
nand U825 (N_825,N_663,N_600);
or U826 (N_826,In_1097,In_1184);
or U827 (N_827,N_226,N_411);
nor U828 (N_828,N_656,In_756);
and U829 (N_829,N_703,N_688);
nand U830 (N_830,In_46,In_846);
xnor U831 (N_831,In_1163,N_202);
xor U832 (N_832,N_629,N_456);
and U833 (N_833,In_607,In_537);
nand U834 (N_834,N_550,N_783);
nor U835 (N_835,In_72,N_72);
and U836 (N_836,N_583,N_690);
or U837 (N_837,N_548,N_544);
nand U838 (N_838,N_300,N_774);
and U839 (N_839,In_292,N_516);
nor U840 (N_840,In_1307,N_565);
xor U841 (N_841,In_260,N_294);
nand U842 (N_842,N_746,N_126);
or U843 (N_843,In_69,In_1176);
and U844 (N_844,In_1325,In_1300);
nor U845 (N_845,N_174,In_68);
nor U846 (N_846,N_712,N_732);
xnor U847 (N_847,In_758,In_371);
nor U848 (N_848,N_683,N_750);
nand U849 (N_849,N_303,N_357);
and U850 (N_850,N_594,In_622);
nor U851 (N_851,N_767,N_709);
nor U852 (N_852,In_1401,N_605);
nand U853 (N_853,In_858,N_609);
nand U854 (N_854,N_743,N_666);
and U855 (N_855,N_677,N_543);
or U856 (N_856,N_771,N_427);
and U857 (N_857,N_491,In_95);
nor U858 (N_858,In_160,N_395);
nor U859 (N_859,In_1236,In_1336);
xnor U860 (N_860,N_742,N_273);
and U861 (N_861,N_283,In_187);
and U862 (N_862,N_275,In_810);
nor U863 (N_863,In_589,N_697);
nand U864 (N_864,In_145,N_601);
nor U865 (N_865,N_669,N_452);
xnor U866 (N_866,N_497,N_235);
or U867 (N_867,N_364,N_751);
xnor U868 (N_868,In_817,N_711);
or U869 (N_869,In_1292,N_329);
xor U870 (N_870,N_679,N_680);
xor U871 (N_871,In_511,In_939);
or U872 (N_872,N_400,N_350);
nand U873 (N_873,N_695,N_533);
nor U874 (N_874,N_323,N_741);
nor U875 (N_875,In_1032,N_722);
xnor U876 (N_876,N_531,In_1159);
and U877 (N_877,In_1063,In_881);
nand U878 (N_878,In_1001,In_271);
and U879 (N_879,In_704,In_19);
xnor U880 (N_880,N_420,N_479);
nor U881 (N_881,N_662,N_418);
nor U882 (N_882,N_713,N_587);
or U883 (N_883,In_425,N_643);
or U884 (N_884,N_397,In_828);
or U885 (N_885,In_364,N_29);
nor U886 (N_886,N_287,In_103);
xor U887 (N_887,N_57,In_621);
xor U888 (N_888,In_86,In_629);
nor U889 (N_889,In_518,N_658);
or U890 (N_890,N_733,In_1004);
nand U891 (N_891,N_290,N_693);
nand U892 (N_892,In_567,N_421);
nand U893 (N_893,N_524,N_493);
nor U894 (N_894,N_526,In_860);
and U895 (N_895,In_1137,In_579);
nor U896 (N_896,In_1387,In_235);
nand U897 (N_897,N_640,In_1406);
xnor U898 (N_898,In_768,N_473);
nand U899 (N_899,N_591,N_698);
or U900 (N_900,N_720,N_793);
or U901 (N_901,N_744,N_619);
nand U902 (N_902,N_686,N_681);
or U903 (N_903,N_780,In_101);
nand U904 (N_904,N_239,N_129);
nand U905 (N_905,N_215,N_568);
xnor U906 (N_906,In_766,In_1198);
nor U907 (N_907,N_573,N_463);
nand U908 (N_908,In_70,In_856);
nor U909 (N_909,N_478,In_1400);
nor U910 (N_910,N_444,N_685);
nand U911 (N_911,N_310,In_1033);
nor U912 (N_912,N_201,N_788);
xor U913 (N_913,In_623,N_451);
or U914 (N_914,In_27,N_261);
nand U915 (N_915,N_315,N_547);
or U916 (N_916,In_448,N_659);
and U917 (N_917,N_545,In_935);
xor U918 (N_918,N_199,N_724);
xnor U919 (N_919,N_170,N_770);
and U920 (N_920,In_551,In_316);
nand U921 (N_921,N_785,N_149);
nand U922 (N_922,N_251,N_217);
nor U923 (N_923,N_5,In_1244);
or U924 (N_924,N_422,N_368);
or U925 (N_925,In_652,N_779);
nor U926 (N_926,N_81,N_721);
and U927 (N_927,N_151,In_473);
or U928 (N_928,N_715,N_595);
nand U929 (N_929,In_601,N_537);
nand U930 (N_930,In_205,In_331);
or U931 (N_931,N_756,N_759);
or U932 (N_932,In_1194,In_1313);
xor U933 (N_933,In_1152,In_1370);
nand U934 (N_934,N_249,N_330);
nor U935 (N_935,In_619,N_648);
xnor U936 (N_936,N_769,In_236);
nand U937 (N_937,N_520,In_1454);
and U938 (N_938,In_979,N_624);
nor U939 (N_939,N_333,In_1170);
or U940 (N_940,N_116,In_305);
nor U941 (N_941,N_611,N_115);
and U942 (N_942,N_292,In_1084);
and U943 (N_943,N_778,In_1384);
or U944 (N_944,N_674,In_561);
or U945 (N_945,In_909,N_424);
xnor U946 (N_946,N_723,N_45);
nand U947 (N_947,In_701,In_1074);
or U948 (N_948,N_412,N_631);
xnor U949 (N_949,N_231,N_22);
nand U950 (N_950,In_874,In_327);
nand U951 (N_951,N_256,N_784);
xnor U952 (N_952,In_1377,N_719);
nand U953 (N_953,N_760,N_621);
and U954 (N_954,In_362,N_729);
or U955 (N_955,N_306,N_295);
nand U956 (N_956,N_749,N_704);
and U957 (N_957,N_519,N_436);
nand U958 (N_958,N_706,N_496);
nor U959 (N_959,N_791,In_1234);
nand U960 (N_960,N_752,N_593);
nand U961 (N_961,N_705,N_646);
or U962 (N_962,N_127,In_378);
nand U963 (N_963,In_1,N_794);
nand U964 (N_964,In_170,In_1251);
nand U965 (N_965,N_440,N_738);
or U966 (N_966,N_650,In_1103);
and U967 (N_967,In_507,N_612);
xor U968 (N_968,N_514,N_317);
xor U969 (N_969,N_561,In_66);
xnor U970 (N_970,In_1293,In_963);
nand U971 (N_971,N_9,In_680);
nor U972 (N_972,N_603,N_781);
or U973 (N_973,N_792,N_247);
nor U974 (N_974,N_795,N_736);
and U975 (N_975,N_467,In_1327);
xor U976 (N_976,In_745,In_1010);
and U977 (N_977,N_500,In_891);
nor U978 (N_978,In_16,In_1213);
nand U979 (N_979,In_1151,N_758);
nor U980 (N_980,In_430,In_929);
or U981 (N_981,In_177,In_666);
nand U982 (N_982,N_687,N_691);
xnor U983 (N_983,N_639,N_678);
nand U984 (N_984,In_234,N_272);
nor U985 (N_985,In_713,N_641);
xor U986 (N_986,N_339,N_409);
or U987 (N_987,N_17,N_374);
xor U988 (N_988,N_312,N_717);
nor U989 (N_989,In_1353,N_730);
xnor U990 (N_990,In_657,N_242);
nor U991 (N_991,In_467,N_443);
xor U992 (N_992,In_303,N_508);
and U993 (N_993,In_563,N_18);
and U994 (N_994,N_160,In_1437);
and U995 (N_995,N_386,In_1371);
xnor U996 (N_996,N_718,In_864);
xnor U997 (N_997,In_310,N_647);
and U998 (N_998,N_714,N_701);
xnor U999 (N_999,In_830,In_747);
and U1000 (N_1000,N_902,N_694);
nor U1001 (N_1001,N_737,N_983);
xor U1002 (N_1002,N_657,In_545);
and U1003 (N_1003,N_807,N_755);
nand U1004 (N_1004,N_846,N_94);
nand U1005 (N_1005,In_1460,N_940);
nand U1006 (N_1006,In_691,In_803);
xnor U1007 (N_1007,N_825,N_911);
or U1008 (N_1008,N_655,N_198);
and U1009 (N_1009,N_748,N_159);
nor U1010 (N_1010,N_38,N_637);
or U1011 (N_1011,N_917,N_836);
xor U1012 (N_1012,N_776,In_743);
nor U1013 (N_1013,N_944,N_616);
or U1014 (N_1014,In_506,N_128);
xor U1015 (N_1015,N_815,N_986);
xnor U1016 (N_1016,N_614,N_480);
nand U1017 (N_1017,N_954,N_880);
nand U1018 (N_1018,N_622,N_606);
and U1019 (N_1019,N_860,In_1203);
xnor U1020 (N_1020,N_811,N_961);
or U1021 (N_1021,In_965,In_700);
nor U1022 (N_1022,N_16,N_503);
nand U1023 (N_1023,In_840,N_821);
xnor U1024 (N_1024,N_897,N_904);
or U1025 (N_1025,N_895,In_44);
nor U1026 (N_1026,N_898,N_877);
or U1027 (N_1027,N_208,N_726);
and U1028 (N_1028,N_684,N_798);
xor U1029 (N_1029,In_257,N_819);
and U1030 (N_1030,N_912,In_402);
nand U1031 (N_1031,N_931,N_908);
or U1032 (N_1032,In_805,N_978);
nand U1033 (N_1033,In_503,N_464);
and U1034 (N_1034,In_988,N_319);
and U1035 (N_1035,N_527,N_892);
nand U1036 (N_1036,N_875,In_852);
nor U1037 (N_1037,N_915,N_955);
xor U1038 (N_1038,N_907,In_581);
and U1039 (N_1039,N_489,N_838);
and U1040 (N_1040,In_853,N_252);
and U1041 (N_1041,N_884,In_395);
and U1042 (N_1042,N_745,In_71);
nor U1043 (N_1043,In_1040,N_812);
and U1044 (N_1044,In_906,N_731);
or U1045 (N_1045,N_301,In_1315);
or U1046 (N_1046,N_992,N_800);
nand U1047 (N_1047,N_276,N_381);
xnor U1048 (N_1048,In_1408,N_982);
nor U1049 (N_1049,N_989,N_632);
nor U1050 (N_1050,N_560,N_747);
nand U1051 (N_1051,N_529,N_484);
and U1052 (N_1052,In_1075,N_849);
or U1053 (N_1053,N_956,N_859);
xor U1054 (N_1054,N_945,In_174);
xnor U1055 (N_1055,In_1304,In_1466);
or U1056 (N_1056,In_462,N_896);
xnor U1057 (N_1057,N_843,N_823);
xor U1058 (N_1058,N_671,N_627);
xnor U1059 (N_1059,N_782,N_920);
xor U1060 (N_1060,N_835,In_1140);
nor U1061 (N_1061,In_393,In_82);
nand U1062 (N_1062,N_557,N_664);
and U1063 (N_1063,N_864,N_354);
and U1064 (N_1064,N_396,N_848);
xnor U1065 (N_1065,In_300,In_148);
nand U1066 (N_1066,N_879,N_399);
nor U1067 (N_1067,N_645,N_809);
xor U1068 (N_1068,N_376,N_682);
and U1069 (N_1069,N_831,N_936);
and U1070 (N_1070,N_445,In_827);
or U1071 (N_1071,N_762,N_689);
and U1072 (N_1072,In_1135,N_935);
nor U1073 (N_1073,N_818,N_164);
or U1074 (N_1074,N_949,N_630);
nand U1075 (N_1075,N_558,N_938);
xnor U1076 (N_1076,N_953,N_620);
xor U1077 (N_1077,In_1177,N_644);
nor U1078 (N_1078,In_9,In_738);
and U1079 (N_1079,N_965,N_810);
nor U1080 (N_1080,In_306,In_188);
xor U1081 (N_1081,N_820,In_750);
xnor U1082 (N_1082,N_513,N_487);
and U1083 (N_1083,N_775,N_710);
or U1084 (N_1084,N_628,N_708);
xor U1085 (N_1085,N_584,N_885);
or U1086 (N_1086,N_262,In_196);
nand U1087 (N_1087,N_891,N_36);
xor U1088 (N_1088,In_389,N_602);
or U1089 (N_1089,N_806,In_889);
and U1090 (N_1090,N_943,N_592);
or U1091 (N_1091,N_899,N_963);
nor U1092 (N_1092,N_692,N_672);
nor U1093 (N_1093,In_1318,N_957);
nand U1094 (N_1094,N_830,N_135);
xor U1095 (N_1095,N_967,N_893);
nand U1096 (N_1096,N_952,N_754);
and U1097 (N_1097,N_869,N_649);
and U1098 (N_1098,In_1331,In_1255);
nor U1099 (N_1099,N_841,In_277);
nand U1100 (N_1100,N_799,N_764);
xor U1101 (N_1101,N_901,In_710);
or U1102 (N_1102,N_889,In_461);
nand U1103 (N_1103,N_635,N_699);
nand U1104 (N_1104,N_850,N_549);
and U1105 (N_1105,N_980,In_1115);
nand U1106 (N_1106,N_932,N_826);
nor U1107 (N_1107,N_834,N_118);
and U1108 (N_1108,N_962,N_62);
nand U1109 (N_1109,N_60,N_471);
nor U1110 (N_1110,N_773,N_28);
and U1111 (N_1111,N_490,N_551);
nand U1112 (N_1112,In_1196,N_623);
nor U1113 (N_1113,N_801,N_857);
nand U1114 (N_1114,N_802,N_852);
xor U1115 (N_1115,In_695,N_937);
and U1116 (N_1116,N_790,N_862);
xor U1117 (N_1117,In_229,N_991);
xnor U1118 (N_1118,N_52,N_886);
and U1119 (N_1119,In_1154,N_867);
and U1120 (N_1120,N_960,N_403);
xor U1121 (N_1121,N_863,N_270);
nor U1122 (N_1122,N_727,In_100);
nor U1123 (N_1123,In_359,N_734);
nand U1124 (N_1124,N_842,In_969);
xor U1125 (N_1125,N_786,N_822);
or U1126 (N_1126,N_419,N_926);
nand U1127 (N_1127,In_528,N_909);
or U1128 (N_1128,N_856,N_851);
and U1129 (N_1129,N_813,N_988);
and U1130 (N_1130,N_285,N_974);
and U1131 (N_1131,N_927,In_133);
nand U1132 (N_1132,N_765,In_136);
and U1133 (N_1133,In_274,N_903);
nand U1134 (N_1134,In_1365,N_948);
xor U1135 (N_1135,In_242,N_236);
nor U1136 (N_1136,N_372,N_336);
nand U1137 (N_1137,N_509,N_578);
nand U1138 (N_1138,N_924,N_725);
xor U1139 (N_1139,N_876,N_868);
and U1140 (N_1140,N_102,In_812);
nor U1141 (N_1141,N_796,N_763);
nand U1142 (N_1142,N_971,In_270);
xor U1143 (N_1143,N_740,In_1156);
nor U1144 (N_1144,In_1044,N_874);
nand U1145 (N_1145,N_827,In_1108);
nor U1146 (N_1146,N_828,N_607);
and U1147 (N_1147,N_872,N_429);
xnor U1148 (N_1148,In_616,N_829);
nand U1149 (N_1149,N_941,N_987);
nor U1150 (N_1150,N_919,N_968);
or U1151 (N_1151,N_279,N_447);
or U1152 (N_1152,In_1368,N_922);
nand U1153 (N_1153,In_910,In_960);
or U1154 (N_1154,In_241,N_777);
and U1155 (N_1155,N_415,In_608);
and U1156 (N_1156,N_958,N_675);
and U1157 (N_1157,N_739,N_934);
or U1158 (N_1158,N_870,N_906);
or U1159 (N_1159,N_855,In_592);
or U1160 (N_1160,N_928,N_343);
xnor U1161 (N_1161,In_85,N_832);
xnor U1162 (N_1162,N_787,In_116);
and U1163 (N_1163,N_716,N_636);
nor U1164 (N_1164,In_901,N_220);
and U1165 (N_1165,N_68,N_652);
nor U1166 (N_1166,N_466,N_707);
nand U1167 (N_1167,N_633,N_858);
or U1168 (N_1168,N_900,N_970);
and U1169 (N_1169,N_905,N_973);
and U1170 (N_1170,In_1171,N_916);
nor U1171 (N_1171,In_1382,N_925);
and U1172 (N_1172,N_608,N_552);
nor U1173 (N_1173,N_998,N_634);
or U1174 (N_1174,N_861,N_702);
nor U1175 (N_1175,N_921,N_939);
nand U1176 (N_1176,In_80,N_349);
nand U1177 (N_1177,N_999,N_181);
nor U1178 (N_1178,In_888,N_881);
and U1179 (N_1179,N_833,N_814);
nor U1180 (N_1180,In_972,N_44);
or U1181 (N_1181,N_761,N_667);
nand U1182 (N_1182,N_979,N_993);
nand U1183 (N_1183,N_413,In_379);
or U1184 (N_1184,N_626,N_969);
nor U1185 (N_1185,N_910,N_972);
or U1186 (N_1186,N_191,N_996);
and U1187 (N_1187,N_933,N_431);
nor U1188 (N_1188,In_582,In_822);
and U1189 (N_1189,In_541,N_914);
and U1190 (N_1190,N_804,N_610);
nand U1191 (N_1191,N_625,N_883);
xor U1192 (N_1192,N_472,N_494);
nor U1193 (N_1193,N_638,N_853);
xnor U1194 (N_1194,N_475,N_816);
nand U1195 (N_1195,N_50,N_661);
xnor U1196 (N_1196,In_199,N_380);
xnor U1197 (N_1197,N_37,N_470);
nor U1198 (N_1198,N_975,In_264);
or U1199 (N_1199,N_486,N_844);
xnor U1200 (N_1200,N_1022,N_1118);
and U1201 (N_1201,N_1035,N_1045);
nand U1202 (N_1202,N_1128,N_990);
or U1203 (N_1203,N_1195,N_541);
nor U1204 (N_1204,N_847,N_1153);
nor U1205 (N_1205,N_995,N_1115);
nand U1206 (N_1206,In_474,N_966);
and U1207 (N_1207,N_1159,N_997);
nor U1208 (N_1208,N_1061,N_878);
nor U1209 (N_1209,N_1091,N_1049);
nor U1210 (N_1210,N_1079,N_1154);
and U1211 (N_1211,N_613,N_959);
xor U1212 (N_1212,N_1139,N_1143);
and U1213 (N_1213,N_1144,N_1105);
xnor U1214 (N_1214,N_839,N_604);
nor U1215 (N_1215,N_1066,N_653);
and U1216 (N_1216,N_1082,N_1103);
nand U1217 (N_1217,N_1181,N_1165);
or U1218 (N_1218,N_1106,N_1059);
nand U1219 (N_1219,N_803,In_169);
or U1220 (N_1220,N_1132,N_1000);
and U1221 (N_1221,N_1039,N_1029);
and U1222 (N_1222,In_585,In_396);
xnor U1223 (N_1223,N_976,In_854);
nand U1224 (N_1224,N_1112,N_1004);
or U1225 (N_1225,N_1080,N_985);
nand U1226 (N_1226,N_918,N_1116);
xor U1227 (N_1227,N_1053,N_1193);
nand U1228 (N_1228,N_1160,N_929);
nor U1229 (N_1229,N_840,N_1094);
or U1230 (N_1230,N_1099,N_1040);
nand U1231 (N_1231,N_1167,N_615);
nand U1232 (N_1232,N_984,N_964);
and U1233 (N_1233,N_1025,N_654);
nand U1234 (N_1234,N_1177,N_1093);
and U1235 (N_1235,N_676,In_926);
xnor U1236 (N_1236,N_1164,N_1090);
or U1237 (N_1237,In_615,N_1068);
nor U1238 (N_1238,N_1083,N_1135);
nor U1239 (N_1239,N_1015,In_213);
nand U1240 (N_1240,N_1155,N_1033);
and U1241 (N_1241,N_1121,N_1174);
xnor U1242 (N_1242,In_1419,N_1011);
or U1243 (N_1243,N_1183,N_642);
and U1244 (N_1244,In_355,N_1109);
xor U1245 (N_1245,N_432,In_857);
nand U1246 (N_1246,N_446,N_1170);
nand U1247 (N_1247,N_1130,N_1017);
xor U1248 (N_1248,N_1085,N_1166);
and U1249 (N_1249,N_1096,N_1137);
and U1250 (N_1250,In_961,N_617);
and U1251 (N_1251,N_1161,N_1072);
xor U1252 (N_1252,N_1032,N_1189);
nand U1253 (N_1253,N_1036,N_1048);
and U1254 (N_1254,N_1101,N_567);
or U1255 (N_1255,N_1037,N_1089);
xnor U1256 (N_1256,N_1184,N_1113);
xnor U1257 (N_1257,N_172,N_1138);
or U1258 (N_1258,N_1041,N_1162);
nor U1259 (N_1259,N_51,N_1108);
nand U1260 (N_1260,N_442,N_1020);
and U1261 (N_1261,N_1010,N_1075);
nor U1262 (N_1262,N_1050,N_887);
and U1263 (N_1263,N_1142,In_1383);
and U1264 (N_1264,N_1084,N_873);
nand U1265 (N_1265,N_1176,N_1058);
and U1266 (N_1266,N_1038,In_776);
nor U1267 (N_1267,N_950,N_696);
or U1268 (N_1268,N_1009,N_1067);
nor U1269 (N_1269,N_1057,N_1188);
or U1270 (N_1270,N_1088,N_1127);
and U1271 (N_1271,N_1179,N_871);
nor U1272 (N_1272,N_1071,N_1007);
or U1273 (N_1273,N_1064,N_670);
nand U1274 (N_1274,N_981,N_1131);
nand U1275 (N_1275,N_882,N_1187);
and U1276 (N_1276,N_1026,N_1182);
xor U1277 (N_1277,N_1173,N_1074);
nor U1278 (N_1278,In_1367,N_1086);
nor U1279 (N_1279,In_1351,N_1180);
or U1280 (N_1280,N_131,N_942);
and U1281 (N_1281,N_1063,N_865);
nand U1282 (N_1282,In_707,N_1190);
and U1283 (N_1283,N_1097,N_1123);
nor U1284 (N_1284,N_1002,N_1056);
xnor U1285 (N_1285,N_1046,N_1133);
or U1286 (N_1286,N_1042,N_453);
xnor U1287 (N_1287,N_837,N_1051);
nand U1288 (N_1288,N_1196,N_854);
nand U1289 (N_1289,N_1065,N_1087);
nand U1290 (N_1290,N_1111,N_1027);
xnor U1291 (N_1291,N_1052,N_1023);
xnor U1292 (N_1292,N_894,N_1043);
and U1293 (N_1293,N_923,N_947);
nor U1294 (N_1294,N_817,N_1003);
nor U1295 (N_1295,N_1006,N_1134);
nand U1296 (N_1296,N_1124,N_1077);
or U1297 (N_1297,N_1014,N_797);
and U1298 (N_1298,N_1069,N_1194);
or U1299 (N_1299,N_1070,N_1157);
nor U1300 (N_1300,N_1152,N_1119);
nor U1301 (N_1301,N_1150,N_1034);
or U1302 (N_1302,In_219,N_1019);
and U1303 (N_1303,In_580,N_1001);
xnor U1304 (N_1304,N_254,N_1031);
nand U1305 (N_1305,N_1055,N_888);
nand U1306 (N_1306,N_1044,N_1178);
nand U1307 (N_1307,N_1125,N_207);
and U1308 (N_1308,In_770,N_1005);
nor U1309 (N_1309,N_913,N_1024);
nor U1310 (N_1310,N_1054,N_1148);
nor U1311 (N_1311,N_1198,N_1172);
xnor U1312 (N_1312,N_1102,N_1192);
xor U1313 (N_1313,N_728,N_1136);
nor U1314 (N_1314,N_890,N_994);
nor U1315 (N_1315,N_1129,N_1141);
xor U1316 (N_1316,N_1140,N_366);
nor U1317 (N_1317,N_438,N_1169);
xor U1318 (N_1318,N_1199,N_1117);
xnor U1319 (N_1319,N_805,N_1122);
nand U1320 (N_1320,N_1171,N_930);
nor U1321 (N_1321,N_1158,N_1047);
nand U1322 (N_1322,N_700,N_1012);
nand U1323 (N_1323,N_1107,N_1197);
nor U1324 (N_1324,N_1126,N_1145);
or U1325 (N_1325,N_98,N_1191);
nor U1326 (N_1326,N_1146,N_977);
xnor U1327 (N_1327,N_1081,N_1156);
xnor U1328 (N_1328,N_1013,N_1163);
nor U1329 (N_1329,N_824,N_1120);
xor U1330 (N_1330,N_1062,N_1110);
or U1331 (N_1331,N_1008,In_1088);
or U1332 (N_1332,N_618,N_1185);
nor U1333 (N_1333,N_1073,N_766);
nor U1334 (N_1334,N_196,N_1114);
nand U1335 (N_1335,N_1030,N_1147);
and U1336 (N_1336,N_1060,N_1151);
or U1337 (N_1337,N_1016,N_866);
and U1338 (N_1338,N_1100,N_772);
nor U1339 (N_1339,N_1104,In_1280);
and U1340 (N_1340,N_1168,N_1078);
nand U1341 (N_1341,N_1021,N_1098);
nor U1342 (N_1342,N_221,N_1186);
nor U1343 (N_1343,N_1095,N_845);
nand U1344 (N_1344,N_1175,N_1149);
or U1345 (N_1345,N_768,N_808);
and U1346 (N_1346,N_1076,In_265);
and U1347 (N_1347,N_951,In_1481);
nor U1348 (N_1348,N_1092,N_946);
or U1349 (N_1349,N_1018,N_1028);
xor U1350 (N_1350,N_1027,N_1186);
nor U1351 (N_1351,N_772,N_959);
xor U1352 (N_1352,N_1119,N_1109);
xnor U1353 (N_1353,N_1138,N_1014);
nand U1354 (N_1354,N_959,N_797);
or U1355 (N_1355,N_1003,N_615);
xor U1356 (N_1356,N_866,In_219);
and U1357 (N_1357,N_1025,N_1035);
nor U1358 (N_1358,N_1145,In_770);
xnor U1359 (N_1359,In_213,N_1128);
nor U1360 (N_1360,N_1172,N_1133);
nor U1361 (N_1361,N_1067,N_1182);
nor U1362 (N_1362,N_1174,N_1126);
nand U1363 (N_1363,In_585,N_1181);
nand U1364 (N_1364,N_1160,N_1074);
nor U1365 (N_1365,N_772,N_1053);
nor U1366 (N_1366,N_913,N_1196);
xor U1367 (N_1367,N_1177,N_1143);
and U1368 (N_1368,N_1192,N_1127);
or U1369 (N_1369,In_707,N_1001);
or U1370 (N_1370,N_1026,N_446);
or U1371 (N_1371,N_1009,N_997);
nand U1372 (N_1372,N_1188,In_585);
nor U1373 (N_1373,N_977,N_1186);
nor U1374 (N_1374,N_1140,N_1051);
xor U1375 (N_1375,N_1199,N_1001);
nand U1376 (N_1376,N_985,In_615);
nand U1377 (N_1377,N_803,N_1117);
nor U1378 (N_1378,N_1095,N_1182);
and U1379 (N_1379,N_1042,N_1158);
xor U1380 (N_1380,In_776,N_1172);
nor U1381 (N_1381,N_670,N_1190);
nor U1382 (N_1382,N_1188,N_1037);
nand U1383 (N_1383,N_1049,N_1034);
xor U1384 (N_1384,N_642,N_207);
nand U1385 (N_1385,N_1110,N_1016);
nand U1386 (N_1386,N_990,N_772);
nor U1387 (N_1387,N_1153,N_1121);
xnor U1388 (N_1388,N_1168,N_642);
and U1389 (N_1389,N_1142,In_1419);
or U1390 (N_1390,N_1106,N_1144);
xor U1391 (N_1391,N_1045,N_1160);
nor U1392 (N_1392,N_1105,N_604);
nor U1393 (N_1393,N_1037,N_1087);
or U1394 (N_1394,In_857,N_1194);
nor U1395 (N_1395,N_1035,N_1063);
nor U1396 (N_1396,N_888,N_1126);
and U1397 (N_1397,N_1049,N_1009);
nand U1398 (N_1398,In_355,N_1015);
and U1399 (N_1399,In_1351,N_1063);
or U1400 (N_1400,N_1359,N_1376);
nand U1401 (N_1401,N_1355,N_1201);
or U1402 (N_1402,N_1260,N_1219);
xor U1403 (N_1403,N_1313,N_1309);
nand U1404 (N_1404,N_1258,N_1269);
xor U1405 (N_1405,N_1364,N_1378);
nor U1406 (N_1406,N_1329,N_1333);
nor U1407 (N_1407,N_1272,N_1291);
xor U1408 (N_1408,N_1342,N_1251);
nand U1409 (N_1409,N_1263,N_1394);
and U1410 (N_1410,N_1233,N_1338);
nand U1411 (N_1411,N_1348,N_1298);
nand U1412 (N_1412,N_1387,N_1239);
and U1413 (N_1413,N_1398,N_1202);
nor U1414 (N_1414,N_1217,N_1312);
and U1415 (N_1415,N_1216,N_1255);
xor U1416 (N_1416,N_1353,N_1344);
or U1417 (N_1417,N_1224,N_1271);
and U1418 (N_1418,N_1274,N_1307);
or U1419 (N_1419,N_1351,N_1372);
and U1420 (N_1420,N_1243,N_1315);
nor U1421 (N_1421,N_1211,N_1297);
xnor U1422 (N_1422,N_1221,N_1273);
nand U1423 (N_1423,N_1393,N_1371);
and U1424 (N_1424,N_1350,N_1324);
and U1425 (N_1425,N_1292,N_1318);
or U1426 (N_1426,N_1383,N_1392);
nor U1427 (N_1427,N_1290,N_1389);
xnor U1428 (N_1428,N_1354,N_1331);
or U1429 (N_1429,N_1214,N_1302);
and U1430 (N_1430,N_1241,N_1294);
nor U1431 (N_1431,N_1340,N_1288);
nand U1432 (N_1432,N_1397,N_1215);
and U1433 (N_1433,N_1254,N_1218);
and U1434 (N_1434,N_1319,N_1235);
xor U1435 (N_1435,N_1304,N_1327);
or U1436 (N_1436,N_1232,N_1287);
xor U1437 (N_1437,N_1311,N_1210);
and U1438 (N_1438,N_1332,N_1231);
nor U1439 (N_1439,N_1270,N_1391);
and U1440 (N_1440,N_1306,N_1384);
nand U1441 (N_1441,N_1339,N_1369);
nor U1442 (N_1442,N_1268,N_1276);
xor U1443 (N_1443,N_1365,N_1301);
and U1444 (N_1444,N_1346,N_1213);
nand U1445 (N_1445,N_1358,N_1293);
and U1446 (N_1446,N_1300,N_1317);
nor U1447 (N_1447,N_1362,N_1222);
nand U1448 (N_1448,N_1328,N_1379);
and U1449 (N_1449,N_1283,N_1382);
and U1450 (N_1450,N_1308,N_1375);
nor U1451 (N_1451,N_1203,N_1226);
nor U1452 (N_1452,N_1284,N_1252);
nand U1453 (N_1453,N_1396,N_1282);
xor U1454 (N_1454,N_1275,N_1316);
nand U1455 (N_1455,N_1386,N_1228);
and U1456 (N_1456,N_1223,N_1326);
or U1457 (N_1457,N_1295,N_1277);
and U1458 (N_1458,N_1380,N_1325);
or U1459 (N_1459,N_1245,N_1381);
xor U1460 (N_1460,N_1238,N_1370);
nand U1461 (N_1461,N_1341,N_1368);
or U1462 (N_1462,N_1209,N_1390);
nor U1463 (N_1463,N_1212,N_1259);
xor U1464 (N_1464,N_1229,N_1261);
or U1465 (N_1465,N_1330,N_1336);
nor U1466 (N_1466,N_1278,N_1227);
and U1467 (N_1467,N_1249,N_1385);
nand U1468 (N_1468,N_1356,N_1321);
or U1469 (N_1469,N_1247,N_1246);
nor U1470 (N_1470,N_1337,N_1314);
nor U1471 (N_1471,N_1237,N_1205);
nand U1472 (N_1472,N_1399,N_1347);
and U1473 (N_1473,N_1323,N_1320);
and U1474 (N_1474,N_1256,N_1257);
xnor U1475 (N_1475,N_1335,N_1225);
nor U1476 (N_1476,N_1296,N_1250);
nand U1477 (N_1477,N_1244,N_1334);
or U1478 (N_1478,N_1281,N_1366);
and U1479 (N_1479,N_1377,N_1299);
nor U1480 (N_1480,N_1289,N_1264);
nand U1481 (N_1481,N_1208,N_1285);
nor U1482 (N_1482,N_1262,N_1200);
nor U1483 (N_1483,N_1265,N_1374);
and U1484 (N_1484,N_1310,N_1395);
nand U1485 (N_1485,N_1267,N_1220);
or U1486 (N_1486,N_1253,N_1204);
or U1487 (N_1487,N_1361,N_1279);
xnor U1488 (N_1488,N_1236,N_1322);
xor U1489 (N_1489,N_1242,N_1360);
nand U1490 (N_1490,N_1343,N_1207);
or U1491 (N_1491,N_1352,N_1349);
nor U1492 (N_1492,N_1367,N_1373);
and U1493 (N_1493,N_1303,N_1357);
or U1494 (N_1494,N_1206,N_1388);
nand U1495 (N_1495,N_1234,N_1345);
or U1496 (N_1496,N_1230,N_1286);
and U1497 (N_1497,N_1266,N_1240);
and U1498 (N_1498,N_1248,N_1363);
xnor U1499 (N_1499,N_1280,N_1305);
xnor U1500 (N_1500,N_1316,N_1267);
nor U1501 (N_1501,N_1272,N_1360);
and U1502 (N_1502,N_1366,N_1369);
nand U1503 (N_1503,N_1308,N_1338);
or U1504 (N_1504,N_1387,N_1224);
nand U1505 (N_1505,N_1317,N_1201);
xnor U1506 (N_1506,N_1209,N_1284);
xnor U1507 (N_1507,N_1238,N_1362);
xor U1508 (N_1508,N_1262,N_1224);
and U1509 (N_1509,N_1329,N_1334);
or U1510 (N_1510,N_1299,N_1239);
nand U1511 (N_1511,N_1319,N_1257);
nand U1512 (N_1512,N_1249,N_1383);
nor U1513 (N_1513,N_1270,N_1243);
or U1514 (N_1514,N_1376,N_1209);
and U1515 (N_1515,N_1243,N_1368);
nand U1516 (N_1516,N_1284,N_1260);
xor U1517 (N_1517,N_1232,N_1220);
or U1518 (N_1518,N_1381,N_1362);
and U1519 (N_1519,N_1209,N_1319);
or U1520 (N_1520,N_1376,N_1374);
and U1521 (N_1521,N_1285,N_1246);
xor U1522 (N_1522,N_1388,N_1243);
nand U1523 (N_1523,N_1268,N_1257);
and U1524 (N_1524,N_1277,N_1346);
xor U1525 (N_1525,N_1389,N_1227);
or U1526 (N_1526,N_1360,N_1243);
xnor U1527 (N_1527,N_1228,N_1265);
or U1528 (N_1528,N_1272,N_1284);
nand U1529 (N_1529,N_1288,N_1232);
nand U1530 (N_1530,N_1339,N_1210);
nor U1531 (N_1531,N_1385,N_1307);
xnor U1532 (N_1532,N_1370,N_1270);
nand U1533 (N_1533,N_1325,N_1303);
xor U1534 (N_1534,N_1349,N_1357);
nand U1535 (N_1535,N_1319,N_1337);
or U1536 (N_1536,N_1312,N_1386);
and U1537 (N_1537,N_1339,N_1333);
nand U1538 (N_1538,N_1205,N_1386);
nand U1539 (N_1539,N_1272,N_1399);
and U1540 (N_1540,N_1300,N_1251);
nand U1541 (N_1541,N_1393,N_1367);
nand U1542 (N_1542,N_1342,N_1203);
xor U1543 (N_1543,N_1343,N_1359);
nand U1544 (N_1544,N_1386,N_1350);
xnor U1545 (N_1545,N_1200,N_1380);
and U1546 (N_1546,N_1308,N_1290);
nor U1547 (N_1547,N_1307,N_1330);
and U1548 (N_1548,N_1372,N_1276);
xor U1549 (N_1549,N_1206,N_1322);
xnor U1550 (N_1550,N_1321,N_1319);
and U1551 (N_1551,N_1260,N_1279);
and U1552 (N_1552,N_1218,N_1367);
xor U1553 (N_1553,N_1347,N_1267);
and U1554 (N_1554,N_1359,N_1349);
nor U1555 (N_1555,N_1377,N_1278);
nor U1556 (N_1556,N_1324,N_1371);
xor U1557 (N_1557,N_1255,N_1393);
or U1558 (N_1558,N_1348,N_1211);
nand U1559 (N_1559,N_1242,N_1358);
nand U1560 (N_1560,N_1354,N_1378);
nor U1561 (N_1561,N_1391,N_1355);
xor U1562 (N_1562,N_1344,N_1375);
and U1563 (N_1563,N_1339,N_1292);
nor U1564 (N_1564,N_1323,N_1243);
and U1565 (N_1565,N_1238,N_1357);
nand U1566 (N_1566,N_1223,N_1273);
or U1567 (N_1567,N_1299,N_1293);
nor U1568 (N_1568,N_1351,N_1276);
and U1569 (N_1569,N_1252,N_1376);
xnor U1570 (N_1570,N_1284,N_1202);
nand U1571 (N_1571,N_1280,N_1263);
nand U1572 (N_1572,N_1347,N_1222);
nand U1573 (N_1573,N_1371,N_1299);
nor U1574 (N_1574,N_1203,N_1231);
nor U1575 (N_1575,N_1279,N_1230);
or U1576 (N_1576,N_1241,N_1380);
nor U1577 (N_1577,N_1220,N_1323);
xnor U1578 (N_1578,N_1263,N_1338);
xnor U1579 (N_1579,N_1237,N_1307);
and U1580 (N_1580,N_1301,N_1352);
or U1581 (N_1581,N_1386,N_1353);
and U1582 (N_1582,N_1340,N_1350);
nand U1583 (N_1583,N_1369,N_1378);
nor U1584 (N_1584,N_1387,N_1256);
and U1585 (N_1585,N_1341,N_1311);
or U1586 (N_1586,N_1202,N_1311);
or U1587 (N_1587,N_1227,N_1302);
nor U1588 (N_1588,N_1390,N_1318);
or U1589 (N_1589,N_1364,N_1220);
xnor U1590 (N_1590,N_1202,N_1205);
nor U1591 (N_1591,N_1352,N_1345);
nor U1592 (N_1592,N_1323,N_1366);
and U1593 (N_1593,N_1349,N_1362);
nor U1594 (N_1594,N_1311,N_1357);
and U1595 (N_1595,N_1204,N_1377);
and U1596 (N_1596,N_1289,N_1387);
and U1597 (N_1597,N_1349,N_1266);
xnor U1598 (N_1598,N_1278,N_1249);
nand U1599 (N_1599,N_1297,N_1368);
and U1600 (N_1600,N_1565,N_1599);
nor U1601 (N_1601,N_1534,N_1552);
xnor U1602 (N_1602,N_1598,N_1563);
nor U1603 (N_1603,N_1463,N_1462);
nor U1604 (N_1604,N_1451,N_1583);
nor U1605 (N_1605,N_1477,N_1512);
or U1606 (N_1606,N_1544,N_1433);
nor U1607 (N_1607,N_1525,N_1516);
xnor U1608 (N_1608,N_1472,N_1495);
nand U1609 (N_1609,N_1474,N_1415);
xnor U1610 (N_1610,N_1483,N_1481);
xnor U1611 (N_1611,N_1427,N_1437);
xnor U1612 (N_1612,N_1569,N_1586);
xor U1613 (N_1613,N_1471,N_1584);
and U1614 (N_1614,N_1424,N_1581);
or U1615 (N_1615,N_1409,N_1504);
xor U1616 (N_1616,N_1466,N_1553);
nor U1617 (N_1617,N_1497,N_1492);
xnor U1618 (N_1618,N_1549,N_1476);
or U1619 (N_1619,N_1468,N_1571);
and U1620 (N_1620,N_1590,N_1426);
xnor U1621 (N_1621,N_1543,N_1442);
nand U1622 (N_1622,N_1489,N_1425);
nor U1623 (N_1623,N_1523,N_1530);
xor U1624 (N_1624,N_1414,N_1555);
or U1625 (N_1625,N_1488,N_1486);
nand U1626 (N_1626,N_1554,N_1502);
xor U1627 (N_1627,N_1545,N_1496);
or U1628 (N_1628,N_1566,N_1469);
or U1629 (N_1629,N_1473,N_1582);
or U1630 (N_1630,N_1467,N_1505);
or U1631 (N_1631,N_1550,N_1561);
nor U1632 (N_1632,N_1570,N_1413);
or U1633 (N_1633,N_1528,N_1490);
and U1634 (N_1634,N_1482,N_1403);
nor U1635 (N_1635,N_1411,N_1568);
nand U1636 (N_1636,N_1589,N_1461);
and U1637 (N_1637,N_1567,N_1597);
or U1638 (N_1638,N_1480,N_1465);
nor U1639 (N_1639,N_1520,N_1591);
xnor U1640 (N_1640,N_1416,N_1594);
nand U1641 (N_1641,N_1576,N_1455);
xor U1642 (N_1642,N_1539,N_1499);
or U1643 (N_1643,N_1408,N_1439);
xnor U1644 (N_1644,N_1518,N_1401);
xnor U1645 (N_1645,N_1460,N_1443);
and U1646 (N_1646,N_1551,N_1453);
nor U1647 (N_1647,N_1519,N_1532);
nand U1648 (N_1648,N_1517,N_1475);
and U1649 (N_1649,N_1547,N_1531);
nand U1650 (N_1650,N_1546,N_1522);
nor U1651 (N_1651,N_1494,N_1470);
and U1652 (N_1652,N_1498,N_1421);
and U1653 (N_1653,N_1441,N_1527);
nand U1654 (N_1654,N_1458,N_1560);
nor U1655 (N_1655,N_1423,N_1418);
or U1656 (N_1656,N_1506,N_1479);
xor U1657 (N_1657,N_1579,N_1542);
or U1658 (N_1658,N_1572,N_1428);
or U1659 (N_1659,N_1573,N_1575);
xor U1660 (N_1660,N_1578,N_1464);
and U1661 (N_1661,N_1448,N_1574);
nor U1662 (N_1662,N_1500,N_1557);
nor U1663 (N_1663,N_1538,N_1407);
nand U1664 (N_1664,N_1540,N_1592);
and U1665 (N_1665,N_1452,N_1417);
or U1666 (N_1666,N_1548,N_1541);
and U1667 (N_1667,N_1432,N_1410);
and U1668 (N_1668,N_1446,N_1402);
nand U1669 (N_1669,N_1580,N_1556);
or U1670 (N_1670,N_1435,N_1400);
or U1671 (N_1671,N_1577,N_1521);
xor U1672 (N_1672,N_1406,N_1491);
and U1673 (N_1673,N_1444,N_1454);
xor U1674 (N_1674,N_1509,N_1485);
and U1675 (N_1675,N_1537,N_1412);
and U1676 (N_1676,N_1459,N_1431);
nand U1677 (N_1677,N_1501,N_1526);
and U1678 (N_1678,N_1429,N_1596);
nand U1679 (N_1679,N_1430,N_1535);
or U1680 (N_1680,N_1533,N_1585);
nor U1681 (N_1681,N_1422,N_1487);
and U1682 (N_1682,N_1438,N_1524);
or U1683 (N_1683,N_1558,N_1436);
xor U1684 (N_1684,N_1513,N_1478);
xnor U1685 (N_1685,N_1456,N_1595);
or U1686 (N_1686,N_1529,N_1503);
and U1687 (N_1687,N_1445,N_1507);
or U1688 (N_1688,N_1405,N_1514);
nor U1689 (N_1689,N_1450,N_1457);
nand U1690 (N_1690,N_1564,N_1511);
nand U1691 (N_1691,N_1562,N_1510);
nand U1692 (N_1692,N_1440,N_1587);
or U1693 (N_1693,N_1447,N_1559);
nor U1694 (N_1694,N_1515,N_1420);
nor U1695 (N_1695,N_1593,N_1434);
and U1696 (N_1696,N_1588,N_1404);
xnor U1697 (N_1697,N_1449,N_1419);
and U1698 (N_1698,N_1508,N_1484);
xnor U1699 (N_1699,N_1536,N_1493);
nor U1700 (N_1700,N_1432,N_1512);
and U1701 (N_1701,N_1573,N_1433);
nor U1702 (N_1702,N_1577,N_1439);
nand U1703 (N_1703,N_1560,N_1580);
nor U1704 (N_1704,N_1589,N_1482);
or U1705 (N_1705,N_1492,N_1560);
xor U1706 (N_1706,N_1440,N_1582);
and U1707 (N_1707,N_1483,N_1546);
nand U1708 (N_1708,N_1575,N_1516);
xnor U1709 (N_1709,N_1471,N_1574);
or U1710 (N_1710,N_1599,N_1475);
and U1711 (N_1711,N_1422,N_1451);
and U1712 (N_1712,N_1428,N_1404);
and U1713 (N_1713,N_1546,N_1467);
xnor U1714 (N_1714,N_1586,N_1527);
and U1715 (N_1715,N_1424,N_1476);
nand U1716 (N_1716,N_1429,N_1492);
nor U1717 (N_1717,N_1521,N_1410);
nor U1718 (N_1718,N_1463,N_1478);
nand U1719 (N_1719,N_1510,N_1443);
and U1720 (N_1720,N_1495,N_1463);
nand U1721 (N_1721,N_1524,N_1580);
or U1722 (N_1722,N_1559,N_1571);
nand U1723 (N_1723,N_1515,N_1579);
and U1724 (N_1724,N_1424,N_1500);
nor U1725 (N_1725,N_1481,N_1457);
nor U1726 (N_1726,N_1457,N_1432);
nor U1727 (N_1727,N_1514,N_1595);
xor U1728 (N_1728,N_1478,N_1533);
nor U1729 (N_1729,N_1595,N_1429);
nand U1730 (N_1730,N_1566,N_1402);
or U1731 (N_1731,N_1573,N_1467);
and U1732 (N_1732,N_1532,N_1452);
and U1733 (N_1733,N_1594,N_1450);
xor U1734 (N_1734,N_1445,N_1509);
nor U1735 (N_1735,N_1500,N_1523);
nand U1736 (N_1736,N_1510,N_1565);
and U1737 (N_1737,N_1402,N_1588);
or U1738 (N_1738,N_1555,N_1583);
and U1739 (N_1739,N_1552,N_1564);
nand U1740 (N_1740,N_1469,N_1498);
xor U1741 (N_1741,N_1573,N_1583);
and U1742 (N_1742,N_1468,N_1464);
xnor U1743 (N_1743,N_1434,N_1414);
xor U1744 (N_1744,N_1425,N_1420);
or U1745 (N_1745,N_1524,N_1556);
and U1746 (N_1746,N_1401,N_1541);
nor U1747 (N_1747,N_1426,N_1435);
nor U1748 (N_1748,N_1596,N_1512);
nand U1749 (N_1749,N_1577,N_1495);
nand U1750 (N_1750,N_1541,N_1451);
nor U1751 (N_1751,N_1528,N_1418);
nand U1752 (N_1752,N_1589,N_1459);
or U1753 (N_1753,N_1474,N_1434);
nand U1754 (N_1754,N_1529,N_1475);
nand U1755 (N_1755,N_1454,N_1528);
nand U1756 (N_1756,N_1536,N_1503);
nor U1757 (N_1757,N_1464,N_1507);
or U1758 (N_1758,N_1474,N_1513);
nor U1759 (N_1759,N_1416,N_1543);
xnor U1760 (N_1760,N_1596,N_1598);
nor U1761 (N_1761,N_1506,N_1487);
nand U1762 (N_1762,N_1584,N_1452);
and U1763 (N_1763,N_1574,N_1430);
and U1764 (N_1764,N_1589,N_1403);
nor U1765 (N_1765,N_1482,N_1475);
or U1766 (N_1766,N_1412,N_1549);
nand U1767 (N_1767,N_1540,N_1532);
xnor U1768 (N_1768,N_1456,N_1455);
nor U1769 (N_1769,N_1538,N_1552);
or U1770 (N_1770,N_1440,N_1592);
or U1771 (N_1771,N_1561,N_1507);
nand U1772 (N_1772,N_1418,N_1554);
nor U1773 (N_1773,N_1495,N_1594);
or U1774 (N_1774,N_1420,N_1418);
or U1775 (N_1775,N_1405,N_1576);
nor U1776 (N_1776,N_1562,N_1502);
nand U1777 (N_1777,N_1453,N_1529);
or U1778 (N_1778,N_1567,N_1419);
or U1779 (N_1779,N_1491,N_1439);
nor U1780 (N_1780,N_1431,N_1532);
nor U1781 (N_1781,N_1563,N_1402);
or U1782 (N_1782,N_1540,N_1450);
and U1783 (N_1783,N_1483,N_1497);
nand U1784 (N_1784,N_1572,N_1436);
and U1785 (N_1785,N_1422,N_1485);
xor U1786 (N_1786,N_1576,N_1506);
xnor U1787 (N_1787,N_1421,N_1453);
xnor U1788 (N_1788,N_1554,N_1547);
nand U1789 (N_1789,N_1557,N_1450);
nand U1790 (N_1790,N_1519,N_1545);
nand U1791 (N_1791,N_1556,N_1543);
or U1792 (N_1792,N_1540,N_1499);
or U1793 (N_1793,N_1474,N_1547);
or U1794 (N_1794,N_1495,N_1557);
xnor U1795 (N_1795,N_1439,N_1465);
nand U1796 (N_1796,N_1492,N_1511);
nand U1797 (N_1797,N_1502,N_1401);
nand U1798 (N_1798,N_1579,N_1580);
nand U1799 (N_1799,N_1497,N_1520);
or U1800 (N_1800,N_1786,N_1684);
nor U1801 (N_1801,N_1642,N_1707);
or U1802 (N_1802,N_1772,N_1657);
nor U1803 (N_1803,N_1637,N_1700);
nor U1804 (N_1804,N_1618,N_1635);
nand U1805 (N_1805,N_1660,N_1658);
or U1806 (N_1806,N_1735,N_1783);
xnor U1807 (N_1807,N_1788,N_1687);
and U1808 (N_1808,N_1621,N_1779);
nor U1809 (N_1809,N_1732,N_1799);
xor U1810 (N_1810,N_1716,N_1787);
or U1811 (N_1811,N_1746,N_1741);
xnor U1812 (N_1812,N_1633,N_1724);
or U1813 (N_1813,N_1720,N_1763);
and U1814 (N_1814,N_1625,N_1714);
nor U1815 (N_1815,N_1774,N_1636);
nand U1816 (N_1816,N_1723,N_1758);
or U1817 (N_1817,N_1639,N_1622);
nor U1818 (N_1818,N_1740,N_1756);
nand U1819 (N_1819,N_1792,N_1781);
nand U1820 (N_1820,N_1793,N_1797);
or U1821 (N_1821,N_1631,N_1722);
and U1822 (N_1822,N_1701,N_1680);
nor U1823 (N_1823,N_1780,N_1683);
nor U1824 (N_1824,N_1685,N_1778);
nand U1825 (N_1825,N_1659,N_1713);
or U1826 (N_1826,N_1769,N_1726);
nor U1827 (N_1827,N_1750,N_1668);
or U1828 (N_1828,N_1616,N_1688);
nand U1829 (N_1829,N_1706,N_1730);
xor U1830 (N_1830,N_1738,N_1754);
and U1831 (N_1831,N_1646,N_1747);
and U1832 (N_1832,N_1753,N_1663);
nor U1833 (N_1833,N_1605,N_1613);
and U1834 (N_1834,N_1640,N_1695);
and U1835 (N_1835,N_1798,N_1785);
xnor U1836 (N_1836,N_1694,N_1692);
xnor U1837 (N_1837,N_1766,N_1734);
and U1838 (N_1838,N_1752,N_1702);
nor U1839 (N_1839,N_1654,N_1665);
nand U1840 (N_1840,N_1782,N_1759);
xnor U1841 (N_1841,N_1727,N_1630);
nor U1842 (N_1842,N_1729,N_1667);
nor U1843 (N_1843,N_1655,N_1608);
nor U1844 (N_1844,N_1617,N_1629);
and U1845 (N_1845,N_1682,N_1719);
and U1846 (N_1846,N_1762,N_1796);
or U1847 (N_1847,N_1760,N_1689);
and U1848 (N_1848,N_1773,N_1674);
or U1849 (N_1849,N_1623,N_1711);
nor U1850 (N_1850,N_1653,N_1691);
nand U1851 (N_1851,N_1661,N_1651);
or U1852 (N_1852,N_1705,N_1696);
xor U1853 (N_1853,N_1632,N_1764);
nor U1854 (N_1854,N_1709,N_1767);
nand U1855 (N_1855,N_1765,N_1673);
and U1856 (N_1856,N_1771,N_1677);
and U1857 (N_1857,N_1690,N_1790);
nor U1858 (N_1858,N_1607,N_1606);
nand U1859 (N_1859,N_1755,N_1645);
nand U1860 (N_1860,N_1610,N_1670);
or U1861 (N_1861,N_1619,N_1679);
or U1862 (N_1862,N_1662,N_1676);
or U1863 (N_1863,N_1656,N_1770);
xor U1864 (N_1864,N_1697,N_1603);
nand U1865 (N_1865,N_1628,N_1733);
nand U1866 (N_1866,N_1601,N_1698);
xor U1867 (N_1867,N_1664,N_1784);
nand U1868 (N_1868,N_1743,N_1717);
or U1869 (N_1869,N_1681,N_1641);
xnor U1870 (N_1870,N_1600,N_1794);
or U1871 (N_1871,N_1736,N_1672);
nor U1872 (N_1872,N_1748,N_1614);
nor U1873 (N_1873,N_1739,N_1777);
or U1874 (N_1874,N_1650,N_1638);
xor U1875 (N_1875,N_1731,N_1620);
and U1876 (N_1876,N_1744,N_1634);
nand U1877 (N_1877,N_1699,N_1712);
or U1878 (N_1878,N_1615,N_1666);
nand U1879 (N_1879,N_1761,N_1757);
or U1880 (N_1880,N_1791,N_1612);
nand U1881 (N_1881,N_1718,N_1675);
nand U1882 (N_1882,N_1609,N_1611);
or U1883 (N_1883,N_1721,N_1643);
and U1884 (N_1884,N_1768,N_1710);
or U1885 (N_1885,N_1604,N_1789);
nor U1886 (N_1886,N_1671,N_1704);
or U1887 (N_1887,N_1644,N_1751);
xnor U1888 (N_1888,N_1649,N_1602);
nor U1889 (N_1889,N_1749,N_1715);
xnor U1890 (N_1890,N_1775,N_1725);
nand U1891 (N_1891,N_1728,N_1742);
and U1892 (N_1892,N_1703,N_1652);
nand U1893 (N_1893,N_1745,N_1795);
and U1894 (N_1894,N_1776,N_1678);
xor U1895 (N_1895,N_1648,N_1708);
xnor U1896 (N_1896,N_1669,N_1647);
nand U1897 (N_1897,N_1686,N_1693);
and U1898 (N_1898,N_1624,N_1627);
or U1899 (N_1899,N_1626,N_1737);
xnor U1900 (N_1900,N_1743,N_1759);
xnor U1901 (N_1901,N_1616,N_1777);
and U1902 (N_1902,N_1627,N_1740);
xnor U1903 (N_1903,N_1614,N_1784);
nor U1904 (N_1904,N_1691,N_1621);
and U1905 (N_1905,N_1795,N_1703);
and U1906 (N_1906,N_1719,N_1741);
or U1907 (N_1907,N_1691,N_1698);
nor U1908 (N_1908,N_1652,N_1645);
or U1909 (N_1909,N_1675,N_1759);
and U1910 (N_1910,N_1739,N_1625);
and U1911 (N_1911,N_1692,N_1684);
and U1912 (N_1912,N_1600,N_1752);
xnor U1913 (N_1913,N_1737,N_1630);
xor U1914 (N_1914,N_1646,N_1769);
or U1915 (N_1915,N_1761,N_1769);
xor U1916 (N_1916,N_1728,N_1650);
and U1917 (N_1917,N_1730,N_1788);
nand U1918 (N_1918,N_1600,N_1746);
or U1919 (N_1919,N_1632,N_1698);
nor U1920 (N_1920,N_1796,N_1672);
or U1921 (N_1921,N_1656,N_1657);
nand U1922 (N_1922,N_1795,N_1763);
nor U1923 (N_1923,N_1780,N_1668);
xor U1924 (N_1924,N_1683,N_1609);
or U1925 (N_1925,N_1627,N_1730);
xor U1926 (N_1926,N_1656,N_1794);
xor U1927 (N_1927,N_1660,N_1685);
nand U1928 (N_1928,N_1608,N_1662);
and U1929 (N_1929,N_1621,N_1795);
and U1930 (N_1930,N_1621,N_1752);
or U1931 (N_1931,N_1791,N_1608);
nor U1932 (N_1932,N_1672,N_1635);
and U1933 (N_1933,N_1607,N_1743);
or U1934 (N_1934,N_1638,N_1680);
and U1935 (N_1935,N_1654,N_1769);
nor U1936 (N_1936,N_1650,N_1768);
nand U1937 (N_1937,N_1776,N_1731);
nor U1938 (N_1938,N_1666,N_1684);
and U1939 (N_1939,N_1633,N_1670);
xor U1940 (N_1940,N_1789,N_1770);
or U1941 (N_1941,N_1688,N_1791);
and U1942 (N_1942,N_1616,N_1644);
nor U1943 (N_1943,N_1615,N_1704);
xor U1944 (N_1944,N_1646,N_1763);
nor U1945 (N_1945,N_1656,N_1686);
nor U1946 (N_1946,N_1698,N_1780);
or U1947 (N_1947,N_1700,N_1775);
or U1948 (N_1948,N_1657,N_1692);
nand U1949 (N_1949,N_1748,N_1650);
and U1950 (N_1950,N_1719,N_1668);
or U1951 (N_1951,N_1629,N_1761);
or U1952 (N_1952,N_1667,N_1650);
and U1953 (N_1953,N_1639,N_1766);
nor U1954 (N_1954,N_1636,N_1795);
xnor U1955 (N_1955,N_1786,N_1623);
or U1956 (N_1956,N_1694,N_1654);
or U1957 (N_1957,N_1769,N_1625);
and U1958 (N_1958,N_1663,N_1770);
nor U1959 (N_1959,N_1603,N_1678);
xnor U1960 (N_1960,N_1635,N_1722);
and U1961 (N_1961,N_1668,N_1756);
or U1962 (N_1962,N_1736,N_1738);
xor U1963 (N_1963,N_1680,N_1725);
xnor U1964 (N_1964,N_1664,N_1693);
and U1965 (N_1965,N_1734,N_1716);
nand U1966 (N_1966,N_1743,N_1795);
xor U1967 (N_1967,N_1794,N_1713);
nand U1968 (N_1968,N_1643,N_1727);
or U1969 (N_1969,N_1621,N_1783);
xor U1970 (N_1970,N_1771,N_1670);
nor U1971 (N_1971,N_1761,N_1763);
xnor U1972 (N_1972,N_1696,N_1683);
xnor U1973 (N_1973,N_1733,N_1691);
xor U1974 (N_1974,N_1635,N_1621);
and U1975 (N_1975,N_1701,N_1675);
xnor U1976 (N_1976,N_1681,N_1717);
xnor U1977 (N_1977,N_1761,N_1726);
and U1978 (N_1978,N_1750,N_1629);
xnor U1979 (N_1979,N_1696,N_1631);
or U1980 (N_1980,N_1654,N_1759);
xnor U1981 (N_1981,N_1703,N_1659);
or U1982 (N_1982,N_1698,N_1645);
or U1983 (N_1983,N_1727,N_1609);
and U1984 (N_1984,N_1600,N_1737);
and U1985 (N_1985,N_1614,N_1794);
xor U1986 (N_1986,N_1733,N_1661);
nor U1987 (N_1987,N_1618,N_1647);
nand U1988 (N_1988,N_1602,N_1684);
and U1989 (N_1989,N_1784,N_1794);
or U1990 (N_1990,N_1737,N_1757);
nand U1991 (N_1991,N_1613,N_1620);
nor U1992 (N_1992,N_1741,N_1718);
or U1993 (N_1993,N_1620,N_1789);
nand U1994 (N_1994,N_1718,N_1767);
xor U1995 (N_1995,N_1602,N_1642);
nand U1996 (N_1996,N_1676,N_1672);
or U1997 (N_1997,N_1734,N_1675);
nor U1998 (N_1998,N_1723,N_1659);
xnor U1999 (N_1999,N_1639,N_1796);
or U2000 (N_2000,N_1831,N_1913);
xnor U2001 (N_2001,N_1800,N_1891);
nor U2002 (N_2002,N_1839,N_1960);
or U2003 (N_2003,N_1927,N_1953);
nor U2004 (N_2004,N_1904,N_1855);
and U2005 (N_2005,N_1849,N_1887);
xnor U2006 (N_2006,N_1914,N_1883);
or U2007 (N_2007,N_1888,N_1947);
xnor U2008 (N_2008,N_1861,N_1840);
and U2009 (N_2009,N_1973,N_1818);
or U2010 (N_2010,N_1827,N_1907);
xor U2011 (N_2011,N_1999,N_1988);
nand U2012 (N_2012,N_1810,N_1903);
nor U2013 (N_2013,N_1983,N_1975);
xor U2014 (N_2014,N_1943,N_1902);
xor U2015 (N_2015,N_1828,N_1823);
nor U2016 (N_2016,N_1928,N_1994);
nor U2017 (N_2017,N_1844,N_1950);
and U2018 (N_2018,N_1972,N_1964);
xnor U2019 (N_2019,N_1857,N_1846);
xor U2020 (N_2020,N_1874,N_1854);
nor U2021 (N_2021,N_1921,N_1954);
xnor U2022 (N_2022,N_1815,N_1880);
nor U2023 (N_2023,N_1935,N_1952);
nor U2024 (N_2024,N_1867,N_1836);
xor U2025 (N_2025,N_1978,N_1872);
nor U2026 (N_2026,N_1982,N_1966);
nand U2027 (N_2027,N_1929,N_1932);
xnor U2028 (N_2028,N_1882,N_1822);
xnor U2029 (N_2029,N_1871,N_1866);
nand U2030 (N_2030,N_1897,N_1924);
nor U2031 (N_2031,N_1826,N_1911);
nand U2032 (N_2032,N_1816,N_1944);
xor U2033 (N_2033,N_1976,N_1915);
and U2034 (N_2034,N_1885,N_1918);
or U2035 (N_2035,N_1884,N_1837);
and U2036 (N_2036,N_1968,N_1958);
and U2037 (N_2037,N_1990,N_1847);
nor U2038 (N_2038,N_1858,N_1959);
xor U2039 (N_2039,N_1895,N_1870);
nor U2040 (N_2040,N_1908,N_1851);
xor U2041 (N_2041,N_1868,N_1808);
or U2042 (N_2042,N_1899,N_1989);
nand U2043 (N_2043,N_1813,N_1946);
or U2044 (N_2044,N_1859,N_1969);
and U2045 (N_2045,N_1949,N_1820);
nand U2046 (N_2046,N_1862,N_1940);
nand U2047 (N_2047,N_1900,N_1951);
and U2048 (N_2048,N_1876,N_1995);
or U2049 (N_2049,N_1869,N_1957);
nor U2050 (N_2050,N_1937,N_1802);
or U2051 (N_2051,N_1805,N_1873);
nand U2052 (N_2052,N_1838,N_1987);
and U2053 (N_2053,N_1925,N_1930);
xnor U2054 (N_2054,N_1910,N_1821);
or U2055 (N_2055,N_1898,N_1878);
nor U2056 (N_2056,N_1890,N_1970);
nor U2057 (N_2057,N_1906,N_1916);
nor U2058 (N_2058,N_1892,N_1830);
and U2059 (N_2059,N_1835,N_1825);
xnor U2060 (N_2060,N_1986,N_1894);
xor U2061 (N_2061,N_1850,N_1931);
and U2062 (N_2062,N_1956,N_1981);
xnor U2063 (N_2063,N_1893,N_1853);
nand U2064 (N_2064,N_1948,N_1991);
nor U2065 (N_2065,N_1967,N_1809);
and U2066 (N_2066,N_1863,N_1992);
nand U2067 (N_2067,N_1814,N_1961);
or U2068 (N_2068,N_1933,N_1997);
nand U2069 (N_2069,N_1905,N_1984);
xor U2070 (N_2070,N_1920,N_1881);
and U2071 (N_2071,N_1980,N_1841);
nor U2072 (N_2072,N_1977,N_1803);
nor U2073 (N_2073,N_1865,N_1834);
or U2074 (N_2074,N_1917,N_1819);
nand U2075 (N_2075,N_1896,N_1945);
nor U2076 (N_2076,N_1955,N_1812);
nand U2077 (N_2077,N_1875,N_1993);
or U2078 (N_2078,N_1806,N_1886);
nand U2079 (N_2079,N_1934,N_1804);
xor U2080 (N_2080,N_1996,N_1912);
xor U2081 (N_2081,N_1807,N_1856);
nor U2082 (N_2082,N_1909,N_1962);
or U2083 (N_2083,N_1963,N_1843);
nor U2084 (N_2084,N_1833,N_1860);
nand U2085 (N_2085,N_1845,N_1879);
nor U2086 (N_2086,N_1832,N_1965);
or U2087 (N_2087,N_1829,N_1842);
or U2088 (N_2088,N_1877,N_1889);
and U2089 (N_2089,N_1923,N_1901);
nand U2090 (N_2090,N_1848,N_1864);
nor U2091 (N_2091,N_1811,N_1801);
nand U2092 (N_2092,N_1942,N_1939);
nand U2093 (N_2093,N_1926,N_1852);
nor U2094 (N_2094,N_1919,N_1941);
nor U2095 (N_2095,N_1979,N_1971);
nand U2096 (N_2096,N_1817,N_1985);
xnor U2097 (N_2097,N_1938,N_1974);
and U2098 (N_2098,N_1824,N_1998);
nor U2099 (N_2099,N_1936,N_1922);
nand U2100 (N_2100,N_1837,N_1849);
nor U2101 (N_2101,N_1895,N_1884);
nand U2102 (N_2102,N_1953,N_1983);
and U2103 (N_2103,N_1924,N_1900);
and U2104 (N_2104,N_1829,N_1915);
nand U2105 (N_2105,N_1871,N_1885);
nor U2106 (N_2106,N_1842,N_1991);
xnor U2107 (N_2107,N_1801,N_1983);
nor U2108 (N_2108,N_1803,N_1875);
nand U2109 (N_2109,N_1881,N_1893);
nand U2110 (N_2110,N_1871,N_1835);
nor U2111 (N_2111,N_1933,N_1945);
nand U2112 (N_2112,N_1974,N_1879);
nor U2113 (N_2113,N_1836,N_1950);
nand U2114 (N_2114,N_1820,N_1876);
or U2115 (N_2115,N_1810,N_1984);
and U2116 (N_2116,N_1861,N_1814);
nand U2117 (N_2117,N_1846,N_1865);
nand U2118 (N_2118,N_1838,N_1814);
xnor U2119 (N_2119,N_1812,N_1854);
or U2120 (N_2120,N_1993,N_1817);
nand U2121 (N_2121,N_1864,N_1826);
nor U2122 (N_2122,N_1820,N_1905);
nor U2123 (N_2123,N_1800,N_1991);
or U2124 (N_2124,N_1984,N_1985);
nor U2125 (N_2125,N_1876,N_1999);
xnor U2126 (N_2126,N_1865,N_1819);
and U2127 (N_2127,N_1986,N_1875);
nand U2128 (N_2128,N_1923,N_1855);
nor U2129 (N_2129,N_1892,N_1951);
or U2130 (N_2130,N_1975,N_1921);
and U2131 (N_2131,N_1816,N_1991);
nand U2132 (N_2132,N_1884,N_1812);
nand U2133 (N_2133,N_1927,N_1981);
xor U2134 (N_2134,N_1800,N_1999);
nor U2135 (N_2135,N_1960,N_1902);
nand U2136 (N_2136,N_1994,N_1944);
nand U2137 (N_2137,N_1859,N_1931);
or U2138 (N_2138,N_1986,N_1933);
nor U2139 (N_2139,N_1927,N_1844);
nand U2140 (N_2140,N_1994,N_1979);
or U2141 (N_2141,N_1959,N_1979);
and U2142 (N_2142,N_1984,N_1971);
nand U2143 (N_2143,N_1995,N_1869);
and U2144 (N_2144,N_1942,N_1818);
nand U2145 (N_2145,N_1905,N_1811);
nor U2146 (N_2146,N_1803,N_1840);
nand U2147 (N_2147,N_1828,N_1829);
nand U2148 (N_2148,N_1942,N_1940);
nand U2149 (N_2149,N_1886,N_1875);
and U2150 (N_2150,N_1809,N_1920);
or U2151 (N_2151,N_1880,N_1970);
or U2152 (N_2152,N_1890,N_1907);
nand U2153 (N_2153,N_1989,N_1853);
nand U2154 (N_2154,N_1815,N_1937);
nor U2155 (N_2155,N_1838,N_1959);
or U2156 (N_2156,N_1819,N_1929);
xor U2157 (N_2157,N_1958,N_1938);
xnor U2158 (N_2158,N_1909,N_1914);
and U2159 (N_2159,N_1878,N_1893);
nand U2160 (N_2160,N_1966,N_1960);
nand U2161 (N_2161,N_1998,N_1909);
xnor U2162 (N_2162,N_1908,N_1902);
nor U2163 (N_2163,N_1868,N_1877);
or U2164 (N_2164,N_1819,N_1822);
nand U2165 (N_2165,N_1827,N_1843);
nor U2166 (N_2166,N_1825,N_1955);
nand U2167 (N_2167,N_1985,N_1915);
xnor U2168 (N_2168,N_1880,N_1809);
and U2169 (N_2169,N_1918,N_1851);
nand U2170 (N_2170,N_1958,N_1810);
nor U2171 (N_2171,N_1809,N_1917);
xnor U2172 (N_2172,N_1864,N_1808);
or U2173 (N_2173,N_1976,N_1866);
and U2174 (N_2174,N_1951,N_1813);
xor U2175 (N_2175,N_1816,N_1841);
or U2176 (N_2176,N_1852,N_1857);
or U2177 (N_2177,N_1884,N_1954);
nor U2178 (N_2178,N_1849,N_1823);
xnor U2179 (N_2179,N_1807,N_1910);
nor U2180 (N_2180,N_1819,N_1942);
xor U2181 (N_2181,N_1805,N_1925);
or U2182 (N_2182,N_1941,N_1907);
nor U2183 (N_2183,N_1996,N_1963);
or U2184 (N_2184,N_1901,N_1885);
xnor U2185 (N_2185,N_1903,N_1805);
or U2186 (N_2186,N_1827,N_1937);
or U2187 (N_2187,N_1996,N_1873);
nor U2188 (N_2188,N_1821,N_1945);
or U2189 (N_2189,N_1919,N_1981);
nor U2190 (N_2190,N_1803,N_1881);
and U2191 (N_2191,N_1883,N_1946);
nand U2192 (N_2192,N_1997,N_1834);
nor U2193 (N_2193,N_1998,N_1941);
or U2194 (N_2194,N_1855,N_1877);
or U2195 (N_2195,N_1804,N_1964);
or U2196 (N_2196,N_1861,N_1960);
xor U2197 (N_2197,N_1809,N_1841);
or U2198 (N_2198,N_1962,N_1986);
nand U2199 (N_2199,N_1860,N_1897);
xnor U2200 (N_2200,N_2123,N_2084);
and U2201 (N_2201,N_2111,N_2106);
xor U2202 (N_2202,N_2082,N_2169);
or U2203 (N_2203,N_2160,N_2051);
xnor U2204 (N_2204,N_2096,N_2011);
or U2205 (N_2205,N_2062,N_2181);
nand U2206 (N_2206,N_2069,N_2012);
or U2207 (N_2207,N_2185,N_2018);
nor U2208 (N_2208,N_2162,N_2146);
xor U2209 (N_2209,N_2014,N_2035);
nor U2210 (N_2210,N_2050,N_2141);
or U2211 (N_2211,N_2030,N_2006);
or U2212 (N_2212,N_2187,N_2139);
nand U2213 (N_2213,N_2191,N_2022);
and U2214 (N_2214,N_2131,N_2075);
and U2215 (N_2215,N_2168,N_2138);
nand U2216 (N_2216,N_2130,N_2193);
xnor U2217 (N_2217,N_2060,N_2180);
or U2218 (N_2218,N_2097,N_2100);
nand U2219 (N_2219,N_2054,N_2026);
xor U2220 (N_2220,N_2170,N_2016);
and U2221 (N_2221,N_2000,N_2017);
and U2222 (N_2222,N_2064,N_2099);
nor U2223 (N_2223,N_2009,N_2145);
nor U2224 (N_2224,N_2110,N_2190);
and U2225 (N_2225,N_2135,N_2116);
nand U2226 (N_2226,N_2189,N_2163);
and U2227 (N_2227,N_2152,N_2118);
nor U2228 (N_2228,N_2129,N_2144);
nor U2229 (N_2229,N_2002,N_2134);
xnor U2230 (N_2230,N_2036,N_2045);
xnor U2231 (N_2231,N_2042,N_2033);
and U2232 (N_2232,N_2098,N_2092);
and U2233 (N_2233,N_2005,N_2056);
xor U2234 (N_2234,N_2159,N_2108);
xnor U2235 (N_2235,N_2117,N_2175);
and U2236 (N_2236,N_2137,N_2028);
or U2237 (N_2237,N_2120,N_2044);
xnor U2238 (N_2238,N_2188,N_2074);
nand U2239 (N_2239,N_2150,N_2133);
nand U2240 (N_2240,N_2156,N_2077);
or U2241 (N_2241,N_2052,N_2085);
or U2242 (N_2242,N_2122,N_2158);
nand U2243 (N_2243,N_2171,N_2031);
nand U2244 (N_2244,N_2010,N_2081);
nand U2245 (N_2245,N_2102,N_2029);
nor U2246 (N_2246,N_2032,N_2182);
and U2247 (N_2247,N_2046,N_2040);
or U2248 (N_2248,N_2184,N_2024);
or U2249 (N_2249,N_2019,N_2015);
xor U2250 (N_2250,N_2073,N_2151);
nand U2251 (N_2251,N_2166,N_2174);
xor U2252 (N_2252,N_2186,N_2065);
or U2253 (N_2253,N_2061,N_2196);
nor U2254 (N_2254,N_2148,N_2067);
nand U2255 (N_2255,N_2004,N_2066);
or U2256 (N_2256,N_2178,N_2027);
xnor U2257 (N_2257,N_2025,N_2078);
nor U2258 (N_2258,N_2173,N_2070);
nand U2259 (N_2259,N_2128,N_2071);
xor U2260 (N_2260,N_2080,N_2199);
xor U2261 (N_2261,N_2104,N_2140);
and U2262 (N_2262,N_2093,N_2149);
nand U2263 (N_2263,N_2127,N_2119);
or U2264 (N_2264,N_2087,N_2124);
xnor U2265 (N_2265,N_2153,N_2109);
or U2266 (N_2266,N_2083,N_2115);
nor U2267 (N_2267,N_2195,N_2089);
nor U2268 (N_2268,N_2086,N_2095);
and U2269 (N_2269,N_2063,N_2001);
nand U2270 (N_2270,N_2079,N_2113);
xnor U2271 (N_2271,N_2101,N_2161);
nor U2272 (N_2272,N_2041,N_2072);
nor U2273 (N_2273,N_2198,N_2157);
nor U2274 (N_2274,N_2176,N_2091);
nand U2275 (N_2275,N_2155,N_2197);
or U2276 (N_2276,N_2039,N_2167);
and U2277 (N_2277,N_2021,N_2132);
nand U2278 (N_2278,N_2112,N_2007);
xnor U2279 (N_2279,N_2142,N_2003);
and U2280 (N_2280,N_2121,N_2103);
and U2281 (N_2281,N_2090,N_2055);
or U2282 (N_2282,N_2023,N_2013);
and U2283 (N_2283,N_2107,N_2154);
nand U2284 (N_2284,N_2047,N_2177);
and U2285 (N_2285,N_2088,N_2038);
nand U2286 (N_2286,N_2114,N_2020);
or U2287 (N_2287,N_2057,N_2105);
xnor U2288 (N_2288,N_2183,N_2059);
xor U2289 (N_2289,N_2147,N_2094);
nand U2290 (N_2290,N_2165,N_2037);
xnor U2291 (N_2291,N_2136,N_2068);
xor U2292 (N_2292,N_2076,N_2172);
xor U2293 (N_2293,N_2164,N_2034);
nor U2294 (N_2294,N_2143,N_2049);
or U2295 (N_2295,N_2058,N_2194);
or U2296 (N_2296,N_2179,N_2126);
and U2297 (N_2297,N_2048,N_2043);
or U2298 (N_2298,N_2008,N_2125);
xor U2299 (N_2299,N_2192,N_2053);
and U2300 (N_2300,N_2091,N_2068);
xor U2301 (N_2301,N_2032,N_2010);
nor U2302 (N_2302,N_2030,N_2066);
or U2303 (N_2303,N_2127,N_2148);
and U2304 (N_2304,N_2076,N_2005);
nor U2305 (N_2305,N_2069,N_2155);
nor U2306 (N_2306,N_2045,N_2013);
xor U2307 (N_2307,N_2052,N_2178);
or U2308 (N_2308,N_2182,N_2090);
nor U2309 (N_2309,N_2061,N_2097);
nand U2310 (N_2310,N_2068,N_2004);
or U2311 (N_2311,N_2062,N_2090);
and U2312 (N_2312,N_2166,N_2137);
and U2313 (N_2313,N_2052,N_2096);
xor U2314 (N_2314,N_2037,N_2016);
xnor U2315 (N_2315,N_2104,N_2011);
or U2316 (N_2316,N_2102,N_2053);
or U2317 (N_2317,N_2134,N_2023);
nor U2318 (N_2318,N_2192,N_2076);
nor U2319 (N_2319,N_2190,N_2128);
nand U2320 (N_2320,N_2069,N_2125);
nor U2321 (N_2321,N_2070,N_2039);
and U2322 (N_2322,N_2180,N_2138);
nand U2323 (N_2323,N_2137,N_2087);
or U2324 (N_2324,N_2100,N_2011);
nand U2325 (N_2325,N_2165,N_2013);
or U2326 (N_2326,N_2021,N_2175);
and U2327 (N_2327,N_2168,N_2009);
xor U2328 (N_2328,N_2191,N_2004);
nor U2329 (N_2329,N_2147,N_2033);
nor U2330 (N_2330,N_2120,N_2032);
and U2331 (N_2331,N_2176,N_2193);
or U2332 (N_2332,N_2185,N_2168);
and U2333 (N_2333,N_2039,N_2175);
nand U2334 (N_2334,N_2067,N_2000);
xor U2335 (N_2335,N_2097,N_2027);
nand U2336 (N_2336,N_2174,N_2172);
or U2337 (N_2337,N_2152,N_2051);
nor U2338 (N_2338,N_2022,N_2121);
nor U2339 (N_2339,N_2030,N_2143);
nand U2340 (N_2340,N_2088,N_2152);
nor U2341 (N_2341,N_2009,N_2086);
or U2342 (N_2342,N_2077,N_2056);
xor U2343 (N_2343,N_2130,N_2001);
and U2344 (N_2344,N_2111,N_2004);
or U2345 (N_2345,N_2064,N_2149);
or U2346 (N_2346,N_2136,N_2007);
nand U2347 (N_2347,N_2009,N_2196);
xnor U2348 (N_2348,N_2000,N_2125);
xnor U2349 (N_2349,N_2102,N_2147);
xor U2350 (N_2350,N_2153,N_2057);
xnor U2351 (N_2351,N_2025,N_2014);
or U2352 (N_2352,N_2093,N_2055);
nand U2353 (N_2353,N_2102,N_2163);
xnor U2354 (N_2354,N_2007,N_2027);
xnor U2355 (N_2355,N_2166,N_2043);
or U2356 (N_2356,N_2172,N_2063);
nor U2357 (N_2357,N_2093,N_2096);
nor U2358 (N_2358,N_2035,N_2163);
nand U2359 (N_2359,N_2155,N_2084);
nor U2360 (N_2360,N_2102,N_2014);
nand U2361 (N_2361,N_2000,N_2181);
nor U2362 (N_2362,N_2169,N_2198);
or U2363 (N_2363,N_2050,N_2167);
xor U2364 (N_2364,N_2192,N_2100);
or U2365 (N_2365,N_2103,N_2059);
and U2366 (N_2366,N_2066,N_2032);
nor U2367 (N_2367,N_2176,N_2166);
xor U2368 (N_2368,N_2150,N_2097);
xnor U2369 (N_2369,N_2074,N_2139);
and U2370 (N_2370,N_2034,N_2135);
xor U2371 (N_2371,N_2004,N_2012);
and U2372 (N_2372,N_2146,N_2037);
and U2373 (N_2373,N_2009,N_2124);
xnor U2374 (N_2374,N_2038,N_2047);
or U2375 (N_2375,N_2183,N_2139);
xnor U2376 (N_2376,N_2144,N_2152);
or U2377 (N_2377,N_2030,N_2078);
nand U2378 (N_2378,N_2190,N_2034);
and U2379 (N_2379,N_2054,N_2005);
or U2380 (N_2380,N_2133,N_2110);
or U2381 (N_2381,N_2108,N_2148);
and U2382 (N_2382,N_2144,N_2078);
and U2383 (N_2383,N_2145,N_2119);
and U2384 (N_2384,N_2069,N_2160);
nand U2385 (N_2385,N_2190,N_2064);
xnor U2386 (N_2386,N_2145,N_2188);
and U2387 (N_2387,N_2039,N_2041);
xnor U2388 (N_2388,N_2183,N_2138);
and U2389 (N_2389,N_2004,N_2073);
or U2390 (N_2390,N_2170,N_2125);
or U2391 (N_2391,N_2037,N_2170);
and U2392 (N_2392,N_2132,N_2041);
and U2393 (N_2393,N_2039,N_2145);
and U2394 (N_2394,N_2159,N_2121);
nor U2395 (N_2395,N_2014,N_2097);
or U2396 (N_2396,N_2131,N_2153);
and U2397 (N_2397,N_2172,N_2140);
nor U2398 (N_2398,N_2053,N_2036);
nor U2399 (N_2399,N_2135,N_2081);
xor U2400 (N_2400,N_2308,N_2255);
xor U2401 (N_2401,N_2243,N_2319);
or U2402 (N_2402,N_2377,N_2359);
and U2403 (N_2403,N_2303,N_2202);
and U2404 (N_2404,N_2291,N_2399);
nand U2405 (N_2405,N_2219,N_2336);
xnor U2406 (N_2406,N_2368,N_2299);
and U2407 (N_2407,N_2387,N_2221);
nand U2408 (N_2408,N_2309,N_2220);
or U2409 (N_2409,N_2206,N_2375);
nor U2410 (N_2410,N_2242,N_2305);
nor U2411 (N_2411,N_2320,N_2208);
xor U2412 (N_2412,N_2313,N_2280);
or U2413 (N_2413,N_2311,N_2223);
xnor U2414 (N_2414,N_2237,N_2371);
or U2415 (N_2415,N_2295,N_2342);
nand U2416 (N_2416,N_2279,N_2355);
and U2417 (N_2417,N_2318,N_2259);
nor U2418 (N_2418,N_2224,N_2276);
and U2419 (N_2419,N_2292,N_2373);
nand U2420 (N_2420,N_2257,N_2290);
or U2421 (N_2421,N_2338,N_2289);
xnor U2422 (N_2422,N_2334,N_2352);
nand U2423 (N_2423,N_2293,N_2235);
or U2424 (N_2424,N_2294,N_2260);
or U2425 (N_2425,N_2356,N_2272);
and U2426 (N_2426,N_2360,N_2332);
nor U2427 (N_2427,N_2370,N_2252);
or U2428 (N_2428,N_2204,N_2391);
or U2429 (N_2429,N_2364,N_2245);
xor U2430 (N_2430,N_2398,N_2273);
nand U2431 (N_2431,N_2265,N_2251);
nor U2432 (N_2432,N_2310,N_2383);
nor U2433 (N_2433,N_2327,N_2358);
nand U2434 (N_2434,N_2315,N_2286);
nand U2435 (N_2435,N_2312,N_2268);
or U2436 (N_2436,N_2306,N_2241);
and U2437 (N_2437,N_2266,N_2393);
or U2438 (N_2438,N_2350,N_2253);
and U2439 (N_2439,N_2304,N_2322);
xor U2440 (N_2440,N_2229,N_2230);
and U2441 (N_2441,N_2250,N_2234);
or U2442 (N_2442,N_2258,N_2329);
xor U2443 (N_2443,N_2264,N_2269);
or U2444 (N_2444,N_2385,N_2307);
or U2445 (N_2445,N_2348,N_2361);
nor U2446 (N_2446,N_2362,N_2381);
xnor U2447 (N_2447,N_2205,N_2382);
xor U2448 (N_2448,N_2366,N_2335);
and U2449 (N_2449,N_2300,N_2228);
xor U2450 (N_2450,N_2261,N_2215);
and U2451 (N_2451,N_2233,N_2270);
and U2452 (N_2452,N_2226,N_2301);
and U2453 (N_2453,N_2285,N_2214);
or U2454 (N_2454,N_2231,N_2324);
nand U2455 (N_2455,N_2248,N_2216);
xor U2456 (N_2456,N_2396,N_2331);
nand U2457 (N_2457,N_2256,N_2282);
and U2458 (N_2458,N_2277,N_2369);
or U2459 (N_2459,N_2351,N_2239);
nand U2460 (N_2460,N_2203,N_2288);
xor U2461 (N_2461,N_2343,N_2225);
or U2462 (N_2462,N_2298,N_2201);
nor U2463 (N_2463,N_2379,N_2394);
nor U2464 (N_2464,N_2314,N_2249);
and U2465 (N_2465,N_2263,N_2212);
nor U2466 (N_2466,N_2367,N_2222);
nand U2467 (N_2467,N_2207,N_2210);
or U2468 (N_2468,N_2341,N_2374);
xor U2469 (N_2469,N_2275,N_2386);
and U2470 (N_2470,N_2353,N_2376);
nor U2471 (N_2471,N_2246,N_2339);
and U2472 (N_2472,N_2213,N_2227);
nand U2473 (N_2473,N_2317,N_2278);
or U2474 (N_2474,N_2325,N_2283);
and U2475 (N_2475,N_2388,N_2232);
and U2476 (N_2476,N_2254,N_2200);
nor U2477 (N_2477,N_2330,N_2372);
or U2478 (N_2478,N_2392,N_2262);
and U2479 (N_2479,N_2247,N_2326);
nor U2480 (N_2480,N_2349,N_2380);
xnor U2481 (N_2481,N_2281,N_2217);
xnor U2482 (N_2482,N_2365,N_2321);
nor U2483 (N_2483,N_2384,N_2238);
nand U2484 (N_2484,N_2267,N_2236);
and U2485 (N_2485,N_2354,N_2302);
nand U2486 (N_2486,N_2218,N_2390);
and U2487 (N_2487,N_2389,N_2297);
nand U2488 (N_2488,N_2378,N_2287);
nor U2489 (N_2489,N_2209,N_2211);
and U2490 (N_2490,N_2347,N_2363);
nand U2491 (N_2491,N_2240,N_2337);
or U2492 (N_2492,N_2333,N_2328);
and U2493 (N_2493,N_2345,N_2395);
nor U2494 (N_2494,N_2244,N_2397);
and U2495 (N_2495,N_2323,N_2271);
and U2496 (N_2496,N_2284,N_2296);
nand U2497 (N_2497,N_2316,N_2274);
xnor U2498 (N_2498,N_2344,N_2340);
or U2499 (N_2499,N_2346,N_2357);
or U2500 (N_2500,N_2288,N_2245);
and U2501 (N_2501,N_2311,N_2217);
xnor U2502 (N_2502,N_2317,N_2313);
nor U2503 (N_2503,N_2295,N_2221);
or U2504 (N_2504,N_2315,N_2343);
or U2505 (N_2505,N_2333,N_2291);
nor U2506 (N_2506,N_2216,N_2267);
nand U2507 (N_2507,N_2378,N_2207);
and U2508 (N_2508,N_2325,N_2392);
xor U2509 (N_2509,N_2314,N_2389);
and U2510 (N_2510,N_2308,N_2339);
nand U2511 (N_2511,N_2312,N_2204);
nand U2512 (N_2512,N_2218,N_2241);
nand U2513 (N_2513,N_2367,N_2221);
xnor U2514 (N_2514,N_2276,N_2346);
nand U2515 (N_2515,N_2241,N_2285);
and U2516 (N_2516,N_2263,N_2236);
xnor U2517 (N_2517,N_2352,N_2209);
or U2518 (N_2518,N_2274,N_2356);
or U2519 (N_2519,N_2365,N_2323);
nor U2520 (N_2520,N_2295,N_2216);
nand U2521 (N_2521,N_2268,N_2347);
nor U2522 (N_2522,N_2275,N_2246);
nor U2523 (N_2523,N_2308,N_2209);
xor U2524 (N_2524,N_2353,N_2276);
and U2525 (N_2525,N_2331,N_2253);
nand U2526 (N_2526,N_2291,N_2321);
nor U2527 (N_2527,N_2326,N_2397);
and U2528 (N_2528,N_2260,N_2267);
xnor U2529 (N_2529,N_2383,N_2279);
nor U2530 (N_2530,N_2220,N_2250);
nor U2531 (N_2531,N_2270,N_2244);
nand U2532 (N_2532,N_2363,N_2384);
and U2533 (N_2533,N_2257,N_2347);
nor U2534 (N_2534,N_2391,N_2224);
nand U2535 (N_2535,N_2255,N_2388);
nor U2536 (N_2536,N_2293,N_2297);
nor U2537 (N_2537,N_2344,N_2295);
nand U2538 (N_2538,N_2388,N_2353);
or U2539 (N_2539,N_2330,N_2269);
nor U2540 (N_2540,N_2209,N_2230);
xnor U2541 (N_2541,N_2283,N_2256);
xor U2542 (N_2542,N_2375,N_2382);
and U2543 (N_2543,N_2338,N_2278);
and U2544 (N_2544,N_2319,N_2370);
nand U2545 (N_2545,N_2316,N_2362);
xnor U2546 (N_2546,N_2347,N_2351);
nor U2547 (N_2547,N_2236,N_2246);
nand U2548 (N_2548,N_2302,N_2305);
and U2549 (N_2549,N_2224,N_2261);
nand U2550 (N_2550,N_2243,N_2298);
and U2551 (N_2551,N_2231,N_2259);
nand U2552 (N_2552,N_2299,N_2267);
and U2553 (N_2553,N_2279,N_2342);
or U2554 (N_2554,N_2200,N_2333);
or U2555 (N_2555,N_2324,N_2245);
xnor U2556 (N_2556,N_2274,N_2230);
xnor U2557 (N_2557,N_2317,N_2375);
xnor U2558 (N_2558,N_2210,N_2363);
xnor U2559 (N_2559,N_2256,N_2356);
and U2560 (N_2560,N_2287,N_2349);
or U2561 (N_2561,N_2328,N_2258);
xnor U2562 (N_2562,N_2259,N_2325);
nand U2563 (N_2563,N_2221,N_2230);
and U2564 (N_2564,N_2385,N_2390);
xor U2565 (N_2565,N_2218,N_2387);
and U2566 (N_2566,N_2310,N_2369);
or U2567 (N_2567,N_2325,N_2237);
xnor U2568 (N_2568,N_2390,N_2212);
xnor U2569 (N_2569,N_2364,N_2341);
nand U2570 (N_2570,N_2322,N_2248);
or U2571 (N_2571,N_2354,N_2298);
or U2572 (N_2572,N_2203,N_2271);
or U2573 (N_2573,N_2274,N_2270);
and U2574 (N_2574,N_2264,N_2227);
or U2575 (N_2575,N_2381,N_2294);
xnor U2576 (N_2576,N_2371,N_2290);
and U2577 (N_2577,N_2281,N_2313);
nor U2578 (N_2578,N_2231,N_2355);
nand U2579 (N_2579,N_2293,N_2386);
and U2580 (N_2580,N_2398,N_2396);
xor U2581 (N_2581,N_2321,N_2397);
nand U2582 (N_2582,N_2229,N_2399);
xnor U2583 (N_2583,N_2224,N_2383);
nand U2584 (N_2584,N_2382,N_2215);
or U2585 (N_2585,N_2267,N_2310);
or U2586 (N_2586,N_2274,N_2238);
nor U2587 (N_2587,N_2338,N_2299);
and U2588 (N_2588,N_2375,N_2311);
nor U2589 (N_2589,N_2375,N_2248);
and U2590 (N_2590,N_2387,N_2382);
and U2591 (N_2591,N_2302,N_2237);
nor U2592 (N_2592,N_2314,N_2296);
or U2593 (N_2593,N_2284,N_2279);
and U2594 (N_2594,N_2390,N_2247);
xnor U2595 (N_2595,N_2374,N_2390);
or U2596 (N_2596,N_2241,N_2397);
xor U2597 (N_2597,N_2234,N_2330);
xnor U2598 (N_2598,N_2354,N_2359);
and U2599 (N_2599,N_2255,N_2234);
or U2600 (N_2600,N_2593,N_2545);
or U2601 (N_2601,N_2410,N_2599);
or U2602 (N_2602,N_2526,N_2565);
xnor U2603 (N_2603,N_2562,N_2552);
nand U2604 (N_2604,N_2491,N_2409);
xor U2605 (N_2605,N_2447,N_2589);
nand U2606 (N_2606,N_2452,N_2448);
and U2607 (N_2607,N_2595,N_2548);
or U2608 (N_2608,N_2551,N_2489);
or U2609 (N_2609,N_2482,N_2594);
and U2610 (N_2610,N_2454,N_2403);
nor U2611 (N_2611,N_2461,N_2525);
nand U2612 (N_2612,N_2431,N_2458);
nand U2613 (N_2613,N_2439,N_2527);
xnor U2614 (N_2614,N_2467,N_2472);
and U2615 (N_2615,N_2494,N_2484);
nor U2616 (N_2616,N_2578,N_2407);
xor U2617 (N_2617,N_2580,N_2419);
nor U2618 (N_2618,N_2415,N_2501);
or U2619 (N_2619,N_2550,N_2518);
and U2620 (N_2620,N_2468,N_2413);
and U2621 (N_2621,N_2505,N_2490);
nor U2622 (N_2622,N_2576,N_2441);
xor U2623 (N_2623,N_2449,N_2426);
or U2624 (N_2624,N_2586,N_2561);
and U2625 (N_2625,N_2559,N_2404);
nor U2626 (N_2626,N_2569,N_2411);
nand U2627 (N_2627,N_2555,N_2408);
nor U2628 (N_2628,N_2572,N_2495);
and U2629 (N_2629,N_2420,N_2522);
or U2630 (N_2630,N_2573,N_2498);
nor U2631 (N_2631,N_2481,N_2438);
nand U2632 (N_2632,N_2584,N_2570);
nand U2633 (N_2633,N_2523,N_2462);
or U2634 (N_2634,N_2400,N_2473);
and U2635 (N_2635,N_2470,N_2566);
or U2636 (N_2636,N_2549,N_2471);
or U2637 (N_2637,N_2487,N_2567);
nand U2638 (N_2638,N_2590,N_2493);
or U2639 (N_2639,N_2503,N_2424);
xnor U2640 (N_2640,N_2564,N_2581);
nor U2641 (N_2641,N_2453,N_2416);
nor U2642 (N_2642,N_2516,N_2577);
or U2643 (N_2643,N_2583,N_2457);
xor U2644 (N_2644,N_2427,N_2499);
or U2645 (N_2645,N_2543,N_2492);
or U2646 (N_2646,N_2460,N_2451);
nand U2647 (N_2647,N_2558,N_2456);
nor U2648 (N_2648,N_2515,N_2496);
nand U2649 (N_2649,N_2446,N_2519);
nor U2650 (N_2650,N_2469,N_2497);
or U2651 (N_2651,N_2588,N_2571);
or U2652 (N_2652,N_2546,N_2510);
nand U2653 (N_2653,N_2429,N_2463);
or U2654 (N_2654,N_2575,N_2402);
xnor U2655 (N_2655,N_2412,N_2435);
and U2656 (N_2656,N_2440,N_2421);
xor U2657 (N_2657,N_2553,N_2433);
xnor U2658 (N_2658,N_2479,N_2459);
or U2659 (N_2659,N_2432,N_2537);
xnor U2660 (N_2660,N_2574,N_2596);
and U2661 (N_2661,N_2541,N_2414);
and U2662 (N_2662,N_2587,N_2428);
nor U2663 (N_2663,N_2557,N_2512);
nor U2664 (N_2664,N_2520,N_2423);
nor U2665 (N_2665,N_2538,N_2568);
xnor U2666 (N_2666,N_2442,N_2436);
or U2667 (N_2667,N_2475,N_2401);
and U2668 (N_2668,N_2425,N_2560);
or U2669 (N_2669,N_2486,N_2539);
nor U2670 (N_2670,N_2466,N_2465);
nor U2671 (N_2671,N_2508,N_2450);
or U2672 (N_2672,N_2511,N_2464);
and U2673 (N_2673,N_2502,N_2544);
xor U2674 (N_2674,N_2422,N_2532);
nor U2675 (N_2675,N_2524,N_2478);
nor U2676 (N_2676,N_2536,N_2514);
or U2677 (N_2677,N_2504,N_2488);
and U2678 (N_2678,N_2513,N_2474);
and U2679 (N_2679,N_2542,N_2563);
nor U2680 (N_2680,N_2591,N_2579);
nand U2681 (N_2681,N_2476,N_2418);
or U2682 (N_2682,N_2554,N_2437);
xnor U2683 (N_2683,N_2443,N_2506);
xnor U2684 (N_2684,N_2477,N_2434);
nand U2685 (N_2685,N_2405,N_2535);
or U2686 (N_2686,N_2417,N_2455);
nor U2687 (N_2687,N_2547,N_2585);
or U2688 (N_2688,N_2500,N_2521);
nand U2689 (N_2689,N_2540,N_2530);
nand U2690 (N_2690,N_2531,N_2485);
nand U2691 (N_2691,N_2598,N_2430);
or U2692 (N_2692,N_2597,N_2483);
nand U2693 (N_2693,N_2444,N_2592);
and U2694 (N_2694,N_2528,N_2445);
xor U2695 (N_2695,N_2480,N_2507);
and U2696 (N_2696,N_2406,N_2582);
or U2697 (N_2697,N_2517,N_2534);
or U2698 (N_2698,N_2533,N_2529);
or U2699 (N_2699,N_2556,N_2509);
nor U2700 (N_2700,N_2505,N_2596);
or U2701 (N_2701,N_2421,N_2404);
or U2702 (N_2702,N_2599,N_2558);
nor U2703 (N_2703,N_2522,N_2471);
xnor U2704 (N_2704,N_2497,N_2517);
nor U2705 (N_2705,N_2593,N_2592);
or U2706 (N_2706,N_2434,N_2500);
xnor U2707 (N_2707,N_2474,N_2524);
xnor U2708 (N_2708,N_2456,N_2509);
xor U2709 (N_2709,N_2575,N_2520);
xor U2710 (N_2710,N_2419,N_2583);
or U2711 (N_2711,N_2504,N_2571);
nand U2712 (N_2712,N_2570,N_2526);
nor U2713 (N_2713,N_2562,N_2432);
nor U2714 (N_2714,N_2501,N_2497);
nor U2715 (N_2715,N_2502,N_2587);
and U2716 (N_2716,N_2461,N_2531);
and U2717 (N_2717,N_2443,N_2400);
and U2718 (N_2718,N_2537,N_2573);
nand U2719 (N_2719,N_2445,N_2489);
and U2720 (N_2720,N_2510,N_2483);
or U2721 (N_2721,N_2444,N_2482);
nand U2722 (N_2722,N_2419,N_2412);
and U2723 (N_2723,N_2403,N_2590);
xnor U2724 (N_2724,N_2438,N_2429);
xnor U2725 (N_2725,N_2514,N_2590);
xnor U2726 (N_2726,N_2508,N_2453);
or U2727 (N_2727,N_2467,N_2441);
and U2728 (N_2728,N_2415,N_2539);
nor U2729 (N_2729,N_2475,N_2542);
nor U2730 (N_2730,N_2437,N_2508);
nor U2731 (N_2731,N_2434,N_2575);
nand U2732 (N_2732,N_2533,N_2541);
xnor U2733 (N_2733,N_2555,N_2526);
nor U2734 (N_2734,N_2544,N_2435);
xor U2735 (N_2735,N_2572,N_2452);
nand U2736 (N_2736,N_2494,N_2549);
xor U2737 (N_2737,N_2471,N_2556);
xnor U2738 (N_2738,N_2595,N_2530);
xor U2739 (N_2739,N_2495,N_2425);
nor U2740 (N_2740,N_2424,N_2426);
nor U2741 (N_2741,N_2466,N_2446);
nor U2742 (N_2742,N_2439,N_2517);
xor U2743 (N_2743,N_2587,N_2452);
or U2744 (N_2744,N_2577,N_2427);
nand U2745 (N_2745,N_2549,N_2520);
and U2746 (N_2746,N_2571,N_2545);
or U2747 (N_2747,N_2421,N_2408);
nand U2748 (N_2748,N_2542,N_2506);
xor U2749 (N_2749,N_2488,N_2424);
and U2750 (N_2750,N_2478,N_2569);
or U2751 (N_2751,N_2561,N_2537);
nor U2752 (N_2752,N_2437,N_2441);
nand U2753 (N_2753,N_2450,N_2410);
nor U2754 (N_2754,N_2566,N_2527);
nand U2755 (N_2755,N_2486,N_2592);
and U2756 (N_2756,N_2526,N_2411);
and U2757 (N_2757,N_2403,N_2467);
nand U2758 (N_2758,N_2590,N_2431);
nand U2759 (N_2759,N_2443,N_2565);
nand U2760 (N_2760,N_2560,N_2496);
or U2761 (N_2761,N_2571,N_2579);
nand U2762 (N_2762,N_2544,N_2413);
nor U2763 (N_2763,N_2560,N_2499);
or U2764 (N_2764,N_2478,N_2424);
and U2765 (N_2765,N_2491,N_2576);
xnor U2766 (N_2766,N_2528,N_2565);
nand U2767 (N_2767,N_2546,N_2400);
or U2768 (N_2768,N_2496,N_2446);
xnor U2769 (N_2769,N_2430,N_2408);
nor U2770 (N_2770,N_2417,N_2403);
xnor U2771 (N_2771,N_2580,N_2511);
or U2772 (N_2772,N_2520,N_2478);
xnor U2773 (N_2773,N_2573,N_2546);
and U2774 (N_2774,N_2586,N_2575);
or U2775 (N_2775,N_2406,N_2487);
nor U2776 (N_2776,N_2524,N_2597);
and U2777 (N_2777,N_2539,N_2495);
xnor U2778 (N_2778,N_2482,N_2529);
nor U2779 (N_2779,N_2480,N_2526);
nor U2780 (N_2780,N_2552,N_2432);
or U2781 (N_2781,N_2437,N_2504);
nor U2782 (N_2782,N_2487,N_2575);
nor U2783 (N_2783,N_2404,N_2593);
or U2784 (N_2784,N_2416,N_2564);
and U2785 (N_2785,N_2464,N_2460);
nand U2786 (N_2786,N_2407,N_2406);
xor U2787 (N_2787,N_2493,N_2463);
nor U2788 (N_2788,N_2434,N_2409);
and U2789 (N_2789,N_2474,N_2463);
xnor U2790 (N_2790,N_2573,N_2496);
nor U2791 (N_2791,N_2563,N_2515);
nor U2792 (N_2792,N_2484,N_2497);
nor U2793 (N_2793,N_2496,N_2444);
or U2794 (N_2794,N_2487,N_2531);
xnor U2795 (N_2795,N_2585,N_2439);
xor U2796 (N_2796,N_2477,N_2547);
or U2797 (N_2797,N_2441,N_2454);
and U2798 (N_2798,N_2569,N_2500);
nor U2799 (N_2799,N_2518,N_2509);
xor U2800 (N_2800,N_2710,N_2713);
and U2801 (N_2801,N_2665,N_2682);
and U2802 (N_2802,N_2783,N_2745);
xnor U2803 (N_2803,N_2630,N_2676);
xor U2804 (N_2804,N_2709,N_2668);
and U2805 (N_2805,N_2723,N_2692);
xnor U2806 (N_2806,N_2769,N_2689);
nor U2807 (N_2807,N_2628,N_2667);
nand U2808 (N_2808,N_2712,N_2655);
xnor U2809 (N_2809,N_2766,N_2660);
xor U2810 (N_2810,N_2601,N_2677);
and U2811 (N_2811,N_2695,N_2728);
and U2812 (N_2812,N_2654,N_2619);
and U2813 (N_2813,N_2672,N_2618);
nor U2814 (N_2814,N_2636,N_2798);
nand U2815 (N_2815,N_2652,N_2678);
and U2816 (N_2816,N_2604,N_2733);
or U2817 (N_2817,N_2686,N_2658);
or U2818 (N_2818,N_2694,N_2736);
or U2819 (N_2819,N_2623,N_2620);
nor U2820 (N_2820,N_2747,N_2753);
xor U2821 (N_2821,N_2663,N_2740);
nand U2822 (N_2822,N_2696,N_2603);
nor U2823 (N_2823,N_2775,N_2719);
nor U2824 (N_2824,N_2782,N_2635);
nor U2825 (N_2825,N_2792,N_2629);
xnor U2826 (N_2826,N_2602,N_2738);
nand U2827 (N_2827,N_2790,N_2780);
or U2828 (N_2828,N_2606,N_2731);
xor U2829 (N_2829,N_2743,N_2679);
xnor U2830 (N_2830,N_2729,N_2772);
and U2831 (N_2831,N_2681,N_2750);
xnor U2832 (N_2832,N_2730,N_2761);
nor U2833 (N_2833,N_2627,N_2700);
nand U2834 (N_2834,N_2645,N_2758);
nor U2835 (N_2835,N_2771,N_2639);
or U2836 (N_2836,N_2787,N_2659);
and U2837 (N_2837,N_2615,N_2774);
and U2838 (N_2838,N_2680,N_2637);
nand U2839 (N_2839,N_2687,N_2647);
xnor U2840 (N_2840,N_2773,N_2794);
nor U2841 (N_2841,N_2751,N_2724);
nand U2842 (N_2842,N_2718,N_2644);
and U2843 (N_2843,N_2742,N_2748);
and U2844 (N_2844,N_2690,N_2737);
nand U2845 (N_2845,N_2779,N_2674);
nor U2846 (N_2846,N_2610,N_2664);
or U2847 (N_2847,N_2617,N_2714);
nor U2848 (N_2848,N_2757,N_2756);
nand U2849 (N_2849,N_2622,N_2614);
nand U2850 (N_2850,N_2781,N_2691);
and U2851 (N_2851,N_2607,N_2760);
or U2852 (N_2852,N_2651,N_2799);
nor U2853 (N_2853,N_2693,N_2685);
and U2854 (N_2854,N_2697,N_2626);
nand U2855 (N_2855,N_2784,N_2721);
nor U2856 (N_2856,N_2778,N_2708);
xor U2857 (N_2857,N_2722,N_2767);
nand U2858 (N_2858,N_2649,N_2749);
nand U2859 (N_2859,N_2641,N_2765);
or U2860 (N_2860,N_2666,N_2701);
and U2861 (N_2861,N_2707,N_2763);
xor U2862 (N_2862,N_2777,N_2640);
xor U2863 (N_2863,N_2702,N_2705);
and U2864 (N_2864,N_2633,N_2785);
xor U2865 (N_2865,N_2616,N_2726);
nor U2866 (N_2866,N_2762,N_2706);
or U2867 (N_2867,N_2795,N_2643);
nand U2868 (N_2868,N_2716,N_2662);
nand U2869 (N_2869,N_2770,N_2791);
or U2870 (N_2870,N_2638,N_2609);
xor U2871 (N_2871,N_2684,N_2683);
nand U2872 (N_2872,N_2711,N_2656);
or U2873 (N_2873,N_2631,N_2648);
nand U2874 (N_2874,N_2739,N_2642);
nand U2875 (N_2875,N_2734,N_2746);
nor U2876 (N_2876,N_2725,N_2669);
and U2877 (N_2877,N_2625,N_2797);
xnor U2878 (N_2878,N_2788,N_2650);
or U2879 (N_2879,N_2624,N_2698);
nand U2880 (N_2880,N_2673,N_2600);
nor U2881 (N_2881,N_2661,N_2612);
nand U2882 (N_2882,N_2670,N_2675);
nand U2883 (N_2883,N_2764,N_2621);
and U2884 (N_2884,N_2793,N_2755);
or U2885 (N_2885,N_2717,N_2754);
xnor U2886 (N_2886,N_2752,N_2703);
and U2887 (N_2887,N_2786,N_2735);
and U2888 (N_2888,N_2720,N_2727);
nor U2889 (N_2889,N_2759,N_2796);
or U2890 (N_2890,N_2768,N_2732);
nand U2891 (N_2891,N_2744,N_2657);
nand U2892 (N_2892,N_2699,N_2646);
and U2893 (N_2893,N_2671,N_2653);
and U2894 (N_2894,N_2632,N_2608);
and U2895 (N_2895,N_2776,N_2605);
nand U2896 (N_2896,N_2704,N_2741);
or U2897 (N_2897,N_2715,N_2634);
xor U2898 (N_2898,N_2688,N_2613);
and U2899 (N_2899,N_2611,N_2789);
xnor U2900 (N_2900,N_2652,N_2748);
nor U2901 (N_2901,N_2773,N_2717);
and U2902 (N_2902,N_2674,N_2740);
or U2903 (N_2903,N_2755,N_2645);
or U2904 (N_2904,N_2712,N_2757);
nand U2905 (N_2905,N_2635,N_2690);
nor U2906 (N_2906,N_2713,N_2693);
nor U2907 (N_2907,N_2662,N_2675);
or U2908 (N_2908,N_2738,N_2659);
or U2909 (N_2909,N_2742,N_2657);
and U2910 (N_2910,N_2680,N_2666);
xor U2911 (N_2911,N_2767,N_2601);
nor U2912 (N_2912,N_2659,N_2770);
or U2913 (N_2913,N_2657,N_2723);
and U2914 (N_2914,N_2651,N_2760);
nor U2915 (N_2915,N_2795,N_2744);
nor U2916 (N_2916,N_2676,N_2687);
or U2917 (N_2917,N_2619,N_2655);
nor U2918 (N_2918,N_2710,N_2622);
or U2919 (N_2919,N_2681,N_2716);
nand U2920 (N_2920,N_2767,N_2723);
and U2921 (N_2921,N_2637,N_2673);
nor U2922 (N_2922,N_2698,N_2792);
nor U2923 (N_2923,N_2694,N_2628);
nand U2924 (N_2924,N_2752,N_2741);
nor U2925 (N_2925,N_2701,N_2615);
and U2926 (N_2926,N_2752,N_2734);
nor U2927 (N_2927,N_2627,N_2778);
nand U2928 (N_2928,N_2641,N_2680);
or U2929 (N_2929,N_2730,N_2720);
nor U2930 (N_2930,N_2656,N_2640);
or U2931 (N_2931,N_2660,N_2736);
and U2932 (N_2932,N_2733,N_2699);
xnor U2933 (N_2933,N_2743,N_2687);
xor U2934 (N_2934,N_2789,N_2790);
xor U2935 (N_2935,N_2646,N_2645);
nand U2936 (N_2936,N_2679,N_2670);
or U2937 (N_2937,N_2757,N_2669);
nor U2938 (N_2938,N_2754,N_2641);
and U2939 (N_2939,N_2700,N_2798);
nand U2940 (N_2940,N_2713,N_2679);
and U2941 (N_2941,N_2684,N_2643);
nand U2942 (N_2942,N_2674,N_2650);
nand U2943 (N_2943,N_2795,N_2678);
or U2944 (N_2944,N_2781,N_2684);
nor U2945 (N_2945,N_2716,N_2612);
nor U2946 (N_2946,N_2785,N_2792);
nand U2947 (N_2947,N_2734,N_2666);
or U2948 (N_2948,N_2731,N_2773);
or U2949 (N_2949,N_2723,N_2682);
or U2950 (N_2950,N_2635,N_2748);
or U2951 (N_2951,N_2746,N_2764);
and U2952 (N_2952,N_2790,N_2600);
nand U2953 (N_2953,N_2687,N_2620);
nand U2954 (N_2954,N_2644,N_2768);
nand U2955 (N_2955,N_2755,N_2743);
or U2956 (N_2956,N_2665,N_2793);
xnor U2957 (N_2957,N_2761,N_2785);
nor U2958 (N_2958,N_2687,N_2649);
nand U2959 (N_2959,N_2630,N_2704);
nor U2960 (N_2960,N_2637,N_2712);
nor U2961 (N_2961,N_2630,N_2795);
and U2962 (N_2962,N_2726,N_2648);
xnor U2963 (N_2963,N_2661,N_2647);
or U2964 (N_2964,N_2677,N_2689);
and U2965 (N_2965,N_2700,N_2674);
nor U2966 (N_2966,N_2609,N_2664);
nand U2967 (N_2967,N_2603,N_2778);
or U2968 (N_2968,N_2685,N_2752);
nor U2969 (N_2969,N_2764,N_2680);
or U2970 (N_2970,N_2676,N_2626);
nor U2971 (N_2971,N_2681,N_2627);
xor U2972 (N_2972,N_2678,N_2620);
nor U2973 (N_2973,N_2745,N_2613);
nand U2974 (N_2974,N_2699,N_2630);
nand U2975 (N_2975,N_2719,N_2627);
nor U2976 (N_2976,N_2641,N_2600);
xnor U2977 (N_2977,N_2675,N_2613);
and U2978 (N_2978,N_2647,N_2703);
xnor U2979 (N_2979,N_2762,N_2615);
and U2980 (N_2980,N_2675,N_2699);
nand U2981 (N_2981,N_2634,N_2790);
or U2982 (N_2982,N_2768,N_2600);
nor U2983 (N_2983,N_2748,N_2712);
nand U2984 (N_2984,N_2750,N_2610);
and U2985 (N_2985,N_2630,N_2789);
and U2986 (N_2986,N_2728,N_2683);
or U2987 (N_2987,N_2602,N_2785);
nor U2988 (N_2988,N_2724,N_2720);
or U2989 (N_2989,N_2737,N_2654);
and U2990 (N_2990,N_2724,N_2713);
and U2991 (N_2991,N_2701,N_2785);
xor U2992 (N_2992,N_2729,N_2605);
nor U2993 (N_2993,N_2758,N_2631);
nor U2994 (N_2994,N_2753,N_2696);
nor U2995 (N_2995,N_2720,N_2798);
and U2996 (N_2996,N_2687,N_2757);
nor U2997 (N_2997,N_2618,N_2647);
nand U2998 (N_2998,N_2638,N_2786);
nand U2999 (N_2999,N_2718,N_2634);
xor U3000 (N_3000,N_2829,N_2917);
nor U3001 (N_3001,N_2872,N_2969);
nand U3002 (N_3002,N_2813,N_2855);
or U3003 (N_3003,N_2819,N_2884);
and U3004 (N_3004,N_2853,N_2898);
nor U3005 (N_3005,N_2802,N_2804);
xor U3006 (N_3006,N_2998,N_2939);
or U3007 (N_3007,N_2970,N_2907);
xor U3008 (N_3008,N_2833,N_2883);
xor U3009 (N_3009,N_2921,N_2910);
nand U3010 (N_3010,N_2942,N_2912);
and U3011 (N_3011,N_2963,N_2977);
xnor U3012 (N_3012,N_2874,N_2827);
nor U3013 (N_3013,N_2806,N_2941);
and U3014 (N_3014,N_2885,N_2914);
xnor U3015 (N_3015,N_2945,N_2851);
or U3016 (N_3016,N_2926,N_2864);
and U3017 (N_3017,N_2915,N_2821);
or U3018 (N_3018,N_2899,N_2920);
and U3019 (N_3019,N_2956,N_2893);
and U3020 (N_3020,N_2801,N_2830);
nor U3021 (N_3021,N_2814,N_2937);
or U3022 (N_3022,N_2900,N_2820);
nor U3023 (N_3023,N_2960,N_2940);
and U3024 (N_3024,N_2894,N_2927);
or U3025 (N_3025,N_2984,N_2962);
xor U3026 (N_3026,N_2825,N_2880);
or U3027 (N_3027,N_2958,N_2892);
nor U3028 (N_3028,N_2965,N_2913);
nor U3029 (N_3029,N_2952,N_2961);
xnor U3030 (N_3030,N_2988,N_2909);
xnor U3031 (N_3031,N_2986,N_2863);
and U3032 (N_3032,N_2826,N_2861);
nand U3033 (N_3033,N_2800,N_2867);
nand U3034 (N_3034,N_2878,N_2823);
or U3035 (N_3035,N_2886,N_2870);
or U3036 (N_3036,N_2879,N_2957);
nand U3037 (N_3037,N_2871,N_2887);
nand U3038 (N_3038,N_2818,N_2889);
nor U3039 (N_3039,N_2866,N_2842);
nand U3040 (N_3040,N_2891,N_2888);
nand U3041 (N_3041,N_2896,N_2934);
and U3042 (N_3042,N_2944,N_2999);
xnor U3043 (N_3043,N_2938,N_2935);
and U3044 (N_3044,N_2950,N_2906);
nor U3045 (N_3045,N_2990,N_2845);
or U3046 (N_3046,N_2955,N_2875);
xnor U3047 (N_3047,N_2876,N_2859);
nand U3048 (N_3048,N_2862,N_2811);
or U3049 (N_3049,N_2837,N_2930);
and U3050 (N_3050,N_2865,N_2897);
xor U3051 (N_3051,N_2996,N_2985);
nor U3052 (N_3052,N_2929,N_2953);
and U3053 (N_3053,N_2847,N_2951);
nand U3054 (N_3054,N_2994,N_2860);
nor U3055 (N_3055,N_2980,N_2931);
nor U3056 (N_3056,N_2982,N_2828);
xor U3057 (N_3057,N_2908,N_2835);
or U3058 (N_3058,N_2848,N_2815);
xnor U3059 (N_3059,N_2895,N_2803);
and U3060 (N_3060,N_2831,N_2844);
xnor U3061 (N_3061,N_2822,N_2839);
and U3062 (N_3062,N_2810,N_2974);
nor U3063 (N_3063,N_2904,N_2809);
or U3064 (N_3064,N_2911,N_2949);
or U3065 (N_3065,N_2902,N_2946);
or U3066 (N_3066,N_2983,N_2971);
and U3067 (N_3067,N_2916,N_2840);
nand U3068 (N_3068,N_2943,N_2868);
xor U3069 (N_3069,N_2975,N_2841);
xnor U3070 (N_3070,N_2993,N_2838);
and U3071 (N_3071,N_2881,N_2852);
nor U3072 (N_3072,N_2846,N_2924);
or U3073 (N_3073,N_2903,N_2901);
nand U3074 (N_3074,N_2997,N_2850);
nor U3075 (N_3075,N_2925,N_2869);
and U3076 (N_3076,N_2948,N_2824);
nor U3077 (N_3077,N_2817,N_2857);
nor U3078 (N_3078,N_2976,N_2981);
or U3079 (N_3079,N_2807,N_2967);
xor U3080 (N_3080,N_2964,N_2922);
xnor U3081 (N_3081,N_2873,N_2858);
and U3082 (N_3082,N_2812,N_2890);
or U3083 (N_3083,N_2834,N_2954);
nor U3084 (N_3084,N_2808,N_2995);
xor U3085 (N_3085,N_2966,N_2849);
and U3086 (N_3086,N_2991,N_2968);
or U3087 (N_3087,N_2856,N_2973);
nand U3088 (N_3088,N_2843,N_2989);
and U3089 (N_3089,N_2854,N_2992);
nand U3090 (N_3090,N_2972,N_2918);
nand U3091 (N_3091,N_2936,N_2905);
nand U3092 (N_3092,N_2959,N_2923);
xnor U3093 (N_3093,N_2933,N_2947);
nor U3094 (N_3094,N_2877,N_2805);
and U3095 (N_3095,N_2882,N_2932);
nand U3096 (N_3096,N_2987,N_2816);
or U3097 (N_3097,N_2919,N_2978);
nor U3098 (N_3098,N_2979,N_2832);
nand U3099 (N_3099,N_2836,N_2928);
xnor U3100 (N_3100,N_2877,N_2826);
nor U3101 (N_3101,N_2801,N_2989);
nand U3102 (N_3102,N_2847,N_2998);
nand U3103 (N_3103,N_2800,N_2841);
and U3104 (N_3104,N_2927,N_2993);
or U3105 (N_3105,N_2881,N_2907);
or U3106 (N_3106,N_2820,N_2942);
or U3107 (N_3107,N_2917,N_2913);
nand U3108 (N_3108,N_2869,N_2853);
nor U3109 (N_3109,N_2817,N_2871);
or U3110 (N_3110,N_2923,N_2969);
and U3111 (N_3111,N_2803,N_2964);
nand U3112 (N_3112,N_2991,N_2802);
xor U3113 (N_3113,N_2959,N_2817);
nor U3114 (N_3114,N_2885,N_2828);
xnor U3115 (N_3115,N_2876,N_2847);
xnor U3116 (N_3116,N_2983,N_2814);
xnor U3117 (N_3117,N_2869,N_2910);
nand U3118 (N_3118,N_2864,N_2824);
nand U3119 (N_3119,N_2931,N_2825);
nand U3120 (N_3120,N_2958,N_2977);
nand U3121 (N_3121,N_2910,N_2857);
or U3122 (N_3122,N_2862,N_2917);
and U3123 (N_3123,N_2826,N_2909);
nand U3124 (N_3124,N_2979,N_2982);
nand U3125 (N_3125,N_2913,N_2959);
and U3126 (N_3126,N_2921,N_2954);
and U3127 (N_3127,N_2859,N_2822);
xnor U3128 (N_3128,N_2992,N_2940);
xor U3129 (N_3129,N_2987,N_2925);
and U3130 (N_3130,N_2801,N_2869);
nor U3131 (N_3131,N_2864,N_2898);
nor U3132 (N_3132,N_2837,N_2892);
nand U3133 (N_3133,N_2813,N_2953);
nor U3134 (N_3134,N_2827,N_2965);
or U3135 (N_3135,N_2882,N_2837);
and U3136 (N_3136,N_2973,N_2927);
nand U3137 (N_3137,N_2901,N_2888);
and U3138 (N_3138,N_2875,N_2900);
nand U3139 (N_3139,N_2987,N_2968);
nor U3140 (N_3140,N_2902,N_2880);
or U3141 (N_3141,N_2827,N_2961);
or U3142 (N_3142,N_2978,N_2965);
nand U3143 (N_3143,N_2948,N_2972);
nor U3144 (N_3144,N_2992,N_2826);
xor U3145 (N_3145,N_2836,N_2894);
nand U3146 (N_3146,N_2917,N_2908);
xor U3147 (N_3147,N_2989,N_2962);
and U3148 (N_3148,N_2849,N_2875);
or U3149 (N_3149,N_2974,N_2905);
nor U3150 (N_3150,N_2993,N_2978);
nand U3151 (N_3151,N_2836,N_2846);
nor U3152 (N_3152,N_2935,N_2819);
nor U3153 (N_3153,N_2937,N_2989);
nor U3154 (N_3154,N_2836,N_2908);
xnor U3155 (N_3155,N_2842,N_2913);
nand U3156 (N_3156,N_2884,N_2975);
nor U3157 (N_3157,N_2812,N_2937);
nor U3158 (N_3158,N_2944,N_2860);
and U3159 (N_3159,N_2874,N_2902);
and U3160 (N_3160,N_2957,N_2995);
xnor U3161 (N_3161,N_2917,N_2929);
xnor U3162 (N_3162,N_2984,N_2982);
nor U3163 (N_3163,N_2843,N_2844);
and U3164 (N_3164,N_2915,N_2886);
and U3165 (N_3165,N_2926,N_2845);
xor U3166 (N_3166,N_2971,N_2925);
nand U3167 (N_3167,N_2837,N_2813);
xor U3168 (N_3168,N_2881,N_2898);
or U3169 (N_3169,N_2892,N_2826);
nor U3170 (N_3170,N_2921,N_2869);
or U3171 (N_3171,N_2997,N_2813);
xor U3172 (N_3172,N_2877,N_2992);
nor U3173 (N_3173,N_2833,N_2933);
nand U3174 (N_3174,N_2962,N_2936);
nand U3175 (N_3175,N_2805,N_2913);
xnor U3176 (N_3176,N_2991,N_2976);
or U3177 (N_3177,N_2819,N_2994);
nand U3178 (N_3178,N_2968,N_2871);
xor U3179 (N_3179,N_2884,N_2843);
nand U3180 (N_3180,N_2866,N_2924);
nor U3181 (N_3181,N_2972,N_2928);
or U3182 (N_3182,N_2802,N_2824);
and U3183 (N_3183,N_2872,N_2935);
nor U3184 (N_3184,N_2906,N_2867);
nor U3185 (N_3185,N_2804,N_2864);
nand U3186 (N_3186,N_2986,N_2857);
xor U3187 (N_3187,N_2936,N_2874);
nand U3188 (N_3188,N_2857,N_2942);
nand U3189 (N_3189,N_2885,N_2834);
nor U3190 (N_3190,N_2845,N_2832);
and U3191 (N_3191,N_2883,N_2871);
and U3192 (N_3192,N_2909,N_2911);
nor U3193 (N_3193,N_2810,N_2923);
xnor U3194 (N_3194,N_2985,N_2920);
or U3195 (N_3195,N_2800,N_2929);
nor U3196 (N_3196,N_2857,N_2893);
or U3197 (N_3197,N_2802,N_2890);
xnor U3198 (N_3198,N_2967,N_2924);
nor U3199 (N_3199,N_2918,N_2839);
and U3200 (N_3200,N_3117,N_3073);
nor U3201 (N_3201,N_3199,N_3029);
xor U3202 (N_3202,N_3115,N_3037);
nor U3203 (N_3203,N_3017,N_3054);
xnor U3204 (N_3204,N_3109,N_3013);
or U3205 (N_3205,N_3153,N_3105);
and U3206 (N_3206,N_3043,N_3044);
and U3207 (N_3207,N_3072,N_3078);
nand U3208 (N_3208,N_3141,N_3001);
or U3209 (N_3209,N_3125,N_3147);
or U3210 (N_3210,N_3127,N_3047);
xnor U3211 (N_3211,N_3134,N_3022);
or U3212 (N_3212,N_3002,N_3007);
xor U3213 (N_3213,N_3130,N_3085);
xnor U3214 (N_3214,N_3041,N_3175);
xor U3215 (N_3215,N_3142,N_3031);
nor U3216 (N_3216,N_3066,N_3040);
and U3217 (N_3217,N_3114,N_3116);
xnor U3218 (N_3218,N_3018,N_3124);
or U3219 (N_3219,N_3068,N_3176);
xnor U3220 (N_3220,N_3048,N_3166);
nor U3221 (N_3221,N_3097,N_3046);
xnor U3222 (N_3222,N_3159,N_3064);
or U3223 (N_3223,N_3191,N_3132);
and U3224 (N_3224,N_3179,N_3143);
xnor U3225 (N_3225,N_3107,N_3102);
or U3226 (N_3226,N_3197,N_3069);
xor U3227 (N_3227,N_3186,N_3099);
xnor U3228 (N_3228,N_3056,N_3196);
nand U3229 (N_3229,N_3121,N_3077);
nand U3230 (N_3230,N_3156,N_3023);
xnor U3231 (N_3231,N_3051,N_3188);
nand U3232 (N_3232,N_3015,N_3027);
nor U3233 (N_3233,N_3092,N_3152);
and U3234 (N_3234,N_3157,N_3016);
nor U3235 (N_3235,N_3106,N_3122);
xnor U3236 (N_3236,N_3065,N_3084);
or U3237 (N_3237,N_3062,N_3032);
xor U3238 (N_3238,N_3138,N_3171);
xor U3239 (N_3239,N_3050,N_3111);
nand U3240 (N_3240,N_3093,N_3168);
or U3241 (N_3241,N_3030,N_3104);
or U3242 (N_3242,N_3151,N_3052);
nand U3243 (N_3243,N_3164,N_3079);
xor U3244 (N_3244,N_3160,N_3014);
xor U3245 (N_3245,N_3194,N_3063);
nor U3246 (N_3246,N_3158,N_3169);
nand U3247 (N_3247,N_3140,N_3128);
xor U3248 (N_3248,N_3019,N_3192);
or U3249 (N_3249,N_3036,N_3012);
or U3250 (N_3250,N_3163,N_3091);
xnor U3251 (N_3251,N_3006,N_3059);
nor U3252 (N_3252,N_3095,N_3089);
nand U3253 (N_3253,N_3183,N_3120);
xnor U3254 (N_3254,N_3139,N_3113);
or U3255 (N_3255,N_3150,N_3024);
nor U3256 (N_3256,N_3033,N_3080);
xor U3257 (N_3257,N_3060,N_3190);
xnor U3258 (N_3258,N_3090,N_3096);
and U3259 (N_3259,N_3133,N_3049);
and U3260 (N_3260,N_3020,N_3126);
xor U3261 (N_3261,N_3045,N_3061);
nand U3262 (N_3262,N_3123,N_3003);
xnor U3263 (N_3263,N_3181,N_3119);
and U3264 (N_3264,N_3055,N_3101);
xnor U3265 (N_3265,N_3025,N_3081);
and U3266 (N_3266,N_3039,N_3178);
nor U3267 (N_3267,N_3087,N_3144);
and U3268 (N_3268,N_3137,N_3195);
xor U3269 (N_3269,N_3004,N_3034);
nand U3270 (N_3270,N_3110,N_3182);
xor U3271 (N_3271,N_3075,N_3146);
nor U3272 (N_3272,N_3011,N_3057);
or U3273 (N_3273,N_3154,N_3086);
and U3274 (N_3274,N_3162,N_3108);
or U3275 (N_3275,N_3010,N_3155);
or U3276 (N_3276,N_3103,N_3067);
nor U3277 (N_3277,N_3129,N_3167);
or U3278 (N_3278,N_3038,N_3174);
xor U3279 (N_3279,N_3193,N_3149);
and U3280 (N_3280,N_3118,N_3136);
nor U3281 (N_3281,N_3026,N_3094);
nor U3282 (N_3282,N_3100,N_3184);
and U3283 (N_3283,N_3008,N_3042);
or U3284 (N_3284,N_3083,N_3187);
or U3285 (N_3285,N_3145,N_3198);
or U3286 (N_3286,N_3148,N_3172);
nor U3287 (N_3287,N_3185,N_3058);
or U3288 (N_3288,N_3028,N_3165);
and U3289 (N_3289,N_3131,N_3112);
nor U3290 (N_3290,N_3009,N_3161);
and U3291 (N_3291,N_3135,N_3071);
nor U3292 (N_3292,N_3170,N_3082);
and U3293 (N_3293,N_3005,N_3021);
nor U3294 (N_3294,N_3053,N_3189);
nand U3295 (N_3295,N_3098,N_3180);
or U3296 (N_3296,N_3177,N_3070);
xor U3297 (N_3297,N_3088,N_3035);
xor U3298 (N_3298,N_3074,N_3173);
nor U3299 (N_3299,N_3000,N_3076);
or U3300 (N_3300,N_3154,N_3091);
nor U3301 (N_3301,N_3139,N_3167);
or U3302 (N_3302,N_3107,N_3010);
xnor U3303 (N_3303,N_3114,N_3151);
xnor U3304 (N_3304,N_3052,N_3114);
nand U3305 (N_3305,N_3066,N_3002);
or U3306 (N_3306,N_3060,N_3083);
or U3307 (N_3307,N_3066,N_3130);
and U3308 (N_3308,N_3186,N_3122);
and U3309 (N_3309,N_3144,N_3005);
and U3310 (N_3310,N_3088,N_3133);
and U3311 (N_3311,N_3018,N_3096);
xor U3312 (N_3312,N_3155,N_3082);
or U3313 (N_3313,N_3078,N_3168);
xor U3314 (N_3314,N_3039,N_3064);
xnor U3315 (N_3315,N_3072,N_3140);
and U3316 (N_3316,N_3082,N_3098);
nor U3317 (N_3317,N_3154,N_3015);
and U3318 (N_3318,N_3019,N_3193);
or U3319 (N_3319,N_3127,N_3130);
nand U3320 (N_3320,N_3066,N_3144);
xor U3321 (N_3321,N_3139,N_3142);
and U3322 (N_3322,N_3130,N_3136);
and U3323 (N_3323,N_3155,N_3085);
nand U3324 (N_3324,N_3065,N_3129);
and U3325 (N_3325,N_3083,N_3072);
nand U3326 (N_3326,N_3122,N_3013);
and U3327 (N_3327,N_3148,N_3139);
or U3328 (N_3328,N_3092,N_3193);
nor U3329 (N_3329,N_3169,N_3116);
nor U3330 (N_3330,N_3092,N_3147);
or U3331 (N_3331,N_3117,N_3028);
or U3332 (N_3332,N_3126,N_3039);
xor U3333 (N_3333,N_3146,N_3110);
xor U3334 (N_3334,N_3000,N_3171);
nand U3335 (N_3335,N_3014,N_3162);
nor U3336 (N_3336,N_3049,N_3032);
and U3337 (N_3337,N_3039,N_3105);
nand U3338 (N_3338,N_3089,N_3112);
or U3339 (N_3339,N_3101,N_3183);
xor U3340 (N_3340,N_3117,N_3023);
and U3341 (N_3341,N_3021,N_3136);
and U3342 (N_3342,N_3182,N_3186);
and U3343 (N_3343,N_3057,N_3147);
nand U3344 (N_3344,N_3143,N_3033);
and U3345 (N_3345,N_3164,N_3052);
or U3346 (N_3346,N_3021,N_3068);
nand U3347 (N_3347,N_3061,N_3193);
nor U3348 (N_3348,N_3003,N_3066);
nor U3349 (N_3349,N_3062,N_3138);
nand U3350 (N_3350,N_3128,N_3055);
nand U3351 (N_3351,N_3185,N_3042);
nor U3352 (N_3352,N_3004,N_3022);
and U3353 (N_3353,N_3147,N_3120);
or U3354 (N_3354,N_3098,N_3099);
xnor U3355 (N_3355,N_3188,N_3029);
nor U3356 (N_3356,N_3030,N_3110);
nand U3357 (N_3357,N_3178,N_3021);
nor U3358 (N_3358,N_3176,N_3198);
nor U3359 (N_3359,N_3103,N_3127);
xnor U3360 (N_3360,N_3048,N_3181);
nor U3361 (N_3361,N_3077,N_3081);
nor U3362 (N_3362,N_3093,N_3009);
nor U3363 (N_3363,N_3111,N_3010);
xnor U3364 (N_3364,N_3022,N_3112);
nand U3365 (N_3365,N_3068,N_3118);
or U3366 (N_3366,N_3056,N_3137);
nand U3367 (N_3367,N_3149,N_3034);
nand U3368 (N_3368,N_3037,N_3124);
xnor U3369 (N_3369,N_3105,N_3020);
nand U3370 (N_3370,N_3142,N_3198);
nor U3371 (N_3371,N_3097,N_3146);
nor U3372 (N_3372,N_3176,N_3043);
nand U3373 (N_3373,N_3086,N_3127);
xnor U3374 (N_3374,N_3051,N_3109);
and U3375 (N_3375,N_3140,N_3024);
and U3376 (N_3376,N_3044,N_3046);
and U3377 (N_3377,N_3099,N_3021);
xor U3378 (N_3378,N_3109,N_3052);
nor U3379 (N_3379,N_3024,N_3058);
nand U3380 (N_3380,N_3121,N_3148);
and U3381 (N_3381,N_3160,N_3022);
nor U3382 (N_3382,N_3032,N_3043);
and U3383 (N_3383,N_3189,N_3001);
nand U3384 (N_3384,N_3011,N_3092);
or U3385 (N_3385,N_3017,N_3032);
nand U3386 (N_3386,N_3152,N_3015);
nor U3387 (N_3387,N_3112,N_3091);
and U3388 (N_3388,N_3181,N_3140);
nand U3389 (N_3389,N_3109,N_3160);
or U3390 (N_3390,N_3127,N_3192);
nor U3391 (N_3391,N_3100,N_3018);
and U3392 (N_3392,N_3172,N_3054);
nand U3393 (N_3393,N_3109,N_3034);
nand U3394 (N_3394,N_3056,N_3189);
xor U3395 (N_3395,N_3056,N_3021);
or U3396 (N_3396,N_3177,N_3064);
nor U3397 (N_3397,N_3034,N_3140);
xor U3398 (N_3398,N_3160,N_3113);
nor U3399 (N_3399,N_3066,N_3016);
xnor U3400 (N_3400,N_3258,N_3201);
or U3401 (N_3401,N_3226,N_3358);
nor U3402 (N_3402,N_3270,N_3248);
xor U3403 (N_3403,N_3251,N_3368);
nor U3404 (N_3404,N_3213,N_3299);
nor U3405 (N_3405,N_3379,N_3269);
nor U3406 (N_3406,N_3285,N_3264);
xor U3407 (N_3407,N_3217,N_3360);
xor U3408 (N_3408,N_3327,N_3315);
and U3409 (N_3409,N_3393,N_3241);
xnor U3410 (N_3410,N_3203,N_3271);
nand U3411 (N_3411,N_3321,N_3260);
xnor U3412 (N_3412,N_3340,N_3253);
or U3413 (N_3413,N_3345,N_3383);
nand U3414 (N_3414,N_3348,N_3371);
or U3415 (N_3415,N_3233,N_3227);
nand U3416 (N_3416,N_3359,N_3295);
nor U3417 (N_3417,N_3362,N_3218);
xor U3418 (N_3418,N_3377,N_3328);
and U3419 (N_3419,N_3289,N_3354);
or U3420 (N_3420,N_3205,N_3313);
and U3421 (N_3421,N_3386,N_3202);
or U3422 (N_3422,N_3214,N_3223);
nand U3423 (N_3423,N_3231,N_3210);
xnor U3424 (N_3424,N_3265,N_3290);
and U3425 (N_3425,N_3247,N_3366);
and U3426 (N_3426,N_3236,N_3263);
nand U3427 (N_3427,N_3230,N_3318);
xnor U3428 (N_3428,N_3303,N_3261);
xnor U3429 (N_3429,N_3361,N_3376);
xor U3430 (N_3430,N_3279,N_3281);
nor U3431 (N_3431,N_3384,N_3336);
and U3432 (N_3432,N_3391,N_3342);
nor U3433 (N_3433,N_3209,N_3294);
and U3434 (N_3434,N_3287,N_3211);
nor U3435 (N_3435,N_3323,N_3319);
xor U3436 (N_3436,N_3304,N_3351);
or U3437 (N_3437,N_3272,N_3365);
or U3438 (N_3438,N_3375,N_3346);
nor U3439 (N_3439,N_3206,N_3308);
and U3440 (N_3440,N_3274,N_3262);
nand U3441 (N_3441,N_3204,N_3257);
nand U3442 (N_3442,N_3317,N_3284);
nand U3443 (N_3443,N_3301,N_3229);
xor U3444 (N_3444,N_3356,N_3283);
and U3445 (N_3445,N_3390,N_3397);
or U3446 (N_3446,N_3266,N_3286);
and U3447 (N_3447,N_3298,N_3344);
or U3448 (N_3448,N_3350,N_3302);
or U3449 (N_3449,N_3394,N_3228);
nand U3450 (N_3450,N_3341,N_3208);
xnor U3451 (N_3451,N_3332,N_3275);
nor U3452 (N_3452,N_3349,N_3268);
nor U3453 (N_3453,N_3200,N_3291);
or U3454 (N_3454,N_3312,N_3326);
xor U3455 (N_3455,N_3364,N_3259);
or U3456 (N_3456,N_3353,N_3238);
and U3457 (N_3457,N_3355,N_3212);
nand U3458 (N_3458,N_3395,N_3357);
nand U3459 (N_3459,N_3278,N_3282);
and U3460 (N_3460,N_3237,N_3389);
or U3461 (N_3461,N_3370,N_3245);
and U3462 (N_3462,N_3207,N_3378);
nor U3463 (N_3463,N_3273,N_3293);
and U3464 (N_3464,N_3373,N_3335);
or U3465 (N_3465,N_3296,N_3280);
or U3466 (N_3466,N_3325,N_3292);
nand U3467 (N_3467,N_3222,N_3300);
nor U3468 (N_3468,N_3232,N_3329);
xnor U3469 (N_3469,N_3352,N_3255);
or U3470 (N_3470,N_3244,N_3374);
nor U3471 (N_3471,N_3388,N_3322);
xor U3472 (N_3472,N_3220,N_3363);
nand U3473 (N_3473,N_3239,N_3225);
or U3474 (N_3474,N_3399,N_3347);
or U3475 (N_3475,N_3305,N_3216);
nand U3476 (N_3476,N_3235,N_3250);
and U3477 (N_3477,N_3367,N_3398);
xor U3478 (N_3478,N_3339,N_3333);
xnor U3479 (N_3479,N_3249,N_3314);
or U3480 (N_3480,N_3338,N_3320);
and U3481 (N_3481,N_3276,N_3337);
or U3482 (N_3482,N_3254,N_3396);
nor U3483 (N_3483,N_3385,N_3331);
or U3484 (N_3484,N_3369,N_3252);
nand U3485 (N_3485,N_3219,N_3306);
xnor U3486 (N_3486,N_3334,N_3242);
and U3487 (N_3487,N_3224,N_3387);
xor U3488 (N_3488,N_3246,N_3316);
xnor U3489 (N_3489,N_3382,N_3243);
xor U3490 (N_3490,N_3256,N_3288);
nor U3491 (N_3491,N_3297,N_3277);
nor U3492 (N_3492,N_3234,N_3392);
nor U3493 (N_3493,N_3324,N_3311);
and U3494 (N_3494,N_3221,N_3215);
or U3495 (N_3495,N_3372,N_3310);
xnor U3496 (N_3496,N_3307,N_3240);
or U3497 (N_3497,N_3381,N_3343);
nor U3498 (N_3498,N_3309,N_3380);
xor U3499 (N_3499,N_3330,N_3267);
and U3500 (N_3500,N_3382,N_3305);
xor U3501 (N_3501,N_3282,N_3314);
nand U3502 (N_3502,N_3268,N_3363);
or U3503 (N_3503,N_3290,N_3303);
or U3504 (N_3504,N_3289,N_3328);
and U3505 (N_3505,N_3243,N_3208);
xnor U3506 (N_3506,N_3233,N_3355);
and U3507 (N_3507,N_3353,N_3399);
nor U3508 (N_3508,N_3287,N_3338);
nand U3509 (N_3509,N_3318,N_3314);
xnor U3510 (N_3510,N_3289,N_3327);
nor U3511 (N_3511,N_3368,N_3268);
xor U3512 (N_3512,N_3238,N_3294);
xor U3513 (N_3513,N_3349,N_3274);
or U3514 (N_3514,N_3202,N_3342);
xnor U3515 (N_3515,N_3256,N_3344);
and U3516 (N_3516,N_3351,N_3355);
xor U3517 (N_3517,N_3257,N_3322);
nand U3518 (N_3518,N_3295,N_3329);
or U3519 (N_3519,N_3259,N_3317);
or U3520 (N_3520,N_3344,N_3234);
or U3521 (N_3521,N_3275,N_3287);
nand U3522 (N_3522,N_3331,N_3340);
nand U3523 (N_3523,N_3200,N_3239);
xor U3524 (N_3524,N_3283,N_3326);
or U3525 (N_3525,N_3314,N_3295);
or U3526 (N_3526,N_3287,N_3286);
or U3527 (N_3527,N_3210,N_3297);
and U3528 (N_3528,N_3212,N_3301);
or U3529 (N_3529,N_3360,N_3287);
or U3530 (N_3530,N_3203,N_3370);
nor U3531 (N_3531,N_3348,N_3295);
xor U3532 (N_3532,N_3382,N_3201);
or U3533 (N_3533,N_3220,N_3324);
or U3534 (N_3534,N_3220,N_3212);
and U3535 (N_3535,N_3335,N_3221);
xor U3536 (N_3536,N_3330,N_3294);
nor U3537 (N_3537,N_3205,N_3277);
nor U3538 (N_3538,N_3357,N_3319);
xnor U3539 (N_3539,N_3217,N_3358);
nand U3540 (N_3540,N_3279,N_3301);
or U3541 (N_3541,N_3294,N_3263);
xor U3542 (N_3542,N_3238,N_3281);
xnor U3543 (N_3543,N_3276,N_3269);
nor U3544 (N_3544,N_3292,N_3226);
nor U3545 (N_3545,N_3306,N_3337);
nor U3546 (N_3546,N_3304,N_3370);
or U3547 (N_3547,N_3250,N_3288);
and U3548 (N_3548,N_3300,N_3235);
or U3549 (N_3549,N_3231,N_3380);
nand U3550 (N_3550,N_3264,N_3229);
xnor U3551 (N_3551,N_3312,N_3396);
nor U3552 (N_3552,N_3366,N_3349);
nand U3553 (N_3553,N_3348,N_3266);
nand U3554 (N_3554,N_3270,N_3261);
or U3555 (N_3555,N_3381,N_3286);
xnor U3556 (N_3556,N_3300,N_3201);
nor U3557 (N_3557,N_3391,N_3330);
xnor U3558 (N_3558,N_3384,N_3230);
nor U3559 (N_3559,N_3314,N_3224);
or U3560 (N_3560,N_3307,N_3202);
nor U3561 (N_3561,N_3271,N_3294);
and U3562 (N_3562,N_3200,N_3296);
and U3563 (N_3563,N_3282,N_3384);
xnor U3564 (N_3564,N_3351,N_3342);
or U3565 (N_3565,N_3334,N_3383);
or U3566 (N_3566,N_3205,N_3299);
and U3567 (N_3567,N_3227,N_3331);
and U3568 (N_3568,N_3300,N_3341);
nand U3569 (N_3569,N_3365,N_3302);
or U3570 (N_3570,N_3381,N_3391);
nand U3571 (N_3571,N_3388,N_3205);
or U3572 (N_3572,N_3301,N_3359);
nor U3573 (N_3573,N_3280,N_3349);
nor U3574 (N_3574,N_3390,N_3238);
and U3575 (N_3575,N_3239,N_3248);
nor U3576 (N_3576,N_3376,N_3349);
nand U3577 (N_3577,N_3253,N_3346);
or U3578 (N_3578,N_3310,N_3208);
nand U3579 (N_3579,N_3325,N_3217);
nand U3580 (N_3580,N_3202,N_3363);
or U3581 (N_3581,N_3299,N_3248);
and U3582 (N_3582,N_3396,N_3314);
xnor U3583 (N_3583,N_3306,N_3263);
and U3584 (N_3584,N_3280,N_3381);
nor U3585 (N_3585,N_3252,N_3272);
or U3586 (N_3586,N_3304,N_3228);
nand U3587 (N_3587,N_3367,N_3378);
and U3588 (N_3588,N_3318,N_3211);
nand U3589 (N_3589,N_3289,N_3389);
and U3590 (N_3590,N_3254,N_3249);
nand U3591 (N_3591,N_3356,N_3252);
nand U3592 (N_3592,N_3213,N_3360);
or U3593 (N_3593,N_3336,N_3326);
xnor U3594 (N_3594,N_3299,N_3385);
nand U3595 (N_3595,N_3302,N_3374);
xor U3596 (N_3596,N_3265,N_3347);
nor U3597 (N_3597,N_3247,N_3244);
nand U3598 (N_3598,N_3258,N_3254);
and U3599 (N_3599,N_3387,N_3234);
nor U3600 (N_3600,N_3565,N_3592);
nand U3601 (N_3601,N_3562,N_3473);
nand U3602 (N_3602,N_3429,N_3522);
and U3603 (N_3603,N_3428,N_3501);
and U3604 (N_3604,N_3558,N_3515);
nand U3605 (N_3605,N_3402,N_3590);
nor U3606 (N_3606,N_3561,N_3455);
and U3607 (N_3607,N_3494,N_3410);
or U3608 (N_3608,N_3456,N_3571);
xnor U3609 (N_3609,N_3405,N_3553);
and U3610 (N_3610,N_3474,N_3491);
nand U3611 (N_3611,N_3564,N_3446);
nand U3612 (N_3612,N_3550,N_3544);
nor U3613 (N_3613,N_3478,N_3548);
xor U3614 (N_3614,N_3425,N_3596);
nand U3615 (N_3615,N_3483,N_3424);
xnor U3616 (N_3616,N_3467,N_3471);
or U3617 (N_3617,N_3400,N_3507);
nand U3618 (N_3618,N_3530,N_3479);
nand U3619 (N_3619,N_3529,N_3447);
or U3620 (N_3620,N_3487,N_3566);
and U3621 (N_3621,N_3427,N_3452);
nor U3622 (N_3622,N_3518,N_3576);
or U3623 (N_3623,N_3586,N_3537);
xnor U3624 (N_3624,N_3431,N_3449);
nor U3625 (N_3625,N_3542,N_3598);
and U3626 (N_3626,N_3572,N_3560);
or U3627 (N_3627,N_3461,N_3458);
or U3628 (N_3628,N_3477,N_3540);
and U3629 (N_3629,N_3510,N_3401);
or U3630 (N_3630,N_3497,N_3573);
nand U3631 (N_3631,N_3519,N_3503);
xnor U3632 (N_3632,N_3442,N_3414);
xnor U3633 (N_3633,N_3523,N_3493);
and U3634 (N_3634,N_3559,N_3408);
xnor U3635 (N_3635,N_3577,N_3450);
or U3636 (N_3636,N_3593,N_3480);
xnor U3637 (N_3637,N_3570,N_3517);
nand U3638 (N_3638,N_3539,N_3505);
nand U3639 (N_3639,N_3422,N_3500);
or U3640 (N_3640,N_3413,N_3437);
nand U3641 (N_3641,N_3541,N_3441);
nand U3642 (N_3642,N_3489,N_3403);
nor U3643 (N_3643,N_3538,N_3569);
or U3644 (N_3644,N_3521,N_3459);
and U3645 (N_3645,N_3587,N_3472);
nand U3646 (N_3646,N_3495,N_3464);
or U3647 (N_3647,N_3526,N_3585);
and U3648 (N_3648,N_3496,N_3490);
and U3649 (N_3649,N_3486,N_3454);
xor U3650 (N_3650,N_3543,N_3504);
xnor U3651 (N_3651,N_3440,N_3545);
nand U3652 (N_3652,N_3568,N_3527);
nand U3653 (N_3653,N_3406,N_3438);
nand U3654 (N_3654,N_3439,N_3580);
or U3655 (N_3655,N_3514,N_3463);
nor U3656 (N_3656,N_3535,N_3445);
nor U3657 (N_3657,N_3426,N_3595);
xnor U3658 (N_3658,N_3546,N_3436);
or U3659 (N_3659,N_3525,N_3420);
nand U3660 (N_3660,N_3448,N_3488);
or U3661 (N_3661,N_3599,N_3407);
nand U3662 (N_3662,N_3502,N_3423);
or U3663 (N_3663,N_3453,N_3582);
nand U3664 (N_3664,N_3597,N_3584);
or U3665 (N_3665,N_3444,N_3591);
xnor U3666 (N_3666,N_3470,N_3520);
and U3667 (N_3667,N_3554,N_3511);
nand U3668 (N_3668,N_3579,N_3524);
or U3669 (N_3669,N_3475,N_3512);
or U3670 (N_3670,N_3555,N_3481);
xor U3671 (N_3671,N_3581,N_3536);
nand U3672 (N_3672,N_3430,N_3415);
xor U3673 (N_3673,N_3508,N_3551);
xnor U3674 (N_3674,N_3575,N_3465);
or U3675 (N_3675,N_3433,N_3443);
nand U3676 (N_3676,N_3589,N_3549);
nor U3677 (N_3677,N_3532,N_3516);
xnor U3678 (N_3678,N_3462,N_3556);
or U3679 (N_3679,N_3513,N_3492);
and U3680 (N_3680,N_3412,N_3509);
nand U3681 (N_3681,N_3419,N_3531);
nor U3682 (N_3682,N_3484,N_3534);
xor U3683 (N_3683,N_3421,N_3404);
and U3684 (N_3684,N_3482,N_3432);
xor U3685 (N_3685,N_3552,N_3466);
or U3686 (N_3686,N_3588,N_3476);
and U3687 (N_3687,N_3583,N_3469);
xnor U3688 (N_3688,N_3411,N_3435);
xor U3689 (N_3689,N_3563,N_3416);
nand U3690 (N_3690,N_3451,N_3528);
or U3691 (N_3691,N_3574,N_3409);
or U3692 (N_3692,N_3460,N_3594);
nand U3693 (N_3693,N_3557,N_3567);
nand U3694 (N_3694,N_3457,N_3498);
nor U3695 (N_3695,N_3485,N_3417);
xnor U3696 (N_3696,N_3499,N_3506);
nor U3697 (N_3697,N_3434,N_3468);
xnor U3698 (N_3698,N_3533,N_3578);
or U3699 (N_3699,N_3418,N_3547);
xor U3700 (N_3700,N_3481,N_3418);
nor U3701 (N_3701,N_3579,N_3598);
and U3702 (N_3702,N_3584,N_3550);
nor U3703 (N_3703,N_3542,N_3443);
nor U3704 (N_3704,N_3565,N_3401);
and U3705 (N_3705,N_3542,N_3470);
nor U3706 (N_3706,N_3421,N_3512);
nor U3707 (N_3707,N_3507,N_3495);
or U3708 (N_3708,N_3431,N_3517);
or U3709 (N_3709,N_3501,N_3448);
xnor U3710 (N_3710,N_3434,N_3566);
or U3711 (N_3711,N_3521,N_3499);
xor U3712 (N_3712,N_3455,N_3501);
nor U3713 (N_3713,N_3499,N_3466);
or U3714 (N_3714,N_3515,N_3492);
and U3715 (N_3715,N_3401,N_3574);
xor U3716 (N_3716,N_3445,N_3465);
and U3717 (N_3717,N_3570,N_3425);
or U3718 (N_3718,N_3469,N_3437);
or U3719 (N_3719,N_3578,N_3568);
nand U3720 (N_3720,N_3465,N_3485);
xnor U3721 (N_3721,N_3569,N_3492);
xnor U3722 (N_3722,N_3448,N_3596);
nor U3723 (N_3723,N_3554,N_3474);
xnor U3724 (N_3724,N_3554,N_3570);
nor U3725 (N_3725,N_3473,N_3456);
or U3726 (N_3726,N_3582,N_3581);
nor U3727 (N_3727,N_3475,N_3593);
xnor U3728 (N_3728,N_3563,N_3555);
nor U3729 (N_3729,N_3441,N_3514);
xnor U3730 (N_3730,N_3492,N_3460);
nor U3731 (N_3731,N_3466,N_3521);
or U3732 (N_3732,N_3512,N_3515);
or U3733 (N_3733,N_3454,N_3423);
and U3734 (N_3734,N_3564,N_3595);
or U3735 (N_3735,N_3501,N_3582);
nor U3736 (N_3736,N_3408,N_3458);
nand U3737 (N_3737,N_3419,N_3568);
and U3738 (N_3738,N_3478,N_3410);
xnor U3739 (N_3739,N_3564,N_3493);
xor U3740 (N_3740,N_3492,N_3468);
or U3741 (N_3741,N_3577,N_3467);
nand U3742 (N_3742,N_3497,N_3554);
nand U3743 (N_3743,N_3507,N_3560);
or U3744 (N_3744,N_3532,N_3512);
xnor U3745 (N_3745,N_3404,N_3456);
nand U3746 (N_3746,N_3484,N_3499);
nand U3747 (N_3747,N_3547,N_3598);
nand U3748 (N_3748,N_3595,N_3521);
or U3749 (N_3749,N_3420,N_3540);
nor U3750 (N_3750,N_3553,N_3512);
nor U3751 (N_3751,N_3417,N_3504);
nand U3752 (N_3752,N_3405,N_3511);
nand U3753 (N_3753,N_3402,N_3538);
or U3754 (N_3754,N_3542,N_3582);
nand U3755 (N_3755,N_3432,N_3592);
xnor U3756 (N_3756,N_3435,N_3416);
xor U3757 (N_3757,N_3481,N_3491);
xor U3758 (N_3758,N_3449,N_3434);
and U3759 (N_3759,N_3564,N_3508);
xnor U3760 (N_3760,N_3475,N_3518);
nand U3761 (N_3761,N_3596,N_3548);
and U3762 (N_3762,N_3526,N_3472);
nor U3763 (N_3763,N_3540,N_3577);
nor U3764 (N_3764,N_3487,N_3554);
nand U3765 (N_3765,N_3449,N_3550);
or U3766 (N_3766,N_3495,N_3584);
and U3767 (N_3767,N_3527,N_3480);
and U3768 (N_3768,N_3479,N_3431);
nand U3769 (N_3769,N_3437,N_3536);
nor U3770 (N_3770,N_3440,N_3543);
or U3771 (N_3771,N_3533,N_3559);
or U3772 (N_3772,N_3525,N_3566);
nand U3773 (N_3773,N_3566,N_3519);
nor U3774 (N_3774,N_3566,N_3561);
xor U3775 (N_3775,N_3485,N_3521);
xor U3776 (N_3776,N_3456,N_3421);
xnor U3777 (N_3777,N_3547,N_3529);
xnor U3778 (N_3778,N_3561,N_3463);
or U3779 (N_3779,N_3514,N_3547);
nor U3780 (N_3780,N_3421,N_3531);
nor U3781 (N_3781,N_3451,N_3588);
or U3782 (N_3782,N_3535,N_3598);
nor U3783 (N_3783,N_3406,N_3562);
nor U3784 (N_3784,N_3520,N_3557);
or U3785 (N_3785,N_3483,N_3489);
xor U3786 (N_3786,N_3506,N_3493);
and U3787 (N_3787,N_3486,N_3565);
nor U3788 (N_3788,N_3569,N_3587);
nand U3789 (N_3789,N_3405,N_3587);
or U3790 (N_3790,N_3504,N_3581);
and U3791 (N_3791,N_3406,N_3470);
or U3792 (N_3792,N_3411,N_3545);
nor U3793 (N_3793,N_3471,N_3579);
nand U3794 (N_3794,N_3408,N_3498);
and U3795 (N_3795,N_3465,N_3483);
xor U3796 (N_3796,N_3540,N_3481);
or U3797 (N_3797,N_3428,N_3486);
nand U3798 (N_3798,N_3480,N_3447);
nand U3799 (N_3799,N_3542,N_3424);
xor U3800 (N_3800,N_3781,N_3722);
xnor U3801 (N_3801,N_3660,N_3784);
xnor U3802 (N_3802,N_3793,N_3750);
and U3803 (N_3803,N_3763,N_3630);
nand U3804 (N_3804,N_3633,N_3651);
xor U3805 (N_3805,N_3770,N_3762);
or U3806 (N_3806,N_3674,N_3614);
nor U3807 (N_3807,N_3625,N_3647);
or U3808 (N_3808,N_3775,N_3726);
nand U3809 (N_3809,N_3759,N_3656);
and U3810 (N_3810,N_3623,N_3659);
nand U3811 (N_3811,N_3635,N_3745);
and U3812 (N_3812,N_3682,N_3730);
or U3813 (N_3813,N_3760,N_3697);
and U3814 (N_3814,N_3714,N_3669);
nand U3815 (N_3815,N_3733,N_3602);
nor U3816 (N_3816,N_3610,N_3641);
nor U3817 (N_3817,N_3799,N_3753);
and U3818 (N_3818,N_3694,N_3672);
xnor U3819 (N_3819,N_3658,N_3600);
nand U3820 (N_3820,N_3665,N_3734);
or U3821 (N_3821,N_3639,N_3649);
and U3822 (N_3822,N_3757,N_3776);
and U3823 (N_3823,N_3678,N_3691);
xnor U3824 (N_3824,N_3792,N_3783);
nor U3825 (N_3825,N_3667,N_3611);
xor U3826 (N_3826,N_3702,N_3715);
and U3827 (N_3827,N_3679,N_3687);
and U3828 (N_3828,N_3657,N_3628);
xor U3829 (N_3829,N_3735,N_3673);
xnor U3830 (N_3830,N_3650,N_3771);
nor U3831 (N_3831,N_3743,N_3744);
xor U3832 (N_3832,N_3703,N_3706);
xnor U3833 (N_3833,N_3725,N_3704);
nand U3834 (N_3834,N_3742,N_3688);
nor U3835 (N_3835,N_3731,N_3746);
xor U3836 (N_3836,N_3609,N_3620);
nand U3837 (N_3837,N_3663,N_3677);
xor U3838 (N_3838,N_3675,N_3720);
nand U3839 (N_3839,N_3699,N_3624);
nand U3840 (N_3840,N_3758,N_3648);
xnor U3841 (N_3841,N_3780,N_3616);
and U3842 (N_3842,N_3728,N_3740);
xnor U3843 (N_3843,N_3779,N_3652);
nand U3844 (N_3844,N_3747,N_3621);
nor U3845 (N_3845,N_3617,N_3676);
xnor U3846 (N_3846,N_3654,N_3768);
xor U3847 (N_3847,N_3769,N_3797);
nand U3848 (N_3848,N_3708,N_3701);
or U3849 (N_3849,N_3786,N_3619);
nand U3850 (N_3850,N_3721,N_3741);
nand U3851 (N_3851,N_3668,N_3790);
nor U3852 (N_3852,N_3789,N_3662);
nor U3853 (N_3853,N_3642,N_3637);
xnor U3854 (N_3854,N_3643,N_3751);
or U3855 (N_3855,N_3622,N_3670);
nor U3856 (N_3856,N_3752,N_3729);
and U3857 (N_3857,N_3613,N_3795);
and U3858 (N_3858,N_3773,N_3724);
or U3859 (N_3859,N_3680,N_3796);
nand U3860 (N_3860,N_3655,N_3664);
nand U3861 (N_3861,N_3705,N_3767);
and U3862 (N_3862,N_3601,N_3774);
and U3863 (N_3863,N_3787,N_3713);
and U3864 (N_3864,N_3718,N_3707);
and U3865 (N_3865,N_3606,N_3719);
nand U3866 (N_3866,N_3712,N_3618);
or U3867 (N_3867,N_3666,N_3794);
nor U3868 (N_3868,N_3754,N_3723);
nor U3869 (N_3869,N_3645,N_3661);
nand U3870 (N_3870,N_3627,N_3671);
and U3871 (N_3871,N_3717,N_3629);
nor U3872 (N_3872,N_3693,N_3709);
nand U3873 (N_3873,N_3727,N_3695);
nor U3874 (N_3874,N_3698,N_3765);
and U3875 (N_3875,N_3612,N_3604);
nor U3876 (N_3876,N_3646,N_3764);
or U3877 (N_3877,N_3653,N_3638);
nor U3878 (N_3878,N_3685,N_3605);
nor U3879 (N_3879,N_3710,N_3772);
xor U3880 (N_3880,N_3748,N_3607);
and U3881 (N_3881,N_3615,N_3700);
or U3882 (N_3882,N_3778,N_3798);
and U3883 (N_3883,N_3785,N_3737);
xnor U3884 (N_3884,N_3777,N_3690);
xor U3885 (N_3885,N_3683,N_3644);
or U3886 (N_3886,N_3634,N_3782);
or U3887 (N_3887,N_3732,N_3692);
and U3888 (N_3888,N_3603,N_3761);
or U3889 (N_3889,N_3788,N_3684);
nand U3890 (N_3890,N_3626,N_3738);
or U3891 (N_3891,N_3640,N_3736);
or U3892 (N_3892,N_3755,N_3716);
xnor U3893 (N_3893,N_3632,N_3608);
nand U3894 (N_3894,N_3756,N_3681);
or U3895 (N_3895,N_3791,N_3696);
nor U3896 (N_3896,N_3689,N_3711);
xnor U3897 (N_3897,N_3739,N_3766);
and U3898 (N_3898,N_3631,N_3636);
and U3899 (N_3899,N_3749,N_3686);
nor U3900 (N_3900,N_3756,N_3662);
xor U3901 (N_3901,N_3746,N_3773);
nand U3902 (N_3902,N_3713,N_3769);
and U3903 (N_3903,N_3771,N_3730);
nand U3904 (N_3904,N_3603,N_3775);
nor U3905 (N_3905,N_3738,N_3767);
or U3906 (N_3906,N_3706,N_3629);
or U3907 (N_3907,N_3632,N_3630);
nand U3908 (N_3908,N_3699,N_3753);
and U3909 (N_3909,N_3646,N_3795);
and U3910 (N_3910,N_3693,N_3696);
and U3911 (N_3911,N_3607,N_3695);
nand U3912 (N_3912,N_3603,N_3680);
xnor U3913 (N_3913,N_3762,N_3700);
nor U3914 (N_3914,N_3647,N_3792);
nand U3915 (N_3915,N_3682,N_3649);
nor U3916 (N_3916,N_3719,N_3660);
xor U3917 (N_3917,N_3649,N_3799);
and U3918 (N_3918,N_3670,N_3746);
nand U3919 (N_3919,N_3750,N_3673);
xnor U3920 (N_3920,N_3742,N_3604);
and U3921 (N_3921,N_3651,N_3744);
nand U3922 (N_3922,N_3653,N_3753);
nor U3923 (N_3923,N_3728,N_3681);
or U3924 (N_3924,N_3764,N_3758);
nor U3925 (N_3925,N_3610,N_3701);
nand U3926 (N_3926,N_3707,N_3783);
or U3927 (N_3927,N_3763,N_3710);
nand U3928 (N_3928,N_3644,N_3741);
or U3929 (N_3929,N_3672,N_3714);
nand U3930 (N_3930,N_3636,N_3707);
and U3931 (N_3931,N_3740,N_3643);
nor U3932 (N_3932,N_3656,N_3756);
nor U3933 (N_3933,N_3784,N_3708);
or U3934 (N_3934,N_3732,N_3799);
or U3935 (N_3935,N_3720,N_3639);
nand U3936 (N_3936,N_3710,N_3750);
nor U3937 (N_3937,N_3768,N_3694);
nand U3938 (N_3938,N_3747,N_3607);
or U3939 (N_3939,N_3723,N_3643);
or U3940 (N_3940,N_3727,N_3652);
or U3941 (N_3941,N_3760,N_3668);
nor U3942 (N_3942,N_3610,N_3627);
nand U3943 (N_3943,N_3665,N_3776);
and U3944 (N_3944,N_3620,N_3761);
xnor U3945 (N_3945,N_3782,N_3638);
and U3946 (N_3946,N_3626,N_3741);
nand U3947 (N_3947,N_3748,N_3600);
and U3948 (N_3948,N_3703,N_3794);
nor U3949 (N_3949,N_3685,N_3676);
and U3950 (N_3950,N_3745,N_3647);
nand U3951 (N_3951,N_3715,N_3774);
or U3952 (N_3952,N_3653,N_3603);
nor U3953 (N_3953,N_3607,N_3742);
or U3954 (N_3954,N_3606,N_3649);
or U3955 (N_3955,N_3738,N_3675);
xnor U3956 (N_3956,N_3632,N_3600);
nor U3957 (N_3957,N_3740,N_3724);
xor U3958 (N_3958,N_3740,N_3721);
xor U3959 (N_3959,N_3678,N_3748);
or U3960 (N_3960,N_3620,N_3760);
xor U3961 (N_3961,N_3675,N_3789);
and U3962 (N_3962,N_3702,N_3638);
xnor U3963 (N_3963,N_3692,N_3673);
or U3964 (N_3964,N_3626,N_3632);
nand U3965 (N_3965,N_3798,N_3746);
nand U3966 (N_3966,N_3701,N_3622);
nor U3967 (N_3967,N_3657,N_3770);
nor U3968 (N_3968,N_3694,N_3745);
and U3969 (N_3969,N_3614,N_3677);
nand U3970 (N_3970,N_3737,N_3623);
nor U3971 (N_3971,N_3611,N_3664);
nor U3972 (N_3972,N_3767,N_3788);
or U3973 (N_3973,N_3759,N_3640);
nor U3974 (N_3974,N_3722,N_3690);
nor U3975 (N_3975,N_3603,N_3694);
nand U3976 (N_3976,N_3744,N_3787);
nor U3977 (N_3977,N_3634,N_3772);
and U3978 (N_3978,N_3613,N_3745);
nor U3979 (N_3979,N_3781,N_3704);
xnor U3980 (N_3980,N_3687,N_3683);
xor U3981 (N_3981,N_3703,N_3605);
or U3982 (N_3982,N_3670,N_3749);
xor U3983 (N_3983,N_3706,N_3699);
and U3984 (N_3984,N_3646,N_3687);
or U3985 (N_3985,N_3741,N_3697);
or U3986 (N_3986,N_3741,N_3685);
xor U3987 (N_3987,N_3695,N_3674);
or U3988 (N_3988,N_3758,N_3716);
nand U3989 (N_3989,N_3781,N_3612);
nor U3990 (N_3990,N_3736,N_3781);
nor U3991 (N_3991,N_3660,N_3721);
nor U3992 (N_3992,N_3683,N_3614);
nor U3993 (N_3993,N_3607,N_3661);
nand U3994 (N_3994,N_3604,N_3721);
xnor U3995 (N_3995,N_3699,N_3752);
or U3996 (N_3996,N_3610,N_3611);
xnor U3997 (N_3997,N_3718,N_3611);
nor U3998 (N_3998,N_3792,N_3643);
nor U3999 (N_3999,N_3670,N_3743);
nand U4000 (N_4000,N_3879,N_3893);
or U4001 (N_4001,N_3861,N_3881);
xnor U4002 (N_4002,N_3832,N_3876);
xnor U4003 (N_4003,N_3947,N_3846);
nor U4004 (N_4004,N_3965,N_3921);
nand U4005 (N_4005,N_3908,N_3910);
xor U4006 (N_4006,N_3951,N_3826);
or U4007 (N_4007,N_3953,N_3806);
xor U4008 (N_4008,N_3877,N_3828);
nand U4009 (N_4009,N_3923,N_3903);
nand U4010 (N_4010,N_3928,N_3853);
nor U4011 (N_4011,N_3834,N_3837);
and U4012 (N_4012,N_3956,N_3823);
nor U4013 (N_4013,N_3969,N_3899);
or U4014 (N_4014,N_3912,N_3831);
and U4015 (N_4015,N_3925,N_3977);
nor U4016 (N_4016,N_3922,N_3855);
and U4017 (N_4017,N_3993,N_3946);
nor U4018 (N_4018,N_3935,N_3984);
nor U4019 (N_4019,N_3962,N_3864);
or U4020 (N_4020,N_3974,N_3992);
and U4021 (N_4021,N_3822,N_3900);
or U4022 (N_4022,N_3952,N_3988);
nor U4023 (N_4023,N_3802,N_3865);
nor U4024 (N_4024,N_3889,N_3886);
nand U4025 (N_4025,N_3820,N_3982);
nor U4026 (N_4026,N_3936,N_3816);
or U4027 (N_4027,N_3960,N_3856);
and U4028 (N_4028,N_3873,N_3959);
nor U4029 (N_4029,N_3887,N_3800);
nand U4030 (N_4030,N_3811,N_3862);
nand U4031 (N_4031,N_3814,N_3851);
or U4032 (N_4032,N_3915,N_3906);
xnor U4033 (N_4033,N_3919,N_3808);
and U4034 (N_4034,N_3938,N_3932);
xnor U4035 (N_4035,N_3849,N_3911);
xor U4036 (N_4036,N_3905,N_3878);
and U4037 (N_4037,N_3942,N_3884);
nand U4038 (N_4038,N_3848,N_3805);
nor U4039 (N_4039,N_3869,N_3989);
nor U4040 (N_4040,N_3863,N_3883);
nor U4041 (N_4041,N_3941,N_3896);
and U4042 (N_4042,N_3839,N_3833);
nor U4043 (N_4043,N_3998,N_3940);
nand U4044 (N_4044,N_3968,N_3819);
or U4045 (N_4045,N_3929,N_3894);
nand U4046 (N_4046,N_3954,N_3990);
xnor U4047 (N_4047,N_3987,N_3892);
xor U4048 (N_4048,N_3857,N_3842);
and U4049 (N_4049,N_3850,N_3815);
nor U4050 (N_4050,N_3909,N_3882);
or U4051 (N_4051,N_3872,N_3888);
or U4052 (N_4052,N_3971,N_3890);
nand U4053 (N_4053,N_3926,N_3854);
and U4054 (N_4054,N_3920,N_3994);
nand U4055 (N_4055,N_3966,N_3867);
nand U4056 (N_4056,N_3976,N_3841);
or U4057 (N_4057,N_3972,N_3866);
nor U4058 (N_4058,N_3817,N_3949);
xnor U4059 (N_4059,N_3948,N_3875);
or U4060 (N_4060,N_3933,N_3897);
xnor U4061 (N_4061,N_3830,N_3858);
nor U4062 (N_4062,N_3803,N_3983);
or U4063 (N_4063,N_3980,N_3918);
xnor U4064 (N_4064,N_3825,N_3985);
and U4065 (N_4065,N_3964,N_3874);
nand U4066 (N_4066,N_3902,N_3810);
or U4067 (N_4067,N_3978,N_3845);
nor U4068 (N_4068,N_3995,N_3907);
nor U4069 (N_4069,N_3945,N_3930);
nand U4070 (N_4070,N_3914,N_3818);
nand U4071 (N_4071,N_3838,N_3973);
or U4072 (N_4072,N_3904,N_3813);
or U4073 (N_4073,N_3852,N_3880);
nor U4074 (N_4074,N_3870,N_3916);
xor U4075 (N_4075,N_3807,N_3961);
xor U4076 (N_4076,N_3809,N_3847);
nor U4077 (N_4077,N_3859,N_3979);
and U4078 (N_4078,N_3937,N_3997);
nand U4079 (N_4079,N_3901,N_3844);
nor U4080 (N_4080,N_3967,N_3996);
nand U4081 (N_4081,N_3991,N_3931);
or U4082 (N_4082,N_3934,N_3958);
nor U4083 (N_4083,N_3975,N_3927);
nor U4084 (N_4084,N_3913,N_3944);
xor U4085 (N_4085,N_3999,N_3970);
xnor U4086 (N_4086,N_3824,N_3836);
xor U4087 (N_4087,N_3981,N_3950);
nor U4088 (N_4088,N_3804,N_3868);
and U4089 (N_4089,N_3955,N_3943);
nor U4090 (N_4090,N_3895,N_3871);
xor U4091 (N_4091,N_3963,N_3801);
or U4092 (N_4092,N_3986,N_3812);
and U4093 (N_4093,N_3885,N_3957);
nor U4094 (N_4094,N_3843,N_3898);
nor U4095 (N_4095,N_3939,N_3860);
nor U4096 (N_4096,N_3917,N_3840);
nor U4097 (N_4097,N_3924,N_3829);
or U4098 (N_4098,N_3827,N_3835);
and U4099 (N_4099,N_3821,N_3891);
nor U4100 (N_4100,N_3986,N_3806);
nor U4101 (N_4101,N_3888,N_3816);
nand U4102 (N_4102,N_3919,N_3814);
and U4103 (N_4103,N_3891,N_3964);
or U4104 (N_4104,N_3867,N_3856);
nand U4105 (N_4105,N_3868,N_3856);
and U4106 (N_4106,N_3817,N_3961);
or U4107 (N_4107,N_3852,N_3962);
or U4108 (N_4108,N_3953,N_3965);
and U4109 (N_4109,N_3917,N_3957);
or U4110 (N_4110,N_3870,N_3969);
and U4111 (N_4111,N_3905,N_3827);
nand U4112 (N_4112,N_3920,N_3857);
nor U4113 (N_4113,N_3943,N_3851);
or U4114 (N_4114,N_3846,N_3819);
nor U4115 (N_4115,N_3984,N_3917);
nor U4116 (N_4116,N_3866,N_3854);
nand U4117 (N_4117,N_3909,N_3863);
or U4118 (N_4118,N_3906,N_3947);
and U4119 (N_4119,N_3894,N_3821);
nand U4120 (N_4120,N_3889,N_3893);
or U4121 (N_4121,N_3979,N_3877);
xnor U4122 (N_4122,N_3922,N_3970);
xnor U4123 (N_4123,N_3962,N_3976);
xnor U4124 (N_4124,N_3995,N_3905);
or U4125 (N_4125,N_3841,N_3928);
xor U4126 (N_4126,N_3902,N_3998);
and U4127 (N_4127,N_3977,N_3926);
xnor U4128 (N_4128,N_3911,N_3973);
nor U4129 (N_4129,N_3968,N_3892);
nand U4130 (N_4130,N_3924,N_3856);
or U4131 (N_4131,N_3944,N_3988);
nor U4132 (N_4132,N_3996,N_3814);
xnor U4133 (N_4133,N_3961,N_3906);
or U4134 (N_4134,N_3961,N_3971);
and U4135 (N_4135,N_3967,N_3878);
nor U4136 (N_4136,N_3873,N_3849);
xnor U4137 (N_4137,N_3842,N_3862);
and U4138 (N_4138,N_3953,N_3884);
nand U4139 (N_4139,N_3976,N_3821);
xor U4140 (N_4140,N_3927,N_3900);
or U4141 (N_4141,N_3843,N_3902);
and U4142 (N_4142,N_3959,N_3919);
nor U4143 (N_4143,N_3830,N_3842);
nand U4144 (N_4144,N_3807,N_3998);
xor U4145 (N_4145,N_3966,N_3846);
or U4146 (N_4146,N_3834,N_3983);
or U4147 (N_4147,N_3800,N_3930);
or U4148 (N_4148,N_3957,N_3812);
nor U4149 (N_4149,N_3817,N_3805);
xnor U4150 (N_4150,N_3822,N_3978);
xnor U4151 (N_4151,N_3973,N_3935);
xor U4152 (N_4152,N_3875,N_3904);
and U4153 (N_4153,N_3958,N_3917);
nor U4154 (N_4154,N_3816,N_3855);
or U4155 (N_4155,N_3966,N_3925);
or U4156 (N_4156,N_3889,N_3895);
and U4157 (N_4157,N_3993,N_3808);
or U4158 (N_4158,N_3863,N_3983);
nor U4159 (N_4159,N_3930,N_3810);
xor U4160 (N_4160,N_3938,N_3804);
nand U4161 (N_4161,N_3841,N_3966);
nand U4162 (N_4162,N_3886,N_3983);
nor U4163 (N_4163,N_3866,N_3992);
and U4164 (N_4164,N_3831,N_3845);
nand U4165 (N_4165,N_3880,N_3839);
and U4166 (N_4166,N_3925,N_3880);
nand U4167 (N_4167,N_3852,N_3989);
nand U4168 (N_4168,N_3831,N_3944);
or U4169 (N_4169,N_3939,N_3931);
xor U4170 (N_4170,N_3897,N_3914);
and U4171 (N_4171,N_3870,N_3945);
nand U4172 (N_4172,N_3893,N_3991);
nor U4173 (N_4173,N_3972,N_3835);
and U4174 (N_4174,N_3808,N_3903);
nor U4175 (N_4175,N_3834,N_3972);
and U4176 (N_4176,N_3943,N_3899);
and U4177 (N_4177,N_3995,N_3807);
nor U4178 (N_4178,N_3839,N_3843);
nor U4179 (N_4179,N_3876,N_3927);
nand U4180 (N_4180,N_3801,N_3961);
xnor U4181 (N_4181,N_3964,N_3968);
nand U4182 (N_4182,N_3927,N_3928);
and U4183 (N_4183,N_3973,N_3881);
nor U4184 (N_4184,N_3872,N_3921);
nand U4185 (N_4185,N_3886,N_3963);
nand U4186 (N_4186,N_3844,N_3914);
nor U4187 (N_4187,N_3900,N_3894);
nor U4188 (N_4188,N_3989,N_3926);
or U4189 (N_4189,N_3943,N_3966);
or U4190 (N_4190,N_3884,N_3893);
or U4191 (N_4191,N_3948,N_3967);
or U4192 (N_4192,N_3822,N_3842);
xor U4193 (N_4193,N_3993,N_3916);
nor U4194 (N_4194,N_3930,N_3964);
nand U4195 (N_4195,N_3806,N_3877);
and U4196 (N_4196,N_3843,N_3812);
nor U4197 (N_4197,N_3812,N_3807);
nand U4198 (N_4198,N_3820,N_3880);
nand U4199 (N_4199,N_3967,N_3889);
or U4200 (N_4200,N_4179,N_4171);
nand U4201 (N_4201,N_4122,N_4100);
nor U4202 (N_4202,N_4069,N_4178);
nor U4203 (N_4203,N_4097,N_4096);
and U4204 (N_4204,N_4057,N_4110);
xor U4205 (N_4205,N_4169,N_4128);
nand U4206 (N_4206,N_4166,N_4083);
nand U4207 (N_4207,N_4176,N_4133);
xnor U4208 (N_4208,N_4117,N_4153);
or U4209 (N_4209,N_4047,N_4199);
nor U4210 (N_4210,N_4186,N_4037);
and U4211 (N_4211,N_4028,N_4078);
nor U4212 (N_4212,N_4061,N_4104);
xor U4213 (N_4213,N_4050,N_4013);
xor U4214 (N_4214,N_4075,N_4024);
nor U4215 (N_4215,N_4058,N_4067);
or U4216 (N_4216,N_4021,N_4015);
nor U4217 (N_4217,N_4158,N_4160);
nor U4218 (N_4218,N_4172,N_4090);
and U4219 (N_4219,N_4027,N_4001);
xnor U4220 (N_4220,N_4018,N_4064);
or U4221 (N_4221,N_4109,N_4073);
or U4222 (N_4222,N_4066,N_4148);
nor U4223 (N_4223,N_4193,N_4146);
nand U4224 (N_4224,N_4164,N_4099);
or U4225 (N_4225,N_4080,N_4114);
xor U4226 (N_4226,N_4065,N_4145);
nor U4227 (N_4227,N_4118,N_4081);
and U4228 (N_4228,N_4119,N_4043);
xnor U4229 (N_4229,N_4184,N_4152);
or U4230 (N_4230,N_4046,N_4054);
and U4231 (N_4231,N_4044,N_4170);
and U4232 (N_4232,N_4007,N_4012);
xnor U4233 (N_4233,N_4130,N_4175);
xor U4234 (N_4234,N_4134,N_4019);
xor U4235 (N_4235,N_4053,N_4036);
xor U4236 (N_4236,N_4198,N_4063);
and U4237 (N_4237,N_4163,N_4173);
nor U4238 (N_4238,N_4004,N_4103);
nand U4239 (N_4239,N_4105,N_4113);
nor U4240 (N_4240,N_4041,N_4154);
or U4241 (N_4241,N_4086,N_4142);
nand U4242 (N_4242,N_4022,N_4143);
nor U4243 (N_4243,N_4031,N_4033);
nor U4244 (N_4244,N_4094,N_4045);
xor U4245 (N_4245,N_4156,N_4077);
nand U4246 (N_4246,N_4111,N_4161);
or U4247 (N_4247,N_4183,N_4196);
nand U4248 (N_4248,N_4026,N_4121);
and U4249 (N_4249,N_4032,N_4010);
nand U4250 (N_4250,N_4115,N_4151);
nand U4251 (N_4251,N_4011,N_4023);
nor U4252 (N_4252,N_4020,N_4074);
nor U4253 (N_4253,N_4182,N_4005);
nand U4254 (N_4254,N_4095,N_4009);
nor U4255 (N_4255,N_4055,N_4008);
nand U4256 (N_4256,N_4189,N_4006);
nor U4257 (N_4257,N_4092,N_4125);
nor U4258 (N_4258,N_4136,N_4167);
or U4259 (N_4259,N_4137,N_4079);
xor U4260 (N_4260,N_4060,N_4070);
and U4261 (N_4261,N_4002,N_4029);
and U4262 (N_4262,N_4174,N_4087);
nand U4263 (N_4263,N_4159,N_4000);
or U4264 (N_4264,N_4042,N_4139);
nand U4265 (N_4265,N_4091,N_4112);
nor U4266 (N_4266,N_4195,N_4030);
or U4267 (N_4267,N_4181,N_4150);
nor U4268 (N_4268,N_4120,N_4016);
xnor U4269 (N_4269,N_4088,N_4072);
nand U4270 (N_4270,N_4056,N_4165);
xor U4271 (N_4271,N_4188,N_4116);
nor U4272 (N_4272,N_4048,N_4082);
or U4273 (N_4273,N_4049,N_4177);
nand U4274 (N_4274,N_4093,N_4068);
nor U4275 (N_4275,N_4123,N_4089);
and U4276 (N_4276,N_4190,N_4102);
nor U4277 (N_4277,N_4085,N_4062);
nand U4278 (N_4278,N_4180,N_4168);
or U4279 (N_4279,N_4144,N_4084);
and U4280 (N_4280,N_4108,N_4197);
or U4281 (N_4281,N_4149,N_4135);
nor U4282 (N_4282,N_4124,N_4194);
nor U4283 (N_4283,N_4106,N_4147);
nand U4284 (N_4284,N_4138,N_4185);
nand U4285 (N_4285,N_4162,N_4039);
xnor U4286 (N_4286,N_4025,N_4003);
or U4287 (N_4287,N_4187,N_4017);
nand U4288 (N_4288,N_4059,N_4129);
nor U4289 (N_4289,N_4192,N_4157);
and U4290 (N_4290,N_4127,N_4071);
or U4291 (N_4291,N_4155,N_4051);
xor U4292 (N_4292,N_4140,N_4101);
and U4293 (N_4293,N_4107,N_4191);
nand U4294 (N_4294,N_4038,N_4035);
nand U4295 (N_4295,N_4141,N_4052);
or U4296 (N_4296,N_4076,N_4131);
xnor U4297 (N_4297,N_4014,N_4126);
nor U4298 (N_4298,N_4040,N_4034);
nand U4299 (N_4299,N_4132,N_4098);
xor U4300 (N_4300,N_4124,N_4183);
nor U4301 (N_4301,N_4108,N_4133);
and U4302 (N_4302,N_4136,N_4033);
xnor U4303 (N_4303,N_4009,N_4043);
nor U4304 (N_4304,N_4121,N_4119);
xnor U4305 (N_4305,N_4039,N_4168);
or U4306 (N_4306,N_4136,N_4150);
nand U4307 (N_4307,N_4037,N_4065);
nand U4308 (N_4308,N_4094,N_4196);
nand U4309 (N_4309,N_4065,N_4053);
nor U4310 (N_4310,N_4047,N_4190);
or U4311 (N_4311,N_4160,N_4105);
nand U4312 (N_4312,N_4051,N_4104);
and U4313 (N_4313,N_4027,N_4004);
nor U4314 (N_4314,N_4175,N_4194);
xor U4315 (N_4315,N_4084,N_4073);
nor U4316 (N_4316,N_4172,N_4142);
xnor U4317 (N_4317,N_4102,N_4048);
or U4318 (N_4318,N_4046,N_4063);
xor U4319 (N_4319,N_4107,N_4077);
xnor U4320 (N_4320,N_4003,N_4073);
nor U4321 (N_4321,N_4006,N_4073);
xor U4322 (N_4322,N_4151,N_4090);
and U4323 (N_4323,N_4089,N_4033);
and U4324 (N_4324,N_4000,N_4104);
nor U4325 (N_4325,N_4136,N_4170);
nand U4326 (N_4326,N_4065,N_4022);
nand U4327 (N_4327,N_4042,N_4149);
nand U4328 (N_4328,N_4145,N_4169);
nor U4329 (N_4329,N_4085,N_4067);
nand U4330 (N_4330,N_4044,N_4034);
and U4331 (N_4331,N_4193,N_4042);
nor U4332 (N_4332,N_4077,N_4060);
nand U4333 (N_4333,N_4190,N_4121);
xor U4334 (N_4334,N_4089,N_4087);
xor U4335 (N_4335,N_4060,N_4115);
nor U4336 (N_4336,N_4068,N_4145);
nand U4337 (N_4337,N_4035,N_4147);
nand U4338 (N_4338,N_4002,N_4007);
and U4339 (N_4339,N_4056,N_4034);
and U4340 (N_4340,N_4107,N_4146);
nand U4341 (N_4341,N_4171,N_4104);
nor U4342 (N_4342,N_4123,N_4133);
and U4343 (N_4343,N_4139,N_4180);
and U4344 (N_4344,N_4117,N_4142);
xnor U4345 (N_4345,N_4079,N_4135);
and U4346 (N_4346,N_4123,N_4042);
or U4347 (N_4347,N_4145,N_4127);
or U4348 (N_4348,N_4132,N_4031);
nor U4349 (N_4349,N_4194,N_4145);
and U4350 (N_4350,N_4027,N_4174);
nor U4351 (N_4351,N_4158,N_4049);
xnor U4352 (N_4352,N_4186,N_4026);
nor U4353 (N_4353,N_4191,N_4186);
nor U4354 (N_4354,N_4076,N_4198);
xnor U4355 (N_4355,N_4073,N_4037);
or U4356 (N_4356,N_4086,N_4186);
xnor U4357 (N_4357,N_4048,N_4045);
and U4358 (N_4358,N_4068,N_4185);
nand U4359 (N_4359,N_4162,N_4101);
nand U4360 (N_4360,N_4017,N_4066);
and U4361 (N_4361,N_4133,N_4157);
nand U4362 (N_4362,N_4088,N_4060);
and U4363 (N_4363,N_4054,N_4072);
xor U4364 (N_4364,N_4009,N_4077);
and U4365 (N_4365,N_4000,N_4152);
xor U4366 (N_4366,N_4109,N_4065);
or U4367 (N_4367,N_4019,N_4012);
xor U4368 (N_4368,N_4094,N_4125);
xnor U4369 (N_4369,N_4053,N_4035);
xor U4370 (N_4370,N_4127,N_4030);
or U4371 (N_4371,N_4175,N_4044);
nand U4372 (N_4372,N_4131,N_4174);
nand U4373 (N_4373,N_4179,N_4060);
xnor U4374 (N_4374,N_4157,N_4014);
nor U4375 (N_4375,N_4072,N_4160);
and U4376 (N_4376,N_4009,N_4011);
and U4377 (N_4377,N_4086,N_4113);
xnor U4378 (N_4378,N_4010,N_4113);
nand U4379 (N_4379,N_4198,N_4169);
or U4380 (N_4380,N_4113,N_4121);
xnor U4381 (N_4381,N_4186,N_4193);
and U4382 (N_4382,N_4075,N_4068);
or U4383 (N_4383,N_4003,N_4110);
nor U4384 (N_4384,N_4105,N_4198);
nor U4385 (N_4385,N_4197,N_4123);
nor U4386 (N_4386,N_4064,N_4066);
nor U4387 (N_4387,N_4098,N_4153);
nor U4388 (N_4388,N_4157,N_4097);
or U4389 (N_4389,N_4082,N_4174);
and U4390 (N_4390,N_4165,N_4143);
and U4391 (N_4391,N_4087,N_4159);
and U4392 (N_4392,N_4129,N_4019);
nand U4393 (N_4393,N_4189,N_4181);
nand U4394 (N_4394,N_4006,N_4151);
xnor U4395 (N_4395,N_4016,N_4057);
or U4396 (N_4396,N_4014,N_4091);
or U4397 (N_4397,N_4153,N_4145);
xnor U4398 (N_4398,N_4043,N_4032);
or U4399 (N_4399,N_4158,N_4157);
nor U4400 (N_4400,N_4321,N_4286);
and U4401 (N_4401,N_4209,N_4295);
and U4402 (N_4402,N_4218,N_4399);
and U4403 (N_4403,N_4262,N_4253);
xnor U4404 (N_4404,N_4367,N_4364);
or U4405 (N_4405,N_4379,N_4393);
nand U4406 (N_4406,N_4330,N_4226);
and U4407 (N_4407,N_4248,N_4341);
or U4408 (N_4408,N_4357,N_4313);
or U4409 (N_4409,N_4351,N_4237);
or U4410 (N_4410,N_4229,N_4352);
and U4411 (N_4411,N_4365,N_4216);
nor U4412 (N_4412,N_4398,N_4245);
or U4413 (N_4413,N_4231,N_4207);
and U4414 (N_4414,N_4247,N_4288);
nor U4415 (N_4415,N_4228,N_4290);
and U4416 (N_4416,N_4240,N_4267);
nor U4417 (N_4417,N_4202,N_4257);
xnor U4418 (N_4418,N_4258,N_4328);
nand U4419 (N_4419,N_4268,N_4235);
nand U4420 (N_4420,N_4389,N_4319);
nor U4421 (N_4421,N_4305,N_4312);
nand U4422 (N_4422,N_4356,N_4390);
nand U4423 (N_4423,N_4287,N_4334);
nand U4424 (N_4424,N_4238,N_4347);
nand U4425 (N_4425,N_4252,N_4336);
xnor U4426 (N_4426,N_4266,N_4339);
nand U4427 (N_4427,N_4396,N_4368);
or U4428 (N_4428,N_4314,N_4333);
nand U4429 (N_4429,N_4210,N_4221);
xnor U4430 (N_4430,N_4222,N_4318);
xor U4431 (N_4431,N_4215,N_4373);
or U4432 (N_4432,N_4392,N_4224);
nand U4433 (N_4433,N_4255,N_4261);
nand U4434 (N_4434,N_4274,N_4244);
nor U4435 (N_4435,N_4350,N_4316);
xor U4436 (N_4436,N_4306,N_4243);
nand U4437 (N_4437,N_4284,N_4346);
and U4438 (N_4438,N_4292,N_4296);
xor U4439 (N_4439,N_4386,N_4359);
or U4440 (N_4440,N_4301,N_4310);
nor U4441 (N_4441,N_4325,N_4382);
or U4442 (N_4442,N_4242,N_4358);
nor U4443 (N_4443,N_4276,N_4323);
or U4444 (N_4444,N_4311,N_4353);
or U4445 (N_4445,N_4377,N_4269);
and U4446 (N_4446,N_4303,N_4384);
and U4447 (N_4447,N_4370,N_4395);
xor U4448 (N_4448,N_4340,N_4348);
or U4449 (N_4449,N_4217,N_4285);
xor U4450 (N_4450,N_4337,N_4214);
nor U4451 (N_4451,N_4291,N_4349);
nor U4452 (N_4452,N_4272,N_4263);
nor U4453 (N_4453,N_4345,N_4283);
or U4454 (N_4454,N_4363,N_4232);
xor U4455 (N_4455,N_4208,N_4338);
nand U4456 (N_4456,N_4374,N_4203);
and U4457 (N_4457,N_4293,N_4200);
nand U4458 (N_4458,N_4360,N_4309);
xnor U4459 (N_4459,N_4264,N_4236);
or U4460 (N_4460,N_4332,N_4320);
nand U4461 (N_4461,N_4304,N_4230);
or U4462 (N_4462,N_4302,N_4246);
and U4463 (N_4463,N_4277,N_4329);
nor U4464 (N_4464,N_4204,N_4241);
nor U4465 (N_4465,N_4315,N_4220);
xor U4466 (N_4466,N_4289,N_4233);
nor U4467 (N_4467,N_4326,N_4227);
and U4468 (N_4468,N_4254,N_4397);
or U4469 (N_4469,N_4223,N_4282);
nor U4470 (N_4470,N_4256,N_4383);
and U4471 (N_4471,N_4294,N_4378);
xnor U4472 (N_4472,N_4317,N_4376);
or U4473 (N_4473,N_4300,N_4343);
or U4474 (N_4474,N_4251,N_4213);
nor U4475 (N_4475,N_4371,N_4381);
xor U4476 (N_4476,N_4362,N_4273);
or U4477 (N_4477,N_4249,N_4327);
or U4478 (N_4478,N_4298,N_4354);
or U4479 (N_4479,N_4385,N_4394);
xor U4480 (N_4480,N_4307,N_4335);
and U4481 (N_4481,N_4372,N_4322);
or U4482 (N_4482,N_4342,N_4201);
nor U4483 (N_4483,N_4344,N_4380);
nand U4484 (N_4484,N_4279,N_4259);
and U4485 (N_4485,N_4388,N_4250);
nand U4486 (N_4486,N_4219,N_4239);
xor U4487 (N_4487,N_4205,N_4234);
xor U4488 (N_4488,N_4212,N_4225);
or U4489 (N_4489,N_4270,N_4278);
xor U4490 (N_4490,N_4308,N_4324);
nand U4491 (N_4491,N_4206,N_4391);
xnor U4492 (N_4492,N_4331,N_4297);
and U4493 (N_4493,N_4275,N_4375);
nor U4494 (N_4494,N_4366,N_4211);
or U4495 (N_4495,N_4260,N_4361);
nor U4496 (N_4496,N_4281,N_4369);
or U4497 (N_4497,N_4280,N_4271);
or U4498 (N_4498,N_4387,N_4265);
and U4499 (N_4499,N_4355,N_4299);
nor U4500 (N_4500,N_4342,N_4389);
and U4501 (N_4501,N_4370,N_4304);
nor U4502 (N_4502,N_4288,N_4266);
and U4503 (N_4503,N_4261,N_4279);
xor U4504 (N_4504,N_4361,N_4259);
xor U4505 (N_4505,N_4214,N_4293);
and U4506 (N_4506,N_4332,N_4301);
xor U4507 (N_4507,N_4300,N_4374);
and U4508 (N_4508,N_4300,N_4350);
nor U4509 (N_4509,N_4259,N_4395);
or U4510 (N_4510,N_4321,N_4303);
and U4511 (N_4511,N_4250,N_4308);
nor U4512 (N_4512,N_4233,N_4245);
xnor U4513 (N_4513,N_4239,N_4354);
xnor U4514 (N_4514,N_4213,N_4294);
and U4515 (N_4515,N_4292,N_4251);
or U4516 (N_4516,N_4303,N_4215);
nand U4517 (N_4517,N_4248,N_4241);
nor U4518 (N_4518,N_4365,N_4258);
nor U4519 (N_4519,N_4201,N_4310);
or U4520 (N_4520,N_4329,N_4328);
nor U4521 (N_4521,N_4234,N_4299);
and U4522 (N_4522,N_4355,N_4274);
nand U4523 (N_4523,N_4233,N_4287);
or U4524 (N_4524,N_4364,N_4397);
nor U4525 (N_4525,N_4257,N_4299);
nor U4526 (N_4526,N_4350,N_4228);
or U4527 (N_4527,N_4326,N_4237);
and U4528 (N_4528,N_4276,N_4277);
and U4529 (N_4529,N_4397,N_4212);
xor U4530 (N_4530,N_4224,N_4289);
nor U4531 (N_4531,N_4350,N_4262);
nor U4532 (N_4532,N_4394,N_4263);
and U4533 (N_4533,N_4237,N_4292);
and U4534 (N_4534,N_4336,N_4393);
and U4535 (N_4535,N_4213,N_4366);
and U4536 (N_4536,N_4269,N_4381);
nor U4537 (N_4537,N_4346,N_4275);
and U4538 (N_4538,N_4359,N_4340);
or U4539 (N_4539,N_4300,N_4331);
xnor U4540 (N_4540,N_4272,N_4244);
xor U4541 (N_4541,N_4314,N_4313);
nor U4542 (N_4542,N_4323,N_4368);
xor U4543 (N_4543,N_4275,N_4385);
or U4544 (N_4544,N_4202,N_4285);
xnor U4545 (N_4545,N_4310,N_4229);
nor U4546 (N_4546,N_4347,N_4385);
xor U4547 (N_4547,N_4256,N_4209);
and U4548 (N_4548,N_4214,N_4211);
xor U4549 (N_4549,N_4331,N_4285);
or U4550 (N_4550,N_4340,N_4389);
or U4551 (N_4551,N_4309,N_4207);
nand U4552 (N_4552,N_4207,N_4298);
and U4553 (N_4553,N_4324,N_4285);
nand U4554 (N_4554,N_4365,N_4344);
xor U4555 (N_4555,N_4280,N_4371);
nor U4556 (N_4556,N_4250,N_4202);
or U4557 (N_4557,N_4258,N_4383);
xnor U4558 (N_4558,N_4221,N_4346);
and U4559 (N_4559,N_4288,N_4377);
nand U4560 (N_4560,N_4322,N_4392);
xor U4561 (N_4561,N_4208,N_4395);
nor U4562 (N_4562,N_4312,N_4229);
nor U4563 (N_4563,N_4273,N_4234);
or U4564 (N_4564,N_4346,N_4297);
nand U4565 (N_4565,N_4245,N_4295);
nand U4566 (N_4566,N_4369,N_4225);
nand U4567 (N_4567,N_4383,N_4282);
nor U4568 (N_4568,N_4388,N_4265);
and U4569 (N_4569,N_4212,N_4279);
xor U4570 (N_4570,N_4365,N_4202);
nor U4571 (N_4571,N_4305,N_4300);
or U4572 (N_4572,N_4290,N_4222);
nand U4573 (N_4573,N_4212,N_4374);
nor U4574 (N_4574,N_4341,N_4222);
nand U4575 (N_4575,N_4212,N_4257);
nand U4576 (N_4576,N_4366,N_4228);
or U4577 (N_4577,N_4297,N_4311);
xnor U4578 (N_4578,N_4398,N_4331);
or U4579 (N_4579,N_4336,N_4231);
xor U4580 (N_4580,N_4217,N_4383);
xor U4581 (N_4581,N_4284,N_4382);
xor U4582 (N_4582,N_4323,N_4392);
nand U4583 (N_4583,N_4284,N_4296);
or U4584 (N_4584,N_4280,N_4236);
nand U4585 (N_4585,N_4223,N_4200);
xor U4586 (N_4586,N_4298,N_4237);
nor U4587 (N_4587,N_4214,N_4226);
or U4588 (N_4588,N_4354,N_4340);
nand U4589 (N_4589,N_4393,N_4344);
xor U4590 (N_4590,N_4254,N_4201);
and U4591 (N_4591,N_4223,N_4351);
xnor U4592 (N_4592,N_4233,N_4344);
nand U4593 (N_4593,N_4206,N_4225);
xor U4594 (N_4594,N_4209,N_4387);
nand U4595 (N_4595,N_4249,N_4247);
xor U4596 (N_4596,N_4281,N_4283);
xnor U4597 (N_4597,N_4204,N_4303);
nor U4598 (N_4598,N_4386,N_4209);
nand U4599 (N_4599,N_4277,N_4337);
or U4600 (N_4600,N_4462,N_4548);
nand U4601 (N_4601,N_4496,N_4402);
xnor U4602 (N_4602,N_4450,N_4498);
and U4603 (N_4603,N_4560,N_4489);
xnor U4604 (N_4604,N_4589,N_4501);
and U4605 (N_4605,N_4456,N_4454);
or U4606 (N_4606,N_4590,N_4538);
nor U4607 (N_4607,N_4470,N_4452);
and U4608 (N_4608,N_4484,N_4566);
xor U4609 (N_4609,N_4591,N_4451);
or U4610 (N_4610,N_4436,N_4431);
and U4611 (N_4611,N_4425,N_4417);
or U4612 (N_4612,N_4408,N_4435);
and U4613 (N_4613,N_4559,N_4532);
and U4614 (N_4614,N_4479,N_4426);
nand U4615 (N_4615,N_4552,N_4563);
nand U4616 (N_4616,N_4445,N_4570);
nor U4617 (N_4617,N_4550,N_4580);
nand U4618 (N_4618,N_4406,N_4473);
nand U4619 (N_4619,N_4593,N_4428);
nand U4620 (N_4620,N_4507,N_4515);
and U4621 (N_4621,N_4578,N_4551);
xnor U4622 (N_4622,N_4586,N_4516);
xor U4623 (N_4623,N_4485,N_4441);
and U4624 (N_4624,N_4467,N_4477);
xor U4625 (N_4625,N_4506,N_4519);
xnor U4626 (N_4626,N_4469,N_4493);
nor U4627 (N_4627,N_4424,N_4541);
and U4628 (N_4628,N_4529,N_4410);
xnor U4629 (N_4629,N_4434,N_4438);
xnor U4630 (N_4630,N_4474,N_4412);
or U4631 (N_4631,N_4416,N_4542);
nand U4632 (N_4632,N_4594,N_4413);
nor U4633 (N_4633,N_4584,N_4429);
xnor U4634 (N_4634,N_4405,N_4500);
or U4635 (N_4635,N_4403,N_4535);
and U4636 (N_4636,N_4433,N_4401);
and U4637 (N_4637,N_4585,N_4511);
nand U4638 (N_4638,N_4569,N_4597);
and U4639 (N_4639,N_4582,N_4508);
xor U4640 (N_4640,N_4531,N_4527);
nand U4641 (N_4641,N_4521,N_4545);
or U4642 (N_4642,N_4581,N_4573);
nand U4643 (N_4643,N_4502,N_4468);
xnor U4644 (N_4644,N_4514,N_4512);
xnor U4645 (N_4645,N_4517,N_4528);
or U4646 (N_4646,N_4430,N_4561);
xor U4647 (N_4647,N_4505,N_4455);
nor U4648 (N_4648,N_4458,N_4494);
xor U4649 (N_4649,N_4547,N_4453);
or U4650 (N_4650,N_4439,N_4557);
nand U4651 (N_4651,N_4504,N_4525);
xor U4652 (N_4652,N_4558,N_4432);
or U4653 (N_4653,N_4556,N_4411);
nand U4654 (N_4654,N_4440,N_4554);
xor U4655 (N_4655,N_4568,N_4419);
or U4656 (N_4656,N_4534,N_4520);
xor U4657 (N_4657,N_4478,N_4421);
and U4658 (N_4658,N_4487,N_4409);
xnor U4659 (N_4659,N_4472,N_4539);
or U4660 (N_4660,N_4464,N_4588);
or U4661 (N_4661,N_4459,N_4457);
nand U4662 (N_4662,N_4526,N_4461);
and U4663 (N_4663,N_4447,N_4481);
xnor U4664 (N_4664,N_4446,N_4510);
or U4665 (N_4665,N_4466,N_4407);
or U4666 (N_4666,N_4476,N_4595);
or U4667 (N_4667,N_4488,N_4444);
or U4668 (N_4668,N_4567,N_4486);
xor U4669 (N_4669,N_4583,N_4443);
nand U4670 (N_4670,N_4490,N_4503);
and U4671 (N_4671,N_4564,N_4449);
nor U4672 (N_4672,N_4579,N_4418);
and U4673 (N_4673,N_4513,N_4483);
nand U4674 (N_4674,N_4442,N_4596);
xor U4675 (N_4675,N_4465,N_4518);
nand U4676 (N_4676,N_4562,N_4460);
and U4677 (N_4677,N_4423,N_4509);
or U4678 (N_4678,N_4599,N_4471);
xnor U4679 (N_4679,N_4524,N_4575);
and U4680 (N_4680,N_4422,N_4544);
nor U4681 (N_4681,N_4530,N_4495);
nor U4682 (N_4682,N_4522,N_4546);
nand U4683 (N_4683,N_4553,N_4414);
and U4684 (N_4684,N_4480,N_4448);
or U4685 (N_4685,N_4565,N_4499);
xor U4686 (N_4686,N_4492,N_4415);
nor U4687 (N_4687,N_4523,N_4587);
nand U4688 (N_4688,N_4536,N_4543);
or U4689 (N_4689,N_4577,N_4475);
or U4690 (N_4690,N_4537,N_4576);
nor U4691 (N_4691,N_4549,N_4540);
or U4692 (N_4692,N_4574,N_4491);
nor U4693 (N_4693,N_4592,N_4427);
and U4694 (N_4694,N_4404,N_4555);
and U4695 (N_4695,N_4482,N_4533);
nor U4696 (N_4696,N_4400,N_4571);
or U4697 (N_4697,N_4497,N_4598);
nor U4698 (N_4698,N_4420,N_4463);
nor U4699 (N_4699,N_4572,N_4437);
and U4700 (N_4700,N_4522,N_4479);
and U4701 (N_4701,N_4436,N_4550);
nand U4702 (N_4702,N_4570,N_4568);
and U4703 (N_4703,N_4459,N_4565);
nand U4704 (N_4704,N_4409,N_4430);
nand U4705 (N_4705,N_4583,N_4480);
nor U4706 (N_4706,N_4454,N_4582);
or U4707 (N_4707,N_4588,N_4557);
nor U4708 (N_4708,N_4422,N_4564);
and U4709 (N_4709,N_4509,N_4584);
nor U4710 (N_4710,N_4524,N_4500);
xor U4711 (N_4711,N_4485,N_4546);
nand U4712 (N_4712,N_4413,N_4440);
and U4713 (N_4713,N_4411,N_4507);
nor U4714 (N_4714,N_4560,N_4471);
xnor U4715 (N_4715,N_4569,N_4590);
xor U4716 (N_4716,N_4470,N_4420);
nand U4717 (N_4717,N_4446,N_4440);
or U4718 (N_4718,N_4517,N_4410);
nand U4719 (N_4719,N_4488,N_4496);
and U4720 (N_4720,N_4526,N_4500);
nor U4721 (N_4721,N_4474,N_4546);
nand U4722 (N_4722,N_4479,N_4470);
and U4723 (N_4723,N_4412,N_4511);
or U4724 (N_4724,N_4435,N_4501);
and U4725 (N_4725,N_4523,N_4558);
nand U4726 (N_4726,N_4491,N_4566);
xor U4727 (N_4727,N_4594,N_4556);
xnor U4728 (N_4728,N_4421,N_4560);
xor U4729 (N_4729,N_4550,N_4431);
or U4730 (N_4730,N_4442,N_4481);
xor U4731 (N_4731,N_4430,N_4421);
or U4732 (N_4732,N_4508,N_4511);
or U4733 (N_4733,N_4518,N_4533);
or U4734 (N_4734,N_4488,N_4593);
or U4735 (N_4735,N_4554,N_4446);
nand U4736 (N_4736,N_4568,N_4533);
or U4737 (N_4737,N_4446,N_4556);
and U4738 (N_4738,N_4534,N_4505);
and U4739 (N_4739,N_4431,N_4598);
xnor U4740 (N_4740,N_4492,N_4504);
xnor U4741 (N_4741,N_4574,N_4423);
nor U4742 (N_4742,N_4493,N_4550);
xnor U4743 (N_4743,N_4583,N_4455);
nor U4744 (N_4744,N_4491,N_4480);
and U4745 (N_4745,N_4462,N_4443);
nor U4746 (N_4746,N_4574,N_4560);
and U4747 (N_4747,N_4405,N_4564);
or U4748 (N_4748,N_4434,N_4478);
nor U4749 (N_4749,N_4546,N_4597);
nor U4750 (N_4750,N_4591,N_4523);
and U4751 (N_4751,N_4549,N_4568);
xnor U4752 (N_4752,N_4423,N_4442);
xor U4753 (N_4753,N_4429,N_4420);
and U4754 (N_4754,N_4451,N_4549);
nor U4755 (N_4755,N_4575,N_4574);
nand U4756 (N_4756,N_4543,N_4417);
or U4757 (N_4757,N_4483,N_4480);
xor U4758 (N_4758,N_4539,N_4469);
and U4759 (N_4759,N_4575,N_4440);
nand U4760 (N_4760,N_4582,N_4561);
and U4761 (N_4761,N_4462,N_4565);
xor U4762 (N_4762,N_4421,N_4543);
xnor U4763 (N_4763,N_4549,N_4556);
xnor U4764 (N_4764,N_4412,N_4445);
nor U4765 (N_4765,N_4581,N_4593);
xor U4766 (N_4766,N_4456,N_4486);
nand U4767 (N_4767,N_4417,N_4414);
nor U4768 (N_4768,N_4410,N_4491);
nor U4769 (N_4769,N_4522,N_4496);
xor U4770 (N_4770,N_4429,N_4520);
nor U4771 (N_4771,N_4483,N_4599);
nor U4772 (N_4772,N_4523,N_4409);
and U4773 (N_4773,N_4533,N_4481);
nand U4774 (N_4774,N_4572,N_4551);
or U4775 (N_4775,N_4550,N_4501);
or U4776 (N_4776,N_4499,N_4444);
nand U4777 (N_4777,N_4588,N_4543);
and U4778 (N_4778,N_4523,N_4566);
xnor U4779 (N_4779,N_4517,N_4462);
and U4780 (N_4780,N_4458,N_4431);
nand U4781 (N_4781,N_4554,N_4506);
nand U4782 (N_4782,N_4523,N_4567);
and U4783 (N_4783,N_4513,N_4557);
xor U4784 (N_4784,N_4453,N_4468);
or U4785 (N_4785,N_4580,N_4514);
xor U4786 (N_4786,N_4407,N_4484);
or U4787 (N_4787,N_4512,N_4421);
nor U4788 (N_4788,N_4577,N_4522);
and U4789 (N_4789,N_4472,N_4459);
xnor U4790 (N_4790,N_4544,N_4522);
and U4791 (N_4791,N_4549,N_4459);
xor U4792 (N_4792,N_4482,N_4505);
or U4793 (N_4793,N_4558,N_4497);
or U4794 (N_4794,N_4468,N_4484);
nor U4795 (N_4795,N_4428,N_4425);
nand U4796 (N_4796,N_4484,N_4408);
xnor U4797 (N_4797,N_4408,N_4547);
nor U4798 (N_4798,N_4517,N_4497);
nand U4799 (N_4799,N_4450,N_4493);
and U4800 (N_4800,N_4765,N_4799);
nand U4801 (N_4801,N_4632,N_4742);
xnor U4802 (N_4802,N_4797,N_4711);
nand U4803 (N_4803,N_4788,N_4717);
xnor U4804 (N_4804,N_4636,N_4787);
nand U4805 (N_4805,N_4624,N_4757);
or U4806 (N_4806,N_4772,N_4657);
or U4807 (N_4807,N_4782,N_4650);
nor U4808 (N_4808,N_4625,N_4667);
nand U4809 (N_4809,N_4732,N_4677);
xor U4810 (N_4810,N_4603,N_4694);
and U4811 (N_4811,N_4722,N_4723);
or U4812 (N_4812,N_4780,N_4708);
nor U4813 (N_4813,N_4674,N_4726);
and U4814 (N_4814,N_4737,N_4704);
and U4815 (N_4815,N_4622,N_4621);
nand U4816 (N_4816,N_4763,N_4796);
nand U4817 (N_4817,N_4658,N_4756);
or U4818 (N_4818,N_4781,N_4750);
nor U4819 (N_4819,N_4664,N_4649);
nor U4820 (N_4820,N_4633,N_4647);
nor U4821 (N_4821,N_4689,N_4612);
nand U4822 (N_4822,N_4734,N_4604);
or U4823 (N_4823,N_4709,N_4776);
nand U4824 (N_4824,N_4699,N_4627);
nand U4825 (N_4825,N_4693,N_4631);
nand U4826 (N_4826,N_4740,N_4754);
or U4827 (N_4827,N_4751,N_4659);
nand U4828 (N_4828,N_4798,N_4638);
xor U4829 (N_4829,N_4626,N_4613);
nor U4830 (N_4830,N_4702,N_4660);
and U4831 (N_4831,N_4630,N_4792);
nand U4832 (N_4832,N_4785,N_4706);
xor U4833 (N_4833,N_4628,N_4645);
and U4834 (N_4834,N_4789,N_4730);
nand U4835 (N_4835,N_4681,N_4771);
nand U4836 (N_4836,N_4703,N_4713);
nand U4837 (N_4837,N_4680,N_4602);
xnor U4838 (N_4838,N_4675,N_4715);
nor U4839 (N_4839,N_4767,N_4769);
nand U4840 (N_4840,N_4768,N_4779);
xnor U4841 (N_4841,N_4774,N_4710);
nor U4842 (N_4842,N_4770,N_4784);
xnor U4843 (N_4843,N_4644,N_4727);
or U4844 (N_4844,N_4705,N_4795);
nand U4845 (N_4845,N_4725,N_4643);
nand U4846 (N_4846,N_4775,N_4696);
nand U4847 (N_4847,N_4718,N_4752);
or U4848 (N_4848,N_4679,N_4669);
nand U4849 (N_4849,N_4648,N_4688);
nand U4850 (N_4850,N_4651,N_4716);
nor U4851 (N_4851,N_4623,N_4684);
and U4852 (N_4852,N_4692,N_4783);
nor U4853 (N_4853,N_4618,N_4791);
and U4854 (N_4854,N_4652,N_4794);
and U4855 (N_4855,N_4668,N_4655);
and U4856 (N_4856,N_4761,N_4637);
nor U4857 (N_4857,N_4665,N_4673);
xnor U4858 (N_4858,N_4685,N_4615);
nor U4859 (N_4859,N_4753,N_4605);
xnor U4860 (N_4860,N_4641,N_4646);
or U4861 (N_4861,N_4707,N_4634);
and U4862 (N_4862,N_4616,N_4642);
nand U4863 (N_4863,N_4639,N_4683);
and U4864 (N_4864,N_4661,N_4629);
nand U4865 (N_4865,N_4608,N_4666);
and U4866 (N_4866,N_4773,N_4720);
xor U4867 (N_4867,N_4676,N_4747);
nand U4868 (N_4868,N_4698,N_4697);
nor U4869 (N_4869,N_4714,N_4728);
nor U4870 (N_4870,N_4620,N_4744);
nor U4871 (N_4871,N_4712,N_4764);
or U4872 (N_4872,N_4724,N_4609);
and U4873 (N_4873,N_4601,N_4741);
and U4874 (N_4874,N_4758,N_4760);
xnor U4875 (N_4875,N_4729,N_4738);
and U4876 (N_4876,N_4653,N_4766);
and U4877 (N_4877,N_4721,N_4619);
or U4878 (N_4878,N_4790,N_4793);
nand U4879 (N_4879,N_4614,N_4762);
or U4880 (N_4880,N_4607,N_4663);
nand U4881 (N_4881,N_4719,N_4686);
and U4882 (N_4882,N_4670,N_4749);
or U4883 (N_4883,N_4748,N_4662);
xnor U4884 (N_4884,N_4640,N_4736);
nor U4885 (N_4885,N_4778,N_4672);
or U4886 (N_4886,N_4735,N_4777);
or U4887 (N_4887,N_4786,N_4700);
nor U4888 (N_4888,N_4755,N_4687);
and U4889 (N_4889,N_4745,N_4654);
nor U4890 (N_4890,N_4611,N_4743);
xnor U4891 (N_4891,N_4682,N_4690);
nor U4892 (N_4892,N_4600,N_4617);
nor U4893 (N_4893,N_4701,N_4635);
nor U4894 (N_4894,N_4759,N_4656);
nor U4895 (N_4895,N_4606,N_4691);
nor U4896 (N_4896,N_4678,N_4731);
nand U4897 (N_4897,N_4733,N_4746);
or U4898 (N_4898,N_4695,N_4739);
or U4899 (N_4899,N_4671,N_4610);
xor U4900 (N_4900,N_4677,N_4656);
or U4901 (N_4901,N_4643,N_4711);
and U4902 (N_4902,N_4788,N_4769);
xnor U4903 (N_4903,N_4654,N_4659);
or U4904 (N_4904,N_4661,N_4767);
and U4905 (N_4905,N_4666,N_4768);
nor U4906 (N_4906,N_4759,N_4799);
nand U4907 (N_4907,N_4736,N_4683);
or U4908 (N_4908,N_4677,N_4660);
or U4909 (N_4909,N_4760,N_4713);
xnor U4910 (N_4910,N_4679,N_4600);
nand U4911 (N_4911,N_4795,N_4622);
and U4912 (N_4912,N_4667,N_4766);
nand U4913 (N_4913,N_4749,N_4613);
xor U4914 (N_4914,N_4739,N_4645);
nand U4915 (N_4915,N_4643,N_4620);
or U4916 (N_4916,N_4600,N_4639);
or U4917 (N_4917,N_4623,N_4788);
nor U4918 (N_4918,N_4715,N_4685);
or U4919 (N_4919,N_4624,N_4628);
and U4920 (N_4920,N_4703,N_4789);
xor U4921 (N_4921,N_4605,N_4760);
nand U4922 (N_4922,N_4734,N_4627);
xnor U4923 (N_4923,N_4759,N_4771);
and U4924 (N_4924,N_4706,N_4705);
and U4925 (N_4925,N_4705,N_4605);
nor U4926 (N_4926,N_4752,N_4648);
xor U4927 (N_4927,N_4680,N_4692);
and U4928 (N_4928,N_4622,N_4752);
or U4929 (N_4929,N_4714,N_4799);
xor U4930 (N_4930,N_4701,N_4716);
nand U4931 (N_4931,N_4747,N_4659);
or U4932 (N_4932,N_4701,N_4736);
nor U4933 (N_4933,N_4605,N_4675);
xnor U4934 (N_4934,N_4680,N_4654);
nand U4935 (N_4935,N_4771,N_4665);
and U4936 (N_4936,N_4789,N_4674);
xor U4937 (N_4937,N_4705,N_4718);
xor U4938 (N_4938,N_4731,N_4616);
nand U4939 (N_4939,N_4617,N_4661);
nand U4940 (N_4940,N_4636,N_4682);
nand U4941 (N_4941,N_4747,N_4664);
or U4942 (N_4942,N_4637,N_4690);
or U4943 (N_4943,N_4778,N_4742);
nand U4944 (N_4944,N_4710,N_4606);
xnor U4945 (N_4945,N_4677,N_4696);
or U4946 (N_4946,N_4717,N_4695);
or U4947 (N_4947,N_4699,N_4762);
or U4948 (N_4948,N_4787,N_4681);
or U4949 (N_4949,N_4669,N_4724);
nor U4950 (N_4950,N_4654,N_4770);
and U4951 (N_4951,N_4706,N_4738);
xnor U4952 (N_4952,N_4719,N_4646);
nand U4953 (N_4953,N_4636,N_4789);
nand U4954 (N_4954,N_4667,N_4779);
and U4955 (N_4955,N_4774,N_4642);
and U4956 (N_4956,N_4637,N_4738);
and U4957 (N_4957,N_4606,N_4628);
nand U4958 (N_4958,N_4618,N_4662);
and U4959 (N_4959,N_4766,N_4798);
xor U4960 (N_4960,N_4706,N_4735);
nand U4961 (N_4961,N_4636,N_4709);
nor U4962 (N_4962,N_4747,N_4662);
or U4963 (N_4963,N_4719,N_4704);
xnor U4964 (N_4964,N_4647,N_4782);
nor U4965 (N_4965,N_4795,N_4654);
and U4966 (N_4966,N_4633,N_4736);
nand U4967 (N_4967,N_4714,N_4639);
xor U4968 (N_4968,N_4709,N_4642);
nor U4969 (N_4969,N_4738,N_4717);
and U4970 (N_4970,N_4683,N_4794);
or U4971 (N_4971,N_4661,N_4643);
or U4972 (N_4972,N_4680,N_4669);
xnor U4973 (N_4973,N_4780,N_4773);
nor U4974 (N_4974,N_4602,N_4613);
and U4975 (N_4975,N_4701,N_4638);
nand U4976 (N_4976,N_4694,N_4605);
and U4977 (N_4977,N_4782,N_4730);
xor U4978 (N_4978,N_4615,N_4645);
xor U4979 (N_4979,N_4609,N_4793);
nor U4980 (N_4980,N_4698,N_4715);
or U4981 (N_4981,N_4795,N_4638);
xnor U4982 (N_4982,N_4600,N_4659);
and U4983 (N_4983,N_4675,N_4691);
nor U4984 (N_4984,N_4779,N_4710);
nor U4985 (N_4985,N_4713,N_4691);
or U4986 (N_4986,N_4653,N_4643);
nor U4987 (N_4987,N_4649,N_4799);
or U4988 (N_4988,N_4607,N_4606);
nor U4989 (N_4989,N_4726,N_4631);
xor U4990 (N_4990,N_4755,N_4749);
nand U4991 (N_4991,N_4754,N_4747);
or U4992 (N_4992,N_4675,N_4629);
and U4993 (N_4993,N_4649,N_4702);
nor U4994 (N_4994,N_4721,N_4635);
and U4995 (N_4995,N_4671,N_4642);
nor U4996 (N_4996,N_4719,N_4635);
or U4997 (N_4997,N_4731,N_4768);
nor U4998 (N_4998,N_4614,N_4671);
and U4999 (N_4999,N_4615,N_4629);
xnor U5000 (N_5000,N_4960,N_4922);
or U5001 (N_5001,N_4987,N_4804);
nand U5002 (N_5002,N_4835,N_4882);
nand U5003 (N_5003,N_4982,N_4891);
or U5004 (N_5004,N_4967,N_4810);
nand U5005 (N_5005,N_4808,N_4876);
xor U5006 (N_5006,N_4895,N_4947);
or U5007 (N_5007,N_4825,N_4873);
and U5008 (N_5008,N_4986,N_4926);
nor U5009 (N_5009,N_4814,N_4829);
xnor U5010 (N_5010,N_4815,N_4856);
xnor U5011 (N_5011,N_4853,N_4910);
and U5012 (N_5012,N_4962,N_4978);
or U5013 (N_5013,N_4937,N_4846);
nor U5014 (N_5014,N_4819,N_4865);
nor U5015 (N_5015,N_4858,N_4953);
or U5016 (N_5016,N_4852,N_4823);
and U5017 (N_5017,N_4948,N_4806);
and U5018 (N_5018,N_4955,N_4870);
and U5019 (N_5019,N_4826,N_4929);
and U5020 (N_5020,N_4924,N_4941);
nand U5021 (N_5021,N_4972,N_4965);
xor U5022 (N_5022,N_4800,N_4921);
nand U5023 (N_5023,N_4887,N_4914);
nor U5024 (N_5024,N_4863,N_4818);
nand U5025 (N_5025,N_4973,N_4862);
xor U5026 (N_5026,N_4899,N_4961);
nor U5027 (N_5027,N_4954,N_4837);
and U5028 (N_5028,N_4822,N_4974);
or U5029 (N_5029,N_4999,N_4970);
xnor U5030 (N_5030,N_4983,N_4904);
xnor U5031 (N_5031,N_4851,N_4908);
and U5032 (N_5032,N_4885,N_4848);
and U5033 (N_5033,N_4913,N_4864);
or U5034 (N_5034,N_4884,N_4945);
and U5035 (N_5035,N_4952,N_4944);
and U5036 (N_5036,N_4838,N_4934);
and U5037 (N_5037,N_4993,N_4812);
nor U5038 (N_5038,N_4989,N_4869);
and U5039 (N_5039,N_4907,N_4988);
xnor U5040 (N_5040,N_4839,N_4919);
nor U5041 (N_5041,N_4963,N_4977);
nand U5042 (N_5042,N_4828,N_4903);
nor U5043 (N_5043,N_4866,N_4992);
or U5044 (N_5044,N_4811,N_4893);
xor U5045 (N_5045,N_4894,N_4824);
and U5046 (N_5046,N_4942,N_4997);
nand U5047 (N_5047,N_4998,N_4832);
and U5048 (N_5048,N_4880,N_4949);
or U5049 (N_5049,N_4816,N_4917);
nor U5050 (N_5050,N_4861,N_4813);
xor U5051 (N_5051,N_4990,N_4860);
and U5052 (N_5052,N_4807,N_4984);
nor U5053 (N_5053,N_4821,N_4896);
or U5054 (N_5054,N_4831,N_4802);
nor U5055 (N_5055,N_4820,N_4902);
and U5056 (N_5056,N_4956,N_4809);
nor U5057 (N_5057,N_4938,N_4971);
nand U5058 (N_5058,N_4918,N_4900);
or U5059 (N_5059,N_4923,N_4901);
nand U5060 (N_5060,N_4964,N_4827);
nand U5061 (N_5061,N_4991,N_4817);
nor U5062 (N_5062,N_4981,N_4927);
nor U5063 (N_5063,N_4881,N_4875);
or U5064 (N_5064,N_4912,N_4878);
or U5065 (N_5065,N_4872,N_4833);
nor U5066 (N_5066,N_4888,N_4975);
or U5067 (N_5067,N_4877,N_4844);
nor U5068 (N_5068,N_4871,N_4957);
and U5069 (N_5069,N_4980,N_4879);
nor U5070 (N_5070,N_4803,N_4946);
or U5071 (N_5071,N_4897,N_4847);
and U5072 (N_5072,N_4976,N_4849);
and U5073 (N_5073,N_4950,N_4905);
or U5074 (N_5074,N_4909,N_4898);
and U5075 (N_5075,N_4841,N_4834);
nand U5076 (N_5076,N_4933,N_4855);
nor U5077 (N_5077,N_4892,N_4936);
nor U5078 (N_5078,N_4925,N_4940);
nor U5079 (N_5079,N_4883,N_4943);
xnor U5080 (N_5080,N_4857,N_4915);
and U5081 (N_5081,N_4836,N_4935);
and U5082 (N_5082,N_4995,N_4868);
and U5083 (N_5083,N_4985,N_4845);
xnor U5084 (N_5084,N_4906,N_4979);
nor U5085 (N_5085,N_4890,N_4959);
or U5086 (N_5086,N_4854,N_4928);
nand U5087 (N_5087,N_4920,N_4911);
nor U5088 (N_5088,N_4931,N_4958);
nor U5089 (N_5089,N_4969,N_4939);
nand U5090 (N_5090,N_4932,N_4930);
xnor U5091 (N_5091,N_4968,N_4805);
and U5092 (N_5092,N_4850,N_4996);
and U5093 (N_5093,N_4916,N_4951);
nor U5094 (N_5094,N_4994,N_4840);
or U5095 (N_5095,N_4859,N_4867);
nand U5096 (N_5096,N_4842,N_4830);
and U5097 (N_5097,N_4801,N_4889);
and U5098 (N_5098,N_4886,N_4874);
nor U5099 (N_5099,N_4843,N_4966);
nand U5100 (N_5100,N_4962,N_4922);
nor U5101 (N_5101,N_4893,N_4803);
nand U5102 (N_5102,N_4927,N_4918);
xor U5103 (N_5103,N_4866,N_4829);
xnor U5104 (N_5104,N_4972,N_4968);
nand U5105 (N_5105,N_4816,N_4985);
nor U5106 (N_5106,N_4959,N_4834);
xnor U5107 (N_5107,N_4820,N_4885);
nor U5108 (N_5108,N_4943,N_4904);
nor U5109 (N_5109,N_4842,N_4934);
and U5110 (N_5110,N_4821,N_4918);
or U5111 (N_5111,N_4821,N_4810);
xor U5112 (N_5112,N_4872,N_4824);
and U5113 (N_5113,N_4936,N_4804);
or U5114 (N_5114,N_4976,N_4971);
nand U5115 (N_5115,N_4924,N_4863);
nand U5116 (N_5116,N_4919,N_4993);
nor U5117 (N_5117,N_4999,N_4951);
nand U5118 (N_5118,N_4836,N_4843);
nand U5119 (N_5119,N_4908,N_4955);
xor U5120 (N_5120,N_4848,N_4831);
or U5121 (N_5121,N_4820,N_4869);
nand U5122 (N_5122,N_4908,N_4863);
and U5123 (N_5123,N_4885,N_4915);
or U5124 (N_5124,N_4806,N_4980);
or U5125 (N_5125,N_4828,N_4944);
xor U5126 (N_5126,N_4863,N_4817);
nor U5127 (N_5127,N_4805,N_4848);
xnor U5128 (N_5128,N_4866,N_4823);
and U5129 (N_5129,N_4953,N_4865);
nor U5130 (N_5130,N_4966,N_4922);
nand U5131 (N_5131,N_4992,N_4831);
and U5132 (N_5132,N_4885,N_4923);
xor U5133 (N_5133,N_4980,N_4889);
nor U5134 (N_5134,N_4828,N_4934);
nand U5135 (N_5135,N_4859,N_4802);
xnor U5136 (N_5136,N_4813,N_4834);
nand U5137 (N_5137,N_4863,N_4865);
nand U5138 (N_5138,N_4853,N_4842);
and U5139 (N_5139,N_4878,N_4857);
nor U5140 (N_5140,N_4829,N_4834);
nand U5141 (N_5141,N_4959,N_4833);
and U5142 (N_5142,N_4834,N_4833);
nor U5143 (N_5143,N_4874,N_4804);
xor U5144 (N_5144,N_4919,N_4805);
nand U5145 (N_5145,N_4860,N_4995);
nand U5146 (N_5146,N_4909,N_4986);
nand U5147 (N_5147,N_4830,N_4961);
nor U5148 (N_5148,N_4911,N_4960);
xnor U5149 (N_5149,N_4899,N_4914);
nor U5150 (N_5150,N_4895,N_4862);
or U5151 (N_5151,N_4885,N_4888);
xnor U5152 (N_5152,N_4819,N_4882);
and U5153 (N_5153,N_4840,N_4935);
nand U5154 (N_5154,N_4908,N_4930);
nor U5155 (N_5155,N_4840,N_4837);
and U5156 (N_5156,N_4923,N_4910);
nor U5157 (N_5157,N_4901,N_4819);
or U5158 (N_5158,N_4979,N_4869);
or U5159 (N_5159,N_4801,N_4962);
nor U5160 (N_5160,N_4941,N_4806);
or U5161 (N_5161,N_4921,N_4955);
nand U5162 (N_5162,N_4879,N_4867);
nor U5163 (N_5163,N_4954,N_4937);
nor U5164 (N_5164,N_4893,N_4935);
nand U5165 (N_5165,N_4934,N_4974);
nor U5166 (N_5166,N_4901,N_4848);
and U5167 (N_5167,N_4887,N_4969);
xor U5168 (N_5168,N_4898,N_4923);
and U5169 (N_5169,N_4814,N_4961);
and U5170 (N_5170,N_4818,N_4934);
nor U5171 (N_5171,N_4866,N_4907);
and U5172 (N_5172,N_4965,N_4923);
nand U5173 (N_5173,N_4923,N_4803);
xor U5174 (N_5174,N_4937,N_4959);
or U5175 (N_5175,N_4822,N_4878);
xor U5176 (N_5176,N_4840,N_4980);
nor U5177 (N_5177,N_4971,N_4880);
or U5178 (N_5178,N_4868,N_4815);
nor U5179 (N_5179,N_4854,N_4824);
or U5180 (N_5180,N_4962,N_4807);
or U5181 (N_5181,N_4938,N_4920);
nor U5182 (N_5182,N_4823,N_4989);
xnor U5183 (N_5183,N_4911,N_4885);
and U5184 (N_5184,N_4892,N_4956);
nand U5185 (N_5185,N_4910,N_4886);
nor U5186 (N_5186,N_4914,N_4863);
and U5187 (N_5187,N_4878,N_4815);
nor U5188 (N_5188,N_4952,N_4922);
or U5189 (N_5189,N_4935,N_4913);
and U5190 (N_5190,N_4841,N_4979);
nor U5191 (N_5191,N_4930,N_4961);
and U5192 (N_5192,N_4863,N_4824);
and U5193 (N_5193,N_4868,N_4829);
nand U5194 (N_5194,N_4917,N_4843);
xnor U5195 (N_5195,N_4983,N_4841);
or U5196 (N_5196,N_4934,N_4933);
xnor U5197 (N_5197,N_4997,N_4800);
nand U5198 (N_5198,N_4819,N_4911);
and U5199 (N_5199,N_4924,N_4950);
nand U5200 (N_5200,N_5189,N_5024);
and U5201 (N_5201,N_5180,N_5140);
and U5202 (N_5202,N_5162,N_5060);
xor U5203 (N_5203,N_5093,N_5037);
or U5204 (N_5204,N_5100,N_5169);
nor U5205 (N_5205,N_5139,N_5161);
nand U5206 (N_5206,N_5195,N_5194);
or U5207 (N_5207,N_5167,N_5111);
xnor U5208 (N_5208,N_5187,N_5062);
and U5209 (N_5209,N_5008,N_5001);
xnor U5210 (N_5210,N_5102,N_5063);
nand U5211 (N_5211,N_5096,N_5020);
and U5212 (N_5212,N_5079,N_5071);
nand U5213 (N_5213,N_5085,N_5122);
nor U5214 (N_5214,N_5154,N_5164);
xnor U5215 (N_5215,N_5192,N_5081);
nand U5216 (N_5216,N_5105,N_5197);
nand U5217 (N_5217,N_5053,N_5070);
nand U5218 (N_5218,N_5023,N_5091);
and U5219 (N_5219,N_5014,N_5098);
nand U5220 (N_5220,N_5087,N_5134);
xor U5221 (N_5221,N_5006,N_5109);
or U5222 (N_5222,N_5160,N_5196);
xor U5223 (N_5223,N_5086,N_5115);
and U5224 (N_5224,N_5147,N_5151);
xnor U5225 (N_5225,N_5009,N_5120);
and U5226 (N_5226,N_5051,N_5157);
or U5227 (N_5227,N_5099,N_5042);
nor U5228 (N_5228,N_5002,N_5004);
nor U5229 (N_5229,N_5121,N_5017);
nor U5230 (N_5230,N_5034,N_5123);
and U5231 (N_5231,N_5144,N_5191);
xor U5232 (N_5232,N_5156,N_5043);
nand U5233 (N_5233,N_5010,N_5097);
nand U5234 (N_5234,N_5084,N_5049);
and U5235 (N_5235,N_5132,N_5103);
nor U5236 (N_5236,N_5107,N_5124);
and U5237 (N_5237,N_5035,N_5118);
xnor U5238 (N_5238,N_5176,N_5059);
nand U5239 (N_5239,N_5128,N_5054);
or U5240 (N_5240,N_5005,N_5150);
nor U5241 (N_5241,N_5031,N_5052);
nor U5242 (N_5242,N_5028,N_5072);
nor U5243 (N_5243,N_5003,N_5044);
nor U5244 (N_5244,N_5074,N_5145);
xnor U5245 (N_5245,N_5050,N_5159);
xor U5246 (N_5246,N_5078,N_5116);
xor U5247 (N_5247,N_5068,N_5090);
xor U5248 (N_5248,N_5033,N_5185);
nor U5249 (N_5249,N_5088,N_5015);
or U5250 (N_5250,N_5061,N_5125);
nand U5251 (N_5251,N_5165,N_5178);
or U5252 (N_5252,N_5025,N_5018);
xor U5253 (N_5253,N_5114,N_5193);
xor U5254 (N_5254,N_5137,N_5146);
xnor U5255 (N_5255,N_5179,N_5141);
or U5256 (N_5256,N_5110,N_5027);
nor U5257 (N_5257,N_5152,N_5127);
and U5258 (N_5258,N_5000,N_5011);
xnor U5259 (N_5259,N_5066,N_5155);
xnor U5260 (N_5260,N_5058,N_5199);
nor U5261 (N_5261,N_5126,N_5065);
nand U5262 (N_5262,N_5198,N_5131);
xor U5263 (N_5263,N_5183,N_5177);
nor U5264 (N_5264,N_5175,N_5013);
nand U5265 (N_5265,N_5092,N_5032);
or U5266 (N_5266,N_5045,N_5046);
nor U5267 (N_5267,N_5184,N_5101);
and U5268 (N_5268,N_5073,N_5026);
nor U5269 (N_5269,N_5036,N_5148);
nor U5270 (N_5270,N_5182,N_5064);
and U5271 (N_5271,N_5158,N_5174);
xnor U5272 (N_5272,N_5048,N_5094);
and U5273 (N_5273,N_5080,N_5047);
and U5274 (N_5274,N_5149,N_5168);
nand U5275 (N_5275,N_5038,N_5112);
xor U5276 (N_5276,N_5119,N_5057);
xor U5277 (N_5277,N_5130,N_5012);
xnor U5278 (N_5278,N_5019,N_5089);
nor U5279 (N_5279,N_5021,N_5083);
xnor U5280 (N_5280,N_5143,N_5163);
and U5281 (N_5281,N_5142,N_5172);
xnor U5282 (N_5282,N_5082,N_5166);
nor U5283 (N_5283,N_5153,N_5040);
nor U5284 (N_5284,N_5181,N_5188);
nor U5285 (N_5285,N_5039,N_5022);
nor U5286 (N_5286,N_5117,N_5056);
nand U5287 (N_5287,N_5030,N_5007);
xnor U5288 (N_5288,N_5076,N_5069);
xor U5289 (N_5289,N_5055,N_5106);
nand U5290 (N_5290,N_5129,N_5135);
nand U5291 (N_5291,N_5075,N_5041);
nor U5292 (N_5292,N_5029,N_5171);
nand U5293 (N_5293,N_5186,N_5170);
xnor U5294 (N_5294,N_5077,N_5016);
nand U5295 (N_5295,N_5190,N_5136);
nor U5296 (N_5296,N_5173,N_5133);
nand U5297 (N_5297,N_5095,N_5104);
nor U5298 (N_5298,N_5108,N_5138);
nor U5299 (N_5299,N_5067,N_5113);
xor U5300 (N_5300,N_5182,N_5010);
or U5301 (N_5301,N_5005,N_5177);
xor U5302 (N_5302,N_5014,N_5085);
xnor U5303 (N_5303,N_5011,N_5161);
or U5304 (N_5304,N_5064,N_5124);
xor U5305 (N_5305,N_5045,N_5031);
and U5306 (N_5306,N_5004,N_5059);
and U5307 (N_5307,N_5019,N_5048);
xor U5308 (N_5308,N_5192,N_5011);
nor U5309 (N_5309,N_5054,N_5028);
nand U5310 (N_5310,N_5188,N_5015);
and U5311 (N_5311,N_5038,N_5178);
nand U5312 (N_5312,N_5190,N_5084);
or U5313 (N_5313,N_5103,N_5199);
xor U5314 (N_5314,N_5111,N_5069);
and U5315 (N_5315,N_5170,N_5182);
or U5316 (N_5316,N_5167,N_5176);
and U5317 (N_5317,N_5092,N_5076);
nor U5318 (N_5318,N_5176,N_5087);
nand U5319 (N_5319,N_5085,N_5136);
nor U5320 (N_5320,N_5056,N_5181);
xnor U5321 (N_5321,N_5162,N_5043);
and U5322 (N_5322,N_5122,N_5024);
and U5323 (N_5323,N_5106,N_5056);
and U5324 (N_5324,N_5084,N_5179);
or U5325 (N_5325,N_5062,N_5146);
nor U5326 (N_5326,N_5107,N_5114);
xor U5327 (N_5327,N_5189,N_5172);
nor U5328 (N_5328,N_5175,N_5102);
or U5329 (N_5329,N_5037,N_5192);
or U5330 (N_5330,N_5124,N_5083);
or U5331 (N_5331,N_5098,N_5181);
nand U5332 (N_5332,N_5192,N_5091);
or U5333 (N_5333,N_5180,N_5021);
and U5334 (N_5334,N_5087,N_5169);
xor U5335 (N_5335,N_5154,N_5007);
nand U5336 (N_5336,N_5169,N_5190);
nand U5337 (N_5337,N_5186,N_5162);
nor U5338 (N_5338,N_5078,N_5176);
nor U5339 (N_5339,N_5137,N_5064);
nand U5340 (N_5340,N_5024,N_5139);
nand U5341 (N_5341,N_5171,N_5177);
nand U5342 (N_5342,N_5178,N_5034);
nand U5343 (N_5343,N_5007,N_5062);
or U5344 (N_5344,N_5088,N_5135);
nand U5345 (N_5345,N_5129,N_5094);
xnor U5346 (N_5346,N_5117,N_5180);
or U5347 (N_5347,N_5143,N_5040);
or U5348 (N_5348,N_5038,N_5196);
or U5349 (N_5349,N_5022,N_5053);
or U5350 (N_5350,N_5193,N_5189);
xor U5351 (N_5351,N_5001,N_5047);
or U5352 (N_5352,N_5147,N_5054);
xor U5353 (N_5353,N_5115,N_5078);
or U5354 (N_5354,N_5166,N_5168);
nor U5355 (N_5355,N_5004,N_5008);
xor U5356 (N_5356,N_5152,N_5060);
or U5357 (N_5357,N_5019,N_5180);
nand U5358 (N_5358,N_5125,N_5108);
or U5359 (N_5359,N_5144,N_5136);
nand U5360 (N_5360,N_5149,N_5170);
and U5361 (N_5361,N_5112,N_5044);
and U5362 (N_5362,N_5083,N_5144);
and U5363 (N_5363,N_5105,N_5052);
and U5364 (N_5364,N_5069,N_5171);
or U5365 (N_5365,N_5093,N_5000);
nor U5366 (N_5366,N_5058,N_5049);
and U5367 (N_5367,N_5058,N_5067);
and U5368 (N_5368,N_5063,N_5129);
xor U5369 (N_5369,N_5148,N_5181);
nor U5370 (N_5370,N_5057,N_5171);
and U5371 (N_5371,N_5156,N_5014);
or U5372 (N_5372,N_5174,N_5080);
and U5373 (N_5373,N_5095,N_5072);
and U5374 (N_5374,N_5181,N_5103);
xnor U5375 (N_5375,N_5165,N_5041);
nand U5376 (N_5376,N_5057,N_5139);
nor U5377 (N_5377,N_5040,N_5176);
and U5378 (N_5378,N_5102,N_5118);
xnor U5379 (N_5379,N_5103,N_5051);
and U5380 (N_5380,N_5166,N_5013);
and U5381 (N_5381,N_5168,N_5145);
nand U5382 (N_5382,N_5162,N_5013);
nand U5383 (N_5383,N_5033,N_5013);
nand U5384 (N_5384,N_5155,N_5010);
nand U5385 (N_5385,N_5021,N_5075);
and U5386 (N_5386,N_5066,N_5125);
nor U5387 (N_5387,N_5189,N_5107);
nor U5388 (N_5388,N_5047,N_5196);
xnor U5389 (N_5389,N_5074,N_5126);
nor U5390 (N_5390,N_5131,N_5113);
and U5391 (N_5391,N_5050,N_5143);
nor U5392 (N_5392,N_5094,N_5078);
nand U5393 (N_5393,N_5045,N_5157);
nor U5394 (N_5394,N_5129,N_5084);
or U5395 (N_5395,N_5133,N_5152);
nor U5396 (N_5396,N_5055,N_5127);
or U5397 (N_5397,N_5171,N_5108);
nand U5398 (N_5398,N_5137,N_5017);
nor U5399 (N_5399,N_5100,N_5141);
or U5400 (N_5400,N_5384,N_5325);
nand U5401 (N_5401,N_5266,N_5399);
xor U5402 (N_5402,N_5295,N_5315);
and U5403 (N_5403,N_5254,N_5236);
nand U5404 (N_5404,N_5354,N_5210);
nand U5405 (N_5405,N_5257,N_5272);
nand U5406 (N_5406,N_5291,N_5264);
nor U5407 (N_5407,N_5246,N_5312);
nand U5408 (N_5408,N_5263,N_5284);
nand U5409 (N_5409,N_5357,N_5378);
xnor U5410 (N_5410,N_5369,N_5248);
xnor U5411 (N_5411,N_5350,N_5339);
xor U5412 (N_5412,N_5390,N_5323);
nand U5413 (N_5413,N_5244,N_5281);
xor U5414 (N_5414,N_5372,N_5258);
or U5415 (N_5415,N_5207,N_5228);
or U5416 (N_5416,N_5376,N_5287);
or U5417 (N_5417,N_5252,N_5290);
nor U5418 (N_5418,N_5214,N_5371);
nand U5419 (N_5419,N_5269,N_5235);
or U5420 (N_5420,N_5392,N_5338);
or U5421 (N_5421,N_5275,N_5368);
nor U5422 (N_5422,N_5270,N_5309);
or U5423 (N_5423,N_5294,N_5231);
or U5424 (N_5424,N_5268,N_5293);
nand U5425 (N_5425,N_5216,N_5277);
or U5426 (N_5426,N_5343,N_5328);
nand U5427 (N_5427,N_5395,N_5299);
nand U5428 (N_5428,N_5249,N_5342);
and U5429 (N_5429,N_5310,N_5363);
nor U5430 (N_5430,N_5320,N_5226);
xor U5431 (N_5431,N_5380,N_5351);
nand U5432 (N_5432,N_5240,N_5253);
and U5433 (N_5433,N_5217,N_5292);
xor U5434 (N_5434,N_5335,N_5382);
or U5435 (N_5435,N_5209,N_5322);
and U5436 (N_5436,N_5330,N_5324);
nand U5437 (N_5437,N_5267,N_5242);
xor U5438 (N_5438,N_5327,N_5233);
and U5439 (N_5439,N_5208,N_5200);
or U5440 (N_5440,N_5301,N_5358);
nor U5441 (N_5441,N_5204,N_5307);
or U5442 (N_5442,N_5261,N_5308);
xnor U5443 (N_5443,N_5305,N_5362);
nor U5444 (N_5444,N_5365,N_5367);
xnor U5445 (N_5445,N_5388,N_5234);
xor U5446 (N_5446,N_5239,N_5241);
or U5447 (N_5447,N_5394,N_5348);
nand U5448 (N_5448,N_5379,N_5206);
and U5449 (N_5449,N_5302,N_5250);
and U5450 (N_5450,N_5353,N_5326);
nor U5451 (N_5451,N_5319,N_5316);
or U5452 (N_5452,N_5243,N_5260);
and U5453 (N_5453,N_5265,N_5313);
nand U5454 (N_5454,N_5355,N_5289);
and U5455 (N_5455,N_5286,N_5262);
nand U5456 (N_5456,N_5389,N_5336);
and U5457 (N_5457,N_5337,N_5245);
and U5458 (N_5458,N_5237,N_5361);
or U5459 (N_5459,N_5385,N_5224);
and U5460 (N_5460,N_5201,N_5359);
and U5461 (N_5461,N_5238,N_5278);
nand U5462 (N_5462,N_5218,N_5247);
and U5463 (N_5463,N_5282,N_5332);
and U5464 (N_5464,N_5306,N_5356);
xor U5465 (N_5465,N_5251,N_5346);
nand U5466 (N_5466,N_5396,N_5349);
xnor U5467 (N_5467,N_5283,N_5285);
xor U5468 (N_5468,N_5397,N_5321);
or U5469 (N_5469,N_5274,N_5317);
nand U5470 (N_5470,N_5375,N_5331);
nor U5471 (N_5471,N_5215,N_5279);
nand U5472 (N_5472,N_5219,N_5220);
and U5473 (N_5473,N_5203,N_5311);
and U5474 (N_5474,N_5223,N_5222);
nand U5475 (N_5475,N_5373,N_5256);
nand U5476 (N_5476,N_5259,N_5227);
nor U5477 (N_5477,N_5329,N_5374);
and U5478 (N_5478,N_5364,N_5205);
and U5479 (N_5479,N_5334,N_5333);
and U5480 (N_5480,N_5296,N_5213);
and U5481 (N_5481,N_5383,N_5211);
nand U5482 (N_5482,N_5297,N_5347);
and U5483 (N_5483,N_5271,N_5280);
nand U5484 (N_5484,N_5377,N_5314);
and U5485 (N_5485,N_5340,N_5381);
xnor U5486 (N_5486,N_5225,N_5360);
nand U5487 (N_5487,N_5345,N_5255);
nor U5488 (N_5488,N_5386,N_5366);
nor U5489 (N_5489,N_5298,N_5318);
xor U5490 (N_5490,N_5370,N_5273);
xnor U5491 (N_5491,N_5229,N_5391);
xor U5492 (N_5492,N_5232,N_5304);
nor U5493 (N_5493,N_5387,N_5303);
or U5494 (N_5494,N_5300,N_5230);
nand U5495 (N_5495,N_5202,N_5352);
xnor U5496 (N_5496,N_5344,N_5341);
and U5497 (N_5497,N_5393,N_5221);
and U5498 (N_5498,N_5276,N_5212);
or U5499 (N_5499,N_5398,N_5288);
and U5500 (N_5500,N_5221,N_5307);
nand U5501 (N_5501,N_5259,N_5397);
nand U5502 (N_5502,N_5275,N_5327);
xor U5503 (N_5503,N_5298,N_5221);
nand U5504 (N_5504,N_5333,N_5275);
and U5505 (N_5505,N_5224,N_5206);
xor U5506 (N_5506,N_5209,N_5293);
or U5507 (N_5507,N_5268,N_5335);
or U5508 (N_5508,N_5212,N_5243);
nor U5509 (N_5509,N_5344,N_5269);
or U5510 (N_5510,N_5393,N_5385);
or U5511 (N_5511,N_5381,N_5260);
nand U5512 (N_5512,N_5310,N_5317);
xor U5513 (N_5513,N_5267,N_5220);
or U5514 (N_5514,N_5255,N_5372);
nand U5515 (N_5515,N_5322,N_5357);
or U5516 (N_5516,N_5316,N_5286);
nor U5517 (N_5517,N_5282,N_5263);
nor U5518 (N_5518,N_5207,N_5273);
nor U5519 (N_5519,N_5340,N_5397);
xnor U5520 (N_5520,N_5235,N_5347);
nand U5521 (N_5521,N_5392,N_5344);
xnor U5522 (N_5522,N_5376,N_5237);
xor U5523 (N_5523,N_5247,N_5296);
and U5524 (N_5524,N_5216,N_5380);
or U5525 (N_5525,N_5202,N_5259);
nor U5526 (N_5526,N_5340,N_5379);
nand U5527 (N_5527,N_5302,N_5315);
or U5528 (N_5528,N_5283,N_5272);
nor U5529 (N_5529,N_5218,N_5336);
nor U5530 (N_5530,N_5318,N_5281);
or U5531 (N_5531,N_5271,N_5331);
nand U5532 (N_5532,N_5336,N_5237);
and U5533 (N_5533,N_5392,N_5341);
nor U5534 (N_5534,N_5379,N_5391);
nand U5535 (N_5535,N_5213,N_5371);
or U5536 (N_5536,N_5216,N_5353);
nor U5537 (N_5537,N_5201,N_5318);
or U5538 (N_5538,N_5285,N_5346);
xor U5539 (N_5539,N_5378,N_5278);
or U5540 (N_5540,N_5326,N_5364);
xnor U5541 (N_5541,N_5229,N_5317);
or U5542 (N_5542,N_5374,N_5275);
and U5543 (N_5543,N_5248,N_5337);
or U5544 (N_5544,N_5396,N_5201);
xnor U5545 (N_5545,N_5278,N_5361);
nor U5546 (N_5546,N_5376,N_5378);
or U5547 (N_5547,N_5339,N_5287);
nand U5548 (N_5548,N_5316,N_5318);
nor U5549 (N_5549,N_5371,N_5237);
xnor U5550 (N_5550,N_5360,N_5252);
and U5551 (N_5551,N_5215,N_5358);
nor U5552 (N_5552,N_5346,N_5297);
or U5553 (N_5553,N_5362,N_5256);
nor U5554 (N_5554,N_5333,N_5204);
xor U5555 (N_5555,N_5265,N_5220);
or U5556 (N_5556,N_5240,N_5257);
or U5557 (N_5557,N_5278,N_5248);
and U5558 (N_5558,N_5341,N_5245);
and U5559 (N_5559,N_5380,N_5235);
xor U5560 (N_5560,N_5302,N_5387);
and U5561 (N_5561,N_5212,N_5217);
nor U5562 (N_5562,N_5216,N_5315);
and U5563 (N_5563,N_5204,N_5388);
or U5564 (N_5564,N_5399,N_5261);
nand U5565 (N_5565,N_5227,N_5201);
and U5566 (N_5566,N_5303,N_5326);
nand U5567 (N_5567,N_5203,N_5271);
xor U5568 (N_5568,N_5350,N_5271);
nor U5569 (N_5569,N_5351,N_5366);
or U5570 (N_5570,N_5276,N_5308);
nor U5571 (N_5571,N_5323,N_5271);
nand U5572 (N_5572,N_5281,N_5243);
nand U5573 (N_5573,N_5306,N_5311);
xor U5574 (N_5574,N_5302,N_5282);
xor U5575 (N_5575,N_5244,N_5359);
or U5576 (N_5576,N_5305,N_5348);
xor U5577 (N_5577,N_5298,N_5274);
or U5578 (N_5578,N_5365,N_5380);
and U5579 (N_5579,N_5291,N_5205);
xnor U5580 (N_5580,N_5309,N_5228);
xor U5581 (N_5581,N_5280,N_5334);
or U5582 (N_5582,N_5247,N_5252);
or U5583 (N_5583,N_5370,N_5307);
or U5584 (N_5584,N_5338,N_5379);
or U5585 (N_5585,N_5398,N_5324);
nor U5586 (N_5586,N_5371,N_5373);
xor U5587 (N_5587,N_5228,N_5211);
and U5588 (N_5588,N_5304,N_5340);
xor U5589 (N_5589,N_5226,N_5217);
nor U5590 (N_5590,N_5397,N_5367);
nor U5591 (N_5591,N_5320,N_5298);
or U5592 (N_5592,N_5219,N_5228);
or U5593 (N_5593,N_5223,N_5300);
nor U5594 (N_5594,N_5275,N_5270);
xnor U5595 (N_5595,N_5295,N_5317);
nand U5596 (N_5596,N_5364,N_5294);
nand U5597 (N_5597,N_5382,N_5242);
nand U5598 (N_5598,N_5241,N_5385);
nor U5599 (N_5599,N_5218,N_5263);
xor U5600 (N_5600,N_5401,N_5443);
nand U5601 (N_5601,N_5410,N_5546);
nand U5602 (N_5602,N_5432,N_5429);
and U5603 (N_5603,N_5516,N_5562);
nand U5604 (N_5604,N_5490,N_5577);
xnor U5605 (N_5605,N_5555,N_5473);
or U5606 (N_5606,N_5487,N_5439);
nand U5607 (N_5607,N_5413,N_5542);
and U5608 (N_5608,N_5552,N_5531);
xor U5609 (N_5609,N_5587,N_5502);
xnor U5610 (N_5610,N_5509,N_5447);
or U5611 (N_5611,N_5431,N_5582);
nor U5612 (N_5612,N_5591,N_5438);
and U5613 (N_5613,N_5455,N_5525);
or U5614 (N_5614,N_5475,N_5427);
and U5615 (N_5615,N_5574,N_5583);
or U5616 (N_5616,N_5507,N_5521);
xnor U5617 (N_5617,N_5476,N_5530);
xor U5618 (N_5618,N_5573,N_5408);
or U5619 (N_5619,N_5456,N_5533);
xor U5620 (N_5620,N_5417,N_5534);
or U5621 (N_5621,N_5549,N_5596);
and U5622 (N_5622,N_5560,N_5474);
nand U5623 (N_5623,N_5508,N_5592);
nand U5624 (N_5624,N_5481,N_5599);
and U5625 (N_5625,N_5598,N_5457);
xor U5626 (N_5626,N_5437,N_5515);
xor U5627 (N_5627,N_5561,N_5557);
or U5628 (N_5628,N_5519,N_5559);
nor U5629 (N_5629,N_5576,N_5567);
and U5630 (N_5630,N_5543,N_5544);
nand U5631 (N_5631,N_5485,N_5460);
nand U5632 (N_5632,N_5436,N_5482);
and U5633 (N_5633,N_5537,N_5514);
nand U5634 (N_5634,N_5588,N_5421);
nand U5635 (N_5635,N_5424,N_5450);
nand U5636 (N_5636,N_5445,N_5469);
nand U5637 (N_5637,N_5480,N_5483);
nand U5638 (N_5638,N_5412,N_5558);
or U5639 (N_5639,N_5400,N_5496);
xor U5640 (N_5640,N_5597,N_5477);
and U5641 (N_5641,N_5548,N_5492);
or U5642 (N_5642,N_5453,N_5538);
nor U5643 (N_5643,N_5568,N_5532);
nor U5644 (N_5644,N_5451,N_5551);
or U5645 (N_5645,N_5500,N_5566);
and U5646 (N_5646,N_5503,N_5467);
xnor U5647 (N_5647,N_5446,N_5471);
and U5648 (N_5648,N_5565,N_5589);
nand U5649 (N_5649,N_5423,N_5522);
nand U5650 (N_5650,N_5479,N_5563);
nand U5651 (N_5651,N_5428,N_5586);
nand U5652 (N_5652,N_5539,N_5518);
xor U5653 (N_5653,N_5569,N_5405);
or U5654 (N_5654,N_5418,N_5575);
xnor U5655 (N_5655,N_5462,N_5425);
xnor U5656 (N_5656,N_5472,N_5550);
nor U5657 (N_5657,N_5498,N_5488);
nand U5658 (N_5658,N_5415,N_5506);
xnor U5659 (N_5659,N_5512,N_5406);
or U5660 (N_5660,N_5556,N_5536);
nor U5661 (N_5661,N_5404,N_5416);
xnor U5662 (N_5662,N_5435,N_5535);
or U5663 (N_5663,N_5442,N_5564);
and U5664 (N_5664,N_5468,N_5458);
and U5665 (N_5665,N_5547,N_5449);
nand U5666 (N_5666,N_5466,N_5441);
xnor U5667 (N_5667,N_5529,N_5584);
nand U5668 (N_5668,N_5422,N_5486);
and U5669 (N_5669,N_5572,N_5493);
and U5670 (N_5670,N_5461,N_5419);
xor U5671 (N_5671,N_5581,N_5520);
nor U5672 (N_5672,N_5407,N_5528);
and U5673 (N_5673,N_5526,N_5523);
nand U5674 (N_5674,N_5464,N_5517);
xnor U5675 (N_5675,N_5527,N_5570);
nor U5676 (N_5676,N_5585,N_5448);
nand U5677 (N_5677,N_5463,N_5571);
and U5678 (N_5678,N_5540,N_5505);
nand U5679 (N_5679,N_5491,N_5553);
nor U5680 (N_5680,N_5578,N_5426);
nand U5681 (N_5681,N_5590,N_5409);
nand U5682 (N_5682,N_5504,N_5510);
xor U5683 (N_5683,N_5541,N_5454);
nand U5684 (N_5684,N_5595,N_5580);
xor U5685 (N_5685,N_5594,N_5484);
nor U5686 (N_5686,N_5499,N_5495);
or U5687 (N_5687,N_5434,N_5403);
and U5688 (N_5688,N_5402,N_5513);
or U5689 (N_5689,N_5433,N_5497);
and U5690 (N_5690,N_5489,N_5465);
and U5691 (N_5691,N_5414,N_5459);
nor U5692 (N_5692,N_5511,N_5420);
nand U5693 (N_5693,N_5579,N_5545);
or U5694 (N_5694,N_5478,N_5494);
or U5695 (N_5695,N_5524,N_5430);
or U5696 (N_5696,N_5593,N_5554);
nand U5697 (N_5697,N_5444,N_5452);
nand U5698 (N_5698,N_5440,N_5411);
or U5699 (N_5699,N_5470,N_5501);
xor U5700 (N_5700,N_5528,N_5543);
xor U5701 (N_5701,N_5453,N_5416);
or U5702 (N_5702,N_5423,N_5428);
xor U5703 (N_5703,N_5425,N_5514);
and U5704 (N_5704,N_5415,N_5529);
nor U5705 (N_5705,N_5466,N_5572);
nand U5706 (N_5706,N_5548,N_5415);
nand U5707 (N_5707,N_5560,N_5411);
xor U5708 (N_5708,N_5496,N_5444);
and U5709 (N_5709,N_5482,N_5586);
nand U5710 (N_5710,N_5523,N_5483);
or U5711 (N_5711,N_5406,N_5549);
nor U5712 (N_5712,N_5447,N_5590);
nor U5713 (N_5713,N_5422,N_5491);
or U5714 (N_5714,N_5583,N_5597);
xor U5715 (N_5715,N_5443,N_5572);
nand U5716 (N_5716,N_5546,N_5451);
and U5717 (N_5717,N_5546,N_5479);
nand U5718 (N_5718,N_5577,N_5480);
and U5719 (N_5719,N_5406,N_5581);
nor U5720 (N_5720,N_5426,N_5596);
nor U5721 (N_5721,N_5453,N_5400);
and U5722 (N_5722,N_5586,N_5552);
nor U5723 (N_5723,N_5564,N_5428);
xnor U5724 (N_5724,N_5400,N_5558);
nor U5725 (N_5725,N_5587,N_5418);
nor U5726 (N_5726,N_5552,N_5483);
xor U5727 (N_5727,N_5419,N_5487);
xnor U5728 (N_5728,N_5403,N_5551);
or U5729 (N_5729,N_5519,N_5572);
and U5730 (N_5730,N_5435,N_5436);
or U5731 (N_5731,N_5406,N_5515);
nor U5732 (N_5732,N_5457,N_5510);
nand U5733 (N_5733,N_5592,N_5544);
nor U5734 (N_5734,N_5512,N_5521);
and U5735 (N_5735,N_5535,N_5439);
or U5736 (N_5736,N_5484,N_5418);
and U5737 (N_5737,N_5453,N_5585);
nand U5738 (N_5738,N_5519,N_5461);
xor U5739 (N_5739,N_5546,N_5598);
or U5740 (N_5740,N_5479,N_5408);
and U5741 (N_5741,N_5502,N_5415);
nand U5742 (N_5742,N_5591,N_5419);
nand U5743 (N_5743,N_5402,N_5497);
xor U5744 (N_5744,N_5495,N_5528);
nor U5745 (N_5745,N_5554,N_5429);
or U5746 (N_5746,N_5565,N_5571);
xnor U5747 (N_5747,N_5435,N_5415);
or U5748 (N_5748,N_5472,N_5545);
and U5749 (N_5749,N_5489,N_5485);
nor U5750 (N_5750,N_5429,N_5599);
nor U5751 (N_5751,N_5496,N_5405);
or U5752 (N_5752,N_5469,N_5580);
or U5753 (N_5753,N_5584,N_5583);
nand U5754 (N_5754,N_5469,N_5553);
or U5755 (N_5755,N_5410,N_5515);
nand U5756 (N_5756,N_5524,N_5584);
nand U5757 (N_5757,N_5480,N_5405);
and U5758 (N_5758,N_5440,N_5482);
or U5759 (N_5759,N_5562,N_5498);
or U5760 (N_5760,N_5498,N_5547);
nor U5761 (N_5761,N_5568,N_5479);
or U5762 (N_5762,N_5583,N_5598);
and U5763 (N_5763,N_5560,N_5432);
nor U5764 (N_5764,N_5436,N_5596);
nor U5765 (N_5765,N_5562,N_5408);
or U5766 (N_5766,N_5573,N_5437);
or U5767 (N_5767,N_5562,N_5561);
nand U5768 (N_5768,N_5489,N_5581);
and U5769 (N_5769,N_5475,N_5542);
or U5770 (N_5770,N_5423,N_5419);
and U5771 (N_5771,N_5542,N_5527);
nor U5772 (N_5772,N_5464,N_5537);
nand U5773 (N_5773,N_5466,N_5514);
xnor U5774 (N_5774,N_5488,N_5473);
nand U5775 (N_5775,N_5586,N_5547);
or U5776 (N_5776,N_5507,N_5431);
nand U5777 (N_5777,N_5549,N_5551);
nor U5778 (N_5778,N_5414,N_5411);
nand U5779 (N_5779,N_5444,N_5457);
xor U5780 (N_5780,N_5536,N_5458);
nand U5781 (N_5781,N_5561,N_5559);
and U5782 (N_5782,N_5445,N_5467);
nor U5783 (N_5783,N_5455,N_5577);
or U5784 (N_5784,N_5521,N_5479);
and U5785 (N_5785,N_5587,N_5410);
nor U5786 (N_5786,N_5457,N_5451);
and U5787 (N_5787,N_5435,N_5467);
xor U5788 (N_5788,N_5536,N_5533);
and U5789 (N_5789,N_5465,N_5587);
nand U5790 (N_5790,N_5473,N_5553);
nor U5791 (N_5791,N_5509,N_5428);
and U5792 (N_5792,N_5585,N_5497);
or U5793 (N_5793,N_5512,N_5414);
nand U5794 (N_5794,N_5559,N_5494);
xnor U5795 (N_5795,N_5469,N_5491);
nor U5796 (N_5796,N_5418,N_5482);
or U5797 (N_5797,N_5483,N_5528);
xor U5798 (N_5798,N_5511,N_5477);
nand U5799 (N_5799,N_5576,N_5569);
nor U5800 (N_5800,N_5659,N_5716);
nor U5801 (N_5801,N_5627,N_5608);
nor U5802 (N_5802,N_5681,N_5617);
nand U5803 (N_5803,N_5763,N_5682);
or U5804 (N_5804,N_5751,N_5637);
and U5805 (N_5805,N_5770,N_5706);
xnor U5806 (N_5806,N_5692,N_5670);
xor U5807 (N_5807,N_5758,N_5623);
nand U5808 (N_5808,N_5641,N_5720);
xor U5809 (N_5809,N_5785,N_5766);
or U5810 (N_5810,N_5779,N_5619);
xnor U5811 (N_5811,N_5648,N_5772);
xnor U5812 (N_5812,N_5738,N_5740);
nand U5813 (N_5813,N_5684,N_5604);
and U5814 (N_5814,N_5680,N_5700);
or U5815 (N_5815,N_5689,N_5728);
nor U5816 (N_5816,N_5739,N_5612);
xnor U5817 (N_5817,N_5775,N_5661);
and U5818 (N_5818,N_5709,N_5695);
and U5819 (N_5819,N_5794,N_5660);
or U5820 (N_5820,N_5694,N_5731);
nand U5821 (N_5821,N_5727,N_5654);
nand U5822 (N_5822,N_5756,N_5656);
and U5823 (N_5823,N_5683,N_5719);
nor U5824 (N_5824,N_5634,N_5703);
and U5825 (N_5825,N_5721,N_5699);
xnor U5826 (N_5826,N_5747,N_5603);
or U5827 (N_5827,N_5626,N_5616);
nor U5828 (N_5828,N_5601,N_5701);
nor U5829 (N_5829,N_5675,N_5714);
xor U5830 (N_5830,N_5786,N_5618);
or U5831 (N_5831,N_5606,N_5639);
or U5832 (N_5832,N_5657,N_5686);
or U5833 (N_5833,N_5759,N_5705);
nor U5834 (N_5834,N_5600,N_5658);
xor U5835 (N_5835,N_5646,N_5613);
or U5836 (N_5836,N_5737,N_5744);
and U5837 (N_5837,N_5762,N_5712);
nand U5838 (N_5838,N_5733,N_5668);
nand U5839 (N_5839,N_5771,N_5726);
nand U5840 (N_5840,N_5696,N_5783);
or U5841 (N_5841,N_5708,N_5602);
xor U5842 (N_5842,N_5678,N_5761);
nand U5843 (N_5843,N_5677,N_5671);
or U5844 (N_5844,N_5723,N_5715);
and U5845 (N_5845,N_5650,N_5638);
xnor U5846 (N_5846,N_5609,N_5636);
nor U5847 (N_5847,N_5798,N_5605);
nor U5848 (N_5848,N_5745,N_5620);
and U5849 (N_5849,N_5614,N_5791);
nor U5850 (N_5850,N_5769,N_5748);
or U5851 (N_5851,N_5743,N_5615);
nand U5852 (N_5852,N_5711,N_5778);
nand U5853 (N_5853,N_5782,N_5746);
and U5854 (N_5854,N_5665,N_5688);
nand U5855 (N_5855,N_5797,N_5741);
or U5856 (N_5856,N_5799,N_5685);
or U5857 (N_5857,N_5679,N_5653);
nor U5858 (N_5858,N_5645,N_5644);
nor U5859 (N_5859,N_5621,N_5767);
or U5860 (N_5860,N_5787,N_5742);
and U5861 (N_5861,N_5640,N_5629);
nor U5862 (N_5862,N_5749,N_5662);
nand U5863 (N_5863,N_5732,N_5784);
and U5864 (N_5864,N_5667,N_5789);
nor U5865 (N_5865,N_5625,N_5750);
nand U5866 (N_5866,N_5633,N_5611);
nand U5867 (N_5867,N_5718,N_5652);
or U5868 (N_5868,N_5768,N_5704);
nand U5869 (N_5869,N_5729,N_5780);
nor U5870 (N_5870,N_5725,N_5735);
or U5871 (N_5871,N_5776,N_5774);
and U5872 (N_5872,N_5655,N_5690);
and U5873 (N_5873,N_5632,N_5676);
xnor U5874 (N_5874,N_5649,N_5792);
xnor U5875 (N_5875,N_5736,N_5734);
or U5876 (N_5876,N_5691,N_5702);
and U5877 (N_5877,N_5630,N_5607);
nor U5878 (N_5878,N_5672,N_5666);
nand U5879 (N_5879,N_5722,N_5764);
or U5880 (N_5880,N_5624,N_5697);
nor U5881 (N_5881,N_5693,N_5669);
xor U5882 (N_5882,N_5674,N_5796);
nor U5883 (N_5883,N_5647,N_5642);
or U5884 (N_5884,N_5781,N_5631);
or U5885 (N_5885,N_5698,N_5730);
and U5886 (N_5886,N_5710,N_5635);
xnor U5887 (N_5887,N_5717,N_5610);
xor U5888 (N_5888,N_5651,N_5622);
nor U5889 (N_5889,N_5793,N_5724);
xor U5890 (N_5890,N_5753,N_5790);
nor U5891 (N_5891,N_5754,N_5628);
nand U5892 (N_5892,N_5752,N_5755);
nand U5893 (N_5893,N_5713,N_5765);
and U5894 (N_5894,N_5664,N_5687);
nor U5895 (N_5895,N_5795,N_5773);
or U5896 (N_5896,N_5643,N_5707);
nor U5897 (N_5897,N_5760,N_5663);
or U5898 (N_5898,N_5788,N_5777);
nor U5899 (N_5899,N_5673,N_5757);
or U5900 (N_5900,N_5624,N_5646);
xnor U5901 (N_5901,N_5618,N_5735);
xnor U5902 (N_5902,N_5607,N_5629);
nand U5903 (N_5903,N_5784,N_5617);
nand U5904 (N_5904,N_5620,N_5650);
or U5905 (N_5905,N_5704,N_5737);
and U5906 (N_5906,N_5679,N_5678);
nor U5907 (N_5907,N_5730,N_5674);
and U5908 (N_5908,N_5682,N_5627);
or U5909 (N_5909,N_5746,N_5626);
nor U5910 (N_5910,N_5676,N_5772);
xnor U5911 (N_5911,N_5721,N_5628);
and U5912 (N_5912,N_5712,N_5745);
or U5913 (N_5913,N_5785,N_5622);
nor U5914 (N_5914,N_5626,N_5728);
or U5915 (N_5915,N_5662,N_5676);
nand U5916 (N_5916,N_5668,N_5652);
or U5917 (N_5917,N_5706,N_5629);
nor U5918 (N_5918,N_5727,N_5621);
or U5919 (N_5919,N_5758,N_5767);
nand U5920 (N_5920,N_5702,N_5757);
nor U5921 (N_5921,N_5709,N_5784);
and U5922 (N_5922,N_5609,N_5666);
or U5923 (N_5923,N_5747,N_5741);
xnor U5924 (N_5924,N_5782,N_5779);
and U5925 (N_5925,N_5733,N_5790);
nor U5926 (N_5926,N_5606,N_5763);
and U5927 (N_5927,N_5635,N_5722);
nor U5928 (N_5928,N_5661,N_5797);
and U5929 (N_5929,N_5704,N_5722);
or U5930 (N_5930,N_5703,N_5620);
xnor U5931 (N_5931,N_5779,N_5628);
or U5932 (N_5932,N_5651,N_5727);
and U5933 (N_5933,N_5750,N_5783);
xnor U5934 (N_5934,N_5772,N_5777);
nor U5935 (N_5935,N_5701,N_5687);
and U5936 (N_5936,N_5600,N_5784);
nor U5937 (N_5937,N_5685,N_5789);
and U5938 (N_5938,N_5669,N_5638);
or U5939 (N_5939,N_5669,N_5761);
nor U5940 (N_5940,N_5724,N_5618);
and U5941 (N_5941,N_5770,N_5695);
or U5942 (N_5942,N_5612,N_5711);
nor U5943 (N_5943,N_5705,N_5751);
and U5944 (N_5944,N_5774,N_5755);
and U5945 (N_5945,N_5633,N_5647);
nand U5946 (N_5946,N_5682,N_5751);
or U5947 (N_5947,N_5769,N_5692);
xnor U5948 (N_5948,N_5759,N_5668);
and U5949 (N_5949,N_5732,N_5683);
xnor U5950 (N_5950,N_5747,N_5671);
nor U5951 (N_5951,N_5798,N_5755);
or U5952 (N_5952,N_5618,N_5751);
xor U5953 (N_5953,N_5786,N_5708);
nor U5954 (N_5954,N_5750,N_5735);
or U5955 (N_5955,N_5681,N_5647);
or U5956 (N_5956,N_5783,N_5770);
xor U5957 (N_5957,N_5603,N_5767);
or U5958 (N_5958,N_5680,N_5609);
nand U5959 (N_5959,N_5707,N_5644);
and U5960 (N_5960,N_5741,N_5627);
or U5961 (N_5961,N_5672,N_5783);
or U5962 (N_5962,N_5678,N_5625);
or U5963 (N_5963,N_5687,N_5722);
and U5964 (N_5964,N_5719,N_5640);
and U5965 (N_5965,N_5773,N_5673);
and U5966 (N_5966,N_5787,N_5704);
or U5967 (N_5967,N_5724,N_5741);
nand U5968 (N_5968,N_5664,N_5607);
and U5969 (N_5969,N_5680,N_5653);
nand U5970 (N_5970,N_5724,N_5783);
and U5971 (N_5971,N_5797,N_5621);
and U5972 (N_5972,N_5699,N_5719);
xnor U5973 (N_5973,N_5763,N_5691);
nor U5974 (N_5974,N_5644,N_5622);
and U5975 (N_5975,N_5745,N_5704);
nor U5976 (N_5976,N_5652,N_5771);
nand U5977 (N_5977,N_5671,N_5625);
nand U5978 (N_5978,N_5713,N_5767);
xor U5979 (N_5979,N_5742,N_5767);
xor U5980 (N_5980,N_5663,N_5609);
nor U5981 (N_5981,N_5714,N_5684);
xor U5982 (N_5982,N_5731,N_5770);
or U5983 (N_5983,N_5786,N_5766);
xnor U5984 (N_5984,N_5697,N_5684);
xor U5985 (N_5985,N_5767,N_5796);
nand U5986 (N_5986,N_5766,N_5780);
nor U5987 (N_5987,N_5763,N_5761);
or U5988 (N_5988,N_5605,N_5616);
nor U5989 (N_5989,N_5726,N_5622);
nor U5990 (N_5990,N_5683,N_5628);
nor U5991 (N_5991,N_5749,N_5630);
or U5992 (N_5992,N_5610,N_5745);
xnor U5993 (N_5993,N_5728,N_5746);
or U5994 (N_5994,N_5655,N_5738);
and U5995 (N_5995,N_5638,N_5661);
or U5996 (N_5996,N_5668,N_5618);
nor U5997 (N_5997,N_5641,N_5678);
and U5998 (N_5998,N_5714,N_5790);
or U5999 (N_5999,N_5653,N_5677);
xor U6000 (N_6000,N_5898,N_5942);
xnor U6001 (N_6001,N_5863,N_5912);
and U6002 (N_6002,N_5804,N_5848);
and U6003 (N_6003,N_5993,N_5864);
and U6004 (N_6004,N_5895,N_5814);
and U6005 (N_6005,N_5940,N_5973);
xnor U6006 (N_6006,N_5997,N_5875);
xor U6007 (N_6007,N_5914,N_5954);
nor U6008 (N_6008,N_5944,N_5913);
nor U6009 (N_6009,N_5858,N_5813);
nand U6010 (N_6010,N_5900,N_5926);
or U6011 (N_6011,N_5809,N_5978);
or U6012 (N_6012,N_5883,N_5932);
nor U6013 (N_6013,N_5995,N_5905);
xnor U6014 (N_6014,N_5921,N_5824);
and U6015 (N_6015,N_5972,N_5806);
and U6016 (N_6016,N_5881,N_5808);
xor U6017 (N_6017,N_5908,N_5843);
nand U6018 (N_6018,N_5839,N_5985);
nor U6019 (N_6019,N_5825,N_5867);
nor U6020 (N_6020,N_5889,N_5817);
and U6021 (N_6021,N_5974,N_5929);
nand U6022 (N_6022,N_5963,N_5847);
nor U6023 (N_6023,N_5807,N_5830);
or U6024 (N_6024,N_5955,N_5994);
and U6025 (N_6025,N_5862,N_5966);
xor U6026 (N_6026,N_5934,N_5840);
xnor U6027 (N_6027,N_5888,N_5968);
xnor U6028 (N_6028,N_5831,N_5918);
xor U6029 (N_6029,N_5854,N_5896);
and U6030 (N_6030,N_5820,N_5981);
nor U6031 (N_6031,N_5937,N_5811);
and U6032 (N_6032,N_5819,N_5826);
or U6033 (N_6033,N_5930,N_5838);
nand U6034 (N_6034,N_5959,N_5936);
nor U6035 (N_6035,N_5935,N_5980);
nand U6036 (N_6036,N_5903,N_5844);
xor U6037 (N_6037,N_5951,N_5953);
nor U6038 (N_6038,N_5938,N_5851);
or U6039 (N_6039,N_5922,N_5902);
nor U6040 (N_6040,N_5871,N_5884);
xor U6041 (N_6041,N_5964,N_5945);
nor U6042 (N_6042,N_5892,N_5958);
nand U6043 (N_6043,N_5880,N_5977);
or U6044 (N_6044,N_5801,N_5841);
and U6045 (N_6045,N_5991,N_5832);
nand U6046 (N_6046,N_5885,N_5961);
or U6047 (N_6047,N_5872,N_5927);
nor U6048 (N_6048,N_5860,N_5986);
xor U6049 (N_6049,N_5984,N_5933);
xor U6050 (N_6050,N_5897,N_5982);
xnor U6051 (N_6051,N_5866,N_5906);
nand U6052 (N_6052,N_5989,N_5803);
nand U6053 (N_6053,N_5917,N_5907);
and U6054 (N_6054,N_5886,N_5810);
nor U6055 (N_6055,N_5971,N_5891);
xor U6056 (N_6056,N_5878,N_5996);
or U6057 (N_6057,N_5845,N_5800);
xnor U6058 (N_6058,N_5822,N_5846);
or U6059 (N_6059,N_5920,N_5915);
xnor U6060 (N_6060,N_5879,N_5979);
or U6061 (N_6061,N_5818,N_5960);
or U6062 (N_6062,N_5957,N_5823);
xnor U6063 (N_6063,N_5952,N_5910);
nor U6064 (N_6064,N_5970,N_5956);
xor U6065 (N_6065,N_5893,N_5887);
nand U6066 (N_6066,N_5924,N_5849);
nand U6067 (N_6067,N_5870,N_5969);
nand U6068 (N_6068,N_5901,N_5948);
nor U6069 (N_6069,N_5909,N_5865);
or U6070 (N_6070,N_5859,N_5877);
nor U6071 (N_6071,N_5941,N_5850);
and U6072 (N_6072,N_5923,N_5853);
and U6073 (N_6073,N_5873,N_5829);
nand U6074 (N_6074,N_5836,N_5983);
nand U6075 (N_6075,N_5827,N_5852);
nor U6076 (N_6076,N_5999,N_5987);
nor U6077 (N_6077,N_5868,N_5855);
or U6078 (N_6078,N_5861,N_5965);
nand U6079 (N_6079,N_5899,N_5894);
or U6080 (N_6080,N_5812,N_5815);
nor U6081 (N_6081,N_5874,N_5856);
xor U6082 (N_6082,N_5837,N_5949);
or U6083 (N_6083,N_5931,N_5992);
or U6084 (N_6084,N_5882,N_5835);
nand U6085 (N_6085,N_5833,N_5842);
or U6086 (N_6086,N_5890,N_5919);
or U6087 (N_6087,N_5925,N_5876);
nand U6088 (N_6088,N_5947,N_5988);
nand U6089 (N_6089,N_5975,N_5939);
nor U6090 (N_6090,N_5916,N_5821);
and U6091 (N_6091,N_5857,N_5998);
nand U6092 (N_6092,N_5911,N_5834);
nor U6093 (N_6093,N_5828,N_5990);
and U6094 (N_6094,N_5869,N_5928);
nor U6095 (N_6095,N_5805,N_5802);
nor U6096 (N_6096,N_5967,N_5816);
or U6097 (N_6097,N_5946,N_5943);
nor U6098 (N_6098,N_5904,N_5976);
nand U6099 (N_6099,N_5962,N_5950);
nor U6100 (N_6100,N_5980,N_5907);
and U6101 (N_6101,N_5978,N_5897);
xnor U6102 (N_6102,N_5868,N_5928);
and U6103 (N_6103,N_5960,N_5997);
nand U6104 (N_6104,N_5920,N_5818);
xnor U6105 (N_6105,N_5947,N_5840);
and U6106 (N_6106,N_5856,N_5910);
nor U6107 (N_6107,N_5947,N_5982);
nor U6108 (N_6108,N_5894,N_5871);
and U6109 (N_6109,N_5998,N_5973);
nand U6110 (N_6110,N_5882,N_5912);
and U6111 (N_6111,N_5872,N_5810);
nand U6112 (N_6112,N_5992,N_5970);
nand U6113 (N_6113,N_5812,N_5854);
and U6114 (N_6114,N_5959,N_5916);
nor U6115 (N_6115,N_5840,N_5872);
or U6116 (N_6116,N_5835,N_5904);
or U6117 (N_6117,N_5851,N_5926);
nand U6118 (N_6118,N_5955,N_5802);
and U6119 (N_6119,N_5996,N_5927);
and U6120 (N_6120,N_5804,N_5944);
nand U6121 (N_6121,N_5802,N_5900);
nor U6122 (N_6122,N_5931,N_5954);
nor U6123 (N_6123,N_5924,N_5869);
nand U6124 (N_6124,N_5963,N_5935);
nor U6125 (N_6125,N_5997,N_5859);
nor U6126 (N_6126,N_5941,N_5803);
nand U6127 (N_6127,N_5956,N_5911);
and U6128 (N_6128,N_5960,N_5840);
nand U6129 (N_6129,N_5927,N_5968);
or U6130 (N_6130,N_5943,N_5853);
and U6131 (N_6131,N_5831,N_5833);
nor U6132 (N_6132,N_5843,N_5808);
nor U6133 (N_6133,N_5889,N_5865);
or U6134 (N_6134,N_5978,N_5965);
xor U6135 (N_6135,N_5803,N_5837);
nor U6136 (N_6136,N_5929,N_5836);
xnor U6137 (N_6137,N_5857,N_5879);
or U6138 (N_6138,N_5977,N_5889);
or U6139 (N_6139,N_5904,N_5964);
nand U6140 (N_6140,N_5925,N_5945);
and U6141 (N_6141,N_5841,N_5958);
or U6142 (N_6142,N_5868,N_5965);
and U6143 (N_6143,N_5892,N_5906);
or U6144 (N_6144,N_5900,N_5941);
nand U6145 (N_6145,N_5914,N_5844);
nand U6146 (N_6146,N_5927,N_5971);
and U6147 (N_6147,N_5844,N_5819);
xor U6148 (N_6148,N_5848,N_5984);
and U6149 (N_6149,N_5906,N_5808);
xor U6150 (N_6150,N_5916,N_5879);
xnor U6151 (N_6151,N_5933,N_5887);
or U6152 (N_6152,N_5895,N_5958);
and U6153 (N_6153,N_5837,N_5825);
nand U6154 (N_6154,N_5961,N_5994);
or U6155 (N_6155,N_5836,N_5883);
nand U6156 (N_6156,N_5985,N_5829);
nor U6157 (N_6157,N_5831,N_5972);
and U6158 (N_6158,N_5997,N_5889);
or U6159 (N_6159,N_5864,N_5880);
and U6160 (N_6160,N_5925,N_5914);
nand U6161 (N_6161,N_5802,N_5819);
nand U6162 (N_6162,N_5930,N_5877);
nor U6163 (N_6163,N_5946,N_5935);
or U6164 (N_6164,N_5833,N_5996);
nor U6165 (N_6165,N_5908,N_5956);
xor U6166 (N_6166,N_5960,N_5925);
nor U6167 (N_6167,N_5843,N_5895);
or U6168 (N_6168,N_5806,N_5885);
and U6169 (N_6169,N_5951,N_5815);
nand U6170 (N_6170,N_5933,N_5821);
and U6171 (N_6171,N_5824,N_5967);
xnor U6172 (N_6172,N_5897,N_5915);
or U6173 (N_6173,N_5952,N_5802);
and U6174 (N_6174,N_5842,N_5959);
or U6175 (N_6175,N_5851,N_5866);
xnor U6176 (N_6176,N_5845,N_5819);
nand U6177 (N_6177,N_5868,N_5809);
or U6178 (N_6178,N_5946,N_5843);
xnor U6179 (N_6179,N_5891,N_5962);
and U6180 (N_6180,N_5811,N_5876);
xor U6181 (N_6181,N_5834,N_5954);
nand U6182 (N_6182,N_5866,N_5912);
nand U6183 (N_6183,N_5962,N_5928);
xnor U6184 (N_6184,N_5945,N_5882);
and U6185 (N_6185,N_5916,N_5880);
xnor U6186 (N_6186,N_5942,N_5856);
nand U6187 (N_6187,N_5920,N_5804);
nand U6188 (N_6188,N_5870,N_5996);
and U6189 (N_6189,N_5935,N_5827);
nand U6190 (N_6190,N_5805,N_5960);
and U6191 (N_6191,N_5824,N_5841);
xnor U6192 (N_6192,N_5914,N_5881);
nand U6193 (N_6193,N_5973,N_5870);
nand U6194 (N_6194,N_5821,N_5863);
nor U6195 (N_6195,N_5912,N_5800);
xnor U6196 (N_6196,N_5848,N_5947);
nor U6197 (N_6197,N_5874,N_5819);
or U6198 (N_6198,N_5864,N_5838);
xor U6199 (N_6199,N_5958,N_5936);
and U6200 (N_6200,N_6166,N_6187);
and U6201 (N_6201,N_6040,N_6115);
nor U6202 (N_6202,N_6043,N_6002);
xnor U6203 (N_6203,N_6135,N_6191);
nand U6204 (N_6204,N_6136,N_6186);
xnor U6205 (N_6205,N_6011,N_6033);
nand U6206 (N_6206,N_6119,N_6104);
or U6207 (N_6207,N_6038,N_6133);
nand U6208 (N_6208,N_6087,N_6060);
or U6209 (N_6209,N_6162,N_6017);
nor U6210 (N_6210,N_6086,N_6059);
and U6211 (N_6211,N_6056,N_6070);
nand U6212 (N_6212,N_6029,N_6013);
nand U6213 (N_6213,N_6152,N_6094);
nor U6214 (N_6214,N_6124,N_6081);
nor U6215 (N_6215,N_6164,N_6092);
or U6216 (N_6216,N_6130,N_6089);
nor U6217 (N_6217,N_6108,N_6053);
nor U6218 (N_6218,N_6116,N_6018);
or U6219 (N_6219,N_6198,N_6068);
and U6220 (N_6220,N_6069,N_6083);
and U6221 (N_6221,N_6167,N_6034);
and U6222 (N_6222,N_6003,N_6022);
nor U6223 (N_6223,N_6126,N_6147);
nand U6224 (N_6224,N_6076,N_6051);
xor U6225 (N_6225,N_6155,N_6122);
nor U6226 (N_6226,N_6182,N_6146);
and U6227 (N_6227,N_6137,N_6010);
and U6228 (N_6228,N_6149,N_6097);
and U6229 (N_6229,N_6020,N_6131);
nand U6230 (N_6230,N_6036,N_6111);
xnor U6231 (N_6231,N_6161,N_6079);
xnor U6232 (N_6232,N_6028,N_6153);
xnor U6233 (N_6233,N_6125,N_6039);
and U6234 (N_6234,N_6192,N_6026);
nor U6235 (N_6235,N_6156,N_6091);
or U6236 (N_6236,N_6165,N_6190);
and U6237 (N_6237,N_6110,N_6129);
xor U6238 (N_6238,N_6168,N_6073);
nor U6239 (N_6239,N_6054,N_6169);
or U6240 (N_6240,N_6012,N_6075);
or U6241 (N_6241,N_6114,N_6151);
and U6242 (N_6242,N_6145,N_6025);
nand U6243 (N_6243,N_6170,N_6046);
or U6244 (N_6244,N_6096,N_6195);
or U6245 (N_6245,N_6100,N_6184);
nor U6246 (N_6246,N_6197,N_6158);
xor U6247 (N_6247,N_6140,N_6128);
nor U6248 (N_6248,N_6024,N_6148);
xor U6249 (N_6249,N_6138,N_6107);
or U6250 (N_6250,N_6078,N_6178);
or U6251 (N_6251,N_6080,N_6142);
and U6252 (N_6252,N_6014,N_6095);
nand U6253 (N_6253,N_6172,N_6090);
nand U6254 (N_6254,N_6199,N_6143);
nand U6255 (N_6255,N_6045,N_6005);
nand U6256 (N_6256,N_6176,N_6181);
or U6257 (N_6257,N_6121,N_6102);
or U6258 (N_6258,N_6196,N_6193);
nor U6259 (N_6259,N_6016,N_6144);
and U6260 (N_6260,N_6042,N_6007);
and U6261 (N_6261,N_6000,N_6027);
nand U6262 (N_6262,N_6037,N_6157);
nor U6263 (N_6263,N_6077,N_6117);
nand U6264 (N_6264,N_6174,N_6139);
or U6265 (N_6265,N_6113,N_6171);
and U6266 (N_6266,N_6004,N_6085);
xnor U6267 (N_6267,N_6071,N_6023);
xor U6268 (N_6268,N_6030,N_6120);
or U6269 (N_6269,N_6185,N_6031);
and U6270 (N_6270,N_6105,N_6065);
and U6271 (N_6271,N_6052,N_6015);
nor U6272 (N_6272,N_6032,N_6189);
xnor U6273 (N_6273,N_6106,N_6066);
or U6274 (N_6274,N_6163,N_6021);
and U6275 (N_6275,N_6188,N_6072);
and U6276 (N_6276,N_6099,N_6063);
and U6277 (N_6277,N_6062,N_6009);
nand U6278 (N_6278,N_6055,N_6084);
nor U6279 (N_6279,N_6118,N_6061);
nand U6280 (N_6280,N_6008,N_6001);
nand U6281 (N_6281,N_6093,N_6127);
nand U6282 (N_6282,N_6074,N_6047);
xnor U6283 (N_6283,N_6194,N_6035);
nand U6284 (N_6284,N_6183,N_6160);
and U6285 (N_6285,N_6082,N_6134);
nor U6286 (N_6286,N_6050,N_6150);
nand U6287 (N_6287,N_6123,N_6044);
or U6288 (N_6288,N_6019,N_6132);
nand U6289 (N_6289,N_6101,N_6057);
and U6290 (N_6290,N_6159,N_6049);
and U6291 (N_6291,N_6098,N_6006);
xnor U6292 (N_6292,N_6180,N_6141);
nor U6293 (N_6293,N_6177,N_6154);
xor U6294 (N_6294,N_6041,N_6058);
and U6295 (N_6295,N_6103,N_6179);
and U6296 (N_6296,N_6064,N_6175);
nor U6297 (N_6297,N_6088,N_6109);
and U6298 (N_6298,N_6067,N_6112);
or U6299 (N_6299,N_6173,N_6048);
nand U6300 (N_6300,N_6166,N_6155);
nor U6301 (N_6301,N_6009,N_6095);
xor U6302 (N_6302,N_6050,N_6134);
nor U6303 (N_6303,N_6114,N_6015);
xor U6304 (N_6304,N_6157,N_6072);
or U6305 (N_6305,N_6121,N_6189);
or U6306 (N_6306,N_6081,N_6156);
nand U6307 (N_6307,N_6054,N_6075);
and U6308 (N_6308,N_6026,N_6097);
nor U6309 (N_6309,N_6011,N_6078);
or U6310 (N_6310,N_6149,N_6152);
and U6311 (N_6311,N_6070,N_6101);
nor U6312 (N_6312,N_6166,N_6025);
nor U6313 (N_6313,N_6151,N_6194);
nand U6314 (N_6314,N_6022,N_6149);
xnor U6315 (N_6315,N_6075,N_6071);
nand U6316 (N_6316,N_6090,N_6049);
nand U6317 (N_6317,N_6160,N_6088);
nand U6318 (N_6318,N_6048,N_6019);
and U6319 (N_6319,N_6030,N_6051);
and U6320 (N_6320,N_6039,N_6175);
nand U6321 (N_6321,N_6138,N_6140);
nand U6322 (N_6322,N_6131,N_6120);
xnor U6323 (N_6323,N_6197,N_6156);
or U6324 (N_6324,N_6165,N_6134);
nor U6325 (N_6325,N_6115,N_6078);
and U6326 (N_6326,N_6009,N_6022);
nor U6327 (N_6327,N_6149,N_6120);
nand U6328 (N_6328,N_6092,N_6126);
xnor U6329 (N_6329,N_6177,N_6117);
or U6330 (N_6330,N_6014,N_6109);
xor U6331 (N_6331,N_6048,N_6168);
nand U6332 (N_6332,N_6131,N_6112);
nor U6333 (N_6333,N_6105,N_6033);
and U6334 (N_6334,N_6054,N_6188);
and U6335 (N_6335,N_6187,N_6037);
nor U6336 (N_6336,N_6054,N_6180);
xor U6337 (N_6337,N_6142,N_6131);
nand U6338 (N_6338,N_6046,N_6058);
xnor U6339 (N_6339,N_6047,N_6054);
and U6340 (N_6340,N_6164,N_6119);
nor U6341 (N_6341,N_6084,N_6178);
xor U6342 (N_6342,N_6190,N_6121);
and U6343 (N_6343,N_6150,N_6060);
xnor U6344 (N_6344,N_6030,N_6053);
and U6345 (N_6345,N_6037,N_6008);
and U6346 (N_6346,N_6015,N_6023);
or U6347 (N_6347,N_6093,N_6005);
xnor U6348 (N_6348,N_6029,N_6076);
and U6349 (N_6349,N_6011,N_6039);
or U6350 (N_6350,N_6119,N_6142);
xor U6351 (N_6351,N_6128,N_6000);
nor U6352 (N_6352,N_6040,N_6181);
or U6353 (N_6353,N_6171,N_6050);
nand U6354 (N_6354,N_6140,N_6079);
nor U6355 (N_6355,N_6039,N_6032);
and U6356 (N_6356,N_6195,N_6128);
or U6357 (N_6357,N_6062,N_6027);
and U6358 (N_6358,N_6149,N_6131);
and U6359 (N_6359,N_6059,N_6064);
xor U6360 (N_6360,N_6008,N_6085);
nor U6361 (N_6361,N_6142,N_6039);
xnor U6362 (N_6362,N_6105,N_6120);
nor U6363 (N_6363,N_6023,N_6073);
or U6364 (N_6364,N_6089,N_6104);
nor U6365 (N_6365,N_6055,N_6110);
nand U6366 (N_6366,N_6018,N_6170);
nor U6367 (N_6367,N_6139,N_6070);
nor U6368 (N_6368,N_6165,N_6183);
and U6369 (N_6369,N_6042,N_6157);
nand U6370 (N_6370,N_6176,N_6036);
or U6371 (N_6371,N_6004,N_6135);
xor U6372 (N_6372,N_6127,N_6117);
nor U6373 (N_6373,N_6096,N_6010);
nor U6374 (N_6374,N_6052,N_6027);
or U6375 (N_6375,N_6093,N_6054);
and U6376 (N_6376,N_6108,N_6158);
and U6377 (N_6377,N_6179,N_6053);
nor U6378 (N_6378,N_6060,N_6077);
and U6379 (N_6379,N_6101,N_6123);
or U6380 (N_6380,N_6136,N_6150);
or U6381 (N_6381,N_6123,N_6140);
or U6382 (N_6382,N_6055,N_6118);
nand U6383 (N_6383,N_6055,N_6150);
or U6384 (N_6384,N_6154,N_6150);
or U6385 (N_6385,N_6032,N_6199);
and U6386 (N_6386,N_6162,N_6100);
and U6387 (N_6387,N_6107,N_6180);
nor U6388 (N_6388,N_6178,N_6039);
nand U6389 (N_6389,N_6085,N_6104);
and U6390 (N_6390,N_6013,N_6028);
nand U6391 (N_6391,N_6183,N_6019);
nor U6392 (N_6392,N_6134,N_6087);
nor U6393 (N_6393,N_6173,N_6121);
xor U6394 (N_6394,N_6153,N_6106);
xnor U6395 (N_6395,N_6164,N_6044);
nand U6396 (N_6396,N_6124,N_6171);
and U6397 (N_6397,N_6119,N_6191);
xnor U6398 (N_6398,N_6068,N_6176);
nor U6399 (N_6399,N_6178,N_6091);
or U6400 (N_6400,N_6398,N_6296);
xnor U6401 (N_6401,N_6231,N_6395);
and U6402 (N_6402,N_6262,N_6328);
or U6403 (N_6403,N_6223,N_6325);
or U6404 (N_6404,N_6373,N_6378);
or U6405 (N_6405,N_6317,N_6265);
nor U6406 (N_6406,N_6238,N_6207);
xnor U6407 (N_6407,N_6200,N_6274);
xor U6408 (N_6408,N_6316,N_6287);
nand U6409 (N_6409,N_6269,N_6235);
and U6410 (N_6410,N_6210,N_6213);
nand U6411 (N_6411,N_6283,N_6326);
or U6412 (N_6412,N_6344,N_6361);
nor U6413 (N_6413,N_6351,N_6365);
nand U6414 (N_6414,N_6346,N_6248);
xor U6415 (N_6415,N_6285,N_6290);
nand U6416 (N_6416,N_6242,N_6389);
or U6417 (N_6417,N_6363,N_6321);
nand U6418 (N_6418,N_6368,N_6237);
xor U6419 (N_6419,N_6301,N_6353);
and U6420 (N_6420,N_6201,N_6270);
xor U6421 (N_6421,N_6203,N_6260);
nor U6422 (N_6422,N_6211,N_6244);
xor U6423 (N_6423,N_6374,N_6202);
nor U6424 (N_6424,N_6228,N_6349);
nor U6425 (N_6425,N_6319,N_6264);
xor U6426 (N_6426,N_6272,N_6247);
or U6427 (N_6427,N_6367,N_6208);
and U6428 (N_6428,N_6281,N_6329);
xor U6429 (N_6429,N_6204,N_6261);
nor U6430 (N_6430,N_6257,N_6371);
nand U6431 (N_6431,N_6256,N_6294);
nand U6432 (N_6432,N_6245,N_6226);
and U6433 (N_6433,N_6302,N_6229);
nand U6434 (N_6434,N_6288,N_6217);
and U6435 (N_6435,N_6286,N_6356);
xnor U6436 (N_6436,N_6307,N_6292);
and U6437 (N_6437,N_6393,N_6318);
xnor U6438 (N_6438,N_6384,N_6216);
and U6439 (N_6439,N_6369,N_6340);
nor U6440 (N_6440,N_6387,N_6249);
xnor U6441 (N_6441,N_6327,N_6336);
xor U6442 (N_6442,N_6370,N_6337);
or U6443 (N_6443,N_6352,N_6215);
nand U6444 (N_6444,N_6320,N_6372);
nor U6445 (N_6445,N_6253,N_6315);
xor U6446 (N_6446,N_6345,N_6366);
and U6447 (N_6447,N_6221,N_6391);
and U6448 (N_6448,N_6394,N_6334);
or U6449 (N_6449,N_6205,N_6392);
xor U6450 (N_6450,N_6343,N_6295);
or U6451 (N_6451,N_6241,N_6278);
nand U6452 (N_6452,N_6390,N_6252);
xor U6453 (N_6453,N_6230,N_6354);
nand U6454 (N_6454,N_6255,N_6324);
and U6455 (N_6455,N_6279,N_6305);
or U6456 (N_6456,N_6299,N_6224);
and U6457 (N_6457,N_6225,N_6322);
or U6458 (N_6458,N_6375,N_6382);
or U6459 (N_6459,N_6251,N_6323);
or U6460 (N_6460,N_6234,N_6341);
and U6461 (N_6461,N_6330,N_6209);
and U6462 (N_6462,N_6271,N_6218);
nor U6463 (N_6463,N_6239,N_6300);
nor U6464 (N_6464,N_6268,N_6227);
and U6465 (N_6465,N_6362,N_6332);
or U6466 (N_6466,N_6219,N_6246);
and U6467 (N_6467,N_6383,N_6212);
nor U6468 (N_6468,N_6308,N_6385);
nor U6469 (N_6469,N_6254,N_6380);
or U6470 (N_6470,N_6309,N_6357);
and U6471 (N_6471,N_6377,N_6291);
or U6472 (N_6472,N_6355,N_6376);
nand U6473 (N_6473,N_6303,N_6250);
and U6474 (N_6474,N_6282,N_6335);
nor U6475 (N_6475,N_6386,N_6236);
xnor U6476 (N_6476,N_6306,N_6333);
or U6477 (N_6477,N_6273,N_6277);
and U6478 (N_6478,N_6396,N_6284);
xor U6479 (N_6479,N_6275,N_6314);
xnor U6480 (N_6480,N_6360,N_6240);
nor U6481 (N_6481,N_6267,N_6379);
nand U6482 (N_6482,N_6259,N_6280);
nor U6483 (N_6483,N_6293,N_6331);
xor U6484 (N_6484,N_6298,N_6347);
and U6485 (N_6485,N_6342,N_6214);
xor U6486 (N_6486,N_6358,N_6388);
nand U6487 (N_6487,N_6266,N_6350);
xor U6488 (N_6488,N_6381,N_6289);
or U6489 (N_6489,N_6263,N_6258);
or U6490 (N_6490,N_6338,N_6364);
nand U6491 (N_6491,N_6304,N_6222);
nor U6492 (N_6492,N_6359,N_6232);
nand U6493 (N_6493,N_6206,N_6348);
xnor U6494 (N_6494,N_6313,N_6310);
xnor U6495 (N_6495,N_6397,N_6243);
or U6496 (N_6496,N_6276,N_6311);
and U6497 (N_6497,N_6339,N_6220);
nor U6498 (N_6498,N_6297,N_6399);
xnor U6499 (N_6499,N_6233,N_6312);
nor U6500 (N_6500,N_6354,N_6328);
nor U6501 (N_6501,N_6347,N_6393);
xor U6502 (N_6502,N_6202,N_6220);
nand U6503 (N_6503,N_6364,N_6227);
or U6504 (N_6504,N_6282,N_6236);
or U6505 (N_6505,N_6206,N_6284);
nand U6506 (N_6506,N_6374,N_6251);
xor U6507 (N_6507,N_6251,N_6218);
or U6508 (N_6508,N_6259,N_6313);
or U6509 (N_6509,N_6218,N_6219);
and U6510 (N_6510,N_6349,N_6385);
or U6511 (N_6511,N_6320,N_6223);
or U6512 (N_6512,N_6298,N_6378);
and U6513 (N_6513,N_6242,N_6368);
or U6514 (N_6514,N_6383,N_6239);
xor U6515 (N_6515,N_6313,N_6321);
or U6516 (N_6516,N_6273,N_6315);
and U6517 (N_6517,N_6237,N_6217);
nor U6518 (N_6518,N_6225,N_6375);
and U6519 (N_6519,N_6219,N_6354);
or U6520 (N_6520,N_6380,N_6225);
and U6521 (N_6521,N_6333,N_6216);
or U6522 (N_6522,N_6370,N_6377);
nand U6523 (N_6523,N_6366,N_6222);
and U6524 (N_6524,N_6293,N_6330);
xor U6525 (N_6525,N_6283,N_6353);
nand U6526 (N_6526,N_6297,N_6222);
and U6527 (N_6527,N_6367,N_6319);
xor U6528 (N_6528,N_6351,N_6350);
or U6529 (N_6529,N_6291,N_6391);
nor U6530 (N_6530,N_6372,N_6362);
xnor U6531 (N_6531,N_6365,N_6247);
nor U6532 (N_6532,N_6269,N_6266);
xnor U6533 (N_6533,N_6343,N_6373);
xnor U6534 (N_6534,N_6211,N_6258);
nor U6535 (N_6535,N_6353,N_6357);
xor U6536 (N_6536,N_6345,N_6374);
nor U6537 (N_6537,N_6354,N_6318);
or U6538 (N_6538,N_6300,N_6245);
or U6539 (N_6539,N_6285,N_6376);
nand U6540 (N_6540,N_6228,N_6210);
and U6541 (N_6541,N_6335,N_6361);
and U6542 (N_6542,N_6355,N_6253);
and U6543 (N_6543,N_6263,N_6383);
and U6544 (N_6544,N_6327,N_6369);
xnor U6545 (N_6545,N_6276,N_6209);
or U6546 (N_6546,N_6364,N_6279);
nor U6547 (N_6547,N_6330,N_6376);
nand U6548 (N_6548,N_6365,N_6385);
nor U6549 (N_6549,N_6313,N_6261);
nor U6550 (N_6550,N_6278,N_6303);
nand U6551 (N_6551,N_6272,N_6206);
xor U6552 (N_6552,N_6376,N_6290);
nand U6553 (N_6553,N_6311,N_6205);
or U6554 (N_6554,N_6242,N_6238);
nor U6555 (N_6555,N_6281,N_6394);
and U6556 (N_6556,N_6255,N_6367);
nor U6557 (N_6557,N_6244,N_6242);
nand U6558 (N_6558,N_6378,N_6344);
or U6559 (N_6559,N_6242,N_6366);
nand U6560 (N_6560,N_6222,N_6301);
nor U6561 (N_6561,N_6358,N_6349);
nor U6562 (N_6562,N_6277,N_6222);
nor U6563 (N_6563,N_6310,N_6355);
nand U6564 (N_6564,N_6338,N_6341);
nor U6565 (N_6565,N_6351,N_6282);
and U6566 (N_6566,N_6251,N_6373);
or U6567 (N_6567,N_6334,N_6318);
xnor U6568 (N_6568,N_6370,N_6381);
nor U6569 (N_6569,N_6316,N_6247);
and U6570 (N_6570,N_6334,N_6357);
nand U6571 (N_6571,N_6295,N_6333);
xor U6572 (N_6572,N_6351,N_6356);
xnor U6573 (N_6573,N_6239,N_6278);
and U6574 (N_6574,N_6260,N_6216);
xnor U6575 (N_6575,N_6332,N_6276);
and U6576 (N_6576,N_6340,N_6234);
nand U6577 (N_6577,N_6204,N_6378);
nand U6578 (N_6578,N_6316,N_6358);
or U6579 (N_6579,N_6289,N_6201);
or U6580 (N_6580,N_6233,N_6295);
nand U6581 (N_6581,N_6279,N_6365);
nand U6582 (N_6582,N_6255,N_6248);
and U6583 (N_6583,N_6313,N_6262);
nor U6584 (N_6584,N_6393,N_6322);
and U6585 (N_6585,N_6224,N_6323);
xor U6586 (N_6586,N_6328,N_6360);
or U6587 (N_6587,N_6219,N_6228);
nand U6588 (N_6588,N_6265,N_6333);
and U6589 (N_6589,N_6256,N_6358);
xnor U6590 (N_6590,N_6234,N_6256);
nand U6591 (N_6591,N_6317,N_6389);
or U6592 (N_6592,N_6274,N_6388);
nand U6593 (N_6593,N_6244,N_6267);
or U6594 (N_6594,N_6383,N_6331);
nand U6595 (N_6595,N_6361,N_6237);
nand U6596 (N_6596,N_6339,N_6279);
and U6597 (N_6597,N_6235,N_6214);
nand U6598 (N_6598,N_6336,N_6335);
nand U6599 (N_6599,N_6351,N_6399);
xnor U6600 (N_6600,N_6579,N_6432);
and U6601 (N_6601,N_6430,N_6511);
nand U6602 (N_6602,N_6505,N_6585);
xnor U6603 (N_6603,N_6552,N_6431);
and U6604 (N_6604,N_6523,N_6529);
xnor U6605 (N_6605,N_6566,N_6416);
xnor U6606 (N_6606,N_6571,N_6447);
nor U6607 (N_6607,N_6503,N_6521);
xnor U6608 (N_6608,N_6551,N_6561);
and U6609 (N_6609,N_6478,N_6509);
or U6610 (N_6610,N_6563,N_6576);
nand U6611 (N_6611,N_6401,N_6567);
xor U6612 (N_6612,N_6510,N_6404);
or U6613 (N_6613,N_6598,N_6547);
or U6614 (N_6614,N_6409,N_6413);
and U6615 (N_6615,N_6480,N_6493);
nand U6616 (N_6616,N_6570,N_6429);
or U6617 (N_6617,N_6513,N_6473);
or U6618 (N_6618,N_6506,N_6422);
or U6619 (N_6619,N_6460,N_6565);
xor U6620 (N_6620,N_6463,N_6483);
nor U6621 (N_6621,N_6491,N_6438);
xnor U6622 (N_6622,N_6540,N_6533);
nor U6623 (N_6623,N_6535,N_6486);
and U6624 (N_6624,N_6449,N_6580);
xnor U6625 (N_6625,N_6470,N_6498);
nand U6626 (N_6626,N_6410,N_6545);
and U6627 (N_6627,N_6402,N_6595);
xor U6628 (N_6628,N_6457,N_6407);
or U6629 (N_6629,N_6559,N_6435);
or U6630 (N_6630,N_6445,N_6536);
and U6631 (N_6631,N_6476,N_6455);
and U6632 (N_6632,N_6412,N_6577);
nand U6633 (N_6633,N_6425,N_6494);
nor U6634 (N_6634,N_6496,N_6538);
or U6635 (N_6635,N_6458,N_6427);
or U6636 (N_6636,N_6514,N_6501);
or U6637 (N_6637,N_6500,N_6419);
and U6638 (N_6638,N_6448,N_6426);
xnor U6639 (N_6639,N_6437,N_6592);
xnor U6640 (N_6640,N_6594,N_6554);
nor U6641 (N_6641,N_6589,N_6466);
and U6642 (N_6642,N_6542,N_6446);
nand U6643 (N_6643,N_6581,N_6564);
and U6644 (N_6644,N_6439,N_6444);
nand U6645 (N_6645,N_6421,N_6502);
nand U6646 (N_6646,N_6572,N_6518);
and U6647 (N_6647,N_6550,N_6515);
nor U6648 (N_6648,N_6417,N_6593);
nand U6649 (N_6649,N_6436,N_6497);
or U6650 (N_6650,N_6451,N_6424);
or U6651 (N_6651,N_6597,N_6588);
xor U6652 (N_6652,N_6548,N_6440);
nor U6653 (N_6653,N_6411,N_6558);
nand U6654 (N_6654,N_6400,N_6482);
nor U6655 (N_6655,N_6467,N_6517);
xnor U6656 (N_6656,N_6406,N_6504);
or U6657 (N_6657,N_6599,N_6557);
and U6658 (N_6658,N_6568,N_6531);
nand U6659 (N_6659,N_6456,N_6587);
xnor U6660 (N_6660,N_6553,N_6528);
nand U6661 (N_6661,N_6462,N_6546);
nor U6662 (N_6662,N_6420,N_6590);
nor U6663 (N_6663,N_6443,N_6441);
or U6664 (N_6664,N_6405,N_6573);
xor U6665 (N_6665,N_6520,N_6465);
nand U6666 (N_6666,N_6453,N_6527);
and U6667 (N_6667,N_6471,N_6512);
and U6668 (N_6668,N_6534,N_6415);
or U6669 (N_6669,N_6526,N_6433);
or U6670 (N_6670,N_6403,N_6428);
or U6671 (N_6671,N_6525,N_6562);
xor U6672 (N_6672,N_6537,N_6539);
xnor U6673 (N_6673,N_6584,N_6522);
or U6674 (N_6674,N_6485,N_6519);
nand U6675 (N_6675,N_6586,N_6452);
or U6676 (N_6676,N_6487,N_6464);
nand U6677 (N_6677,N_6474,N_6508);
or U6678 (N_6678,N_6408,N_6479);
xnor U6679 (N_6679,N_6477,N_6423);
nand U6680 (N_6680,N_6544,N_6543);
or U6681 (N_6681,N_6468,N_6475);
xor U6682 (N_6682,N_6499,N_6549);
nand U6683 (N_6683,N_6434,N_6414);
and U6684 (N_6684,N_6524,N_6481);
and U6685 (N_6685,N_6418,N_6530);
nand U6686 (N_6686,N_6578,N_6489);
xnor U6687 (N_6687,N_6596,N_6442);
nand U6688 (N_6688,N_6454,N_6560);
xor U6689 (N_6689,N_6492,N_6574);
or U6690 (N_6690,N_6450,N_6569);
and U6691 (N_6691,N_6461,N_6472);
or U6692 (N_6692,N_6495,N_6507);
nand U6693 (N_6693,N_6591,N_6556);
or U6694 (N_6694,N_6469,N_6555);
nor U6695 (N_6695,N_6575,N_6583);
or U6696 (N_6696,N_6459,N_6484);
xor U6697 (N_6697,N_6488,N_6532);
or U6698 (N_6698,N_6582,N_6516);
xnor U6699 (N_6699,N_6490,N_6541);
or U6700 (N_6700,N_6562,N_6494);
or U6701 (N_6701,N_6467,N_6585);
nor U6702 (N_6702,N_6427,N_6489);
nand U6703 (N_6703,N_6537,N_6594);
nor U6704 (N_6704,N_6560,N_6491);
xor U6705 (N_6705,N_6468,N_6588);
nand U6706 (N_6706,N_6556,N_6436);
or U6707 (N_6707,N_6520,N_6563);
xnor U6708 (N_6708,N_6579,N_6503);
nor U6709 (N_6709,N_6479,N_6477);
or U6710 (N_6710,N_6574,N_6595);
xor U6711 (N_6711,N_6409,N_6527);
or U6712 (N_6712,N_6508,N_6480);
nor U6713 (N_6713,N_6501,N_6444);
nor U6714 (N_6714,N_6596,N_6592);
nand U6715 (N_6715,N_6597,N_6419);
or U6716 (N_6716,N_6406,N_6437);
xnor U6717 (N_6717,N_6419,N_6536);
xnor U6718 (N_6718,N_6586,N_6403);
nor U6719 (N_6719,N_6516,N_6545);
nand U6720 (N_6720,N_6462,N_6475);
and U6721 (N_6721,N_6486,N_6413);
xnor U6722 (N_6722,N_6551,N_6569);
nor U6723 (N_6723,N_6428,N_6439);
and U6724 (N_6724,N_6445,N_6564);
xor U6725 (N_6725,N_6412,N_6571);
or U6726 (N_6726,N_6564,N_6569);
or U6727 (N_6727,N_6568,N_6514);
and U6728 (N_6728,N_6422,N_6497);
xor U6729 (N_6729,N_6452,N_6476);
and U6730 (N_6730,N_6478,N_6400);
xor U6731 (N_6731,N_6444,N_6457);
nand U6732 (N_6732,N_6487,N_6598);
or U6733 (N_6733,N_6425,N_6553);
xnor U6734 (N_6734,N_6436,N_6424);
nor U6735 (N_6735,N_6575,N_6408);
or U6736 (N_6736,N_6498,N_6539);
xor U6737 (N_6737,N_6509,N_6547);
nor U6738 (N_6738,N_6457,N_6414);
xor U6739 (N_6739,N_6541,N_6515);
xor U6740 (N_6740,N_6512,N_6444);
xnor U6741 (N_6741,N_6547,N_6558);
and U6742 (N_6742,N_6487,N_6496);
and U6743 (N_6743,N_6562,N_6585);
or U6744 (N_6744,N_6570,N_6466);
xnor U6745 (N_6745,N_6581,N_6416);
or U6746 (N_6746,N_6400,N_6524);
and U6747 (N_6747,N_6501,N_6423);
and U6748 (N_6748,N_6599,N_6528);
nor U6749 (N_6749,N_6468,N_6467);
xor U6750 (N_6750,N_6419,N_6530);
nor U6751 (N_6751,N_6517,N_6535);
and U6752 (N_6752,N_6543,N_6595);
and U6753 (N_6753,N_6586,N_6523);
nor U6754 (N_6754,N_6461,N_6541);
nor U6755 (N_6755,N_6581,N_6557);
nand U6756 (N_6756,N_6522,N_6473);
and U6757 (N_6757,N_6546,N_6570);
and U6758 (N_6758,N_6409,N_6580);
or U6759 (N_6759,N_6501,N_6559);
nand U6760 (N_6760,N_6535,N_6402);
nand U6761 (N_6761,N_6495,N_6440);
nand U6762 (N_6762,N_6492,N_6439);
and U6763 (N_6763,N_6573,N_6531);
xnor U6764 (N_6764,N_6439,N_6593);
nor U6765 (N_6765,N_6422,N_6460);
nand U6766 (N_6766,N_6526,N_6543);
nor U6767 (N_6767,N_6509,N_6508);
or U6768 (N_6768,N_6548,N_6435);
or U6769 (N_6769,N_6407,N_6596);
or U6770 (N_6770,N_6538,N_6439);
xnor U6771 (N_6771,N_6442,N_6531);
and U6772 (N_6772,N_6420,N_6513);
nor U6773 (N_6773,N_6574,N_6592);
nor U6774 (N_6774,N_6517,N_6547);
or U6775 (N_6775,N_6592,N_6514);
xor U6776 (N_6776,N_6428,N_6464);
nor U6777 (N_6777,N_6450,N_6447);
nand U6778 (N_6778,N_6435,N_6418);
nor U6779 (N_6779,N_6481,N_6541);
or U6780 (N_6780,N_6462,N_6401);
nor U6781 (N_6781,N_6499,N_6521);
xnor U6782 (N_6782,N_6592,N_6483);
xor U6783 (N_6783,N_6498,N_6490);
xor U6784 (N_6784,N_6425,N_6514);
xor U6785 (N_6785,N_6465,N_6458);
nor U6786 (N_6786,N_6507,N_6467);
and U6787 (N_6787,N_6523,N_6484);
nor U6788 (N_6788,N_6582,N_6432);
xnor U6789 (N_6789,N_6558,N_6522);
xnor U6790 (N_6790,N_6554,N_6504);
nor U6791 (N_6791,N_6550,N_6598);
or U6792 (N_6792,N_6537,N_6438);
or U6793 (N_6793,N_6562,N_6545);
xnor U6794 (N_6794,N_6511,N_6592);
xnor U6795 (N_6795,N_6469,N_6574);
xor U6796 (N_6796,N_6558,N_6434);
or U6797 (N_6797,N_6493,N_6575);
nand U6798 (N_6798,N_6569,N_6562);
nor U6799 (N_6799,N_6478,N_6588);
xor U6800 (N_6800,N_6624,N_6759);
and U6801 (N_6801,N_6727,N_6601);
nor U6802 (N_6802,N_6777,N_6616);
and U6803 (N_6803,N_6756,N_6744);
nor U6804 (N_6804,N_6700,N_6717);
xnor U6805 (N_6805,N_6668,N_6607);
and U6806 (N_6806,N_6741,N_6724);
nand U6807 (N_6807,N_6602,N_6653);
or U6808 (N_6808,N_6618,N_6775);
and U6809 (N_6809,N_6651,N_6694);
and U6810 (N_6810,N_6675,N_6630);
nor U6811 (N_6811,N_6726,N_6712);
or U6812 (N_6812,N_6695,N_6768);
xnor U6813 (N_6813,N_6797,N_6626);
or U6814 (N_6814,N_6605,N_6677);
and U6815 (N_6815,N_6764,N_6765);
or U6816 (N_6816,N_6696,N_6687);
nor U6817 (N_6817,N_6753,N_6705);
xor U6818 (N_6818,N_6662,N_6736);
nand U6819 (N_6819,N_6725,N_6609);
or U6820 (N_6820,N_6690,N_6779);
and U6821 (N_6821,N_6711,N_6789);
nor U6822 (N_6822,N_6722,N_6785);
nand U6823 (N_6823,N_6621,N_6782);
and U6824 (N_6824,N_6676,N_6619);
nand U6825 (N_6825,N_6629,N_6663);
xor U6826 (N_6826,N_6702,N_6778);
nor U6827 (N_6827,N_6754,N_6718);
or U6828 (N_6828,N_6732,N_6612);
nor U6829 (N_6829,N_6666,N_6661);
xnor U6830 (N_6830,N_6739,N_6790);
nand U6831 (N_6831,N_6650,N_6640);
xnor U6832 (N_6832,N_6706,N_6610);
nand U6833 (N_6833,N_6615,N_6699);
xor U6834 (N_6834,N_6625,N_6709);
nor U6835 (N_6835,N_6637,N_6784);
nand U6836 (N_6836,N_6781,N_6620);
nand U6837 (N_6837,N_6792,N_6600);
or U6838 (N_6838,N_6787,N_6627);
nor U6839 (N_6839,N_6762,N_6691);
xnor U6840 (N_6840,N_6667,N_6755);
or U6841 (N_6841,N_6780,N_6721);
or U6842 (N_6842,N_6758,N_6730);
and U6843 (N_6843,N_6632,N_6728);
nor U6844 (N_6844,N_6684,N_6798);
nor U6845 (N_6845,N_6611,N_6652);
or U6846 (N_6846,N_6643,N_6763);
nand U6847 (N_6847,N_6740,N_6751);
or U6848 (N_6848,N_6719,N_6729);
nor U6849 (N_6849,N_6664,N_6743);
nand U6850 (N_6850,N_6704,N_6688);
nor U6851 (N_6851,N_6760,N_6654);
nand U6852 (N_6852,N_6681,N_6749);
xnor U6853 (N_6853,N_6686,N_6701);
or U6854 (N_6854,N_6660,N_6669);
or U6855 (N_6855,N_6613,N_6670);
or U6856 (N_6856,N_6693,N_6734);
nand U6857 (N_6857,N_6772,N_6748);
nand U6858 (N_6858,N_6648,N_6707);
and U6859 (N_6859,N_6692,N_6647);
xor U6860 (N_6860,N_6769,N_6634);
or U6861 (N_6861,N_6794,N_6622);
and U6862 (N_6862,N_6714,N_6606);
nand U6863 (N_6863,N_6678,N_6680);
nand U6864 (N_6864,N_6703,N_6671);
and U6865 (N_6865,N_6731,N_6655);
nand U6866 (N_6866,N_6710,N_6673);
nand U6867 (N_6867,N_6766,N_6635);
nor U6868 (N_6868,N_6665,N_6672);
nor U6869 (N_6869,N_6715,N_6708);
nor U6870 (N_6870,N_6747,N_6776);
nor U6871 (N_6871,N_6656,N_6738);
nand U6872 (N_6872,N_6657,N_6761);
xor U6873 (N_6873,N_6604,N_6639);
nand U6874 (N_6874,N_6659,N_6698);
or U6875 (N_6875,N_6791,N_6771);
or U6876 (N_6876,N_6737,N_6644);
nand U6877 (N_6877,N_6716,N_6735);
and U6878 (N_6878,N_6603,N_6750);
nand U6879 (N_6879,N_6679,N_6742);
xor U6880 (N_6880,N_6689,N_6649);
nor U6881 (N_6881,N_6793,N_6642);
or U6882 (N_6882,N_6633,N_6788);
nor U6883 (N_6883,N_6773,N_6631);
and U6884 (N_6884,N_6723,N_6733);
nand U6885 (N_6885,N_6623,N_6799);
or U6886 (N_6886,N_6697,N_6770);
nor U6887 (N_6887,N_6617,N_6746);
xor U6888 (N_6888,N_6645,N_6614);
xnor U6889 (N_6889,N_6641,N_6636);
and U6890 (N_6890,N_6685,N_6638);
nor U6891 (N_6891,N_6674,N_6713);
nand U6892 (N_6892,N_6783,N_6745);
and U6893 (N_6893,N_6608,N_6767);
nand U6894 (N_6894,N_6796,N_6683);
nand U6895 (N_6895,N_6628,N_6752);
and U6896 (N_6896,N_6774,N_6682);
nand U6897 (N_6897,N_6720,N_6757);
xor U6898 (N_6898,N_6658,N_6786);
and U6899 (N_6899,N_6795,N_6646);
and U6900 (N_6900,N_6608,N_6644);
and U6901 (N_6901,N_6656,N_6726);
and U6902 (N_6902,N_6656,N_6701);
nand U6903 (N_6903,N_6701,N_6728);
nand U6904 (N_6904,N_6690,N_6643);
nand U6905 (N_6905,N_6620,N_6658);
xor U6906 (N_6906,N_6761,N_6721);
or U6907 (N_6907,N_6707,N_6710);
nand U6908 (N_6908,N_6672,N_6662);
and U6909 (N_6909,N_6617,N_6680);
xnor U6910 (N_6910,N_6749,N_6652);
and U6911 (N_6911,N_6662,N_6659);
xor U6912 (N_6912,N_6621,N_6795);
nor U6913 (N_6913,N_6730,N_6702);
and U6914 (N_6914,N_6796,N_6700);
or U6915 (N_6915,N_6673,N_6653);
xor U6916 (N_6916,N_6797,N_6714);
nor U6917 (N_6917,N_6668,N_6729);
and U6918 (N_6918,N_6677,N_6622);
xor U6919 (N_6919,N_6641,N_6603);
or U6920 (N_6920,N_6610,N_6651);
or U6921 (N_6921,N_6611,N_6610);
nand U6922 (N_6922,N_6756,N_6776);
xor U6923 (N_6923,N_6730,N_6733);
xor U6924 (N_6924,N_6685,N_6661);
and U6925 (N_6925,N_6748,N_6607);
or U6926 (N_6926,N_6692,N_6739);
or U6927 (N_6927,N_6675,N_6605);
and U6928 (N_6928,N_6713,N_6632);
nor U6929 (N_6929,N_6781,N_6663);
xor U6930 (N_6930,N_6617,N_6762);
nor U6931 (N_6931,N_6709,N_6762);
nand U6932 (N_6932,N_6736,N_6626);
nor U6933 (N_6933,N_6667,N_6631);
or U6934 (N_6934,N_6771,N_6613);
nor U6935 (N_6935,N_6727,N_6742);
nand U6936 (N_6936,N_6779,N_6650);
nand U6937 (N_6937,N_6720,N_6727);
xnor U6938 (N_6938,N_6612,N_6739);
and U6939 (N_6939,N_6710,N_6609);
nor U6940 (N_6940,N_6604,N_6788);
and U6941 (N_6941,N_6691,N_6730);
xnor U6942 (N_6942,N_6685,N_6715);
nor U6943 (N_6943,N_6607,N_6747);
nand U6944 (N_6944,N_6775,N_6772);
or U6945 (N_6945,N_6624,N_6747);
nand U6946 (N_6946,N_6682,N_6702);
nor U6947 (N_6947,N_6622,N_6750);
nand U6948 (N_6948,N_6724,N_6668);
and U6949 (N_6949,N_6618,N_6696);
or U6950 (N_6950,N_6604,N_6778);
or U6951 (N_6951,N_6645,N_6729);
nor U6952 (N_6952,N_6655,N_6600);
or U6953 (N_6953,N_6684,N_6661);
or U6954 (N_6954,N_6754,N_6687);
and U6955 (N_6955,N_6760,N_6634);
nor U6956 (N_6956,N_6782,N_6647);
xor U6957 (N_6957,N_6705,N_6782);
and U6958 (N_6958,N_6654,N_6682);
nand U6959 (N_6959,N_6767,N_6765);
nand U6960 (N_6960,N_6600,N_6612);
nor U6961 (N_6961,N_6778,N_6728);
xor U6962 (N_6962,N_6708,N_6621);
or U6963 (N_6963,N_6738,N_6795);
nor U6964 (N_6964,N_6759,N_6645);
and U6965 (N_6965,N_6706,N_6623);
nor U6966 (N_6966,N_6652,N_6798);
xnor U6967 (N_6967,N_6681,N_6797);
and U6968 (N_6968,N_6670,N_6797);
nor U6969 (N_6969,N_6770,N_6708);
or U6970 (N_6970,N_6635,N_6760);
nand U6971 (N_6971,N_6652,N_6711);
nand U6972 (N_6972,N_6669,N_6620);
and U6973 (N_6973,N_6788,N_6786);
xor U6974 (N_6974,N_6670,N_6750);
or U6975 (N_6975,N_6624,N_6775);
nor U6976 (N_6976,N_6767,N_6777);
xor U6977 (N_6977,N_6728,N_6742);
xnor U6978 (N_6978,N_6640,N_6737);
and U6979 (N_6979,N_6655,N_6610);
nand U6980 (N_6980,N_6732,N_6707);
xor U6981 (N_6981,N_6655,N_6675);
or U6982 (N_6982,N_6693,N_6743);
or U6983 (N_6983,N_6661,N_6656);
or U6984 (N_6984,N_6628,N_6780);
nand U6985 (N_6985,N_6659,N_6733);
xor U6986 (N_6986,N_6720,N_6722);
nand U6987 (N_6987,N_6717,N_6750);
or U6988 (N_6988,N_6708,N_6745);
nand U6989 (N_6989,N_6645,N_6707);
xnor U6990 (N_6990,N_6715,N_6723);
and U6991 (N_6991,N_6688,N_6709);
and U6992 (N_6992,N_6685,N_6798);
or U6993 (N_6993,N_6760,N_6636);
nor U6994 (N_6994,N_6777,N_6621);
nand U6995 (N_6995,N_6742,N_6763);
or U6996 (N_6996,N_6691,N_6729);
or U6997 (N_6997,N_6656,N_6737);
and U6998 (N_6998,N_6731,N_6723);
nand U6999 (N_6999,N_6642,N_6667);
or U7000 (N_7000,N_6983,N_6979);
or U7001 (N_7001,N_6914,N_6810);
or U7002 (N_7002,N_6833,N_6921);
and U7003 (N_7003,N_6895,N_6869);
and U7004 (N_7004,N_6875,N_6959);
and U7005 (N_7005,N_6879,N_6864);
xnor U7006 (N_7006,N_6840,N_6847);
or U7007 (N_7007,N_6872,N_6988);
nand U7008 (N_7008,N_6962,N_6993);
xor U7009 (N_7009,N_6890,N_6876);
xor U7010 (N_7010,N_6984,N_6897);
nor U7011 (N_7011,N_6991,N_6995);
and U7012 (N_7012,N_6965,N_6853);
and U7013 (N_7013,N_6913,N_6968);
xnor U7014 (N_7014,N_6807,N_6849);
and U7015 (N_7015,N_6923,N_6973);
nand U7016 (N_7016,N_6905,N_6911);
xnor U7017 (N_7017,N_6883,N_6850);
or U7018 (N_7018,N_6801,N_6811);
xnor U7019 (N_7019,N_6990,N_6892);
and U7020 (N_7020,N_6867,N_6824);
xnor U7021 (N_7021,N_6981,N_6814);
or U7022 (N_7022,N_6842,N_6808);
xor U7023 (N_7023,N_6956,N_6975);
xnor U7024 (N_7024,N_6932,N_6936);
nand U7025 (N_7025,N_6951,N_6955);
or U7026 (N_7026,N_6865,N_6862);
nor U7027 (N_7027,N_6907,N_6901);
nand U7028 (N_7028,N_6925,N_6917);
or U7029 (N_7029,N_6896,N_6976);
nor U7030 (N_7030,N_6947,N_6967);
nand U7031 (N_7031,N_6845,N_6848);
nor U7032 (N_7032,N_6891,N_6916);
and U7033 (N_7033,N_6885,N_6819);
and U7034 (N_7034,N_6858,N_6929);
xnor U7035 (N_7035,N_6812,N_6945);
xnor U7036 (N_7036,N_6823,N_6860);
xnor U7037 (N_7037,N_6884,N_6871);
xnor U7038 (N_7038,N_6974,N_6870);
nor U7039 (N_7039,N_6886,N_6894);
xnor U7040 (N_7040,N_6924,N_6844);
and U7041 (N_7041,N_6934,N_6903);
nand U7042 (N_7042,N_6828,N_6822);
nand U7043 (N_7043,N_6900,N_6971);
and U7044 (N_7044,N_6994,N_6928);
or U7045 (N_7045,N_6950,N_6857);
or U7046 (N_7046,N_6904,N_6941);
xor U7047 (N_7047,N_6852,N_6989);
nor U7048 (N_7048,N_6922,N_6918);
and U7049 (N_7049,N_6826,N_6966);
nand U7050 (N_7050,N_6952,N_6832);
and U7051 (N_7051,N_6818,N_6957);
nor U7052 (N_7052,N_6898,N_6958);
or U7053 (N_7053,N_6915,N_6909);
or U7054 (N_7054,N_6863,N_6882);
nor U7055 (N_7055,N_6809,N_6821);
nor U7056 (N_7056,N_6825,N_6873);
nand U7057 (N_7057,N_6972,N_6817);
nand U7058 (N_7058,N_6881,N_6888);
or U7059 (N_7059,N_6940,N_6838);
nand U7060 (N_7060,N_6906,N_6953);
nand U7061 (N_7061,N_6893,N_6815);
and U7062 (N_7062,N_6946,N_6910);
nand U7063 (N_7063,N_6987,N_6887);
xnor U7064 (N_7064,N_6943,N_6927);
nor U7065 (N_7065,N_6949,N_6980);
nand U7066 (N_7066,N_6912,N_6839);
nor U7067 (N_7067,N_6859,N_6837);
nor U7068 (N_7068,N_6816,N_6834);
or U7069 (N_7069,N_6964,N_6830);
or U7070 (N_7070,N_6954,N_6846);
or U7071 (N_7071,N_6942,N_6866);
nor U7072 (N_7072,N_6829,N_6899);
or U7073 (N_7073,N_6986,N_6803);
nor U7074 (N_7074,N_6970,N_6982);
or U7075 (N_7075,N_6856,N_6868);
or U7076 (N_7076,N_6841,N_6806);
xor U7077 (N_7077,N_6919,N_6935);
or U7078 (N_7078,N_6938,N_6851);
or U7079 (N_7079,N_6835,N_6861);
nor U7080 (N_7080,N_6939,N_6937);
and U7081 (N_7081,N_6978,N_6800);
and U7082 (N_7082,N_6855,N_6963);
and U7083 (N_7083,N_6969,N_6908);
or U7084 (N_7084,N_6985,N_6960);
nand U7085 (N_7085,N_6992,N_6854);
and U7086 (N_7086,N_6802,N_6944);
xor U7087 (N_7087,N_6977,N_6933);
and U7088 (N_7088,N_6880,N_6930);
or U7089 (N_7089,N_6813,N_6831);
or U7090 (N_7090,N_6804,N_6827);
xnor U7091 (N_7091,N_6961,N_6997);
nor U7092 (N_7092,N_6998,N_6889);
nor U7093 (N_7093,N_6902,N_6820);
and U7094 (N_7094,N_6948,N_6836);
nor U7095 (N_7095,N_6843,N_6805);
nor U7096 (N_7096,N_6931,N_6877);
or U7097 (N_7097,N_6878,N_6874);
or U7098 (N_7098,N_6999,N_6996);
nand U7099 (N_7099,N_6926,N_6920);
nor U7100 (N_7100,N_6843,N_6893);
nor U7101 (N_7101,N_6884,N_6994);
xnor U7102 (N_7102,N_6966,N_6976);
nor U7103 (N_7103,N_6953,N_6963);
nand U7104 (N_7104,N_6902,N_6914);
nand U7105 (N_7105,N_6920,N_6921);
nor U7106 (N_7106,N_6829,N_6861);
and U7107 (N_7107,N_6990,N_6830);
nand U7108 (N_7108,N_6802,N_6989);
or U7109 (N_7109,N_6978,N_6899);
nand U7110 (N_7110,N_6885,N_6973);
or U7111 (N_7111,N_6869,N_6853);
nand U7112 (N_7112,N_6960,N_6903);
nand U7113 (N_7113,N_6810,N_6806);
and U7114 (N_7114,N_6967,N_6849);
nand U7115 (N_7115,N_6876,N_6871);
nand U7116 (N_7116,N_6819,N_6992);
nor U7117 (N_7117,N_6912,N_6841);
or U7118 (N_7118,N_6900,N_6995);
nand U7119 (N_7119,N_6824,N_6868);
nand U7120 (N_7120,N_6814,N_6908);
and U7121 (N_7121,N_6923,N_6842);
nor U7122 (N_7122,N_6870,N_6959);
xor U7123 (N_7123,N_6822,N_6840);
or U7124 (N_7124,N_6804,N_6894);
nor U7125 (N_7125,N_6865,N_6934);
xor U7126 (N_7126,N_6835,N_6916);
or U7127 (N_7127,N_6821,N_6879);
nor U7128 (N_7128,N_6968,N_6903);
or U7129 (N_7129,N_6962,N_6940);
nor U7130 (N_7130,N_6897,N_6842);
and U7131 (N_7131,N_6844,N_6822);
nand U7132 (N_7132,N_6870,N_6901);
and U7133 (N_7133,N_6981,N_6998);
or U7134 (N_7134,N_6940,N_6993);
nor U7135 (N_7135,N_6827,N_6853);
nand U7136 (N_7136,N_6869,N_6863);
nand U7137 (N_7137,N_6924,N_6806);
xnor U7138 (N_7138,N_6869,N_6847);
nor U7139 (N_7139,N_6924,N_6941);
and U7140 (N_7140,N_6950,N_6847);
xor U7141 (N_7141,N_6859,N_6897);
or U7142 (N_7142,N_6803,N_6844);
nor U7143 (N_7143,N_6896,N_6878);
and U7144 (N_7144,N_6834,N_6882);
and U7145 (N_7145,N_6952,N_6895);
xor U7146 (N_7146,N_6952,N_6800);
and U7147 (N_7147,N_6900,N_6859);
nor U7148 (N_7148,N_6860,N_6815);
nor U7149 (N_7149,N_6976,N_6811);
nand U7150 (N_7150,N_6887,N_6818);
and U7151 (N_7151,N_6969,N_6856);
nor U7152 (N_7152,N_6902,N_6951);
nand U7153 (N_7153,N_6994,N_6963);
and U7154 (N_7154,N_6853,N_6839);
nor U7155 (N_7155,N_6993,N_6898);
nor U7156 (N_7156,N_6804,N_6874);
xnor U7157 (N_7157,N_6866,N_6834);
or U7158 (N_7158,N_6812,N_6820);
xnor U7159 (N_7159,N_6960,N_6818);
xnor U7160 (N_7160,N_6910,N_6964);
nor U7161 (N_7161,N_6979,N_6986);
and U7162 (N_7162,N_6882,N_6835);
and U7163 (N_7163,N_6820,N_6992);
xnor U7164 (N_7164,N_6992,N_6973);
nor U7165 (N_7165,N_6979,N_6931);
and U7166 (N_7166,N_6934,N_6911);
or U7167 (N_7167,N_6959,N_6803);
xor U7168 (N_7168,N_6909,N_6812);
xnor U7169 (N_7169,N_6899,N_6950);
nand U7170 (N_7170,N_6968,N_6844);
nor U7171 (N_7171,N_6871,N_6863);
xor U7172 (N_7172,N_6908,N_6953);
and U7173 (N_7173,N_6939,N_6990);
nor U7174 (N_7174,N_6903,N_6973);
nand U7175 (N_7175,N_6864,N_6963);
and U7176 (N_7176,N_6939,N_6968);
nand U7177 (N_7177,N_6824,N_6903);
nor U7178 (N_7178,N_6984,N_6817);
nor U7179 (N_7179,N_6862,N_6802);
nor U7180 (N_7180,N_6979,N_6815);
and U7181 (N_7181,N_6810,N_6878);
and U7182 (N_7182,N_6808,N_6896);
nor U7183 (N_7183,N_6938,N_6899);
and U7184 (N_7184,N_6893,N_6958);
and U7185 (N_7185,N_6990,N_6885);
and U7186 (N_7186,N_6863,N_6804);
nand U7187 (N_7187,N_6863,N_6995);
xor U7188 (N_7188,N_6837,N_6948);
nand U7189 (N_7189,N_6817,N_6895);
nand U7190 (N_7190,N_6864,N_6924);
xor U7191 (N_7191,N_6921,N_6953);
nand U7192 (N_7192,N_6914,N_6822);
nor U7193 (N_7193,N_6970,N_6831);
or U7194 (N_7194,N_6965,N_6895);
nor U7195 (N_7195,N_6872,N_6938);
nor U7196 (N_7196,N_6891,N_6808);
nor U7197 (N_7197,N_6847,N_6856);
nand U7198 (N_7198,N_6859,N_6817);
nor U7199 (N_7199,N_6913,N_6840);
xor U7200 (N_7200,N_7015,N_7081);
or U7201 (N_7201,N_7151,N_7135);
nand U7202 (N_7202,N_7193,N_7107);
and U7203 (N_7203,N_7000,N_7053);
and U7204 (N_7204,N_7089,N_7019);
nor U7205 (N_7205,N_7162,N_7097);
xor U7206 (N_7206,N_7144,N_7103);
and U7207 (N_7207,N_7030,N_7154);
nor U7208 (N_7208,N_7042,N_7014);
or U7209 (N_7209,N_7029,N_7186);
nand U7210 (N_7210,N_7190,N_7141);
nor U7211 (N_7211,N_7159,N_7163);
and U7212 (N_7212,N_7018,N_7196);
nand U7213 (N_7213,N_7001,N_7013);
xor U7214 (N_7214,N_7062,N_7026);
nand U7215 (N_7215,N_7145,N_7056);
nand U7216 (N_7216,N_7198,N_7124);
nand U7217 (N_7217,N_7038,N_7058);
xor U7218 (N_7218,N_7007,N_7125);
nor U7219 (N_7219,N_7118,N_7130);
or U7220 (N_7220,N_7121,N_7132);
nand U7221 (N_7221,N_7104,N_7101);
xnor U7222 (N_7222,N_7067,N_7194);
or U7223 (N_7223,N_7158,N_7192);
xor U7224 (N_7224,N_7037,N_7075);
xnor U7225 (N_7225,N_7040,N_7137);
nor U7226 (N_7226,N_7028,N_7105);
nand U7227 (N_7227,N_7108,N_7100);
xor U7228 (N_7228,N_7073,N_7178);
or U7229 (N_7229,N_7087,N_7168);
or U7230 (N_7230,N_7150,N_7164);
xnor U7231 (N_7231,N_7115,N_7091);
nand U7232 (N_7232,N_7039,N_7094);
or U7233 (N_7233,N_7191,N_7183);
nor U7234 (N_7234,N_7140,N_7012);
nor U7235 (N_7235,N_7063,N_7035);
nand U7236 (N_7236,N_7195,N_7139);
xor U7237 (N_7237,N_7057,N_7070);
and U7238 (N_7238,N_7156,N_7123);
nor U7239 (N_7239,N_7043,N_7095);
or U7240 (N_7240,N_7021,N_7004);
xor U7241 (N_7241,N_7051,N_7093);
nand U7242 (N_7242,N_7110,N_7120);
xnor U7243 (N_7243,N_7086,N_7134);
nand U7244 (N_7244,N_7016,N_7047);
nand U7245 (N_7245,N_7003,N_7061);
or U7246 (N_7246,N_7082,N_7020);
nor U7247 (N_7247,N_7024,N_7076);
or U7248 (N_7248,N_7153,N_7055);
xor U7249 (N_7249,N_7128,N_7078);
and U7250 (N_7250,N_7175,N_7098);
and U7251 (N_7251,N_7152,N_7023);
and U7252 (N_7252,N_7079,N_7165);
nor U7253 (N_7253,N_7011,N_7117);
or U7254 (N_7254,N_7064,N_7069);
and U7255 (N_7255,N_7025,N_7199);
or U7256 (N_7256,N_7188,N_7032);
nor U7257 (N_7257,N_7169,N_7109);
nor U7258 (N_7258,N_7072,N_7142);
or U7259 (N_7259,N_7092,N_7197);
and U7260 (N_7260,N_7189,N_7049);
nand U7261 (N_7261,N_7031,N_7155);
and U7262 (N_7262,N_7147,N_7184);
nand U7263 (N_7263,N_7090,N_7002);
and U7264 (N_7264,N_7041,N_7113);
nor U7265 (N_7265,N_7022,N_7084);
nor U7266 (N_7266,N_7046,N_7157);
xor U7267 (N_7267,N_7114,N_7085);
xnor U7268 (N_7268,N_7182,N_7096);
nor U7269 (N_7269,N_7080,N_7112);
and U7270 (N_7270,N_7181,N_7111);
xor U7271 (N_7271,N_7008,N_7172);
and U7272 (N_7272,N_7045,N_7102);
or U7273 (N_7273,N_7033,N_7074);
nor U7274 (N_7274,N_7177,N_7127);
xnor U7275 (N_7275,N_7170,N_7116);
or U7276 (N_7276,N_7167,N_7060);
nor U7277 (N_7277,N_7068,N_7143);
nor U7278 (N_7278,N_7166,N_7174);
nor U7279 (N_7279,N_7083,N_7148);
nand U7280 (N_7280,N_7131,N_7050);
or U7281 (N_7281,N_7005,N_7149);
xor U7282 (N_7282,N_7034,N_7146);
or U7283 (N_7283,N_7106,N_7133);
and U7284 (N_7284,N_7187,N_7044);
nor U7285 (N_7285,N_7010,N_7129);
and U7286 (N_7286,N_7071,N_7138);
and U7287 (N_7287,N_7179,N_7054);
nand U7288 (N_7288,N_7122,N_7017);
or U7289 (N_7289,N_7059,N_7173);
nor U7290 (N_7290,N_7077,N_7160);
nor U7291 (N_7291,N_7088,N_7006);
nand U7292 (N_7292,N_7066,N_7176);
or U7293 (N_7293,N_7119,N_7036);
xor U7294 (N_7294,N_7126,N_7065);
and U7295 (N_7295,N_7009,N_7180);
and U7296 (N_7296,N_7161,N_7027);
and U7297 (N_7297,N_7099,N_7052);
and U7298 (N_7298,N_7136,N_7171);
nand U7299 (N_7299,N_7185,N_7048);
xnor U7300 (N_7300,N_7157,N_7034);
xnor U7301 (N_7301,N_7194,N_7098);
or U7302 (N_7302,N_7125,N_7005);
and U7303 (N_7303,N_7018,N_7076);
nor U7304 (N_7304,N_7042,N_7118);
or U7305 (N_7305,N_7087,N_7018);
nand U7306 (N_7306,N_7120,N_7053);
xor U7307 (N_7307,N_7175,N_7089);
nor U7308 (N_7308,N_7101,N_7070);
xnor U7309 (N_7309,N_7017,N_7052);
nand U7310 (N_7310,N_7166,N_7178);
xnor U7311 (N_7311,N_7077,N_7177);
or U7312 (N_7312,N_7027,N_7185);
or U7313 (N_7313,N_7084,N_7095);
and U7314 (N_7314,N_7159,N_7079);
nor U7315 (N_7315,N_7083,N_7062);
nor U7316 (N_7316,N_7094,N_7090);
and U7317 (N_7317,N_7180,N_7054);
nor U7318 (N_7318,N_7041,N_7002);
and U7319 (N_7319,N_7115,N_7118);
xor U7320 (N_7320,N_7061,N_7139);
nand U7321 (N_7321,N_7001,N_7100);
and U7322 (N_7322,N_7133,N_7115);
nand U7323 (N_7323,N_7117,N_7010);
or U7324 (N_7324,N_7082,N_7141);
and U7325 (N_7325,N_7144,N_7148);
nand U7326 (N_7326,N_7075,N_7181);
nand U7327 (N_7327,N_7023,N_7025);
nor U7328 (N_7328,N_7184,N_7089);
nor U7329 (N_7329,N_7114,N_7188);
nor U7330 (N_7330,N_7129,N_7087);
and U7331 (N_7331,N_7145,N_7177);
xnor U7332 (N_7332,N_7045,N_7130);
and U7333 (N_7333,N_7159,N_7015);
and U7334 (N_7334,N_7096,N_7106);
and U7335 (N_7335,N_7186,N_7052);
nor U7336 (N_7336,N_7183,N_7099);
and U7337 (N_7337,N_7153,N_7035);
xnor U7338 (N_7338,N_7006,N_7066);
nand U7339 (N_7339,N_7043,N_7194);
nor U7340 (N_7340,N_7076,N_7127);
nand U7341 (N_7341,N_7082,N_7173);
or U7342 (N_7342,N_7000,N_7008);
or U7343 (N_7343,N_7044,N_7026);
or U7344 (N_7344,N_7010,N_7136);
xnor U7345 (N_7345,N_7116,N_7007);
xor U7346 (N_7346,N_7143,N_7196);
or U7347 (N_7347,N_7020,N_7153);
nand U7348 (N_7348,N_7085,N_7187);
or U7349 (N_7349,N_7125,N_7049);
xor U7350 (N_7350,N_7088,N_7044);
xnor U7351 (N_7351,N_7055,N_7050);
nand U7352 (N_7352,N_7131,N_7058);
or U7353 (N_7353,N_7119,N_7030);
xnor U7354 (N_7354,N_7015,N_7169);
or U7355 (N_7355,N_7009,N_7082);
nor U7356 (N_7356,N_7074,N_7128);
nand U7357 (N_7357,N_7092,N_7042);
and U7358 (N_7358,N_7118,N_7038);
nand U7359 (N_7359,N_7007,N_7179);
and U7360 (N_7360,N_7076,N_7148);
or U7361 (N_7361,N_7123,N_7188);
or U7362 (N_7362,N_7101,N_7022);
nor U7363 (N_7363,N_7059,N_7011);
or U7364 (N_7364,N_7183,N_7149);
nor U7365 (N_7365,N_7124,N_7191);
nand U7366 (N_7366,N_7005,N_7012);
xnor U7367 (N_7367,N_7156,N_7013);
and U7368 (N_7368,N_7082,N_7076);
xor U7369 (N_7369,N_7032,N_7115);
or U7370 (N_7370,N_7006,N_7097);
nand U7371 (N_7371,N_7125,N_7128);
xnor U7372 (N_7372,N_7086,N_7044);
xor U7373 (N_7373,N_7025,N_7154);
xnor U7374 (N_7374,N_7039,N_7103);
nor U7375 (N_7375,N_7110,N_7135);
or U7376 (N_7376,N_7135,N_7012);
and U7377 (N_7377,N_7048,N_7040);
nor U7378 (N_7378,N_7067,N_7172);
and U7379 (N_7379,N_7187,N_7024);
xnor U7380 (N_7380,N_7179,N_7055);
or U7381 (N_7381,N_7072,N_7076);
nand U7382 (N_7382,N_7061,N_7152);
nor U7383 (N_7383,N_7098,N_7013);
nor U7384 (N_7384,N_7107,N_7089);
nor U7385 (N_7385,N_7141,N_7075);
nand U7386 (N_7386,N_7103,N_7153);
xnor U7387 (N_7387,N_7105,N_7010);
and U7388 (N_7388,N_7176,N_7079);
nand U7389 (N_7389,N_7080,N_7177);
xor U7390 (N_7390,N_7177,N_7078);
and U7391 (N_7391,N_7032,N_7168);
and U7392 (N_7392,N_7067,N_7047);
nand U7393 (N_7393,N_7068,N_7112);
and U7394 (N_7394,N_7067,N_7031);
nand U7395 (N_7395,N_7177,N_7021);
xor U7396 (N_7396,N_7091,N_7063);
and U7397 (N_7397,N_7183,N_7161);
or U7398 (N_7398,N_7017,N_7176);
xor U7399 (N_7399,N_7061,N_7164);
and U7400 (N_7400,N_7341,N_7271);
or U7401 (N_7401,N_7331,N_7325);
nor U7402 (N_7402,N_7311,N_7279);
xnor U7403 (N_7403,N_7301,N_7300);
or U7404 (N_7404,N_7295,N_7309);
nand U7405 (N_7405,N_7242,N_7314);
nor U7406 (N_7406,N_7231,N_7210);
nor U7407 (N_7407,N_7267,N_7332);
nor U7408 (N_7408,N_7336,N_7322);
and U7409 (N_7409,N_7282,N_7204);
or U7410 (N_7410,N_7294,N_7348);
xor U7411 (N_7411,N_7389,N_7392);
xnor U7412 (N_7412,N_7219,N_7237);
or U7413 (N_7413,N_7304,N_7258);
nand U7414 (N_7414,N_7251,N_7357);
and U7415 (N_7415,N_7216,N_7225);
nor U7416 (N_7416,N_7306,N_7288);
and U7417 (N_7417,N_7283,N_7214);
xor U7418 (N_7418,N_7256,N_7303);
and U7419 (N_7419,N_7375,N_7324);
xnor U7420 (N_7420,N_7380,N_7327);
nand U7421 (N_7421,N_7291,N_7265);
nor U7422 (N_7422,N_7373,N_7272);
nor U7423 (N_7423,N_7395,N_7248);
nand U7424 (N_7424,N_7330,N_7253);
and U7425 (N_7425,N_7293,N_7211);
nor U7426 (N_7426,N_7245,N_7270);
nand U7427 (N_7427,N_7203,N_7366);
or U7428 (N_7428,N_7218,N_7312);
and U7429 (N_7429,N_7278,N_7305);
or U7430 (N_7430,N_7257,N_7289);
and U7431 (N_7431,N_7338,N_7208);
nor U7432 (N_7432,N_7232,N_7205);
nor U7433 (N_7433,N_7223,N_7310);
and U7434 (N_7434,N_7226,N_7246);
nand U7435 (N_7435,N_7254,N_7290);
and U7436 (N_7436,N_7321,N_7388);
xnor U7437 (N_7437,N_7372,N_7234);
or U7438 (N_7438,N_7222,N_7281);
nand U7439 (N_7439,N_7264,N_7386);
nor U7440 (N_7440,N_7399,N_7284);
or U7441 (N_7441,N_7224,N_7261);
and U7442 (N_7442,N_7376,N_7356);
nor U7443 (N_7443,N_7384,N_7362);
or U7444 (N_7444,N_7221,N_7266);
and U7445 (N_7445,N_7343,N_7280);
nand U7446 (N_7446,N_7363,N_7263);
xor U7447 (N_7447,N_7398,N_7238);
nand U7448 (N_7448,N_7287,N_7274);
nor U7449 (N_7449,N_7354,N_7359);
nand U7450 (N_7450,N_7317,N_7365);
and U7451 (N_7451,N_7353,N_7259);
xor U7452 (N_7452,N_7358,N_7374);
xnor U7453 (N_7453,N_7390,N_7276);
and U7454 (N_7454,N_7334,N_7250);
nand U7455 (N_7455,N_7315,N_7367);
and U7456 (N_7456,N_7207,N_7220);
nor U7457 (N_7457,N_7342,N_7350);
nor U7458 (N_7458,N_7368,N_7240);
nand U7459 (N_7459,N_7382,N_7328);
and U7460 (N_7460,N_7233,N_7239);
and U7461 (N_7461,N_7379,N_7313);
or U7462 (N_7462,N_7377,N_7370);
xnor U7463 (N_7463,N_7255,N_7393);
nor U7464 (N_7464,N_7345,N_7308);
xor U7465 (N_7465,N_7228,N_7349);
and U7466 (N_7466,N_7262,N_7352);
or U7467 (N_7467,N_7260,N_7252);
nand U7468 (N_7468,N_7249,N_7236);
nand U7469 (N_7469,N_7206,N_7292);
and U7470 (N_7470,N_7299,N_7339);
or U7471 (N_7471,N_7302,N_7273);
nand U7472 (N_7472,N_7333,N_7200);
nand U7473 (N_7473,N_7275,N_7351);
nor U7474 (N_7474,N_7307,N_7212);
xor U7475 (N_7475,N_7241,N_7337);
nand U7476 (N_7476,N_7297,N_7201);
nand U7477 (N_7477,N_7285,N_7391);
nand U7478 (N_7478,N_7244,N_7277);
and U7479 (N_7479,N_7347,N_7316);
or U7480 (N_7480,N_7340,N_7247);
nor U7481 (N_7481,N_7355,N_7326);
xnor U7482 (N_7482,N_7298,N_7269);
xnor U7483 (N_7483,N_7383,N_7378);
nand U7484 (N_7484,N_7335,N_7235);
and U7485 (N_7485,N_7215,N_7369);
and U7486 (N_7486,N_7202,N_7329);
and U7487 (N_7487,N_7296,N_7320);
or U7488 (N_7488,N_7360,N_7344);
nor U7489 (N_7489,N_7387,N_7268);
nand U7490 (N_7490,N_7243,N_7394);
or U7491 (N_7491,N_7217,N_7364);
and U7492 (N_7492,N_7286,N_7229);
nor U7493 (N_7493,N_7396,N_7346);
nand U7494 (N_7494,N_7385,N_7227);
and U7495 (N_7495,N_7361,N_7319);
or U7496 (N_7496,N_7209,N_7397);
nor U7497 (N_7497,N_7230,N_7381);
or U7498 (N_7498,N_7323,N_7371);
xor U7499 (N_7499,N_7318,N_7213);
xnor U7500 (N_7500,N_7371,N_7256);
nor U7501 (N_7501,N_7383,N_7355);
nor U7502 (N_7502,N_7257,N_7347);
nand U7503 (N_7503,N_7208,N_7378);
xnor U7504 (N_7504,N_7382,N_7364);
xor U7505 (N_7505,N_7214,N_7396);
xor U7506 (N_7506,N_7280,N_7331);
nand U7507 (N_7507,N_7389,N_7264);
nor U7508 (N_7508,N_7256,N_7310);
nor U7509 (N_7509,N_7249,N_7210);
and U7510 (N_7510,N_7346,N_7244);
nor U7511 (N_7511,N_7388,N_7383);
xnor U7512 (N_7512,N_7312,N_7380);
nand U7513 (N_7513,N_7327,N_7384);
nand U7514 (N_7514,N_7360,N_7309);
nand U7515 (N_7515,N_7347,N_7286);
nor U7516 (N_7516,N_7302,N_7237);
nand U7517 (N_7517,N_7322,N_7337);
or U7518 (N_7518,N_7398,N_7313);
and U7519 (N_7519,N_7249,N_7228);
and U7520 (N_7520,N_7330,N_7221);
or U7521 (N_7521,N_7208,N_7359);
or U7522 (N_7522,N_7274,N_7254);
nor U7523 (N_7523,N_7373,N_7324);
and U7524 (N_7524,N_7356,N_7365);
nor U7525 (N_7525,N_7379,N_7256);
nand U7526 (N_7526,N_7212,N_7390);
and U7527 (N_7527,N_7211,N_7200);
nand U7528 (N_7528,N_7226,N_7341);
and U7529 (N_7529,N_7201,N_7354);
nand U7530 (N_7530,N_7217,N_7322);
xor U7531 (N_7531,N_7352,N_7304);
nand U7532 (N_7532,N_7258,N_7284);
nor U7533 (N_7533,N_7370,N_7330);
nor U7534 (N_7534,N_7323,N_7394);
or U7535 (N_7535,N_7226,N_7223);
nor U7536 (N_7536,N_7286,N_7335);
or U7537 (N_7537,N_7275,N_7333);
nand U7538 (N_7538,N_7314,N_7216);
and U7539 (N_7539,N_7266,N_7337);
nand U7540 (N_7540,N_7259,N_7276);
and U7541 (N_7541,N_7311,N_7307);
xnor U7542 (N_7542,N_7340,N_7368);
xnor U7543 (N_7543,N_7382,N_7363);
nand U7544 (N_7544,N_7345,N_7282);
xor U7545 (N_7545,N_7399,N_7320);
or U7546 (N_7546,N_7214,N_7326);
and U7547 (N_7547,N_7235,N_7365);
and U7548 (N_7548,N_7326,N_7303);
nand U7549 (N_7549,N_7204,N_7341);
xnor U7550 (N_7550,N_7334,N_7359);
or U7551 (N_7551,N_7201,N_7399);
nor U7552 (N_7552,N_7339,N_7328);
or U7553 (N_7553,N_7335,N_7220);
nand U7554 (N_7554,N_7390,N_7203);
or U7555 (N_7555,N_7219,N_7398);
nor U7556 (N_7556,N_7253,N_7220);
nor U7557 (N_7557,N_7398,N_7362);
nand U7558 (N_7558,N_7243,N_7315);
nand U7559 (N_7559,N_7204,N_7292);
nor U7560 (N_7560,N_7232,N_7322);
and U7561 (N_7561,N_7218,N_7281);
xor U7562 (N_7562,N_7230,N_7342);
nor U7563 (N_7563,N_7297,N_7384);
or U7564 (N_7564,N_7340,N_7332);
and U7565 (N_7565,N_7276,N_7308);
and U7566 (N_7566,N_7392,N_7227);
nand U7567 (N_7567,N_7308,N_7233);
or U7568 (N_7568,N_7314,N_7275);
xor U7569 (N_7569,N_7358,N_7314);
nand U7570 (N_7570,N_7322,N_7249);
nor U7571 (N_7571,N_7346,N_7392);
and U7572 (N_7572,N_7345,N_7235);
nor U7573 (N_7573,N_7341,N_7246);
xnor U7574 (N_7574,N_7238,N_7203);
or U7575 (N_7575,N_7286,N_7250);
and U7576 (N_7576,N_7304,N_7288);
and U7577 (N_7577,N_7253,N_7289);
or U7578 (N_7578,N_7286,N_7231);
xnor U7579 (N_7579,N_7224,N_7354);
and U7580 (N_7580,N_7268,N_7238);
xor U7581 (N_7581,N_7383,N_7203);
and U7582 (N_7582,N_7272,N_7233);
and U7583 (N_7583,N_7365,N_7240);
xnor U7584 (N_7584,N_7210,N_7357);
and U7585 (N_7585,N_7294,N_7370);
xnor U7586 (N_7586,N_7360,N_7341);
or U7587 (N_7587,N_7343,N_7325);
nor U7588 (N_7588,N_7207,N_7331);
nand U7589 (N_7589,N_7247,N_7255);
or U7590 (N_7590,N_7384,N_7213);
nand U7591 (N_7591,N_7242,N_7247);
or U7592 (N_7592,N_7260,N_7321);
nor U7593 (N_7593,N_7390,N_7375);
and U7594 (N_7594,N_7248,N_7286);
nand U7595 (N_7595,N_7344,N_7295);
or U7596 (N_7596,N_7365,N_7263);
and U7597 (N_7597,N_7249,N_7272);
xor U7598 (N_7598,N_7375,N_7229);
or U7599 (N_7599,N_7318,N_7214);
and U7600 (N_7600,N_7491,N_7474);
nand U7601 (N_7601,N_7576,N_7403);
xor U7602 (N_7602,N_7481,N_7581);
and U7603 (N_7603,N_7456,N_7484);
or U7604 (N_7604,N_7473,N_7565);
or U7605 (N_7605,N_7503,N_7404);
xor U7606 (N_7606,N_7550,N_7502);
nand U7607 (N_7607,N_7477,N_7422);
nor U7608 (N_7608,N_7588,N_7500);
xor U7609 (N_7609,N_7419,N_7570);
nand U7610 (N_7610,N_7489,N_7505);
nor U7611 (N_7611,N_7467,N_7430);
and U7612 (N_7612,N_7447,N_7480);
nand U7613 (N_7613,N_7584,N_7560);
nand U7614 (N_7614,N_7461,N_7439);
and U7615 (N_7615,N_7498,N_7518);
nor U7616 (N_7616,N_7425,N_7548);
and U7617 (N_7617,N_7412,N_7547);
or U7618 (N_7618,N_7415,N_7408);
and U7619 (N_7619,N_7564,N_7438);
nand U7620 (N_7620,N_7558,N_7431);
or U7621 (N_7621,N_7520,N_7407);
or U7622 (N_7622,N_7435,N_7492);
and U7623 (N_7623,N_7544,N_7437);
xnor U7624 (N_7624,N_7551,N_7554);
nand U7625 (N_7625,N_7524,N_7434);
nor U7626 (N_7626,N_7442,N_7531);
nor U7627 (N_7627,N_7469,N_7496);
xor U7628 (N_7628,N_7466,N_7450);
nand U7629 (N_7629,N_7413,N_7596);
nand U7630 (N_7630,N_7427,N_7420);
nand U7631 (N_7631,N_7533,N_7455);
or U7632 (N_7632,N_7465,N_7487);
or U7633 (N_7633,N_7532,N_7510);
xor U7634 (N_7634,N_7515,N_7457);
or U7635 (N_7635,N_7525,N_7433);
or U7636 (N_7636,N_7535,N_7471);
nand U7637 (N_7637,N_7569,N_7538);
xor U7638 (N_7638,N_7589,N_7566);
nand U7639 (N_7639,N_7598,N_7472);
nor U7640 (N_7640,N_7454,N_7509);
nand U7641 (N_7641,N_7562,N_7542);
xnor U7642 (N_7642,N_7462,N_7468);
or U7643 (N_7643,N_7426,N_7536);
or U7644 (N_7644,N_7414,N_7549);
xor U7645 (N_7645,N_7561,N_7572);
or U7646 (N_7646,N_7527,N_7599);
nor U7647 (N_7647,N_7546,N_7580);
xnor U7648 (N_7648,N_7406,N_7514);
nand U7649 (N_7649,N_7488,N_7446);
nor U7650 (N_7650,N_7543,N_7522);
nand U7651 (N_7651,N_7410,N_7553);
or U7652 (N_7652,N_7539,N_7423);
and U7653 (N_7653,N_7575,N_7523);
and U7654 (N_7654,N_7595,N_7464);
nand U7655 (N_7655,N_7594,N_7541);
and U7656 (N_7656,N_7499,N_7511);
or U7657 (N_7657,N_7490,N_7555);
or U7658 (N_7658,N_7453,N_7585);
xor U7659 (N_7659,N_7530,N_7578);
or U7660 (N_7660,N_7459,N_7516);
nand U7661 (N_7661,N_7440,N_7537);
and U7662 (N_7662,N_7495,N_7592);
nand U7663 (N_7663,N_7497,N_7521);
or U7664 (N_7664,N_7483,N_7421);
or U7665 (N_7665,N_7448,N_7476);
xor U7666 (N_7666,N_7441,N_7571);
or U7667 (N_7667,N_7409,N_7429);
or U7668 (N_7668,N_7526,N_7485);
nand U7669 (N_7669,N_7597,N_7479);
and U7670 (N_7670,N_7445,N_7436);
and U7671 (N_7671,N_7577,N_7573);
xnor U7672 (N_7672,N_7556,N_7540);
nand U7673 (N_7673,N_7557,N_7458);
nor U7674 (N_7674,N_7583,N_7418);
or U7675 (N_7675,N_7493,N_7451);
and U7676 (N_7676,N_7432,N_7587);
xor U7677 (N_7677,N_7563,N_7482);
nor U7678 (N_7678,N_7545,N_7519);
nor U7679 (N_7679,N_7528,N_7529);
nor U7680 (N_7680,N_7486,N_7416);
nand U7681 (N_7681,N_7579,N_7517);
nand U7682 (N_7682,N_7494,N_7475);
nor U7683 (N_7683,N_7504,N_7400);
or U7684 (N_7684,N_7449,N_7508);
xnor U7685 (N_7685,N_7513,N_7501);
or U7686 (N_7686,N_7506,N_7591);
and U7687 (N_7687,N_7402,N_7401);
nor U7688 (N_7688,N_7586,N_7463);
nor U7689 (N_7689,N_7534,N_7428);
or U7690 (N_7690,N_7567,N_7568);
or U7691 (N_7691,N_7559,N_7444);
xnor U7692 (N_7692,N_7460,N_7405);
and U7693 (N_7693,N_7452,N_7478);
nor U7694 (N_7694,N_7552,N_7411);
and U7695 (N_7695,N_7590,N_7417);
nand U7696 (N_7696,N_7424,N_7470);
xnor U7697 (N_7697,N_7507,N_7443);
or U7698 (N_7698,N_7574,N_7582);
xnor U7699 (N_7699,N_7512,N_7593);
or U7700 (N_7700,N_7506,N_7586);
and U7701 (N_7701,N_7530,N_7466);
nor U7702 (N_7702,N_7594,N_7524);
xor U7703 (N_7703,N_7550,N_7463);
or U7704 (N_7704,N_7558,N_7472);
or U7705 (N_7705,N_7561,N_7549);
and U7706 (N_7706,N_7423,N_7556);
nand U7707 (N_7707,N_7510,N_7437);
nor U7708 (N_7708,N_7562,N_7553);
nor U7709 (N_7709,N_7482,N_7593);
xor U7710 (N_7710,N_7475,N_7429);
xor U7711 (N_7711,N_7575,N_7447);
xnor U7712 (N_7712,N_7516,N_7527);
or U7713 (N_7713,N_7423,N_7424);
nor U7714 (N_7714,N_7515,N_7409);
and U7715 (N_7715,N_7471,N_7556);
and U7716 (N_7716,N_7473,N_7408);
or U7717 (N_7717,N_7402,N_7560);
nand U7718 (N_7718,N_7482,N_7541);
nand U7719 (N_7719,N_7463,N_7556);
nor U7720 (N_7720,N_7447,N_7432);
nor U7721 (N_7721,N_7417,N_7497);
nand U7722 (N_7722,N_7473,N_7433);
and U7723 (N_7723,N_7446,N_7554);
xor U7724 (N_7724,N_7558,N_7405);
nand U7725 (N_7725,N_7456,N_7535);
xor U7726 (N_7726,N_7514,N_7456);
nand U7727 (N_7727,N_7450,N_7516);
and U7728 (N_7728,N_7493,N_7534);
nand U7729 (N_7729,N_7491,N_7592);
nor U7730 (N_7730,N_7426,N_7597);
or U7731 (N_7731,N_7582,N_7405);
nor U7732 (N_7732,N_7593,N_7584);
xor U7733 (N_7733,N_7571,N_7533);
and U7734 (N_7734,N_7471,N_7530);
nand U7735 (N_7735,N_7428,N_7495);
nand U7736 (N_7736,N_7559,N_7504);
and U7737 (N_7737,N_7588,N_7515);
xnor U7738 (N_7738,N_7472,N_7574);
xor U7739 (N_7739,N_7415,N_7495);
and U7740 (N_7740,N_7445,N_7444);
nor U7741 (N_7741,N_7446,N_7467);
or U7742 (N_7742,N_7482,N_7515);
xnor U7743 (N_7743,N_7401,N_7547);
nor U7744 (N_7744,N_7553,N_7431);
or U7745 (N_7745,N_7499,N_7484);
or U7746 (N_7746,N_7468,N_7582);
nor U7747 (N_7747,N_7534,N_7510);
or U7748 (N_7748,N_7567,N_7507);
xor U7749 (N_7749,N_7586,N_7496);
and U7750 (N_7750,N_7562,N_7447);
nand U7751 (N_7751,N_7512,N_7566);
nor U7752 (N_7752,N_7420,N_7527);
nand U7753 (N_7753,N_7496,N_7571);
and U7754 (N_7754,N_7423,N_7518);
nor U7755 (N_7755,N_7501,N_7418);
and U7756 (N_7756,N_7405,N_7509);
nor U7757 (N_7757,N_7432,N_7475);
nor U7758 (N_7758,N_7526,N_7553);
xnor U7759 (N_7759,N_7472,N_7473);
and U7760 (N_7760,N_7407,N_7570);
and U7761 (N_7761,N_7572,N_7413);
or U7762 (N_7762,N_7571,N_7457);
or U7763 (N_7763,N_7428,N_7431);
nor U7764 (N_7764,N_7481,N_7400);
xnor U7765 (N_7765,N_7425,N_7576);
xor U7766 (N_7766,N_7566,N_7508);
nor U7767 (N_7767,N_7555,N_7471);
or U7768 (N_7768,N_7535,N_7566);
nor U7769 (N_7769,N_7405,N_7583);
xnor U7770 (N_7770,N_7574,N_7597);
xnor U7771 (N_7771,N_7403,N_7532);
nor U7772 (N_7772,N_7578,N_7541);
xor U7773 (N_7773,N_7534,N_7576);
and U7774 (N_7774,N_7453,N_7455);
or U7775 (N_7775,N_7501,N_7423);
or U7776 (N_7776,N_7492,N_7466);
nor U7777 (N_7777,N_7451,N_7517);
nand U7778 (N_7778,N_7493,N_7465);
xor U7779 (N_7779,N_7427,N_7517);
nor U7780 (N_7780,N_7590,N_7552);
nor U7781 (N_7781,N_7438,N_7514);
nor U7782 (N_7782,N_7565,N_7517);
xor U7783 (N_7783,N_7456,N_7496);
or U7784 (N_7784,N_7588,N_7446);
nand U7785 (N_7785,N_7438,N_7408);
nor U7786 (N_7786,N_7504,N_7456);
or U7787 (N_7787,N_7433,N_7526);
nand U7788 (N_7788,N_7573,N_7563);
xor U7789 (N_7789,N_7502,N_7596);
nor U7790 (N_7790,N_7443,N_7442);
and U7791 (N_7791,N_7561,N_7535);
or U7792 (N_7792,N_7538,N_7530);
xnor U7793 (N_7793,N_7485,N_7568);
nand U7794 (N_7794,N_7564,N_7403);
and U7795 (N_7795,N_7571,N_7520);
nand U7796 (N_7796,N_7552,N_7481);
nand U7797 (N_7797,N_7520,N_7495);
nor U7798 (N_7798,N_7440,N_7459);
or U7799 (N_7799,N_7462,N_7452);
and U7800 (N_7800,N_7779,N_7638);
nand U7801 (N_7801,N_7767,N_7694);
nor U7802 (N_7802,N_7662,N_7736);
and U7803 (N_7803,N_7785,N_7697);
nand U7804 (N_7804,N_7787,N_7602);
and U7805 (N_7805,N_7632,N_7668);
xor U7806 (N_7806,N_7795,N_7761);
and U7807 (N_7807,N_7728,N_7763);
nor U7808 (N_7808,N_7745,N_7760);
nor U7809 (N_7809,N_7670,N_7611);
nand U7810 (N_7810,N_7714,N_7724);
and U7811 (N_7811,N_7713,N_7790);
xor U7812 (N_7812,N_7727,N_7667);
and U7813 (N_7813,N_7762,N_7609);
xnor U7814 (N_7814,N_7721,N_7684);
nand U7815 (N_7815,N_7748,N_7679);
nor U7816 (N_7816,N_7676,N_7650);
or U7817 (N_7817,N_7648,N_7620);
xor U7818 (N_7818,N_7606,N_7778);
xor U7819 (N_7819,N_7643,N_7675);
nand U7820 (N_7820,N_7665,N_7765);
nor U7821 (N_7821,N_7616,N_7623);
xor U7822 (N_7822,N_7604,N_7744);
nand U7823 (N_7823,N_7674,N_7749);
or U7824 (N_7824,N_7772,N_7708);
and U7825 (N_7825,N_7738,N_7746);
nor U7826 (N_7826,N_7773,N_7726);
nor U7827 (N_7827,N_7678,N_7758);
nand U7828 (N_7828,N_7686,N_7711);
or U7829 (N_7829,N_7729,N_7751);
nand U7830 (N_7830,N_7631,N_7653);
nand U7831 (N_7831,N_7698,N_7725);
nor U7832 (N_7832,N_7747,N_7699);
nand U7833 (N_7833,N_7797,N_7630);
nand U7834 (N_7834,N_7644,N_7703);
and U7835 (N_7835,N_7659,N_7757);
and U7836 (N_7836,N_7622,N_7646);
or U7837 (N_7837,N_7601,N_7640);
xor U7838 (N_7838,N_7704,N_7723);
or U7839 (N_7839,N_7691,N_7682);
nand U7840 (N_7840,N_7782,N_7756);
nor U7841 (N_7841,N_7702,N_7783);
nand U7842 (N_7842,N_7781,N_7759);
or U7843 (N_7843,N_7656,N_7605);
xor U7844 (N_7844,N_7712,N_7755);
and U7845 (N_7845,N_7626,N_7799);
nor U7846 (N_7846,N_7780,N_7617);
nor U7847 (N_7847,N_7798,N_7775);
nand U7848 (N_7848,N_7701,N_7695);
nand U7849 (N_7849,N_7614,N_7625);
xor U7850 (N_7850,N_7651,N_7716);
and U7851 (N_7851,N_7705,N_7658);
nor U7852 (N_7852,N_7720,N_7776);
or U7853 (N_7853,N_7685,N_7673);
xnor U7854 (N_7854,N_7693,N_7608);
or U7855 (N_7855,N_7717,N_7731);
xor U7856 (N_7856,N_7766,N_7734);
nor U7857 (N_7857,N_7769,N_7770);
nor U7858 (N_7858,N_7664,N_7796);
or U7859 (N_7859,N_7603,N_7621);
xnor U7860 (N_7860,N_7610,N_7791);
and U7861 (N_7861,N_7635,N_7661);
and U7862 (N_7862,N_7788,N_7777);
or U7863 (N_7863,N_7737,N_7672);
and U7864 (N_7864,N_7690,N_7652);
and U7865 (N_7865,N_7794,N_7612);
and U7866 (N_7866,N_7774,N_7677);
and U7867 (N_7867,N_7750,N_7634);
xor U7868 (N_7868,N_7666,N_7733);
nand U7869 (N_7869,N_7793,N_7636);
xor U7870 (N_7870,N_7771,N_7706);
xor U7871 (N_7871,N_7742,N_7789);
or U7872 (N_7872,N_7683,N_7655);
xnor U7873 (N_7873,N_7740,N_7639);
nor U7874 (N_7874,N_7764,N_7752);
xnor U7875 (N_7875,N_7669,N_7730);
or U7876 (N_7876,N_7619,N_7600);
nor U7877 (N_7877,N_7645,N_7687);
nor U7878 (N_7878,N_7657,N_7613);
nor U7879 (N_7879,N_7753,N_7784);
nand U7880 (N_7880,N_7642,N_7719);
or U7881 (N_7881,N_7722,N_7792);
or U7882 (N_7882,N_7707,N_7688);
xor U7883 (N_7883,N_7629,N_7607);
nor U7884 (N_7884,N_7692,N_7633);
nand U7885 (N_7885,N_7689,N_7739);
or U7886 (N_7886,N_7627,N_7768);
or U7887 (N_7887,N_7654,N_7660);
nand U7888 (N_7888,N_7637,N_7735);
and U7889 (N_7889,N_7743,N_7709);
nand U7890 (N_7890,N_7624,N_7615);
and U7891 (N_7891,N_7649,N_7700);
nand U7892 (N_7892,N_7647,N_7681);
and U7893 (N_7893,N_7628,N_7715);
xnor U7894 (N_7894,N_7671,N_7754);
xor U7895 (N_7895,N_7732,N_7786);
nand U7896 (N_7896,N_7710,N_7663);
nor U7897 (N_7897,N_7641,N_7741);
nor U7898 (N_7898,N_7680,N_7696);
xnor U7899 (N_7899,N_7618,N_7718);
nor U7900 (N_7900,N_7643,N_7752);
and U7901 (N_7901,N_7700,N_7740);
and U7902 (N_7902,N_7608,N_7641);
and U7903 (N_7903,N_7666,N_7637);
or U7904 (N_7904,N_7622,N_7638);
xor U7905 (N_7905,N_7764,N_7771);
xnor U7906 (N_7906,N_7797,N_7660);
nor U7907 (N_7907,N_7656,N_7615);
and U7908 (N_7908,N_7619,N_7738);
or U7909 (N_7909,N_7746,N_7745);
xor U7910 (N_7910,N_7719,N_7793);
xnor U7911 (N_7911,N_7724,N_7785);
nand U7912 (N_7912,N_7621,N_7716);
or U7913 (N_7913,N_7620,N_7605);
and U7914 (N_7914,N_7758,N_7609);
nand U7915 (N_7915,N_7795,N_7738);
nor U7916 (N_7916,N_7662,N_7634);
xor U7917 (N_7917,N_7748,N_7666);
and U7918 (N_7918,N_7671,N_7769);
nor U7919 (N_7919,N_7614,N_7715);
or U7920 (N_7920,N_7617,N_7649);
xor U7921 (N_7921,N_7610,N_7790);
or U7922 (N_7922,N_7640,N_7617);
and U7923 (N_7923,N_7681,N_7653);
and U7924 (N_7924,N_7659,N_7780);
nand U7925 (N_7925,N_7655,N_7796);
nor U7926 (N_7926,N_7623,N_7601);
or U7927 (N_7927,N_7645,N_7721);
xnor U7928 (N_7928,N_7739,N_7633);
nand U7929 (N_7929,N_7682,N_7667);
nor U7930 (N_7930,N_7642,N_7788);
xnor U7931 (N_7931,N_7798,N_7637);
or U7932 (N_7932,N_7638,N_7796);
and U7933 (N_7933,N_7711,N_7698);
xor U7934 (N_7934,N_7643,N_7770);
or U7935 (N_7935,N_7705,N_7792);
or U7936 (N_7936,N_7735,N_7746);
and U7937 (N_7937,N_7773,N_7720);
and U7938 (N_7938,N_7721,N_7739);
xnor U7939 (N_7939,N_7718,N_7712);
nor U7940 (N_7940,N_7664,N_7770);
nor U7941 (N_7941,N_7625,N_7645);
nand U7942 (N_7942,N_7735,N_7700);
and U7943 (N_7943,N_7778,N_7637);
xor U7944 (N_7944,N_7630,N_7757);
xor U7945 (N_7945,N_7616,N_7741);
nor U7946 (N_7946,N_7660,N_7679);
nor U7947 (N_7947,N_7685,N_7631);
xnor U7948 (N_7948,N_7719,N_7694);
nand U7949 (N_7949,N_7777,N_7688);
or U7950 (N_7950,N_7647,N_7699);
nor U7951 (N_7951,N_7689,N_7717);
nor U7952 (N_7952,N_7728,N_7761);
and U7953 (N_7953,N_7743,N_7648);
nand U7954 (N_7954,N_7718,N_7723);
xor U7955 (N_7955,N_7679,N_7774);
or U7956 (N_7956,N_7762,N_7661);
xor U7957 (N_7957,N_7707,N_7681);
and U7958 (N_7958,N_7791,N_7602);
or U7959 (N_7959,N_7794,N_7622);
nor U7960 (N_7960,N_7780,N_7642);
and U7961 (N_7961,N_7764,N_7615);
nor U7962 (N_7962,N_7721,N_7669);
nand U7963 (N_7963,N_7764,N_7788);
and U7964 (N_7964,N_7607,N_7762);
or U7965 (N_7965,N_7740,N_7694);
nand U7966 (N_7966,N_7638,N_7688);
nor U7967 (N_7967,N_7762,N_7646);
xor U7968 (N_7968,N_7698,N_7672);
nand U7969 (N_7969,N_7663,N_7605);
nor U7970 (N_7970,N_7768,N_7672);
xor U7971 (N_7971,N_7643,N_7648);
nand U7972 (N_7972,N_7744,N_7714);
nand U7973 (N_7973,N_7707,N_7662);
or U7974 (N_7974,N_7764,N_7664);
or U7975 (N_7975,N_7691,N_7636);
and U7976 (N_7976,N_7613,N_7767);
and U7977 (N_7977,N_7744,N_7673);
or U7978 (N_7978,N_7712,N_7744);
xor U7979 (N_7979,N_7690,N_7753);
and U7980 (N_7980,N_7766,N_7717);
nor U7981 (N_7981,N_7740,N_7776);
or U7982 (N_7982,N_7677,N_7648);
nand U7983 (N_7983,N_7663,N_7742);
and U7984 (N_7984,N_7608,N_7765);
nor U7985 (N_7985,N_7709,N_7694);
and U7986 (N_7986,N_7790,N_7669);
or U7987 (N_7987,N_7670,N_7681);
and U7988 (N_7988,N_7761,N_7781);
nand U7989 (N_7989,N_7769,N_7688);
nand U7990 (N_7990,N_7699,N_7633);
or U7991 (N_7991,N_7750,N_7719);
and U7992 (N_7992,N_7763,N_7714);
and U7993 (N_7993,N_7697,N_7668);
and U7994 (N_7994,N_7747,N_7612);
xor U7995 (N_7995,N_7723,N_7627);
and U7996 (N_7996,N_7747,N_7623);
xnor U7997 (N_7997,N_7702,N_7780);
nor U7998 (N_7998,N_7615,N_7797);
and U7999 (N_7999,N_7628,N_7619);
or U8000 (N_8000,N_7845,N_7809);
nand U8001 (N_8001,N_7872,N_7918);
or U8002 (N_8002,N_7905,N_7936);
and U8003 (N_8003,N_7839,N_7893);
and U8004 (N_8004,N_7824,N_7900);
nor U8005 (N_8005,N_7883,N_7841);
or U8006 (N_8006,N_7982,N_7899);
nand U8007 (N_8007,N_7870,N_7993);
nand U8008 (N_8008,N_7821,N_7980);
nor U8009 (N_8009,N_7838,N_7862);
nand U8010 (N_8010,N_7814,N_7922);
xnor U8011 (N_8011,N_7969,N_7871);
or U8012 (N_8012,N_7805,N_7984);
xor U8013 (N_8013,N_7853,N_7807);
nor U8014 (N_8014,N_7926,N_7965);
or U8015 (N_8015,N_7825,N_7929);
nand U8016 (N_8016,N_7834,N_7874);
xor U8017 (N_8017,N_7860,N_7806);
or U8018 (N_8018,N_7995,N_7920);
xnor U8019 (N_8019,N_7950,N_7810);
nand U8020 (N_8020,N_7844,N_7878);
xnor U8021 (N_8021,N_7815,N_7849);
and U8022 (N_8022,N_7879,N_7817);
nor U8023 (N_8023,N_7831,N_7949);
nor U8024 (N_8024,N_7962,N_7867);
or U8025 (N_8025,N_7912,N_7863);
nor U8026 (N_8026,N_7803,N_7859);
nand U8027 (N_8027,N_7868,N_7966);
and U8028 (N_8028,N_7819,N_7985);
nor U8029 (N_8029,N_7943,N_7895);
nand U8030 (N_8030,N_7861,N_7972);
nand U8031 (N_8031,N_7932,N_7818);
or U8032 (N_8032,N_7945,N_7832);
or U8033 (N_8033,N_7935,N_7842);
nand U8034 (N_8034,N_7963,N_7873);
or U8035 (N_8035,N_7992,N_7971);
nand U8036 (N_8036,N_7991,N_7858);
xor U8037 (N_8037,N_7916,N_7908);
nand U8038 (N_8038,N_7811,N_7975);
nand U8039 (N_8039,N_7856,N_7970);
and U8040 (N_8040,N_7958,N_7989);
and U8041 (N_8041,N_7851,N_7829);
or U8042 (N_8042,N_7813,N_7956);
nor U8043 (N_8043,N_7892,N_7865);
nor U8044 (N_8044,N_7830,N_7974);
nor U8045 (N_8045,N_7919,N_7968);
and U8046 (N_8046,N_7977,N_7875);
and U8047 (N_8047,N_7979,N_7959);
nor U8048 (N_8048,N_7801,N_7934);
or U8049 (N_8049,N_7957,N_7927);
or U8050 (N_8050,N_7826,N_7915);
or U8051 (N_8051,N_7903,N_7850);
and U8052 (N_8052,N_7976,N_7928);
xor U8053 (N_8053,N_7930,N_7866);
nand U8054 (N_8054,N_7973,N_7944);
or U8055 (N_8055,N_7907,N_7906);
nor U8056 (N_8056,N_7931,N_7960);
nand U8057 (N_8057,N_7887,N_7828);
xnor U8058 (N_8058,N_7967,N_7852);
nor U8059 (N_8059,N_7843,N_7951);
nor U8060 (N_8060,N_7802,N_7888);
and U8061 (N_8061,N_7964,N_7990);
and U8062 (N_8062,N_7880,N_7983);
or U8063 (N_8063,N_7836,N_7835);
xor U8064 (N_8064,N_7896,N_7808);
xnor U8065 (N_8065,N_7885,N_7877);
or U8066 (N_8066,N_7864,N_7946);
xor U8067 (N_8067,N_7952,N_7996);
nand U8068 (N_8068,N_7981,N_7882);
or U8069 (N_8069,N_7997,N_7933);
or U8070 (N_8070,N_7823,N_7820);
xor U8071 (N_8071,N_7816,N_7942);
or U8072 (N_8072,N_7999,N_7855);
or U8073 (N_8073,N_7869,N_7847);
nand U8074 (N_8074,N_7938,N_7901);
xnor U8075 (N_8075,N_7917,N_7904);
and U8076 (N_8076,N_7948,N_7857);
or U8077 (N_8077,N_7827,N_7881);
xnor U8078 (N_8078,N_7955,N_7889);
and U8079 (N_8079,N_7840,N_7954);
or U8080 (N_8080,N_7848,N_7924);
xor U8081 (N_8081,N_7898,N_7961);
and U8082 (N_8082,N_7902,N_7921);
or U8083 (N_8083,N_7876,N_7994);
nand U8084 (N_8084,N_7998,N_7854);
or U8085 (N_8085,N_7822,N_7884);
or U8086 (N_8086,N_7846,N_7953);
xnor U8087 (N_8087,N_7886,N_7940);
and U8088 (N_8088,N_7833,N_7986);
and U8089 (N_8089,N_7800,N_7913);
xnor U8090 (N_8090,N_7812,N_7941);
nor U8091 (N_8091,N_7891,N_7987);
nor U8092 (N_8092,N_7937,N_7923);
nand U8093 (N_8093,N_7894,N_7978);
nor U8094 (N_8094,N_7804,N_7947);
nand U8095 (N_8095,N_7909,N_7890);
or U8096 (N_8096,N_7925,N_7837);
nor U8097 (N_8097,N_7897,N_7910);
and U8098 (N_8098,N_7939,N_7988);
nand U8099 (N_8099,N_7914,N_7911);
or U8100 (N_8100,N_7964,N_7947);
xor U8101 (N_8101,N_7933,N_7848);
or U8102 (N_8102,N_7859,N_7923);
nand U8103 (N_8103,N_7883,N_7866);
or U8104 (N_8104,N_7924,N_7956);
nand U8105 (N_8105,N_7857,N_7848);
xnor U8106 (N_8106,N_7985,N_7883);
xor U8107 (N_8107,N_7903,N_7837);
xnor U8108 (N_8108,N_7915,N_7905);
and U8109 (N_8109,N_7806,N_7972);
nor U8110 (N_8110,N_7942,N_7823);
nor U8111 (N_8111,N_7852,N_7987);
nand U8112 (N_8112,N_7910,N_7868);
nand U8113 (N_8113,N_7881,N_7979);
or U8114 (N_8114,N_7811,N_7832);
or U8115 (N_8115,N_7945,N_7948);
nand U8116 (N_8116,N_7941,N_7863);
nand U8117 (N_8117,N_7855,N_7899);
and U8118 (N_8118,N_7800,N_7851);
nand U8119 (N_8119,N_7844,N_7976);
nor U8120 (N_8120,N_7908,N_7815);
xnor U8121 (N_8121,N_7902,N_7997);
xnor U8122 (N_8122,N_7967,N_7903);
xor U8123 (N_8123,N_7944,N_7963);
or U8124 (N_8124,N_7981,N_7919);
xnor U8125 (N_8125,N_7847,N_7928);
or U8126 (N_8126,N_7838,N_7966);
xnor U8127 (N_8127,N_7933,N_7926);
xor U8128 (N_8128,N_7974,N_7914);
xor U8129 (N_8129,N_7841,N_7936);
nor U8130 (N_8130,N_7969,N_7856);
and U8131 (N_8131,N_7990,N_7986);
xnor U8132 (N_8132,N_7887,N_7946);
and U8133 (N_8133,N_7874,N_7898);
xor U8134 (N_8134,N_7853,N_7856);
nand U8135 (N_8135,N_7854,N_7944);
and U8136 (N_8136,N_7887,N_7938);
and U8137 (N_8137,N_7971,N_7955);
nand U8138 (N_8138,N_7961,N_7976);
xnor U8139 (N_8139,N_7891,N_7831);
nor U8140 (N_8140,N_7918,N_7807);
and U8141 (N_8141,N_7837,N_7979);
or U8142 (N_8142,N_7843,N_7815);
nor U8143 (N_8143,N_7831,N_7942);
or U8144 (N_8144,N_7913,N_7864);
and U8145 (N_8145,N_7869,N_7968);
xnor U8146 (N_8146,N_7880,N_7912);
nor U8147 (N_8147,N_7986,N_7885);
xor U8148 (N_8148,N_7965,N_7817);
nand U8149 (N_8149,N_7808,N_7844);
xnor U8150 (N_8150,N_7990,N_7852);
nor U8151 (N_8151,N_7902,N_7917);
nor U8152 (N_8152,N_7950,N_7836);
nor U8153 (N_8153,N_7890,N_7815);
nand U8154 (N_8154,N_7906,N_7836);
and U8155 (N_8155,N_7898,N_7832);
xnor U8156 (N_8156,N_7802,N_7863);
or U8157 (N_8157,N_7857,N_7861);
xnor U8158 (N_8158,N_7946,N_7838);
or U8159 (N_8159,N_7937,N_7883);
xnor U8160 (N_8160,N_7831,N_7972);
nand U8161 (N_8161,N_7951,N_7882);
and U8162 (N_8162,N_7844,N_7963);
nor U8163 (N_8163,N_7912,N_7808);
xor U8164 (N_8164,N_7916,N_7918);
nor U8165 (N_8165,N_7926,N_7954);
nand U8166 (N_8166,N_7898,N_7881);
nand U8167 (N_8167,N_7906,N_7892);
xor U8168 (N_8168,N_7841,N_7975);
and U8169 (N_8169,N_7964,N_7817);
and U8170 (N_8170,N_7843,N_7908);
xor U8171 (N_8171,N_7834,N_7825);
xor U8172 (N_8172,N_7950,N_7939);
nor U8173 (N_8173,N_7929,N_7810);
nor U8174 (N_8174,N_7915,N_7958);
nand U8175 (N_8175,N_7923,N_7808);
and U8176 (N_8176,N_7894,N_7843);
and U8177 (N_8177,N_7895,N_7921);
nand U8178 (N_8178,N_7865,N_7904);
nor U8179 (N_8179,N_7809,N_7932);
xor U8180 (N_8180,N_7880,N_7943);
and U8181 (N_8181,N_7800,N_7877);
and U8182 (N_8182,N_7828,N_7809);
xor U8183 (N_8183,N_7878,N_7895);
and U8184 (N_8184,N_7920,N_7914);
and U8185 (N_8185,N_7898,N_7947);
nand U8186 (N_8186,N_7830,N_7997);
and U8187 (N_8187,N_7913,N_7906);
and U8188 (N_8188,N_7802,N_7920);
xor U8189 (N_8189,N_7916,N_7889);
xor U8190 (N_8190,N_7956,N_7892);
or U8191 (N_8191,N_7886,N_7919);
and U8192 (N_8192,N_7827,N_7922);
nor U8193 (N_8193,N_7909,N_7959);
or U8194 (N_8194,N_7872,N_7820);
or U8195 (N_8195,N_7875,N_7963);
nand U8196 (N_8196,N_7962,N_7990);
and U8197 (N_8197,N_7818,N_7958);
nor U8198 (N_8198,N_7880,N_7889);
xor U8199 (N_8199,N_7968,N_7959);
nand U8200 (N_8200,N_8197,N_8118);
nor U8201 (N_8201,N_8148,N_8108);
nor U8202 (N_8202,N_8101,N_8135);
nand U8203 (N_8203,N_8151,N_8027);
or U8204 (N_8204,N_8089,N_8165);
or U8205 (N_8205,N_8069,N_8053);
xnor U8206 (N_8206,N_8061,N_8037);
nand U8207 (N_8207,N_8103,N_8100);
nor U8208 (N_8208,N_8075,N_8087);
xor U8209 (N_8209,N_8175,N_8187);
nor U8210 (N_8210,N_8147,N_8133);
and U8211 (N_8211,N_8048,N_8038);
nor U8212 (N_8212,N_8000,N_8113);
and U8213 (N_8213,N_8097,N_8042);
nor U8214 (N_8214,N_8188,N_8153);
nand U8215 (N_8215,N_8039,N_8119);
or U8216 (N_8216,N_8074,N_8049);
nor U8217 (N_8217,N_8025,N_8009);
and U8218 (N_8218,N_8137,N_8046);
xnor U8219 (N_8219,N_8082,N_8195);
nor U8220 (N_8220,N_8043,N_8160);
nor U8221 (N_8221,N_8007,N_8057);
xnor U8222 (N_8222,N_8115,N_8117);
or U8223 (N_8223,N_8124,N_8077);
nor U8224 (N_8224,N_8081,N_8098);
or U8225 (N_8225,N_8020,N_8092);
nand U8226 (N_8226,N_8062,N_8141);
or U8227 (N_8227,N_8123,N_8035);
xor U8228 (N_8228,N_8126,N_8186);
nand U8229 (N_8229,N_8033,N_8159);
and U8230 (N_8230,N_8105,N_8199);
or U8231 (N_8231,N_8162,N_8182);
or U8232 (N_8232,N_8173,N_8129);
nand U8233 (N_8233,N_8060,N_8152);
and U8234 (N_8234,N_8122,N_8116);
and U8235 (N_8235,N_8161,N_8189);
nor U8236 (N_8236,N_8176,N_8030);
and U8237 (N_8237,N_8104,N_8168);
and U8238 (N_8238,N_8073,N_8149);
nor U8239 (N_8239,N_8095,N_8180);
nand U8240 (N_8240,N_8093,N_8070);
nor U8241 (N_8241,N_8001,N_8065);
xnor U8242 (N_8242,N_8066,N_8196);
or U8243 (N_8243,N_8004,N_8078);
and U8244 (N_8244,N_8181,N_8112);
nand U8245 (N_8245,N_8170,N_8138);
nor U8246 (N_8246,N_8174,N_8067);
nand U8247 (N_8247,N_8084,N_8080);
and U8248 (N_8248,N_8127,N_8008);
or U8249 (N_8249,N_8079,N_8094);
and U8250 (N_8250,N_8088,N_8010);
nand U8251 (N_8251,N_8017,N_8169);
or U8252 (N_8252,N_8006,N_8085);
or U8253 (N_8253,N_8091,N_8155);
or U8254 (N_8254,N_8194,N_8096);
and U8255 (N_8255,N_8106,N_8072);
nand U8256 (N_8256,N_8058,N_8090);
or U8257 (N_8257,N_8055,N_8011);
nor U8258 (N_8258,N_8032,N_8034);
nor U8259 (N_8259,N_8190,N_8052);
nor U8260 (N_8260,N_8036,N_8191);
xnor U8261 (N_8261,N_8198,N_8158);
xnor U8262 (N_8262,N_8145,N_8193);
and U8263 (N_8263,N_8045,N_8192);
and U8264 (N_8264,N_8177,N_8156);
nor U8265 (N_8265,N_8121,N_8056);
or U8266 (N_8266,N_8018,N_8185);
nand U8267 (N_8267,N_8068,N_8114);
and U8268 (N_8268,N_8128,N_8041);
xor U8269 (N_8269,N_8166,N_8023);
or U8270 (N_8270,N_8015,N_8143);
nor U8271 (N_8271,N_8099,N_8183);
nand U8272 (N_8272,N_8164,N_8167);
xor U8273 (N_8273,N_8003,N_8050);
nor U8274 (N_8274,N_8012,N_8111);
or U8275 (N_8275,N_8014,N_8071);
nor U8276 (N_8276,N_8047,N_8139);
xor U8277 (N_8277,N_8044,N_8059);
nor U8278 (N_8278,N_8021,N_8150);
or U8279 (N_8279,N_8028,N_8178);
nand U8280 (N_8280,N_8063,N_8134);
nand U8281 (N_8281,N_8054,N_8031);
xnor U8282 (N_8282,N_8132,N_8024);
or U8283 (N_8283,N_8163,N_8157);
xor U8284 (N_8284,N_8086,N_8130);
and U8285 (N_8285,N_8002,N_8171);
and U8286 (N_8286,N_8016,N_8179);
nor U8287 (N_8287,N_8142,N_8140);
and U8288 (N_8288,N_8083,N_8146);
and U8289 (N_8289,N_8102,N_8026);
nor U8290 (N_8290,N_8136,N_8172);
and U8291 (N_8291,N_8022,N_8040);
nand U8292 (N_8292,N_8154,N_8013);
or U8293 (N_8293,N_8125,N_8110);
xnor U8294 (N_8294,N_8144,N_8076);
nor U8295 (N_8295,N_8107,N_8051);
xnor U8296 (N_8296,N_8064,N_8109);
nor U8297 (N_8297,N_8019,N_8131);
and U8298 (N_8298,N_8120,N_8184);
and U8299 (N_8299,N_8029,N_8005);
and U8300 (N_8300,N_8187,N_8080);
and U8301 (N_8301,N_8158,N_8181);
nand U8302 (N_8302,N_8088,N_8081);
and U8303 (N_8303,N_8073,N_8065);
nor U8304 (N_8304,N_8100,N_8185);
nor U8305 (N_8305,N_8186,N_8053);
nor U8306 (N_8306,N_8171,N_8060);
or U8307 (N_8307,N_8179,N_8149);
nand U8308 (N_8308,N_8096,N_8115);
xnor U8309 (N_8309,N_8018,N_8001);
and U8310 (N_8310,N_8054,N_8119);
or U8311 (N_8311,N_8061,N_8093);
and U8312 (N_8312,N_8161,N_8197);
xor U8313 (N_8313,N_8124,N_8178);
nor U8314 (N_8314,N_8046,N_8062);
or U8315 (N_8315,N_8019,N_8060);
nor U8316 (N_8316,N_8192,N_8020);
nand U8317 (N_8317,N_8124,N_8005);
nor U8318 (N_8318,N_8047,N_8027);
xor U8319 (N_8319,N_8136,N_8065);
and U8320 (N_8320,N_8178,N_8116);
nor U8321 (N_8321,N_8182,N_8102);
xor U8322 (N_8322,N_8059,N_8122);
and U8323 (N_8323,N_8112,N_8028);
xor U8324 (N_8324,N_8080,N_8193);
nand U8325 (N_8325,N_8004,N_8128);
xor U8326 (N_8326,N_8007,N_8101);
nand U8327 (N_8327,N_8097,N_8099);
nand U8328 (N_8328,N_8018,N_8169);
and U8329 (N_8329,N_8065,N_8039);
nand U8330 (N_8330,N_8086,N_8046);
or U8331 (N_8331,N_8199,N_8095);
nand U8332 (N_8332,N_8174,N_8164);
or U8333 (N_8333,N_8151,N_8098);
nand U8334 (N_8334,N_8084,N_8188);
xor U8335 (N_8335,N_8130,N_8094);
or U8336 (N_8336,N_8035,N_8167);
xor U8337 (N_8337,N_8011,N_8099);
nand U8338 (N_8338,N_8007,N_8109);
or U8339 (N_8339,N_8023,N_8127);
nand U8340 (N_8340,N_8021,N_8081);
and U8341 (N_8341,N_8057,N_8177);
nand U8342 (N_8342,N_8006,N_8022);
and U8343 (N_8343,N_8000,N_8172);
or U8344 (N_8344,N_8089,N_8050);
nand U8345 (N_8345,N_8084,N_8017);
or U8346 (N_8346,N_8011,N_8119);
and U8347 (N_8347,N_8051,N_8102);
nor U8348 (N_8348,N_8020,N_8081);
xnor U8349 (N_8349,N_8014,N_8194);
nor U8350 (N_8350,N_8038,N_8017);
nand U8351 (N_8351,N_8140,N_8120);
nand U8352 (N_8352,N_8193,N_8048);
nor U8353 (N_8353,N_8069,N_8084);
or U8354 (N_8354,N_8091,N_8150);
and U8355 (N_8355,N_8101,N_8164);
xor U8356 (N_8356,N_8112,N_8099);
nor U8357 (N_8357,N_8127,N_8002);
nor U8358 (N_8358,N_8163,N_8186);
or U8359 (N_8359,N_8165,N_8028);
or U8360 (N_8360,N_8002,N_8148);
nor U8361 (N_8361,N_8153,N_8176);
and U8362 (N_8362,N_8051,N_8004);
nor U8363 (N_8363,N_8056,N_8043);
and U8364 (N_8364,N_8063,N_8152);
nand U8365 (N_8365,N_8130,N_8156);
or U8366 (N_8366,N_8028,N_8020);
nand U8367 (N_8367,N_8189,N_8128);
and U8368 (N_8368,N_8161,N_8113);
xnor U8369 (N_8369,N_8031,N_8044);
nand U8370 (N_8370,N_8138,N_8049);
nand U8371 (N_8371,N_8050,N_8036);
and U8372 (N_8372,N_8136,N_8127);
or U8373 (N_8373,N_8149,N_8090);
xnor U8374 (N_8374,N_8083,N_8162);
nand U8375 (N_8375,N_8005,N_8198);
nand U8376 (N_8376,N_8161,N_8048);
xor U8377 (N_8377,N_8138,N_8012);
xnor U8378 (N_8378,N_8056,N_8197);
xor U8379 (N_8379,N_8147,N_8146);
or U8380 (N_8380,N_8121,N_8190);
xor U8381 (N_8381,N_8141,N_8176);
or U8382 (N_8382,N_8062,N_8137);
and U8383 (N_8383,N_8152,N_8048);
nor U8384 (N_8384,N_8086,N_8009);
nand U8385 (N_8385,N_8113,N_8060);
or U8386 (N_8386,N_8108,N_8040);
xor U8387 (N_8387,N_8072,N_8070);
nor U8388 (N_8388,N_8027,N_8152);
nor U8389 (N_8389,N_8031,N_8199);
or U8390 (N_8390,N_8116,N_8099);
nor U8391 (N_8391,N_8184,N_8074);
or U8392 (N_8392,N_8110,N_8111);
nor U8393 (N_8393,N_8134,N_8189);
or U8394 (N_8394,N_8127,N_8046);
and U8395 (N_8395,N_8046,N_8164);
and U8396 (N_8396,N_8104,N_8024);
or U8397 (N_8397,N_8113,N_8171);
and U8398 (N_8398,N_8079,N_8151);
nor U8399 (N_8399,N_8116,N_8023);
or U8400 (N_8400,N_8272,N_8356);
or U8401 (N_8401,N_8308,N_8284);
xnor U8402 (N_8402,N_8303,N_8217);
xnor U8403 (N_8403,N_8215,N_8366);
or U8404 (N_8404,N_8363,N_8261);
or U8405 (N_8405,N_8386,N_8315);
nand U8406 (N_8406,N_8210,N_8357);
nor U8407 (N_8407,N_8388,N_8282);
and U8408 (N_8408,N_8281,N_8376);
xor U8409 (N_8409,N_8227,N_8263);
nand U8410 (N_8410,N_8360,N_8289);
xnor U8411 (N_8411,N_8393,N_8211);
or U8412 (N_8412,N_8352,N_8270);
nor U8413 (N_8413,N_8321,N_8382);
or U8414 (N_8414,N_8390,N_8374);
and U8415 (N_8415,N_8209,N_8239);
and U8416 (N_8416,N_8257,N_8395);
nor U8417 (N_8417,N_8229,N_8365);
and U8418 (N_8418,N_8234,N_8245);
nor U8419 (N_8419,N_8293,N_8206);
nor U8420 (N_8420,N_8280,N_8320);
and U8421 (N_8421,N_8236,N_8219);
nand U8422 (N_8422,N_8380,N_8277);
and U8423 (N_8423,N_8364,N_8299);
nand U8424 (N_8424,N_8319,N_8231);
nor U8425 (N_8425,N_8342,N_8397);
and U8426 (N_8426,N_8240,N_8396);
nand U8427 (N_8427,N_8331,N_8248);
or U8428 (N_8428,N_8324,N_8249);
nor U8429 (N_8429,N_8333,N_8302);
nand U8430 (N_8430,N_8233,N_8246);
nand U8431 (N_8431,N_8335,N_8255);
nor U8432 (N_8432,N_8312,N_8351);
or U8433 (N_8433,N_8332,N_8346);
nor U8434 (N_8434,N_8225,N_8273);
xnor U8435 (N_8435,N_8200,N_8305);
nand U8436 (N_8436,N_8290,N_8330);
and U8437 (N_8437,N_8317,N_8337);
or U8438 (N_8438,N_8218,N_8325);
nor U8439 (N_8439,N_8349,N_8221);
xor U8440 (N_8440,N_8262,N_8264);
nor U8441 (N_8441,N_8220,N_8253);
nand U8442 (N_8442,N_8329,N_8328);
nor U8443 (N_8443,N_8361,N_8226);
or U8444 (N_8444,N_8347,N_8201);
or U8445 (N_8445,N_8367,N_8381);
xnor U8446 (N_8446,N_8230,N_8286);
xor U8447 (N_8447,N_8399,N_8216);
nor U8448 (N_8448,N_8327,N_8336);
nor U8449 (N_8449,N_8398,N_8295);
or U8450 (N_8450,N_8259,N_8223);
nor U8451 (N_8451,N_8222,N_8298);
nand U8452 (N_8452,N_8345,N_8278);
and U8453 (N_8453,N_8322,N_8256);
or U8454 (N_8454,N_8334,N_8268);
xor U8455 (N_8455,N_8297,N_8343);
nand U8456 (N_8456,N_8355,N_8387);
or U8457 (N_8457,N_8339,N_8274);
nand U8458 (N_8458,N_8244,N_8313);
xnor U8459 (N_8459,N_8285,N_8314);
xnor U8460 (N_8460,N_8348,N_8271);
or U8461 (N_8461,N_8232,N_8344);
nand U8462 (N_8462,N_8301,N_8247);
nor U8463 (N_8463,N_8237,N_8238);
and U8464 (N_8464,N_8241,N_8269);
and U8465 (N_8465,N_8311,N_8276);
xor U8466 (N_8466,N_8318,N_8260);
nor U8467 (N_8467,N_8212,N_8370);
nor U8468 (N_8468,N_8251,N_8267);
or U8469 (N_8469,N_8283,N_8300);
xor U8470 (N_8470,N_8250,N_8207);
nor U8471 (N_8471,N_8291,N_8304);
or U8472 (N_8472,N_8254,N_8307);
nor U8473 (N_8473,N_8306,N_8243);
xor U8474 (N_8474,N_8292,N_8316);
or U8475 (N_8475,N_8353,N_8202);
or U8476 (N_8476,N_8354,N_8242);
xnor U8477 (N_8477,N_8341,N_8214);
nand U8478 (N_8478,N_8326,N_8394);
or U8479 (N_8479,N_8208,N_8359);
and U8480 (N_8480,N_8235,N_8203);
and U8481 (N_8481,N_8275,N_8358);
nor U8482 (N_8482,N_8378,N_8288);
nor U8483 (N_8483,N_8266,N_8372);
or U8484 (N_8484,N_8375,N_8279);
nor U8485 (N_8485,N_8258,N_8224);
and U8486 (N_8486,N_8384,N_8205);
nor U8487 (N_8487,N_8385,N_8252);
nand U8488 (N_8488,N_8369,N_8294);
xnor U8489 (N_8489,N_8392,N_8368);
xor U8490 (N_8490,N_8340,N_8213);
nor U8491 (N_8491,N_8383,N_8309);
xor U8492 (N_8492,N_8389,N_8204);
nor U8493 (N_8493,N_8310,N_8323);
nand U8494 (N_8494,N_8373,N_8287);
and U8495 (N_8495,N_8379,N_8371);
xnor U8496 (N_8496,N_8265,N_8391);
and U8497 (N_8497,N_8362,N_8350);
nand U8498 (N_8498,N_8228,N_8338);
and U8499 (N_8499,N_8377,N_8296);
xor U8500 (N_8500,N_8235,N_8359);
nor U8501 (N_8501,N_8229,N_8258);
nor U8502 (N_8502,N_8208,N_8231);
nor U8503 (N_8503,N_8297,N_8309);
and U8504 (N_8504,N_8201,N_8227);
nor U8505 (N_8505,N_8321,N_8267);
nand U8506 (N_8506,N_8375,N_8244);
nor U8507 (N_8507,N_8340,N_8268);
nand U8508 (N_8508,N_8318,N_8374);
and U8509 (N_8509,N_8217,N_8203);
xor U8510 (N_8510,N_8229,N_8275);
nor U8511 (N_8511,N_8337,N_8281);
or U8512 (N_8512,N_8245,N_8373);
xor U8513 (N_8513,N_8382,N_8312);
or U8514 (N_8514,N_8297,N_8384);
nand U8515 (N_8515,N_8286,N_8372);
or U8516 (N_8516,N_8375,N_8388);
xor U8517 (N_8517,N_8326,N_8319);
and U8518 (N_8518,N_8361,N_8215);
nor U8519 (N_8519,N_8241,N_8245);
nor U8520 (N_8520,N_8328,N_8376);
and U8521 (N_8521,N_8266,N_8328);
xor U8522 (N_8522,N_8395,N_8271);
and U8523 (N_8523,N_8208,N_8378);
xor U8524 (N_8524,N_8222,N_8212);
and U8525 (N_8525,N_8307,N_8240);
nand U8526 (N_8526,N_8277,N_8248);
or U8527 (N_8527,N_8244,N_8391);
nand U8528 (N_8528,N_8245,N_8385);
xnor U8529 (N_8529,N_8255,N_8309);
and U8530 (N_8530,N_8355,N_8391);
and U8531 (N_8531,N_8295,N_8284);
and U8532 (N_8532,N_8218,N_8388);
or U8533 (N_8533,N_8204,N_8237);
xor U8534 (N_8534,N_8285,N_8225);
and U8535 (N_8535,N_8210,N_8372);
or U8536 (N_8536,N_8385,N_8283);
or U8537 (N_8537,N_8389,N_8315);
nor U8538 (N_8538,N_8337,N_8283);
nor U8539 (N_8539,N_8249,N_8279);
or U8540 (N_8540,N_8273,N_8283);
and U8541 (N_8541,N_8358,N_8345);
xnor U8542 (N_8542,N_8394,N_8324);
nor U8543 (N_8543,N_8370,N_8368);
nand U8544 (N_8544,N_8256,N_8391);
xor U8545 (N_8545,N_8362,N_8302);
or U8546 (N_8546,N_8389,N_8236);
nand U8547 (N_8547,N_8301,N_8295);
nor U8548 (N_8548,N_8303,N_8306);
or U8549 (N_8549,N_8254,N_8395);
or U8550 (N_8550,N_8351,N_8344);
nor U8551 (N_8551,N_8286,N_8284);
nand U8552 (N_8552,N_8269,N_8242);
nand U8553 (N_8553,N_8233,N_8315);
and U8554 (N_8554,N_8386,N_8348);
xnor U8555 (N_8555,N_8233,N_8318);
nor U8556 (N_8556,N_8256,N_8243);
nor U8557 (N_8557,N_8282,N_8247);
nor U8558 (N_8558,N_8205,N_8212);
nand U8559 (N_8559,N_8375,N_8374);
nand U8560 (N_8560,N_8263,N_8261);
or U8561 (N_8561,N_8295,N_8384);
and U8562 (N_8562,N_8322,N_8278);
or U8563 (N_8563,N_8371,N_8271);
and U8564 (N_8564,N_8343,N_8358);
nor U8565 (N_8565,N_8340,N_8222);
xnor U8566 (N_8566,N_8370,N_8282);
and U8567 (N_8567,N_8356,N_8323);
xnor U8568 (N_8568,N_8271,N_8238);
nor U8569 (N_8569,N_8221,N_8208);
nor U8570 (N_8570,N_8201,N_8267);
nor U8571 (N_8571,N_8290,N_8221);
xor U8572 (N_8572,N_8307,N_8297);
nand U8573 (N_8573,N_8300,N_8252);
and U8574 (N_8574,N_8215,N_8327);
xor U8575 (N_8575,N_8254,N_8272);
xor U8576 (N_8576,N_8358,N_8351);
xor U8577 (N_8577,N_8280,N_8318);
and U8578 (N_8578,N_8340,N_8302);
xnor U8579 (N_8579,N_8300,N_8296);
xor U8580 (N_8580,N_8319,N_8301);
nor U8581 (N_8581,N_8249,N_8225);
nand U8582 (N_8582,N_8380,N_8221);
and U8583 (N_8583,N_8224,N_8222);
xor U8584 (N_8584,N_8372,N_8338);
nor U8585 (N_8585,N_8216,N_8275);
or U8586 (N_8586,N_8229,N_8325);
xor U8587 (N_8587,N_8295,N_8275);
nand U8588 (N_8588,N_8221,N_8241);
xor U8589 (N_8589,N_8308,N_8242);
or U8590 (N_8590,N_8204,N_8233);
and U8591 (N_8591,N_8270,N_8321);
nand U8592 (N_8592,N_8348,N_8368);
or U8593 (N_8593,N_8354,N_8291);
nand U8594 (N_8594,N_8246,N_8339);
nand U8595 (N_8595,N_8288,N_8303);
or U8596 (N_8596,N_8213,N_8342);
nand U8597 (N_8597,N_8375,N_8360);
or U8598 (N_8598,N_8249,N_8268);
xor U8599 (N_8599,N_8387,N_8275);
or U8600 (N_8600,N_8455,N_8492);
nand U8601 (N_8601,N_8486,N_8525);
nor U8602 (N_8602,N_8528,N_8553);
xor U8603 (N_8603,N_8438,N_8567);
xnor U8604 (N_8604,N_8511,N_8459);
or U8605 (N_8605,N_8465,N_8470);
nand U8606 (N_8606,N_8504,N_8566);
xor U8607 (N_8607,N_8508,N_8558);
xnor U8608 (N_8608,N_8419,N_8480);
nor U8609 (N_8609,N_8513,N_8457);
nand U8610 (N_8610,N_8417,N_8533);
nor U8611 (N_8611,N_8440,N_8569);
or U8612 (N_8612,N_8412,N_8491);
xor U8613 (N_8613,N_8559,N_8561);
or U8614 (N_8614,N_8404,N_8434);
xnor U8615 (N_8615,N_8416,N_8531);
nor U8616 (N_8616,N_8532,N_8427);
or U8617 (N_8617,N_8414,N_8571);
or U8618 (N_8618,N_8517,N_8503);
nor U8619 (N_8619,N_8460,N_8501);
xnor U8620 (N_8620,N_8564,N_8599);
xor U8621 (N_8621,N_8496,N_8590);
xor U8622 (N_8622,N_8436,N_8595);
nand U8623 (N_8623,N_8518,N_8441);
nand U8624 (N_8624,N_8444,N_8497);
nand U8625 (N_8625,N_8529,N_8520);
or U8626 (N_8626,N_8439,N_8406);
xor U8627 (N_8627,N_8554,N_8542);
or U8628 (N_8628,N_8422,N_8579);
and U8629 (N_8629,N_8489,N_8562);
or U8630 (N_8630,N_8550,N_8487);
and U8631 (N_8631,N_8587,N_8410);
and U8632 (N_8632,N_8585,N_8546);
nand U8633 (N_8633,N_8573,N_8428);
xnor U8634 (N_8634,N_8583,N_8495);
or U8635 (N_8635,N_8452,N_8537);
or U8636 (N_8636,N_8424,N_8471);
nand U8637 (N_8637,N_8442,N_8538);
nand U8638 (N_8638,N_8556,N_8512);
xor U8639 (N_8639,N_8401,N_8402);
nand U8640 (N_8640,N_8431,N_8456);
or U8641 (N_8641,N_8478,N_8481);
or U8642 (N_8642,N_8475,N_8549);
nor U8643 (N_8643,N_8453,N_8530);
nor U8644 (N_8644,N_8548,N_8473);
and U8645 (N_8645,N_8499,N_8514);
and U8646 (N_8646,N_8403,N_8407);
and U8647 (N_8647,N_8461,N_8469);
xor U8648 (N_8648,N_8462,N_8575);
nor U8649 (N_8649,N_8433,N_8474);
xnor U8650 (N_8650,N_8408,N_8588);
nand U8651 (N_8651,N_8418,N_8448);
nand U8652 (N_8652,N_8420,N_8498);
and U8653 (N_8653,N_8409,N_8454);
or U8654 (N_8654,N_8540,N_8584);
and U8655 (N_8655,N_8527,N_8446);
nand U8656 (N_8656,N_8545,N_8415);
or U8657 (N_8657,N_8477,N_8581);
nand U8658 (N_8658,N_8524,N_8582);
or U8659 (N_8659,N_8464,N_8432);
nand U8660 (N_8660,N_8458,N_8502);
nand U8661 (N_8661,N_8534,N_8463);
or U8662 (N_8662,N_8572,N_8466);
nand U8663 (N_8663,N_8506,N_8577);
xnor U8664 (N_8664,N_8500,N_8536);
nand U8665 (N_8665,N_8543,N_8445);
or U8666 (N_8666,N_8560,N_8490);
nor U8667 (N_8667,N_8526,N_8598);
and U8668 (N_8668,N_8519,N_8488);
or U8669 (N_8669,N_8467,N_8535);
nand U8670 (N_8670,N_8426,N_8484);
xnor U8671 (N_8671,N_8443,N_8555);
and U8672 (N_8672,N_8578,N_8423);
nand U8673 (N_8673,N_8447,N_8565);
and U8674 (N_8674,N_8400,N_8509);
nor U8675 (N_8675,N_8476,N_8574);
xor U8676 (N_8676,N_8479,N_8586);
and U8677 (N_8677,N_8405,N_8435);
or U8678 (N_8678,N_8451,N_8449);
nor U8679 (N_8679,N_8516,N_8468);
or U8680 (N_8680,N_8594,N_8576);
xor U8681 (N_8681,N_8563,N_8437);
nand U8682 (N_8682,N_8570,N_8510);
and U8683 (N_8683,N_8591,N_8413);
and U8684 (N_8684,N_8557,N_8547);
or U8685 (N_8685,N_8515,N_8552);
or U8686 (N_8686,N_8485,N_8544);
or U8687 (N_8687,N_8589,N_8411);
xor U8688 (N_8688,N_8522,N_8580);
xnor U8689 (N_8689,N_8472,N_8551);
nand U8690 (N_8690,N_8505,N_8430);
or U8691 (N_8691,N_8592,N_8425);
or U8692 (N_8692,N_8507,N_8494);
xnor U8693 (N_8693,N_8482,N_8539);
nor U8694 (N_8694,N_8483,N_8523);
or U8695 (N_8695,N_8597,N_8596);
nor U8696 (N_8696,N_8450,N_8493);
nand U8697 (N_8697,N_8421,N_8593);
xnor U8698 (N_8698,N_8429,N_8541);
xor U8699 (N_8699,N_8521,N_8568);
nand U8700 (N_8700,N_8572,N_8479);
nor U8701 (N_8701,N_8439,N_8589);
xor U8702 (N_8702,N_8411,N_8466);
nor U8703 (N_8703,N_8421,N_8591);
and U8704 (N_8704,N_8458,N_8440);
or U8705 (N_8705,N_8422,N_8416);
nor U8706 (N_8706,N_8433,N_8461);
xnor U8707 (N_8707,N_8567,N_8537);
nor U8708 (N_8708,N_8458,N_8401);
nor U8709 (N_8709,N_8505,N_8462);
nor U8710 (N_8710,N_8539,N_8565);
and U8711 (N_8711,N_8496,N_8460);
or U8712 (N_8712,N_8443,N_8510);
nor U8713 (N_8713,N_8520,N_8468);
nand U8714 (N_8714,N_8416,N_8409);
or U8715 (N_8715,N_8576,N_8557);
nand U8716 (N_8716,N_8543,N_8443);
or U8717 (N_8717,N_8461,N_8595);
xor U8718 (N_8718,N_8436,N_8465);
and U8719 (N_8719,N_8401,N_8480);
nand U8720 (N_8720,N_8442,N_8428);
xor U8721 (N_8721,N_8528,N_8513);
nand U8722 (N_8722,N_8543,N_8467);
nor U8723 (N_8723,N_8561,N_8520);
nor U8724 (N_8724,N_8424,N_8454);
and U8725 (N_8725,N_8494,N_8552);
and U8726 (N_8726,N_8510,N_8432);
nand U8727 (N_8727,N_8408,N_8405);
nor U8728 (N_8728,N_8581,N_8567);
or U8729 (N_8729,N_8587,N_8480);
nor U8730 (N_8730,N_8426,N_8535);
xnor U8731 (N_8731,N_8579,N_8425);
xnor U8732 (N_8732,N_8455,N_8572);
and U8733 (N_8733,N_8565,N_8530);
and U8734 (N_8734,N_8596,N_8463);
xor U8735 (N_8735,N_8477,N_8534);
nand U8736 (N_8736,N_8560,N_8403);
nand U8737 (N_8737,N_8480,N_8538);
or U8738 (N_8738,N_8567,N_8422);
or U8739 (N_8739,N_8460,N_8509);
nor U8740 (N_8740,N_8578,N_8512);
and U8741 (N_8741,N_8584,N_8513);
and U8742 (N_8742,N_8595,N_8550);
xnor U8743 (N_8743,N_8412,N_8567);
or U8744 (N_8744,N_8589,N_8582);
nand U8745 (N_8745,N_8554,N_8425);
nor U8746 (N_8746,N_8422,N_8578);
and U8747 (N_8747,N_8494,N_8558);
nand U8748 (N_8748,N_8435,N_8460);
nand U8749 (N_8749,N_8516,N_8476);
xnor U8750 (N_8750,N_8542,N_8432);
nand U8751 (N_8751,N_8456,N_8401);
or U8752 (N_8752,N_8587,N_8569);
and U8753 (N_8753,N_8410,N_8526);
and U8754 (N_8754,N_8476,N_8474);
nand U8755 (N_8755,N_8461,N_8440);
or U8756 (N_8756,N_8582,N_8465);
and U8757 (N_8757,N_8434,N_8535);
or U8758 (N_8758,N_8481,N_8530);
nand U8759 (N_8759,N_8511,N_8562);
and U8760 (N_8760,N_8499,N_8406);
nor U8761 (N_8761,N_8517,N_8538);
and U8762 (N_8762,N_8429,N_8496);
xnor U8763 (N_8763,N_8438,N_8404);
nand U8764 (N_8764,N_8580,N_8596);
or U8765 (N_8765,N_8589,N_8576);
nand U8766 (N_8766,N_8417,N_8458);
or U8767 (N_8767,N_8578,N_8424);
xnor U8768 (N_8768,N_8572,N_8415);
and U8769 (N_8769,N_8451,N_8526);
or U8770 (N_8770,N_8518,N_8411);
nand U8771 (N_8771,N_8450,N_8462);
xnor U8772 (N_8772,N_8559,N_8525);
and U8773 (N_8773,N_8414,N_8543);
xnor U8774 (N_8774,N_8493,N_8586);
xnor U8775 (N_8775,N_8520,N_8586);
nor U8776 (N_8776,N_8440,N_8455);
xnor U8777 (N_8777,N_8471,N_8541);
and U8778 (N_8778,N_8445,N_8460);
and U8779 (N_8779,N_8503,N_8402);
xnor U8780 (N_8780,N_8401,N_8545);
nor U8781 (N_8781,N_8467,N_8402);
and U8782 (N_8782,N_8573,N_8445);
nand U8783 (N_8783,N_8462,N_8482);
or U8784 (N_8784,N_8442,N_8503);
nand U8785 (N_8785,N_8514,N_8532);
and U8786 (N_8786,N_8561,N_8578);
xor U8787 (N_8787,N_8581,N_8413);
nand U8788 (N_8788,N_8595,N_8466);
or U8789 (N_8789,N_8541,N_8424);
nor U8790 (N_8790,N_8462,N_8582);
or U8791 (N_8791,N_8581,N_8474);
nor U8792 (N_8792,N_8592,N_8463);
nand U8793 (N_8793,N_8466,N_8434);
and U8794 (N_8794,N_8425,N_8430);
and U8795 (N_8795,N_8507,N_8577);
xor U8796 (N_8796,N_8433,N_8558);
or U8797 (N_8797,N_8526,N_8415);
nor U8798 (N_8798,N_8517,N_8536);
and U8799 (N_8799,N_8516,N_8532);
or U8800 (N_8800,N_8673,N_8781);
nor U8801 (N_8801,N_8710,N_8670);
nor U8802 (N_8802,N_8602,N_8647);
or U8803 (N_8803,N_8649,N_8656);
nand U8804 (N_8804,N_8719,N_8745);
or U8805 (N_8805,N_8771,N_8623);
nor U8806 (N_8806,N_8757,N_8680);
xor U8807 (N_8807,N_8732,N_8629);
and U8808 (N_8808,N_8759,N_8603);
xor U8809 (N_8809,N_8788,N_8607);
nor U8810 (N_8810,N_8600,N_8690);
xor U8811 (N_8811,N_8679,N_8717);
xnor U8812 (N_8812,N_8702,N_8688);
xnor U8813 (N_8813,N_8659,N_8770);
or U8814 (N_8814,N_8753,N_8644);
nor U8815 (N_8815,N_8696,N_8733);
or U8816 (N_8816,N_8726,N_8618);
xor U8817 (N_8817,N_8638,N_8783);
nor U8818 (N_8818,N_8744,N_8764);
or U8819 (N_8819,N_8739,N_8798);
xor U8820 (N_8820,N_8677,N_8632);
nand U8821 (N_8821,N_8756,N_8791);
xnor U8822 (N_8822,N_8751,N_8766);
nor U8823 (N_8823,N_8635,N_8777);
xnor U8824 (N_8824,N_8691,N_8605);
nor U8825 (N_8825,N_8678,N_8760);
nor U8826 (N_8826,N_8620,N_8721);
and U8827 (N_8827,N_8650,N_8676);
nand U8828 (N_8828,N_8619,N_8708);
nand U8829 (N_8829,N_8754,N_8606);
xnor U8830 (N_8830,N_8707,N_8712);
nor U8831 (N_8831,N_8633,N_8713);
or U8832 (N_8832,N_8660,N_8748);
nor U8833 (N_8833,N_8682,N_8609);
nor U8834 (N_8834,N_8684,N_8686);
nand U8835 (N_8835,N_8630,N_8782);
or U8836 (N_8836,N_8703,N_8790);
nor U8837 (N_8837,N_8674,N_8625);
and U8838 (N_8838,N_8627,N_8740);
nor U8839 (N_8839,N_8742,N_8665);
nand U8840 (N_8840,N_8767,N_8731);
nand U8841 (N_8841,N_8768,N_8769);
or U8842 (N_8842,N_8683,N_8792);
nor U8843 (N_8843,N_8785,N_8615);
nand U8844 (N_8844,N_8709,N_8750);
and U8845 (N_8845,N_8755,N_8737);
and U8846 (N_8846,N_8761,N_8648);
or U8847 (N_8847,N_8711,N_8700);
nor U8848 (N_8848,N_8714,N_8669);
or U8849 (N_8849,N_8734,N_8720);
xor U8850 (N_8850,N_8786,N_8765);
and U8851 (N_8851,N_8773,N_8672);
xor U8852 (N_8852,N_8749,N_8657);
nor U8853 (N_8853,N_8701,N_8794);
or U8854 (N_8854,N_8653,N_8780);
nor U8855 (N_8855,N_8741,N_8675);
or U8856 (N_8856,N_8687,N_8774);
and U8857 (N_8857,N_8637,N_8671);
and U8858 (N_8858,N_8705,N_8692);
and U8859 (N_8859,N_8746,N_8730);
nand U8860 (N_8860,N_8735,N_8795);
nand U8861 (N_8861,N_8784,N_8747);
nor U8862 (N_8862,N_8729,N_8614);
nand U8863 (N_8863,N_8601,N_8645);
or U8864 (N_8864,N_8681,N_8642);
and U8865 (N_8865,N_8695,N_8778);
nand U8866 (N_8866,N_8654,N_8662);
xor U8867 (N_8867,N_8722,N_8736);
nor U8868 (N_8868,N_8789,N_8631);
and U8869 (N_8869,N_8636,N_8706);
xnor U8870 (N_8870,N_8697,N_8775);
and U8871 (N_8871,N_8758,N_8655);
or U8872 (N_8872,N_8698,N_8664);
nor U8873 (N_8873,N_8715,N_8793);
nand U8874 (N_8874,N_8704,N_8616);
xnor U8875 (N_8875,N_8752,N_8652);
xor U8876 (N_8876,N_8689,N_8661);
and U8877 (N_8877,N_8762,N_8694);
nand U8878 (N_8878,N_8699,N_8628);
or U8879 (N_8879,N_8763,N_8718);
and U8880 (N_8880,N_8621,N_8738);
xnor U8881 (N_8881,N_8643,N_8796);
nand U8882 (N_8882,N_8613,N_8622);
xnor U8883 (N_8883,N_8626,N_8723);
nand U8884 (N_8884,N_8772,N_8685);
and U8885 (N_8885,N_8639,N_8640);
nor U8886 (N_8886,N_8604,N_8667);
nor U8887 (N_8887,N_8641,N_8617);
nand U8888 (N_8888,N_8797,N_8651);
nor U8889 (N_8889,N_8608,N_8724);
nor U8890 (N_8890,N_8668,N_8728);
nor U8891 (N_8891,N_8716,N_8634);
and U8892 (N_8892,N_8663,N_8743);
nor U8893 (N_8893,N_8658,N_8799);
and U8894 (N_8894,N_8610,N_8646);
or U8895 (N_8895,N_8779,N_8693);
or U8896 (N_8896,N_8612,N_8611);
and U8897 (N_8897,N_8624,N_8787);
or U8898 (N_8898,N_8776,N_8666);
or U8899 (N_8899,N_8727,N_8725);
nor U8900 (N_8900,N_8626,N_8632);
and U8901 (N_8901,N_8724,N_8674);
nor U8902 (N_8902,N_8796,N_8737);
or U8903 (N_8903,N_8681,N_8671);
xnor U8904 (N_8904,N_8643,N_8684);
or U8905 (N_8905,N_8693,N_8704);
nor U8906 (N_8906,N_8637,N_8720);
or U8907 (N_8907,N_8688,N_8753);
xnor U8908 (N_8908,N_8741,N_8728);
xor U8909 (N_8909,N_8749,N_8697);
nand U8910 (N_8910,N_8729,N_8793);
or U8911 (N_8911,N_8690,N_8796);
or U8912 (N_8912,N_8706,N_8686);
xor U8913 (N_8913,N_8724,N_8651);
and U8914 (N_8914,N_8651,N_8693);
or U8915 (N_8915,N_8711,N_8759);
and U8916 (N_8916,N_8664,N_8638);
xnor U8917 (N_8917,N_8734,N_8672);
or U8918 (N_8918,N_8715,N_8655);
xnor U8919 (N_8919,N_8620,N_8756);
nand U8920 (N_8920,N_8714,N_8645);
xnor U8921 (N_8921,N_8604,N_8630);
or U8922 (N_8922,N_8746,N_8600);
and U8923 (N_8923,N_8606,N_8797);
nor U8924 (N_8924,N_8750,N_8653);
nand U8925 (N_8925,N_8614,N_8780);
nor U8926 (N_8926,N_8730,N_8683);
nor U8927 (N_8927,N_8609,N_8615);
and U8928 (N_8928,N_8785,N_8641);
or U8929 (N_8929,N_8756,N_8669);
and U8930 (N_8930,N_8763,N_8794);
nor U8931 (N_8931,N_8717,N_8632);
xnor U8932 (N_8932,N_8745,N_8605);
or U8933 (N_8933,N_8722,N_8650);
xor U8934 (N_8934,N_8742,N_8600);
nand U8935 (N_8935,N_8774,N_8661);
xnor U8936 (N_8936,N_8634,N_8735);
nand U8937 (N_8937,N_8643,N_8752);
nor U8938 (N_8938,N_8658,N_8607);
xnor U8939 (N_8939,N_8624,N_8623);
nor U8940 (N_8940,N_8788,N_8643);
or U8941 (N_8941,N_8744,N_8616);
nor U8942 (N_8942,N_8697,N_8620);
nor U8943 (N_8943,N_8767,N_8790);
and U8944 (N_8944,N_8650,N_8633);
nand U8945 (N_8945,N_8765,N_8653);
nand U8946 (N_8946,N_8638,N_8707);
nand U8947 (N_8947,N_8768,N_8766);
and U8948 (N_8948,N_8693,N_8645);
or U8949 (N_8949,N_8615,N_8641);
nor U8950 (N_8950,N_8685,N_8644);
or U8951 (N_8951,N_8698,N_8682);
or U8952 (N_8952,N_8655,N_8788);
nand U8953 (N_8953,N_8713,N_8790);
and U8954 (N_8954,N_8654,N_8715);
nor U8955 (N_8955,N_8789,N_8647);
xnor U8956 (N_8956,N_8736,N_8701);
and U8957 (N_8957,N_8734,N_8660);
nor U8958 (N_8958,N_8698,N_8639);
xor U8959 (N_8959,N_8773,N_8739);
xor U8960 (N_8960,N_8680,N_8750);
or U8961 (N_8961,N_8770,N_8610);
nor U8962 (N_8962,N_8662,N_8717);
or U8963 (N_8963,N_8607,N_8670);
nand U8964 (N_8964,N_8667,N_8673);
and U8965 (N_8965,N_8735,N_8760);
xnor U8966 (N_8966,N_8771,N_8688);
xor U8967 (N_8967,N_8796,N_8745);
or U8968 (N_8968,N_8608,N_8643);
and U8969 (N_8969,N_8760,N_8625);
nor U8970 (N_8970,N_8792,N_8691);
or U8971 (N_8971,N_8725,N_8665);
and U8972 (N_8972,N_8744,N_8645);
and U8973 (N_8973,N_8675,N_8638);
nor U8974 (N_8974,N_8727,N_8776);
nor U8975 (N_8975,N_8662,N_8640);
or U8976 (N_8976,N_8772,N_8760);
nor U8977 (N_8977,N_8721,N_8609);
nor U8978 (N_8978,N_8625,N_8701);
nand U8979 (N_8979,N_8791,N_8731);
and U8980 (N_8980,N_8629,N_8746);
xor U8981 (N_8981,N_8720,N_8616);
xor U8982 (N_8982,N_8705,N_8769);
xnor U8983 (N_8983,N_8738,N_8637);
and U8984 (N_8984,N_8741,N_8779);
nor U8985 (N_8985,N_8747,N_8600);
nor U8986 (N_8986,N_8610,N_8618);
nand U8987 (N_8987,N_8614,N_8747);
nand U8988 (N_8988,N_8738,N_8790);
or U8989 (N_8989,N_8647,N_8720);
and U8990 (N_8990,N_8704,N_8724);
xnor U8991 (N_8991,N_8616,N_8746);
nor U8992 (N_8992,N_8640,N_8729);
or U8993 (N_8993,N_8760,N_8734);
or U8994 (N_8994,N_8621,N_8736);
and U8995 (N_8995,N_8796,N_8601);
or U8996 (N_8996,N_8669,N_8683);
or U8997 (N_8997,N_8710,N_8774);
xor U8998 (N_8998,N_8758,N_8739);
and U8999 (N_8999,N_8762,N_8646);
or U9000 (N_9000,N_8900,N_8934);
xor U9001 (N_9001,N_8924,N_8842);
or U9002 (N_9002,N_8894,N_8948);
and U9003 (N_9003,N_8880,N_8888);
and U9004 (N_9004,N_8884,N_8913);
nor U9005 (N_9005,N_8930,N_8808);
or U9006 (N_9006,N_8921,N_8856);
or U9007 (N_9007,N_8833,N_8803);
nor U9008 (N_9008,N_8931,N_8836);
or U9009 (N_9009,N_8974,N_8994);
and U9010 (N_9010,N_8818,N_8889);
nand U9011 (N_9011,N_8867,N_8824);
and U9012 (N_9012,N_8862,N_8831);
or U9013 (N_9013,N_8855,N_8935);
xor U9014 (N_9014,N_8834,N_8812);
and U9015 (N_9015,N_8910,N_8835);
nand U9016 (N_9016,N_8852,N_8807);
xor U9017 (N_9017,N_8901,N_8904);
xor U9018 (N_9018,N_8967,N_8866);
nor U9019 (N_9019,N_8999,N_8980);
nand U9020 (N_9020,N_8938,N_8919);
or U9021 (N_9021,N_8987,N_8928);
or U9022 (N_9022,N_8870,N_8979);
nor U9023 (N_9023,N_8861,N_8827);
nor U9024 (N_9024,N_8922,N_8874);
and U9025 (N_9025,N_8925,N_8939);
and U9026 (N_9026,N_8860,N_8891);
or U9027 (N_9027,N_8973,N_8848);
nand U9028 (N_9028,N_8850,N_8876);
or U9029 (N_9029,N_8964,N_8975);
nor U9030 (N_9030,N_8943,N_8918);
xnor U9031 (N_9031,N_8929,N_8896);
xor U9032 (N_9032,N_8817,N_8877);
and U9033 (N_9033,N_8906,N_8909);
nor U9034 (N_9034,N_8816,N_8970);
xor U9035 (N_9035,N_8957,N_8941);
xor U9036 (N_9036,N_8926,N_8840);
nor U9037 (N_9037,N_8813,N_8996);
or U9038 (N_9038,N_8841,N_8912);
xnor U9039 (N_9039,N_8832,N_8917);
or U9040 (N_9040,N_8956,N_8905);
xor U9041 (N_9041,N_8998,N_8985);
nand U9042 (N_9042,N_8819,N_8871);
nand U9043 (N_9043,N_8863,N_8971);
or U9044 (N_9044,N_8950,N_8826);
and U9045 (N_9045,N_8969,N_8893);
nand U9046 (N_9046,N_8959,N_8927);
xor U9047 (N_9047,N_8875,N_8864);
xnor U9048 (N_9048,N_8993,N_8997);
xor U9049 (N_9049,N_8873,N_8991);
and U9050 (N_9050,N_8823,N_8945);
or U9051 (N_9051,N_8898,N_8839);
xor U9052 (N_9052,N_8857,N_8853);
and U9053 (N_9053,N_8802,N_8854);
or U9054 (N_9054,N_8811,N_8953);
xor U9055 (N_9055,N_8830,N_8890);
nor U9056 (N_9056,N_8962,N_8806);
or U9057 (N_9057,N_8892,N_8878);
nand U9058 (N_9058,N_8859,N_8966);
nor U9059 (N_9059,N_8984,N_8915);
or U9060 (N_9060,N_8820,N_8887);
and U9061 (N_9061,N_8988,N_8911);
xor U9062 (N_9062,N_8828,N_8940);
and U9063 (N_9063,N_8804,N_8849);
xor U9064 (N_9064,N_8937,N_8825);
nand U9065 (N_9065,N_8879,N_8989);
nor U9066 (N_9066,N_8872,N_8936);
or U9067 (N_9067,N_8903,N_8844);
or U9068 (N_9068,N_8978,N_8965);
nor U9069 (N_9069,N_8932,N_8983);
nand U9070 (N_9070,N_8810,N_8829);
nand U9071 (N_9071,N_8951,N_8869);
nor U9072 (N_9072,N_8881,N_8986);
or U9073 (N_9073,N_8837,N_8920);
nor U9074 (N_9074,N_8846,N_8809);
and U9075 (N_9075,N_8982,N_8851);
and U9076 (N_9076,N_8963,N_8883);
nor U9077 (N_9077,N_8899,N_8995);
nand U9078 (N_9078,N_8805,N_8845);
xor U9079 (N_9079,N_8858,N_8946);
and U9080 (N_9080,N_8908,N_8990);
and U9081 (N_9081,N_8960,N_8885);
and U9082 (N_9082,N_8843,N_8821);
or U9083 (N_9083,N_8952,N_8907);
and U9084 (N_9084,N_8801,N_8897);
or U9085 (N_9085,N_8958,N_8800);
nor U9086 (N_9086,N_8976,N_8949);
nor U9087 (N_9087,N_8972,N_8955);
or U9088 (N_9088,N_8902,N_8822);
or U9089 (N_9089,N_8886,N_8914);
nor U9090 (N_9090,N_8868,N_8981);
nand U9091 (N_9091,N_8968,N_8977);
nand U9092 (N_9092,N_8814,N_8933);
xor U9093 (N_9093,N_8815,N_8954);
and U9094 (N_9094,N_8947,N_8865);
xnor U9095 (N_9095,N_8923,N_8961);
xnor U9096 (N_9096,N_8838,N_8847);
xor U9097 (N_9097,N_8895,N_8944);
or U9098 (N_9098,N_8916,N_8942);
xnor U9099 (N_9099,N_8882,N_8992);
xnor U9100 (N_9100,N_8879,N_8928);
xor U9101 (N_9101,N_8811,N_8815);
nand U9102 (N_9102,N_8801,N_8841);
nand U9103 (N_9103,N_8913,N_8896);
and U9104 (N_9104,N_8814,N_8867);
or U9105 (N_9105,N_8883,N_8839);
or U9106 (N_9106,N_8973,N_8951);
nor U9107 (N_9107,N_8902,N_8994);
xor U9108 (N_9108,N_8890,N_8828);
nor U9109 (N_9109,N_8872,N_8963);
xor U9110 (N_9110,N_8822,N_8910);
nand U9111 (N_9111,N_8938,N_8846);
xnor U9112 (N_9112,N_8964,N_8869);
and U9113 (N_9113,N_8820,N_8926);
nor U9114 (N_9114,N_8928,N_8995);
nand U9115 (N_9115,N_8823,N_8954);
or U9116 (N_9116,N_8833,N_8922);
nor U9117 (N_9117,N_8885,N_8979);
nor U9118 (N_9118,N_8995,N_8923);
nand U9119 (N_9119,N_8973,N_8870);
or U9120 (N_9120,N_8978,N_8866);
or U9121 (N_9121,N_8904,N_8876);
and U9122 (N_9122,N_8989,N_8987);
nand U9123 (N_9123,N_8890,N_8996);
nor U9124 (N_9124,N_8905,N_8862);
xnor U9125 (N_9125,N_8953,N_8840);
and U9126 (N_9126,N_8910,N_8991);
xor U9127 (N_9127,N_8820,N_8877);
or U9128 (N_9128,N_8827,N_8871);
xnor U9129 (N_9129,N_8906,N_8998);
xnor U9130 (N_9130,N_8935,N_8827);
or U9131 (N_9131,N_8936,N_8987);
nand U9132 (N_9132,N_8854,N_8841);
nand U9133 (N_9133,N_8897,N_8904);
or U9134 (N_9134,N_8966,N_8861);
nand U9135 (N_9135,N_8818,N_8823);
nand U9136 (N_9136,N_8979,N_8916);
xnor U9137 (N_9137,N_8991,N_8901);
xnor U9138 (N_9138,N_8873,N_8903);
nor U9139 (N_9139,N_8820,N_8861);
nand U9140 (N_9140,N_8819,N_8831);
nand U9141 (N_9141,N_8941,N_8872);
xor U9142 (N_9142,N_8901,N_8997);
nor U9143 (N_9143,N_8902,N_8861);
or U9144 (N_9144,N_8949,N_8825);
or U9145 (N_9145,N_8927,N_8840);
and U9146 (N_9146,N_8952,N_8836);
and U9147 (N_9147,N_8834,N_8936);
or U9148 (N_9148,N_8994,N_8943);
nand U9149 (N_9149,N_8923,N_8921);
nor U9150 (N_9150,N_8822,N_8909);
xor U9151 (N_9151,N_8931,N_8868);
nand U9152 (N_9152,N_8828,N_8918);
nor U9153 (N_9153,N_8905,N_8871);
xnor U9154 (N_9154,N_8919,N_8911);
and U9155 (N_9155,N_8879,N_8949);
or U9156 (N_9156,N_8927,N_8831);
and U9157 (N_9157,N_8895,N_8996);
or U9158 (N_9158,N_8889,N_8959);
and U9159 (N_9159,N_8940,N_8813);
xor U9160 (N_9160,N_8983,N_8937);
or U9161 (N_9161,N_8823,N_8871);
xnor U9162 (N_9162,N_8983,N_8984);
nand U9163 (N_9163,N_8976,N_8988);
or U9164 (N_9164,N_8846,N_8856);
and U9165 (N_9165,N_8906,N_8904);
and U9166 (N_9166,N_8804,N_8867);
or U9167 (N_9167,N_8976,N_8935);
nor U9168 (N_9168,N_8824,N_8845);
and U9169 (N_9169,N_8966,N_8958);
and U9170 (N_9170,N_8965,N_8934);
nor U9171 (N_9171,N_8923,N_8864);
xnor U9172 (N_9172,N_8976,N_8892);
xor U9173 (N_9173,N_8904,N_8921);
and U9174 (N_9174,N_8909,N_8975);
and U9175 (N_9175,N_8829,N_8811);
nor U9176 (N_9176,N_8948,N_8883);
nor U9177 (N_9177,N_8839,N_8818);
and U9178 (N_9178,N_8879,N_8852);
nand U9179 (N_9179,N_8959,N_8819);
or U9180 (N_9180,N_8859,N_8953);
xor U9181 (N_9181,N_8806,N_8935);
nand U9182 (N_9182,N_8949,N_8947);
or U9183 (N_9183,N_8884,N_8970);
nor U9184 (N_9184,N_8913,N_8872);
and U9185 (N_9185,N_8863,N_8827);
or U9186 (N_9186,N_8931,N_8967);
nand U9187 (N_9187,N_8861,N_8926);
xnor U9188 (N_9188,N_8983,N_8805);
and U9189 (N_9189,N_8893,N_8867);
or U9190 (N_9190,N_8830,N_8807);
nand U9191 (N_9191,N_8851,N_8904);
xor U9192 (N_9192,N_8805,N_8910);
and U9193 (N_9193,N_8996,N_8800);
xnor U9194 (N_9194,N_8869,N_8918);
xor U9195 (N_9195,N_8946,N_8830);
nor U9196 (N_9196,N_8904,N_8891);
nand U9197 (N_9197,N_8818,N_8899);
xnor U9198 (N_9198,N_8995,N_8851);
or U9199 (N_9199,N_8882,N_8972);
nand U9200 (N_9200,N_9137,N_9167);
xor U9201 (N_9201,N_9071,N_9132);
and U9202 (N_9202,N_9171,N_9007);
xnor U9203 (N_9203,N_9063,N_9002);
or U9204 (N_9204,N_9060,N_9178);
nor U9205 (N_9205,N_9086,N_9028);
or U9206 (N_9206,N_9116,N_9089);
and U9207 (N_9207,N_9062,N_9075);
or U9208 (N_9208,N_9164,N_9168);
or U9209 (N_9209,N_9038,N_9103);
or U9210 (N_9210,N_9154,N_9165);
nand U9211 (N_9211,N_9070,N_9117);
xnor U9212 (N_9212,N_9022,N_9072);
and U9213 (N_9213,N_9145,N_9140);
or U9214 (N_9214,N_9162,N_9026);
or U9215 (N_9215,N_9073,N_9106);
xnor U9216 (N_9216,N_9199,N_9149);
xor U9217 (N_9217,N_9064,N_9045);
xnor U9218 (N_9218,N_9197,N_9081);
and U9219 (N_9219,N_9047,N_9151);
xor U9220 (N_9220,N_9015,N_9100);
nor U9221 (N_9221,N_9169,N_9025);
xor U9222 (N_9222,N_9156,N_9146);
nor U9223 (N_9223,N_9041,N_9125);
nand U9224 (N_9224,N_9166,N_9195);
nand U9225 (N_9225,N_9068,N_9061);
nand U9226 (N_9226,N_9010,N_9190);
and U9227 (N_9227,N_9191,N_9055);
and U9228 (N_9228,N_9155,N_9127);
nor U9229 (N_9229,N_9067,N_9054);
nor U9230 (N_9230,N_9076,N_9153);
or U9231 (N_9231,N_9194,N_9152);
and U9232 (N_9232,N_9115,N_9148);
xnor U9233 (N_9233,N_9131,N_9113);
nor U9234 (N_9234,N_9193,N_9079);
nand U9235 (N_9235,N_9069,N_9035);
nand U9236 (N_9236,N_9094,N_9129);
nor U9237 (N_9237,N_9024,N_9180);
nor U9238 (N_9238,N_9143,N_9056);
nor U9239 (N_9239,N_9017,N_9179);
nor U9240 (N_9240,N_9001,N_9074);
and U9241 (N_9241,N_9078,N_9130);
or U9242 (N_9242,N_9059,N_9107);
nor U9243 (N_9243,N_9181,N_9021);
or U9244 (N_9244,N_9098,N_9009);
nor U9245 (N_9245,N_9049,N_9088);
xnor U9246 (N_9246,N_9008,N_9095);
and U9247 (N_9247,N_9192,N_9004);
xnor U9248 (N_9248,N_9150,N_9034);
nor U9249 (N_9249,N_9003,N_9039);
nand U9250 (N_9250,N_9011,N_9087);
xnor U9251 (N_9251,N_9093,N_9048);
xor U9252 (N_9252,N_9083,N_9046);
xnor U9253 (N_9253,N_9027,N_9033);
nand U9254 (N_9254,N_9018,N_9160);
xor U9255 (N_9255,N_9013,N_9043);
xnor U9256 (N_9256,N_9092,N_9044);
nor U9257 (N_9257,N_9114,N_9198);
xor U9258 (N_9258,N_9090,N_9097);
or U9259 (N_9259,N_9030,N_9066);
xnor U9260 (N_9260,N_9112,N_9020);
or U9261 (N_9261,N_9108,N_9082);
nand U9262 (N_9262,N_9172,N_9111);
xor U9263 (N_9263,N_9173,N_9144);
nand U9264 (N_9264,N_9184,N_9105);
xor U9265 (N_9265,N_9077,N_9109);
nand U9266 (N_9266,N_9120,N_9005);
xnor U9267 (N_9267,N_9000,N_9012);
nand U9268 (N_9268,N_9029,N_9136);
nor U9269 (N_9269,N_9158,N_9157);
or U9270 (N_9270,N_9182,N_9189);
nor U9271 (N_9271,N_9177,N_9176);
nor U9272 (N_9272,N_9186,N_9118);
or U9273 (N_9273,N_9174,N_9040);
or U9274 (N_9274,N_9096,N_9187);
or U9275 (N_9275,N_9019,N_9124);
or U9276 (N_9276,N_9123,N_9147);
or U9277 (N_9277,N_9052,N_9091);
nor U9278 (N_9278,N_9104,N_9037);
or U9279 (N_9279,N_9185,N_9175);
xor U9280 (N_9280,N_9080,N_9138);
or U9281 (N_9281,N_9036,N_9119);
and U9282 (N_9282,N_9042,N_9050);
or U9283 (N_9283,N_9128,N_9053);
or U9284 (N_9284,N_9183,N_9196);
xor U9285 (N_9285,N_9084,N_9121);
and U9286 (N_9286,N_9099,N_9134);
nand U9287 (N_9287,N_9102,N_9133);
xor U9288 (N_9288,N_9101,N_9065);
xor U9289 (N_9289,N_9141,N_9161);
and U9290 (N_9290,N_9135,N_9032);
nand U9291 (N_9291,N_9016,N_9110);
xnor U9292 (N_9292,N_9031,N_9139);
or U9293 (N_9293,N_9023,N_9142);
xnor U9294 (N_9294,N_9051,N_9122);
xnor U9295 (N_9295,N_9159,N_9188);
xnor U9296 (N_9296,N_9170,N_9014);
nor U9297 (N_9297,N_9058,N_9006);
and U9298 (N_9298,N_9126,N_9085);
xor U9299 (N_9299,N_9163,N_9057);
and U9300 (N_9300,N_9131,N_9015);
or U9301 (N_9301,N_9195,N_9088);
nor U9302 (N_9302,N_9169,N_9074);
or U9303 (N_9303,N_9067,N_9014);
and U9304 (N_9304,N_9080,N_9184);
and U9305 (N_9305,N_9028,N_9080);
xor U9306 (N_9306,N_9078,N_9198);
nor U9307 (N_9307,N_9161,N_9197);
and U9308 (N_9308,N_9199,N_9179);
and U9309 (N_9309,N_9090,N_9052);
and U9310 (N_9310,N_9002,N_9194);
nand U9311 (N_9311,N_9058,N_9086);
and U9312 (N_9312,N_9005,N_9009);
or U9313 (N_9313,N_9020,N_9039);
and U9314 (N_9314,N_9025,N_9122);
xnor U9315 (N_9315,N_9040,N_9190);
nor U9316 (N_9316,N_9071,N_9093);
nand U9317 (N_9317,N_9083,N_9142);
or U9318 (N_9318,N_9195,N_9101);
or U9319 (N_9319,N_9016,N_9042);
nand U9320 (N_9320,N_9169,N_9122);
xnor U9321 (N_9321,N_9191,N_9035);
and U9322 (N_9322,N_9009,N_9176);
nand U9323 (N_9323,N_9141,N_9042);
or U9324 (N_9324,N_9143,N_9147);
xor U9325 (N_9325,N_9194,N_9091);
xor U9326 (N_9326,N_9167,N_9134);
nand U9327 (N_9327,N_9071,N_9080);
nand U9328 (N_9328,N_9047,N_9187);
nor U9329 (N_9329,N_9050,N_9139);
or U9330 (N_9330,N_9139,N_9013);
and U9331 (N_9331,N_9122,N_9001);
and U9332 (N_9332,N_9125,N_9178);
nor U9333 (N_9333,N_9001,N_9041);
nand U9334 (N_9334,N_9190,N_9117);
xnor U9335 (N_9335,N_9175,N_9117);
and U9336 (N_9336,N_9049,N_9180);
nor U9337 (N_9337,N_9050,N_9188);
nor U9338 (N_9338,N_9140,N_9114);
or U9339 (N_9339,N_9166,N_9162);
nand U9340 (N_9340,N_9198,N_9190);
xor U9341 (N_9341,N_9175,N_9105);
nor U9342 (N_9342,N_9062,N_9002);
nand U9343 (N_9343,N_9028,N_9152);
and U9344 (N_9344,N_9046,N_9044);
and U9345 (N_9345,N_9050,N_9012);
nor U9346 (N_9346,N_9148,N_9167);
and U9347 (N_9347,N_9190,N_9062);
xor U9348 (N_9348,N_9036,N_9191);
or U9349 (N_9349,N_9132,N_9013);
or U9350 (N_9350,N_9043,N_9050);
xnor U9351 (N_9351,N_9015,N_9057);
xor U9352 (N_9352,N_9014,N_9126);
or U9353 (N_9353,N_9080,N_9112);
and U9354 (N_9354,N_9121,N_9159);
nand U9355 (N_9355,N_9128,N_9169);
xnor U9356 (N_9356,N_9130,N_9153);
or U9357 (N_9357,N_9168,N_9064);
nor U9358 (N_9358,N_9007,N_9040);
and U9359 (N_9359,N_9172,N_9178);
or U9360 (N_9360,N_9070,N_9163);
nor U9361 (N_9361,N_9121,N_9047);
nor U9362 (N_9362,N_9030,N_9065);
or U9363 (N_9363,N_9022,N_9181);
nor U9364 (N_9364,N_9121,N_9048);
and U9365 (N_9365,N_9103,N_9108);
nand U9366 (N_9366,N_9029,N_9178);
and U9367 (N_9367,N_9073,N_9118);
nor U9368 (N_9368,N_9078,N_9017);
or U9369 (N_9369,N_9114,N_9030);
nor U9370 (N_9370,N_9049,N_9001);
nor U9371 (N_9371,N_9067,N_9174);
and U9372 (N_9372,N_9151,N_9090);
xor U9373 (N_9373,N_9097,N_9119);
or U9374 (N_9374,N_9021,N_9119);
and U9375 (N_9375,N_9039,N_9144);
and U9376 (N_9376,N_9199,N_9182);
and U9377 (N_9377,N_9024,N_9037);
nor U9378 (N_9378,N_9158,N_9035);
nor U9379 (N_9379,N_9001,N_9124);
nor U9380 (N_9380,N_9084,N_9072);
or U9381 (N_9381,N_9157,N_9075);
and U9382 (N_9382,N_9083,N_9082);
xor U9383 (N_9383,N_9068,N_9089);
nor U9384 (N_9384,N_9182,N_9192);
xnor U9385 (N_9385,N_9031,N_9068);
xnor U9386 (N_9386,N_9031,N_9189);
or U9387 (N_9387,N_9170,N_9187);
nor U9388 (N_9388,N_9172,N_9006);
xor U9389 (N_9389,N_9125,N_9175);
xor U9390 (N_9390,N_9190,N_9130);
or U9391 (N_9391,N_9057,N_9026);
and U9392 (N_9392,N_9046,N_9085);
nor U9393 (N_9393,N_9172,N_9171);
and U9394 (N_9394,N_9076,N_9149);
and U9395 (N_9395,N_9079,N_9063);
and U9396 (N_9396,N_9000,N_9001);
and U9397 (N_9397,N_9129,N_9156);
or U9398 (N_9398,N_9056,N_9063);
nand U9399 (N_9399,N_9095,N_9048);
or U9400 (N_9400,N_9387,N_9352);
nand U9401 (N_9401,N_9367,N_9386);
or U9402 (N_9402,N_9339,N_9200);
xnor U9403 (N_9403,N_9249,N_9300);
and U9404 (N_9404,N_9329,N_9284);
or U9405 (N_9405,N_9356,N_9395);
nor U9406 (N_9406,N_9354,N_9326);
nor U9407 (N_9407,N_9266,N_9269);
or U9408 (N_9408,N_9226,N_9327);
and U9409 (N_9409,N_9325,N_9260);
or U9410 (N_9410,N_9212,N_9308);
xor U9411 (N_9411,N_9231,N_9285);
or U9412 (N_9412,N_9365,N_9235);
nand U9413 (N_9413,N_9241,N_9273);
xnor U9414 (N_9414,N_9382,N_9384);
or U9415 (N_9415,N_9370,N_9224);
or U9416 (N_9416,N_9385,N_9360);
and U9417 (N_9417,N_9363,N_9394);
or U9418 (N_9418,N_9351,N_9345);
nor U9419 (N_9419,N_9310,N_9248);
nor U9420 (N_9420,N_9344,N_9259);
nand U9421 (N_9421,N_9380,N_9247);
nor U9422 (N_9422,N_9228,N_9230);
and U9423 (N_9423,N_9294,N_9261);
nand U9424 (N_9424,N_9361,N_9319);
or U9425 (N_9425,N_9256,N_9304);
and U9426 (N_9426,N_9292,N_9368);
nand U9427 (N_9427,N_9376,N_9398);
nand U9428 (N_9428,N_9221,N_9373);
nor U9429 (N_9429,N_9348,N_9306);
or U9430 (N_9430,N_9378,N_9298);
or U9431 (N_9431,N_9202,N_9372);
nor U9432 (N_9432,N_9263,N_9320);
nor U9433 (N_9433,N_9393,N_9207);
or U9434 (N_9434,N_9383,N_9270);
nand U9435 (N_9435,N_9302,N_9227);
and U9436 (N_9436,N_9331,N_9214);
xnor U9437 (N_9437,N_9333,N_9239);
nor U9438 (N_9438,N_9281,N_9279);
nand U9439 (N_9439,N_9201,N_9366);
xor U9440 (N_9440,N_9397,N_9211);
or U9441 (N_9441,N_9286,N_9290);
nor U9442 (N_9442,N_9229,N_9388);
or U9443 (N_9443,N_9208,N_9346);
nor U9444 (N_9444,N_9357,N_9359);
nor U9445 (N_9445,N_9377,N_9299);
nand U9446 (N_9446,N_9350,N_9343);
nand U9447 (N_9447,N_9204,N_9317);
nand U9448 (N_9448,N_9213,N_9246);
or U9449 (N_9449,N_9234,N_9347);
nor U9450 (N_9450,N_9210,N_9289);
and U9451 (N_9451,N_9355,N_9280);
or U9452 (N_9452,N_9297,N_9291);
or U9453 (N_9453,N_9309,N_9392);
nand U9454 (N_9454,N_9271,N_9244);
nand U9455 (N_9455,N_9240,N_9338);
or U9456 (N_9456,N_9251,N_9243);
nor U9457 (N_9457,N_9264,N_9369);
nand U9458 (N_9458,N_9362,N_9287);
nor U9459 (N_9459,N_9301,N_9257);
or U9460 (N_9460,N_9295,N_9283);
or U9461 (N_9461,N_9332,N_9216);
or U9462 (N_9462,N_9335,N_9220);
and U9463 (N_9463,N_9250,N_9399);
or U9464 (N_9464,N_9318,N_9305);
xor U9465 (N_9465,N_9381,N_9334);
and U9466 (N_9466,N_9209,N_9265);
or U9467 (N_9467,N_9272,N_9222);
or U9468 (N_9468,N_9203,N_9307);
xnor U9469 (N_9469,N_9349,N_9323);
and U9470 (N_9470,N_9330,N_9321);
nand U9471 (N_9471,N_9358,N_9245);
xnor U9472 (N_9472,N_9277,N_9303);
nand U9473 (N_9473,N_9371,N_9225);
xor U9474 (N_9474,N_9206,N_9215);
nand U9475 (N_9475,N_9328,N_9293);
nand U9476 (N_9476,N_9312,N_9217);
xnor U9477 (N_9477,N_9282,N_9242);
nor U9478 (N_9478,N_9288,N_9253);
or U9479 (N_9479,N_9238,N_9223);
nand U9480 (N_9480,N_9274,N_9268);
nand U9481 (N_9481,N_9341,N_9390);
or U9482 (N_9482,N_9374,N_9296);
or U9483 (N_9483,N_9252,N_9218);
nand U9484 (N_9484,N_9337,N_9379);
nor U9485 (N_9485,N_9276,N_9205);
and U9486 (N_9486,N_9336,N_9311);
xnor U9487 (N_9487,N_9322,N_9278);
or U9488 (N_9488,N_9364,N_9262);
xor U9489 (N_9489,N_9389,N_9237);
nand U9490 (N_9490,N_9340,N_9342);
or U9491 (N_9491,N_9254,N_9258);
and U9492 (N_9492,N_9275,N_9236);
xor U9493 (N_9493,N_9375,N_9313);
nand U9494 (N_9494,N_9353,N_9324);
xor U9495 (N_9495,N_9315,N_9255);
nor U9496 (N_9496,N_9316,N_9396);
and U9497 (N_9497,N_9267,N_9314);
xnor U9498 (N_9498,N_9233,N_9391);
nor U9499 (N_9499,N_9219,N_9232);
xnor U9500 (N_9500,N_9243,N_9254);
nand U9501 (N_9501,N_9358,N_9373);
xnor U9502 (N_9502,N_9233,N_9354);
or U9503 (N_9503,N_9272,N_9353);
nand U9504 (N_9504,N_9313,N_9243);
or U9505 (N_9505,N_9320,N_9397);
nor U9506 (N_9506,N_9223,N_9395);
and U9507 (N_9507,N_9249,N_9377);
and U9508 (N_9508,N_9317,N_9344);
nor U9509 (N_9509,N_9215,N_9241);
xor U9510 (N_9510,N_9212,N_9276);
nor U9511 (N_9511,N_9346,N_9342);
and U9512 (N_9512,N_9345,N_9360);
nand U9513 (N_9513,N_9315,N_9214);
xnor U9514 (N_9514,N_9252,N_9330);
or U9515 (N_9515,N_9332,N_9377);
or U9516 (N_9516,N_9388,N_9363);
xnor U9517 (N_9517,N_9387,N_9339);
nor U9518 (N_9518,N_9251,N_9228);
and U9519 (N_9519,N_9319,N_9390);
nand U9520 (N_9520,N_9240,N_9268);
nor U9521 (N_9521,N_9352,N_9351);
and U9522 (N_9522,N_9248,N_9315);
nor U9523 (N_9523,N_9237,N_9333);
and U9524 (N_9524,N_9246,N_9375);
nor U9525 (N_9525,N_9385,N_9249);
and U9526 (N_9526,N_9389,N_9220);
xnor U9527 (N_9527,N_9347,N_9318);
or U9528 (N_9528,N_9217,N_9210);
nand U9529 (N_9529,N_9258,N_9324);
nor U9530 (N_9530,N_9293,N_9347);
and U9531 (N_9531,N_9229,N_9318);
or U9532 (N_9532,N_9372,N_9256);
and U9533 (N_9533,N_9369,N_9213);
xor U9534 (N_9534,N_9293,N_9397);
and U9535 (N_9535,N_9261,N_9284);
xor U9536 (N_9536,N_9275,N_9366);
and U9537 (N_9537,N_9340,N_9246);
or U9538 (N_9538,N_9235,N_9301);
xor U9539 (N_9539,N_9310,N_9335);
and U9540 (N_9540,N_9348,N_9245);
nor U9541 (N_9541,N_9225,N_9247);
xor U9542 (N_9542,N_9358,N_9336);
xnor U9543 (N_9543,N_9262,N_9299);
and U9544 (N_9544,N_9398,N_9390);
nor U9545 (N_9545,N_9261,N_9335);
and U9546 (N_9546,N_9304,N_9211);
nand U9547 (N_9547,N_9257,N_9380);
nand U9548 (N_9548,N_9368,N_9326);
nand U9549 (N_9549,N_9213,N_9209);
and U9550 (N_9550,N_9212,N_9229);
or U9551 (N_9551,N_9335,N_9327);
or U9552 (N_9552,N_9288,N_9356);
and U9553 (N_9553,N_9282,N_9287);
or U9554 (N_9554,N_9288,N_9273);
nand U9555 (N_9555,N_9384,N_9301);
nor U9556 (N_9556,N_9368,N_9282);
and U9557 (N_9557,N_9303,N_9312);
or U9558 (N_9558,N_9267,N_9283);
xnor U9559 (N_9559,N_9322,N_9223);
nor U9560 (N_9560,N_9213,N_9264);
nor U9561 (N_9561,N_9266,N_9201);
and U9562 (N_9562,N_9308,N_9370);
nand U9563 (N_9563,N_9359,N_9340);
nor U9564 (N_9564,N_9399,N_9327);
nand U9565 (N_9565,N_9327,N_9252);
or U9566 (N_9566,N_9269,N_9218);
nand U9567 (N_9567,N_9309,N_9301);
or U9568 (N_9568,N_9304,N_9227);
nor U9569 (N_9569,N_9290,N_9360);
and U9570 (N_9570,N_9233,N_9263);
or U9571 (N_9571,N_9208,N_9215);
and U9572 (N_9572,N_9308,N_9378);
xnor U9573 (N_9573,N_9282,N_9265);
xnor U9574 (N_9574,N_9270,N_9370);
and U9575 (N_9575,N_9204,N_9240);
and U9576 (N_9576,N_9348,N_9295);
or U9577 (N_9577,N_9227,N_9294);
or U9578 (N_9578,N_9330,N_9287);
nor U9579 (N_9579,N_9345,N_9336);
xor U9580 (N_9580,N_9272,N_9210);
or U9581 (N_9581,N_9283,N_9356);
nand U9582 (N_9582,N_9315,N_9247);
nor U9583 (N_9583,N_9261,N_9372);
or U9584 (N_9584,N_9243,N_9224);
xnor U9585 (N_9585,N_9241,N_9250);
xor U9586 (N_9586,N_9341,N_9395);
nor U9587 (N_9587,N_9360,N_9294);
or U9588 (N_9588,N_9376,N_9367);
or U9589 (N_9589,N_9386,N_9258);
and U9590 (N_9590,N_9237,N_9295);
and U9591 (N_9591,N_9377,N_9263);
nor U9592 (N_9592,N_9319,N_9318);
nor U9593 (N_9593,N_9214,N_9283);
and U9594 (N_9594,N_9226,N_9303);
nor U9595 (N_9595,N_9202,N_9294);
xnor U9596 (N_9596,N_9245,N_9251);
nand U9597 (N_9597,N_9207,N_9304);
xor U9598 (N_9598,N_9248,N_9201);
or U9599 (N_9599,N_9376,N_9399);
nand U9600 (N_9600,N_9558,N_9447);
xor U9601 (N_9601,N_9407,N_9534);
and U9602 (N_9602,N_9441,N_9414);
nor U9603 (N_9603,N_9461,N_9579);
nand U9604 (N_9604,N_9499,N_9425);
or U9605 (N_9605,N_9501,N_9521);
nand U9606 (N_9606,N_9446,N_9436);
and U9607 (N_9607,N_9475,N_9406);
xnor U9608 (N_9608,N_9575,N_9493);
xnor U9609 (N_9609,N_9474,N_9549);
nand U9610 (N_9610,N_9566,N_9463);
nor U9611 (N_9611,N_9427,N_9513);
or U9612 (N_9612,N_9535,N_9443);
or U9613 (N_9613,N_9538,N_9510);
nand U9614 (N_9614,N_9401,N_9458);
or U9615 (N_9615,N_9484,N_9413);
nor U9616 (N_9616,N_9551,N_9487);
and U9617 (N_9617,N_9462,N_9528);
or U9618 (N_9618,N_9509,N_9404);
nor U9619 (N_9619,N_9418,N_9589);
and U9620 (N_9620,N_9573,N_9564);
or U9621 (N_9621,N_9569,N_9502);
nand U9622 (N_9622,N_9586,N_9400);
or U9623 (N_9623,N_9433,N_9592);
nor U9624 (N_9624,N_9581,N_9587);
nand U9625 (N_9625,N_9578,N_9491);
xor U9626 (N_9626,N_9561,N_9431);
nand U9627 (N_9627,N_9480,N_9449);
nand U9628 (N_9628,N_9426,N_9559);
nor U9629 (N_9629,N_9460,N_9405);
nand U9630 (N_9630,N_9503,N_9428);
xnor U9631 (N_9631,N_9434,N_9507);
xor U9632 (N_9632,N_9500,N_9488);
nor U9633 (N_9633,N_9508,N_9523);
nand U9634 (N_9634,N_9504,N_9497);
nand U9635 (N_9635,N_9481,N_9553);
nand U9636 (N_9636,N_9454,N_9547);
and U9637 (N_9637,N_9542,N_9482);
xnor U9638 (N_9638,N_9483,N_9471);
or U9639 (N_9639,N_9448,N_9479);
xor U9640 (N_9640,N_9432,N_9469);
or U9641 (N_9641,N_9596,N_9512);
and U9642 (N_9642,N_9537,N_9554);
xnor U9643 (N_9643,N_9598,N_9456);
and U9644 (N_9644,N_9533,N_9473);
nor U9645 (N_9645,N_9459,N_9560);
xnor U9646 (N_9646,N_9588,N_9595);
or U9647 (N_9647,N_9444,N_9416);
nor U9648 (N_9648,N_9563,N_9593);
nor U9649 (N_9649,N_9437,N_9530);
and U9650 (N_9650,N_9402,N_9590);
nand U9651 (N_9651,N_9464,N_9498);
xnor U9652 (N_9652,N_9457,N_9529);
or U9653 (N_9653,N_9516,N_9570);
nor U9654 (N_9654,N_9415,N_9477);
nor U9655 (N_9655,N_9545,N_9571);
and U9656 (N_9656,N_9557,N_9411);
nand U9657 (N_9657,N_9518,N_9453);
and U9658 (N_9658,N_9429,N_9438);
xor U9659 (N_9659,N_9472,N_9582);
xor U9660 (N_9660,N_9543,N_9532);
or U9661 (N_9661,N_9562,N_9580);
and U9662 (N_9662,N_9597,N_9565);
nand U9663 (N_9663,N_9568,N_9591);
and U9664 (N_9664,N_9594,N_9511);
or U9665 (N_9665,N_9408,N_9490);
nor U9666 (N_9666,N_9478,N_9419);
nor U9667 (N_9667,N_9476,N_9525);
or U9668 (N_9668,N_9599,N_9495);
nand U9669 (N_9669,N_9515,N_9423);
and U9670 (N_9670,N_9465,N_9576);
xor U9671 (N_9671,N_9496,N_9584);
xor U9672 (N_9672,N_9524,N_9485);
and U9673 (N_9673,N_9522,N_9410);
and U9674 (N_9674,N_9550,N_9536);
nor U9675 (N_9675,N_9424,N_9556);
or U9676 (N_9676,N_9422,N_9466);
xnor U9677 (N_9677,N_9527,N_9430);
nand U9678 (N_9678,N_9555,N_9583);
and U9679 (N_9679,N_9574,N_9468);
nor U9680 (N_9680,N_9409,N_9412);
nor U9681 (N_9681,N_9452,N_9505);
nor U9682 (N_9682,N_9403,N_9417);
xor U9683 (N_9683,N_9520,N_9577);
xor U9684 (N_9684,N_9439,N_9489);
and U9685 (N_9685,N_9450,N_9445);
nand U9686 (N_9686,N_9552,N_9585);
and U9687 (N_9687,N_9531,N_9494);
or U9688 (N_9688,N_9420,N_9540);
and U9689 (N_9689,N_9435,N_9572);
or U9690 (N_9690,N_9517,N_9526);
nor U9691 (N_9691,N_9492,N_9455);
or U9692 (N_9692,N_9442,N_9514);
nor U9693 (N_9693,N_9440,N_9539);
xnor U9694 (N_9694,N_9467,N_9470);
and U9695 (N_9695,N_9519,N_9567);
or U9696 (N_9696,N_9541,N_9546);
xnor U9697 (N_9697,N_9544,N_9451);
nor U9698 (N_9698,N_9421,N_9486);
xnor U9699 (N_9699,N_9506,N_9548);
or U9700 (N_9700,N_9408,N_9498);
and U9701 (N_9701,N_9523,N_9505);
xor U9702 (N_9702,N_9445,N_9539);
xor U9703 (N_9703,N_9433,N_9589);
xnor U9704 (N_9704,N_9413,N_9424);
nand U9705 (N_9705,N_9401,N_9492);
nor U9706 (N_9706,N_9581,N_9565);
nor U9707 (N_9707,N_9436,N_9424);
nand U9708 (N_9708,N_9553,N_9467);
and U9709 (N_9709,N_9493,N_9485);
xnor U9710 (N_9710,N_9459,N_9586);
nor U9711 (N_9711,N_9595,N_9529);
nand U9712 (N_9712,N_9597,N_9581);
and U9713 (N_9713,N_9427,N_9432);
nand U9714 (N_9714,N_9423,N_9412);
nor U9715 (N_9715,N_9466,N_9582);
and U9716 (N_9716,N_9415,N_9513);
xnor U9717 (N_9717,N_9505,N_9481);
nor U9718 (N_9718,N_9507,N_9469);
or U9719 (N_9719,N_9418,N_9598);
and U9720 (N_9720,N_9500,N_9539);
nor U9721 (N_9721,N_9433,N_9437);
or U9722 (N_9722,N_9548,N_9543);
nor U9723 (N_9723,N_9596,N_9493);
xnor U9724 (N_9724,N_9566,N_9576);
nand U9725 (N_9725,N_9551,N_9517);
or U9726 (N_9726,N_9457,N_9463);
nand U9727 (N_9727,N_9410,N_9562);
or U9728 (N_9728,N_9503,N_9516);
or U9729 (N_9729,N_9490,N_9567);
nor U9730 (N_9730,N_9520,N_9448);
and U9731 (N_9731,N_9496,N_9571);
nand U9732 (N_9732,N_9492,N_9410);
nor U9733 (N_9733,N_9467,N_9528);
nor U9734 (N_9734,N_9485,N_9510);
nand U9735 (N_9735,N_9510,N_9400);
nor U9736 (N_9736,N_9524,N_9417);
or U9737 (N_9737,N_9517,N_9455);
nand U9738 (N_9738,N_9514,N_9512);
nor U9739 (N_9739,N_9527,N_9409);
xor U9740 (N_9740,N_9504,N_9537);
nor U9741 (N_9741,N_9473,N_9440);
or U9742 (N_9742,N_9519,N_9471);
and U9743 (N_9743,N_9570,N_9585);
xnor U9744 (N_9744,N_9512,N_9517);
xnor U9745 (N_9745,N_9534,N_9536);
or U9746 (N_9746,N_9447,N_9488);
or U9747 (N_9747,N_9485,N_9437);
nand U9748 (N_9748,N_9584,N_9497);
and U9749 (N_9749,N_9542,N_9416);
xnor U9750 (N_9750,N_9417,N_9480);
nor U9751 (N_9751,N_9516,N_9457);
and U9752 (N_9752,N_9524,N_9542);
xor U9753 (N_9753,N_9549,N_9466);
nor U9754 (N_9754,N_9461,N_9505);
xor U9755 (N_9755,N_9590,N_9548);
nand U9756 (N_9756,N_9549,N_9542);
nand U9757 (N_9757,N_9584,N_9434);
nor U9758 (N_9758,N_9535,N_9538);
or U9759 (N_9759,N_9556,N_9578);
and U9760 (N_9760,N_9457,N_9449);
nor U9761 (N_9761,N_9464,N_9435);
and U9762 (N_9762,N_9519,N_9407);
nand U9763 (N_9763,N_9516,N_9588);
xnor U9764 (N_9764,N_9591,N_9422);
nor U9765 (N_9765,N_9443,N_9447);
and U9766 (N_9766,N_9507,N_9568);
nor U9767 (N_9767,N_9532,N_9503);
or U9768 (N_9768,N_9472,N_9455);
nor U9769 (N_9769,N_9513,N_9504);
or U9770 (N_9770,N_9400,N_9419);
nand U9771 (N_9771,N_9534,N_9525);
nor U9772 (N_9772,N_9493,N_9567);
nor U9773 (N_9773,N_9546,N_9537);
and U9774 (N_9774,N_9589,N_9574);
and U9775 (N_9775,N_9451,N_9460);
xnor U9776 (N_9776,N_9467,N_9479);
or U9777 (N_9777,N_9469,N_9595);
nor U9778 (N_9778,N_9565,N_9418);
or U9779 (N_9779,N_9460,N_9539);
or U9780 (N_9780,N_9406,N_9593);
nand U9781 (N_9781,N_9444,N_9479);
nor U9782 (N_9782,N_9468,N_9533);
and U9783 (N_9783,N_9434,N_9404);
nand U9784 (N_9784,N_9416,N_9521);
xnor U9785 (N_9785,N_9411,N_9591);
nor U9786 (N_9786,N_9580,N_9552);
xor U9787 (N_9787,N_9436,N_9547);
and U9788 (N_9788,N_9506,N_9509);
xor U9789 (N_9789,N_9570,N_9568);
xnor U9790 (N_9790,N_9586,N_9483);
nor U9791 (N_9791,N_9470,N_9581);
xnor U9792 (N_9792,N_9549,N_9510);
xnor U9793 (N_9793,N_9588,N_9582);
nand U9794 (N_9794,N_9416,N_9510);
nand U9795 (N_9795,N_9501,N_9435);
nor U9796 (N_9796,N_9572,N_9574);
or U9797 (N_9797,N_9412,N_9419);
nand U9798 (N_9798,N_9567,N_9553);
and U9799 (N_9799,N_9497,N_9569);
or U9800 (N_9800,N_9792,N_9764);
nor U9801 (N_9801,N_9745,N_9645);
nand U9802 (N_9802,N_9607,N_9760);
or U9803 (N_9803,N_9650,N_9746);
nor U9804 (N_9804,N_9710,N_9732);
xor U9805 (N_9805,N_9711,N_9608);
and U9806 (N_9806,N_9601,N_9680);
and U9807 (N_9807,N_9664,N_9653);
and U9808 (N_9808,N_9733,N_9708);
and U9809 (N_9809,N_9610,N_9699);
xnor U9810 (N_9810,N_9744,N_9755);
nor U9811 (N_9811,N_9621,N_9788);
or U9812 (N_9812,N_9790,N_9615);
and U9813 (N_9813,N_9696,N_9604);
and U9814 (N_9814,N_9759,N_9751);
nand U9815 (N_9815,N_9712,N_9734);
nand U9816 (N_9816,N_9725,N_9706);
and U9817 (N_9817,N_9781,N_9637);
and U9818 (N_9818,N_9667,N_9682);
nor U9819 (N_9819,N_9616,N_9747);
or U9820 (N_9820,N_9627,N_9662);
nand U9821 (N_9821,N_9721,N_9668);
nand U9822 (N_9822,N_9756,N_9773);
xor U9823 (N_9823,N_9758,N_9681);
nand U9824 (N_9824,N_9738,N_9688);
nor U9825 (N_9825,N_9737,N_9705);
or U9826 (N_9826,N_9686,N_9740);
nor U9827 (N_9827,N_9613,N_9789);
or U9828 (N_9828,N_9640,N_9634);
and U9829 (N_9829,N_9735,N_9641);
nor U9830 (N_9830,N_9619,N_9612);
nor U9831 (N_9831,N_9643,N_9633);
nor U9832 (N_9832,N_9769,N_9661);
and U9833 (N_9833,N_9693,N_9635);
nand U9834 (N_9834,N_9652,N_9656);
nand U9835 (N_9835,N_9793,N_9690);
xnor U9836 (N_9836,N_9786,N_9692);
and U9837 (N_9837,N_9685,N_9605);
nor U9838 (N_9838,N_9767,N_9753);
nor U9839 (N_9839,N_9600,N_9603);
and U9840 (N_9840,N_9739,N_9624);
nor U9841 (N_9841,N_9724,N_9632);
nor U9842 (N_9842,N_9776,N_9784);
and U9843 (N_9843,N_9674,N_9727);
nand U9844 (N_9844,N_9614,N_9799);
nor U9845 (N_9845,N_9684,N_9660);
xor U9846 (N_9846,N_9715,N_9741);
xnor U9847 (N_9847,N_9774,N_9642);
and U9848 (N_9848,N_9683,N_9709);
nand U9849 (N_9849,N_9698,N_9625);
or U9850 (N_9850,N_9730,N_9630);
and U9851 (N_9851,N_9602,N_9761);
nor U9852 (N_9852,N_9676,N_9798);
nor U9853 (N_9853,N_9765,N_9731);
nor U9854 (N_9854,N_9678,N_9718);
nor U9855 (N_9855,N_9677,N_9729);
and U9856 (N_9856,N_9675,N_9611);
xnor U9857 (N_9857,N_9754,N_9763);
xnor U9858 (N_9858,N_9750,N_9639);
or U9859 (N_9859,N_9782,N_9651);
or U9860 (N_9860,N_9772,N_9778);
and U9861 (N_9861,N_9771,N_9654);
xnor U9862 (N_9862,N_9702,N_9636);
or U9863 (N_9863,N_9762,N_9757);
nand U9864 (N_9864,N_9794,N_9779);
nor U9865 (N_9865,N_9797,N_9671);
nor U9866 (N_9866,N_9701,N_9673);
xnor U9867 (N_9867,N_9655,N_9687);
xnor U9868 (N_9868,N_9623,N_9626);
and U9869 (N_9869,N_9722,N_9638);
xor U9870 (N_9870,N_9736,N_9666);
nand U9871 (N_9871,N_9795,N_9659);
or U9872 (N_9872,N_9665,N_9728);
nand U9873 (N_9873,N_9628,N_9663);
and U9874 (N_9874,N_9694,N_9689);
or U9875 (N_9875,N_9629,N_9691);
nand U9876 (N_9876,N_9720,N_9669);
or U9877 (N_9877,N_9657,N_9726);
nor U9878 (N_9878,N_9777,N_9714);
xor U9879 (N_9879,N_9785,N_9697);
or U9880 (N_9880,N_9704,N_9748);
or U9881 (N_9881,N_9719,N_9713);
nor U9882 (N_9882,N_9783,N_9707);
or U9883 (N_9883,N_9618,N_9617);
nor U9884 (N_9884,N_9695,N_9749);
nor U9885 (N_9885,N_9700,N_9770);
and U9886 (N_9886,N_9703,N_9743);
nand U9887 (N_9887,N_9791,N_9716);
nor U9888 (N_9888,N_9670,N_9658);
and U9889 (N_9889,N_9646,N_9672);
or U9890 (N_9890,N_9766,N_9609);
nor U9891 (N_9891,N_9717,N_9649);
nor U9892 (N_9892,N_9679,N_9796);
nor U9893 (N_9893,N_9606,N_9787);
or U9894 (N_9894,N_9780,N_9620);
and U9895 (N_9895,N_9631,N_9742);
and U9896 (N_9896,N_9723,N_9752);
or U9897 (N_9897,N_9622,N_9648);
nor U9898 (N_9898,N_9644,N_9768);
xor U9899 (N_9899,N_9647,N_9775);
nor U9900 (N_9900,N_9643,N_9698);
nand U9901 (N_9901,N_9723,N_9656);
and U9902 (N_9902,N_9778,N_9744);
xnor U9903 (N_9903,N_9693,N_9720);
or U9904 (N_9904,N_9759,N_9747);
nand U9905 (N_9905,N_9771,N_9702);
xor U9906 (N_9906,N_9670,N_9710);
xnor U9907 (N_9907,N_9780,N_9774);
xor U9908 (N_9908,N_9695,N_9789);
or U9909 (N_9909,N_9766,N_9789);
nor U9910 (N_9910,N_9758,N_9648);
or U9911 (N_9911,N_9688,N_9600);
or U9912 (N_9912,N_9622,N_9609);
or U9913 (N_9913,N_9762,N_9626);
nor U9914 (N_9914,N_9711,N_9686);
or U9915 (N_9915,N_9769,N_9717);
and U9916 (N_9916,N_9644,N_9706);
and U9917 (N_9917,N_9751,N_9710);
or U9918 (N_9918,N_9647,N_9631);
xnor U9919 (N_9919,N_9651,N_9634);
nor U9920 (N_9920,N_9641,N_9741);
or U9921 (N_9921,N_9720,N_9792);
xnor U9922 (N_9922,N_9702,N_9693);
nand U9923 (N_9923,N_9754,N_9687);
xor U9924 (N_9924,N_9637,N_9676);
or U9925 (N_9925,N_9773,N_9625);
and U9926 (N_9926,N_9708,N_9726);
and U9927 (N_9927,N_9785,N_9654);
nand U9928 (N_9928,N_9748,N_9658);
or U9929 (N_9929,N_9651,N_9710);
and U9930 (N_9930,N_9730,N_9695);
nor U9931 (N_9931,N_9606,N_9717);
nand U9932 (N_9932,N_9643,N_9731);
and U9933 (N_9933,N_9672,N_9602);
and U9934 (N_9934,N_9745,N_9668);
and U9935 (N_9935,N_9600,N_9713);
and U9936 (N_9936,N_9617,N_9767);
and U9937 (N_9937,N_9639,N_9731);
nand U9938 (N_9938,N_9725,N_9729);
nor U9939 (N_9939,N_9657,N_9618);
and U9940 (N_9940,N_9614,N_9620);
nor U9941 (N_9941,N_9692,N_9774);
nand U9942 (N_9942,N_9775,N_9780);
xor U9943 (N_9943,N_9793,N_9656);
or U9944 (N_9944,N_9619,N_9622);
nand U9945 (N_9945,N_9631,N_9760);
nand U9946 (N_9946,N_9782,N_9643);
or U9947 (N_9947,N_9783,N_9648);
xnor U9948 (N_9948,N_9611,N_9760);
nor U9949 (N_9949,N_9769,N_9609);
or U9950 (N_9950,N_9749,N_9765);
and U9951 (N_9951,N_9782,N_9683);
nand U9952 (N_9952,N_9687,N_9658);
nor U9953 (N_9953,N_9656,N_9621);
or U9954 (N_9954,N_9745,N_9600);
xnor U9955 (N_9955,N_9664,N_9735);
nor U9956 (N_9956,N_9706,N_9705);
xnor U9957 (N_9957,N_9734,N_9787);
and U9958 (N_9958,N_9737,N_9729);
nand U9959 (N_9959,N_9773,N_9790);
or U9960 (N_9960,N_9783,N_9797);
and U9961 (N_9961,N_9799,N_9693);
xnor U9962 (N_9962,N_9687,N_9688);
or U9963 (N_9963,N_9796,N_9715);
xnor U9964 (N_9964,N_9631,N_9663);
xor U9965 (N_9965,N_9689,N_9757);
or U9966 (N_9966,N_9727,N_9782);
xnor U9967 (N_9967,N_9776,N_9612);
nor U9968 (N_9968,N_9624,N_9615);
xor U9969 (N_9969,N_9722,N_9765);
and U9970 (N_9970,N_9741,N_9675);
or U9971 (N_9971,N_9622,N_9799);
nand U9972 (N_9972,N_9708,N_9799);
and U9973 (N_9973,N_9766,N_9749);
or U9974 (N_9974,N_9689,N_9620);
or U9975 (N_9975,N_9733,N_9723);
nor U9976 (N_9976,N_9605,N_9630);
or U9977 (N_9977,N_9661,N_9686);
nor U9978 (N_9978,N_9772,N_9642);
xor U9979 (N_9979,N_9616,N_9629);
nand U9980 (N_9980,N_9716,N_9666);
nor U9981 (N_9981,N_9613,N_9780);
nand U9982 (N_9982,N_9686,N_9660);
xnor U9983 (N_9983,N_9731,N_9718);
nand U9984 (N_9984,N_9601,N_9731);
and U9985 (N_9985,N_9635,N_9645);
nor U9986 (N_9986,N_9743,N_9608);
or U9987 (N_9987,N_9653,N_9774);
or U9988 (N_9988,N_9610,N_9659);
or U9989 (N_9989,N_9786,N_9666);
nor U9990 (N_9990,N_9708,N_9784);
or U9991 (N_9991,N_9676,N_9642);
nor U9992 (N_9992,N_9632,N_9716);
nor U9993 (N_9993,N_9704,N_9662);
xor U9994 (N_9994,N_9636,N_9674);
nand U9995 (N_9995,N_9626,N_9697);
nand U9996 (N_9996,N_9692,N_9643);
nor U9997 (N_9997,N_9782,N_9698);
nor U9998 (N_9998,N_9692,N_9731);
nor U9999 (N_9999,N_9638,N_9639);
nor U10000 (N_10000,N_9929,N_9816);
or U10001 (N_10001,N_9825,N_9931);
nor U10002 (N_10002,N_9801,N_9815);
xor U10003 (N_10003,N_9885,N_9987);
and U10004 (N_10004,N_9813,N_9973);
xnor U10005 (N_10005,N_9865,N_9912);
and U10006 (N_10006,N_9952,N_9978);
xor U10007 (N_10007,N_9947,N_9823);
or U10008 (N_10008,N_9842,N_9872);
nor U10009 (N_10009,N_9868,N_9869);
xor U10010 (N_10010,N_9806,N_9986);
and U10011 (N_10011,N_9915,N_9976);
or U10012 (N_10012,N_9920,N_9911);
nand U10013 (N_10013,N_9817,N_9848);
or U10014 (N_10014,N_9910,N_9961);
xnor U10015 (N_10015,N_9821,N_9950);
xnor U10016 (N_10016,N_9901,N_9831);
xnor U10017 (N_10017,N_9836,N_9875);
nand U10018 (N_10018,N_9991,N_9917);
nor U10019 (N_10019,N_9919,N_9838);
or U10020 (N_10020,N_9894,N_9803);
xnor U10021 (N_10021,N_9932,N_9877);
and U10022 (N_10022,N_9982,N_9841);
or U10023 (N_10023,N_9851,N_9804);
xor U10024 (N_10024,N_9940,N_9936);
nand U10025 (N_10025,N_9914,N_9994);
nor U10026 (N_10026,N_9913,N_9941);
xor U10027 (N_10027,N_9923,N_9992);
and U10028 (N_10028,N_9820,N_9907);
and U10029 (N_10029,N_9918,N_9857);
nand U10030 (N_10030,N_9988,N_9967);
nand U10031 (N_10031,N_9984,N_9863);
nand U10032 (N_10032,N_9859,N_9899);
xnor U10033 (N_10033,N_9945,N_9873);
or U10034 (N_10034,N_9985,N_9926);
and U10035 (N_10035,N_9951,N_9802);
nor U10036 (N_10036,N_9828,N_9965);
or U10037 (N_10037,N_9960,N_9898);
nor U10038 (N_10038,N_9997,N_9959);
and U10039 (N_10039,N_9856,N_9916);
nand U10040 (N_10040,N_9888,N_9900);
or U10041 (N_10041,N_9963,N_9822);
or U10042 (N_10042,N_9843,N_9981);
xor U10043 (N_10043,N_9924,N_9890);
nor U10044 (N_10044,N_9904,N_9860);
nor U10045 (N_10045,N_9834,N_9905);
and U10046 (N_10046,N_9895,N_9939);
and U10047 (N_10047,N_9812,N_9922);
and U10048 (N_10048,N_9927,N_9990);
nand U10049 (N_10049,N_9980,N_9808);
xor U10050 (N_10050,N_9897,N_9896);
or U10051 (N_10051,N_9955,N_9845);
and U10052 (N_10052,N_9884,N_9977);
nand U10053 (N_10053,N_9809,N_9824);
xnor U10054 (N_10054,N_9906,N_9953);
nor U10055 (N_10055,N_9948,N_9878);
and U10056 (N_10056,N_9861,N_9935);
and U10057 (N_10057,N_9930,N_9983);
and U10058 (N_10058,N_9956,N_9807);
or U10059 (N_10059,N_9864,N_9946);
nor U10060 (N_10060,N_9852,N_9979);
nor U10061 (N_10061,N_9902,N_9829);
nand U10062 (N_10062,N_9954,N_9969);
and U10063 (N_10063,N_9847,N_9810);
and U10064 (N_10064,N_9943,N_9995);
and U10065 (N_10065,N_9974,N_9964);
nand U10066 (N_10066,N_9993,N_9826);
or U10067 (N_10067,N_9949,N_9866);
nand U10068 (N_10068,N_9999,N_9887);
nor U10069 (N_10069,N_9921,N_9933);
nor U10070 (N_10070,N_9958,N_9942);
or U10071 (N_10071,N_9862,N_9934);
nand U10072 (N_10072,N_9800,N_9938);
or U10073 (N_10073,N_9854,N_9879);
nand U10074 (N_10074,N_9819,N_9883);
and U10075 (N_10075,N_9839,N_9962);
and U10076 (N_10076,N_9892,N_9996);
nand U10077 (N_10077,N_9840,N_9876);
and U10078 (N_10078,N_9889,N_9814);
and U10079 (N_10079,N_9966,N_9827);
nor U10080 (N_10080,N_9849,N_9850);
or U10081 (N_10081,N_9909,N_9805);
nor U10082 (N_10082,N_9870,N_9833);
xor U10083 (N_10083,N_9972,N_9832);
nand U10084 (N_10084,N_9989,N_9925);
nand U10085 (N_10085,N_9844,N_9871);
and U10086 (N_10086,N_9881,N_9971);
xnor U10087 (N_10087,N_9893,N_9830);
or U10088 (N_10088,N_9835,N_9886);
and U10089 (N_10089,N_9968,N_9855);
or U10090 (N_10090,N_9944,N_9957);
and U10091 (N_10091,N_9837,N_9874);
nand U10092 (N_10092,N_9975,N_9880);
and U10093 (N_10093,N_9882,N_9846);
or U10094 (N_10094,N_9811,N_9998);
and U10095 (N_10095,N_9903,N_9858);
nand U10096 (N_10096,N_9818,N_9891);
xor U10097 (N_10097,N_9867,N_9970);
nand U10098 (N_10098,N_9908,N_9853);
and U10099 (N_10099,N_9937,N_9928);
xor U10100 (N_10100,N_9912,N_9908);
nor U10101 (N_10101,N_9894,N_9838);
or U10102 (N_10102,N_9819,N_9901);
nor U10103 (N_10103,N_9976,N_9972);
nand U10104 (N_10104,N_9988,N_9915);
nand U10105 (N_10105,N_9933,N_9892);
nand U10106 (N_10106,N_9991,N_9939);
or U10107 (N_10107,N_9985,N_9853);
xor U10108 (N_10108,N_9895,N_9874);
or U10109 (N_10109,N_9867,N_9882);
nor U10110 (N_10110,N_9926,N_9955);
and U10111 (N_10111,N_9826,N_9807);
xor U10112 (N_10112,N_9948,N_9994);
nor U10113 (N_10113,N_9982,N_9826);
nor U10114 (N_10114,N_9967,N_9996);
and U10115 (N_10115,N_9891,N_9981);
nor U10116 (N_10116,N_9888,N_9816);
xnor U10117 (N_10117,N_9961,N_9897);
nor U10118 (N_10118,N_9844,N_9856);
or U10119 (N_10119,N_9816,N_9898);
nand U10120 (N_10120,N_9911,N_9866);
nor U10121 (N_10121,N_9935,N_9963);
or U10122 (N_10122,N_9891,N_9984);
nor U10123 (N_10123,N_9815,N_9982);
or U10124 (N_10124,N_9968,N_9999);
nor U10125 (N_10125,N_9861,N_9855);
xor U10126 (N_10126,N_9906,N_9842);
or U10127 (N_10127,N_9972,N_9993);
nor U10128 (N_10128,N_9823,N_9941);
nand U10129 (N_10129,N_9953,N_9946);
xor U10130 (N_10130,N_9819,N_9937);
xor U10131 (N_10131,N_9911,N_9951);
and U10132 (N_10132,N_9888,N_9832);
xor U10133 (N_10133,N_9858,N_9808);
or U10134 (N_10134,N_9935,N_9908);
nand U10135 (N_10135,N_9891,N_9945);
or U10136 (N_10136,N_9904,N_9880);
xor U10137 (N_10137,N_9992,N_9850);
nor U10138 (N_10138,N_9838,N_9885);
nor U10139 (N_10139,N_9973,N_9985);
or U10140 (N_10140,N_9802,N_9960);
or U10141 (N_10141,N_9889,N_9945);
nor U10142 (N_10142,N_9969,N_9837);
xor U10143 (N_10143,N_9898,N_9878);
xor U10144 (N_10144,N_9866,N_9881);
or U10145 (N_10145,N_9878,N_9924);
nor U10146 (N_10146,N_9891,N_9919);
and U10147 (N_10147,N_9951,N_9835);
nor U10148 (N_10148,N_9916,N_9843);
and U10149 (N_10149,N_9905,N_9966);
nand U10150 (N_10150,N_9858,N_9828);
xor U10151 (N_10151,N_9931,N_9866);
or U10152 (N_10152,N_9885,N_9825);
or U10153 (N_10153,N_9950,N_9979);
nor U10154 (N_10154,N_9938,N_9962);
xnor U10155 (N_10155,N_9886,N_9915);
nor U10156 (N_10156,N_9908,N_9901);
nand U10157 (N_10157,N_9817,N_9909);
nand U10158 (N_10158,N_9870,N_9903);
or U10159 (N_10159,N_9936,N_9882);
xor U10160 (N_10160,N_9840,N_9996);
nand U10161 (N_10161,N_9853,N_9873);
or U10162 (N_10162,N_9806,N_9890);
nand U10163 (N_10163,N_9833,N_9814);
and U10164 (N_10164,N_9906,N_9903);
and U10165 (N_10165,N_9949,N_9952);
xnor U10166 (N_10166,N_9972,N_9901);
and U10167 (N_10167,N_9984,N_9809);
or U10168 (N_10168,N_9939,N_9987);
or U10169 (N_10169,N_9976,N_9839);
nor U10170 (N_10170,N_9985,N_9852);
and U10171 (N_10171,N_9978,N_9971);
xnor U10172 (N_10172,N_9968,N_9948);
xnor U10173 (N_10173,N_9853,N_9807);
nor U10174 (N_10174,N_9959,N_9918);
xnor U10175 (N_10175,N_9800,N_9820);
or U10176 (N_10176,N_9951,N_9897);
xnor U10177 (N_10177,N_9969,N_9959);
and U10178 (N_10178,N_9892,N_9936);
nand U10179 (N_10179,N_9954,N_9943);
nor U10180 (N_10180,N_9971,N_9832);
and U10181 (N_10181,N_9840,N_9902);
nor U10182 (N_10182,N_9910,N_9856);
nor U10183 (N_10183,N_9946,N_9857);
nor U10184 (N_10184,N_9957,N_9869);
nor U10185 (N_10185,N_9809,N_9834);
nand U10186 (N_10186,N_9962,N_9998);
nand U10187 (N_10187,N_9903,N_9971);
and U10188 (N_10188,N_9829,N_9883);
xnor U10189 (N_10189,N_9908,N_9951);
xnor U10190 (N_10190,N_9807,N_9817);
or U10191 (N_10191,N_9853,N_9953);
and U10192 (N_10192,N_9961,N_9817);
nor U10193 (N_10193,N_9872,N_9843);
and U10194 (N_10194,N_9848,N_9951);
nand U10195 (N_10195,N_9864,N_9998);
and U10196 (N_10196,N_9803,N_9984);
nor U10197 (N_10197,N_9955,N_9910);
xor U10198 (N_10198,N_9889,N_9877);
xor U10199 (N_10199,N_9812,N_9823);
and U10200 (N_10200,N_10026,N_10195);
nor U10201 (N_10201,N_10177,N_10116);
or U10202 (N_10202,N_10197,N_10170);
nor U10203 (N_10203,N_10181,N_10131);
xnor U10204 (N_10204,N_10047,N_10183);
or U10205 (N_10205,N_10013,N_10049);
xnor U10206 (N_10206,N_10123,N_10067);
and U10207 (N_10207,N_10095,N_10097);
xor U10208 (N_10208,N_10021,N_10016);
nand U10209 (N_10209,N_10122,N_10008);
nand U10210 (N_10210,N_10165,N_10017);
and U10211 (N_10211,N_10088,N_10115);
and U10212 (N_10212,N_10023,N_10092);
nand U10213 (N_10213,N_10150,N_10168);
nand U10214 (N_10214,N_10127,N_10164);
nor U10215 (N_10215,N_10079,N_10101);
or U10216 (N_10216,N_10107,N_10100);
xor U10217 (N_10217,N_10153,N_10033);
xor U10218 (N_10218,N_10185,N_10069);
and U10219 (N_10219,N_10172,N_10178);
and U10220 (N_10220,N_10042,N_10176);
nor U10221 (N_10221,N_10158,N_10010);
or U10222 (N_10222,N_10137,N_10140);
nand U10223 (N_10223,N_10055,N_10082);
xnor U10224 (N_10224,N_10138,N_10161);
nor U10225 (N_10225,N_10083,N_10000);
and U10226 (N_10226,N_10139,N_10105);
or U10227 (N_10227,N_10040,N_10098);
and U10228 (N_10228,N_10077,N_10147);
nor U10229 (N_10229,N_10003,N_10070);
or U10230 (N_10230,N_10074,N_10086);
or U10231 (N_10231,N_10191,N_10006);
nor U10232 (N_10232,N_10112,N_10031);
or U10233 (N_10233,N_10059,N_10128);
and U10234 (N_10234,N_10125,N_10103);
nor U10235 (N_10235,N_10198,N_10136);
or U10236 (N_10236,N_10154,N_10130);
xor U10237 (N_10237,N_10096,N_10066);
or U10238 (N_10238,N_10048,N_10179);
xor U10239 (N_10239,N_10064,N_10155);
nand U10240 (N_10240,N_10029,N_10126);
nor U10241 (N_10241,N_10052,N_10051);
nor U10242 (N_10242,N_10002,N_10114);
nand U10243 (N_10243,N_10011,N_10044);
nand U10244 (N_10244,N_10143,N_10159);
xor U10245 (N_10245,N_10053,N_10027);
and U10246 (N_10246,N_10166,N_10032);
and U10247 (N_10247,N_10175,N_10078);
xor U10248 (N_10248,N_10057,N_10020);
xnor U10249 (N_10249,N_10144,N_10056);
xor U10250 (N_10250,N_10169,N_10072);
nor U10251 (N_10251,N_10121,N_10146);
xnor U10252 (N_10252,N_10180,N_10090);
or U10253 (N_10253,N_10073,N_10038);
nand U10254 (N_10254,N_10065,N_10174);
xnor U10255 (N_10255,N_10062,N_10124);
and U10256 (N_10256,N_10134,N_10156);
nand U10257 (N_10257,N_10080,N_10132);
and U10258 (N_10258,N_10068,N_10007);
or U10259 (N_10259,N_10054,N_10025);
or U10260 (N_10260,N_10199,N_10036);
or U10261 (N_10261,N_10012,N_10094);
nor U10262 (N_10262,N_10045,N_10093);
and U10263 (N_10263,N_10009,N_10087);
nor U10264 (N_10264,N_10084,N_10035);
or U10265 (N_10265,N_10163,N_10028);
and U10266 (N_10266,N_10050,N_10148);
and U10267 (N_10267,N_10110,N_10117);
and U10268 (N_10268,N_10160,N_10005);
xor U10269 (N_10269,N_10058,N_10129);
and U10270 (N_10270,N_10118,N_10142);
or U10271 (N_10271,N_10034,N_10106);
xor U10272 (N_10272,N_10119,N_10145);
xor U10273 (N_10273,N_10167,N_10184);
or U10274 (N_10274,N_10120,N_10018);
nor U10275 (N_10275,N_10063,N_10149);
nor U10276 (N_10276,N_10171,N_10060);
and U10277 (N_10277,N_10162,N_10141);
nor U10278 (N_10278,N_10151,N_10104);
nor U10279 (N_10279,N_10037,N_10173);
nand U10280 (N_10280,N_10061,N_10196);
xor U10281 (N_10281,N_10075,N_10019);
nor U10282 (N_10282,N_10015,N_10022);
or U10283 (N_10283,N_10111,N_10099);
nand U10284 (N_10284,N_10085,N_10041);
nor U10285 (N_10285,N_10135,N_10014);
nor U10286 (N_10286,N_10024,N_10113);
nor U10287 (N_10287,N_10189,N_10188);
and U10288 (N_10288,N_10186,N_10108);
xor U10289 (N_10289,N_10109,N_10192);
nor U10290 (N_10290,N_10102,N_10081);
xor U10291 (N_10291,N_10194,N_10193);
nand U10292 (N_10292,N_10043,N_10046);
xnor U10293 (N_10293,N_10091,N_10001);
nand U10294 (N_10294,N_10089,N_10039);
or U10295 (N_10295,N_10030,N_10182);
nand U10296 (N_10296,N_10190,N_10071);
and U10297 (N_10297,N_10004,N_10152);
and U10298 (N_10298,N_10076,N_10187);
nand U10299 (N_10299,N_10157,N_10133);
or U10300 (N_10300,N_10078,N_10012);
and U10301 (N_10301,N_10065,N_10169);
and U10302 (N_10302,N_10049,N_10156);
nor U10303 (N_10303,N_10111,N_10192);
or U10304 (N_10304,N_10022,N_10080);
nand U10305 (N_10305,N_10117,N_10039);
or U10306 (N_10306,N_10054,N_10105);
nand U10307 (N_10307,N_10050,N_10103);
nand U10308 (N_10308,N_10173,N_10043);
nand U10309 (N_10309,N_10016,N_10062);
nand U10310 (N_10310,N_10068,N_10011);
nand U10311 (N_10311,N_10131,N_10100);
xor U10312 (N_10312,N_10169,N_10101);
nor U10313 (N_10313,N_10044,N_10173);
nor U10314 (N_10314,N_10134,N_10150);
xnor U10315 (N_10315,N_10190,N_10055);
nor U10316 (N_10316,N_10176,N_10152);
nand U10317 (N_10317,N_10012,N_10070);
xnor U10318 (N_10318,N_10162,N_10183);
nor U10319 (N_10319,N_10087,N_10032);
nand U10320 (N_10320,N_10068,N_10117);
xnor U10321 (N_10321,N_10098,N_10034);
xor U10322 (N_10322,N_10004,N_10067);
nor U10323 (N_10323,N_10062,N_10169);
xnor U10324 (N_10324,N_10181,N_10110);
nor U10325 (N_10325,N_10175,N_10054);
and U10326 (N_10326,N_10058,N_10040);
nand U10327 (N_10327,N_10003,N_10048);
or U10328 (N_10328,N_10182,N_10004);
nand U10329 (N_10329,N_10140,N_10013);
xor U10330 (N_10330,N_10148,N_10164);
and U10331 (N_10331,N_10177,N_10122);
and U10332 (N_10332,N_10064,N_10154);
xor U10333 (N_10333,N_10121,N_10036);
and U10334 (N_10334,N_10105,N_10041);
nand U10335 (N_10335,N_10149,N_10114);
or U10336 (N_10336,N_10173,N_10108);
and U10337 (N_10337,N_10089,N_10163);
or U10338 (N_10338,N_10120,N_10021);
nand U10339 (N_10339,N_10091,N_10047);
nor U10340 (N_10340,N_10022,N_10053);
nor U10341 (N_10341,N_10198,N_10199);
xor U10342 (N_10342,N_10170,N_10036);
xor U10343 (N_10343,N_10091,N_10039);
xnor U10344 (N_10344,N_10191,N_10115);
xor U10345 (N_10345,N_10118,N_10049);
and U10346 (N_10346,N_10064,N_10194);
xor U10347 (N_10347,N_10127,N_10141);
xnor U10348 (N_10348,N_10157,N_10019);
nor U10349 (N_10349,N_10139,N_10122);
or U10350 (N_10350,N_10125,N_10017);
or U10351 (N_10351,N_10019,N_10149);
nand U10352 (N_10352,N_10094,N_10132);
xor U10353 (N_10353,N_10187,N_10167);
or U10354 (N_10354,N_10154,N_10133);
nor U10355 (N_10355,N_10173,N_10028);
xnor U10356 (N_10356,N_10001,N_10009);
or U10357 (N_10357,N_10002,N_10030);
nand U10358 (N_10358,N_10165,N_10038);
and U10359 (N_10359,N_10059,N_10022);
nor U10360 (N_10360,N_10022,N_10018);
or U10361 (N_10361,N_10021,N_10188);
nor U10362 (N_10362,N_10021,N_10191);
nand U10363 (N_10363,N_10079,N_10145);
nand U10364 (N_10364,N_10178,N_10121);
nor U10365 (N_10365,N_10149,N_10095);
nor U10366 (N_10366,N_10156,N_10017);
xnor U10367 (N_10367,N_10022,N_10098);
nand U10368 (N_10368,N_10093,N_10130);
nor U10369 (N_10369,N_10016,N_10035);
nand U10370 (N_10370,N_10079,N_10121);
xor U10371 (N_10371,N_10040,N_10008);
and U10372 (N_10372,N_10151,N_10046);
nor U10373 (N_10373,N_10090,N_10022);
or U10374 (N_10374,N_10096,N_10102);
or U10375 (N_10375,N_10178,N_10107);
or U10376 (N_10376,N_10080,N_10160);
or U10377 (N_10377,N_10103,N_10099);
and U10378 (N_10378,N_10158,N_10106);
and U10379 (N_10379,N_10003,N_10146);
xnor U10380 (N_10380,N_10079,N_10183);
nand U10381 (N_10381,N_10091,N_10038);
nor U10382 (N_10382,N_10027,N_10065);
nor U10383 (N_10383,N_10037,N_10069);
nor U10384 (N_10384,N_10107,N_10102);
xnor U10385 (N_10385,N_10075,N_10065);
or U10386 (N_10386,N_10097,N_10070);
nand U10387 (N_10387,N_10091,N_10062);
xor U10388 (N_10388,N_10042,N_10197);
nor U10389 (N_10389,N_10148,N_10192);
and U10390 (N_10390,N_10019,N_10159);
nand U10391 (N_10391,N_10022,N_10193);
or U10392 (N_10392,N_10082,N_10083);
xor U10393 (N_10393,N_10012,N_10188);
and U10394 (N_10394,N_10194,N_10124);
nand U10395 (N_10395,N_10173,N_10154);
nor U10396 (N_10396,N_10128,N_10036);
xor U10397 (N_10397,N_10049,N_10166);
nand U10398 (N_10398,N_10138,N_10180);
nand U10399 (N_10399,N_10108,N_10063);
nor U10400 (N_10400,N_10375,N_10380);
or U10401 (N_10401,N_10326,N_10363);
or U10402 (N_10402,N_10398,N_10301);
or U10403 (N_10403,N_10340,N_10306);
or U10404 (N_10404,N_10284,N_10245);
nand U10405 (N_10405,N_10236,N_10349);
nor U10406 (N_10406,N_10343,N_10342);
and U10407 (N_10407,N_10206,N_10378);
nand U10408 (N_10408,N_10290,N_10385);
nand U10409 (N_10409,N_10319,N_10270);
or U10410 (N_10410,N_10230,N_10285);
nor U10411 (N_10411,N_10280,N_10260);
xor U10412 (N_10412,N_10318,N_10391);
xor U10413 (N_10413,N_10209,N_10376);
or U10414 (N_10414,N_10242,N_10231);
or U10415 (N_10415,N_10365,N_10307);
and U10416 (N_10416,N_10327,N_10325);
xnor U10417 (N_10417,N_10238,N_10333);
and U10418 (N_10418,N_10395,N_10295);
xnor U10419 (N_10419,N_10292,N_10392);
xnor U10420 (N_10420,N_10399,N_10249);
nand U10421 (N_10421,N_10202,N_10294);
and U10422 (N_10422,N_10227,N_10369);
and U10423 (N_10423,N_10255,N_10210);
or U10424 (N_10424,N_10360,N_10220);
nand U10425 (N_10425,N_10311,N_10350);
and U10426 (N_10426,N_10314,N_10269);
or U10427 (N_10427,N_10348,N_10372);
or U10428 (N_10428,N_10339,N_10286);
nand U10429 (N_10429,N_10237,N_10213);
and U10430 (N_10430,N_10321,N_10346);
or U10431 (N_10431,N_10297,N_10323);
or U10432 (N_10432,N_10254,N_10276);
nand U10433 (N_10433,N_10259,N_10384);
nand U10434 (N_10434,N_10324,N_10267);
and U10435 (N_10435,N_10264,N_10257);
nor U10436 (N_10436,N_10338,N_10222);
and U10437 (N_10437,N_10396,N_10358);
nor U10438 (N_10438,N_10374,N_10345);
xor U10439 (N_10439,N_10312,N_10268);
or U10440 (N_10440,N_10386,N_10207);
xor U10441 (N_10441,N_10235,N_10214);
nor U10442 (N_10442,N_10383,N_10215);
nand U10443 (N_10443,N_10322,N_10313);
and U10444 (N_10444,N_10201,N_10250);
xor U10445 (N_10445,N_10351,N_10291);
nor U10446 (N_10446,N_10388,N_10357);
or U10447 (N_10447,N_10389,N_10379);
and U10448 (N_10448,N_10273,N_10226);
xor U10449 (N_10449,N_10356,N_10233);
and U10450 (N_10450,N_10223,N_10243);
nor U10451 (N_10451,N_10332,N_10211);
nand U10452 (N_10452,N_10364,N_10232);
nor U10453 (N_10453,N_10287,N_10283);
xnor U10454 (N_10454,N_10328,N_10221);
or U10455 (N_10455,N_10205,N_10296);
or U10456 (N_10456,N_10335,N_10278);
or U10457 (N_10457,N_10299,N_10302);
and U10458 (N_10458,N_10217,N_10281);
xnor U10459 (N_10459,N_10337,N_10382);
and U10460 (N_10460,N_10308,N_10224);
xor U10461 (N_10461,N_10234,N_10394);
and U10462 (N_10462,N_10303,N_10288);
nor U10463 (N_10463,N_10225,N_10266);
nand U10464 (N_10464,N_10336,N_10241);
nor U10465 (N_10465,N_10393,N_10248);
and U10466 (N_10466,N_10208,N_10275);
xnor U10467 (N_10467,N_10304,N_10361);
or U10468 (N_10468,N_10247,N_10203);
nor U10469 (N_10469,N_10329,N_10352);
or U10470 (N_10470,N_10334,N_10387);
or U10471 (N_10471,N_10359,N_10354);
xnor U10472 (N_10472,N_10253,N_10244);
xor U10473 (N_10473,N_10261,N_10355);
xor U10474 (N_10474,N_10300,N_10390);
xor U10475 (N_10475,N_10366,N_10320);
xnor U10476 (N_10476,N_10246,N_10272);
xnor U10477 (N_10477,N_10228,N_10397);
nand U10478 (N_10478,N_10262,N_10341);
and U10479 (N_10479,N_10218,N_10289);
and U10480 (N_10480,N_10279,N_10381);
nand U10481 (N_10481,N_10258,N_10293);
nand U10482 (N_10482,N_10282,N_10331);
nand U10483 (N_10483,N_10216,N_10316);
or U10484 (N_10484,N_10298,N_10265);
or U10485 (N_10485,N_10309,N_10347);
and U10486 (N_10486,N_10305,N_10277);
and U10487 (N_10487,N_10315,N_10353);
xnor U10488 (N_10488,N_10274,N_10373);
or U10489 (N_10489,N_10219,N_10239);
xnor U10490 (N_10490,N_10212,N_10229);
and U10491 (N_10491,N_10367,N_10251);
and U10492 (N_10492,N_10330,N_10344);
and U10493 (N_10493,N_10271,N_10204);
xor U10494 (N_10494,N_10256,N_10371);
nor U10495 (N_10495,N_10317,N_10200);
and U10496 (N_10496,N_10252,N_10377);
nand U10497 (N_10497,N_10368,N_10240);
nor U10498 (N_10498,N_10370,N_10310);
and U10499 (N_10499,N_10263,N_10362);
or U10500 (N_10500,N_10370,N_10281);
nand U10501 (N_10501,N_10217,N_10380);
and U10502 (N_10502,N_10307,N_10260);
nor U10503 (N_10503,N_10217,N_10366);
nand U10504 (N_10504,N_10277,N_10244);
xor U10505 (N_10505,N_10305,N_10243);
or U10506 (N_10506,N_10331,N_10361);
nor U10507 (N_10507,N_10260,N_10239);
xor U10508 (N_10508,N_10217,N_10382);
and U10509 (N_10509,N_10386,N_10374);
nor U10510 (N_10510,N_10292,N_10220);
and U10511 (N_10511,N_10352,N_10297);
nand U10512 (N_10512,N_10311,N_10365);
nor U10513 (N_10513,N_10200,N_10391);
or U10514 (N_10514,N_10284,N_10314);
xor U10515 (N_10515,N_10313,N_10253);
xor U10516 (N_10516,N_10315,N_10239);
xnor U10517 (N_10517,N_10323,N_10262);
or U10518 (N_10518,N_10307,N_10348);
nand U10519 (N_10519,N_10264,N_10309);
nor U10520 (N_10520,N_10338,N_10224);
xnor U10521 (N_10521,N_10366,N_10390);
xor U10522 (N_10522,N_10262,N_10360);
nor U10523 (N_10523,N_10246,N_10260);
and U10524 (N_10524,N_10313,N_10352);
nor U10525 (N_10525,N_10293,N_10339);
or U10526 (N_10526,N_10224,N_10334);
xor U10527 (N_10527,N_10246,N_10380);
nand U10528 (N_10528,N_10317,N_10275);
nor U10529 (N_10529,N_10335,N_10315);
xor U10530 (N_10530,N_10376,N_10207);
and U10531 (N_10531,N_10332,N_10334);
nand U10532 (N_10532,N_10375,N_10341);
xor U10533 (N_10533,N_10229,N_10256);
xor U10534 (N_10534,N_10265,N_10390);
or U10535 (N_10535,N_10351,N_10201);
and U10536 (N_10536,N_10374,N_10370);
nor U10537 (N_10537,N_10284,N_10312);
nor U10538 (N_10538,N_10311,N_10334);
nor U10539 (N_10539,N_10309,N_10222);
xnor U10540 (N_10540,N_10294,N_10304);
xor U10541 (N_10541,N_10339,N_10370);
and U10542 (N_10542,N_10292,N_10231);
xnor U10543 (N_10543,N_10338,N_10205);
xnor U10544 (N_10544,N_10255,N_10284);
or U10545 (N_10545,N_10398,N_10307);
or U10546 (N_10546,N_10298,N_10375);
nor U10547 (N_10547,N_10239,N_10313);
nand U10548 (N_10548,N_10213,N_10214);
and U10549 (N_10549,N_10390,N_10374);
xor U10550 (N_10550,N_10347,N_10396);
and U10551 (N_10551,N_10269,N_10313);
nand U10552 (N_10552,N_10253,N_10262);
nand U10553 (N_10553,N_10309,N_10228);
nor U10554 (N_10554,N_10247,N_10311);
and U10555 (N_10555,N_10391,N_10233);
nor U10556 (N_10556,N_10271,N_10303);
and U10557 (N_10557,N_10264,N_10260);
xor U10558 (N_10558,N_10375,N_10243);
and U10559 (N_10559,N_10200,N_10263);
and U10560 (N_10560,N_10330,N_10205);
and U10561 (N_10561,N_10291,N_10299);
xnor U10562 (N_10562,N_10327,N_10303);
nor U10563 (N_10563,N_10267,N_10346);
nor U10564 (N_10564,N_10291,N_10363);
nor U10565 (N_10565,N_10303,N_10227);
nor U10566 (N_10566,N_10331,N_10294);
nand U10567 (N_10567,N_10297,N_10307);
nor U10568 (N_10568,N_10258,N_10327);
nand U10569 (N_10569,N_10351,N_10294);
and U10570 (N_10570,N_10388,N_10228);
and U10571 (N_10571,N_10389,N_10247);
and U10572 (N_10572,N_10287,N_10205);
nor U10573 (N_10573,N_10269,N_10302);
and U10574 (N_10574,N_10311,N_10236);
xor U10575 (N_10575,N_10354,N_10292);
nor U10576 (N_10576,N_10310,N_10340);
or U10577 (N_10577,N_10384,N_10303);
or U10578 (N_10578,N_10277,N_10202);
or U10579 (N_10579,N_10393,N_10223);
nand U10580 (N_10580,N_10292,N_10311);
xnor U10581 (N_10581,N_10303,N_10245);
nor U10582 (N_10582,N_10338,N_10228);
nor U10583 (N_10583,N_10387,N_10304);
nor U10584 (N_10584,N_10302,N_10348);
xor U10585 (N_10585,N_10231,N_10232);
and U10586 (N_10586,N_10361,N_10287);
xor U10587 (N_10587,N_10288,N_10347);
or U10588 (N_10588,N_10308,N_10309);
xnor U10589 (N_10589,N_10375,N_10229);
or U10590 (N_10590,N_10253,N_10226);
and U10591 (N_10591,N_10311,N_10280);
nand U10592 (N_10592,N_10333,N_10324);
nand U10593 (N_10593,N_10226,N_10243);
nand U10594 (N_10594,N_10397,N_10209);
or U10595 (N_10595,N_10302,N_10314);
and U10596 (N_10596,N_10228,N_10273);
nand U10597 (N_10597,N_10273,N_10264);
or U10598 (N_10598,N_10247,N_10321);
and U10599 (N_10599,N_10327,N_10299);
nor U10600 (N_10600,N_10588,N_10505);
xor U10601 (N_10601,N_10557,N_10409);
and U10602 (N_10602,N_10489,N_10440);
and U10603 (N_10603,N_10425,N_10568);
nand U10604 (N_10604,N_10551,N_10576);
and U10605 (N_10605,N_10584,N_10547);
xnor U10606 (N_10606,N_10437,N_10495);
nand U10607 (N_10607,N_10436,N_10535);
nor U10608 (N_10608,N_10561,N_10564);
or U10609 (N_10609,N_10514,N_10593);
xor U10610 (N_10610,N_10468,N_10527);
nand U10611 (N_10611,N_10504,N_10571);
xnor U10612 (N_10612,N_10497,N_10528);
nand U10613 (N_10613,N_10506,N_10507);
xnor U10614 (N_10614,N_10502,N_10487);
or U10615 (N_10615,N_10525,N_10471);
nor U10616 (N_10616,N_10493,N_10444);
and U10617 (N_10617,N_10476,N_10474);
nand U10618 (N_10618,N_10524,N_10598);
nor U10619 (N_10619,N_10582,N_10407);
nand U10620 (N_10620,N_10591,N_10509);
or U10621 (N_10621,N_10555,N_10431);
nor U10622 (N_10622,N_10473,N_10516);
nor U10623 (N_10623,N_10549,N_10542);
and U10624 (N_10624,N_10475,N_10481);
nor U10625 (N_10625,N_10567,N_10586);
xnor U10626 (N_10626,N_10494,N_10556);
xor U10627 (N_10627,N_10403,N_10408);
nor U10628 (N_10628,N_10450,N_10522);
nor U10629 (N_10629,N_10491,N_10523);
xor U10630 (N_10630,N_10424,N_10415);
or U10631 (N_10631,N_10590,N_10530);
and U10632 (N_10632,N_10455,N_10460);
nor U10633 (N_10633,N_10581,N_10447);
and U10634 (N_10634,N_10410,N_10483);
and U10635 (N_10635,N_10463,N_10526);
nand U10636 (N_10636,N_10537,N_10445);
nand U10637 (N_10637,N_10416,N_10470);
xnor U10638 (N_10638,N_10429,N_10559);
and U10639 (N_10639,N_10540,N_10421);
nand U10640 (N_10640,N_10400,N_10417);
xor U10641 (N_10641,N_10404,N_10480);
or U10642 (N_10642,N_10521,N_10578);
or U10643 (N_10643,N_10513,N_10402);
nor U10644 (N_10644,N_10461,N_10466);
nor U10645 (N_10645,N_10577,N_10550);
nand U10646 (N_10646,N_10519,N_10496);
xor U10647 (N_10647,N_10478,N_10454);
and U10648 (N_10648,N_10511,N_10512);
and U10649 (N_10649,N_10401,N_10405);
xnor U10650 (N_10650,N_10548,N_10456);
xnor U10651 (N_10651,N_10482,N_10569);
and U10652 (N_10652,N_10565,N_10414);
nand U10653 (N_10653,N_10465,N_10413);
nor U10654 (N_10654,N_10448,N_10587);
nand U10655 (N_10655,N_10510,N_10443);
nor U10656 (N_10656,N_10426,N_10420);
nand U10657 (N_10657,N_10543,N_10490);
xor U10658 (N_10658,N_10427,N_10477);
nor U10659 (N_10659,N_10566,N_10563);
and U10660 (N_10660,N_10438,N_10595);
xnor U10661 (N_10661,N_10518,N_10486);
nand U10662 (N_10662,N_10508,N_10498);
nand U10663 (N_10663,N_10422,N_10579);
or U10664 (N_10664,N_10501,N_10594);
xnor U10665 (N_10665,N_10467,N_10485);
xnor U10666 (N_10666,N_10589,N_10599);
or U10667 (N_10667,N_10580,N_10458);
nor U10668 (N_10668,N_10552,N_10517);
nor U10669 (N_10669,N_10531,N_10453);
nand U10670 (N_10670,N_10435,N_10544);
nand U10671 (N_10671,N_10529,N_10558);
xor U10672 (N_10672,N_10539,N_10575);
nand U10673 (N_10673,N_10574,N_10464);
xor U10674 (N_10674,N_10553,N_10449);
xnor U10675 (N_10675,N_10541,N_10441);
nand U10676 (N_10676,N_10446,N_10585);
and U10677 (N_10677,N_10534,N_10442);
or U10678 (N_10678,N_10423,N_10492);
nor U10679 (N_10679,N_10452,N_10419);
nor U10680 (N_10680,N_10462,N_10432);
nor U10681 (N_10681,N_10545,N_10538);
xor U10682 (N_10682,N_10592,N_10433);
xnor U10683 (N_10683,N_10488,N_10451);
xnor U10684 (N_10684,N_10570,N_10546);
or U10685 (N_10685,N_10434,N_10469);
nand U10686 (N_10686,N_10520,N_10532);
nor U10687 (N_10687,N_10573,N_10560);
xor U10688 (N_10688,N_10484,N_10515);
and U10689 (N_10689,N_10406,N_10499);
nor U10690 (N_10690,N_10536,N_10596);
nor U10691 (N_10691,N_10503,N_10411);
or U10692 (N_10692,N_10597,N_10418);
xnor U10693 (N_10693,N_10533,N_10459);
nand U10694 (N_10694,N_10572,N_10583);
and U10695 (N_10695,N_10472,N_10430);
and U10696 (N_10696,N_10412,N_10562);
xnor U10697 (N_10697,N_10428,N_10457);
or U10698 (N_10698,N_10479,N_10500);
nor U10699 (N_10699,N_10439,N_10554);
or U10700 (N_10700,N_10528,N_10492);
or U10701 (N_10701,N_10454,N_10577);
xor U10702 (N_10702,N_10448,N_10481);
nand U10703 (N_10703,N_10412,N_10576);
xor U10704 (N_10704,N_10531,N_10471);
nand U10705 (N_10705,N_10595,N_10507);
nor U10706 (N_10706,N_10583,N_10511);
xor U10707 (N_10707,N_10592,N_10557);
nand U10708 (N_10708,N_10504,N_10503);
nor U10709 (N_10709,N_10542,N_10595);
nor U10710 (N_10710,N_10542,N_10474);
nor U10711 (N_10711,N_10447,N_10443);
xnor U10712 (N_10712,N_10543,N_10415);
xnor U10713 (N_10713,N_10573,N_10534);
nor U10714 (N_10714,N_10516,N_10580);
or U10715 (N_10715,N_10457,N_10484);
or U10716 (N_10716,N_10562,N_10451);
or U10717 (N_10717,N_10454,N_10422);
xnor U10718 (N_10718,N_10483,N_10501);
nor U10719 (N_10719,N_10427,N_10532);
or U10720 (N_10720,N_10492,N_10580);
nor U10721 (N_10721,N_10416,N_10404);
xor U10722 (N_10722,N_10430,N_10480);
and U10723 (N_10723,N_10428,N_10591);
or U10724 (N_10724,N_10406,N_10566);
xor U10725 (N_10725,N_10580,N_10594);
nor U10726 (N_10726,N_10437,N_10527);
or U10727 (N_10727,N_10584,N_10444);
and U10728 (N_10728,N_10479,N_10427);
nand U10729 (N_10729,N_10565,N_10448);
xor U10730 (N_10730,N_10548,N_10539);
and U10731 (N_10731,N_10480,N_10524);
xnor U10732 (N_10732,N_10584,N_10494);
and U10733 (N_10733,N_10458,N_10438);
or U10734 (N_10734,N_10556,N_10453);
nor U10735 (N_10735,N_10574,N_10555);
and U10736 (N_10736,N_10445,N_10441);
and U10737 (N_10737,N_10418,N_10529);
nand U10738 (N_10738,N_10578,N_10463);
nand U10739 (N_10739,N_10595,N_10445);
xnor U10740 (N_10740,N_10598,N_10571);
nand U10741 (N_10741,N_10519,N_10444);
nor U10742 (N_10742,N_10576,N_10436);
nor U10743 (N_10743,N_10414,N_10436);
nand U10744 (N_10744,N_10560,N_10400);
or U10745 (N_10745,N_10422,N_10472);
nor U10746 (N_10746,N_10407,N_10464);
nor U10747 (N_10747,N_10566,N_10428);
or U10748 (N_10748,N_10501,N_10543);
nor U10749 (N_10749,N_10526,N_10499);
xnor U10750 (N_10750,N_10483,N_10551);
and U10751 (N_10751,N_10496,N_10521);
and U10752 (N_10752,N_10420,N_10467);
or U10753 (N_10753,N_10427,N_10562);
and U10754 (N_10754,N_10405,N_10488);
xnor U10755 (N_10755,N_10409,N_10472);
xor U10756 (N_10756,N_10465,N_10475);
and U10757 (N_10757,N_10568,N_10583);
or U10758 (N_10758,N_10490,N_10536);
nand U10759 (N_10759,N_10579,N_10509);
nor U10760 (N_10760,N_10564,N_10421);
nand U10761 (N_10761,N_10492,N_10502);
nand U10762 (N_10762,N_10518,N_10536);
or U10763 (N_10763,N_10590,N_10416);
xor U10764 (N_10764,N_10451,N_10596);
nand U10765 (N_10765,N_10552,N_10448);
and U10766 (N_10766,N_10534,N_10465);
nand U10767 (N_10767,N_10496,N_10464);
or U10768 (N_10768,N_10507,N_10592);
and U10769 (N_10769,N_10545,N_10502);
or U10770 (N_10770,N_10500,N_10448);
xor U10771 (N_10771,N_10445,N_10418);
xnor U10772 (N_10772,N_10440,N_10476);
xor U10773 (N_10773,N_10508,N_10533);
nand U10774 (N_10774,N_10502,N_10427);
nor U10775 (N_10775,N_10528,N_10549);
nand U10776 (N_10776,N_10427,N_10528);
nand U10777 (N_10777,N_10468,N_10426);
nor U10778 (N_10778,N_10556,N_10504);
nand U10779 (N_10779,N_10574,N_10479);
nor U10780 (N_10780,N_10522,N_10565);
xnor U10781 (N_10781,N_10512,N_10569);
xor U10782 (N_10782,N_10500,N_10474);
xnor U10783 (N_10783,N_10560,N_10516);
nor U10784 (N_10784,N_10469,N_10574);
or U10785 (N_10785,N_10528,N_10593);
and U10786 (N_10786,N_10524,N_10587);
nor U10787 (N_10787,N_10449,N_10459);
and U10788 (N_10788,N_10553,N_10534);
nor U10789 (N_10789,N_10561,N_10518);
nand U10790 (N_10790,N_10467,N_10547);
nand U10791 (N_10791,N_10535,N_10454);
xor U10792 (N_10792,N_10424,N_10410);
nand U10793 (N_10793,N_10486,N_10580);
xor U10794 (N_10794,N_10412,N_10487);
and U10795 (N_10795,N_10439,N_10526);
or U10796 (N_10796,N_10449,N_10559);
or U10797 (N_10797,N_10555,N_10416);
and U10798 (N_10798,N_10489,N_10431);
xnor U10799 (N_10799,N_10410,N_10429);
or U10800 (N_10800,N_10667,N_10688);
xor U10801 (N_10801,N_10659,N_10745);
xnor U10802 (N_10802,N_10689,N_10655);
nor U10803 (N_10803,N_10680,N_10799);
nand U10804 (N_10804,N_10768,N_10629);
xor U10805 (N_10805,N_10706,N_10735);
or U10806 (N_10806,N_10737,N_10767);
nand U10807 (N_10807,N_10726,N_10711);
and U10808 (N_10808,N_10698,N_10707);
xnor U10809 (N_10809,N_10662,N_10666);
xor U10810 (N_10810,N_10676,N_10686);
nor U10811 (N_10811,N_10732,N_10777);
xor U10812 (N_10812,N_10741,N_10634);
xor U10813 (N_10813,N_10715,N_10644);
nand U10814 (N_10814,N_10759,N_10675);
xor U10815 (N_10815,N_10791,N_10635);
nand U10816 (N_10816,N_10673,N_10646);
xnor U10817 (N_10817,N_10754,N_10758);
xor U10818 (N_10818,N_10690,N_10625);
or U10819 (N_10819,N_10751,N_10624);
and U10820 (N_10820,N_10749,N_10782);
or U10821 (N_10821,N_10660,N_10691);
or U10822 (N_10822,N_10653,N_10752);
nor U10823 (N_10823,N_10795,N_10720);
nor U10824 (N_10824,N_10613,N_10772);
nor U10825 (N_10825,N_10658,N_10652);
and U10826 (N_10826,N_10731,N_10786);
nand U10827 (N_10827,N_10610,N_10612);
and U10828 (N_10828,N_10779,N_10748);
nor U10829 (N_10829,N_10616,N_10778);
and U10830 (N_10830,N_10702,N_10746);
nand U10831 (N_10831,N_10723,N_10770);
nand U10832 (N_10832,N_10716,N_10774);
or U10833 (N_10833,N_10750,N_10605);
and U10834 (N_10834,N_10794,N_10760);
nor U10835 (N_10835,N_10651,N_10722);
and U10836 (N_10836,N_10641,N_10609);
or U10837 (N_10837,N_10661,N_10600);
or U10838 (N_10838,N_10684,N_10733);
xnor U10839 (N_10839,N_10717,N_10674);
nor U10840 (N_10840,N_10643,N_10788);
nor U10841 (N_10841,N_10704,N_10623);
nand U10842 (N_10842,N_10650,N_10769);
or U10843 (N_10843,N_10739,N_10725);
and U10844 (N_10844,N_10695,N_10763);
xor U10845 (N_10845,N_10789,N_10796);
or U10846 (N_10846,N_10626,N_10649);
nor U10847 (N_10847,N_10742,N_10632);
nor U10848 (N_10848,N_10756,N_10678);
nor U10849 (N_10849,N_10679,N_10743);
nor U10850 (N_10850,N_10633,N_10614);
xnor U10851 (N_10851,N_10622,N_10645);
xor U10852 (N_10852,N_10700,N_10697);
or U10853 (N_10853,N_10773,N_10714);
nor U10854 (N_10854,N_10738,N_10683);
xnor U10855 (N_10855,N_10656,N_10757);
and U10856 (N_10856,N_10775,N_10640);
and U10857 (N_10857,N_10618,N_10730);
nor U10858 (N_10858,N_10708,N_10607);
and U10859 (N_10859,N_10712,N_10761);
and U10860 (N_10860,N_10669,N_10630);
xnor U10861 (N_10861,N_10639,N_10718);
and U10862 (N_10862,N_10764,N_10628);
nor U10863 (N_10863,N_10664,N_10766);
nor U10864 (N_10864,N_10699,N_10710);
and U10865 (N_10865,N_10703,N_10780);
xor U10866 (N_10866,N_10642,N_10719);
nor U10867 (N_10867,N_10696,N_10736);
and U10868 (N_10868,N_10665,N_10681);
nand U10869 (N_10869,N_10747,N_10621);
nand U10870 (N_10870,N_10762,N_10734);
nand U10871 (N_10871,N_10617,N_10755);
nand U10872 (N_10872,N_10663,N_10627);
or U10873 (N_10873,N_10787,N_10728);
nor U10874 (N_10874,N_10685,N_10672);
and U10875 (N_10875,N_10729,N_10765);
and U10876 (N_10876,N_10631,N_10771);
nor U10877 (N_10877,N_10784,N_10647);
xnor U10878 (N_10878,N_10790,N_10694);
nor U10879 (N_10879,N_10636,N_10753);
nor U10880 (N_10880,N_10783,N_10606);
xor U10881 (N_10881,N_10693,N_10608);
and U10882 (N_10882,N_10602,N_10721);
nor U10883 (N_10883,N_10744,N_10619);
nor U10884 (N_10884,N_10677,N_10668);
nand U10885 (N_10885,N_10713,N_10781);
nand U10886 (N_10886,N_10657,N_10740);
nor U10887 (N_10887,N_10670,N_10638);
and U10888 (N_10888,N_10615,N_10682);
nand U10889 (N_10889,N_10724,N_10620);
nor U10890 (N_10890,N_10687,N_10604);
nor U10891 (N_10891,N_10792,N_10798);
nor U10892 (N_10892,N_10603,N_10727);
xor U10893 (N_10893,N_10705,N_10601);
xor U10894 (N_10894,N_10648,N_10654);
and U10895 (N_10895,N_10793,N_10637);
nor U10896 (N_10896,N_10611,N_10701);
and U10897 (N_10897,N_10709,N_10692);
nand U10898 (N_10898,N_10776,N_10797);
nand U10899 (N_10899,N_10785,N_10671);
nor U10900 (N_10900,N_10714,N_10625);
and U10901 (N_10901,N_10621,N_10675);
nand U10902 (N_10902,N_10617,N_10754);
and U10903 (N_10903,N_10695,N_10751);
nor U10904 (N_10904,N_10779,N_10642);
or U10905 (N_10905,N_10620,N_10711);
or U10906 (N_10906,N_10715,N_10766);
or U10907 (N_10907,N_10766,N_10637);
or U10908 (N_10908,N_10622,N_10737);
and U10909 (N_10909,N_10727,N_10763);
nand U10910 (N_10910,N_10663,N_10664);
and U10911 (N_10911,N_10727,N_10674);
xor U10912 (N_10912,N_10710,N_10642);
nand U10913 (N_10913,N_10703,N_10736);
nor U10914 (N_10914,N_10631,N_10675);
nor U10915 (N_10915,N_10738,N_10785);
xor U10916 (N_10916,N_10743,N_10660);
or U10917 (N_10917,N_10764,N_10776);
and U10918 (N_10918,N_10657,N_10721);
nand U10919 (N_10919,N_10709,N_10635);
nand U10920 (N_10920,N_10726,N_10776);
nor U10921 (N_10921,N_10744,N_10643);
nand U10922 (N_10922,N_10615,N_10632);
nand U10923 (N_10923,N_10684,N_10601);
or U10924 (N_10924,N_10693,N_10768);
nor U10925 (N_10925,N_10609,N_10618);
or U10926 (N_10926,N_10653,N_10741);
xor U10927 (N_10927,N_10719,N_10733);
or U10928 (N_10928,N_10654,N_10705);
xnor U10929 (N_10929,N_10740,N_10769);
and U10930 (N_10930,N_10777,N_10796);
or U10931 (N_10931,N_10654,N_10730);
and U10932 (N_10932,N_10732,N_10627);
xnor U10933 (N_10933,N_10774,N_10648);
and U10934 (N_10934,N_10713,N_10732);
nand U10935 (N_10935,N_10693,N_10783);
nor U10936 (N_10936,N_10701,N_10707);
or U10937 (N_10937,N_10736,N_10632);
nor U10938 (N_10938,N_10601,N_10741);
xnor U10939 (N_10939,N_10749,N_10623);
xor U10940 (N_10940,N_10786,N_10665);
nand U10941 (N_10941,N_10606,N_10734);
or U10942 (N_10942,N_10776,N_10791);
nand U10943 (N_10943,N_10685,N_10727);
and U10944 (N_10944,N_10688,N_10650);
nand U10945 (N_10945,N_10695,N_10653);
or U10946 (N_10946,N_10715,N_10710);
or U10947 (N_10947,N_10731,N_10601);
and U10948 (N_10948,N_10620,N_10758);
and U10949 (N_10949,N_10664,N_10666);
xnor U10950 (N_10950,N_10660,N_10622);
xnor U10951 (N_10951,N_10778,N_10794);
xnor U10952 (N_10952,N_10745,N_10618);
nor U10953 (N_10953,N_10748,N_10790);
nand U10954 (N_10954,N_10679,N_10655);
xnor U10955 (N_10955,N_10781,N_10679);
nor U10956 (N_10956,N_10738,N_10719);
nor U10957 (N_10957,N_10656,N_10781);
nand U10958 (N_10958,N_10716,N_10618);
nor U10959 (N_10959,N_10663,N_10687);
or U10960 (N_10960,N_10620,N_10785);
nor U10961 (N_10961,N_10616,N_10625);
and U10962 (N_10962,N_10658,N_10649);
and U10963 (N_10963,N_10657,N_10746);
nand U10964 (N_10964,N_10770,N_10630);
xnor U10965 (N_10965,N_10694,N_10754);
nand U10966 (N_10966,N_10717,N_10737);
or U10967 (N_10967,N_10683,N_10761);
xor U10968 (N_10968,N_10726,N_10768);
xnor U10969 (N_10969,N_10715,N_10773);
and U10970 (N_10970,N_10742,N_10757);
nand U10971 (N_10971,N_10760,N_10676);
or U10972 (N_10972,N_10609,N_10633);
nor U10973 (N_10973,N_10611,N_10636);
nand U10974 (N_10974,N_10675,N_10763);
nand U10975 (N_10975,N_10794,N_10691);
xnor U10976 (N_10976,N_10786,N_10677);
or U10977 (N_10977,N_10677,N_10757);
or U10978 (N_10978,N_10681,N_10776);
and U10979 (N_10979,N_10680,N_10780);
xor U10980 (N_10980,N_10613,N_10697);
nor U10981 (N_10981,N_10701,N_10711);
or U10982 (N_10982,N_10705,N_10630);
nand U10983 (N_10983,N_10604,N_10693);
nand U10984 (N_10984,N_10732,N_10776);
xor U10985 (N_10985,N_10658,N_10702);
nand U10986 (N_10986,N_10659,N_10703);
nor U10987 (N_10987,N_10647,N_10765);
nand U10988 (N_10988,N_10680,N_10703);
or U10989 (N_10989,N_10669,N_10614);
xnor U10990 (N_10990,N_10700,N_10656);
and U10991 (N_10991,N_10723,N_10708);
and U10992 (N_10992,N_10730,N_10653);
or U10993 (N_10993,N_10630,N_10721);
xnor U10994 (N_10994,N_10629,N_10733);
or U10995 (N_10995,N_10730,N_10792);
and U10996 (N_10996,N_10697,N_10635);
or U10997 (N_10997,N_10617,N_10631);
nor U10998 (N_10998,N_10714,N_10686);
nand U10999 (N_10999,N_10699,N_10641);
or U11000 (N_11000,N_10877,N_10909);
xnor U11001 (N_11001,N_10945,N_10912);
nor U11002 (N_11002,N_10808,N_10905);
or U11003 (N_11003,N_10911,N_10817);
or U11004 (N_11004,N_10851,N_10848);
nor U11005 (N_11005,N_10875,N_10862);
xor U11006 (N_11006,N_10828,N_10842);
xnor U11007 (N_11007,N_10918,N_10929);
or U11008 (N_11008,N_10984,N_10972);
and U11009 (N_11009,N_10947,N_10873);
xor U11010 (N_11010,N_10809,N_10993);
or U11011 (N_11011,N_10802,N_10902);
nand U11012 (N_11012,N_10950,N_10879);
or U11013 (N_11013,N_10805,N_10895);
and U11014 (N_11014,N_10932,N_10910);
xnor U11015 (N_11015,N_10846,N_10840);
xor U11016 (N_11016,N_10983,N_10874);
or U11017 (N_11017,N_10847,N_10922);
xnor U11018 (N_11018,N_10974,N_10948);
and U11019 (N_11019,N_10927,N_10944);
or U11020 (N_11020,N_10959,N_10903);
nor U11021 (N_11021,N_10941,N_10928);
and U11022 (N_11022,N_10931,N_10892);
nand U11023 (N_11023,N_10855,N_10819);
xor U11024 (N_11024,N_10966,N_10853);
or U11025 (N_11025,N_10878,N_10955);
or U11026 (N_11026,N_10890,N_10998);
nand U11027 (N_11027,N_10858,N_10963);
or U11028 (N_11028,N_10867,N_10889);
nor U11029 (N_11029,N_10881,N_10872);
or U11030 (N_11030,N_10813,N_10990);
nor U11031 (N_11031,N_10982,N_10801);
nor U11032 (N_11032,N_10830,N_10876);
nand U11033 (N_11033,N_10859,N_10991);
nand U11034 (N_11034,N_10917,N_10899);
nor U11035 (N_11035,N_10898,N_10829);
and U11036 (N_11036,N_10852,N_10882);
and U11037 (N_11037,N_10836,N_10961);
or U11038 (N_11038,N_10850,N_10967);
xor U11039 (N_11039,N_10865,N_10854);
xnor U11040 (N_11040,N_10832,N_10958);
xor U11041 (N_11041,N_10915,N_10921);
and U11042 (N_11042,N_10887,N_10893);
or U11043 (N_11043,N_10996,N_10936);
and U11044 (N_11044,N_10841,N_10886);
or U11045 (N_11045,N_10926,N_10952);
nand U11046 (N_11046,N_10992,N_10821);
nand U11047 (N_11047,N_10839,N_10976);
nand U11048 (N_11048,N_10834,N_10951);
or U11049 (N_11049,N_10980,N_10897);
and U11050 (N_11050,N_10816,N_10975);
nand U11051 (N_11051,N_10815,N_10934);
nor U11052 (N_11052,N_10940,N_10857);
xnor U11053 (N_11053,N_10985,N_10870);
and U11054 (N_11054,N_10826,N_10986);
nor U11055 (N_11055,N_10949,N_10837);
nand U11056 (N_11056,N_10919,N_10856);
nand U11057 (N_11057,N_10885,N_10920);
xor U11058 (N_11058,N_10962,N_10994);
xor U11059 (N_11059,N_10888,N_10861);
or U11060 (N_11060,N_10880,N_10868);
or U11061 (N_11061,N_10891,N_10849);
nor U11062 (N_11062,N_10954,N_10900);
xnor U11063 (N_11063,N_10864,N_10823);
xnor U11064 (N_11064,N_10894,N_10866);
xor U11065 (N_11065,N_10973,N_10933);
nand U11066 (N_11066,N_10968,N_10981);
nor U11067 (N_11067,N_10906,N_10925);
or U11068 (N_11068,N_10814,N_10969);
or U11069 (N_11069,N_10844,N_10939);
or U11070 (N_11070,N_10824,N_10970);
or U11071 (N_11071,N_10971,N_10937);
and U11072 (N_11072,N_10822,N_10965);
and U11073 (N_11073,N_10884,N_10913);
nand U11074 (N_11074,N_10883,N_10953);
xor U11075 (N_11075,N_10978,N_10979);
and U11076 (N_11076,N_10935,N_10871);
nand U11077 (N_11077,N_10827,N_10916);
or U11078 (N_11078,N_10803,N_10838);
or U11079 (N_11079,N_10820,N_10989);
xor U11080 (N_11080,N_10818,N_10831);
xor U11081 (N_11081,N_10812,N_10908);
nor U11082 (N_11082,N_10942,N_10901);
and U11083 (N_11083,N_10964,N_10863);
xor U11084 (N_11084,N_10999,N_10930);
or U11085 (N_11085,N_10988,N_10811);
or U11086 (N_11086,N_10806,N_10807);
and U11087 (N_11087,N_10977,N_10896);
xor U11088 (N_11088,N_10987,N_10907);
nor U11089 (N_11089,N_10860,N_10938);
and U11090 (N_11090,N_10943,N_10946);
or U11091 (N_11091,N_10914,N_10997);
xor U11092 (N_11092,N_10869,N_10800);
nor U11093 (N_11093,N_10960,N_10810);
nor U11094 (N_11094,N_10804,N_10923);
nor U11095 (N_11095,N_10835,N_10845);
or U11096 (N_11096,N_10957,N_10833);
and U11097 (N_11097,N_10904,N_10956);
nor U11098 (N_11098,N_10995,N_10843);
xor U11099 (N_11099,N_10825,N_10924);
and U11100 (N_11100,N_10810,N_10813);
nand U11101 (N_11101,N_10985,N_10842);
nor U11102 (N_11102,N_10824,N_10943);
or U11103 (N_11103,N_10892,N_10854);
or U11104 (N_11104,N_10802,N_10965);
nor U11105 (N_11105,N_10951,N_10803);
nand U11106 (N_11106,N_10856,N_10983);
and U11107 (N_11107,N_10857,N_10963);
and U11108 (N_11108,N_10831,N_10980);
nand U11109 (N_11109,N_10983,N_10806);
or U11110 (N_11110,N_10873,N_10834);
xnor U11111 (N_11111,N_10951,N_10920);
and U11112 (N_11112,N_10816,N_10800);
xnor U11113 (N_11113,N_10979,N_10934);
xor U11114 (N_11114,N_10941,N_10855);
xor U11115 (N_11115,N_10986,N_10802);
xor U11116 (N_11116,N_10827,N_10947);
nand U11117 (N_11117,N_10982,N_10812);
and U11118 (N_11118,N_10815,N_10841);
xor U11119 (N_11119,N_10976,N_10994);
xnor U11120 (N_11120,N_10902,N_10874);
or U11121 (N_11121,N_10867,N_10921);
nor U11122 (N_11122,N_10910,N_10835);
xnor U11123 (N_11123,N_10891,N_10967);
and U11124 (N_11124,N_10937,N_10868);
or U11125 (N_11125,N_10948,N_10850);
nand U11126 (N_11126,N_10820,N_10900);
nand U11127 (N_11127,N_10995,N_10893);
xnor U11128 (N_11128,N_10917,N_10903);
nor U11129 (N_11129,N_10968,N_10858);
and U11130 (N_11130,N_10814,N_10919);
or U11131 (N_11131,N_10994,N_10970);
nor U11132 (N_11132,N_10937,N_10805);
and U11133 (N_11133,N_10874,N_10885);
nand U11134 (N_11134,N_10850,N_10913);
and U11135 (N_11135,N_10860,N_10828);
nor U11136 (N_11136,N_10884,N_10927);
or U11137 (N_11137,N_10812,N_10814);
nand U11138 (N_11138,N_10835,N_10941);
nand U11139 (N_11139,N_10943,N_10922);
or U11140 (N_11140,N_10876,N_10918);
xor U11141 (N_11141,N_10996,N_10870);
xnor U11142 (N_11142,N_10837,N_10891);
or U11143 (N_11143,N_10894,N_10848);
or U11144 (N_11144,N_10982,N_10959);
nor U11145 (N_11145,N_10809,N_10969);
nor U11146 (N_11146,N_10828,N_10877);
nor U11147 (N_11147,N_10837,N_10964);
xor U11148 (N_11148,N_10854,N_10870);
nor U11149 (N_11149,N_10954,N_10878);
xnor U11150 (N_11150,N_10820,N_10828);
or U11151 (N_11151,N_10845,N_10890);
and U11152 (N_11152,N_10802,N_10858);
nand U11153 (N_11153,N_10804,N_10882);
nand U11154 (N_11154,N_10993,N_10882);
nor U11155 (N_11155,N_10878,N_10893);
and U11156 (N_11156,N_10803,N_10898);
nor U11157 (N_11157,N_10856,N_10980);
nand U11158 (N_11158,N_10816,N_10959);
or U11159 (N_11159,N_10917,N_10991);
or U11160 (N_11160,N_10971,N_10994);
nor U11161 (N_11161,N_10877,N_10891);
and U11162 (N_11162,N_10986,N_10901);
or U11163 (N_11163,N_10948,N_10817);
or U11164 (N_11164,N_10824,N_10964);
or U11165 (N_11165,N_10806,N_10955);
xor U11166 (N_11166,N_10923,N_10928);
and U11167 (N_11167,N_10928,N_10956);
xor U11168 (N_11168,N_10800,N_10849);
nand U11169 (N_11169,N_10975,N_10952);
and U11170 (N_11170,N_10959,N_10968);
or U11171 (N_11171,N_10953,N_10929);
and U11172 (N_11172,N_10808,N_10854);
or U11173 (N_11173,N_10819,N_10908);
nand U11174 (N_11174,N_10928,N_10998);
nor U11175 (N_11175,N_10938,N_10842);
and U11176 (N_11176,N_10937,N_10860);
nand U11177 (N_11177,N_10800,N_10858);
or U11178 (N_11178,N_10900,N_10927);
and U11179 (N_11179,N_10855,N_10800);
and U11180 (N_11180,N_10840,N_10949);
nand U11181 (N_11181,N_10898,N_10993);
nor U11182 (N_11182,N_10822,N_10840);
or U11183 (N_11183,N_10849,N_10890);
or U11184 (N_11184,N_10912,N_10871);
nand U11185 (N_11185,N_10978,N_10958);
nand U11186 (N_11186,N_10850,N_10978);
and U11187 (N_11187,N_10922,N_10814);
or U11188 (N_11188,N_10809,N_10951);
nor U11189 (N_11189,N_10938,N_10898);
nor U11190 (N_11190,N_10896,N_10804);
nand U11191 (N_11191,N_10842,N_10853);
nor U11192 (N_11192,N_10936,N_10914);
xnor U11193 (N_11193,N_10872,N_10900);
or U11194 (N_11194,N_10914,N_10896);
nor U11195 (N_11195,N_10907,N_10917);
nand U11196 (N_11196,N_10958,N_10922);
and U11197 (N_11197,N_10872,N_10991);
nor U11198 (N_11198,N_10919,N_10838);
or U11199 (N_11199,N_10857,N_10864);
nand U11200 (N_11200,N_11157,N_11098);
xor U11201 (N_11201,N_11173,N_11124);
or U11202 (N_11202,N_11144,N_11026);
nand U11203 (N_11203,N_11082,N_11051);
nor U11204 (N_11204,N_11185,N_11145);
or U11205 (N_11205,N_11078,N_11190);
xor U11206 (N_11206,N_11084,N_11132);
xor U11207 (N_11207,N_11116,N_11104);
nor U11208 (N_11208,N_11014,N_11161);
nand U11209 (N_11209,N_11058,N_11034);
nor U11210 (N_11210,N_11071,N_11008);
or U11211 (N_11211,N_11126,N_11075);
and U11212 (N_11212,N_11148,N_11167);
or U11213 (N_11213,N_11041,N_11138);
nand U11214 (N_11214,N_11088,N_11068);
or U11215 (N_11215,N_11069,N_11196);
nand U11216 (N_11216,N_11007,N_11150);
and U11217 (N_11217,N_11015,N_11044);
or U11218 (N_11218,N_11010,N_11127);
xnor U11219 (N_11219,N_11159,N_11181);
xnor U11220 (N_11220,N_11067,N_11012);
nand U11221 (N_11221,N_11095,N_11101);
xnor U11222 (N_11222,N_11178,N_11057);
xor U11223 (N_11223,N_11062,N_11146);
xor U11224 (N_11224,N_11176,N_11121);
or U11225 (N_11225,N_11093,N_11042);
or U11226 (N_11226,N_11056,N_11184);
xor U11227 (N_11227,N_11166,N_11091);
and U11228 (N_11228,N_11153,N_11179);
nand U11229 (N_11229,N_11103,N_11073);
and U11230 (N_11230,N_11003,N_11013);
nand U11231 (N_11231,N_11165,N_11152);
xnor U11232 (N_11232,N_11183,N_11081);
nand U11233 (N_11233,N_11032,N_11050);
nand U11234 (N_11234,N_11059,N_11024);
nand U11235 (N_11235,N_11100,N_11065);
or U11236 (N_11236,N_11049,N_11072);
and U11237 (N_11237,N_11137,N_11115);
or U11238 (N_11238,N_11187,N_11035);
nor U11239 (N_11239,N_11142,N_11037);
or U11240 (N_11240,N_11096,N_11197);
and U11241 (N_11241,N_11143,N_11054);
and U11242 (N_11242,N_11122,N_11195);
nor U11243 (N_11243,N_11106,N_11135);
nand U11244 (N_11244,N_11114,N_11099);
nor U11245 (N_11245,N_11079,N_11182);
nor U11246 (N_11246,N_11193,N_11011);
and U11247 (N_11247,N_11021,N_11188);
and U11248 (N_11248,N_11117,N_11005);
nor U11249 (N_11249,N_11000,N_11060);
and U11250 (N_11250,N_11023,N_11199);
or U11251 (N_11251,N_11118,N_11040);
nand U11252 (N_11252,N_11017,N_11194);
or U11253 (N_11253,N_11141,N_11052);
nand U11254 (N_11254,N_11149,N_11076);
or U11255 (N_11255,N_11047,N_11033);
or U11256 (N_11256,N_11027,N_11154);
nor U11257 (N_11257,N_11109,N_11186);
xor U11258 (N_11258,N_11112,N_11006);
or U11259 (N_11259,N_11070,N_11134);
nand U11260 (N_11260,N_11139,N_11043);
nand U11261 (N_11261,N_11198,N_11036);
nor U11262 (N_11262,N_11066,N_11077);
xor U11263 (N_11263,N_11048,N_11158);
nand U11264 (N_11264,N_11031,N_11022);
or U11265 (N_11265,N_11151,N_11002);
nor U11266 (N_11266,N_11192,N_11001);
or U11267 (N_11267,N_11140,N_11162);
or U11268 (N_11268,N_11180,N_11174);
and U11269 (N_11269,N_11063,N_11029);
nand U11270 (N_11270,N_11053,N_11092);
nor U11271 (N_11271,N_11085,N_11080);
xor U11272 (N_11272,N_11136,N_11163);
or U11273 (N_11273,N_11020,N_11130);
nor U11274 (N_11274,N_11061,N_11120);
nor U11275 (N_11275,N_11046,N_11083);
nor U11276 (N_11276,N_11171,N_11175);
xnor U11277 (N_11277,N_11133,N_11170);
and U11278 (N_11278,N_11131,N_11016);
nor U11279 (N_11279,N_11074,N_11156);
xor U11280 (N_11280,N_11105,N_11097);
or U11281 (N_11281,N_11160,N_11087);
and U11282 (N_11282,N_11125,N_11086);
xnor U11283 (N_11283,N_11164,N_11111);
nand U11284 (N_11284,N_11191,N_11168);
nor U11285 (N_11285,N_11107,N_11055);
nand U11286 (N_11286,N_11045,N_11064);
nor U11287 (N_11287,N_11018,N_11177);
xor U11288 (N_11288,N_11102,N_11089);
xnor U11289 (N_11289,N_11039,N_11113);
nor U11290 (N_11290,N_11169,N_11172);
xnor U11291 (N_11291,N_11025,N_11108);
and U11292 (N_11292,N_11009,N_11128);
nor U11293 (N_11293,N_11147,N_11155);
or U11294 (N_11294,N_11030,N_11129);
and U11295 (N_11295,N_11189,N_11038);
xor U11296 (N_11296,N_11110,N_11004);
nand U11297 (N_11297,N_11028,N_11123);
or U11298 (N_11298,N_11019,N_11094);
nand U11299 (N_11299,N_11090,N_11119);
or U11300 (N_11300,N_11022,N_11173);
and U11301 (N_11301,N_11145,N_11130);
and U11302 (N_11302,N_11046,N_11165);
nor U11303 (N_11303,N_11011,N_11120);
nand U11304 (N_11304,N_11074,N_11059);
nor U11305 (N_11305,N_11116,N_11111);
xor U11306 (N_11306,N_11082,N_11073);
and U11307 (N_11307,N_11049,N_11177);
nand U11308 (N_11308,N_11180,N_11133);
xor U11309 (N_11309,N_11109,N_11025);
xor U11310 (N_11310,N_11040,N_11094);
xor U11311 (N_11311,N_11127,N_11059);
xnor U11312 (N_11312,N_11121,N_11074);
xnor U11313 (N_11313,N_11061,N_11082);
and U11314 (N_11314,N_11089,N_11023);
and U11315 (N_11315,N_11065,N_11076);
or U11316 (N_11316,N_11004,N_11057);
or U11317 (N_11317,N_11085,N_11128);
nor U11318 (N_11318,N_11181,N_11149);
xor U11319 (N_11319,N_11051,N_11101);
xor U11320 (N_11320,N_11126,N_11124);
nor U11321 (N_11321,N_11047,N_11190);
and U11322 (N_11322,N_11127,N_11069);
nor U11323 (N_11323,N_11193,N_11161);
nand U11324 (N_11324,N_11167,N_11042);
or U11325 (N_11325,N_11130,N_11022);
nor U11326 (N_11326,N_11050,N_11109);
nor U11327 (N_11327,N_11067,N_11198);
or U11328 (N_11328,N_11151,N_11112);
nand U11329 (N_11329,N_11061,N_11068);
or U11330 (N_11330,N_11059,N_11071);
xnor U11331 (N_11331,N_11061,N_11180);
and U11332 (N_11332,N_11061,N_11168);
or U11333 (N_11333,N_11066,N_11028);
and U11334 (N_11334,N_11019,N_11043);
xnor U11335 (N_11335,N_11024,N_11156);
nand U11336 (N_11336,N_11078,N_11007);
and U11337 (N_11337,N_11119,N_11192);
xor U11338 (N_11338,N_11030,N_11070);
or U11339 (N_11339,N_11098,N_11075);
or U11340 (N_11340,N_11176,N_11009);
xnor U11341 (N_11341,N_11158,N_11020);
nand U11342 (N_11342,N_11098,N_11197);
or U11343 (N_11343,N_11065,N_11059);
nand U11344 (N_11344,N_11165,N_11029);
and U11345 (N_11345,N_11185,N_11174);
or U11346 (N_11346,N_11032,N_11097);
nor U11347 (N_11347,N_11168,N_11138);
nor U11348 (N_11348,N_11123,N_11149);
nand U11349 (N_11349,N_11092,N_11198);
and U11350 (N_11350,N_11031,N_11089);
or U11351 (N_11351,N_11092,N_11081);
and U11352 (N_11352,N_11048,N_11197);
nand U11353 (N_11353,N_11191,N_11173);
xnor U11354 (N_11354,N_11026,N_11182);
or U11355 (N_11355,N_11194,N_11092);
nor U11356 (N_11356,N_11171,N_11185);
and U11357 (N_11357,N_11009,N_11142);
xnor U11358 (N_11358,N_11109,N_11081);
and U11359 (N_11359,N_11069,N_11102);
or U11360 (N_11360,N_11068,N_11154);
and U11361 (N_11361,N_11037,N_11157);
and U11362 (N_11362,N_11014,N_11051);
xnor U11363 (N_11363,N_11083,N_11014);
nor U11364 (N_11364,N_11134,N_11136);
and U11365 (N_11365,N_11033,N_11074);
nor U11366 (N_11366,N_11112,N_11152);
or U11367 (N_11367,N_11123,N_11124);
nor U11368 (N_11368,N_11129,N_11109);
nor U11369 (N_11369,N_11027,N_11114);
nor U11370 (N_11370,N_11097,N_11194);
nand U11371 (N_11371,N_11158,N_11107);
xnor U11372 (N_11372,N_11129,N_11166);
nor U11373 (N_11373,N_11012,N_11199);
or U11374 (N_11374,N_11109,N_11194);
or U11375 (N_11375,N_11120,N_11161);
nor U11376 (N_11376,N_11093,N_11103);
and U11377 (N_11377,N_11141,N_11177);
nand U11378 (N_11378,N_11170,N_11094);
or U11379 (N_11379,N_11151,N_11126);
or U11380 (N_11380,N_11037,N_11066);
nand U11381 (N_11381,N_11155,N_11030);
nand U11382 (N_11382,N_11151,N_11044);
nand U11383 (N_11383,N_11060,N_11068);
or U11384 (N_11384,N_11070,N_11145);
nor U11385 (N_11385,N_11193,N_11148);
nor U11386 (N_11386,N_11155,N_11185);
xnor U11387 (N_11387,N_11119,N_11059);
nor U11388 (N_11388,N_11057,N_11017);
and U11389 (N_11389,N_11121,N_11007);
and U11390 (N_11390,N_11084,N_11051);
nor U11391 (N_11391,N_11190,N_11137);
and U11392 (N_11392,N_11025,N_11049);
or U11393 (N_11393,N_11197,N_11185);
and U11394 (N_11394,N_11060,N_11156);
nor U11395 (N_11395,N_11198,N_11133);
nand U11396 (N_11396,N_11083,N_11049);
nor U11397 (N_11397,N_11065,N_11168);
nand U11398 (N_11398,N_11069,N_11183);
nor U11399 (N_11399,N_11046,N_11119);
nand U11400 (N_11400,N_11268,N_11346);
nand U11401 (N_11401,N_11306,N_11328);
or U11402 (N_11402,N_11333,N_11313);
or U11403 (N_11403,N_11315,N_11254);
xnor U11404 (N_11404,N_11266,N_11275);
xor U11405 (N_11405,N_11235,N_11335);
or U11406 (N_11406,N_11385,N_11301);
xor U11407 (N_11407,N_11290,N_11365);
or U11408 (N_11408,N_11340,N_11256);
or U11409 (N_11409,N_11317,N_11241);
xnor U11410 (N_11410,N_11223,N_11305);
nand U11411 (N_11411,N_11259,N_11386);
nand U11412 (N_11412,N_11249,N_11347);
nand U11413 (N_11413,N_11248,N_11334);
and U11414 (N_11414,N_11286,N_11208);
or U11415 (N_11415,N_11279,N_11281);
nor U11416 (N_11416,N_11211,N_11360);
nor U11417 (N_11417,N_11350,N_11204);
xnor U11418 (N_11418,N_11302,N_11273);
and U11419 (N_11419,N_11250,N_11314);
nand U11420 (N_11420,N_11376,N_11351);
or U11421 (N_11421,N_11338,N_11319);
nor U11422 (N_11422,N_11221,N_11252);
nor U11423 (N_11423,N_11382,N_11206);
or U11424 (N_11424,N_11298,N_11258);
xor U11425 (N_11425,N_11332,N_11261);
or U11426 (N_11426,N_11312,N_11354);
nand U11427 (N_11427,N_11231,N_11348);
and U11428 (N_11428,N_11209,N_11371);
nand U11429 (N_11429,N_11295,N_11270);
xnor U11430 (N_11430,N_11368,N_11205);
nand U11431 (N_11431,N_11228,N_11329);
or U11432 (N_11432,N_11233,N_11239);
and U11433 (N_11433,N_11276,N_11324);
or U11434 (N_11434,N_11242,N_11336);
xor U11435 (N_11435,N_11257,N_11307);
nand U11436 (N_11436,N_11269,N_11323);
and U11437 (N_11437,N_11391,N_11245);
and U11438 (N_11438,N_11215,N_11381);
xnor U11439 (N_11439,N_11364,N_11217);
nor U11440 (N_11440,N_11264,N_11311);
nor U11441 (N_11441,N_11395,N_11299);
nor U11442 (N_11442,N_11237,N_11247);
or U11443 (N_11443,N_11296,N_11331);
nand U11444 (N_11444,N_11370,N_11358);
or U11445 (N_11445,N_11308,N_11253);
xor U11446 (N_11446,N_11234,N_11289);
xnor U11447 (N_11447,N_11397,N_11322);
xor U11448 (N_11448,N_11352,N_11251);
or U11449 (N_11449,N_11341,N_11325);
nor U11450 (N_11450,N_11292,N_11272);
nand U11451 (N_11451,N_11377,N_11262);
nand U11452 (N_11452,N_11398,N_11310);
xnor U11453 (N_11453,N_11379,N_11366);
nor U11454 (N_11454,N_11203,N_11297);
nand U11455 (N_11455,N_11384,N_11246);
or U11456 (N_11456,N_11349,N_11287);
nor U11457 (N_11457,N_11339,N_11359);
nor U11458 (N_11458,N_11271,N_11316);
nand U11459 (N_11459,N_11399,N_11390);
xor U11460 (N_11460,N_11355,N_11378);
nor U11461 (N_11461,N_11300,N_11243);
and U11462 (N_11462,N_11274,N_11367);
or U11463 (N_11463,N_11222,N_11214);
nand U11464 (N_11464,N_11294,N_11232);
nand U11465 (N_11465,N_11387,N_11212);
xor U11466 (N_11466,N_11229,N_11219);
nand U11467 (N_11467,N_11230,N_11200);
xnor U11468 (N_11468,N_11374,N_11369);
xor U11469 (N_11469,N_11330,N_11284);
or U11470 (N_11470,N_11383,N_11394);
xnor U11471 (N_11471,N_11373,N_11362);
nor U11472 (N_11472,N_11201,N_11388);
or U11473 (N_11473,N_11216,N_11285);
nand U11474 (N_11474,N_11327,N_11320);
nand U11475 (N_11475,N_11260,N_11380);
nor U11476 (N_11476,N_11282,N_11396);
nor U11477 (N_11477,N_11356,N_11240);
xor U11478 (N_11478,N_11353,N_11218);
and U11479 (N_11479,N_11226,N_11337);
nor U11480 (N_11480,N_11321,N_11357);
and U11481 (N_11481,N_11342,N_11304);
or U11482 (N_11482,N_11263,N_11363);
nand U11483 (N_11483,N_11202,N_11227);
xor U11484 (N_11484,N_11344,N_11225);
xor U11485 (N_11485,N_11280,N_11244);
and U11486 (N_11486,N_11375,N_11293);
nand U11487 (N_11487,N_11291,N_11326);
xor U11488 (N_11488,N_11283,N_11278);
and U11489 (N_11489,N_11303,N_11345);
or U11490 (N_11490,N_11255,N_11343);
xor U11491 (N_11491,N_11267,N_11288);
and U11492 (N_11492,N_11277,N_11309);
and U11493 (N_11493,N_11393,N_11213);
nor U11494 (N_11494,N_11265,N_11210);
nand U11495 (N_11495,N_11207,N_11392);
nor U11496 (N_11496,N_11389,N_11372);
nor U11497 (N_11497,N_11361,N_11318);
or U11498 (N_11498,N_11238,N_11224);
xor U11499 (N_11499,N_11220,N_11236);
and U11500 (N_11500,N_11365,N_11227);
nor U11501 (N_11501,N_11303,N_11259);
nand U11502 (N_11502,N_11304,N_11340);
xnor U11503 (N_11503,N_11357,N_11325);
nand U11504 (N_11504,N_11342,N_11343);
or U11505 (N_11505,N_11347,N_11225);
or U11506 (N_11506,N_11312,N_11365);
or U11507 (N_11507,N_11260,N_11362);
nor U11508 (N_11508,N_11224,N_11383);
nand U11509 (N_11509,N_11204,N_11384);
nor U11510 (N_11510,N_11240,N_11380);
or U11511 (N_11511,N_11253,N_11228);
nor U11512 (N_11512,N_11269,N_11394);
and U11513 (N_11513,N_11357,N_11246);
xnor U11514 (N_11514,N_11216,N_11207);
and U11515 (N_11515,N_11252,N_11376);
and U11516 (N_11516,N_11392,N_11208);
nor U11517 (N_11517,N_11229,N_11210);
or U11518 (N_11518,N_11307,N_11228);
or U11519 (N_11519,N_11287,N_11248);
nor U11520 (N_11520,N_11393,N_11312);
xnor U11521 (N_11521,N_11268,N_11343);
nand U11522 (N_11522,N_11339,N_11297);
xnor U11523 (N_11523,N_11377,N_11225);
nor U11524 (N_11524,N_11399,N_11369);
xnor U11525 (N_11525,N_11241,N_11285);
nor U11526 (N_11526,N_11398,N_11362);
and U11527 (N_11527,N_11254,N_11380);
or U11528 (N_11528,N_11248,N_11339);
or U11529 (N_11529,N_11365,N_11358);
xnor U11530 (N_11530,N_11201,N_11336);
and U11531 (N_11531,N_11284,N_11379);
nand U11532 (N_11532,N_11295,N_11378);
nand U11533 (N_11533,N_11302,N_11201);
nand U11534 (N_11534,N_11298,N_11229);
or U11535 (N_11535,N_11328,N_11301);
nor U11536 (N_11536,N_11359,N_11249);
nor U11537 (N_11537,N_11395,N_11367);
nor U11538 (N_11538,N_11287,N_11230);
and U11539 (N_11539,N_11354,N_11255);
and U11540 (N_11540,N_11260,N_11303);
nand U11541 (N_11541,N_11247,N_11381);
nand U11542 (N_11542,N_11303,N_11285);
and U11543 (N_11543,N_11289,N_11260);
nor U11544 (N_11544,N_11349,N_11270);
nand U11545 (N_11545,N_11333,N_11271);
nor U11546 (N_11546,N_11300,N_11266);
xor U11547 (N_11547,N_11211,N_11393);
or U11548 (N_11548,N_11323,N_11359);
nor U11549 (N_11549,N_11271,N_11289);
or U11550 (N_11550,N_11346,N_11324);
or U11551 (N_11551,N_11391,N_11305);
xor U11552 (N_11552,N_11329,N_11207);
and U11553 (N_11553,N_11214,N_11343);
nand U11554 (N_11554,N_11373,N_11389);
nor U11555 (N_11555,N_11325,N_11397);
and U11556 (N_11556,N_11355,N_11210);
or U11557 (N_11557,N_11316,N_11347);
xnor U11558 (N_11558,N_11295,N_11362);
nor U11559 (N_11559,N_11376,N_11270);
nor U11560 (N_11560,N_11222,N_11299);
or U11561 (N_11561,N_11207,N_11286);
and U11562 (N_11562,N_11337,N_11369);
nand U11563 (N_11563,N_11232,N_11308);
nand U11564 (N_11564,N_11247,N_11291);
nor U11565 (N_11565,N_11240,N_11371);
xor U11566 (N_11566,N_11277,N_11246);
and U11567 (N_11567,N_11244,N_11393);
xor U11568 (N_11568,N_11281,N_11221);
nor U11569 (N_11569,N_11324,N_11323);
xor U11570 (N_11570,N_11240,N_11202);
nand U11571 (N_11571,N_11258,N_11334);
xnor U11572 (N_11572,N_11399,N_11275);
and U11573 (N_11573,N_11311,N_11223);
nor U11574 (N_11574,N_11269,N_11253);
and U11575 (N_11575,N_11277,N_11396);
nand U11576 (N_11576,N_11277,N_11385);
nor U11577 (N_11577,N_11299,N_11295);
xnor U11578 (N_11578,N_11369,N_11263);
xor U11579 (N_11579,N_11262,N_11203);
and U11580 (N_11580,N_11206,N_11259);
nor U11581 (N_11581,N_11398,N_11387);
or U11582 (N_11582,N_11361,N_11385);
nor U11583 (N_11583,N_11200,N_11270);
or U11584 (N_11584,N_11326,N_11223);
and U11585 (N_11585,N_11326,N_11233);
and U11586 (N_11586,N_11351,N_11395);
xnor U11587 (N_11587,N_11378,N_11213);
nor U11588 (N_11588,N_11232,N_11399);
xnor U11589 (N_11589,N_11200,N_11307);
or U11590 (N_11590,N_11268,N_11334);
xor U11591 (N_11591,N_11222,N_11355);
xor U11592 (N_11592,N_11229,N_11323);
xor U11593 (N_11593,N_11388,N_11392);
and U11594 (N_11594,N_11294,N_11239);
and U11595 (N_11595,N_11386,N_11347);
nand U11596 (N_11596,N_11248,N_11391);
nor U11597 (N_11597,N_11221,N_11236);
nand U11598 (N_11598,N_11310,N_11304);
and U11599 (N_11599,N_11252,N_11310);
and U11600 (N_11600,N_11402,N_11438);
and U11601 (N_11601,N_11563,N_11419);
xnor U11602 (N_11602,N_11595,N_11592);
or U11603 (N_11603,N_11479,N_11467);
and U11604 (N_11604,N_11437,N_11581);
or U11605 (N_11605,N_11526,N_11527);
nand U11606 (N_11606,N_11593,N_11544);
nor U11607 (N_11607,N_11520,N_11597);
xnor U11608 (N_11608,N_11589,N_11497);
nor U11609 (N_11609,N_11405,N_11401);
xnor U11610 (N_11610,N_11456,N_11586);
nor U11611 (N_11611,N_11484,N_11573);
nand U11612 (N_11612,N_11599,N_11548);
and U11613 (N_11613,N_11558,N_11473);
or U11614 (N_11614,N_11511,N_11565);
xor U11615 (N_11615,N_11491,N_11449);
xnor U11616 (N_11616,N_11461,N_11412);
xor U11617 (N_11617,N_11471,N_11427);
xnor U11618 (N_11618,N_11505,N_11448);
and U11619 (N_11619,N_11521,N_11553);
xnor U11620 (N_11620,N_11556,N_11441);
nor U11621 (N_11621,N_11578,N_11562);
nand U11622 (N_11622,N_11570,N_11429);
xor U11623 (N_11623,N_11434,N_11446);
and U11624 (N_11624,N_11410,N_11583);
nand U11625 (N_11625,N_11470,N_11535);
or U11626 (N_11626,N_11546,N_11481);
or U11627 (N_11627,N_11557,N_11406);
and U11628 (N_11628,N_11504,N_11569);
nor U11629 (N_11629,N_11492,N_11432);
xor U11630 (N_11630,N_11460,N_11512);
and U11631 (N_11631,N_11494,N_11502);
nor U11632 (N_11632,N_11537,N_11483);
or U11633 (N_11633,N_11571,N_11580);
xor U11634 (N_11634,N_11525,N_11472);
and U11635 (N_11635,N_11478,N_11498);
xor U11636 (N_11636,N_11503,N_11531);
nor U11637 (N_11637,N_11561,N_11555);
xnor U11638 (N_11638,N_11407,N_11591);
xor U11639 (N_11639,N_11513,N_11480);
xor U11640 (N_11640,N_11530,N_11559);
nor U11641 (N_11641,N_11543,N_11426);
and U11642 (N_11642,N_11564,N_11485);
or U11643 (N_11643,N_11457,N_11540);
nor U11644 (N_11644,N_11487,N_11482);
and U11645 (N_11645,N_11545,N_11445);
and U11646 (N_11646,N_11418,N_11598);
nor U11647 (N_11647,N_11428,N_11509);
or U11648 (N_11648,N_11510,N_11463);
or U11649 (N_11649,N_11524,N_11550);
nor U11650 (N_11650,N_11590,N_11422);
nor U11651 (N_11651,N_11420,N_11501);
nand U11652 (N_11652,N_11452,N_11495);
nand U11653 (N_11653,N_11572,N_11435);
and U11654 (N_11654,N_11514,N_11596);
and U11655 (N_11655,N_11486,N_11538);
and U11656 (N_11656,N_11587,N_11518);
nand U11657 (N_11657,N_11541,N_11574);
nor U11658 (N_11658,N_11508,N_11517);
nand U11659 (N_11659,N_11417,N_11500);
nor U11660 (N_11660,N_11400,N_11560);
and U11661 (N_11661,N_11489,N_11408);
and U11662 (N_11662,N_11549,N_11421);
nor U11663 (N_11663,N_11442,N_11522);
nor U11664 (N_11664,N_11477,N_11507);
or U11665 (N_11665,N_11454,N_11499);
and U11666 (N_11666,N_11488,N_11403);
or U11667 (N_11667,N_11575,N_11585);
nand U11668 (N_11668,N_11528,N_11424);
or U11669 (N_11669,N_11566,N_11551);
xnor U11670 (N_11670,N_11447,N_11431);
nand U11671 (N_11671,N_11413,N_11415);
nor U11672 (N_11672,N_11425,N_11519);
nor U11673 (N_11673,N_11529,N_11423);
and U11674 (N_11674,N_11547,N_11411);
nor U11675 (N_11675,N_11433,N_11542);
or U11676 (N_11676,N_11462,N_11490);
or U11677 (N_11677,N_11523,N_11496);
or U11678 (N_11678,N_11516,N_11453);
or U11679 (N_11679,N_11539,N_11458);
nand U11680 (N_11680,N_11582,N_11443);
nor U11681 (N_11681,N_11451,N_11469);
nor U11682 (N_11682,N_11588,N_11464);
nor U11683 (N_11683,N_11536,N_11552);
xnor U11684 (N_11684,N_11534,N_11594);
xnor U11685 (N_11685,N_11554,N_11568);
xnor U11686 (N_11686,N_11404,N_11532);
or U11687 (N_11687,N_11576,N_11567);
xor U11688 (N_11688,N_11533,N_11439);
or U11689 (N_11689,N_11430,N_11579);
and U11690 (N_11690,N_11465,N_11577);
xnor U11691 (N_11691,N_11474,N_11459);
or U11692 (N_11692,N_11436,N_11416);
nor U11693 (N_11693,N_11455,N_11414);
nor U11694 (N_11694,N_11409,N_11584);
and U11695 (N_11695,N_11506,N_11493);
nor U11696 (N_11696,N_11475,N_11515);
xor U11697 (N_11697,N_11468,N_11476);
xor U11698 (N_11698,N_11450,N_11466);
or U11699 (N_11699,N_11440,N_11444);
and U11700 (N_11700,N_11464,N_11452);
xor U11701 (N_11701,N_11464,N_11582);
and U11702 (N_11702,N_11402,N_11567);
nor U11703 (N_11703,N_11486,N_11487);
and U11704 (N_11704,N_11402,N_11425);
nor U11705 (N_11705,N_11486,N_11591);
nor U11706 (N_11706,N_11550,N_11576);
and U11707 (N_11707,N_11513,N_11545);
xnor U11708 (N_11708,N_11529,N_11450);
nor U11709 (N_11709,N_11574,N_11536);
nor U11710 (N_11710,N_11592,N_11520);
or U11711 (N_11711,N_11549,N_11418);
and U11712 (N_11712,N_11563,N_11530);
nand U11713 (N_11713,N_11424,N_11548);
and U11714 (N_11714,N_11569,N_11455);
and U11715 (N_11715,N_11502,N_11477);
or U11716 (N_11716,N_11539,N_11594);
xnor U11717 (N_11717,N_11482,N_11560);
and U11718 (N_11718,N_11467,N_11494);
nor U11719 (N_11719,N_11583,N_11440);
nor U11720 (N_11720,N_11569,N_11537);
xor U11721 (N_11721,N_11467,N_11490);
xor U11722 (N_11722,N_11425,N_11433);
nand U11723 (N_11723,N_11447,N_11443);
and U11724 (N_11724,N_11500,N_11543);
xor U11725 (N_11725,N_11440,N_11484);
nor U11726 (N_11726,N_11401,N_11477);
nand U11727 (N_11727,N_11454,N_11561);
nor U11728 (N_11728,N_11513,N_11590);
or U11729 (N_11729,N_11424,N_11503);
xnor U11730 (N_11730,N_11446,N_11599);
or U11731 (N_11731,N_11592,N_11449);
or U11732 (N_11732,N_11593,N_11545);
or U11733 (N_11733,N_11598,N_11442);
or U11734 (N_11734,N_11543,N_11438);
or U11735 (N_11735,N_11527,N_11406);
or U11736 (N_11736,N_11586,N_11429);
or U11737 (N_11737,N_11547,N_11597);
nand U11738 (N_11738,N_11550,N_11435);
nand U11739 (N_11739,N_11489,N_11516);
and U11740 (N_11740,N_11427,N_11477);
xor U11741 (N_11741,N_11562,N_11488);
xor U11742 (N_11742,N_11507,N_11429);
or U11743 (N_11743,N_11597,N_11489);
nor U11744 (N_11744,N_11405,N_11531);
nand U11745 (N_11745,N_11484,N_11414);
nor U11746 (N_11746,N_11480,N_11515);
nand U11747 (N_11747,N_11445,N_11410);
nor U11748 (N_11748,N_11421,N_11428);
nor U11749 (N_11749,N_11563,N_11464);
and U11750 (N_11750,N_11468,N_11560);
xor U11751 (N_11751,N_11518,N_11553);
and U11752 (N_11752,N_11468,N_11512);
nand U11753 (N_11753,N_11487,N_11450);
nor U11754 (N_11754,N_11537,N_11447);
and U11755 (N_11755,N_11455,N_11581);
nand U11756 (N_11756,N_11494,N_11456);
or U11757 (N_11757,N_11563,N_11411);
nand U11758 (N_11758,N_11424,N_11515);
nand U11759 (N_11759,N_11404,N_11575);
or U11760 (N_11760,N_11566,N_11425);
nor U11761 (N_11761,N_11461,N_11538);
and U11762 (N_11762,N_11545,N_11469);
or U11763 (N_11763,N_11448,N_11526);
nand U11764 (N_11764,N_11455,N_11400);
or U11765 (N_11765,N_11535,N_11478);
and U11766 (N_11766,N_11449,N_11439);
xnor U11767 (N_11767,N_11449,N_11424);
nand U11768 (N_11768,N_11460,N_11476);
nand U11769 (N_11769,N_11557,N_11512);
nor U11770 (N_11770,N_11452,N_11553);
nor U11771 (N_11771,N_11510,N_11563);
or U11772 (N_11772,N_11560,N_11537);
and U11773 (N_11773,N_11506,N_11448);
and U11774 (N_11774,N_11581,N_11498);
nor U11775 (N_11775,N_11535,N_11508);
xnor U11776 (N_11776,N_11424,N_11436);
nand U11777 (N_11777,N_11503,N_11550);
nor U11778 (N_11778,N_11444,N_11582);
and U11779 (N_11779,N_11403,N_11411);
nor U11780 (N_11780,N_11522,N_11507);
nand U11781 (N_11781,N_11551,N_11581);
or U11782 (N_11782,N_11428,N_11584);
xor U11783 (N_11783,N_11452,N_11404);
nor U11784 (N_11784,N_11428,N_11534);
nand U11785 (N_11785,N_11551,N_11574);
xnor U11786 (N_11786,N_11493,N_11588);
and U11787 (N_11787,N_11404,N_11523);
nor U11788 (N_11788,N_11524,N_11533);
xor U11789 (N_11789,N_11533,N_11583);
and U11790 (N_11790,N_11485,N_11478);
or U11791 (N_11791,N_11519,N_11451);
and U11792 (N_11792,N_11417,N_11557);
and U11793 (N_11793,N_11485,N_11493);
or U11794 (N_11794,N_11502,N_11511);
nor U11795 (N_11795,N_11527,N_11458);
nor U11796 (N_11796,N_11591,N_11552);
nand U11797 (N_11797,N_11512,N_11491);
and U11798 (N_11798,N_11469,N_11407);
nor U11799 (N_11799,N_11421,N_11450);
or U11800 (N_11800,N_11796,N_11645);
xnor U11801 (N_11801,N_11607,N_11793);
nand U11802 (N_11802,N_11733,N_11627);
and U11803 (N_11803,N_11718,N_11771);
and U11804 (N_11804,N_11703,N_11695);
xor U11805 (N_11805,N_11656,N_11794);
nand U11806 (N_11806,N_11697,N_11610);
nor U11807 (N_11807,N_11626,N_11661);
xnor U11808 (N_11808,N_11777,N_11600);
nor U11809 (N_11809,N_11712,N_11609);
nand U11810 (N_11810,N_11784,N_11786);
nor U11811 (N_11811,N_11620,N_11705);
or U11812 (N_11812,N_11783,N_11633);
or U11813 (N_11813,N_11644,N_11662);
nand U11814 (N_11814,N_11778,N_11624);
xor U11815 (N_11815,N_11754,N_11650);
nand U11816 (N_11816,N_11734,N_11696);
nor U11817 (N_11817,N_11710,N_11728);
and U11818 (N_11818,N_11735,N_11757);
or U11819 (N_11819,N_11659,N_11779);
nor U11820 (N_11820,N_11789,N_11686);
and U11821 (N_11821,N_11640,N_11630);
and U11822 (N_11822,N_11635,N_11629);
or U11823 (N_11823,N_11719,N_11671);
nor U11824 (N_11824,N_11622,N_11688);
nand U11825 (N_11825,N_11660,N_11792);
nor U11826 (N_11826,N_11611,N_11738);
nor U11827 (N_11827,N_11722,N_11636);
nand U11828 (N_11828,N_11693,N_11670);
xnor U11829 (N_11829,N_11678,N_11724);
nand U11830 (N_11830,N_11727,N_11651);
nor U11831 (N_11831,N_11641,N_11603);
nor U11832 (N_11832,N_11788,N_11744);
or U11833 (N_11833,N_11745,N_11782);
or U11834 (N_11834,N_11787,N_11772);
nand U11835 (N_11835,N_11642,N_11648);
and U11836 (N_11836,N_11657,N_11785);
or U11837 (N_11837,N_11666,N_11691);
xor U11838 (N_11838,N_11692,N_11740);
nor U11839 (N_11839,N_11639,N_11653);
or U11840 (N_11840,N_11618,N_11752);
xor U11841 (N_11841,N_11658,N_11761);
or U11842 (N_11842,N_11760,N_11781);
and U11843 (N_11843,N_11720,N_11643);
and U11844 (N_11844,N_11677,N_11755);
xnor U11845 (N_11845,N_11773,N_11685);
and U11846 (N_11846,N_11619,N_11631);
and U11847 (N_11847,N_11751,N_11614);
or U11848 (N_11848,N_11654,N_11770);
or U11849 (N_11849,N_11775,N_11684);
and U11850 (N_11850,N_11725,N_11604);
nor U11851 (N_11851,N_11664,N_11743);
xor U11852 (N_11852,N_11665,N_11682);
nand U11853 (N_11853,N_11749,N_11759);
and U11854 (N_11854,N_11638,N_11681);
or U11855 (N_11855,N_11736,N_11732);
xor U11856 (N_11856,N_11742,N_11767);
or U11857 (N_11857,N_11780,N_11694);
nand U11858 (N_11858,N_11676,N_11737);
xnor U11859 (N_11859,N_11699,N_11790);
nor U11860 (N_11860,N_11704,N_11674);
and U11861 (N_11861,N_11608,N_11621);
nor U11862 (N_11862,N_11726,N_11702);
xnor U11863 (N_11863,N_11701,N_11700);
or U11864 (N_11864,N_11709,N_11669);
nand U11865 (N_11865,N_11748,N_11715);
or U11866 (N_11866,N_11762,N_11729);
xor U11867 (N_11867,N_11646,N_11713);
or U11868 (N_11868,N_11606,N_11628);
xor U11869 (N_11869,N_11690,N_11689);
nand U11870 (N_11870,N_11797,N_11675);
nor U11871 (N_11871,N_11764,N_11632);
nand U11872 (N_11872,N_11731,N_11663);
and U11873 (N_11873,N_11756,N_11680);
xnor U11874 (N_11874,N_11747,N_11679);
xnor U11875 (N_11875,N_11672,N_11776);
xor U11876 (N_11876,N_11714,N_11746);
nor U11877 (N_11877,N_11634,N_11617);
xnor U11878 (N_11878,N_11708,N_11774);
and U11879 (N_11879,N_11698,N_11687);
or U11880 (N_11880,N_11758,N_11766);
and U11881 (N_11881,N_11753,N_11798);
nor U11882 (N_11882,N_11706,N_11716);
nand U11883 (N_11883,N_11625,N_11765);
nand U11884 (N_11884,N_11605,N_11769);
or U11885 (N_11885,N_11717,N_11601);
xnor U11886 (N_11886,N_11750,N_11637);
or U11887 (N_11887,N_11795,N_11707);
xnor U11888 (N_11888,N_11623,N_11683);
nand U11889 (N_11889,N_11652,N_11768);
and U11890 (N_11890,N_11612,N_11655);
nor U11891 (N_11891,N_11730,N_11649);
and U11892 (N_11892,N_11613,N_11739);
nand U11893 (N_11893,N_11673,N_11616);
or U11894 (N_11894,N_11721,N_11602);
nor U11895 (N_11895,N_11668,N_11647);
xnor U11896 (N_11896,N_11791,N_11711);
nand U11897 (N_11897,N_11763,N_11723);
xor U11898 (N_11898,N_11615,N_11741);
nand U11899 (N_11899,N_11667,N_11799);
nand U11900 (N_11900,N_11604,N_11691);
or U11901 (N_11901,N_11669,N_11607);
xor U11902 (N_11902,N_11665,N_11650);
and U11903 (N_11903,N_11674,N_11652);
nor U11904 (N_11904,N_11729,N_11635);
and U11905 (N_11905,N_11669,N_11725);
nor U11906 (N_11906,N_11712,N_11701);
nand U11907 (N_11907,N_11666,N_11742);
and U11908 (N_11908,N_11743,N_11738);
nand U11909 (N_11909,N_11766,N_11734);
and U11910 (N_11910,N_11741,N_11602);
and U11911 (N_11911,N_11636,N_11672);
or U11912 (N_11912,N_11763,N_11608);
nand U11913 (N_11913,N_11790,N_11669);
and U11914 (N_11914,N_11730,N_11737);
xor U11915 (N_11915,N_11774,N_11768);
nor U11916 (N_11916,N_11738,N_11787);
xnor U11917 (N_11917,N_11733,N_11767);
or U11918 (N_11918,N_11600,N_11760);
and U11919 (N_11919,N_11678,N_11662);
and U11920 (N_11920,N_11608,N_11674);
nor U11921 (N_11921,N_11796,N_11758);
and U11922 (N_11922,N_11609,N_11661);
nor U11923 (N_11923,N_11709,N_11764);
and U11924 (N_11924,N_11703,N_11778);
and U11925 (N_11925,N_11755,N_11604);
nand U11926 (N_11926,N_11748,N_11721);
nand U11927 (N_11927,N_11776,N_11693);
nand U11928 (N_11928,N_11729,N_11666);
or U11929 (N_11929,N_11688,N_11705);
xor U11930 (N_11930,N_11711,N_11784);
nor U11931 (N_11931,N_11673,N_11660);
nand U11932 (N_11932,N_11753,N_11708);
xnor U11933 (N_11933,N_11658,N_11793);
nand U11934 (N_11934,N_11649,N_11719);
and U11935 (N_11935,N_11754,N_11646);
and U11936 (N_11936,N_11640,N_11739);
xor U11937 (N_11937,N_11759,N_11739);
nand U11938 (N_11938,N_11653,N_11685);
nand U11939 (N_11939,N_11693,N_11770);
xnor U11940 (N_11940,N_11771,N_11722);
nand U11941 (N_11941,N_11797,N_11672);
or U11942 (N_11942,N_11733,N_11641);
or U11943 (N_11943,N_11707,N_11659);
and U11944 (N_11944,N_11768,N_11677);
or U11945 (N_11945,N_11796,N_11772);
nor U11946 (N_11946,N_11794,N_11785);
or U11947 (N_11947,N_11734,N_11618);
nand U11948 (N_11948,N_11755,N_11733);
nor U11949 (N_11949,N_11746,N_11726);
or U11950 (N_11950,N_11775,N_11655);
and U11951 (N_11951,N_11684,N_11659);
and U11952 (N_11952,N_11712,N_11615);
or U11953 (N_11953,N_11654,N_11766);
and U11954 (N_11954,N_11734,N_11623);
nor U11955 (N_11955,N_11608,N_11645);
xor U11956 (N_11956,N_11647,N_11690);
and U11957 (N_11957,N_11720,N_11743);
nand U11958 (N_11958,N_11612,N_11724);
xnor U11959 (N_11959,N_11717,N_11778);
xor U11960 (N_11960,N_11671,N_11794);
nand U11961 (N_11961,N_11719,N_11672);
or U11962 (N_11962,N_11731,N_11677);
nand U11963 (N_11963,N_11650,N_11731);
and U11964 (N_11964,N_11753,N_11712);
nand U11965 (N_11965,N_11692,N_11707);
and U11966 (N_11966,N_11679,N_11726);
xnor U11967 (N_11967,N_11791,N_11600);
nor U11968 (N_11968,N_11638,N_11656);
or U11969 (N_11969,N_11661,N_11600);
and U11970 (N_11970,N_11708,N_11737);
xnor U11971 (N_11971,N_11648,N_11764);
nand U11972 (N_11972,N_11633,N_11625);
nor U11973 (N_11973,N_11673,N_11620);
or U11974 (N_11974,N_11679,N_11635);
nand U11975 (N_11975,N_11743,N_11650);
xnor U11976 (N_11976,N_11614,N_11631);
xnor U11977 (N_11977,N_11637,N_11660);
nor U11978 (N_11978,N_11686,N_11655);
and U11979 (N_11979,N_11632,N_11751);
nor U11980 (N_11980,N_11768,N_11723);
xor U11981 (N_11981,N_11601,N_11762);
xnor U11982 (N_11982,N_11767,N_11715);
or U11983 (N_11983,N_11715,N_11626);
xor U11984 (N_11984,N_11731,N_11781);
xnor U11985 (N_11985,N_11622,N_11725);
nor U11986 (N_11986,N_11666,N_11747);
nand U11987 (N_11987,N_11752,N_11700);
nor U11988 (N_11988,N_11724,N_11694);
xor U11989 (N_11989,N_11668,N_11793);
xnor U11990 (N_11990,N_11783,N_11688);
xor U11991 (N_11991,N_11623,N_11700);
xor U11992 (N_11992,N_11664,N_11678);
xnor U11993 (N_11993,N_11630,N_11762);
xnor U11994 (N_11994,N_11656,N_11767);
xor U11995 (N_11995,N_11698,N_11772);
xnor U11996 (N_11996,N_11797,N_11693);
and U11997 (N_11997,N_11713,N_11791);
nand U11998 (N_11998,N_11787,N_11710);
nor U11999 (N_11999,N_11776,N_11654);
or U12000 (N_12000,N_11862,N_11967);
nand U12001 (N_12001,N_11995,N_11952);
and U12002 (N_12002,N_11873,N_11980);
nor U12003 (N_12003,N_11885,N_11993);
nand U12004 (N_12004,N_11902,N_11963);
nand U12005 (N_12005,N_11845,N_11803);
and U12006 (N_12006,N_11867,N_11820);
xnor U12007 (N_12007,N_11932,N_11912);
nor U12008 (N_12008,N_11946,N_11988);
nand U12009 (N_12009,N_11954,N_11962);
xnor U12010 (N_12010,N_11865,N_11928);
xor U12011 (N_12011,N_11832,N_11838);
nor U12012 (N_12012,N_11859,N_11884);
and U12013 (N_12013,N_11921,N_11812);
and U12014 (N_12014,N_11828,N_11800);
xor U12015 (N_12015,N_11934,N_11856);
xor U12016 (N_12016,N_11807,N_11936);
xor U12017 (N_12017,N_11985,N_11805);
xnor U12018 (N_12018,N_11833,N_11931);
or U12019 (N_12019,N_11846,N_11907);
and U12020 (N_12020,N_11958,N_11910);
nor U12021 (N_12021,N_11919,N_11899);
nor U12022 (N_12022,N_11887,N_11965);
or U12023 (N_12023,N_11830,N_11900);
xor U12024 (N_12024,N_11864,N_11990);
nor U12025 (N_12025,N_11904,N_11829);
or U12026 (N_12026,N_11938,N_11827);
nand U12027 (N_12027,N_11999,N_11978);
nor U12028 (N_12028,N_11850,N_11986);
and U12029 (N_12029,N_11992,N_11964);
or U12030 (N_12030,N_11972,N_11969);
and U12031 (N_12031,N_11841,N_11960);
and U12032 (N_12032,N_11950,N_11863);
and U12033 (N_12033,N_11808,N_11976);
or U12034 (N_12034,N_11840,N_11888);
nor U12035 (N_12035,N_11903,N_11835);
xnor U12036 (N_12036,N_11922,N_11861);
xnor U12037 (N_12037,N_11806,N_11817);
xnor U12038 (N_12038,N_11870,N_11914);
or U12039 (N_12039,N_11983,N_11831);
and U12040 (N_12040,N_11918,N_11897);
nor U12041 (N_12041,N_11961,N_11891);
nor U12042 (N_12042,N_11948,N_11854);
xnor U12043 (N_12043,N_11804,N_11984);
and U12044 (N_12044,N_11809,N_11937);
xnor U12045 (N_12045,N_11896,N_11810);
or U12046 (N_12046,N_11957,N_11882);
xnor U12047 (N_12047,N_11947,N_11801);
nor U12048 (N_12048,N_11920,N_11927);
nand U12049 (N_12049,N_11945,N_11834);
xor U12050 (N_12050,N_11814,N_11869);
and U12051 (N_12051,N_11811,N_11822);
or U12052 (N_12052,N_11816,N_11959);
xor U12053 (N_12053,N_11973,N_11880);
xor U12054 (N_12054,N_11935,N_11839);
and U12055 (N_12055,N_11898,N_11956);
or U12056 (N_12056,N_11889,N_11943);
or U12057 (N_12057,N_11924,N_11824);
and U12058 (N_12058,N_11875,N_11979);
xnor U12059 (N_12059,N_11982,N_11901);
or U12060 (N_12060,N_11977,N_11930);
xor U12061 (N_12061,N_11975,N_11923);
xor U12062 (N_12062,N_11837,N_11929);
xor U12063 (N_12063,N_11966,N_11815);
xor U12064 (N_12064,N_11892,N_11877);
nor U12065 (N_12065,N_11908,N_11925);
nand U12066 (N_12066,N_11852,N_11953);
nor U12067 (N_12067,N_11941,N_11994);
nor U12068 (N_12068,N_11858,N_11853);
or U12069 (N_12069,N_11987,N_11886);
xnor U12070 (N_12070,N_11883,N_11917);
xnor U12071 (N_12071,N_11942,N_11848);
nor U12072 (N_12072,N_11951,N_11971);
or U12073 (N_12073,N_11872,N_11968);
and U12074 (N_12074,N_11868,N_11989);
and U12075 (N_12075,N_11851,N_11847);
and U12076 (N_12076,N_11855,N_11916);
xnor U12077 (N_12077,N_11876,N_11844);
nor U12078 (N_12078,N_11939,N_11915);
nand U12079 (N_12079,N_11836,N_11895);
xor U12080 (N_12080,N_11906,N_11821);
nor U12081 (N_12081,N_11860,N_11991);
nand U12082 (N_12082,N_11823,N_11911);
and U12083 (N_12083,N_11997,N_11881);
nor U12084 (N_12084,N_11940,N_11818);
xor U12085 (N_12085,N_11874,N_11949);
and U12086 (N_12086,N_11825,N_11998);
and U12087 (N_12087,N_11857,N_11819);
nand U12088 (N_12088,N_11955,N_11944);
xor U12089 (N_12089,N_11879,N_11878);
nor U12090 (N_12090,N_11813,N_11866);
nand U12091 (N_12091,N_11849,N_11842);
xor U12092 (N_12092,N_11996,N_11893);
xnor U12093 (N_12093,N_11905,N_11926);
or U12094 (N_12094,N_11890,N_11826);
nand U12095 (N_12095,N_11802,N_11933);
xnor U12096 (N_12096,N_11843,N_11913);
or U12097 (N_12097,N_11909,N_11974);
nor U12098 (N_12098,N_11981,N_11970);
and U12099 (N_12099,N_11871,N_11894);
xor U12100 (N_12100,N_11820,N_11910);
xnor U12101 (N_12101,N_11979,N_11882);
nor U12102 (N_12102,N_11850,N_11992);
nand U12103 (N_12103,N_11991,N_11816);
xor U12104 (N_12104,N_11978,N_11845);
nand U12105 (N_12105,N_11948,N_11879);
xor U12106 (N_12106,N_11965,N_11809);
xnor U12107 (N_12107,N_11804,N_11945);
xor U12108 (N_12108,N_11995,N_11942);
nand U12109 (N_12109,N_11993,N_11882);
or U12110 (N_12110,N_11878,N_11942);
and U12111 (N_12111,N_11847,N_11883);
nand U12112 (N_12112,N_11968,N_11929);
and U12113 (N_12113,N_11815,N_11805);
xnor U12114 (N_12114,N_11986,N_11916);
and U12115 (N_12115,N_11880,N_11897);
nor U12116 (N_12116,N_11946,N_11812);
and U12117 (N_12117,N_11985,N_11866);
or U12118 (N_12118,N_11958,N_11988);
or U12119 (N_12119,N_11823,N_11806);
and U12120 (N_12120,N_11862,N_11938);
nor U12121 (N_12121,N_11884,N_11985);
or U12122 (N_12122,N_11811,N_11802);
nand U12123 (N_12123,N_11936,N_11954);
xnor U12124 (N_12124,N_11854,N_11810);
and U12125 (N_12125,N_11886,N_11883);
and U12126 (N_12126,N_11817,N_11960);
nand U12127 (N_12127,N_11927,N_11810);
xor U12128 (N_12128,N_11936,N_11814);
xor U12129 (N_12129,N_11889,N_11869);
or U12130 (N_12130,N_11976,N_11809);
nand U12131 (N_12131,N_11950,N_11882);
and U12132 (N_12132,N_11836,N_11973);
or U12133 (N_12133,N_11923,N_11981);
or U12134 (N_12134,N_11882,N_11821);
and U12135 (N_12135,N_11802,N_11827);
nand U12136 (N_12136,N_11975,N_11892);
and U12137 (N_12137,N_11933,N_11874);
nand U12138 (N_12138,N_11835,N_11946);
nor U12139 (N_12139,N_11939,N_11916);
nor U12140 (N_12140,N_11834,N_11993);
nand U12141 (N_12141,N_11851,N_11814);
xnor U12142 (N_12142,N_11855,N_11841);
xor U12143 (N_12143,N_11838,N_11830);
xor U12144 (N_12144,N_11951,N_11948);
and U12145 (N_12145,N_11821,N_11956);
nor U12146 (N_12146,N_11976,N_11843);
and U12147 (N_12147,N_11867,N_11986);
nand U12148 (N_12148,N_11952,N_11802);
nor U12149 (N_12149,N_11844,N_11809);
and U12150 (N_12150,N_11987,N_11859);
nor U12151 (N_12151,N_11974,N_11884);
nor U12152 (N_12152,N_11896,N_11940);
and U12153 (N_12153,N_11993,N_11864);
and U12154 (N_12154,N_11976,N_11837);
nor U12155 (N_12155,N_11814,N_11957);
and U12156 (N_12156,N_11938,N_11858);
or U12157 (N_12157,N_11942,N_11921);
nand U12158 (N_12158,N_11821,N_11800);
and U12159 (N_12159,N_11873,N_11999);
or U12160 (N_12160,N_11808,N_11997);
xor U12161 (N_12161,N_11860,N_11936);
nand U12162 (N_12162,N_11836,N_11845);
and U12163 (N_12163,N_11992,N_11853);
or U12164 (N_12164,N_11884,N_11977);
nand U12165 (N_12165,N_11853,N_11860);
nand U12166 (N_12166,N_11913,N_11829);
nor U12167 (N_12167,N_11872,N_11995);
and U12168 (N_12168,N_11952,N_11924);
nand U12169 (N_12169,N_11871,N_11815);
nand U12170 (N_12170,N_11820,N_11931);
nor U12171 (N_12171,N_11875,N_11858);
and U12172 (N_12172,N_11960,N_11839);
nor U12173 (N_12173,N_11928,N_11866);
nor U12174 (N_12174,N_11947,N_11887);
or U12175 (N_12175,N_11845,N_11940);
nand U12176 (N_12176,N_11921,N_11875);
or U12177 (N_12177,N_11987,N_11944);
nor U12178 (N_12178,N_11864,N_11923);
or U12179 (N_12179,N_11956,N_11803);
xor U12180 (N_12180,N_11881,N_11952);
xnor U12181 (N_12181,N_11815,N_11901);
or U12182 (N_12182,N_11901,N_11911);
nor U12183 (N_12183,N_11931,N_11840);
xor U12184 (N_12184,N_11855,N_11928);
nor U12185 (N_12185,N_11834,N_11957);
and U12186 (N_12186,N_11851,N_11914);
nor U12187 (N_12187,N_11913,N_11832);
nor U12188 (N_12188,N_11901,N_11907);
and U12189 (N_12189,N_11833,N_11927);
or U12190 (N_12190,N_11948,N_11825);
nand U12191 (N_12191,N_11970,N_11858);
nand U12192 (N_12192,N_11873,N_11867);
xor U12193 (N_12193,N_11922,N_11972);
xnor U12194 (N_12194,N_11985,N_11907);
or U12195 (N_12195,N_11977,N_11823);
or U12196 (N_12196,N_11865,N_11921);
or U12197 (N_12197,N_11956,N_11808);
and U12198 (N_12198,N_11996,N_11828);
and U12199 (N_12199,N_11972,N_11858);
xor U12200 (N_12200,N_12190,N_12074);
nand U12201 (N_12201,N_12172,N_12091);
nand U12202 (N_12202,N_12192,N_12082);
and U12203 (N_12203,N_12046,N_12108);
xor U12204 (N_12204,N_12150,N_12007);
xnor U12205 (N_12205,N_12106,N_12038);
xnor U12206 (N_12206,N_12037,N_12017);
or U12207 (N_12207,N_12195,N_12128);
xor U12208 (N_12208,N_12054,N_12073);
nand U12209 (N_12209,N_12187,N_12080);
or U12210 (N_12210,N_12168,N_12121);
nor U12211 (N_12211,N_12133,N_12199);
nand U12212 (N_12212,N_12024,N_12023);
xnor U12213 (N_12213,N_12158,N_12065);
nor U12214 (N_12214,N_12105,N_12099);
nand U12215 (N_12215,N_12135,N_12022);
nor U12216 (N_12216,N_12160,N_12002);
xnor U12217 (N_12217,N_12039,N_12112);
xor U12218 (N_12218,N_12178,N_12020);
nor U12219 (N_12219,N_12173,N_12126);
or U12220 (N_12220,N_12120,N_12087);
nand U12221 (N_12221,N_12071,N_12010);
or U12222 (N_12222,N_12115,N_12095);
nand U12223 (N_12223,N_12101,N_12030);
nand U12224 (N_12224,N_12110,N_12185);
and U12225 (N_12225,N_12147,N_12097);
and U12226 (N_12226,N_12051,N_12182);
nand U12227 (N_12227,N_12067,N_12191);
xor U12228 (N_12228,N_12188,N_12033);
xor U12229 (N_12229,N_12040,N_12144);
and U12230 (N_12230,N_12155,N_12084);
and U12231 (N_12231,N_12053,N_12186);
or U12232 (N_12232,N_12181,N_12109);
nor U12233 (N_12233,N_12193,N_12124);
nor U12234 (N_12234,N_12148,N_12003);
nor U12235 (N_12235,N_12153,N_12163);
nand U12236 (N_12236,N_12011,N_12146);
and U12237 (N_12237,N_12090,N_12159);
xor U12238 (N_12238,N_12085,N_12130);
and U12239 (N_12239,N_12004,N_12117);
nand U12240 (N_12240,N_12131,N_12127);
and U12241 (N_12241,N_12025,N_12058);
nor U12242 (N_12242,N_12161,N_12092);
and U12243 (N_12243,N_12089,N_12012);
nor U12244 (N_12244,N_12122,N_12064);
xor U12245 (N_12245,N_12057,N_12139);
nor U12246 (N_12246,N_12183,N_12196);
or U12247 (N_12247,N_12170,N_12138);
xor U12248 (N_12248,N_12018,N_12140);
and U12249 (N_12249,N_12156,N_12048);
nand U12250 (N_12250,N_12098,N_12157);
xor U12251 (N_12251,N_12045,N_12145);
or U12252 (N_12252,N_12179,N_12102);
or U12253 (N_12253,N_12184,N_12069);
nor U12254 (N_12254,N_12151,N_12125);
and U12255 (N_12255,N_12119,N_12032);
nand U12256 (N_12256,N_12072,N_12169);
nand U12257 (N_12257,N_12197,N_12076);
and U12258 (N_12258,N_12044,N_12008);
nand U12259 (N_12259,N_12149,N_12165);
and U12260 (N_12260,N_12047,N_12118);
nor U12261 (N_12261,N_12198,N_12041);
nand U12262 (N_12262,N_12129,N_12001);
nor U12263 (N_12263,N_12083,N_12050);
or U12264 (N_12264,N_12021,N_12123);
xor U12265 (N_12265,N_12176,N_12049);
nand U12266 (N_12266,N_12094,N_12136);
xor U12267 (N_12267,N_12029,N_12060);
or U12268 (N_12268,N_12114,N_12175);
xor U12269 (N_12269,N_12162,N_12174);
xnor U12270 (N_12270,N_12068,N_12009);
nor U12271 (N_12271,N_12075,N_12061);
nor U12272 (N_12272,N_12035,N_12164);
xnor U12273 (N_12273,N_12107,N_12113);
or U12274 (N_12274,N_12152,N_12081);
nand U12275 (N_12275,N_12070,N_12189);
or U12276 (N_12276,N_12059,N_12042);
or U12277 (N_12277,N_12132,N_12103);
and U12278 (N_12278,N_12116,N_12078);
and U12279 (N_12279,N_12016,N_12015);
and U12280 (N_12280,N_12027,N_12052);
and U12281 (N_12281,N_12167,N_12180);
xor U12282 (N_12282,N_12194,N_12066);
nand U12283 (N_12283,N_12077,N_12031);
nand U12284 (N_12284,N_12134,N_12062);
or U12285 (N_12285,N_12056,N_12043);
or U12286 (N_12286,N_12019,N_12100);
nand U12287 (N_12287,N_12104,N_12079);
or U12288 (N_12288,N_12137,N_12154);
and U12289 (N_12289,N_12013,N_12036);
and U12290 (N_12290,N_12028,N_12142);
nand U12291 (N_12291,N_12000,N_12034);
nor U12292 (N_12292,N_12086,N_12111);
nor U12293 (N_12293,N_12177,N_12166);
and U12294 (N_12294,N_12141,N_12014);
xor U12295 (N_12295,N_12026,N_12093);
or U12296 (N_12296,N_12006,N_12096);
or U12297 (N_12297,N_12055,N_12088);
xor U12298 (N_12298,N_12171,N_12063);
nand U12299 (N_12299,N_12005,N_12143);
and U12300 (N_12300,N_12015,N_12061);
and U12301 (N_12301,N_12057,N_12140);
nand U12302 (N_12302,N_12140,N_12080);
and U12303 (N_12303,N_12184,N_12151);
or U12304 (N_12304,N_12031,N_12161);
nor U12305 (N_12305,N_12143,N_12051);
nand U12306 (N_12306,N_12182,N_12006);
nand U12307 (N_12307,N_12189,N_12075);
or U12308 (N_12308,N_12145,N_12001);
xnor U12309 (N_12309,N_12085,N_12050);
nand U12310 (N_12310,N_12013,N_12195);
or U12311 (N_12311,N_12044,N_12162);
nor U12312 (N_12312,N_12044,N_12197);
nand U12313 (N_12313,N_12066,N_12096);
or U12314 (N_12314,N_12114,N_12174);
nand U12315 (N_12315,N_12036,N_12019);
xor U12316 (N_12316,N_12184,N_12121);
and U12317 (N_12317,N_12028,N_12044);
nor U12318 (N_12318,N_12161,N_12029);
xnor U12319 (N_12319,N_12109,N_12050);
nand U12320 (N_12320,N_12092,N_12005);
nand U12321 (N_12321,N_12063,N_12175);
xor U12322 (N_12322,N_12090,N_12064);
or U12323 (N_12323,N_12076,N_12006);
or U12324 (N_12324,N_12009,N_12184);
or U12325 (N_12325,N_12149,N_12025);
or U12326 (N_12326,N_12094,N_12093);
or U12327 (N_12327,N_12150,N_12167);
nand U12328 (N_12328,N_12192,N_12104);
xor U12329 (N_12329,N_12059,N_12074);
and U12330 (N_12330,N_12023,N_12081);
nor U12331 (N_12331,N_12143,N_12096);
nor U12332 (N_12332,N_12104,N_12080);
and U12333 (N_12333,N_12175,N_12051);
xnor U12334 (N_12334,N_12006,N_12058);
nor U12335 (N_12335,N_12182,N_12113);
or U12336 (N_12336,N_12108,N_12164);
xor U12337 (N_12337,N_12042,N_12107);
or U12338 (N_12338,N_12156,N_12145);
nor U12339 (N_12339,N_12057,N_12120);
nor U12340 (N_12340,N_12053,N_12146);
nand U12341 (N_12341,N_12113,N_12004);
nand U12342 (N_12342,N_12125,N_12170);
or U12343 (N_12343,N_12150,N_12020);
and U12344 (N_12344,N_12076,N_12011);
nand U12345 (N_12345,N_12185,N_12129);
nor U12346 (N_12346,N_12178,N_12088);
nor U12347 (N_12347,N_12092,N_12159);
xnor U12348 (N_12348,N_12158,N_12086);
and U12349 (N_12349,N_12127,N_12099);
nor U12350 (N_12350,N_12100,N_12178);
and U12351 (N_12351,N_12023,N_12064);
or U12352 (N_12352,N_12030,N_12123);
nor U12353 (N_12353,N_12082,N_12183);
and U12354 (N_12354,N_12015,N_12089);
and U12355 (N_12355,N_12163,N_12123);
nand U12356 (N_12356,N_12185,N_12107);
and U12357 (N_12357,N_12146,N_12021);
xnor U12358 (N_12358,N_12138,N_12009);
nand U12359 (N_12359,N_12171,N_12001);
nand U12360 (N_12360,N_12035,N_12053);
or U12361 (N_12361,N_12142,N_12192);
or U12362 (N_12362,N_12050,N_12033);
or U12363 (N_12363,N_12031,N_12108);
or U12364 (N_12364,N_12187,N_12102);
nand U12365 (N_12365,N_12059,N_12115);
and U12366 (N_12366,N_12046,N_12024);
nor U12367 (N_12367,N_12022,N_12168);
xnor U12368 (N_12368,N_12163,N_12030);
xnor U12369 (N_12369,N_12017,N_12082);
xor U12370 (N_12370,N_12015,N_12050);
and U12371 (N_12371,N_12054,N_12113);
xor U12372 (N_12372,N_12068,N_12187);
nor U12373 (N_12373,N_12018,N_12051);
and U12374 (N_12374,N_12012,N_12137);
xnor U12375 (N_12375,N_12069,N_12102);
nor U12376 (N_12376,N_12188,N_12162);
and U12377 (N_12377,N_12094,N_12100);
xnor U12378 (N_12378,N_12040,N_12127);
xnor U12379 (N_12379,N_12127,N_12156);
nor U12380 (N_12380,N_12098,N_12125);
or U12381 (N_12381,N_12145,N_12051);
xnor U12382 (N_12382,N_12182,N_12164);
and U12383 (N_12383,N_12077,N_12037);
nor U12384 (N_12384,N_12075,N_12100);
or U12385 (N_12385,N_12062,N_12043);
and U12386 (N_12386,N_12158,N_12189);
and U12387 (N_12387,N_12126,N_12059);
or U12388 (N_12388,N_12051,N_12193);
nand U12389 (N_12389,N_12003,N_12095);
nand U12390 (N_12390,N_12065,N_12012);
and U12391 (N_12391,N_12027,N_12020);
nand U12392 (N_12392,N_12065,N_12035);
nand U12393 (N_12393,N_12169,N_12114);
xor U12394 (N_12394,N_12015,N_12116);
and U12395 (N_12395,N_12004,N_12094);
nor U12396 (N_12396,N_12101,N_12108);
nand U12397 (N_12397,N_12046,N_12002);
nor U12398 (N_12398,N_12111,N_12139);
or U12399 (N_12399,N_12149,N_12100);
and U12400 (N_12400,N_12236,N_12399);
and U12401 (N_12401,N_12345,N_12332);
nor U12402 (N_12402,N_12309,N_12256);
nand U12403 (N_12403,N_12348,N_12331);
xnor U12404 (N_12404,N_12229,N_12304);
nand U12405 (N_12405,N_12346,N_12206);
nand U12406 (N_12406,N_12214,N_12392);
xnor U12407 (N_12407,N_12370,N_12344);
and U12408 (N_12408,N_12360,N_12371);
nor U12409 (N_12409,N_12283,N_12209);
xor U12410 (N_12410,N_12245,N_12350);
nor U12411 (N_12411,N_12250,N_12340);
and U12412 (N_12412,N_12267,N_12203);
xor U12413 (N_12413,N_12217,N_12338);
or U12414 (N_12414,N_12367,N_12328);
and U12415 (N_12415,N_12326,N_12311);
or U12416 (N_12416,N_12204,N_12202);
nor U12417 (N_12417,N_12298,N_12231);
xnor U12418 (N_12418,N_12307,N_12211);
xnor U12419 (N_12419,N_12275,N_12270);
and U12420 (N_12420,N_12384,N_12366);
nor U12421 (N_12421,N_12276,N_12274);
or U12422 (N_12422,N_12335,N_12334);
and U12423 (N_12423,N_12244,N_12213);
or U12424 (N_12424,N_12354,N_12319);
nand U12425 (N_12425,N_12339,N_12258);
nor U12426 (N_12426,N_12385,N_12249);
nor U12427 (N_12427,N_12312,N_12296);
or U12428 (N_12428,N_12306,N_12329);
xnor U12429 (N_12429,N_12361,N_12308);
xor U12430 (N_12430,N_12232,N_12394);
nand U12431 (N_12431,N_12284,N_12260);
xnor U12432 (N_12432,N_12221,N_12246);
xor U12433 (N_12433,N_12321,N_12292);
or U12434 (N_12434,N_12286,N_12255);
xnor U12435 (N_12435,N_12356,N_12386);
xnor U12436 (N_12436,N_12397,N_12277);
or U12437 (N_12437,N_12281,N_12314);
nand U12438 (N_12438,N_12376,N_12337);
nor U12439 (N_12439,N_12240,N_12347);
or U12440 (N_12440,N_12271,N_12359);
nor U12441 (N_12441,N_12353,N_12374);
nand U12442 (N_12442,N_12342,N_12252);
nand U12443 (N_12443,N_12288,N_12238);
nand U12444 (N_12444,N_12282,N_12253);
xnor U12445 (N_12445,N_12272,N_12264);
xnor U12446 (N_12446,N_12382,N_12285);
and U12447 (N_12447,N_12222,N_12225);
nand U12448 (N_12448,N_12263,N_12302);
nand U12449 (N_12449,N_12218,N_12318);
or U12450 (N_12450,N_12220,N_12362);
nand U12451 (N_12451,N_12278,N_12317);
nand U12452 (N_12452,N_12320,N_12233);
nor U12453 (N_12453,N_12248,N_12259);
xor U12454 (N_12454,N_12310,N_12254);
nor U12455 (N_12455,N_12352,N_12216);
nand U12456 (N_12456,N_12303,N_12243);
nor U12457 (N_12457,N_12269,N_12294);
nand U12458 (N_12458,N_12235,N_12390);
nor U12459 (N_12459,N_12262,N_12389);
nor U12460 (N_12460,N_12230,N_12387);
or U12461 (N_12461,N_12379,N_12290);
nor U12462 (N_12462,N_12369,N_12299);
xnor U12463 (N_12463,N_12330,N_12372);
or U12464 (N_12464,N_12375,N_12393);
xnor U12465 (N_12465,N_12363,N_12313);
nand U12466 (N_12466,N_12242,N_12324);
or U12467 (N_12467,N_12223,N_12295);
and U12468 (N_12468,N_12381,N_12287);
or U12469 (N_12469,N_12391,N_12357);
or U12470 (N_12470,N_12323,N_12266);
nand U12471 (N_12471,N_12336,N_12279);
and U12472 (N_12472,N_12237,N_12200);
or U12473 (N_12473,N_12349,N_12273);
nor U12474 (N_12474,N_12293,N_12239);
and U12475 (N_12475,N_12378,N_12388);
nor U12476 (N_12476,N_12291,N_12343);
or U12477 (N_12477,N_12300,N_12224);
or U12478 (N_12478,N_12207,N_12355);
or U12479 (N_12479,N_12289,N_12398);
and U12480 (N_12480,N_12265,N_12201);
nor U12481 (N_12481,N_12212,N_12251);
nor U12482 (N_12482,N_12380,N_12341);
or U12483 (N_12483,N_12333,N_12297);
xor U12484 (N_12484,N_12268,N_12257);
and U12485 (N_12485,N_12365,N_12261);
and U12486 (N_12486,N_12247,N_12316);
or U12487 (N_12487,N_12301,N_12305);
or U12488 (N_12488,N_12358,N_12377);
and U12489 (N_12489,N_12368,N_12327);
xor U12490 (N_12490,N_12395,N_12208);
nor U12491 (N_12491,N_12227,N_12280);
nor U12492 (N_12492,N_12325,N_12351);
and U12493 (N_12493,N_12383,N_12226);
xnor U12494 (N_12494,N_12215,N_12373);
and U12495 (N_12495,N_12234,N_12205);
nand U12496 (N_12496,N_12210,N_12322);
and U12497 (N_12497,N_12315,N_12219);
nor U12498 (N_12498,N_12396,N_12364);
nand U12499 (N_12499,N_12228,N_12241);
nand U12500 (N_12500,N_12331,N_12352);
nor U12501 (N_12501,N_12243,N_12259);
xor U12502 (N_12502,N_12392,N_12383);
or U12503 (N_12503,N_12286,N_12246);
xnor U12504 (N_12504,N_12361,N_12337);
or U12505 (N_12505,N_12247,N_12324);
and U12506 (N_12506,N_12311,N_12393);
or U12507 (N_12507,N_12360,N_12243);
or U12508 (N_12508,N_12319,N_12225);
nand U12509 (N_12509,N_12215,N_12249);
or U12510 (N_12510,N_12382,N_12253);
nand U12511 (N_12511,N_12390,N_12303);
and U12512 (N_12512,N_12384,N_12297);
and U12513 (N_12513,N_12278,N_12283);
nand U12514 (N_12514,N_12226,N_12354);
xnor U12515 (N_12515,N_12292,N_12248);
nand U12516 (N_12516,N_12316,N_12366);
nor U12517 (N_12517,N_12359,N_12276);
and U12518 (N_12518,N_12308,N_12346);
or U12519 (N_12519,N_12206,N_12287);
nand U12520 (N_12520,N_12316,N_12389);
or U12521 (N_12521,N_12276,N_12202);
or U12522 (N_12522,N_12226,N_12396);
xnor U12523 (N_12523,N_12249,N_12307);
xnor U12524 (N_12524,N_12339,N_12315);
nand U12525 (N_12525,N_12206,N_12349);
xor U12526 (N_12526,N_12302,N_12218);
or U12527 (N_12527,N_12221,N_12345);
nand U12528 (N_12528,N_12315,N_12325);
and U12529 (N_12529,N_12204,N_12314);
nor U12530 (N_12530,N_12319,N_12340);
xor U12531 (N_12531,N_12362,N_12269);
nor U12532 (N_12532,N_12238,N_12296);
xnor U12533 (N_12533,N_12321,N_12218);
and U12534 (N_12534,N_12339,N_12245);
or U12535 (N_12535,N_12275,N_12209);
nand U12536 (N_12536,N_12352,N_12263);
xor U12537 (N_12537,N_12356,N_12387);
nor U12538 (N_12538,N_12367,N_12308);
and U12539 (N_12539,N_12284,N_12269);
nor U12540 (N_12540,N_12392,N_12290);
nand U12541 (N_12541,N_12362,N_12394);
and U12542 (N_12542,N_12273,N_12261);
or U12543 (N_12543,N_12232,N_12379);
and U12544 (N_12544,N_12224,N_12278);
and U12545 (N_12545,N_12273,N_12351);
and U12546 (N_12546,N_12351,N_12350);
nand U12547 (N_12547,N_12309,N_12255);
nand U12548 (N_12548,N_12234,N_12338);
or U12549 (N_12549,N_12281,N_12265);
or U12550 (N_12550,N_12308,N_12391);
nor U12551 (N_12551,N_12230,N_12225);
or U12552 (N_12552,N_12293,N_12299);
or U12553 (N_12553,N_12203,N_12239);
or U12554 (N_12554,N_12234,N_12317);
nand U12555 (N_12555,N_12238,N_12338);
or U12556 (N_12556,N_12257,N_12379);
nand U12557 (N_12557,N_12306,N_12275);
nand U12558 (N_12558,N_12202,N_12256);
nor U12559 (N_12559,N_12207,N_12391);
nor U12560 (N_12560,N_12338,N_12212);
xnor U12561 (N_12561,N_12272,N_12265);
nor U12562 (N_12562,N_12313,N_12299);
nand U12563 (N_12563,N_12278,N_12254);
and U12564 (N_12564,N_12360,N_12251);
or U12565 (N_12565,N_12243,N_12239);
nand U12566 (N_12566,N_12312,N_12392);
nand U12567 (N_12567,N_12274,N_12208);
nand U12568 (N_12568,N_12282,N_12399);
nand U12569 (N_12569,N_12363,N_12323);
nor U12570 (N_12570,N_12233,N_12355);
nor U12571 (N_12571,N_12245,N_12345);
and U12572 (N_12572,N_12247,N_12311);
xor U12573 (N_12573,N_12392,N_12266);
xor U12574 (N_12574,N_12352,N_12379);
nor U12575 (N_12575,N_12231,N_12305);
nor U12576 (N_12576,N_12343,N_12233);
or U12577 (N_12577,N_12364,N_12207);
nand U12578 (N_12578,N_12355,N_12336);
nor U12579 (N_12579,N_12314,N_12229);
nand U12580 (N_12580,N_12268,N_12215);
or U12581 (N_12581,N_12306,N_12334);
or U12582 (N_12582,N_12272,N_12299);
nand U12583 (N_12583,N_12379,N_12289);
and U12584 (N_12584,N_12254,N_12367);
and U12585 (N_12585,N_12367,N_12336);
and U12586 (N_12586,N_12259,N_12368);
nor U12587 (N_12587,N_12384,N_12335);
nand U12588 (N_12588,N_12232,N_12309);
or U12589 (N_12589,N_12215,N_12278);
nor U12590 (N_12590,N_12289,N_12247);
nor U12591 (N_12591,N_12366,N_12333);
nor U12592 (N_12592,N_12347,N_12282);
xnor U12593 (N_12593,N_12366,N_12335);
xnor U12594 (N_12594,N_12292,N_12329);
and U12595 (N_12595,N_12302,N_12219);
or U12596 (N_12596,N_12263,N_12248);
nand U12597 (N_12597,N_12263,N_12379);
xor U12598 (N_12598,N_12302,N_12227);
or U12599 (N_12599,N_12306,N_12205);
nor U12600 (N_12600,N_12429,N_12487);
xor U12601 (N_12601,N_12507,N_12420);
or U12602 (N_12602,N_12570,N_12529);
nand U12603 (N_12603,N_12588,N_12480);
or U12604 (N_12604,N_12556,N_12521);
xor U12605 (N_12605,N_12592,N_12539);
and U12606 (N_12606,N_12585,N_12542);
xor U12607 (N_12607,N_12426,N_12454);
nand U12608 (N_12608,N_12533,N_12575);
nor U12609 (N_12609,N_12477,N_12497);
xor U12610 (N_12610,N_12590,N_12442);
or U12611 (N_12611,N_12517,N_12560);
and U12612 (N_12612,N_12441,N_12464);
and U12613 (N_12613,N_12526,N_12433);
nand U12614 (N_12614,N_12485,N_12407);
and U12615 (N_12615,N_12536,N_12460);
nand U12616 (N_12616,N_12413,N_12565);
or U12617 (N_12617,N_12548,N_12427);
and U12618 (N_12618,N_12405,N_12523);
nor U12619 (N_12619,N_12597,N_12522);
nand U12620 (N_12620,N_12421,N_12409);
or U12621 (N_12621,N_12438,N_12567);
nor U12622 (N_12622,N_12532,N_12436);
nand U12623 (N_12623,N_12439,N_12538);
or U12624 (N_12624,N_12551,N_12596);
nand U12625 (N_12625,N_12492,N_12572);
nor U12626 (N_12626,N_12466,N_12525);
or U12627 (N_12627,N_12450,N_12555);
nand U12628 (N_12628,N_12453,N_12414);
or U12629 (N_12629,N_12554,N_12528);
and U12630 (N_12630,N_12591,N_12424);
xnor U12631 (N_12631,N_12490,N_12573);
and U12632 (N_12632,N_12550,N_12562);
nand U12633 (N_12633,N_12514,N_12474);
nand U12634 (N_12634,N_12440,N_12563);
nor U12635 (N_12635,N_12443,N_12534);
and U12636 (N_12636,N_12545,N_12465);
nand U12637 (N_12637,N_12401,N_12473);
nor U12638 (N_12638,N_12574,N_12559);
nand U12639 (N_12639,N_12584,N_12494);
nor U12640 (N_12640,N_12417,N_12557);
or U12641 (N_12641,N_12408,N_12520);
nor U12642 (N_12642,N_12411,N_12491);
xnor U12643 (N_12643,N_12552,N_12455);
and U12644 (N_12644,N_12541,N_12416);
or U12645 (N_12645,N_12484,N_12467);
nor U12646 (N_12646,N_12415,N_12505);
or U12647 (N_12647,N_12461,N_12568);
xnor U12648 (N_12648,N_12400,N_12457);
nor U12649 (N_12649,N_12459,N_12543);
and U12650 (N_12650,N_12499,N_12583);
and U12651 (N_12651,N_12403,N_12599);
and U12652 (N_12652,N_12462,N_12430);
nand U12653 (N_12653,N_12553,N_12531);
xor U12654 (N_12654,N_12540,N_12432);
nor U12655 (N_12655,N_12475,N_12434);
nor U12656 (N_12656,N_12530,N_12431);
nor U12657 (N_12657,N_12435,N_12452);
or U12658 (N_12658,N_12447,N_12511);
xnor U12659 (N_12659,N_12537,N_12468);
nor U12660 (N_12660,N_12501,N_12509);
xnor U12661 (N_12661,N_12502,N_12581);
nand U12662 (N_12662,N_12512,N_12476);
nor U12663 (N_12663,N_12472,N_12524);
or U12664 (N_12664,N_12594,N_12493);
and U12665 (N_12665,N_12515,N_12451);
xnor U12666 (N_12666,N_12412,N_12445);
or U12667 (N_12667,N_12463,N_12469);
xnor U12668 (N_12668,N_12402,N_12549);
xor U12669 (N_12669,N_12422,N_12576);
or U12670 (N_12670,N_12496,N_12544);
or U12671 (N_12671,N_12513,N_12589);
and U12672 (N_12672,N_12587,N_12481);
nor U12673 (N_12673,N_12488,N_12437);
nor U12674 (N_12674,N_12504,N_12593);
and U12675 (N_12675,N_12498,N_12489);
nor U12676 (N_12676,N_12578,N_12503);
xor U12677 (N_12677,N_12479,N_12579);
or U12678 (N_12678,N_12486,N_12406);
or U12679 (N_12679,N_12482,N_12449);
or U12680 (N_12680,N_12418,N_12410);
and U12681 (N_12681,N_12564,N_12448);
or U12682 (N_12682,N_12478,N_12558);
xnor U12683 (N_12683,N_12506,N_12516);
nor U12684 (N_12684,N_12571,N_12577);
or U12685 (N_12685,N_12404,N_12566);
nand U12686 (N_12686,N_12495,N_12561);
xor U12687 (N_12687,N_12546,N_12483);
or U12688 (N_12688,N_12519,N_12595);
nor U12689 (N_12689,N_12471,N_12582);
xor U12690 (N_12690,N_12419,N_12580);
nor U12691 (N_12691,N_12425,N_12598);
and U12692 (N_12692,N_12586,N_12428);
nand U12693 (N_12693,N_12423,N_12444);
nand U12694 (N_12694,N_12547,N_12527);
or U12695 (N_12695,N_12470,N_12535);
xor U12696 (N_12696,N_12569,N_12446);
nand U12697 (N_12697,N_12508,N_12510);
and U12698 (N_12698,N_12456,N_12500);
and U12699 (N_12699,N_12518,N_12458);
nor U12700 (N_12700,N_12589,N_12519);
xor U12701 (N_12701,N_12519,N_12432);
xor U12702 (N_12702,N_12598,N_12562);
or U12703 (N_12703,N_12407,N_12408);
or U12704 (N_12704,N_12486,N_12556);
nor U12705 (N_12705,N_12487,N_12563);
nand U12706 (N_12706,N_12511,N_12407);
xnor U12707 (N_12707,N_12420,N_12569);
and U12708 (N_12708,N_12462,N_12533);
and U12709 (N_12709,N_12575,N_12568);
and U12710 (N_12710,N_12511,N_12437);
nor U12711 (N_12711,N_12437,N_12448);
or U12712 (N_12712,N_12523,N_12427);
xor U12713 (N_12713,N_12429,N_12458);
nor U12714 (N_12714,N_12495,N_12590);
and U12715 (N_12715,N_12596,N_12561);
xnor U12716 (N_12716,N_12483,N_12559);
or U12717 (N_12717,N_12401,N_12440);
nor U12718 (N_12718,N_12515,N_12561);
xor U12719 (N_12719,N_12467,N_12495);
xor U12720 (N_12720,N_12492,N_12410);
xnor U12721 (N_12721,N_12422,N_12434);
and U12722 (N_12722,N_12591,N_12437);
nor U12723 (N_12723,N_12477,N_12431);
nor U12724 (N_12724,N_12421,N_12526);
and U12725 (N_12725,N_12404,N_12440);
nor U12726 (N_12726,N_12440,N_12497);
nand U12727 (N_12727,N_12544,N_12477);
nor U12728 (N_12728,N_12500,N_12477);
and U12729 (N_12729,N_12573,N_12453);
and U12730 (N_12730,N_12422,N_12585);
and U12731 (N_12731,N_12482,N_12433);
or U12732 (N_12732,N_12577,N_12460);
nand U12733 (N_12733,N_12574,N_12401);
or U12734 (N_12734,N_12570,N_12538);
or U12735 (N_12735,N_12455,N_12459);
and U12736 (N_12736,N_12584,N_12408);
and U12737 (N_12737,N_12515,N_12436);
and U12738 (N_12738,N_12548,N_12531);
nor U12739 (N_12739,N_12566,N_12473);
nor U12740 (N_12740,N_12535,N_12402);
xor U12741 (N_12741,N_12565,N_12422);
or U12742 (N_12742,N_12409,N_12519);
or U12743 (N_12743,N_12454,N_12583);
nand U12744 (N_12744,N_12529,N_12568);
nor U12745 (N_12745,N_12541,N_12482);
xor U12746 (N_12746,N_12519,N_12407);
or U12747 (N_12747,N_12456,N_12471);
nor U12748 (N_12748,N_12400,N_12509);
nand U12749 (N_12749,N_12512,N_12514);
xnor U12750 (N_12750,N_12456,N_12484);
nand U12751 (N_12751,N_12566,N_12453);
nor U12752 (N_12752,N_12456,N_12514);
nor U12753 (N_12753,N_12512,N_12402);
xor U12754 (N_12754,N_12529,N_12511);
or U12755 (N_12755,N_12574,N_12561);
nor U12756 (N_12756,N_12446,N_12445);
nand U12757 (N_12757,N_12456,N_12452);
nand U12758 (N_12758,N_12481,N_12413);
and U12759 (N_12759,N_12423,N_12506);
nor U12760 (N_12760,N_12529,N_12414);
nand U12761 (N_12761,N_12413,N_12459);
or U12762 (N_12762,N_12587,N_12509);
xor U12763 (N_12763,N_12509,N_12599);
and U12764 (N_12764,N_12471,N_12439);
nor U12765 (N_12765,N_12440,N_12585);
or U12766 (N_12766,N_12540,N_12528);
xor U12767 (N_12767,N_12419,N_12510);
xnor U12768 (N_12768,N_12545,N_12538);
nor U12769 (N_12769,N_12438,N_12545);
nor U12770 (N_12770,N_12455,N_12512);
and U12771 (N_12771,N_12551,N_12414);
or U12772 (N_12772,N_12488,N_12426);
and U12773 (N_12773,N_12503,N_12580);
or U12774 (N_12774,N_12460,N_12540);
nor U12775 (N_12775,N_12402,N_12526);
or U12776 (N_12776,N_12547,N_12439);
and U12777 (N_12777,N_12402,N_12450);
nor U12778 (N_12778,N_12408,N_12450);
or U12779 (N_12779,N_12570,N_12419);
and U12780 (N_12780,N_12486,N_12580);
and U12781 (N_12781,N_12581,N_12404);
and U12782 (N_12782,N_12455,N_12598);
nand U12783 (N_12783,N_12400,N_12478);
nor U12784 (N_12784,N_12530,N_12453);
nor U12785 (N_12785,N_12455,N_12414);
or U12786 (N_12786,N_12509,N_12551);
or U12787 (N_12787,N_12479,N_12464);
or U12788 (N_12788,N_12494,N_12542);
and U12789 (N_12789,N_12539,N_12513);
or U12790 (N_12790,N_12502,N_12445);
nand U12791 (N_12791,N_12509,N_12558);
and U12792 (N_12792,N_12532,N_12565);
nor U12793 (N_12793,N_12507,N_12422);
nor U12794 (N_12794,N_12565,N_12415);
nand U12795 (N_12795,N_12569,N_12429);
nor U12796 (N_12796,N_12467,N_12426);
xnor U12797 (N_12797,N_12582,N_12518);
and U12798 (N_12798,N_12415,N_12506);
nor U12799 (N_12799,N_12566,N_12541);
or U12800 (N_12800,N_12766,N_12733);
or U12801 (N_12801,N_12625,N_12608);
nor U12802 (N_12802,N_12749,N_12639);
nor U12803 (N_12803,N_12774,N_12666);
and U12804 (N_12804,N_12669,N_12640);
xnor U12805 (N_12805,N_12650,N_12752);
nor U12806 (N_12806,N_12792,N_12701);
xnor U12807 (N_12807,N_12641,N_12755);
nor U12808 (N_12808,N_12611,N_12620);
and U12809 (N_12809,N_12748,N_12692);
and U12810 (N_12810,N_12722,N_12797);
or U12811 (N_12811,N_12730,N_12778);
xnor U12812 (N_12812,N_12783,N_12760);
and U12813 (N_12813,N_12699,N_12679);
xor U12814 (N_12814,N_12762,N_12614);
nand U12815 (N_12815,N_12784,N_12646);
nor U12816 (N_12816,N_12768,N_12612);
xnor U12817 (N_12817,N_12659,N_12775);
nand U12818 (N_12818,N_12782,N_12719);
or U12819 (N_12819,N_12616,N_12697);
or U12820 (N_12820,N_12601,N_12770);
or U12821 (N_12821,N_12607,N_12724);
xnor U12822 (N_12822,N_12713,N_12763);
and U12823 (N_12823,N_12729,N_12773);
xor U12824 (N_12824,N_12676,N_12683);
nand U12825 (N_12825,N_12725,N_12765);
or U12826 (N_12826,N_12746,N_12694);
nand U12827 (N_12827,N_12658,N_12734);
nor U12828 (N_12828,N_12745,N_12671);
and U12829 (N_12829,N_12623,N_12624);
nor U12830 (N_12830,N_12772,N_12657);
xnor U12831 (N_12831,N_12781,N_12718);
nor U12832 (N_12832,N_12794,N_12753);
and U12833 (N_12833,N_12708,N_12715);
or U12834 (N_12834,N_12720,N_12700);
nor U12835 (N_12835,N_12710,N_12735);
xor U12836 (N_12836,N_12702,N_12617);
or U12837 (N_12837,N_12675,N_12740);
or U12838 (N_12838,N_12736,N_12648);
xor U12839 (N_12839,N_12788,N_12712);
and U12840 (N_12840,N_12795,N_12677);
and U12841 (N_12841,N_12727,N_12779);
nand U12842 (N_12842,N_12603,N_12731);
nor U12843 (N_12843,N_12610,N_12622);
nor U12844 (N_12844,N_12742,N_12696);
nand U12845 (N_12845,N_12786,N_12796);
nand U12846 (N_12846,N_12703,N_12661);
nand U12847 (N_12847,N_12787,N_12709);
nor U12848 (N_12848,N_12631,N_12618);
xor U12849 (N_12849,N_12728,N_12714);
nand U12850 (N_12850,N_12759,N_12769);
and U12851 (N_12851,N_12600,N_12653);
nor U12852 (N_12852,N_12673,N_12695);
or U12853 (N_12853,N_12758,N_12663);
nand U12854 (N_12854,N_12652,N_12723);
or U12855 (N_12855,N_12739,N_12726);
and U12856 (N_12856,N_12680,N_12785);
nor U12857 (N_12857,N_12721,N_12757);
or U12858 (N_12858,N_12629,N_12602);
and U12859 (N_12859,N_12799,N_12649);
xnor U12860 (N_12860,N_12651,N_12647);
nand U12861 (N_12861,N_12754,N_12798);
nor U12862 (N_12862,N_12642,N_12732);
nor U12863 (N_12863,N_12630,N_12662);
and U12864 (N_12864,N_12665,N_12604);
or U12865 (N_12865,N_12627,N_12678);
xor U12866 (N_12866,N_12756,N_12717);
xor U12867 (N_12867,N_12606,N_12693);
or U12868 (N_12868,N_12668,N_12672);
xnor U12869 (N_12869,N_12705,N_12767);
nand U12870 (N_12870,N_12688,N_12761);
and U12871 (N_12871,N_12689,N_12691);
or U12872 (N_12872,N_12686,N_12764);
xor U12873 (N_12873,N_12777,N_12670);
nor U12874 (N_12874,N_12790,N_12643);
or U12875 (N_12875,N_12789,N_12660);
xnor U12876 (N_12876,N_12637,N_12780);
nand U12877 (N_12877,N_12776,N_12698);
nor U12878 (N_12878,N_12793,N_12706);
nand U12879 (N_12879,N_12635,N_12613);
nor U12880 (N_12880,N_12628,N_12638);
or U12881 (N_12881,N_12687,N_12738);
or U12882 (N_12882,N_12771,N_12791);
nand U12883 (N_12883,N_12645,N_12636);
and U12884 (N_12884,N_12656,N_12681);
xnor U12885 (N_12885,N_12674,N_12632);
and U12886 (N_12886,N_12655,N_12619);
nand U12887 (N_12887,N_12626,N_12621);
xnor U12888 (N_12888,N_12743,N_12737);
or U12889 (N_12889,N_12711,N_12704);
nand U12890 (N_12890,N_12644,N_12707);
and U12891 (N_12891,N_12716,N_12609);
and U12892 (N_12892,N_12605,N_12664);
or U12893 (N_12893,N_12741,N_12654);
or U12894 (N_12894,N_12684,N_12750);
xnor U12895 (N_12895,N_12685,N_12751);
xor U12896 (N_12896,N_12744,N_12615);
nand U12897 (N_12897,N_12747,N_12690);
nand U12898 (N_12898,N_12633,N_12667);
nor U12899 (N_12899,N_12634,N_12682);
xor U12900 (N_12900,N_12701,N_12604);
xor U12901 (N_12901,N_12726,N_12797);
nor U12902 (N_12902,N_12738,N_12647);
xor U12903 (N_12903,N_12721,N_12756);
and U12904 (N_12904,N_12607,N_12608);
xnor U12905 (N_12905,N_12794,N_12781);
and U12906 (N_12906,N_12704,N_12773);
and U12907 (N_12907,N_12760,N_12711);
or U12908 (N_12908,N_12773,N_12619);
and U12909 (N_12909,N_12753,N_12682);
and U12910 (N_12910,N_12756,N_12775);
nand U12911 (N_12911,N_12606,N_12756);
xor U12912 (N_12912,N_12761,N_12747);
nor U12913 (N_12913,N_12635,N_12772);
nor U12914 (N_12914,N_12773,N_12655);
and U12915 (N_12915,N_12789,N_12715);
nor U12916 (N_12916,N_12746,N_12631);
or U12917 (N_12917,N_12752,N_12680);
and U12918 (N_12918,N_12756,N_12750);
or U12919 (N_12919,N_12736,N_12705);
and U12920 (N_12920,N_12767,N_12796);
and U12921 (N_12921,N_12649,N_12662);
nand U12922 (N_12922,N_12751,N_12628);
nor U12923 (N_12923,N_12608,N_12670);
xor U12924 (N_12924,N_12736,N_12671);
and U12925 (N_12925,N_12794,N_12718);
nand U12926 (N_12926,N_12728,N_12795);
nor U12927 (N_12927,N_12669,N_12763);
and U12928 (N_12928,N_12609,N_12798);
xnor U12929 (N_12929,N_12788,N_12678);
xnor U12930 (N_12930,N_12671,N_12693);
xnor U12931 (N_12931,N_12657,N_12771);
xnor U12932 (N_12932,N_12673,N_12660);
or U12933 (N_12933,N_12652,N_12642);
nand U12934 (N_12934,N_12729,N_12704);
nand U12935 (N_12935,N_12769,N_12625);
nor U12936 (N_12936,N_12634,N_12788);
or U12937 (N_12937,N_12735,N_12722);
and U12938 (N_12938,N_12799,N_12628);
xor U12939 (N_12939,N_12773,N_12690);
nand U12940 (N_12940,N_12739,N_12703);
nor U12941 (N_12941,N_12677,N_12793);
or U12942 (N_12942,N_12763,N_12785);
nor U12943 (N_12943,N_12723,N_12693);
nor U12944 (N_12944,N_12664,N_12680);
or U12945 (N_12945,N_12761,N_12695);
nand U12946 (N_12946,N_12667,N_12762);
xor U12947 (N_12947,N_12733,N_12739);
and U12948 (N_12948,N_12776,N_12738);
nor U12949 (N_12949,N_12739,N_12732);
nand U12950 (N_12950,N_12603,N_12707);
nor U12951 (N_12951,N_12709,N_12766);
nor U12952 (N_12952,N_12797,N_12629);
xnor U12953 (N_12953,N_12721,N_12602);
or U12954 (N_12954,N_12710,N_12695);
or U12955 (N_12955,N_12720,N_12623);
or U12956 (N_12956,N_12693,N_12670);
nand U12957 (N_12957,N_12701,N_12769);
and U12958 (N_12958,N_12677,N_12630);
and U12959 (N_12959,N_12624,N_12756);
and U12960 (N_12960,N_12759,N_12689);
or U12961 (N_12961,N_12684,N_12767);
or U12962 (N_12962,N_12639,N_12732);
nand U12963 (N_12963,N_12753,N_12720);
nor U12964 (N_12964,N_12785,N_12622);
and U12965 (N_12965,N_12767,N_12627);
xor U12966 (N_12966,N_12633,N_12747);
nand U12967 (N_12967,N_12759,N_12641);
xnor U12968 (N_12968,N_12795,N_12764);
nand U12969 (N_12969,N_12719,N_12743);
or U12970 (N_12970,N_12676,N_12613);
nor U12971 (N_12971,N_12795,N_12727);
nand U12972 (N_12972,N_12714,N_12742);
nand U12973 (N_12973,N_12623,N_12724);
or U12974 (N_12974,N_12654,N_12789);
xnor U12975 (N_12975,N_12690,N_12667);
nor U12976 (N_12976,N_12666,N_12732);
and U12977 (N_12977,N_12745,N_12699);
nand U12978 (N_12978,N_12662,N_12777);
nand U12979 (N_12979,N_12608,N_12700);
nor U12980 (N_12980,N_12683,N_12631);
nor U12981 (N_12981,N_12708,N_12709);
xor U12982 (N_12982,N_12648,N_12642);
xnor U12983 (N_12983,N_12611,N_12722);
xor U12984 (N_12984,N_12711,N_12644);
and U12985 (N_12985,N_12734,N_12784);
nor U12986 (N_12986,N_12685,N_12632);
and U12987 (N_12987,N_12740,N_12692);
or U12988 (N_12988,N_12780,N_12788);
nand U12989 (N_12989,N_12684,N_12761);
nor U12990 (N_12990,N_12679,N_12609);
or U12991 (N_12991,N_12798,N_12642);
nor U12992 (N_12992,N_12711,N_12751);
nand U12993 (N_12993,N_12734,N_12681);
and U12994 (N_12994,N_12667,N_12796);
and U12995 (N_12995,N_12641,N_12792);
nand U12996 (N_12996,N_12718,N_12612);
or U12997 (N_12997,N_12732,N_12762);
nor U12998 (N_12998,N_12752,N_12750);
xnor U12999 (N_12999,N_12655,N_12786);
nor U13000 (N_13000,N_12838,N_12926);
xnor U13001 (N_13001,N_12930,N_12892);
or U13002 (N_13002,N_12928,N_12921);
or U13003 (N_13003,N_12963,N_12998);
nand U13004 (N_13004,N_12865,N_12956);
xor U13005 (N_13005,N_12933,N_12853);
nor U13006 (N_13006,N_12828,N_12811);
xor U13007 (N_13007,N_12941,N_12942);
or U13008 (N_13008,N_12946,N_12925);
nand U13009 (N_13009,N_12821,N_12902);
nor U13010 (N_13010,N_12891,N_12982);
xnor U13011 (N_13011,N_12958,N_12988);
and U13012 (N_13012,N_12857,N_12992);
nor U13013 (N_13013,N_12849,N_12929);
nand U13014 (N_13014,N_12852,N_12911);
xnor U13015 (N_13015,N_12949,N_12801);
and U13016 (N_13016,N_12945,N_12850);
xnor U13017 (N_13017,N_12806,N_12979);
xor U13018 (N_13018,N_12848,N_12954);
or U13019 (N_13019,N_12965,N_12832);
or U13020 (N_13020,N_12989,N_12904);
xnor U13021 (N_13021,N_12987,N_12914);
xnor U13022 (N_13022,N_12923,N_12996);
nand U13023 (N_13023,N_12844,N_12819);
nor U13024 (N_13024,N_12916,N_12886);
or U13025 (N_13025,N_12815,N_12964);
nor U13026 (N_13026,N_12836,N_12855);
xor U13027 (N_13027,N_12820,N_12972);
xnor U13028 (N_13028,N_12910,N_12858);
nor U13029 (N_13029,N_12968,N_12953);
or U13030 (N_13030,N_12903,N_12974);
nor U13031 (N_13031,N_12837,N_12931);
xor U13032 (N_13032,N_12802,N_12950);
or U13033 (N_13033,N_12981,N_12901);
xor U13034 (N_13034,N_12814,N_12879);
xnor U13035 (N_13035,N_12851,N_12990);
or U13036 (N_13036,N_12969,N_12980);
or U13037 (N_13037,N_12908,N_12876);
nor U13038 (N_13038,N_12948,N_12919);
or U13039 (N_13039,N_12875,N_12835);
and U13040 (N_13040,N_12805,N_12840);
or U13041 (N_13041,N_12888,N_12924);
nor U13042 (N_13042,N_12807,N_12822);
nand U13043 (N_13043,N_12845,N_12962);
xor U13044 (N_13044,N_12859,N_12861);
nor U13045 (N_13045,N_12983,N_12939);
or U13046 (N_13046,N_12842,N_12986);
xnor U13047 (N_13047,N_12947,N_12804);
nor U13048 (N_13048,N_12864,N_12995);
xnor U13049 (N_13049,N_12809,N_12994);
nor U13050 (N_13050,N_12833,N_12882);
xnor U13051 (N_13051,N_12977,N_12863);
nand U13052 (N_13052,N_12831,N_12934);
or U13053 (N_13053,N_12862,N_12913);
nand U13054 (N_13054,N_12889,N_12922);
and U13055 (N_13055,N_12866,N_12967);
or U13056 (N_13056,N_12829,N_12800);
nand U13057 (N_13057,N_12847,N_12884);
or U13058 (N_13058,N_12878,N_12912);
and U13059 (N_13059,N_12810,N_12940);
xnor U13060 (N_13060,N_12854,N_12834);
nor U13061 (N_13061,N_12970,N_12872);
or U13062 (N_13062,N_12915,N_12984);
nor U13063 (N_13063,N_12896,N_12976);
nor U13064 (N_13064,N_12966,N_12997);
and U13065 (N_13065,N_12971,N_12827);
or U13066 (N_13066,N_12943,N_12951);
and U13067 (N_13067,N_12808,N_12909);
xor U13068 (N_13068,N_12871,N_12841);
or U13069 (N_13069,N_12816,N_12920);
or U13070 (N_13070,N_12874,N_12839);
nand U13071 (N_13071,N_12830,N_12868);
or U13072 (N_13072,N_12813,N_12973);
nand U13073 (N_13073,N_12906,N_12927);
and U13074 (N_13074,N_12880,N_12900);
or U13075 (N_13075,N_12917,N_12824);
nand U13076 (N_13076,N_12856,N_12860);
or U13077 (N_13077,N_12817,N_12978);
xnor U13078 (N_13078,N_12826,N_12895);
or U13079 (N_13079,N_12961,N_12823);
and U13080 (N_13080,N_12803,N_12959);
xor U13081 (N_13081,N_12825,N_12905);
or U13082 (N_13082,N_12873,N_12867);
nor U13083 (N_13083,N_12957,N_12818);
and U13084 (N_13084,N_12932,N_12812);
and U13085 (N_13085,N_12991,N_12869);
and U13086 (N_13086,N_12885,N_12897);
nor U13087 (N_13087,N_12877,N_12893);
nand U13088 (N_13088,N_12898,N_12881);
xor U13089 (N_13089,N_12993,N_12935);
xnor U13090 (N_13090,N_12937,N_12936);
and U13091 (N_13091,N_12890,N_12975);
nor U13092 (N_13092,N_12883,N_12985);
or U13093 (N_13093,N_12894,N_12944);
nor U13094 (N_13094,N_12870,N_12899);
and U13095 (N_13095,N_12938,N_12999);
nand U13096 (N_13096,N_12843,N_12952);
nor U13097 (N_13097,N_12918,N_12960);
xnor U13098 (N_13098,N_12846,N_12955);
nor U13099 (N_13099,N_12887,N_12907);
nor U13100 (N_13100,N_12951,N_12851);
xnor U13101 (N_13101,N_12878,N_12980);
nor U13102 (N_13102,N_12800,N_12991);
and U13103 (N_13103,N_12894,N_12890);
nand U13104 (N_13104,N_12895,N_12952);
xnor U13105 (N_13105,N_12917,N_12802);
xnor U13106 (N_13106,N_12847,N_12883);
xor U13107 (N_13107,N_12888,N_12901);
or U13108 (N_13108,N_12898,N_12801);
xnor U13109 (N_13109,N_12958,N_12879);
or U13110 (N_13110,N_12904,N_12853);
or U13111 (N_13111,N_12958,N_12851);
nor U13112 (N_13112,N_12890,N_12835);
xor U13113 (N_13113,N_12932,N_12911);
xor U13114 (N_13114,N_12974,N_12855);
xor U13115 (N_13115,N_12940,N_12824);
and U13116 (N_13116,N_12967,N_12981);
xor U13117 (N_13117,N_12982,N_12819);
and U13118 (N_13118,N_12820,N_12855);
xnor U13119 (N_13119,N_12836,N_12822);
nor U13120 (N_13120,N_12950,N_12921);
and U13121 (N_13121,N_12813,N_12887);
xnor U13122 (N_13122,N_12905,N_12809);
nand U13123 (N_13123,N_12985,N_12810);
nand U13124 (N_13124,N_12823,N_12812);
xnor U13125 (N_13125,N_12880,N_12814);
and U13126 (N_13126,N_12883,N_12975);
nand U13127 (N_13127,N_12921,N_12809);
xnor U13128 (N_13128,N_12808,N_12881);
or U13129 (N_13129,N_12817,N_12825);
nand U13130 (N_13130,N_12828,N_12931);
nor U13131 (N_13131,N_12975,N_12986);
nand U13132 (N_13132,N_12992,N_12856);
nand U13133 (N_13133,N_12899,N_12838);
or U13134 (N_13134,N_12908,N_12988);
nand U13135 (N_13135,N_12952,N_12975);
nor U13136 (N_13136,N_12945,N_12819);
nor U13137 (N_13137,N_12888,N_12846);
and U13138 (N_13138,N_12942,N_12812);
and U13139 (N_13139,N_12869,N_12926);
and U13140 (N_13140,N_12926,N_12892);
nand U13141 (N_13141,N_12841,N_12974);
nand U13142 (N_13142,N_12953,N_12955);
or U13143 (N_13143,N_12921,N_12889);
xnor U13144 (N_13144,N_12812,N_12888);
and U13145 (N_13145,N_12869,N_12988);
and U13146 (N_13146,N_12978,N_12975);
and U13147 (N_13147,N_12923,N_12976);
and U13148 (N_13148,N_12991,N_12932);
and U13149 (N_13149,N_12940,N_12943);
nand U13150 (N_13150,N_12980,N_12853);
nor U13151 (N_13151,N_12940,N_12863);
xor U13152 (N_13152,N_12972,N_12999);
or U13153 (N_13153,N_12906,N_12846);
xnor U13154 (N_13154,N_12890,N_12823);
and U13155 (N_13155,N_12946,N_12969);
or U13156 (N_13156,N_12839,N_12969);
nand U13157 (N_13157,N_12886,N_12801);
nand U13158 (N_13158,N_12965,N_12801);
and U13159 (N_13159,N_12973,N_12868);
nand U13160 (N_13160,N_12816,N_12910);
xnor U13161 (N_13161,N_12876,N_12983);
or U13162 (N_13162,N_12963,N_12886);
nor U13163 (N_13163,N_12903,N_12963);
xnor U13164 (N_13164,N_12846,N_12935);
nor U13165 (N_13165,N_12939,N_12867);
nor U13166 (N_13166,N_12983,N_12862);
nand U13167 (N_13167,N_12826,N_12927);
and U13168 (N_13168,N_12831,N_12953);
xnor U13169 (N_13169,N_12862,N_12869);
or U13170 (N_13170,N_12882,N_12900);
nand U13171 (N_13171,N_12882,N_12811);
nand U13172 (N_13172,N_12818,N_12961);
and U13173 (N_13173,N_12835,N_12837);
nor U13174 (N_13174,N_12869,N_12848);
or U13175 (N_13175,N_12811,N_12852);
and U13176 (N_13176,N_12923,N_12839);
nor U13177 (N_13177,N_12848,N_12901);
and U13178 (N_13178,N_12984,N_12998);
xor U13179 (N_13179,N_12918,N_12991);
and U13180 (N_13180,N_12895,N_12911);
or U13181 (N_13181,N_12853,N_12843);
nand U13182 (N_13182,N_12882,N_12960);
nor U13183 (N_13183,N_12886,N_12934);
nand U13184 (N_13184,N_12866,N_12915);
nor U13185 (N_13185,N_12841,N_12910);
xor U13186 (N_13186,N_12903,N_12916);
nand U13187 (N_13187,N_12968,N_12806);
nor U13188 (N_13188,N_12976,N_12963);
nor U13189 (N_13189,N_12868,N_12889);
and U13190 (N_13190,N_12826,N_12989);
xnor U13191 (N_13191,N_12894,N_12900);
nand U13192 (N_13192,N_12971,N_12908);
and U13193 (N_13193,N_12840,N_12864);
xnor U13194 (N_13194,N_12837,N_12913);
and U13195 (N_13195,N_12901,N_12870);
xor U13196 (N_13196,N_12853,N_12966);
nand U13197 (N_13197,N_12877,N_12869);
and U13198 (N_13198,N_12915,N_12845);
xor U13199 (N_13199,N_12896,N_12853);
nand U13200 (N_13200,N_13080,N_13040);
or U13201 (N_13201,N_13030,N_13055);
nand U13202 (N_13202,N_13120,N_13065);
xnor U13203 (N_13203,N_13028,N_13002);
nand U13204 (N_13204,N_13059,N_13003);
nand U13205 (N_13205,N_13125,N_13052);
xor U13206 (N_13206,N_13182,N_13013);
and U13207 (N_13207,N_13064,N_13095);
and U13208 (N_13208,N_13026,N_13086);
or U13209 (N_13209,N_13142,N_13049);
nor U13210 (N_13210,N_13169,N_13104);
and U13211 (N_13211,N_13093,N_13078);
xor U13212 (N_13212,N_13072,N_13155);
nor U13213 (N_13213,N_13074,N_13138);
and U13214 (N_13214,N_13186,N_13046);
and U13215 (N_13215,N_13196,N_13191);
xnor U13216 (N_13216,N_13134,N_13004);
and U13217 (N_13217,N_13033,N_13185);
xnor U13218 (N_13218,N_13114,N_13041);
and U13219 (N_13219,N_13197,N_13039);
and U13220 (N_13220,N_13009,N_13170);
nand U13221 (N_13221,N_13061,N_13024);
or U13222 (N_13222,N_13171,N_13076);
nand U13223 (N_13223,N_13113,N_13101);
or U13224 (N_13224,N_13147,N_13129);
or U13225 (N_13225,N_13122,N_13157);
and U13226 (N_13226,N_13044,N_13015);
and U13227 (N_13227,N_13192,N_13035);
nor U13228 (N_13228,N_13190,N_13012);
nor U13229 (N_13229,N_13115,N_13133);
nand U13230 (N_13230,N_13089,N_13108);
and U13231 (N_13231,N_13181,N_13016);
nand U13232 (N_13232,N_13067,N_13139);
or U13233 (N_13233,N_13184,N_13118);
xor U13234 (N_13234,N_13137,N_13132);
nor U13235 (N_13235,N_13116,N_13130);
and U13236 (N_13236,N_13032,N_13048);
nor U13237 (N_13237,N_13167,N_13094);
xnor U13238 (N_13238,N_13023,N_13057);
nand U13239 (N_13239,N_13090,N_13031);
or U13240 (N_13240,N_13193,N_13097);
or U13241 (N_13241,N_13121,N_13177);
nand U13242 (N_13242,N_13198,N_13178);
or U13243 (N_13243,N_13005,N_13152);
and U13244 (N_13244,N_13098,N_13084);
and U13245 (N_13245,N_13109,N_13183);
xor U13246 (N_13246,N_13085,N_13143);
or U13247 (N_13247,N_13077,N_13162);
and U13248 (N_13248,N_13001,N_13091);
nand U13249 (N_13249,N_13063,N_13053);
xnor U13250 (N_13250,N_13087,N_13047);
nand U13251 (N_13251,N_13069,N_13168);
and U13252 (N_13252,N_13099,N_13038);
or U13253 (N_13253,N_13022,N_13082);
nor U13254 (N_13254,N_13075,N_13021);
and U13255 (N_13255,N_13158,N_13100);
xnor U13256 (N_13256,N_13079,N_13194);
xor U13257 (N_13257,N_13060,N_13092);
nand U13258 (N_13258,N_13054,N_13160);
nand U13259 (N_13259,N_13037,N_13103);
nor U13260 (N_13260,N_13135,N_13019);
nand U13261 (N_13261,N_13175,N_13163);
nand U13262 (N_13262,N_13111,N_13027);
xor U13263 (N_13263,N_13161,N_13180);
nand U13264 (N_13264,N_13124,N_13051);
nor U13265 (N_13265,N_13106,N_13189);
xnor U13266 (N_13266,N_13020,N_13126);
nor U13267 (N_13267,N_13071,N_13179);
nand U13268 (N_13268,N_13172,N_13066);
nor U13269 (N_13269,N_13173,N_13165);
xnor U13270 (N_13270,N_13148,N_13014);
nor U13271 (N_13271,N_13123,N_13010);
nand U13272 (N_13272,N_13145,N_13011);
nor U13273 (N_13273,N_13107,N_13050);
nand U13274 (N_13274,N_13149,N_13164);
nor U13275 (N_13275,N_13017,N_13029);
xor U13276 (N_13276,N_13110,N_13117);
nand U13277 (N_13277,N_13058,N_13088);
and U13278 (N_13278,N_13007,N_13006);
nand U13279 (N_13279,N_13073,N_13102);
nor U13280 (N_13280,N_13105,N_13018);
and U13281 (N_13281,N_13195,N_13045);
and U13282 (N_13282,N_13070,N_13042);
nand U13283 (N_13283,N_13136,N_13062);
nor U13284 (N_13284,N_13150,N_13154);
nor U13285 (N_13285,N_13151,N_13083);
or U13286 (N_13286,N_13128,N_13166);
xor U13287 (N_13287,N_13188,N_13127);
and U13288 (N_13288,N_13056,N_13140);
nor U13289 (N_13289,N_13146,N_13176);
nor U13290 (N_13290,N_13153,N_13112);
or U13291 (N_13291,N_13141,N_13081);
nor U13292 (N_13292,N_13034,N_13131);
and U13293 (N_13293,N_13144,N_13025);
or U13294 (N_13294,N_13159,N_13043);
or U13295 (N_13295,N_13187,N_13096);
nor U13296 (N_13296,N_13119,N_13008);
nand U13297 (N_13297,N_13156,N_13068);
xnor U13298 (N_13298,N_13036,N_13000);
nand U13299 (N_13299,N_13199,N_13174);
nor U13300 (N_13300,N_13158,N_13167);
xor U13301 (N_13301,N_13156,N_13075);
nand U13302 (N_13302,N_13038,N_13110);
nor U13303 (N_13303,N_13037,N_13026);
nor U13304 (N_13304,N_13103,N_13144);
nand U13305 (N_13305,N_13050,N_13177);
and U13306 (N_13306,N_13050,N_13033);
nor U13307 (N_13307,N_13035,N_13196);
nor U13308 (N_13308,N_13085,N_13037);
nand U13309 (N_13309,N_13022,N_13131);
xor U13310 (N_13310,N_13003,N_13089);
xnor U13311 (N_13311,N_13175,N_13180);
nor U13312 (N_13312,N_13179,N_13117);
xor U13313 (N_13313,N_13081,N_13062);
or U13314 (N_13314,N_13048,N_13073);
or U13315 (N_13315,N_13180,N_13107);
nor U13316 (N_13316,N_13180,N_13144);
nor U13317 (N_13317,N_13011,N_13028);
nor U13318 (N_13318,N_13001,N_13090);
nand U13319 (N_13319,N_13082,N_13164);
nand U13320 (N_13320,N_13143,N_13133);
nor U13321 (N_13321,N_13088,N_13152);
or U13322 (N_13322,N_13095,N_13176);
nor U13323 (N_13323,N_13072,N_13081);
or U13324 (N_13324,N_13009,N_13001);
or U13325 (N_13325,N_13098,N_13178);
nor U13326 (N_13326,N_13125,N_13010);
or U13327 (N_13327,N_13054,N_13052);
nand U13328 (N_13328,N_13118,N_13099);
nor U13329 (N_13329,N_13171,N_13093);
and U13330 (N_13330,N_13188,N_13167);
or U13331 (N_13331,N_13002,N_13081);
or U13332 (N_13332,N_13042,N_13091);
nor U13333 (N_13333,N_13141,N_13020);
or U13334 (N_13334,N_13050,N_13098);
and U13335 (N_13335,N_13103,N_13158);
xor U13336 (N_13336,N_13148,N_13141);
and U13337 (N_13337,N_13034,N_13166);
or U13338 (N_13338,N_13172,N_13090);
nand U13339 (N_13339,N_13159,N_13124);
nor U13340 (N_13340,N_13185,N_13107);
or U13341 (N_13341,N_13155,N_13143);
or U13342 (N_13342,N_13110,N_13040);
or U13343 (N_13343,N_13065,N_13185);
and U13344 (N_13344,N_13057,N_13076);
or U13345 (N_13345,N_13103,N_13114);
xnor U13346 (N_13346,N_13052,N_13161);
nand U13347 (N_13347,N_13104,N_13096);
or U13348 (N_13348,N_13129,N_13059);
or U13349 (N_13349,N_13158,N_13099);
xnor U13350 (N_13350,N_13118,N_13167);
or U13351 (N_13351,N_13125,N_13098);
nor U13352 (N_13352,N_13011,N_13138);
nand U13353 (N_13353,N_13089,N_13167);
nor U13354 (N_13354,N_13085,N_13191);
and U13355 (N_13355,N_13101,N_13068);
nand U13356 (N_13356,N_13013,N_13021);
nor U13357 (N_13357,N_13027,N_13097);
xor U13358 (N_13358,N_13120,N_13156);
or U13359 (N_13359,N_13041,N_13110);
and U13360 (N_13360,N_13029,N_13166);
nor U13361 (N_13361,N_13089,N_13192);
nand U13362 (N_13362,N_13077,N_13157);
nand U13363 (N_13363,N_13158,N_13140);
or U13364 (N_13364,N_13016,N_13021);
xor U13365 (N_13365,N_13089,N_13093);
or U13366 (N_13366,N_13139,N_13159);
or U13367 (N_13367,N_13183,N_13099);
nand U13368 (N_13368,N_13094,N_13150);
nand U13369 (N_13369,N_13179,N_13009);
nor U13370 (N_13370,N_13045,N_13078);
or U13371 (N_13371,N_13016,N_13062);
nand U13372 (N_13372,N_13060,N_13120);
and U13373 (N_13373,N_13033,N_13078);
nand U13374 (N_13374,N_13104,N_13085);
xnor U13375 (N_13375,N_13017,N_13124);
and U13376 (N_13376,N_13102,N_13032);
or U13377 (N_13377,N_13080,N_13008);
xnor U13378 (N_13378,N_13100,N_13133);
xnor U13379 (N_13379,N_13115,N_13127);
or U13380 (N_13380,N_13138,N_13094);
xnor U13381 (N_13381,N_13169,N_13187);
xnor U13382 (N_13382,N_13027,N_13082);
nand U13383 (N_13383,N_13013,N_13193);
or U13384 (N_13384,N_13033,N_13193);
nand U13385 (N_13385,N_13057,N_13125);
and U13386 (N_13386,N_13022,N_13112);
nor U13387 (N_13387,N_13076,N_13177);
nor U13388 (N_13388,N_13194,N_13191);
or U13389 (N_13389,N_13186,N_13164);
xor U13390 (N_13390,N_13110,N_13060);
xnor U13391 (N_13391,N_13094,N_13027);
nor U13392 (N_13392,N_13012,N_13134);
xnor U13393 (N_13393,N_13043,N_13106);
nand U13394 (N_13394,N_13119,N_13198);
xor U13395 (N_13395,N_13163,N_13024);
xnor U13396 (N_13396,N_13012,N_13005);
xnor U13397 (N_13397,N_13069,N_13125);
or U13398 (N_13398,N_13124,N_13187);
nor U13399 (N_13399,N_13175,N_13032);
or U13400 (N_13400,N_13363,N_13304);
and U13401 (N_13401,N_13374,N_13235);
and U13402 (N_13402,N_13330,N_13393);
nor U13403 (N_13403,N_13368,N_13337);
xor U13404 (N_13404,N_13341,N_13358);
nand U13405 (N_13405,N_13208,N_13205);
nand U13406 (N_13406,N_13340,N_13200);
nand U13407 (N_13407,N_13316,N_13280);
xor U13408 (N_13408,N_13252,N_13229);
xnor U13409 (N_13409,N_13317,N_13241);
nand U13410 (N_13410,N_13262,N_13357);
and U13411 (N_13411,N_13321,N_13231);
or U13412 (N_13412,N_13333,N_13238);
or U13413 (N_13413,N_13266,N_13286);
xor U13414 (N_13414,N_13242,N_13339);
and U13415 (N_13415,N_13251,N_13294);
and U13416 (N_13416,N_13350,N_13276);
nand U13417 (N_13417,N_13293,N_13343);
or U13418 (N_13418,N_13388,N_13232);
nand U13419 (N_13419,N_13298,N_13222);
and U13420 (N_13420,N_13297,N_13360);
or U13421 (N_13421,N_13212,N_13320);
and U13422 (N_13422,N_13201,N_13322);
nand U13423 (N_13423,N_13254,N_13285);
nand U13424 (N_13424,N_13275,N_13364);
nand U13425 (N_13425,N_13326,N_13268);
or U13426 (N_13426,N_13290,N_13224);
nand U13427 (N_13427,N_13240,N_13325);
and U13428 (N_13428,N_13203,N_13389);
xor U13429 (N_13429,N_13303,N_13269);
nand U13430 (N_13430,N_13216,N_13292);
and U13431 (N_13431,N_13265,N_13394);
nor U13432 (N_13432,N_13239,N_13291);
and U13433 (N_13433,N_13335,N_13253);
and U13434 (N_13434,N_13261,N_13207);
or U13435 (N_13435,N_13354,N_13277);
nor U13436 (N_13436,N_13271,N_13225);
or U13437 (N_13437,N_13399,N_13259);
nor U13438 (N_13438,N_13305,N_13234);
nor U13439 (N_13439,N_13307,N_13273);
nand U13440 (N_13440,N_13328,N_13384);
or U13441 (N_13441,N_13356,N_13308);
nand U13442 (N_13442,N_13382,N_13383);
or U13443 (N_13443,N_13366,N_13211);
xor U13444 (N_13444,N_13386,N_13352);
or U13445 (N_13445,N_13347,N_13362);
nand U13446 (N_13446,N_13376,N_13295);
nor U13447 (N_13447,N_13323,N_13355);
nand U13448 (N_13448,N_13313,N_13218);
nor U13449 (N_13449,N_13267,N_13215);
nor U13450 (N_13450,N_13209,N_13221);
xor U13451 (N_13451,N_13296,N_13248);
and U13452 (N_13452,N_13338,N_13284);
or U13453 (N_13453,N_13349,N_13217);
nand U13454 (N_13454,N_13237,N_13367);
xor U13455 (N_13455,N_13219,N_13289);
and U13456 (N_13456,N_13391,N_13381);
xnor U13457 (N_13457,N_13282,N_13331);
nand U13458 (N_13458,N_13392,N_13396);
or U13459 (N_13459,N_13233,N_13373);
xnor U13460 (N_13460,N_13310,N_13255);
xor U13461 (N_13461,N_13306,N_13214);
xnor U13462 (N_13462,N_13227,N_13245);
and U13463 (N_13463,N_13365,N_13250);
nor U13464 (N_13464,N_13380,N_13309);
and U13465 (N_13465,N_13345,N_13370);
and U13466 (N_13466,N_13260,N_13371);
nand U13467 (N_13467,N_13287,N_13281);
nor U13468 (N_13468,N_13398,N_13324);
or U13469 (N_13469,N_13206,N_13351);
and U13470 (N_13470,N_13390,N_13379);
nand U13471 (N_13471,N_13270,N_13243);
or U13472 (N_13472,N_13264,N_13378);
nor U13473 (N_13473,N_13369,N_13223);
nand U13474 (N_13474,N_13226,N_13336);
and U13475 (N_13475,N_13332,N_13257);
xnor U13476 (N_13476,N_13315,N_13230);
and U13477 (N_13477,N_13327,N_13213);
and U13478 (N_13478,N_13395,N_13244);
nand U13479 (N_13479,N_13258,N_13348);
and U13480 (N_13480,N_13302,N_13278);
xor U13481 (N_13481,N_13359,N_13283);
nand U13482 (N_13482,N_13314,N_13204);
or U13483 (N_13483,N_13256,N_13279);
and U13484 (N_13484,N_13301,N_13228);
or U13485 (N_13485,N_13334,N_13319);
xor U13486 (N_13486,N_13312,N_13377);
and U13487 (N_13487,N_13300,N_13263);
and U13488 (N_13488,N_13202,N_13353);
nor U13489 (N_13489,N_13274,N_13288);
or U13490 (N_13490,N_13385,N_13249);
nand U13491 (N_13491,N_13236,N_13220);
nand U13492 (N_13492,N_13346,N_13210);
nand U13493 (N_13493,N_13318,N_13387);
nand U13494 (N_13494,N_13246,N_13329);
nor U13495 (N_13495,N_13272,N_13311);
nand U13496 (N_13496,N_13375,N_13247);
or U13497 (N_13497,N_13299,N_13397);
nand U13498 (N_13498,N_13361,N_13342);
xnor U13499 (N_13499,N_13372,N_13344);
nor U13500 (N_13500,N_13287,N_13235);
or U13501 (N_13501,N_13283,N_13248);
nand U13502 (N_13502,N_13213,N_13374);
xor U13503 (N_13503,N_13298,N_13204);
nand U13504 (N_13504,N_13271,N_13335);
and U13505 (N_13505,N_13216,N_13229);
and U13506 (N_13506,N_13274,N_13236);
xor U13507 (N_13507,N_13359,N_13394);
nor U13508 (N_13508,N_13225,N_13324);
xor U13509 (N_13509,N_13257,N_13320);
nor U13510 (N_13510,N_13335,N_13277);
xnor U13511 (N_13511,N_13348,N_13269);
nand U13512 (N_13512,N_13253,N_13383);
xnor U13513 (N_13513,N_13272,N_13324);
nand U13514 (N_13514,N_13341,N_13246);
xnor U13515 (N_13515,N_13217,N_13333);
and U13516 (N_13516,N_13399,N_13375);
xnor U13517 (N_13517,N_13389,N_13364);
and U13518 (N_13518,N_13371,N_13250);
and U13519 (N_13519,N_13285,N_13380);
nand U13520 (N_13520,N_13267,N_13376);
nand U13521 (N_13521,N_13210,N_13203);
or U13522 (N_13522,N_13229,N_13282);
xor U13523 (N_13523,N_13398,N_13376);
nand U13524 (N_13524,N_13202,N_13302);
nand U13525 (N_13525,N_13285,N_13341);
and U13526 (N_13526,N_13304,N_13246);
and U13527 (N_13527,N_13320,N_13230);
nor U13528 (N_13528,N_13308,N_13272);
and U13529 (N_13529,N_13271,N_13266);
nor U13530 (N_13530,N_13203,N_13376);
xnor U13531 (N_13531,N_13385,N_13273);
or U13532 (N_13532,N_13259,N_13220);
or U13533 (N_13533,N_13393,N_13387);
and U13534 (N_13534,N_13200,N_13381);
nand U13535 (N_13535,N_13378,N_13321);
xor U13536 (N_13536,N_13259,N_13215);
and U13537 (N_13537,N_13367,N_13268);
nor U13538 (N_13538,N_13216,N_13319);
nand U13539 (N_13539,N_13309,N_13279);
nand U13540 (N_13540,N_13248,N_13301);
and U13541 (N_13541,N_13361,N_13234);
or U13542 (N_13542,N_13345,N_13258);
nand U13543 (N_13543,N_13316,N_13297);
or U13544 (N_13544,N_13372,N_13308);
and U13545 (N_13545,N_13224,N_13392);
nor U13546 (N_13546,N_13388,N_13360);
and U13547 (N_13547,N_13388,N_13356);
nor U13548 (N_13548,N_13230,N_13269);
and U13549 (N_13549,N_13281,N_13306);
xnor U13550 (N_13550,N_13339,N_13399);
nor U13551 (N_13551,N_13282,N_13221);
or U13552 (N_13552,N_13311,N_13267);
or U13553 (N_13553,N_13324,N_13231);
nand U13554 (N_13554,N_13310,N_13330);
and U13555 (N_13555,N_13297,N_13240);
and U13556 (N_13556,N_13313,N_13320);
and U13557 (N_13557,N_13291,N_13391);
nand U13558 (N_13558,N_13366,N_13308);
or U13559 (N_13559,N_13232,N_13345);
nand U13560 (N_13560,N_13238,N_13384);
xor U13561 (N_13561,N_13260,N_13304);
nor U13562 (N_13562,N_13378,N_13344);
or U13563 (N_13563,N_13250,N_13311);
or U13564 (N_13564,N_13296,N_13240);
xor U13565 (N_13565,N_13350,N_13352);
nand U13566 (N_13566,N_13315,N_13263);
and U13567 (N_13567,N_13235,N_13224);
or U13568 (N_13568,N_13340,N_13250);
nor U13569 (N_13569,N_13215,N_13378);
and U13570 (N_13570,N_13218,N_13210);
or U13571 (N_13571,N_13272,N_13328);
nor U13572 (N_13572,N_13297,N_13356);
or U13573 (N_13573,N_13230,N_13256);
and U13574 (N_13574,N_13385,N_13218);
nor U13575 (N_13575,N_13239,N_13252);
and U13576 (N_13576,N_13267,N_13357);
nand U13577 (N_13577,N_13272,N_13294);
nand U13578 (N_13578,N_13333,N_13241);
and U13579 (N_13579,N_13398,N_13208);
and U13580 (N_13580,N_13261,N_13352);
xnor U13581 (N_13581,N_13248,N_13221);
nor U13582 (N_13582,N_13304,N_13318);
nor U13583 (N_13583,N_13206,N_13377);
and U13584 (N_13584,N_13384,N_13282);
and U13585 (N_13585,N_13291,N_13259);
nor U13586 (N_13586,N_13372,N_13333);
nand U13587 (N_13587,N_13346,N_13211);
nor U13588 (N_13588,N_13207,N_13227);
xnor U13589 (N_13589,N_13300,N_13249);
nand U13590 (N_13590,N_13236,N_13254);
nand U13591 (N_13591,N_13380,N_13367);
nand U13592 (N_13592,N_13329,N_13238);
xor U13593 (N_13593,N_13317,N_13214);
nand U13594 (N_13594,N_13243,N_13297);
nand U13595 (N_13595,N_13226,N_13249);
or U13596 (N_13596,N_13215,N_13270);
and U13597 (N_13597,N_13294,N_13320);
xnor U13598 (N_13598,N_13336,N_13262);
nand U13599 (N_13599,N_13270,N_13242);
xnor U13600 (N_13600,N_13593,N_13565);
or U13601 (N_13601,N_13428,N_13442);
nor U13602 (N_13602,N_13569,N_13458);
nor U13603 (N_13603,N_13500,N_13534);
nor U13604 (N_13604,N_13556,N_13437);
nor U13605 (N_13605,N_13579,N_13444);
and U13606 (N_13606,N_13594,N_13403);
nand U13607 (N_13607,N_13554,N_13468);
nor U13608 (N_13608,N_13485,N_13581);
nor U13609 (N_13609,N_13598,N_13411);
and U13610 (N_13610,N_13409,N_13573);
or U13611 (N_13611,N_13563,N_13432);
or U13612 (N_13612,N_13502,N_13517);
and U13613 (N_13613,N_13491,N_13460);
nor U13614 (N_13614,N_13465,N_13533);
nand U13615 (N_13615,N_13482,N_13404);
nand U13616 (N_13616,N_13507,N_13541);
or U13617 (N_13617,N_13431,N_13481);
and U13618 (N_13618,N_13558,N_13443);
xnor U13619 (N_13619,N_13483,N_13514);
and U13620 (N_13620,N_13503,N_13511);
or U13621 (N_13621,N_13542,N_13414);
xnor U13622 (N_13622,N_13597,N_13523);
or U13623 (N_13623,N_13497,N_13464);
xor U13624 (N_13624,N_13400,N_13474);
xnor U13625 (N_13625,N_13509,N_13548);
or U13626 (N_13626,N_13498,N_13518);
nand U13627 (N_13627,N_13596,N_13552);
or U13628 (N_13628,N_13478,N_13504);
or U13629 (N_13629,N_13557,N_13567);
or U13630 (N_13630,N_13587,N_13592);
and U13631 (N_13631,N_13476,N_13425);
xor U13632 (N_13632,N_13440,N_13433);
and U13633 (N_13633,N_13574,N_13520);
and U13634 (N_13634,N_13493,N_13577);
or U13635 (N_13635,N_13501,N_13412);
or U13636 (N_13636,N_13549,N_13510);
nor U13637 (N_13637,N_13560,N_13599);
or U13638 (N_13638,N_13457,N_13405);
nor U13639 (N_13639,N_13551,N_13401);
nand U13640 (N_13640,N_13423,N_13408);
nand U13641 (N_13641,N_13480,N_13462);
xor U13642 (N_13642,N_13516,N_13453);
and U13643 (N_13643,N_13540,N_13562);
nand U13644 (N_13644,N_13568,N_13459);
nor U13645 (N_13645,N_13529,N_13492);
nand U13646 (N_13646,N_13447,N_13434);
and U13647 (N_13647,N_13530,N_13463);
or U13648 (N_13648,N_13449,N_13439);
and U13649 (N_13649,N_13450,N_13477);
xnor U13650 (N_13650,N_13436,N_13546);
or U13651 (N_13651,N_13410,N_13572);
or U13652 (N_13652,N_13564,N_13531);
and U13653 (N_13653,N_13580,N_13583);
nor U13654 (N_13654,N_13589,N_13575);
xnor U13655 (N_13655,N_13513,N_13470);
and U13656 (N_13656,N_13535,N_13435);
and U13657 (N_13657,N_13471,N_13488);
xnor U13658 (N_13658,N_13545,N_13595);
xor U13659 (N_13659,N_13469,N_13406);
nand U13660 (N_13660,N_13489,N_13475);
nor U13661 (N_13661,N_13527,N_13588);
and U13662 (N_13662,N_13578,N_13416);
nand U13663 (N_13663,N_13495,N_13487);
and U13664 (N_13664,N_13537,N_13415);
or U13665 (N_13665,N_13559,N_13521);
nor U13666 (N_13666,N_13582,N_13484);
xnor U13667 (N_13667,N_13566,N_13499);
nand U13668 (N_13668,N_13438,N_13550);
nand U13669 (N_13669,N_13528,N_13570);
xor U13670 (N_13670,N_13422,N_13424);
and U13671 (N_13671,N_13418,N_13506);
nand U13672 (N_13672,N_13585,N_13525);
xor U13673 (N_13673,N_13539,N_13584);
and U13674 (N_13674,N_13486,N_13413);
xor U13675 (N_13675,N_13448,N_13456);
or U13676 (N_13676,N_13446,N_13590);
nand U13677 (N_13677,N_13441,N_13466);
nand U13678 (N_13678,N_13591,N_13420);
nand U13679 (N_13679,N_13536,N_13494);
xor U13680 (N_13680,N_13429,N_13454);
and U13681 (N_13681,N_13402,N_13544);
nand U13682 (N_13682,N_13553,N_13417);
nand U13683 (N_13683,N_13445,N_13519);
nand U13684 (N_13684,N_13407,N_13524);
and U13685 (N_13685,N_13561,N_13455);
xnor U13686 (N_13686,N_13473,N_13461);
and U13687 (N_13687,N_13526,N_13452);
xnor U13688 (N_13688,N_13451,N_13576);
or U13689 (N_13689,N_13543,N_13571);
and U13690 (N_13690,N_13547,N_13427);
and U13691 (N_13691,N_13490,N_13505);
xnor U13692 (N_13692,N_13472,N_13522);
nor U13693 (N_13693,N_13430,N_13515);
nor U13694 (N_13694,N_13496,N_13426);
nand U13695 (N_13695,N_13538,N_13467);
and U13696 (N_13696,N_13508,N_13512);
xnor U13697 (N_13697,N_13555,N_13419);
nand U13698 (N_13698,N_13586,N_13421);
nor U13699 (N_13699,N_13479,N_13532);
and U13700 (N_13700,N_13552,N_13544);
nor U13701 (N_13701,N_13430,N_13429);
nor U13702 (N_13702,N_13583,N_13451);
nand U13703 (N_13703,N_13462,N_13530);
nor U13704 (N_13704,N_13543,N_13550);
and U13705 (N_13705,N_13445,N_13488);
and U13706 (N_13706,N_13516,N_13496);
xor U13707 (N_13707,N_13589,N_13509);
or U13708 (N_13708,N_13562,N_13470);
nor U13709 (N_13709,N_13442,N_13538);
xnor U13710 (N_13710,N_13463,N_13508);
nor U13711 (N_13711,N_13510,N_13589);
nand U13712 (N_13712,N_13461,N_13597);
or U13713 (N_13713,N_13455,N_13586);
xor U13714 (N_13714,N_13413,N_13502);
xnor U13715 (N_13715,N_13555,N_13564);
nand U13716 (N_13716,N_13496,N_13440);
xnor U13717 (N_13717,N_13506,N_13488);
and U13718 (N_13718,N_13552,N_13426);
nand U13719 (N_13719,N_13568,N_13503);
and U13720 (N_13720,N_13443,N_13564);
xnor U13721 (N_13721,N_13421,N_13556);
xnor U13722 (N_13722,N_13405,N_13428);
or U13723 (N_13723,N_13543,N_13493);
xnor U13724 (N_13724,N_13438,N_13599);
nand U13725 (N_13725,N_13415,N_13420);
nor U13726 (N_13726,N_13465,N_13594);
or U13727 (N_13727,N_13514,N_13430);
xor U13728 (N_13728,N_13407,N_13430);
or U13729 (N_13729,N_13421,N_13485);
nand U13730 (N_13730,N_13471,N_13406);
and U13731 (N_13731,N_13429,N_13584);
nor U13732 (N_13732,N_13468,N_13458);
xnor U13733 (N_13733,N_13493,N_13538);
and U13734 (N_13734,N_13419,N_13514);
nor U13735 (N_13735,N_13532,N_13517);
xnor U13736 (N_13736,N_13471,N_13517);
nand U13737 (N_13737,N_13488,N_13501);
and U13738 (N_13738,N_13480,N_13586);
xnor U13739 (N_13739,N_13470,N_13565);
nor U13740 (N_13740,N_13451,N_13515);
nand U13741 (N_13741,N_13484,N_13437);
nand U13742 (N_13742,N_13544,N_13442);
or U13743 (N_13743,N_13404,N_13420);
nand U13744 (N_13744,N_13434,N_13559);
nor U13745 (N_13745,N_13465,N_13516);
and U13746 (N_13746,N_13473,N_13415);
and U13747 (N_13747,N_13480,N_13584);
or U13748 (N_13748,N_13583,N_13424);
or U13749 (N_13749,N_13574,N_13463);
nand U13750 (N_13750,N_13464,N_13434);
nand U13751 (N_13751,N_13465,N_13592);
nand U13752 (N_13752,N_13596,N_13592);
nor U13753 (N_13753,N_13509,N_13492);
nand U13754 (N_13754,N_13504,N_13529);
xnor U13755 (N_13755,N_13405,N_13592);
xnor U13756 (N_13756,N_13440,N_13478);
xnor U13757 (N_13757,N_13476,N_13496);
xor U13758 (N_13758,N_13520,N_13522);
xnor U13759 (N_13759,N_13555,N_13471);
nor U13760 (N_13760,N_13497,N_13435);
xnor U13761 (N_13761,N_13542,N_13438);
or U13762 (N_13762,N_13595,N_13429);
or U13763 (N_13763,N_13450,N_13474);
xnor U13764 (N_13764,N_13563,N_13426);
or U13765 (N_13765,N_13424,N_13463);
nand U13766 (N_13766,N_13424,N_13494);
and U13767 (N_13767,N_13455,N_13577);
and U13768 (N_13768,N_13431,N_13474);
and U13769 (N_13769,N_13449,N_13467);
or U13770 (N_13770,N_13551,N_13523);
xnor U13771 (N_13771,N_13520,N_13498);
and U13772 (N_13772,N_13443,N_13471);
or U13773 (N_13773,N_13409,N_13411);
xnor U13774 (N_13774,N_13461,N_13586);
nor U13775 (N_13775,N_13415,N_13445);
nor U13776 (N_13776,N_13524,N_13512);
nor U13777 (N_13777,N_13431,N_13521);
and U13778 (N_13778,N_13523,N_13561);
and U13779 (N_13779,N_13441,N_13425);
and U13780 (N_13780,N_13409,N_13519);
nand U13781 (N_13781,N_13432,N_13508);
nand U13782 (N_13782,N_13593,N_13490);
nor U13783 (N_13783,N_13556,N_13483);
xor U13784 (N_13784,N_13593,N_13411);
nand U13785 (N_13785,N_13437,N_13442);
nor U13786 (N_13786,N_13445,N_13521);
or U13787 (N_13787,N_13541,N_13448);
nor U13788 (N_13788,N_13433,N_13449);
nand U13789 (N_13789,N_13482,N_13485);
nor U13790 (N_13790,N_13560,N_13558);
nand U13791 (N_13791,N_13536,N_13510);
and U13792 (N_13792,N_13588,N_13539);
nand U13793 (N_13793,N_13417,N_13504);
or U13794 (N_13794,N_13483,N_13423);
xor U13795 (N_13795,N_13420,N_13443);
xor U13796 (N_13796,N_13453,N_13473);
nor U13797 (N_13797,N_13517,N_13432);
or U13798 (N_13798,N_13537,N_13440);
xor U13799 (N_13799,N_13483,N_13447);
nand U13800 (N_13800,N_13698,N_13788);
xor U13801 (N_13801,N_13646,N_13773);
nand U13802 (N_13802,N_13716,N_13743);
or U13803 (N_13803,N_13730,N_13668);
and U13804 (N_13804,N_13778,N_13651);
nand U13805 (N_13805,N_13750,N_13798);
xnor U13806 (N_13806,N_13794,N_13747);
and U13807 (N_13807,N_13634,N_13739);
and U13808 (N_13808,N_13767,N_13649);
xnor U13809 (N_13809,N_13728,N_13702);
nand U13810 (N_13810,N_13602,N_13642);
nand U13811 (N_13811,N_13627,N_13638);
nand U13812 (N_13812,N_13618,N_13608);
or U13813 (N_13813,N_13701,N_13640);
or U13814 (N_13814,N_13697,N_13683);
nand U13815 (N_13815,N_13601,N_13658);
nand U13816 (N_13816,N_13790,N_13774);
nor U13817 (N_13817,N_13754,N_13738);
nand U13818 (N_13818,N_13636,N_13763);
nand U13819 (N_13819,N_13660,N_13674);
and U13820 (N_13820,N_13734,N_13741);
xor U13821 (N_13821,N_13619,N_13665);
and U13822 (N_13822,N_13735,N_13779);
nand U13823 (N_13823,N_13706,N_13623);
nor U13824 (N_13824,N_13709,N_13755);
nand U13825 (N_13825,N_13748,N_13784);
nand U13826 (N_13826,N_13662,N_13717);
nand U13827 (N_13827,N_13729,N_13704);
nor U13828 (N_13828,N_13617,N_13737);
xor U13829 (N_13829,N_13605,N_13791);
and U13830 (N_13830,N_13652,N_13705);
nand U13831 (N_13831,N_13687,N_13757);
xnor U13832 (N_13832,N_13693,N_13609);
nor U13833 (N_13833,N_13615,N_13688);
nor U13834 (N_13834,N_13639,N_13770);
nor U13835 (N_13835,N_13696,N_13726);
or U13836 (N_13836,N_13679,N_13742);
nand U13837 (N_13837,N_13795,N_13644);
and U13838 (N_13838,N_13699,N_13607);
nor U13839 (N_13839,N_13733,N_13732);
nor U13840 (N_13840,N_13657,N_13682);
or U13841 (N_13841,N_13710,N_13677);
nor U13842 (N_13842,N_13764,N_13744);
nor U13843 (N_13843,N_13797,N_13678);
and U13844 (N_13844,N_13719,N_13690);
xor U13845 (N_13845,N_13695,N_13723);
or U13846 (N_13846,N_13789,N_13633);
or U13847 (N_13847,N_13659,N_13783);
or U13848 (N_13848,N_13653,N_13648);
nand U13849 (N_13849,N_13606,N_13661);
xnor U13850 (N_13850,N_13758,N_13720);
nand U13851 (N_13851,N_13759,N_13727);
nor U13852 (N_13852,N_13655,N_13670);
or U13853 (N_13853,N_13746,N_13721);
nand U13854 (N_13854,N_13613,N_13664);
nor U13855 (N_13855,N_13685,N_13708);
nand U13856 (N_13856,N_13793,N_13624);
nor U13857 (N_13857,N_13756,N_13780);
nor U13858 (N_13858,N_13629,N_13614);
xor U13859 (N_13859,N_13771,N_13632);
xnor U13860 (N_13860,N_13772,N_13666);
nand U13861 (N_13861,N_13603,N_13680);
or U13862 (N_13862,N_13777,N_13761);
xor U13863 (N_13863,N_13782,N_13715);
nor U13864 (N_13864,N_13672,N_13625);
nor U13865 (N_13865,N_13760,N_13616);
or U13866 (N_13866,N_13786,N_13753);
and U13867 (N_13867,N_13676,N_13673);
nor U13868 (N_13868,N_13612,N_13630);
and U13869 (N_13869,N_13671,N_13643);
or U13870 (N_13870,N_13703,N_13628);
nor U13871 (N_13871,N_13654,N_13637);
xor U13872 (N_13872,N_13740,N_13684);
nor U13873 (N_13873,N_13745,N_13787);
and U13874 (N_13874,N_13762,N_13796);
nand U13875 (N_13875,N_13611,N_13641);
or U13876 (N_13876,N_13781,N_13718);
or U13877 (N_13877,N_13631,N_13656);
nand U13878 (N_13878,N_13621,N_13751);
xnor U13879 (N_13879,N_13620,N_13711);
and U13880 (N_13880,N_13667,N_13722);
or U13881 (N_13881,N_13635,N_13785);
and U13882 (N_13882,N_13600,N_13736);
and U13883 (N_13883,N_13766,N_13604);
nor U13884 (N_13884,N_13776,N_13681);
xor U13885 (N_13885,N_13663,N_13692);
or U13886 (N_13886,N_13650,N_13645);
or U13887 (N_13887,N_13765,N_13731);
nand U13888 (N_13888,N_13775,N_13769);
xor U13889 (N_13889,N_13622,N_13725);
or U13890 (N_13890,N_13669,N_13752);
xnor U13891 (N_13891,N_13647,N_13749);
nand U13892 (N_13892,N_13707,N_13694);
nor U13893 (N_13893,N_13689,N_13610);
xnor U13894 (N_13894,N_13626,N_13712);
and U13895 (N_13895,N_13724,N_13713);
nand U13896 (N_13896,N_13768,N_13799);
and U13897 (N_13897,N_13686,N_13700);
xor U13898 (N_13898,N_13792,N_13675);
xor U13899 (N_13899,N_13714,N_13691);
xor U13900 (N_13900,N_13767,N_13659);
nand U13901 (N_13901,N_13606,N_13704);
nor U13902 (N_13902,N_13705,N_13738);
or U13903 (N_13903,N_13667,N_13695);
xnor U13904 (N_13904,N_13756,N_13661);
xnor U13905 (N_13905,N_13738,N_13752);
nor U13906 (N_13906,N_13738,N_13664);
and U13907 (N_13907,N_13650,N_13797);
and U13908 (N_13908,N_13670,N_13749);
nand U13909 (N_13909,N_13647,N_13743);
or U13910 (N_13910,N_13770,N_13686);
xor U13911 (N_13911,N_13652,N_13661);
or U13912 (N_13912,N_13739,N_13716);
and U13913 (N_13913,N_13602,N_13623);
xor U13914 (N_13914,N_13605,N_13627);
xor U13915 (N_13915,N_13634,N_13690);
xnor U13916 (N_13916,N_13791,N_13788);
or U13917 (N_13917,N_13671,N_13774);
nand U13918 (N_13918,N_13658,N_13606);
nand U13919 (N_13919,N_13790,N_13650);
xor U13920 (N_13920,N_13654,N_13604);
or U13921 (N_13921,N_13721,N_13754);
xor U13922 (N_13922,N_13763,N_13771);
nand U13923 (N_13923,N_13611,N_13658);
xnor U13924 (N_13924,N_13774,N_13792);
and U13925 (N_13925,N_13668,N_13707);
or U13926 (N_13926,N_13707,N_13638);
xor U13927 (N_13927,N_13679,N_13750);
xnor U13928 (N_13928,N_13626,N_13795);
and U13929 (N_13929,N_13685,N_13750);
nor U13930 (N_13930,N_13796,N_13798);
nor U13931 (N_13931,N_13716,N_13692);
xor U13932 (N_13932,N_13758,N_13786);
nand U13933 (N_13933,N_13785,N_13611);
xnor U13934 (N_13934,N_13752,N_13721);
xnor U13935 (N_13935,N_13743,N_13728);
nand U13936 (N_13936,N_13775,N_13622);
and U13937 (N_13937,N_13761,N_13780);
nor U13938 (N_13938,N_13797,N_13789);
nor U13939 (N_13939,N_13652,N_13628);
xor U13940 (N_13940,N_13773,N_13671);
or U13941 (N_13941,N_13626,N_13781);
nand U13942 (N_13942,N_13718,N_13655);
nor U13943 (N_13943,N_13686,N_13607);
or U13944 (N_13944,N_13722,N_13641);
nand U13945 (N_13945,N_13638,N_13687);
or U13946 (N_13946,N_13723,N_13779);
xnor U13947 (N_13947,N_13735,N_13642);
xor U13948 (N_13948,N_13738,N_13770);
xnor U13949 (N_13949,N_13680,N_13656);
or U13950 (N_13950,N_13713,N_13696);
xnor U13951 (N_13951,N_13661,N_13629);
xor U13952 (N_13952,N_13758,N_13646);
nand U13953 (N_13953,N_13708,N_13707);
nor U13954 (N_13954,N_13774,N_13631);
and U13955 (N_13955,N_13685,N_13602);
or U13956 (N_13956,N_13799,N_13660);
nor U13957 (N_13957,N_13646,N_13717);
xnor U13958 (N_13958,N_13738,N_13776);
nand U13959 (N_13959,N_13706,N_13617);
or U13960 (N_13960,N_13745,N_13682);
nor U13961 (N_13961,N_13757,N_13603);
xnor U13962 (N_13962,N_13756,N_13772);
and U13963 (N_13963,N_13616,N_13627);
nand U13964 (N_13964,N_13681,N_13704);
and U13965 (N_13965,N_13767,N_13729);
nor U13966 (N_13966,N_13649,N_13708);
nor U13967 (N_13967,N_13658,N_13663);
and U13968 (N_13968,N_13725,N_13655);
and U13969 (N_13969,N_13637,N_13709);
nand U13970 (N_13970,N_13723,N_13691);
and U13971 (N_13971,N_13692,N_13751);
nand U13972 (N_13972,N_13743,N_13796);
or U13973 (N_13973,N_13666,N_13667);
nand U13974 (N_13974,N_13777,N_13757);
nor U13975 (N_13975,N_13737,N_13652);
xnor U13976 (N_13976,N_13710,N_13739);
nor U13977 (N_13977,N_13780,N_13646);
nor U13978 (N_13978,N_13634,N_13781);
nor U13979 (N_13979,N_13652,N_13693);
and U13980 (N_13980,N_13758,N_13670);
xnor U13981 (N_13981,N_13691,N_13705);
and U13982 (N_13982,N_13616,N_13751);
xor U13983 (N_13983,N_13776,N_13717);
and U13984 (N_13984,N_13751,N_13640);
and U13985 (N_13985,N_13619,N_13608);
xor U13986 (N_13986,N_13789,N_13717);
or U13987 (N_13987,N_13697,N_13735);
nor U13988 (N_13988,N_13671,N_13776);
or U13989 (N_13989,N_13639,N_13686);
and U13990 (N_13990,N_13769,N_13620);
nand U13991 (N_13991,N_13705,N_13669);
and U13992 (N_13992,N_13685,N_13660);
nand U13993 (N_13993,N_13611,N_13612);
nor U13994 (N_13994,N_13695,N_13771);
nand U13995 (N_13995,N_13743,N_13673);
or U13996 (N_13996,N_13641,N_13657);
xnor U13997 (N_13997,N_13775,N_13709);
nor U13998 (N_13998,N_13763,N_13754);
nor U13999 (N_13999,N_13684,N_13778);
nor U14000 (N_14000,N_13802,N_13931);
nor U14001 (N_14001,N_13973,N_13801);
or U14002 (N_14002,N_13882,N_13969);
xnor U14003 (N_14003,N_13938,N_13976);
xnor U14004 (N_14004,N_13897,N_13998);
or U14005 (N_14005,N_13831,N_13849);
or U14006 (N_14006,N_13966,N_13820);
nor U14007 (N_14007,N_13985,N_13928);
and U14008 (N_14008,N_13906,N_13933);
nand U14009 (N_14009,N_13816,N_13834);
nand U14010 (N_14010,N_13884,N_13946);
nand U14011 (N_14011,N_13919,N_13952);
nor U14012 (N_14012,N_13999,N_13807);
and U14013 (N_14013,N_13850,N_13949);
or U14014 (N_14014,N_13824,N_13874);
nor U14015 (N_14015,N_13865,N_13803);
xnor U14016 (N_14016,N_13868,N_13947);
xnor U14017 (N_14017,N_13830,N_13904);
nor U14018 (N_14018,N_13920,N_13908);
nand U14019 (N_14019,N_13854,N_13987);
and U14020 (N_14020,N_13826,N_13875);
and U14021 (N_14021,N_13932,N_13996);
xnor U14022 (N_14022,N_13907,N_13980);
xor U14023 (N_14023,N_13846,N_13909);
nand U14024 (N_14024,N_13841,N_13956);
and U14025 (N_14025,N_13978,N_13936);
xor U14026 (N_14026,N_13898,N_13859);
nand U14027 (N_14027,N_13892,N_13876);
nor U14028 (N_14028,N_13886,N_13871);
and U14029 (N_14029,N_13900,N_13883);
xnor U14030 (N_14030,N_13974,N_13829);
nand U14031 (N_14031,N_13893,N_13986);
nand U14032 (N_14032,N_13843,N_13948);
or U14033 (N_14033,N_13852,N_13923);
or U14034 (N_14034,N_13839,N_13962);
nor U14035 (N_14035,N_13961,N_13945);
nor U14036 (N_14036,N_13845,N_13842);
nand U14037 (N_14037,N_13917,N_13942);
or U14038 (N_14038,N_13914,N_13862);
and U14039 (N_14039,N_13915,N_13922);
nor U14040 (N_14040,N_13885,N_13995);
nand U14041 (N_14041,N_13815,N_13983);
nor U14042 (N_14042,N_13913,N_13958);
xor U14043 (N_14043,N_13997,N_13954);
nor U14044 (N_14044,N_13895,N_13870);
nor U14045 (N_14045,N_13814,N_13927);
and U14046 (N_14046,N_13937,N_13869);
nand U14047 (N_14047,N_13805,N_13889);
or U14048 (N_14048,N_13877,N_13992);
xnor U14049 (N_14049,N_13990,N_13890);
xor U14050 (N_14050,N_13848,N_13896);
xnor U14051 (N_14051,N_13988,N_13951);
nand U14052 (N_14052,N_13899,N_13856);
xor U14053 (N_14053,N_13838,N_13918);
nor U14054 (N_14054,N_13991,N_13836);
nor U14055 (N_14055,N_13943,N_13925);
and U14056 (N_14056,N_13894,N_13964);
xor U14057 (N_14057,N_13860,N_13910);
nor U14058 (N_14058,N_13866,N_13800);
or U14059 (N_14059,N_13994,N_13953);
nand U14060 (N_14060,N_13823,N_13955);
xor U14061 (N_14061,N_13858,N_13929);
nor U14062 (N_14062,N_13891,N_13873);
nor U14063 (N_14063,N_13828,N_13982);
or U14064 (N_14064,N_13903,N_13959);
nor U14065 (N_14065,N_13905,N_13861);
and U14066 (N_14066,N_13960,N_13911);
xor U14067 (N_14067,N_13993,N_13963);
nand U14068 (N_14068,N_13939,N_13981);
or U14069 (N_14069,N_13880,N_13804);
or U14070 (N_14070,N_13818,N_13902);
nand U14071 (N_14071,N_13810,N_13821);
nand U14072 (N_14072,N_13835,N_13965);
nor U14073 (N_14073,N_13881,N_13822);
nand U14074 (N_14074,N_13901,N_13935);
xor U14075 (N_14075,N_13832,N_13817);
nor U14076 (N_14076,N_13872,N_13809);
nand U14077 (N_14077,N_13968,N_13851);
nor U14078 (N_14078,N_13888,N_13979);
or U14079 (N_14079,N_13853,N_13819);
or U14080 (N_14080,N_13879,N_13855);
xnor U14081 (N_14081,N_13921,N_13808);
xnor U14082 (N_14082,N_13957,N_13867);
nand U14083 (N_14083,N_13813,N_13827);
and U14084 (N_14084,N_13989,N_13916);
nand U14085 (N_14085,N_13971,N_13972);
and U14086 (N_14086,N_13837,N_13825);
or U14087 (N_14087,N_13844,N_13811);
nor U14088 (N_14088,N_13812,N_13941);
nor U14089 (N_14089,N_13857,N_13984);
nor U14090 (N_14090,N_13944,N_13975);
or U14091 (N_14091,N_13878,N_13950);
and U14092 (N_14092,N_13887,N_13863);
or U14093 (N_14093,N_13926,N_13864);
nand U14094 (N_14094,N_13806,N_13970);
nand U14095 (N_14095,N_13977,N_13967);
nand U14096 (N_14096,N_13930,N_13924);
xor U14097 (N_14097,N_13940,N_13833);
and U14098 (N_14098,N_13840,N_13847);
nand U14099 (N_14099,N_13934,N_13912);
nand U14100 (N_14100,N_13900,N_13952);
nand U14101 (N_14101,N_13862,N_13875);
nor U14102 (N_14102,N_13954,N_13902);
and U14103 (N_14103,N_13891,N_13954);
nor U14104 (N_14104,N_13917,N_13843);
nand U14105 (N_14105,N_13849,N_13993);
nor U14106 (N_14106,N_13839,N_13912);
or U14107 (N_14107,N_13839,N_13996);
and U14108 (N_14108,N_13882,N_13933);
nor U14109 (N_14109,N_13971,N_13999);
xnor U14110 (N_14110,N_13805,N_13868);
or U14111 (N_14111,N_13879,N_13991);
nor U14112 (N_14112,N_13858,N_13995);
and U14113 (N_14113,N_13982,N_13838);
xnor U14114 (N_14114,N_13877,N_13818);
nand U14115 (N_14115,N_13833,N_13929);
and U14116 (N_14116,N_13962,N_13831);
or U14117 (N_14117,N_13832,N_13847);
or U14118 (N_14118,N_13920,N_13814);
xor U14119 (N_14119,N_13925,N_13992);
or U14120 (N_14120,N_13976,N_13931);
nand U14121 (N_14121,N_13934,N_13805);
or U14122 (N_14122,N_13929,N_13994);
and U14123 (N_14123,N_13825,N_13810);
and U14124 (N_14124,N_13909,N_13924);
or U14125 (N_14125,N_13901,N_13805);
xnor U14126 (N_14126,N_13843,N_13845);
nor U14127 (N_14127,N_13947,N_13844);
nor U14128 (N_14128,N_13939,N_13837);
and U14129 (N_14129,N_13920,N_13895);
or U14130 (N_14130,N_13848,N_13839);
nor U14131 (N_14131,N_13889,N_13868);
nand U14132 (N_14132,N_13956,N_13949);
nand U14133 (N_14133,N_13971,N_13932);
nand U14134 (N_14134,N_13913,N_13808);
xnor U14135 (N_14135,N_13950,N_13970);
or U14136 (N_14136,N_13818,N_13976);
xor U14137 (N_14137,N_13940,N_13995);
and U14138 (N_14138,N_13821,N_13958);
xor U14139 (N_14139,N_13991,N_13803);
or U14140 (N_14140,N_13900,N_13922);
and U14141 (N_14141,N_13864,N_13947);
and U14142 (N_14142,N_13973,N_13921);
xnor U14143 (N_14143,N_13804,N_13816);
or U14144 (N_14144,N_13835,N_13913);
or U14145 (N_14145,N_13987,N_13904);
nor U14146 (N_14146,N_13923,N_13832);
nand U14147 (N_14147,N_13947,N_13940);
and U14148 (N_14148,N_13820,N_13895);
and U14149 (N_14149,N_13960,N_13943);
xor U14150 (N_14150,N_13929,N_13862);
and U14151 (N_14151,N_13862,N_13825);
and U14152 (N_14152,N_13848,N_13804);
nand U14153 (N_14153,N_13807,N_13933);
nor U14154 (N_14154,N_13900,N_13832);
xnor U14155 (N_14155,N_13946,N_13885);
and U14156 (N_14156,N_13915,N_13858);
and U14157 (N_14157,N_13955,N_13832);
xnor U14158 (N_14158,N_13805,N_13949);
or U14159 (N_14159,N_13808,N_13874);
nand U14160 (N_14160,N_13904,N_13975);
or U14161 (N_14161,N_13903,N_13981);
xor U14162 (N_14162,N_13856,N_13975);
xor U14163 (N_14163,N_13889,N_13956);
nor U14164 (N_14164,N_13837,N_13881);
xnor U14165 (N_14165,N_13994,N_13908);
nor U14166 (N_14166,N_13960,N_13981);
and U14167 (N_14167,N_13817,N_13831);
nor U14168 (N_14168,N_13838,N_13905);
nor U14169 (N_14169,N_13973,N_13803);
and U14170 (N_14170,N_13839,N_13805);
xor U14171 (N_14171,N_13957,N_13992);
xnor U14172 (N_14172,N_13826,N_13831);
or U14173 (N_14173,N_13804,N_13958);
or U14174 (N_14174,N_13885,N_13972);
and U14175 (N_14175,N_13805,N_13821);
or U14176 (N_14176,N_13969,N_13966);
nor U14177 (N_14177,N_13888,N_13833);
xnor U14178 (N_14178,N_13857,N_13874);
nor U14179 (N_14179,N_13936,N_13876);
or U14180 (N_14180,N_13893,N_13833);
or U14181 (N_14181,N_13890,N_13874);
nand U14182 (N_14182,N_13957,N_13817);
nor U14183 (N_14183,N_13912,N_13834);
or U14184 (N_14184,N_13943,N_13949);
nor U14185 (N_14185,N_13938,N_13808);
nand U14186 (N_14186,N_13963,N_13859);
nand U14187 (N_14187,N_13852,N_13907);
nor U14188 (N_14188,N_13820,N_13806);
nand U14189 (N_14189,N_13805,N_13952);
and U14190 (N_14190,N_13831,N_13840);
nor U14191 (N_14191,N_13843,N_13808);
nor U14192 (N_14192,N_13814,N_13973);
nor U14193 (N_14193,N_13933,N_13844);
nand U14194 (N_14194,N_13801,N_13888);
or U14195 (N_14195,N_13921,N_13915);
nor U14196 (N_14196,N_13968,N_13996);
xnor U14197 (N_14197,N_13816,N_13847);
or U14198 (N_14198,N_13890,N_13961);
or U14199 (N_14199,N_13802,N_13912);
nor U14200 (N_14200,N_14177,N_14163);
nand U14201 (N_14201,N_14054,N_14039);
or U14202 (N_14202,N_14183,N_14176);
nand U14203 (N_14203,N_14047,N_14118);
and U14204 (N_14204,N_14157,N_14065);
nand U14205 (N_14205,N_14015,N_14166);
xnor U14206 (N_14206,N_14044,N_14161);
and U14207 (N_14207,N_14007,N_14092);
xnor U14208 (N_14208,N_14142,N_14071);
nand U14209 (N_14209,N_14095,N_14067);
xnor U14210 (N_14210,N_14072,N_14005);
nand U14211 (N_14211,N_14091,N_14094);
or U14212 (N_14212,N_14050,N_14045);
and U14213 (N_14213,N_14162,N_14178);
and U14214 (N_14214,N_14035,N_14154);
and U14215 (N_14215,N_14002,N_14073);
nor U14216 (N_14216,N_14084,N_14048);
or U14217 (N_14217,N_14131,N_14099);
nand U14218 (N_14218,N_14160,N_14187);
and U14219 (N_14219,N_14025,N_14165);
xor U14220 (N_14220,N_14119,N_14192);
nand U14221 (N_14221,N_14128,N_14182);
or U14222 (N_14222,N_14129,N_14149);
nand U14223 (N_14223,N_14158,N_14138);
nand U14224 (N_14224,N_14191,N_14055);
nor U14225 (N_14225,N_14169,N_14133);
or U14226 (N_14226,N_14085,N_14125);
nand U14227 (N_14227,N_14179,N_14083);
and U14228 (N_14228,N_14031,N_14089);
nor U14229 (N_14229,N_14023,N_14021);
or U14230 (N_14230,N_14196,N_14051);
and U14231 (N_14231,N_14195,N_14028);
and U14232 (N_14232,N_14114,N_14103);
xnor U14233 (N_14233,N_14043,N_14074);
nor U14234 (N_14234,N_14136,N_14116);
and U14235 (N_14235,N_14170,N_14121);
nand U14236 (N_14236,N_14009,N_14061);
nand U14237 (N_14237,N_14145,N_14040);
and U14238 (N_14238,N_14171,N_14027);
xnor U14239 (N_14239,N_14020,N_14122);
or U14240 (N_14240,N_14042,N_14167);
or U14241 (N_14241,N_14175,N_14110);
nor U14242 (N_14242,N_14126,N_14102);
and U14243 (N_14243,N_14029,N_14077);
xnor U14244 (N_14244,N_14088,N_14150);
nand U14245 (N_14245,N_14198,N_14096);
nor U14246 (N_14246,N_14168,N_14033);
xor U14247 (N_14247,N_14185,N_14086);
or U14248 (N_14248,N_14057,N_14141);
or U14249 (N_14249,N_14014,N_14174);
nor U14250 (N_14250,N_14001,N_14069);
nand U14251 (N_14251,N_14004,N_14101);
nor U14252 (N_14252,N_14197,N_14063);
nor U14253 (N_14253,N_14107,N_14068);
nor U14254 (N_14254,N_14194,N_14013);
nor U14255 (N_14255,N_14104,N_14017);
xor U14256 (N_14256,N_14080,N_14180);
and U14257 (N_14257,N_14059,N_14036);
or U14258 (N_14258,N_14060,N_14124);
nand U14259 (N_14259,N_14159,N_14134);
xnor U14260 (N_14260,N_14010,N_14018);
xnor U14261 (N_14261,N_14115,N_14140);
and U14262 (N_14262,N_14112,N_14105);
and U14263 (N_14263,N_14032,N_14098);
nand U14264 (N_14264,N_14123,N_14144);
nor U14265 (N_14265,N_14082,N_14012);
xor U14266 (N_14266,N_14053,N_14111);
and U14267 (N_14267,N_14148,N_14188);
nand U14268 (N_14268,N_14070,N_14193);
and U14269 (N_14269,N_14135,N_14153);
and U14270 (N_14270,N_14143,N_14011);
or U14271 (N_14271,N_14147,N_14120);
nor U14272 (N_14272,N_14113,N_14041);
or U14273 (N_14273,N_14024,N_14189);
nand U14274 (N_14274,N_14156,N_14127);
xnor U14275 (N_14275,N_14130,N_14173);
nand U14276 (N_14276,N_14132,N_14003);
and U14277 (N_14277,N_14064,N_14181);
or U14278 (N_14278,N_14062,N_14037);
nor U14279 (N_14279,N_14038,N_14034);
or U14280 (N_14280,N_14093,N_14090);
nand U14281 (N_14281,N_14186,N_14058);
or U14282 (N_14282,N_14152,N_14076);
nand U14283 (N_14283,N_14078,N_14106);
and U14284 (N_14284,N_14155,N_14199);
nand U14285 (N_14285,N_14087,N_14172);
nor U14286 (N_14286,N_14146,N_14117);
or U14287 (N_14287,N_14164,N_14139);
nor U14288 (N_14288,N_14019,N_14056);
and U14289 (N_14289,N_14006,N_14097);
nand U14290 (N_14290,N_14046,N_14022);
nand U14291 (N_14291,N_14137,N_14052);
or U14292 (N_14292,N_14108,N_14075);
and U14293 (N_14293,N_14049,N_14079);
xnor U14294 (N_14294,N_14190,N_14000);
nor U14295 (N_14295,N_14184,N_14151);
and U14296 (N_14296,N_14081,N_14100);
xnor U14297 (N_14297,N_14066,N_14016);
nand U14298 (N_14298,N_14008,N_14030);
and U14299 (N_14299,N_14109,N_14026);
or U14300 (N_14300,N_14155,N_14170);
nor U14301 (N_14301,N_14010,N_14127);
and U14302 (N_14302,N_14154,N_14174);
nor U14303 (N_14303,N_14006,N_14188);
nor U14304 (N_14304,N_14076,N_14040);
or U14305 (N_14305,N_14043,N_14195);
or U14306 (N_14306,N_14026,N_14014);
and U14307 (N_14307,N_14065,N_14095);
or U14308 (N_14308,N_14027,N_14189);
nand U14309 (N_14309,N_14017,N_14172);
or U14310 (N_14310,N_14044,N_14177);
nor U14311 (N_14311,N_14110,N_14098);
nor U14312 (N_14312,N_14189,N_14026);
nor U14313 (N_14313,N_14025,N_14178);
nand U14314 (N_14314,N_14038,N_14061);
nand U14315 (N_14315,N_14095,N_14076);
or U14316 (N_14316,N_14115,N_14108);
nand U14317 (N_14317,N_14068,N_14123);
and U14318 (N_14318,N_14165,N_14190);
or U14319 (N_14319,N_14080,N_14079);
nand U14320 (N_14320,N_14004,N_14087);
or U14321 (N_14321,N_14071,N_14045);
nor U14322 (N_14322,N_14180,N_14058);
nor U14323 (N_14323,N_14042,N_14103);
xnor U14324 (N_14324,N_14159,N_14001);
nand U14325 (N_14325,N_14026,N_14119);
nor U14326 (N_14326,N_14079,N_14022);
or U14327 (N_14327,N_14122,N_14178);
and U14328 (N_14328,N_14152,N_14015);
xnor U14329 (N_14329,N_14086,N_14097);
nand U14330 (N_14330,N_14144,N_14039);
and U14331 (N_14331,N_14003,N_14155);
xnor U14332 (N_14332,N_14082,N_14001);
nor U14333 (N_14333,N_14060,N_14155);
and U14334 (N_14334,N_14011,N_14033);
or U14335 (N_14335,N_14007,N_14097);
nand U14336 (N_14336,N_14148,N_14083);
xnor U14337 (N_14337,N_14090,N_14086);
nand U14338 (N_14338,N_14037,N_14119);
or U14339 (N_14339,N_14133,N_14095);
xnor U14340 (N_14340,N_14063,N_14099);
xor U14341 (N_14341,N_14028,N_14031);
nand U14342 (N_14342,N_14012,N_14068);
nand U14343 (N_14343,N_14195,N_14181);
and U14344 (N_14344,N_14131,N_14070);
nand U14345 (N_14345,N_14068,N_14004);
nor U14346 (N_14346,N_14068,N_14031);
nor U14347 (N_14347,N_14080,N_14086);
nor U14348 (N_14348,N_14065,N_14167);
nand U14349 (N_14349,N_14074,N_14123);
nand U14350 (N_14350,N_14109,N_14066);
xor U14351 (N_14351,N_14185,N_14191);
and U14352 (N_14352,N_14143,N_14044);
xor U14353 (N_14353,N_14175,N_14181);
and U14354 (N_14354,N_14091,N_14003);
nand U14355 (N_14355,N_14101,N_14190);
xnor U14356 (N_14356,N_14090,N_14071);
xnor U14357 (N_14357,N_14048,N_14172);
and U14358 (N_14358,N_14108,N_14100);
and U14359 (N_14359,N_14028,N_14114);
nor U14360 (N_14360,N_14177,N_14063);
or U14361 (N_14361,N_14052,N_14149);
and U14362 (N_14362,N_14039,N_14068);
xor U14363 (N_14363,N_14109,N_14149);
xor U14364 (N_14364,N_14099,N_14082);
nor U14365 (N_14365,N_14134,N_14131);
or U14366 (N_14366,N_14131,N_14080);
or U14367 (N_14367,N_14096,N_14008);
and U14368 (N_14368,N_14098,N_14120);
nand U14369 (N_14369,N_14013,N_14075);
or U14370 (N_14370,N_14091,N_14048);
and U14371 (N_14371,N_14182,N_14097);
and U14372 (N_14372,N_14133,N_14128);
or U14373 (N_14373,N_14072,N_14071);
xnor U14374 (N_14374,N_14043,N_14099);
xor U14375 (N_14375,N_14102,N_14015);
nand U14376 (N_14376,N_14017,N_14049);
nand U14377 (N_14377,N_14160,N_14172);
xor U14378 (N_14378,N_14137,N_14158);
xnor U14379 (N_14379,N_14031,N_14032);
nor U14380 (N_14380,N_14073,N_14027);
nand U14381 (N_14381,N_14171,N_14102);
xor U14382 (N_14382,N_14032,N_14103);
xnor U14383 (N_14383,N_14054,N_14113);
and U14384 (N_14384,N_14098,N_14022);
and U14385 (N_14385,N_14086,N_14118);
nand U14386 (N_14386,N_14073,N_14159);
and U14387 (N_14387,N_14154,N_14031);
or U14388 (N_14388,N_14009,N_14114);
nand U14389 (N_14389,N_14133,N_14064);
xnor U14390 (N_14390,N_14075,N_14172);
or U14391 (N_14391,N_14139,N_14004);
xnor U14392 (N_14392,N_14034,N_14119);
or U14393 (N_14393,N_14157,N_14001);
or U14394 (N_14394,N_14124,N_14083);
xor U14395 (N_14395,N_14092,N_14099);
or U14396 (N_14396,N_14029,N_14064);
and U14397 (N_14397,N_14174,N_14148);
or U14398 (N_14398,N_14039,N_14147);
nand U14399 (N_14399,N_14107,N_14124);
or U14400 (N_14400,N_14288,N_14326);
and U14401 (N_14401,N_14366,N_14232);
or U14402 (N_14402,N_14221,N_14234);
nor U14403 (N_14403,N_14220,N_14299);
nor U14404 (N_14404,N_14292,N_14228);
and U14405 (N_14405,N_14338,N_14345);
xnor U14406 (N_14406,N_14357,N_14208);
and U14407 (N_14407,N_14371,N_14282);
or U14408 (N_14408,N_14304,N_14249);
xor U14409 (N_14409,N_14356,N_14364);
nand U14410 (N_14410,N_14312,N_14362);
nor U14411 (N_14411,N_14233,N_14311);
or U14412 (N_14412,N_14353,N_14397);
nor U14413 (N_14413,N_14358,N_14335);
xnor U14414 (N_14414,N_14274,N_14306);
or U14415 (N_14415,N_14206,N_14272);
nand U14416 (N_14416,N_14339,N_14333);
xor U14417 (N_14417,N_14226,N_14344);
nand U14418 (N_14418,N_14239,N_14201);
or U14419 (N_14419,N_14348,N_14278);
or U14420 (N_14420,N_14252,N_14260);
nor U14421 (N_14421,N_14317,N_14303);
xnor U14422 (N_14422,N_14385,N_14395);
nand U14423 (N_14423,N_14265,N_14238);
nand U14424 (N_14424,N_14396,N_14351);
xnor U14425 (N_14425,N_14318,N_14399);
or U14426 (N_14426,N_14286,N_14354);
or U14427 (N_14427,N_14222,N_14263);
or U14428 (N_14428,N_14322,N_14355);
or U14429 (N_14429,N_14219,N_14349);
and U14430 (N_14430,N_14380,N_14394);
nor U14431 (N_14431,N_14313,N_14264);
nand U14432 (N_14432,N_14370,N_14218);
and U14433 (N_14433,N_14331,N_14204);
or U14434 (N_14434,N_14393,N_14281);
or U14435 (N_14435,N_14254,N_14307);
xor U14436 (N_14436,N_14291,N_14375);
or U14437 (N_14437,N_14368,N_14310);
nor U14438 (N_14438,N_14323,N_14276);
or U14439 (N_14439,N_14308,N_14334);
nor U14440 (N_14440,N_14332,N_14285);
and U14441 (N_14441,N_14235,N_14301);
nor U14442 (N_14442,N_14298,N_14279);
or U14443 (N_14443,N_14329,N_14297);
xor U14444 (N_14444,N_14378,N_14256);
or U14445 (N_14445,N_14342,N_14271);
and U14446 (N_14446,N_14374,N_14365);
xor U14447 (N_14447,N_14248,N_14324);
or U14448 (N_14448,N_14215,N_14277);
nor U14449 (N_14449,N_14302,N_14346);
nand U14450 (N_14450,N_14316,N_14207);
nand U14451 (N_14451,N_14314,N_14259);
nor U14452 (N_14452,N_14245,N_14261);
and U14453 (N_14453,N_14305,N_14361);
nor U14454 (N_14454,N_14255,N_14360);
xor U14455 (N_14455,N_14251,N_14262);
nor U14456 (N_14456,N_14376,N_14379);
nor U14457 (N_14457,N_14347,N_14266);
nand U14458 (N_14458,N_14367,N_14283);
xnor U14459 (N_14459,N_14328,N_14389);
xor U14460 (N_14460,N_14216,N_14212);
nor U14461 (N_14461,N_14381,N_14223);
and U14462 (N_14462,N_14227,N_14398);
nor U14463 (N_14463,N_14315,N_14372);
nor U14464 (N_14464,N_14280,N_14236);
and U14465 (N_14465,N_14203,N_14242);
or U14466 (N_14466,N_14273,N_14294);
or U14467 (N_14467,N_14268,N_14341);
nand U14468 (N_14468,N_14296,N_14246);
and U14469 (N_14469,N_14267,N_14230);
nand U14470 (N_14470,N_14247,N_14244);
xnor U14471 (N_14471,N_14373,N_14386);
and U14472 (N_14472,N_14388,N_14391);
nor U14473 (N_14473,N_14257,N_14213);
and U14474 (N_14474,N_14340,N_14327);
nand U14475 (N_14475,N_14295,N_14319);
nor U14476 (N_14476,N_14224,N_14231);
nand U14477 (N_14477,N_14336,N_14337);
nand U14478 (N_14478,N_14211,N_14275);
nand U14479 (N_14479,N_14377,N_14320);
nand U14480 (N_14480,N_14350,N_14250);
or U14481 (N_14481,N_14321,N_14392);
nor U14482 (N_14482,N_14383,N_14258);
or U14483 (N_14483,N_14229,N_14343);
and U14484 (N_14484,N_14205,N_14359);
and U14485 (N_14485,N_14225,N_14243);
and U14486 (N_14486,N_14330,N_14210);
and U14487 (N_14487,N_14202,N_14269);
and U14488 (N_14488,N_14309,N_14382);
nor U14489 (N_14489,N_14352,N_14387);
xor U14490 (N_14490,N_14237,N_14284);
and U14491 (N_14491,N_14270,N_14287);
nand U14492 (N_14492,N_14325,N_14369);
nor U14493 (N_14493,N_14240,N_14217);
nor U14494 (N_14494,N_14290,N_14390);
or U14495 (N_14495,N_14209,N_14300);
nand U14496 (N_14496,N_14241,N_14363);
xor U14497 (N_14497,N_14289,N_14253);
or U14498 (N_14498,N_14384,N_14200);
or U14499 (N_14499,N_14214,N_14293);
or U14500 (N_14500,N_14375,N_14299);
xnor U14501 (N_14501,N_14331,N_14303);
or U14502 (N_14502,N_14205,N_14349);
and U14503 (N_14503,N_14213,N_14295);
nand U14504 (N_14504,N_14320,N_14339);
xor U14505 (N_14505,N_14386,N_14358);
xnor U14506 (N_14506,N_14301,N_14354);
and U14507 (N_14507,N_14250,N_14345);
nand U14508 (N_14508,N_14247,N_14238);
nand U14509 (N_14509,N_14335,N_14251);
or U14510 (N_14510,N_14252,N_14291);
xnor U14511 (N_14511,N_14241,N_14201);
or U14512 (N_14512,N_14390,N_14224);
or U14513 (N_14513,N_14396,N_14335);
and U14514 (N_14514,N_14357,N_14367);
nand U14515 (N_14515,N_14396,N_14237);
or U14516 (N_14516,N_14268,N_14378);
or U14517 (N_14517,N_14299,N_14221);
nor U14518 (N_14518,N_14305,N_14379);
nor U14519 (N_14519,N_14331,N_14335);
nor U14520 (N_14520,N_14332,N_14334);
nand U14521 (N_14521,N_14310,N_14231);
and U14522 (N_14522,N_14214,N_14271);
xor U14523 (N_14523,N_14352,N_14336);
and U14524 (N_14524,N_14328,N_14369);
or U14525 (N_14525,N_14361,N_14395);
or U14526 (N_14526,N_14290,N_14264);
nor U14527 (N_14527,N_14218,N_14242);
nor U14528 (N_14528,N_14296,N_14208);
and U14529 (N_14529,N_14392,N_14387);
and U14530 (N_14530,N_14224,N_14308);
xnor U14531 (N_14531,N_14200,N_14220);
xor U14532 (N_14532,N_14266,N_14238);
or U14533 (N_14533,N_14209,N_14311);
nand U14534 (N_14534,N_14299,N_14393);
nand U14535 (N_14535,N_14377,N_14317);
xor U14536 (N_14536,N_14229,N_14359);
nor U14537 (N_14537,N_14394,N_14270);
xnor U14538 (N_14538,N_14271,N_14333);
nor U14539 (N_14539,N_14287,N_14265);
nand U14540 (N_14540,N_14335,N_14391);
nor U14541 (N_14541,N_14234,N_14397);
nand U14542 (N_14542,N_14203,N_14285);
xor U14543 (N_14543,N_14258,N_14366);
or U14544 (N_14544,N_14278,N_14374);
xnor U14545 (N_14545,N_14287,N_14340);
or U14546 (N_14546,N_14259,N_14369);
or U14547 (N_14547,N_14356,N_14387);
and U14548 (N_14548,N_14229,N_14296);
nand U14549 (N_14549,N_14395,N_14277);
or U14550 (N_14550,N_14335,N_14387);
nand U14551 (N_14551,N_14397,N_14268);
nor U14552 (N_14552,N_14358,N_14227);
and U14553 (N_14553,N_14311,N_14344);
xor U14554 (N_14554,N_14316,N_14375);
nor U14555 (N_14555,N_14356,N_14346);
or U14556 (N_14556,N_14220,N_14388);
xnor U14557 (N_14557,N_14285,N_14290);
nor U14558 (N_14558,N_14273,N_14340);
and U14559 (N_14559,N_14228,N_14238);
or U14560 (N_14560,N_14246,N_14331);
nand U14561 (N_14561,N_14244,N_14214);
nand U14562 (N_14562,N_14355,N_14253);
and U14563 (N_14563,N_14293,N_14381);
or U14564 (N_14564,N_14316,N_14338);
xor U14565 (N_14565,N_14335,N_14257);
and U14566 (N_14566,N_14200,N_14266);
nor U14567 (N_14567,N_14337,N_14328);
xor U14568 (N_14568,N_14234,N_14207);
or U14569 (N_14569,N_14260,N_14223);
and U14570 (N_14570,N_14383,N_14343);
xor U14571 (N_14571,N_14303,N_14230);
and U14572 (N_14572,N_14317,N_14339);
or U14573 (N_14573,N_14218,N_14303);
or U14574 (N_14574,N_14349,N_14376);
nor U14575 (N_14575,N_14261,N_14343);
or U14576 (N_14576,N_14314,N_14297);
xor U14577 (N_14577,N_14365,N_14338);
nand U14578 (N_14578,N_14352,N_14368);
or U14579 (N_14579,N_14267,N_14273);
or U14580 (N_14580,N_14334,N_14242);
nand U14581 (N_14581,N_14387,N_14360);
or U14582 (N_14582,N_14276,N_14259);
nand U14583 (N_14583,N_14260,N_14229);
or U14584 (N_14584,N_14261,N_14288);
and U14585 (N_14585,N_14341,N_14350);
and U14586 (N_14586,N_14305,N_14277);
and U14587 (N_14587,N_14204,N_14384);
nand U14588 (N_14588,N_14238,N_14257);
xor U14589 (N_14589,N_14388,N_14240);
and U14590 (N_14590,N_14318,N_14236);
nand U14591 (N_14591,N_14332,N_14333);
xor U14592 (N_14592,N_14269,N_14399);
nor U14593 (N_14593,N_14231,N_14356);
nand U14594 (N_14594,N_14259,N_14364);
nand U14595 (N_14595,N_14295,N_14332);
nand U14596 (N_14596,N_14208,N_14379);
or U14597 (N_14597,N_14238,N_14395);
or U14598 (N_14598,N_14209,N_14240);
and U14599 (N_14599,N_14242,N_14336);
nor U14600 (N_14600,N_14496,N_14548);
xnor U14601 (N_14601,N_14526,N_14454);
and U14602 (N_14602,N_14457,N_14512);
and U14603 (N_14603,N_14467,N_14460);
or U14604 (N_14604,N_14596,N_14519);
nor U14605 (N_14605,N_14417,N_14456);
nor U14606 (N_14606,N_14589,N_14546);
xor U14607 (N_14607,N_14579,N_14432);
nor U14608 (N_14608,N_14573,N_14483);
or U14609 (N_14609,N_14464,N_14592);
or U14610 (N_14610,N_14488,N_14420);
and U14611 (N_14611,N_14451,N_14528);
xnor U14612 (N_14612,N_14449,N_14470);
and U14613 (N_14613,N_14561,N_14510);
nor U14614 (N_14614,N_14490,N_14511);
xnor U14615 (N_14615,N_14495,N_14473);
nand U14616 (N_14616,N_14506,N_14503);
or U14617 (N_14617,N_14431,N_14418);
and U14618 (N_14618,N_14499,N_14577);
and U14619 (N_14619,N_14400,N_14582);
xnor U14620 (N_14620,N_14500,N_14494);
and U14621 (N_14621,N_14481,N_14521);
xnor U14622 (N_14622,N_14446,N_14474);
xnor U14623 (N_14623,N_14547,N_14448);
or U14624 (N_14624,N_14513,N_14586);
and U14625 (N_14625,N_14404,N_14437);
or U14626 (N_14626,N_14566,N_14529);
and U14627 (N_14627,N_14476,N_14570);
and U14628 (N_14628,N_14416,N_14421);
nand U14629 (N_14629,N_14556,N_14405);
or U14630 (N_14630,N_14507,N_14508);
xnor U14631 (N_14631,N_14563,N_14537);
nand U14632 (N_14632,N_14409,N_14591);
nor U14633 (N_14633,N_14514,N_14518);
xor U14634 (N_14634,N_14434,N_14545);
or U14635 (N_14635,N_14465,N_14455);
nand U14636 (N_14636,N_14452,N_14433);
and U14637 (N_14637,N_14584,N_14410);
xnor U14638 (N_14638,N_14472,N_14462);
xnor U14639 (N_14639,N_14402,N_14539);
and U14640 (N_14640,N_14517,N_14498);
nand U14641 (N_14641,N_14492,N_14453);
nor U14642 (N_14642,N_14493,N_14558);
or U14643 (N_14643,N_14590,N_14485);
and U14644 (N_14644,N_14530,N_14542);
or U14645 (N_14645,N_14435,N_14594);
nand U14646 (N_14646,N_14466,N_14569);
nor U14647 (N_14647,N_14543,N_14536);
or U14648 (N_14648,N_14475,N_14480);
nand U14649 (N_14649,N_14436,N_14599);
nand U14650 (N_14650,N_14580,N_14430);
and U14651 (N_14651,N_14497,N_14427);
nand U14652 (N_14652,N_14549,N_14585);
nor U14653 (N_14653,N_14415,N_14560);
xnor U14654 (N_14654,N_14422,N_14419);
xnor U14655 (N_14655,N_14444,N_14524);
nor U14656 (N_14656,N_14406,N_14438);
and U14657 (N_14657,N_14450,N_14403);
nor U14658 (N_14658,N_14571,N_14552);
or U14659 (N_14659,N_14491,N_14443);
or U14660 (N_14660,N_14550,N_14505);
and U14661 (N_14661,N_14463,N_14482);
or U14662 (N_14662,N_14534,N_14429);
and U14663 (N_14663,N_14414,N_14554);
xor U14664 (N_14664,N_14559,N_14544);
xnor U14665 (N_14665,N_14595,N_14515);
nand U14666 (N_14666,N_14447,N_14562);
nor U14667 (N_14667,N_14459,N_14413);
xor U14668 (N_14668,N_14442,N_14535);
nor U14669 (N_14669,N_14441,N_14531);
or U14670 (N_14670,N_14458,N_14479);
nor U14671 (N_14671,N_14557,N_14461);
and U14672 (N_14672,N_14407,N_14439);
and U14673 (N_14673,N_14471,N_14408);
and U14674 (N_14674,N_14587,N_14489);
nand U14675 (N_14675,N_14551,N_14581);
nand U14676 (N_14676,N_14525,N_14477);
and U14677 (N_14677,N_14541,N_14469);
or U14678 (N_14678,N_14574,N_14423);
xnor U14679 (N_14679,N_14411,N_14468);
nor U14680 (N_14680,N_14401,N_14440);
xnor U14681 (N_14681,N_14598,N_14538);
xnor U14682 (N_14682,N_14568,N_14578);
nand U14683 (N_14683,N_14553,N_14509);
nor U14684 (N_14684,N_14588,N_14478);
or U14685 (N_14685,N_14564,N_14501);
nand U14686 (N_14686,N_14425,N_14487);
nand U14687 (N_14687,N_14576,N_14565);
and U14688 (N_14688,N_14502,N_14412);
or U14689 (N_14689,N_14424,N_14567);
nand U14690 (N_14690,N_14428,N_14523);
xor U14691 (N_14691,N_14593,N_14504);
and U14692 (N_14692,N_14516,N_14540);
nor U14693 (N_14693,N_14445,N_14575);
nand U14694 (N_14694,N_14583,N_14532);
xor U14695 (N_14695,N_14486,N_14522);
and U14696 (N_14696,N_14555,N_14533);
nand U14697 (N_14697,N_14520,N_14527);
nand U14698 (N_14698,N_14426,N_14597);
nand U14699 (N_14699,N_14572,N_14484);
and U14700 (N_14700,N_14523,N_14492);
xnor U14701 (N_14701,N_14567,N_14517);
xnor U14702 (N_14702,N_14543,N_14582);
nand U14703 (N_14703,N_14500,N_14506);
nor U14704 (N_14704,N_14597,N_14414);
nor U14705 (N_14705,N_14530,N_14480);
xor U14706 (N_14706,N_14572,N_14524);
nor U14707 (N_14707,N_14562,N_14551);
nand U14708 (N_14708,N_14556,N_14422);
nand U14709 (N_14709,N_14434,N_14596);
nand U14710 (N_14710,N_14500,N_14544);
nor U14711 (N_14711,N_14452,N_14535);
nand U14712 (N_14712,N_14402,N_14583);
nor U14713 (N_14713,N_14471,N_14586);
xnor U14714 (N_14714,N_14400,N_14487);
and U14715 (N_14715,N_14498,N_14580);
xor U14716 (N_14716,N_14552,N_14541);
or U14717 (N_14717,N_14440,N_14499);
nor U14718 (N_14718,N_14511,N_14504);
nor U14719 (N_14719,N_14528,N_14468);
nor U14720 (N_14720,N_14563,N_14419);
xnor U14721 (N_14721,N_14550,N_14461);
and U14722 (N_14722,N_14546,N_14407);
nand U14723 (N_14723,N_14477,N_14567);
nand U14724 (N_14724,N_14433,N_14510);
or U14725 (N_14725,N_14440,N_14443);
nand U14726 (N_14726,N_14408,N_14430);
or U14727 (N_14727,N_14523,N_14463);
xor U14728 (N_14728,N_14560,N_14458);
xor U14729 (N_14729,N_14503,N_14546);
nand U14730 (N_14730,N_14499,N_14543);
and U14731 (N_14731,N_14557,N_14494);
or U14732 (N_14732,N_14435,N_14595);
or U14733 (N_14733,N_14582,N_14523);
nand U14734 (N_14734,N_14421,N_14579);
and U14735 (N_14735,N_14467,N_14576);
nand U14736 (N_14736,N_14563,N_14462);
nand U14737 (N_14737,N_14465,N_14577);
and U14738 (N_14738,N_14502,N_14559);
and U14739 (N_14739,N_14558,N_14502);
nor U14740 (N_14740,N_14557,N_14427);
or U14741 (N_14741,N_14496,N_14515);
or U14742 (N_14742,N_14419,N_14400);
xor U14743 (N_14743,N_14584,N_14428);
nor U14744 (N_14744,N_14427,N_14561);
nand U14745 (N_14745,N_14479,N_14493);
nand U14746 (N_14746,N_14400,N_14511);
or U14747 (N_14747,N_14575,N_14560);
nor U14748 (N_14748,N_14459,N_14418);
or U14749 (N_14749,N_14564,N_14511);
nand U14750 (N_14750,N_14441,N_14455);
nor U14751 (N_14751,N_14549,N_14554);
or U14752 (N_14752,N_14543,N_14574);
or U14753 (N_14753,N_14519,N_14574);
and U14754 (N_14754,N_14544,N_14442);
or U14755 (N_14755,N_14542,N_14471);
or U14756 (N_14756,N_14525,N_14423);
and U14757 (N_14757,N_14573,N_14443);
and U14758 (N_14758,N_14541,N_14564);
nand U14759 (N_14759,N_14403,N_14495);
nor U14760 (N_14760,N_14462,N_14525);
nor U14761 (N_14761,N_14459,N_14495);
nor U14762 (N_14762,N_14400,N_14569);
and U14763 (N_14763,N_14509,N_14568);
nand U14764 (N_14764,N_14572,N_14515);
nand U14765 (N_14765,N_14557,N_14567);
nor U14766 (N_14766,N_14570,N_14482);
nor U14767 (N_14767,N_14433,N_14482);
nor U14768 (N_14768,N_14414,N_14431);
or U14769 (N_14769,N_14513,N_14518);
nand U14770 (N_14770,N_14464,N_14539);
xnor U14771 (N_14771,N_14480,N_14516);
nor U14772 (N_14772,N_14424,N_14437);
nand U14773 (N_14773,N_14438,N_14548);
nand U14774 (N_14774,N_14550,N_14543);
nor U14775 (N_14775,N_14409,N_14554);
and U14776 (N_14776,N_14513,N_14401);
xor U14777 (N_14777,N_14531,N_14592);
and U14778 (N_14778,N_14493,N_14457);
or U14779 (N_14779,N_14596,N_14590);
xor U14780 (N_14780,N_14568,N_14495);
nand U14781 (N_14781,N_14505,N_14514);
nand U14782 (N_14782,N_14509,N_14413);
nand U14783 (N_14783,N_14521,N_14439);
nand U14784 (N_14784,N_14537,N_14453);
nor U14785 (N_14785,N_14567,N_14417);
xnor U14786 (N_14786,N_14430,N_14558);
nor U14787 (N_14787,N_14495,N_14578);
nand U14788 (N_14788,N_14572,N_14414);
and U14789 (N_14789,N_14448,N_14596);
nand U14790 (N_14790,N_14415,N_14517);
and U14791 (N_14791,N_14483,N_14519);
and U14792 (N_14792,N_14492,N_14558);
and U14793 (N_14793,N_14426,N_14451);
or U14794 (N_14794,N_14485,N_14517);
nor U14795 (N_14795,N_14599,N_14476);
and U14796 (N_14796,N_14587,N_14493);
or U14797 (N_14797,N_14473,N_14590);
and U14798 (N_14798,N_14486,N_14561);
xor U14799 (N_14799,N_14537,N_14526);
and U14800 (N_14800,N_14666,N_14765);
and U14801 (N_14801,N_14726,N_14774);
xor U14802 (N_14802,N_14766,N_14636);
nor U14803 (N_14803,N_14788,N_14735);
and U14804 (N_14804,N_14678,N_14684);
nand U14805 (N_14805,N_14694,N_14600);
or U14806 (N_14806,N_14629,N_14702);
xor U14807 (N_14807,N_14653,N_14752);
and U14808 (N_14808,N_14637,N_14606);
or U14809 (N_14809,N_14633,N_14767);
xor U14810 (N_14810,N_14796,N_14623);
and U14811 (N_14811,N_14727,N_14621);
nor U14812 (N_14812,N_14772,N_14614);
and U14813 (N_14813,N_14649,N_14618);
nand U14814 (N_14814,N_14696,N_14699);
or U14815 (N_14815,N_14622,N_14603);
nor U14816 (N_14816,N_14660,N_14758);
nand U14817 (N_14817,N_14697,N_14707);
or U14818 (N_14818,N_14646,N_14680);
nand U14819 (N_14819,N_14668,N_14651);
and U14820 (N_14820,N_14741,N_14672);
nand U14821 (N_14821,N_14626,N_14683);
or U14822 (N_14822,N_14768,N_14676);
nor U14823 (N_14823,N_14662,N_14799);
and U14824 (N_14824,N_14777,N_14793);
or U14825 (N_14825,N_14643,N_14756);
or U14826 (N_14826,N_14703,N_14748);
xnor U14827 (N_14827,N_14700,N_14667);
or U14828 (N_14828,N_14740,N_14632);
xor U14829 (N_14829,N_14721,N_14784);
nor U14830 (N_14830,N_14719,N_14785);
and U14831 (N_14831,N_14664,N_14717);
xor U14832 (N_14832,N_14640,N_14731);
or U14833 (N_14833,N_14779,N_14620);
and U14834 (N_14834,N_14677,N_14709);
nor U14835 (N_14835,N_14669,N_14624);
nor U14836 (N_14836,N_14608,N_14751);
xnor U14837 (N_14837,N_14628,N_14760);
or U14838 (N_14838,N_14745,N_14659);
and U14839 (N_14839,N_14671,N_14638);
nor U14840 (N_14840,N_14790,N_14673);
nand U14841 (N_14841,N_14698,N_14795);
nor U14842 (N_14842,N_14681,N_14786);
xnor U14843 (N_14843,N_14607,N_14674);
nor U14844 (N_14844,N_14687,N_14647);
and U14845 (N_14845,N_14754,N_14782);
nor U14846 (N_14846,N_14652,N_14729);
xor U14847 (N_14847,N_14743,N_14613);
or U14848 (N_14848,N_14794,N_14757);
xnor U14849 (N_14849,N_14797,N_14675);
nand U14850 (N_14850,N_14690,N_14691);
xor U14851 (N_14851,N_14755,N_14693);
xor U14852 (N_14852,N_14711,N_14761);
and U14853 (N_14853,N_14789,N_14645);
and U14854 (N_14854,N_14686,N_14715);
and U14855 (N_14855,N_14712,N_14734);
nand U14856 (N_14856,N_14695,N_14737);
xor U14857 (N_14857,N_14762,N_14612);
nand U14858 (N_14858,N_14625,N_14769);
and U14859 (N_14859,N_14639,N_14778);
nand U14860 (N_14860,N_14724,N_14749);
nor U14861 (N_14861,N_14601,N_14764);
nand U14862 (N_14862,N_14641,N_14630);
xnor U14863 (N_14863,N_14609,N_14776);
and U14864 (N_14864,N_14615,N_14663);
nor U14865 (N_14865,N_14605,N_14661);
or U14866 (N_14866,N_14736,N_14720);
xnor U14867 (N_14867,N_14656,N_14705);
and U14868 (N_14868,N_14679,N_14708);
nand U14869 (N_14869,N_14792,N_14682);
nor U14870 (N_14870,N_14723,N_14791);
nor U14871 (N_14871,N_14604,N_14798);
xor U14872 (N_14872,N_14617,N_14710);
nor U14873 (N_14873,N_14732,N_14718);
nand U14874 (N_14874,N_14773,N_14787);
nor U14875 (N_14875,N_14689,N_14739);
or U14876 (N_14876,N_14714,N_14619);
nand U14877 (N_14877,N_14750,N_14781);
nand U14878 (N_14878,N_14627,N_14610);
or U14879 (N_14879,N_14692,N_14780);
and U14880 (N_14880,N_14763,N_14611);
or U14881 (N_14881,N_14706,N_14701);
and U14882 (N_14882,N_14704,N_14733);
nand U14883 (N_14883,N_14747,N_14713);
and U14884 (N_14884,N_14730,N_14644);
nor U14885 (N_14885,N_14658,N_14771);
nor U14886 (N_14886,N_14746,N_14616);
nor U14887 (N_14887,N_14670,N_14770);
nand U14888 (N_14888,N_14602,N_14655);
xnor U14889 (N_14889,N_14744,N_14631);
xnor U14890 (N_14890,N_14759,N_14738);
nor U14891 (N_14891,N_14634,N_14725);
xnor U14892 (N_14892,N_14783,N_14742);
nand U14893 (N_14893,N_14635,N_14688);
xor U14894 (N_14894,N_14654,N_14775);
nand U14895 (N_14895,N_14665,N_14728);
or U14896 (N_14896,N_14642,N_14657);
nand U14897 (N_14897,N_14685,N_14650);
or U14898 (N_14898,N_14716,N_14648);
nand U14899 (N_14899,N_14722,N_14753);
nand U14900 (N_14900,N_14600,N_14783);
xnor U14901 (N_14901,N_14628,N_14681);
xnor U14902 (N_14902,N_14611,N_14738);
nand U14903 (N_14903,N_14635,N_14754);
nand U14904 (N_14904,N_14794,N_14626);
and U14905 (N_14905,N_14740,N_14607);
xnor U14906 (N_14906,N_14701,N_14764);
xnor U14907 (N_14907,N_14756,N_14613);
nor U14908 (N_14908,N_14703,N_14662);
nor U14909 (N_14909,N_14787,N_14669);
nand U14910 (N_14910,N_14624,N_14714);
xnor U14911 (N_14911,N_14723,N_14637);
or U14912 (N_14912,N_14797,N_14629);
nor U14913 (N_14913,N_14608,N_14619);
or U14914 (N_14914,N_14636,N_14610);
or U14915 (N_14915,N_14797,N_14799);
nand U14916 (N_14916,N_14687,N_14646);
nand U14917 (N_14917,N_14746,N_14695);
xor U14918 (N_14918,N_14630,N_14780);
and U14919 (N_14919,N_14740,N_14725);
xnor U14920 (N_14920,N_14762,N_14640);
nor U14921 (N_14921,N_14708,N_14686);
xor U14922 (N_14922,N_14790,N_14758);
xnor U14923 (N_14923,N_14767,N_14662);
xnor U14924 (N_14924,N_14743,N_14736);
and U14925 (N_14925,N_14641,N_14773);
nand U14926 (N_14926,N_14733,N_14743);
xor U14927 (N_14927,N_14638,N_14695);
xnor U14928 (N_14928,N_14681,N_14768);
nor U14929 (N_14929,N_14621,N_14667);
or U14930 (N_14930,N_14707,N_14757);
nand U14931 (N_14931,N_14603,N_14651);
and U14932 (N_14932,N_14612,N_14631);
or U14933 (N_14933,N_14600,N_14765);
xnor U14934 (N_14934,N_14641,N_14622);
or U14935 (N_14935,N_14691,N_14706);
nand U14936 (N_14936,N_14644,N_14610);
nand U14937 (N_14937,N_14655,N_14680);
xnor U14938 (N_14938,N_14725,N_14649);
and U14939 (N_14939,N_14603,N_14701);
and U14940 (N_14940,N_14731,N_14649);
and U14941 (N_14941,N_14725,N_14647);
and U14942 (N_14942,N_14753,N_14713);
nand U14943 (N_14943,N_14772,N_14745);
nor U14944 (N_14944,N_14760,N_14724);
and U14945 (N_14945,N_14625,N_14718);
nand U14946 (N_14946,N_14617,N_14668);
nand U14947 (N_14947,N_14664,N_14762);
nor U14948 (N_14948,N_14618,N_14622);
and U14949 (N_14949,N_14649,N_14796);
xnor U14950 (N_14950,N_14765,N_14745);
nand U14951 (N_14951,N_14782,N_14734);
xor U14952 (N_14952,N_14633,N_14677);
or U14953 (N_14953,N_14705,N_14626);
nand U14954 (N_14954,N_14695,N_14618);
or U14955 (N_14955,N_14754,N_14785);
or U14956 (N_14956,N_14643,N_14600);
or U14957 (N_14957,N_14749,N_14650);
nand U14958 (N_14958,N_14683,N_14624);
nor U14959 (N_14959,N_14680,N_14662);
xor U14960 (N_14960,N_14695,N_14674);
or U14961 (N_14961,N_14716,N_14607);
and U14962 (N_14962,N_14705,N_14799);
nand U14963 (N_14963,N_14603,N_14745);
or U14964 (N_14964,N_14642,N_14704);
and U14965 (N_14965,N_14764,N_14647);
xor U14966 (N_14966,N_14775,N_14612);
and U14967 (N_14967,N_14756,N_14647);
or U14968 (N_14968,N_14697,N_14656);
nand U14969 (N_14969,N_14605,N_14755);
and U14970 (N_14970,N_14651,N_14699);
nand U14971 (N_14971,N_14763,N_14681);
nor U14972 (N_14972,N_14710,N_14643);
xnor U14973 (N_14973,N_14784,N_14793);
nor U14974 (N_14974,N_14616,N_14727);
or U14975 (N_14975,N_14746,N_14622);
or U14976 (N_14976,N_14705,N_14679);
or U14977 (N_14977,N_14787,N_14659);
nand U14978 (N_14978,N_14738,N_14794);
nor U14979 (N_14979,N_14600,N_14636);
xnor U14980 (N_14980,N_14751,N_14605);
nand U14981 (N_14981,N_14794,N_14643);
or U14982 (N_14982,N_14701,N_14688);
nor U14983 (N_14983,N_14692,N_14661);
or U14984 (N_14984,N_14790,N_14708);
xnor U14985 (N_14985,N_14677,N_14771);
nor U14986 (N_14986,N_14658,N_14619);
or U14987 (N_14987,N_14614,N_14717);
nor U14988 (N_14988,N_14664,N_14637);
and U14989 (N_14989,N_14615,N_14724);
or U14990 (N_14990,N_14745,N_14712);
nor U14991 (N_14991,N_14672,N_14700);
nand U14992 (N_14992,N_14625,N_14780);
xor U14993 (N_14993,N_14698,N_14793);
and U14994 (N_14994,N_14796,N_14752);
nand U14995 (N_14995,N_14716,N_14686);
or U14996 (N_14996,N_14739,N_14658);
and U14997 (N_14997,N_14776,N_14742);
or U14998 (N_14998,N_14743,N_14609);
nand U14999 (N_14999,N_14604,N_14651);
and UO_0 (O_0,N_14965,N_14906);
and UO_1 (O_1,N_14988,N_14838);
nor UO_2 (O_2,N_14928,N_14954);
and UO_3 (O_3,N_14829,N_14995);
nand UO_4 (O_4,N_14827,N_14972);
and UO_5 (O_5,N_14914,N_14835);
or UO_6 (O_6,N_14953,N_14824);
xnor UO_7 (O_7,N_14861,N_14854);
or UO_8 (O_8,N_14911,N_14934);
or UO_9 (O_9,N_14918,N_14933);
and UO_10 (O_10,N_14804,N_14836);
xnor UO_11 (O_11,N_14971,N_14922);
xor UO_12 (O_12,N_14974,N_14999);
nand UO_13 (O_13,N_14980,N_14812);
nor UO_14 (O_14,N_14832,N_14864);
nor UO_15 (O_15,N_14927,N_14975);
nand UO_16 (O_16,N_14917,N_14948);
or UO_17 (O_17,N_14963,N_14936);
and UO_18 (O_18,N_14913,N_14968);
xor UO_19 (O_19,N_14805,N_14970);
xnor UO_20 (O_20,N_14895,N_14900);
or UO_21 (O_21,N_14935,N_14855);
or UO_22 (O_22,N_14820,N_14811);
or UO_23 (O_23,N_14964,N_14976);
nor UO_24 (O_24,N_14857,N_14881);
xor UO_25 (O_25,N_14916,N_14834);
and UO_26 (O_26,N_14956,N_14991);
xor UO_27 (O_27,N_14915,N_14908);
or UO_28 (O_28,N_14808,N_14907);
xor UO_29 (O_29,N_14890,N_14880);
and UO_30 (O_30,N_14868,N_14875);
xnor UO_31 (O_31,N_14951,N_14990);
or UO_32 (O_32,N_14982,N_14967);
and UO_33 (O_33,N_14831,N_14814);
xnor UO_34 (O_34,N_14940,N_14958);
nand UO_35 (O_35,N_14941,N_14952);
or UO_36 (O_36,N_14874,N_14978);
or UO_37 (O_37,N_14993,N_14893);
xor UO_38 (O_38,N_14889,N_14830);
nor UO_39 (O_39,N_14984,N_14858);
or UO_40 (O_40,N_14870,N_14803);
nor UO_41 (O_41,N_14939,N_14949);
xor UO_42 (O_42,N_14816,N_14866);
or UO_43 (O_43,N_14871,N_14960);
and UO_44 (O_44,N_14903,N_14989);
and UO_45 (O_45,N_14878,N_14986);
nand UO_46 (O_46,N_14801,N_14846);
nand UO_47 (O_47,N_14912,N_14959);
and UO_48 (O_48,N_14902,N_14886);
xnor UO_49 (O_49,N_14867,N_14942);
or UO_50 (O_50,N_14904,N_14810);
or UO_51 (O_51,N_14969,N_14894);
nand UO_52 (O_52,N_14840,N_14802);
and UO_53 (O_53,N_14966,N_14909);
and UO_54 (O_54,N_14845,N_14828);
and UO_55 (O_55,N_14926,N_14821);
nand UO_56 (O_56,N_14979,N_14947);
or UO_57 (O_57,N_14925,N_14860);
and UO_58 (O_58,N_14872,N_14937);
nand UO_59 (O_59,N_14806,N_14882);
and UO_60 (O_60,N_14851,N_14932);
nand UO_61 (O_61,N_14887,N_14961);
xor UO_62 (O_62,N_14877,N_14849);
or UO_63 (O_63,N_14847,N_14823);
nor UO_64 (O_64,N_14957,N_14873);
nand UO_65 (O_65,N_14833,N_14899);
nor UO_66 (O_66,N_14891,N_14837);
xor UO_67 (O_67,N_14905,N_14946);
and UO_68 (O_68,N_14930,N_14992);
xnor UO_69 (O_69,N_14910,N_14973);
and UO_70 (O_70,N_14862,N_14825);
xor UO_71 (O_71,N_14997,N_14852);
xor UO_72 (O_72,N_14998,N_14839);
or UO_73 (O_73,N_14843,N_14955);
nor UO_74 (O_74,N_14817,N_14885);
and UO_75 (O_75,N_14938,N_14931);
xor UO_76 (O_76,N_14853,N_14841);
nor UO_77 (O_77,N_14818,N_14856);
nor UO_78 (O_78,N_14994,N_14859);
xnor UO_79 (O_79,N_14815,N_14985);
xnor UO_80 (O_80,N_14924,N_14896);
xnor UO_81 (O_81,N_14883,N_14923);
nor UO_82 (O_82,N_14983,N_14865);
nor UO_83 (O_83,N_14897,N_14842);
or UO_84 (O_84,N_14879,N_14950);
and UO_85 (O_85,N_14826,N_14807);
xor UO_86 (O_86,N_14876,N_14929);
or UO_87 (O_87,N_14850,N_14863);
nor UO_88 (O_88,N_14848,N_14981);
or UO_89 (O_89,N_14987,N_14844);
or UO_90 (O_90,N_14888,N_14901);
xnor UO_91 (O_91,N_14819,N_14920);
xor UO_92 (O_92,N_14800,N_14884);
nand UO_93 (O_93,N_14892,N_14822);
nor UO_94 (O_94,N_14943,N_14898);
and UO_95 (O_95,N_14869,N_14962);
xor UO_96 (O_96,N_14945,N_14919);
nor UO_97 (O_97,N_14921,N_14996);
or UO_98 (O_98,N_14809,N_14813);
or UO_99 (O_99,N_14977,N_14944);
nand UO_100 (O_100,N_14895,N_14953);
nor UO_101 (O_101,N_14972,N_14894);
or UO_102 (O_102,N_14928,N_14851);
xor UO_103 (O_103,N_14823,N_14849);
or UO_104 (O_104,N_14912,N_14988);
nand UO_105 (O_105,N_14992,N_14998);
nand UO_106 (O_106,N_14951,N_14817);
or UO_107 (O_107,N_14858,N_14979);
nand UO_108 (O_108,N_14924,N_14935);
nand UO_109 (O_109,N_14993,N_14875);
or UO_110 (O_110,N_14827,N_14976);
or UO_111 (O_111,N_14844,N_14961);
xnor UO_112 (O_112,N_14830,N_14812);
xor UO_113 (O_113,N_14857,N_14905);
nor UO_114 (O_114,N_14854,N_14870);
xnor UO_115 (O_115,N_14988,N_14871);
or UO_116 (O_116,N_14953,N_14932);
and UO_117 (O_117,N_14900,N_14923);
and UO_118 (O_118,N_14928,N_14995);
nor UO_119 (O_119,N_14910,N_14990);
nor UO_120 (O_120,N_14868,N_14903);
nor UO_121 (O_121,N_14924,N_14818);
or UO_122 (O_122,N_14829,N_14854);
nand UO_123 (O_123,N_14868,N_14827);
xnor UO_124 (O_124,N_14996,N_14935);
and UO_125 (O_125,N_14911,N_14996);
or UO_126 (O_126,N_14931,N_14939);
xor UO_127 (O_127,N_14821,N_14996);
and UO_128 (O_128,N_14958,N_14933);
and UO_129 (O_129,N_14954,N_14881);
nand UO_130 (O_130,N_14938,N_14952);
or UO_131 (O_131,N_14875,N_14991);
and UO_132 (O_132,N_14919,N_14992);
xnor UO_133 (O_133,N_14999,N_14895);
xnor UO_134 (O_134,N_14929,N_14920);
or UO_135 (O_135,N_14923,N_14913);
xnor UO_136 (O_136,N_14984,N_14868);
and UO_137 (O_137,N_14885,N_14811);
and UO_138 (O_138,N_14818,N_14829);
and UO_139 (O_139,N_14802,N_14867);
nand UO_140 (O_140,N_14877,N_14884);
xor UO_141 (O_141,N_14908,N_14944);
or UO_142 (O_142,N_14908,N_14884);
nor UO_143 (O_143,N_14847,N_14859);
nor UO_144 (O_144,N_14872,N_14932);
nor UO_145 (O_145,N_14982,N_14823);
or UO_146 (O_146,N_14928,N_14949);
or UO_147 (O_147,N_14991,N_14852);
nand UO_148 (O_148,N_14875,N_14816);
nor UO_149 (O_149,N_14983,N_14892);
nor UO_150 (O_150,N_14843,N_14845);
nand UO_151 (O_151,N_14868,N_14874);
xnor UO_152 (O_152,N_14912,N_14832);
and UO_153 (O_153,N_14893,N_14836);
and UO_154 (O_154,N_14816,N_14935);
nor UO_155 (O_155,N_14920,N_14925);
and UO_156 (O_156,N_14951,N_14934);
nand UO_157 (O_157,N_14818,N_14966);
nor UO_158 (O_158,N_14917,N_14997);
or UO_159 (O_159,N_14861,N_14868);
xor UO_160 (O_160,N_14890,N_14900);
nand UO_161 (O_161,N_14974,N_14882);
nand UO_162 (O_162,N_14995,N_14958);
and UO_163 (O_163,N_14800,N_14886);
nor UO_164 (O_164,N_14859,N_14945);
and UO_165 (O_165,N_14982,N_14839);
xnor UO_166 (O_166,N_14956,N_14889);
nor UO_167 (O_167,N_14806,N_14938);
nand UO_168 (O_168,N_14838,N_14867);
or UO_169 (O_169,N_14839,N_14976);
or UO_170 (O_170,N_14927,N_14821);
or UO_171 (O_171,N_14960,N_14874);
and UO_172 (O_172,N_14858,N_14827);
nand UO_173 (O_173,N_14811,N_14947);
and UO_174 (O_174,N_14839,N_14968);
or UO_175 (O_175,N_14992,N_14886);
and UO_176 (O_176,N_14828,N_14923);
xnor UO_177 (O_177,N_14838,N_14918);
and UO_178 (O_178,N_14925,N_14907);
and UO_179 (O_179,N_14902,N_14881);
xnor UO_180 (O_180,N_14928,N_14870);
and UO_181 (O_181,N_14930,N_14847);
nor UO_182 (O_182,N_14802,N_14862);
and UO_183 (O_183,N_14975,N_14843);
or UO_184 (O_184,N_14961,N_14929);
nand UO_185 (O_185,N_14955,N_14803);
nand UO_186 (O_186,N_14983,N_14860);
xor UO_187 (O_187,N_14826,N_14965);
nand UO_188 (O_188,N_14958,N_14978);
nand UO_189 (O_189,N_14888,N_14840);
nor UO_190 (O_190,N_14902,N_14981);
xor UO_191 (O_191,N_14808,N_14857);
or UO_192 (O_192,N_14848,N_14978);
xnor UO_193 (O_193,N_14846,N_14800);
nand UO_194 (O_194,N_14847,N_14822);
xnor UO_195 (O_195,N_14827,N_14918);
or UO_196 (O_196,N_14891,N_14836);
nand UO_197 (O_197,N_14870,N_14873);
and UO_198 (O_198,N_14849,N_14850);
nor UO_199 (O_199,N_14973,N_14882);
xor UO_200 (O_200,N_14807,N_14865);
xor UO_201 (O_201,N_14855,N_14865);
and UO_202 (O_202,N_14814,N_14823);
and UO_203 (O_203,N_14837,N_14991);
or UO_204 (O_204,N_14837,N_14881);
nand UO_205 (O_205,N_14806,N_14935);
nor UO_206 (O_206,N_14942,N_14992);
nand UO_207 (O_207,N_14830,N_14826);
or UO_208 (O_208,N_14940,N_14991);
and UO_209 (O_209,N_14948,N_14988);
nor UO_210 (O_210,N_14894,N_14993);
or UO_211 (O_211,N_14922,N_14950);
nand UO_212 (O_212,N_14978,N_14901);
nor UO_213 (O_213,N_14918,N_14996);
nor UO_214 (O_214,N_14911,N_14900);
xor UO_215 (O_215,N_14860,N_14840);
nand UO_216 (O_216,N_14871,N_14963);
xnor UO_217 (O_217,N_14977,N_14967);
nor UO_218 (O_218,N_14902,N_14946);
nor UO_219 (O_219,N_14846,N_14909);
nor UO_220 (O_220,N_14876,N_14841);
or UO_221 (O_221,N_14829,N_14937);
nand UO_222 (O_222,N_14859,N_14954);
nand UO_223 (O_223,N_14906,N_14971);
nand UO_224 (O_224,N_14959,N_14820);
xnor UO_225 (O_225,N_14916,N_14837);
or UO_226 (O_226,N_14999,N_14978);
xnor UO_227 (O_227,N_14811,N_14945);
or UO_228 (O_228,N_14815,N_14898);
nor UO_229 (O_229,N_14977,N_14978);
and UO_230 (O_230,N_14909,N_14934);
or UO_231 (O_231,N_14830,N_14800);
and UO_232 (O_232,N_14847,N_14835);
xnor UO_233 (O_233,N_14944,N_14954);
nand UO_234 (O_234,N_14887,N_14865);
nand UO_235 (O_235,N_14825,N_14950);
nor UO_236 (O_236,N_14946,N_14846);
and UO_237 (O_237,N_14934,N_14912);
or UO_238 (O_238,N_14925,N_14984);
and UO_239 (O_239,N_14945,N_14926);
and UO_240 (O_240,N_14994,N_14836);
xor UO_241 (O_241,N_14922,N_14877);
xor UO_242 (O_242,N_14890,N_14946);
nand UO_243 (O_243,N_14883,N_14843);
or UO_244 (O_244,N_14986,N_14939);
nand UO_245 (O_245,N_14928,N_14828);
or UO_246 (O_246,N_14956,N_14891);
and UO_247 (O_247,N_14830,N_14882);
and UO_248 (O_248,N_14923,N_14979);
nor UO_249 (O_249,N_14893,N_14813);
nor UO_250 (O_250,N_14867,N_14928);
xnor UO_251 (O_251,N_14800,N_14858);
and UO_252 (O_252,N_14815,N_14877);
or UO_253 (O_253,N_14920,N_14885);
and UO_254 (O_254,N_14957,N_14893);
or UO_255 (O_255,N_14983,N_14820);
nand UO_256 (O_256,N_14882,N_14992);
nor UO_257 (O_257,N_14847,N_14885);
or UO_258 (O_258,N_14837,N_14867);
or UO_259 (O_259,N_14803,N_14992);
and UO_260 (O_260,N_14970,N_14823);
nand UO_261 (O_261,N_14977,N_14997);
and UO_262 (O_262,N_14984,N_14942);
or UO_263 (O_263,N_14993,N_14814);
nand UO_264 (O_264,N_14905,N_14819);
and UO_265 (O_265,N_14895,N_14851);
and UO_266 (O_266,N_14842,N_14892);
and UO_267 (O_267,N_14816,N_14872);
and UO_268 (O_268,N_14839,N_14820);
or UO_269 (O_269,N_14986,N_14942);
nand UO_270 (O_270,N_14893,N_14844);
nor UO_271 (O_271,N_14976,N_14841);
or UO_272 (O_272,N_14859,N_14810);
nor UO_273 (O_273,N_14933,N_14846);
or UO_274 (O_274,N_14972,N_14928);
or UO_275 (O_275,N_14850,N_14919);
or UO_276 (O_276,N_14802,N_14820);
xnor UO_277 (O_277,N_14887,N_14974);
xor UO_278 (O_278,N_14925,N_14994);
nand UO_279 (O_279,N_14804,N_14961);
xor UO_280 (O_280,N_14992,N_14916);
nor UO_281 (O_281,N_14878,N_14930);
or UO_282 (O_282,N_14839,N_14800);
nor UO_283 (O_283,N_14800,N_14892);
nor UO_284 (O_284,N_14938,N_14853);
nor UO_285 (O_285,N_14961,N_14805);
or UO_286 (O_286,N_14958,N_14923);
nor UO_287 (O_287,N_14954,N_14965);
or UO_288 (O_288,N_14858,N_14801);
nor UO_289 (O_289,N_14936,N_14855);
or UO_290 (O_290,N_14877,N_14887);
nor UO_291 (O_291,N_14989,N_14838);
or UO_292 (O_292,N_14973,N_14812);
nor UO_293 (O_293,N_14891,N_14823);
nor UO_294 (O_294,N_14899,N_14872);
nor UO_295 (O_295,N_14885,N_14846);
xor UO_296 (O_296,N_14805,N_14806);
nand UO_297 (O_297,N_14982,N_14998);
or UO_298 (O_298,N_14914,N_14845);
nor UO_299 (O_299,N_14803,N_14846);
xnor UO_300 (O_300,N_14915,N_14912);
or UO_301 (O_301,N_14879,N_14808);
xor UO_302 (O_302,N_14828,N_14892);
or UO_303 (O_303,N_14906,N_14877);
and UO_304 (O_304,N_14966,N_14981);
and UO_305 (O_305,N_14995,N_14863);
or UO_306 (O_306,N_14839,N_14905);
or UO_307 (O_307,N_14890,N_14869);
nor UO_308 (O_308,N_14983,N_14895);
xor UO_309 (O_309,N_14837,N_14983);
and UO_310 (O_310,N_14932,N_14907);
nand UO_311 (O_311,N_14838,N_14903);
nand UO_312 (O_312,N_14904,N_14804);
nand UO_313 (O_313,N_14823,N_14919);
xnor UO_314 (O_314,N_14822,N_14845);
or UO_315 (O_315,N_14814,N_14916);
xor UO_316 (O_316,N_14915,N_14969);
xor UO_317 (O_317,N_14840,N_14930);
xnor UO_318 (O_318,N_14926,N_14962);
or UO_319 (O_319,N_14905,N_14853);
xnor UO_320 (O_320,N_14816,N_14979);
and UO_321 (O_321,N_14838,N_14911);
nand UO_322 (O_322,N_14813,N_14815);
nand UO_323 (O_323,N_14833,N_14913);
xor UO_324 (O_324,N_14856,N_14990);
xor UO_325 (O_325,N_14944,N_14803);
xnor UO_326 (O_326,N_14890,N_14895);
nand UO_327 (O_327,N_14890,N_14876);
xor UO_328 (O_328,N_14831,N_14908);
and UO_329 (O_329,N_14992,N_14876);
xnor UO_330 (O_330,N_14831,N_14998);
nand UO_331 (O_331,N_14850,N_14827);
nor UO_332 (O_332,N_14985,N_14910);
and UO_333 (O_333,N_14846,N_14980);
nor UO_334 (O_334,N_14990,N_14934);
xnor UO_335 (O_335,N_14846,N_14932);
or UO_336 (O_336,N_14854,N_14819);
nand UO_337 (O_337,N_14934,N_14991);
xnor UO_338 (O_338,N_14916,N_14835);
xnor UO_339 (O_339,N_14874,N_14824);
and UO_340 (O_340,N_14865,N_14905);
nand UO_341 (O_341,N_14801,N_14820);
nor UO_342 (O_342,N_14945,N_14958);
nand UO_343 (O_343,N_14995,N_14809);
or UO_344 (O_344,N_14963,N_14998);
and UO_345 (O_345,N_14806,N_14941);
xnor UO_346 (O_346,N_14801,N_14825);
nand UO_347 (O_347,N_14916,N_14924);
and UO_348 (O_348,N_14878,N_14919);
and UO_349 (O_349,N_14891,N_14847);
xnor UO_350 (O_350,N_14808,N_14924);
xnor UO_351 (O_351,N_14951,N_14967);
nor UO_352 (O_352,N_14823,N_14934);
and UO_353 (O_353,N_14975,N_14959);
nand UO_354 (O_354,N_14877,N_14988);
nand UO_355 (O_355,N_14996,N_14992);
nor UO_356 (O_356,N_14866,N_14855);
and UO_357 (O_357,N_14950,N_14965);
or UO_358 (O_358,N_14974,N_14895);
and UO_359 (O_359,N_14915,N_14853);
and UO_360 (O_360,N_14845,N_14919);
nand UO_361 (O_361,N_14874,N_14930);
or UO_362 (O_362,N_14886,N_14909);
or UO_363 (O_363,N_14805,N_14800);
xor UO_364 (O_364,N_14918,N_14948);
nor UO_365 (O_365,N_14870,N_14828);
and UO_366 (O_366,N_14883,N_14990);
or UO_367 (O_367,N_14994,N_14977);
and UO_368 (O_368,N_14926,N_14912);
xor UO_369 (O_369,N_14859,N_14906);
nand UO_370 (O_370,N_14853,N_14801);
and UO_371 (O_371,N_14888,N_14827);
xnor UO_372 (O_372,N_14831,N_14917);
xor UO_373 (O_373,N_14894,N_14836);
or UO_374 (O_374,N_14960,N_14908);
or UO_375 (O_375,N_14931,N_14987);
xor UO_376 (O_376,N_14818,N_14891);
and UO_377 (O_377,N_14820,N_14886);
xnor UO_378 (O_378,N_14896,N_14898);
and UO_379 (O_379,N_14884,N_14913);
xnor UO_380 (O_380,N_14838,N_14815);
and UO_381 (O_381,N_14854,N_14983);
or UO_382 (O_382,N_14975,N_14916);
nand UO_383 (O_383,N_14865,N_14860);
nand UO_384 (O_384,N_14824,N_14888);
and UO_385 (O_385,N_14800,N_14989);
and UO_386 (O_386,N_14819,N_14850);
nand UO_387 (O_387,N_14902,N_14968);
or UO_388 (O_388,N_14939,N_14858);
or UO_389 (O_389,N_14970,N_14829);
and UO_390 (O_390,N_14815,N_14953);
nand UO_391 (O_391,N_14937,N_14919);
nor UO_392 (O_392,N_14903,N_14946);
or UO_393 (O_393,N_14992,N_14850);
xnor UO_394 (O_394,N_14944,N_14901);
or UO_395 (O_395,N_14804,N_14937);
nand UO_396 (O_396,N_14959,N_14870);
nand UO_397 (O_397,N_14842,N_14943);
nand UO_398 (O_398,N_14899,N_14997);
nand UO_399 (O_399,N_14926,N_14815);
and UO_400 (O_400,N_14942,N_14853);
nor UO_401 (O_401,N_14826,N_14957);
or UO_402 (O_402,N_14951,N_14877);
and UO_403 (O_403,N_14965,N_14917);
or UO_404 (O_404,N_14983,N_14842);
nor UO_405 (O_405,N_14867,N_14861);
xor UO_406 (O_406,N_14861,N_14966);
nor UO_407 (O_407,N_14955,N_14929);
or UO_408 (O_408,N_14858,N_14812);
and UO_409 (O_409,N_14970,N_14804);
and UO_410 (O_410,N_14911,N_14971);
xor UO_411 (O_411,N_14839,N_14985);
or UO_412 (O_412,N_14968,N_14899);
or UO_413 (O_413,N_14825,N_14959);
nand UO_414 (O_414,N_14980,N_14822);
xor UO_415 (O_415,N_14973,N_14907);
or UO_416 (O_416,N_14913,N_14880);
nor UO_417 (O_417,N_14997,N_14853);
and UO_418 (O_418,N_14811,N_14955);
xnor UO_419 (O_419,N_14879,N_14924);
and UO_420 (O_420,N_14805,N_14850);
and UO_421 (O_421,N_14806,N_14888);
nor UO_422 (O_422,N_14995,N_14906);
or UO_423 (O_423,N_14909,N_14853);
xor UO_424 (O_424,N_14932,N_14971);
or UO_425 (O_425,N_14962,N_14808);
xor UO_426 (O_426,N_14882,N_14934);
or UO_427 (O_427,N_14861,N_14841);
and UO_428 (O_428,N_14979,N_14856);
nand UO_429 (O_429,N_14995,N_14952);
nor UO_430 (O_430,N_14853,N_14831);
nand UO_431 (O_431,N_14966,N_14934);
or UO_432 (O_432,N_14929,N_14932);
nand UO_433 (O_433,N_14869,N_14937);
and UO_434 (O_434,N_14955,N_14890);
nor UO_435 (O_435,N_14954,N_14952);
nor UO_436 (O_436,N_14921,N_14979);
nor UO_437 (O_437,N_14976,N_14851);
xor UO_438 (O_438,N_14971,N_14997);
xor UO_439 (O_439,N_14997,N_14849);
or UO_440 (O_440,N_14892,N_14871);
or UO_441 (O_441,N_14825,N_14821);
xnor UO_442 (O_442,N_14948,N_14855);
and UO_443 (O_443,N_14924,N_14862);
nand UO_444 (O_444,N_14831,N_14897);
xor UO_445 (O_445,N_14974,N_14975);
and UO_446 (O_446,N_14891,N_14802);
xnor UO_447 (O_447,N_14852,N_14922);
or UO_448 (O_448,N_14997,N_14861);
or UO_449 (O_449,N_14927,N_14904);
nand UO_450 (O_450,N_14929,N_14826);
or UO_451 (O_451,N_14957,N_14962);
and UO_452 (O_452,N_14864,N_14885);
and UO_453 (O_453,N_14858,N_14853);
xnor UO_454 (O_454,N_14818,N_14893);
xnor UO_455 (O_455,N_14966,N_14983);
and UO_456 (O_456,N_14865,N_14852);
nor UO_457 (O_457,N_14996,N_14891);
xor UO_458 (O_458,N_14870,N_14979);
nor UO_459 (O_459,N_14844,N_14831);
nand UO_460 (O_460,N_14836,N_14882);
or UO_461 (O_461,N_14993,N_14800);
xor UO_462 (O_462,N_14809,N_14979);
or UO_463 (O_463,N_14976,N_14804);
or UO_464 (O_464,N_14827,N_14942);
xor UO_465 (O_465,N_14823,N_14842);
nor UO_466 (O_466,N_14961,N_14870);
nor UO_467 (O_467,N_14846,N_14870);
nor UO_468 (O_468,N_14953,N_14899);
xor UO_469 (O_469,N_14815,N_14809);
xor UO_470 (O_470,N_14963,N_14959);
nor UO_471 (O_471,N_14889,N_14848);
or UO_472 (O_472,N_14854,N_14996);
and UO_473 (O_473,N_14957,N_14853);
xor UO_474 (O_474,N_14993,N_14911);
nor UO_475 (O_475,N_14874,N_14985);
nand UO_476 (O_476,N_14908,N_14999);
xnor UO_477 (O_477,N_14957,N_14970);
and UO_478 (O_478,N_14988,N_14850);
xor UO_479 (O_479,N_14909,N_14900);
or UO_480 (O_480,N_14803,N_14972);
nor UO_481 (O_481,N_14903,N_14921);
and UO_482 (O_482,N_14959,N_14856);
nor UO_483 (O_483,N_14877,N_14942);
nor UO_484 (O_484,N_14950,N_14839);
or UO_485 (O_485,N_14925,N_14995);
nand UO_486 (O_486,N_14986,N_14901);
xor UO_487 (O_487,N_14826,N_14859);
and UO_488 (O_488,N_14961,N_14996);
nor UO_489 (O_489,N_14847,N_14998);
and UO_490 (O_490,N_14968,N_14980);
or UO_491 (O_491,N_14961,N_14901);
xnor UO_492 (O_492,N_14997,N_14996);
or UO_493 (O_493,N_14812,N_14806);
nand UO_494 (O_494,N_14828,N_14949);
or UO_495 (O_495,N_14979,N_14826);
and UO_496 (O_496,N_14915,N_14893);
nand UO_497 (O_497,N_14800,N_14986);
nand UO_498 (O_498,N_14811,N_14867);
xor UO_499 (O_499,N_14982,N_14898);
xor UO_500 (O_500,N_14838,N_14958);
and UO_501 (O_501,N_14818,N_14861);
nor UO_502 (O_502,N_14805,N_14819);
nand UO_503 (O_503,N_14913,N_14981);
nand UO_504 (O_504,N_14946,N_14844);
nand UO_505 (O_505,N_14952,N_14858);
xnor UO_506 (O_506,N_14883,N_14851);
and UO_507 (O_507,N_14859,N_14853);
xnor UO_508 (O_508,N_14863,N_14958);
or UO_509 (O_509,N_14875,N_14855);
nand UO_510 (O_510,N_14932,N_14813);
and UO_511 (O_511,N_14966,N_14961);
nand UO_512 (O_512,N_14947,N_14916);
nand UO_513 (O_513,N_14954,N_14822);
xor UO_514 (O_514,N_14835,N_14959);
or UO_515 (O_515,N_14943,N_14942);
nor UO_516 (O_516,N_14993,N_14886);
nand UO_517 (O_517,N_14809,N_14927);
nand UO_518 (O_518,N_14870,N_14888);
nor UO_519 (O_519,N_14999,N_14871);
nor UO_520 (O_520,N_14883,N_14900);
xnor UO_521 (O_521,N_14815,N_14925);
or UO_522 (O_522,N_14801,N_14864);
xnor UO_523 (O_523,N_14959,N_14922);
xor UO_524 (O_524,N_14912,N_14846);
and UO_525 (O_525,N_14941,N_14814);
nand UO_526 (O_526,N_14915,N_14845);
and UO_527 (O_527,N_14950,N_14975);
nand UO_528 (O_528,N_14976,N_14960);
nand UO_529 (O_529,N_14888,N_14936);
or UO_530 (O_530,N_14949,N_14863);
and UO_531 (O_531,N_14893,N_14816);
or UO_532 (O_532,N_14894,N_14949);
or UO_533 (O_533,N_14874,N_14869);
or UO_534 (O_534,N_14942,N_14896);
nor UO_535 (O_535,N_14834,N_14981);
or UO_536 (O_536,N_14891,N_14984);
and UO_537 (O_537,N_14853,N_14889);
or UO_538 (O_538,N_14882,N_14869);
nand UO_539 (O_539,N_14952,N_14991);
and UO_540 (O_540,N_14838,N_14847);
or UO_541 (O_541,N_14882,N_14903);
xnor UO_542 (O_542,N_14925,N_14833);
or UO_543 (O_543,N_14965,N_14874);
xor UO_544 (O_544,N_14967,N_14913);
nor UO_545 (O_545,N_14929,N_14962);
and UO_546 (O_546,N_14853,N_14982);
xnor UO_547 (O_547,N_14916,N_14900);
or UO_548 (O_548,N_14878,N_14957);
xor UO_549 (O_549,N_14816,N_14817);
or UO_550 (O_550,N_14931,N_14899);
nand UO_551 (O_551,N_14926,N_14896);
nand UO_552 (O_552,N_14979,N_14949);
nor UO_553 (O_553,N_14806,N_14881);
or UO_554 (O_554,N_14889,N_14986);
nand UO_555 (O_555,N_14817,N_14966);
or UO_556 (O_556,N_14811,N_14822);
nor UO_557 (O_557,N_14999,N_14801);
or UO_558 (O_558,N_14835,N_14911);
nor UO_559 (O_559,N_14958,N_14824);
or UO_560 (O_560,N_14805,N_14857);
nand UO_561 (O_561,N_14883,N_14853);
and UO_562 (O_562,N_14917,N_14991);
xor UO_563 (O_563,N_14878,N_14966);
and UO_564 (O_564,N_14991,N_14808);
nor UO_565 (O_565,N_14824,N_14961);
xor UO_566 (O_566,N_14948,N_14835);
nor UO_567 (O_567,N_14823,N_14840);
nor UO_568 (O_568,N_14872,N_14841);
nor UO_569 (O_569,N_14887,N_14932);
nor UO_570 (O_570,N_14970,N_14949);
nor UO_571 (O_571,N_14821,N_14961);
xor UO_572 (O_572,N_14941,N_14961);
nand UO_573 (O_573,N_14862,N_14909);
xnor UO_574 (O_574,N_14932,N_14883);
nor UO_575 (O_575,N_14896,N_14950);
or UO_576 (O_576,N_14957,N_14816);
or UO_577 (O_577,N_14804,N_14800);
or UO_578 (O_578,N_14824,N_14833);
nor UO_579 (O_579,N_14851,N_14896);
nand UO_580 (O_580,N_14991,N_14933);
xor UO_581 (O_581,N_14816,N_14894);
and UO_582 (O_582,N_14803,N_14948);
and UO_583 (O_583,N_14852,N_14879);
nor UO_584 (O_584,N_14857,N_14984);
and UO_585 (O_585,N_14872,N_14854);
xnor UO_586 (O_586,N_14804,N_14899);
xnor UO_587 (O_587,N_14804,N_14811);
nor UO_588 (O_588,N_14853,N_14861);
and UO_589 (O_589,N_14876,N_14935);
nor UO_590 (O_590,N_14924,N_14871);
and UO_591 (O_591,N_14875,N_14920);
or UO_592 (O_592,N_14969,N_14997);
xor UO_593 (O_593,N_14981,N_14876);
or UO_594 (O_594,N_14827,N_14807);
nand UO_595 (O_595,N_14917,N_14989);
xor UO_596 (O_596,N_14852,N_14968);
nand UO_597 (O_597,N_14943,N_14968);
nand UO_598 (O_598,N_14889,N_14878);
and UO_599 (O_599,N_14989,N_14995);
nor UO_600 (O_600,N_14969,N_14829);
or UO_601 (O_601,N_14846,N_14830);
nand UO_602 (O_602,N_14984,N_14804);
nand UO_603 (O_603,N_14967,N_14829);
or UO_604 (O_604,N_14874,N_14914);
nand UO_605 (O_605,N_14835,N_14832);
nor UO_606 (O_606,N_14870,N_14949);
or UO_607 (O_607,N_14861,N_14973);
nand UO_608 (O_608,N_14935,N_14846);
nand UO_609 (O_609,N_14944,N_14815);
nor UO_610 (O_610,N_14984,N_14803);
nor UO_611 (O_611,N_14916,N_14803);
xnor UO_612 (O_612,N_14913,N_14803);
nand UO_613 (O_613,N_14929,N_14956);
and UO_614 (O_614,N_14834,N_14996);
nand UO_615 (O_615,N_14841,N_14987);
nor UO_616 (O_616,N_14949,N_14803);
nand UO_617 (O_617,N_14809,N_14992);
nor UO_618 (O_618,N_14935,N_14933);
nand UO_619 (O_619,N_14951,N_14914);
nor UO_620 (O_620,N_14839,N_14904);
or UO_621 (O_621,N_14957,N_14871);
and UO_622 (O_622,N_14907,N_14852);
nand UO_623 (O_623,N_14821,N_14905);
or UO_624 (O_624,N_14866,N_14899);
or UO_625 (O_625,N_14812,N_14998);
or UO_626 (O_626,N_14961,N_14867);
xnor UO_627 (O_627,N_14869,N_14833);
xor UO_628 (O_628,N_14816,N_14986);
and UO_629 (O_629,N_14922,N_14988);
and UO_630 (O_630,N_14976,N_14830);
xor UO_631 (O_631,N_14867,N_14862);
nor UO_632 (O_632,N_14998,N_14918);
nand UO_633 (O_633,N_14978,N_14802);
nor UO_634 (O_634,N_14810,N_14998);
nand UO_635 (O_635,N_14835,N_14840);
nor UO_636 (O_636,N_14956,N_14878);
and UO_637 (O_637,N_14963,N_14878);
nor UO_638 (O_638,N_14999,N_14884);
nand UO_639 (O_639,N_14846,N_14896);
xnor UO_640 (O_640,N_14820,N_14827);
and UO_641 (O_641,N_14801,N_14878);
nand UO_642 (O_642,N_14834,N_14912);
or UO_643 (O_643,N_14924,N_14931);
or UO_644 (O_644,N_14836,N_14878);
xor UO_645 (O_645,N_14935,N_14815);
nand UO_646 (O_646,N_14923,N_14976);
nor UO_647 (O_647,N_14812,N_14924);
nand UO_648 (O_648,N_14954,N_14873);
xor UO_649 (O_649,N_14925,N_14914);
and UO_650 (O_650,N_14991,N_14872);
nor UO_651 (O_651,N_14913,N_14808);
xor UO_652 (O_652,N_14879,N_14986);
xnor UO_653 (O_653,N_14873,N_14970);
or UO_654 (O_654,N_14920,N_14854);
nor UO_655 (O_655,N_14948,N_14916);
nand UO_656 (O_656,N_14827,N_14871);
nand UO_657 (O_657,N_14925,N_14817);
xnor UO_658 (O_658,N_14828,N_14887);
and UO_659 (O_659,N_14932,N_14961);
and UO_660 (O_660,N_14957,N_14989);
or UO_661 (O_661,N_14946,N_14979);
xnor UO_662 (O_662,N_14842,N_14820);
xnor UO_663 (O_663,N_14916,N_14849);
or UO_664 (O_664,N_14932,N_14912);
nand UO_665 (O_665,N_14900,N_14939);
and UO_666 (O_666,N_14915,N_14850);
xor UO_667 (O_667,N_14876,N_14968);
or UO_668 (O_668,N_14875,N_14927);
xor UO_669 (O_669,N_14831,N_14895);
xor UO_670 (O_670,N_14828,N_14994);
and UO_671 (O_671,N_14952,N_14972);
or UO_672 (O_672,N_14854,N_14977);
or UO_673 (O_673,N_14939,N_14860);
or UO_674 (O_674,N_14891,N_14875);
nor UO_675 (O_675,N_14947,N_14929);
and UO_676 (O_676,N_14821,N_14822);
nor UO_677 (O_677,N_14998,N_14965);
nand UO_678 (O_678,N_14976,N_14983);
or UO_679 (O_679,N_14834,N_14939);
nand UO_680 (O_680,N_14923,N_14831);
and UO_681 (O_681,N_14805,N_14925);
nor UO_682 (O_682,N_14967,N_14883);
nor UO_683 (O_683,N_14983,N_14864);
nor UO_684 (O_684,N_14879,N_14891);
xnor UO_685 (O_685,N_14806,N_14845);
nand UO_686 (O_686,N_14903,N_14937);
xor UO_687 (O_687,N_14897,N_14915);
and UO_688 (O_688,N_14814,N_14853);
nor UO_689 (O_689,N_14808,N_14946);
or UO_690 (O_690,N_14999,N_14833);
nor UO_691 (O_691,N_14833,N_14903);
or UO_692 (O_692,N_14967,N_14852);
xor UO_693 (O_693,N_14965,N_14825);
or UO_694 (O_694,N_14908,N_14835);
or UO_695 (O_695,N_14856,N_14828);
xnor UO_696 (O_696,N_14830,N_14873);
nand UO_697 (O_697,N_14802,N_14921);
or UO_698 (O_698,N_14880,N_14847);
xor UO_699 (O_699,N_14908,N_14851);
nand UO_700 (O_700,N_14869,N_14812);
and UO_701 (O_701,N_14976,N_14967);
xnor UO_702 (O_702,N_14977,N_14894);
xnor UO_703 (O_703,N_14884,N_14803);
nor UO_704 (O_704,N_14982,N_14840);
nor UO_705 (O_705,N_14987,N_14944);
nand UO_706 (O_706,N_14919,N_14811);
nand UO_707 (O_707,N_14998,N_14894);
nand UO_708 (O_708,N_14831,N_14852);
or UO_709 (O_709,N_14948,N_14992);
nor UO_710 (O_710,N_14932,N_14834);
and UO_711 (O_711,N_14938,N_14971);
xnor UO_712 (O_712,N_14815,N_14835);
xnor UO_713 (O_713,N_14926,N_14809);
nand UO_714 (O_714,N_14827,N_14971);
and UO_715 (O_715,N_14944,N_14899);
and UO_716 (O_716,N_14823,N_14800);
xor UO_717 (O_717,N_14878,N_14896);
nand UO_718 (O_718,N_14800,N_14983);
xor UO_719 (O_719,N_14989,N_14915);
nand UO_720 (O_720,N_14801,N_14852);
nor UO_721 (O_721,N_14971,N_14936);
nand UO_722 (O_722,N_14894,N_14805);
nor UO_723 (O_723,N_14917,N_14885);
nor UO_724 (O_724,N_14940,N_14981);
xor UO_725 (O_725,N_14947,N_14936);
nand UO_726 (O_726,N_14827,N_14815);
or UO_727 (O_727,N_14952,N_14967);
or UO_728 (O_728,N_14898,N_14916);
or UO_729 (O_729,N_14866,N_14994);
nand UO_730 (O_730,N_14886,N_14831);
xnor UO_731 (O_731,N_14850,N_14998);
xor UO_732 (O_732,N_14863,N_14860);
nand UO_733 (O_733,N_14819,N_14941);
and UO_734 (O_734,N_14920,N_14802);
xor UO_735 (O_735,N_14978,N_14864);
nand UO_736 (O_736,N_14914,N_14908);
and UO_737 (O_737,N_14849,N_14881);
or UO_738 (O_738,N_14813,N_14851);
and UO_739 (O_739,N_14895,N_14807);
and UO_740 (O_740,N_14959,N_14876);
and UO_741 (O_741,N_14838,N_14816);
or UO_742 (O_742,N_14860,N_14806);
nor UO_743 (O_743,N_14989,N_14865);
or UO_744 (O_744,N_14818,N_14949);
nor UO_745 (O_745,N_14878,N_14841);
and UO_746 (O_746,N_14867,N_14934);
and UO_747 (O_747,N_14868,N_14853);
and UO_748 (O_748,N_14801,N_14842);
and UO_749 (O_749,N_14854,N_14963);
nand UO_750 (O_750,N_14962,N_14995);
nor UO_751 (O_751,N_14852,N_14926);
xnor UO_752 (O_752,N_14971,N_14809);
nor UO_753 (O_753,N_14886,N_14915);
nand UO_754 (O_754,N_14842,N_14864);
xor UO_755 (O_755,N_14876,N_14972);
nor UO_756 (O_756,N_14929,N_14814);
and UO_757 (O_757,N_14889,N_14850);
and UO_758 (O_758,N_14993,N_14842);
xnor UO_759 (O_759,N_14880,N_14832);
xor UO_760 (O_760,N_14803,N_14817);
xnor UO_761 (O_761,N_14996,N_14835);
and UO_762 (O_762,N_14859,N_14809);
nand UO_763 (O_763,N_14876,N_14914);
nand UO_764 (O_764,N_14968,N_14924);
xor UO_765 (O_765,N_14955,N_14938);
nand UO_766 (O_766,N_14803,N_14882);
xor UO_767 (O_767,N_14870,N_14915);
nand UO_768 (O_768,N_14954,N_14956);
nand UO_769 (O_769,N_14822,N_14879);
xor UO_770 (O_770,N_14815,N_14995);
nand UO_771 (O_771,N_14934,N_14822);
and UO_772 (O_772,N_14990,N_14920);
nor UO_773 (O_773,N_14977,N_14835);
nand UO_774 (O_774,N_14933,N_14845);
nor UO_775 (O_775,N_14979,N_14892);
and UO_776 (O_776,N_14810,N_14857);
xnor UO_777 (O_777,N_14981,N_14889);
or UO_778 (O_778,N_14878,N_14989);
or UO_779 (O_779,N_14997,N_14870);
nor UO_780 (O_780,N_14885,N_14982);
or UO_781 (O_781,N_14856,N_14934);
nand UO_782 (O_782,N_14853,N_14816);
nand UO_783 (O_783,N_14824,N_14814);
xor UO_784 (O_784,N_14930,N_14801);
and UO_785 (O_785,N_14950,N_14917);
nor UO_786 (O_786,N_14873,N_14883);
and UO_787 (O_787,N_14915,N_14843);
or UO_788 (O_788,N_14820,N_14877);
and UO_789 (O_789,N_14916,N_14821);
xor UO_790 (O_790,N_14961,N_14911);
nor UO_791 (O_791,N_14851,N_14872);
nand UO_792 (O_792,N_14966,N_14913);
xor UO_793 (O_793,N_14961,N_14907);
nor UO_794 (O_794,N_14803,N_14847);
nand UO_795 (O_795,N_14817,N_14894);
or UO_796 (O_796,N_14889,N_14910);
and UO_797 (O_797,N_14963,N_14897);
xnor UO_798 (O_798,N_14862,N_14818);
or UO_799 (O_799,N_14879,N_14856);
or UO_800 (O_800,N_14876,N_14975);
and UO_801 (O_801,N_14994,N_14872);
or UO_802 (O_802,N_14905,N_14872);
xor UO_803 (O_803,N_14978,N_14860);
nor UO_804 (O_804,N_14813,N_14822);
nand UO_805 (O_805,N_14807,N_14916);
or UO_806 (O_806,N_14908,N_14956);
nor UO_807 (O_807,N_14801,N_14834);
and UO_808 (O_808,N_14921,N_14868);
and UO_809 (O_809,N_14945,N_14928);
nand UO_810 (O_810,N_14977,N_14892);
nor UO_811 (O_811,N_14845,N_14942);
nand UO_812 (O_812,N_14904,N_14949);
or UO_813 (O_813,N_14886,N_14876);
or UO_814 (O_814,N_14969,N_14937);
and UO_815 (O_815,N_14986,N_14963);
and UO_816 (O_816,N_14953,N_14896);
and UO_817 (O_817,N_14929,N_14893);
nand UO_818 (O_818,N_14864,N_14918);
xor UO_819 (O_819,N_14817,N_14933);
nand UO_820 (O_820,N_14959,N_14838);
nand UO_821 (O_821,N_14818,N_14805);
and UO_822 (O_822,N_14963,N_14869);
nor UO_823 (O_823,N_14809,N_14864);
nor UO_824 (O_824,N_14979,N_14908);
nand UO_825 (O_825,N_14913,N_14995);
xnor UO_826 (O_826,N_14838,N_14915);
or UO_827 (O_827,N_14818,N_14904);
xnor UO_828 (O_828,N_14808,N_14998);
and UO_829 (O_829,N_14916,N_14995);
and UO_830 (O_830,N_14816,N_14832);
nor UO_831 (O_831,N_14902,N_14844);
xor UO_832 (O_832,N_14979,N_14975);
and UO_833 (O_833,N_14955,N_14854);
nand UO_834 (O_834,N_14832,N_14985);
and UO_835 (O_835,N_14838,N_14820);
xor UO_836 (O_836,N_14828,N_14829);
or UO_837 (O_837,N_14931,N_14912);
nand UO_838 (O_838,N_14834,N_14904);
xor UO_839 (O_839,N_14942,N_14901);
nor UO_840 (O_840,N_14844,N_14826);
xnor UO_841 (O_841,N_14876,N_14896);
nand UO_842 (O_842,N_14960,N_14948);
or UO_843 (O_843,N_14966,N_14843);
nor UO_844 (O_844,N_14997,N_14856);
nand UO_845 (O_845,N_14909,N_14929);
nand UO_846 (O_846,N_14909,N_14893);
nor UO_847 (O_847,N_14983,N_14819);
nand UO_848 (O_848,N_14916,N_14810);
and UO_849 (O_849,N_14993,N_14941);
and UO_850 (O_850,N_14822,N_14855);
or UO_851 (O_851,N_14891,N_14892);
and UO_852 (O_852,N_14941,N_14944);
or UO_853 (O_853,N_14816,N_14882);
xor UO_854 (O_854,N_14858,N_14891);
xor UO_855 (O_855,N_14887,N_14986);
xnor UO_856 (O_856,N_14908,N_14904);
xnor UO_857 (O_857,N_14857,N_14978);
nand UO_858 (O_858,N_14814,N_14838);
xnor UO_859 (O_859,N_14917,N_14888);
and UO_860 (O_860,N_14802,N_14883);
and UO_861 (O_861,N_14999,N_14841);
nand UO_862 (O_862,N_14846,N_14983);
nor UO_863 (O_863,N_14831,N_14994);
nor UO_864 (O_864,N_14995,N_14849);
nor UO_865 (O_865,N_14921,N_14905);
xor UO_866 (O_866,N_14951,N_14920);
nor UO_867 (O_867,N_14815,N_14929);
xor UO_868 (O_868,N_14968,N_14811);
nand UO_869 (O_869,N_14878,N_14904);
nor UO_870 (O_870,N_14829,N_14954);
nor UO_871 (O_871,N_14900,N_14838);
or UO_872 (O_872,N_14945,N_14942);
nor UO_873 (O_873,N_14816,N_14925);
xor UO_874 (O_874,N_14871,N_14816);
xnor UO_875 (O_875,N_14957,N_14886);
and UO_876 (O_876,N_14990,N_14804);
xor UO_877 (O_877,N_14879,N_14825);
nand UO_878 (O_878,N_14901,N_14891);
or UO_879 (O_879,N_14962,N_14890);
and UO_880 (O_880,N_14979,N_14959);
nand UO_881 (O_881,N_14927,N_14978);
nand UO_882 (O_882,N_14924,N_14914);
nor UO_883 (O_883,N_14928,N_14868);
and UO_884 (O_884,N_14834,N_14818);
and UO_885 (O_885,N_14970,N_14986);
xor UO_886 (O_886,N_14837,N_14967);
nand UO_887 (O_887,N_14977,N_14941);
xnor UO_888 (O_888,N_14826,N_14918);
or UO_889 (O_889,N_14896,N_14828);
nand UO_890 (O_890,N_14840,N_14868);
nand UO_891 (O_891,N_14995,N_14823);
nor UO_892 (O_892,N_14800,N_14894);
nor UO_893 (O_893,N_14948,N_14903);
or UO_894 (O_894,N_14808,N_14863);
nor UO_895 (O_895,N_14932,N_14829);
nor UO_896 (O_896,N_14972,N_14932);
xor UO_897 (O_897,N_14957,N_14828);
xnor UO_898 (O_898,N_14863,N_14903);
or UO_899 (O_899,N_14924,N_14870);
and UO_900 (O_900,N_14912,N_14805);
or UO_901 (O_901,N_14887,N_14924);
nand UO_902 (O_902,N_14804,N_14889);
nor UO_903 (O_903,N_14877,N_14819);
xor UO_904 (O_904,N_14830,N_14813);
xnor UO_905 (O_905,N_14976,N_14896);
or UO_906 (O_906,N_14905,N_14900);
xnor UO_907 (O_907,N_14866,N_14901);
xor UO_908 (O_908,N_14951,N_14873);
or UO_909 (O_909,N_14997,N_14932);
nor UO_910 (O_910,N_14965,N_14860);
or UO_911 (O_911,N_14912,N_14856);
nand UO_912 (O_912,N_14810,N_14965);
xnor UO_913 (O_913,N_14970,N_14802);
and UO_914 (O_914,N_14906,N_14836);
or UO_915 (O_915,N_14896,N_14860);
nor UO_916 (O_916,N_14861,N_14894);
and UO_917 (O_917,N_14960,N_14978);
nand UO_918 (O_918,N_14923,N_14891);
xnor UO_919 (O_919,N_14922,N_14880);
xnor UO_920 (O_920,N_14821,N_14824);
nor UO_921 (O_921,N_14974,N_14957);
and UO_922 (O_922,N_14932,N_14863);
nand UO_923 (O_923,N_14971,N_14874);
nor UO_924 (O_924,N_14996,N_14974);
nor UO_925 (O_925,N_14958,N_14955);
xor UO_926 (O_926,N_14937,N_14922);
nor UO_927 (O_927,N_14873,N_14890);
nor UO_928 (O_928,N_14968,N_14843);
or UO_929 (O_929,N_14897,N_14826);
nand UO_930 (O_930,N_14855,N_14916);
and UO_931 (O_931,N_14952,N_14872);
nor UO_932 (O_932,N_14930,N_14916);
and UO_933 (O_933,N_14902,N_14943);
or UO_934 (O_934,N_14927,N_14997);
xor UO_935 (O_935,N_14839,N_14826);
nand UO_936 (O_936,N_14937,N_14957);
xnor UO_937 (O_937,N_14809,N_14847);
and UO_938 (O_938,N_14920,N_14883);
xnor UO_939 (O_939,N_14978,N_14840);
xor UO_940 (O_940,N_14809,N_14872);
or UO_941 (O_941,N_14907,N_14937);
and UO_942 (O_942,N_14845,N_14888);
nand UO_943 (O_943,N_14851,N_14885);
xnor UO_944 (O_944,N_14843,N_14977);
or UO_945 (O_945,N_14935,N_14943);
or UO_946 (O_946,N_14986,N_14928);
or UO_947 (O_947,N_14864,N_14976);
and UO_948 (O_948,N_14868,N_14931);
nand UO_949 (O_949,N_14969,N_14841);
nand UO_950 (O_950,N_14917,N_14968);
or UO_951 (O_951,N_14954,N_14806);
xnor UO_952 (O_952,N_14889,N_14871);
nand UO_953 (O_953,N_14856,N_14954);
and UO_954 (O_954,N_14986,N_14865);
and UO_955 (O_955,N_14893,N_14874);
and UO_956 (O_956,N_14843,N_14936);
or UO_957 (O_957,N_14851,N_14802);
nand UO_958 (O_958,N_14953,N_14999);
and UO_959 (O_959,N_14871,N_14881);
xnor UO_960 (O_960,N_14878,N_14902);
nor UO_961 (O_961,N_14960,N_14987);
nor UO_962 (O_962,N_14988,N_14929);
xnor UO_963 (O_963,N_14810,N_14892);
nand UO_964 (O_964,N_14978,N_14926);
xor UO_965 (O_965,N_14817,N_14921);
nor UO_966 (O_966,N_14878,N_14884);
nor UO_967 (O_967,N_14922,N_14842);
nand UO_968 (O_968,N_14861,N_14951);
xor UO_969 (O_969,N_14838,N_14876);
and UO_970 (O_970,N_14959,N_14810);
nand UO_971 (O_971,N_14807,N_14842);
xor UO_972 (O_972,N_14928,N_14859);
xor UO_973 (O_973,N_14908,N_14917);
nand UO_974 (O_974,N_14987,N_14971);
and UO_975 (O_975,N_14913,N_14906);
and UO_976 (O_976,N_14875,N_14997);
xor UO_977 (O_977,N_14870,N_14970);
nor UO_978 (O_978,N_14809,N_14905);
or UO_979 (O_979,N_14938,N_14982);
xor UO_980 (O_980,N_14989,N_14889);
or UO_981 (O_981,N_14855,N_14848);
nand UO_982 (O_982,N_14858,N_14961);
and UO_983 (O_983,N_14825,N_14944);
nor UO_984 (O_984,N_14894,N_14908);
nor UO_985 (O_985,N_14806,N_14937);
and UO_986 (O_986,N_14853,N_14874);
or UO_987 (O_987,N_14866,N_14958);
xnor UO_988 (O_988,N_14911,N_14909);
nor UO_989 (O_989,N_14881,N_14822);
or UO_990 (O_990,N_14951,N_14870);
and UO_991 (O_991,N_14856,N_14859);
and UO_992 (O_992,N_14918,N_14878);
or UO_993 (O_993,N_14985,N_14939);
xnor UO_994 (O_994,N_14842,N_14883);
or UO_995 (O_995,N_14946,N_14885);
nor UO_996 (O_996,N_14816,N_14902);
and UO_997 (O_997,N_14892,N_14864);
nand UO_998 (O_998,N_14890,N_14935);
xor UO_999 (O_999,N_14965,N_14987);
or UO_1000 (O_1000,N_14815,N_14902);
and UO_1001 (O_1001,N_14935,N_14962);
nor UO_1002 (O_1002,N_14819,N_14899);
nand UO_1003 (O_1003,N_14988,N_14829);
or UO_1004 (O_1004,N_14818,N_14879);
xor UO_1005 (O_1005,N_14802,N_14937);
nor UO_1006 (O_1006,N_14933,N_14839);
xor UO_1007 (O_1007,N_14831,N_14861);
and UO_1008 (O_1008,N_14938,N_14945);
and UO_1009 (O_1009,N_14849,N_14920);
and UO_1010 (O_1010,N_14943,N_14946);
nand UO_1011 (O_1011,N_14812,N_14927);
xnor UO_1012 (O_1012,N_14970,N_14903);
nand UO_1013 (O_1013,N_14848,N_14947);
nand UO_1014 (O_1014,N_14951,N_14801);
and UO_1015 (O_1015,N_14858,N_14954);
xnor UO_1016 (O_1016,N_14957,N_14829);
and UO_1017 (O_1017,N_14802,N_14827);
and UO_1018 (O_1018,N_14942,N_14911);
or UO_1019 (O_1019,N_14884,N_14864);
nand UO_1020 (O_1020,N_14989,N_14840);
xor UO_1021 (O_1021,N_14804,N_14843);
and UO_1022 (O_1022,N_14976,N_14977);
nor UO_1023 (O_1023,N_14837,N_14861);
nand UO_1024 (O_1024,N_14805,N_14872);
xor UO_1025 (O_1025,N_14820,N_14832);
and UO_1026 (O_1026,N_14951,N_14947);
xor UO_1027 (O_1027,N_14848,N_14866);
xnor UO_1028 (O_1028,N_14881,N_14949);
or UO_1029 (O_1029,N_14921,N_14867);
nor UO_1030 (O_1030,N_14908,N_14880);
nand UO_1031 (O_1031,N_14985,N_14937);
and UO_1032 (O_1032,N_14927,N_14903);
and UO_1033 (O_1033,N_14844,N_14977);
xnor UO_1034 (O_1034,N_14862,N_14815);
nor UO_1035 (O_1035,N_14805,N_14910);
or UO_1036 (O_1036,N_14819,N_14898);
and UO_1037 (O_1037,N_14841,N_14993);
nor UO_1038 (O_1038,N_14917,N_14977);
nor UO_1039 (O_1039,N_14906,N_14801);
nor UO_1040 (O_1040,N_14931,N_14925);
and UO_1041 (O_1041,N_14974,N_14866);
nor UO_1042 (O_1042,N_14907,N_14999);
nor UO_1043 (O_1043,N_14874,N_14804);
xor UO_1044 (O_1044,N_14933,N_14936);
nand UO_1045 (O_1045,N_14830,N_14802);
or UO_1046 (O_1046,N_14861,N_14848);
xor UO_1047 (O_1047,N_14974,N_14854);
nor UO_1048 (O_1048,N_14836,N_14997);
nand UO_1049 (O_1049,N_14821,N_14954);
nand UO_1050 (O_1050,N_14921,N_14984);
and UO_1051 (O_1051,N_14972,N_14917);
or UO_1052 (O_1052,N_14924,N_14908);
and UO_1053 (O_1053,N_14909,N_14842);
nand UO_1054 (O_1054,N_14861,N_14864);
or UO_1055 (O_1055,N_14831,N_14822);
or UO_1056 (O_1056,N_14990,N_14850);
nor UO_1057 (O_1057,N_14855,N_14853);
and UO_1058 (O_1058,N_14820,N_14882);
or UO_1059 (O_1059,N_14810,N_14925);
xnor UO_1060 (O_1060,N_14837,N_14895);
nor UO_1061 (O_1061,N_14959,N_14827);
nor UO_1062 (O_1062,N_14953,N_14974);
nand UO_1063 (O_1063,N_14841,N_14806);
xor UO_1064 (O_1064,N_14874,N_14838);
xor UO_1065 (O_1065,N_14897,N_14845);
nor UO_1066 (O_1066,N_14909,N_14894);
xor UO_1067 (O_1067,N_14991,N_14857);
xnor UO_1068 (O_1068,N_14971,N_14877);
or UO_1069 (O_1069,N_14906,N_14891);
nand UO_1070 (O_1070,N_14955,N_14884);
xor UO_1071 (O_1071,N_14984,N_14867);
or UO_1072 (O_1072,N_14865,N_14906);
nor UO_1073 (O_1073,N_14974,N_14867);
nand UO_1074 (O_1074,N_14854,N_14941);
nand UO_1075 (O_1075,N_14862,N_14950);
or UO_1076 (O_1076,N_14998,N_14923);
and UO_1077 (O_1077,N_14988,N_14960);
nand UO_1078 (O_1078,N_14890,N_14954);
xnor UO_1079 (O_1079,N_14822,N_14851);
xnor UO_1080 (O_1080,N_14933,N_14996);
and UO_1081 (O_1081,N_14951,N_14983);
nand UO_1082 (O_1082,N_14894,N_14982);
nand UO_1083 (O_1083,N_14845,N_14861);
or UO_1084 (O_1084,N_14989,N_14923);
and UO_1085 (O_1085,N_14963,N_14844);
xnor UO_1086 (O_1086,N_14968,N_14997);
nand UO_1087 (O_1087,N_14869,N_14918);
nand UO_1088 (O_1088,N_14846,N_14977);
nor UO_1089 (O_1089,N_14920,N_14817);
and UO_1090 (O_1090,N_14899,N_14932);
and UO_1091 (O_1091,N_14821,N_14977);
nand UO_1092 (O_1092,N_14902,N_14937);
xor UO_1093 (O_1093,N_14872,N_14856);
or UO_1094 (O_1094,N_14847,N_14853);
nor UO_1095 (O_1095,N_14948,N_14939);
or UO_1096 (O_1096,N_14999,N_14819);
xnor UO_1097 (O_1097,N_14869,N_14871);
nor UO_1098 (O_1098,N_14989,N_14977);
nand UO_1099 (O_1099,N_14955,N_14815);
or UO_1100 (O_1100,N_14802,N_14816);
nor UO_1101 (O_1101,N_14957,N_14946);
xor UO_1102 (O_1102,N_14885,N_14839);
and UO_1103 (O_1103,N_14952,N_14888);
or UO_1104 (O_1104,N_14975,N_14934);
and UO_1105 (O_1105,N_14923,N_14948);
nand UO_1106 (O_1106,N_14834,N_14914);
and UO_1107 (O_1107,N_14951,N_14982);
nand UO_1108 (O_1108,N_14864,N_14993);
or UO_1109 (O_1109,N_14971,N_14908);
nor UO_1110 (O_1110,N_14908,N_14876);
and UO_1111 (O_1111,N_14803,N_14982);
xnor UO_1112 (O_1112,N_14985,N_14935);
or UO_1113 (O_1113,N_14869,N_14824);
nand UO_1114 (O_1114,N_14923,N_14870);
nor UO_1115 (O_1115,N_14855,N_14899);
nand UO_1116 (O_1116,N_14889,N_14872);
nor UO_1117 (O_1117,N_14996,N_14983);
or UO_1118 (O_1118,N_14910,N_14916);
xnor UO_1119 (O_1119,N_14890,N_14996);
nor UO_1120 (O_1120,N_14864,N_14844);
or UO_1121 (O_1121,N_14947,N_14890);
or UO_1122 (O_1122,N_14819,N_14948);
and UO_1123 (O_1123,N_14943,N_14820);
nand UO_1124 (O_1124,N_14832,N_14833);
nand UO_1125 (O_1125,N_14895,N_14976);
nand UO_1126 (O_1126,N_14853,N_14932);
xor UO_1127 (O_1127,N_14910,N_14855);
xnor UO_1128 (O_1128,N_14996,N_14977);
xnor UO_1129 (O_1129,N_14926,N_14931);
or UO_1130 (O_1130,N_14814,N_14927);
nor UO_1131 (O_1131,N_14812,N_14885);
nand UO_1132 (O_1132,N_14959,N_14850);
xor UO_1133 (O_1133,N_14837,N_14820);
nand UO_1134 (O_1134,N_14801,N_14899);
xnor UO_1135 (O_1135,N_14858,N_14908);
xnor UO_1136 (O_1136,N_14843,N_14934);
and UO_1137 (O_1137,N_14902,N_14803);
xor UO_1138 (O_1138,N_14949,N_14869);
or UO_1139 (O_1139,N_14824,N_14846);
and UO_1140 (O_1140,N_14979,N_14968);
nand UO_1141 (O_1141,N_14827,N_14878);
nor UO_1142 (O_1142,N_14824,N_14998);
nand UO_1143 (O_1143,N_14999,N_14816);
nand UO_1144 (O_1144,N_14941,N_14811);
or UO_1145 (O_1145,N_14913,N_14964);
nand UO_1146 (O_1146,N_14944,N_14990);
and UO_1147 (O_1147,N_14825,N_14931);
nand UO_1148 (O_1148,N_14837,N_14800);
nor UO_1149 (O_1149,N_14800,N_14920);
or UO_1150 (O_1150,N_14840,N_14910);
nand UO_1151 (O_1151,N_14899,N_14915);
or UO_1152 (O_1152,N_14955,N_14848);
xnor UO_1153 (O_1153,N_14848,N_14906);
xor UO_1154 (O_1154,N_14909,N_14872);
and UO_1155 (O_1155,N_14930,N_14952);
and UO_1156 (O_1156,N_14835,N_14810);
nor UO_1157 (O_1157,N_14973,N_14825);
and UO_1158 (O_1158,N_14988,N_14862);
or UO_1159 (O_1159,N_14806,N_14968);
or UO_1160 (O_1160,N_14860,N_14870);
or UO_1161 (O_1161,N_14926,N_14908);
nand UO_1162 (O_1162,N_14915,N_14866);
nand UO_1163 (O_1163,N_14920,N_14821);
xnor UO_1164 (O_1164,N_14932,N_14982);
or UO_1165 (O_1165,N_14974,N_14902);
nor UO_1166 (O_1166,N_14869,N_14850);
xnor UO_1167 (O_1167,N_14848,N_14879);
and UO_1168 (O_1168,N_14810,N_14988);
xnor UO_1169 (O_1169,N_14911,N_14949);
and UO_1170 (O_1170,N_14855,N_14870);
nor UO_1171 (O_1171,N_14985,N_14915);
and UO_1172 (O_1172,N_14896,N_14987);
and UO_1173 (O_1173,N_14872,N_14957);
and UO_1174 (O_1174,N_14876,N_14963);
or UO_1175 (O_1175,N_14955,N_14898);
nand UO_1176 (O_1176,N_14944,N_14876);
or UO_1177 (O_1177,N_14845,N_14974);
or UO_1178 (O_1178,N_14958,N_14873);
nor UO_1179 (O_1179,N_14965,N_14879);
or UO_1180 (O_1180,N_14899,N_14843);
or UO_1181 (O_1181,N_14817,N_14971);
or UO_1182 (O_1182,N_14890,N_14997);
nor UO_1183 (O_1183,N_14841,N_14983);
and UO_1184 (O_1184,N_14937,N_14994);
or UO_1185 (O_1185,N_14968,N_14960);
xor UO_1186 (O_1186,N_14948,N_14875);
or UO_1187 (O_1187,N_14879,N_14884);
xnor UO_1188 (O_1188,N_14826,N_14857);
nand UO_1189 (O_1189,N_14894,N_14927);
and UO_1190 (O_1190,N_14978,N_14952);
or UO_1191 (O_1191,N_14936,N_14967);
xnor UO_1192 (O_1192,N_14838,N_14829);
xor UO_1193 (O_1193,N_14911,N_14984);
and UO_1194 (O_1194,N_14953,N_14955);
nand UO_1195 (O_1195,N_14982,N_14899);
nand UO_1196 (O_1196,N_14864,N_14849);
nand UO_1197 (O_1197,N_14875,N_14950);
nand UO_1198 (O_1198,N_14847,N_14863);
and UO_1199 (O_1199,N_14934,N_14802);
nor UO_1200 (O_1200,N_14883,N_14840);
nor UO_1201 (O_1201,N_14976,N_14904);
or UO_1202 (O_1202,N_14822,N_14907);
nand UO_1203 (O_1203,N_14935,N_14946);
or UO_1204 (O_1204,N_14906,N_14827);
and UO_1205 (O_1205,N_14916,N_14973);
nor UO_1206 (O_1206,N_14961,N_14884);
xnor UO_1207 (O_1207,N_14910,N_14800);
nor UO_1208 (O_1208,N_14974,N_14894);
nand UO_1209 (O_1209,N_14811,N_14825);
and UO_1210 (O_1210,N_14927,N_14973);
nand UO_1211 (O_1211,N_14973,N_14807);
nand UO_1212 (O_1212,N_14992,N_14833);
and UO_1213 (O_1213,N_14973,N_14863);
nand UO_1214 (O_1214,N_14879,N_14827);
xnor UO_1215 (O_1215,N_14961,N_14859);
or UO_1216 (O_1216,N_14807,N_14871);
or UO_1217 (O_1217,N_14890,N_14978);
nand UO_1218 (O_1218,N_14884,N_14819);
nor UO_1219 (O_1219,N_14985,N_14818);
and UO_1220 (O_1220,N_14895,N_14844);
xor UO_1221 (O_1221,N_14990,N_14869);
nor UO_1222 (O_1222,N_14930,N_14871);
or UO_1223 (O_1223,N_14819,N_14910);
xor UO_1224 (O_1224,N_14952,N_14927);
and UO_1225 (O_1225,N_14825,N_14836);
nand UO_1226 (O_1226,N_14866,N_14882);
and UO_1227 (O_1227,N_14919,N_14977);
nand UO_1228 (O_1228,N_14876,N_14921);
and UO_1229 (O_1229,N_14876,N_14812);
nand UO_1230 (O_1230,N_14890,N_14840);
nor UO_1231 (O_1231,N_14875,N_14850);
xor UO_1232 (O_1232,N_14862,N_14806);
or UO_1233 (O_1233,N_14897,N_14967);
xor UO_1234 (O_1234,N_14938,N_14940);
nor UO_1235 (O_1235,N_14867,N_14933);
nand UO_1236 (O_1236,N_14806,N_14893);
nand UO_1237 (O_1237,N_14825,N_14850);
or UO_1238 (O_1238,N_14854,N_14915);
nand UO_1239 (O_1239,N_14858,N_14909);
xor UO_1240 (O_1240,N_14847,N_14923);
nor UO_1241 (O_1241,N_14879,N_14992);
xnor UO_1242 (O_1242,N_14836,N_14828);
nor UO_1243 (O_1243,N_14928,N_14913);
nand UO_1244 (O_1244,N_14883,N_14909);
nor UO_1245 (O_1245,N_14928,N_14817);
or UO_1246 (O_1246,N_14805,N_14915);
and UO_1247 (O_1247,N_14869,N_14926);
or UO_1248 (O_1248,N_14992,N_14898);
nor UO_1249 (O_1249,N_14828,N_14955);
and UO_1250 (O_1250,N_14944,N_14961);
nand UO_1251 (O_1251,N_14876,N_14916);
nor UO_1252 (O_1252,N_14998,N_14986);
or UO_1253 (O_1253,N_14867,N_14965);
and UO_1254 (O_1254,N_14984,N_14882);
nor UO_1255 (O_1255,N_14807,N_14878);
or UO_1256 (O_1256,N_14885,N_14830);
xnor UO_1257 (O_1257,N_14829,N_14978);
nand UO_1258 (O_1258,N_14814,N_14835);
nor UO_1259 (O_1259,N_14963,N_14833);
or UO_1260 (O_1260,N_14878,N_14952);
nand UO_1261 (O_1261,N_14874,N_14855);
nor UO_1262 (O_1262,N_14921,N_14845);
or UO_1263 (O_1263,N_14806,N_14956);
nand UO_1264 (O_1264,N_14924,N_14826);
xnor UO_1265 (O_1265,N_14888,N_14892);
nand UO_1266 (O_1266,N_14890,N_14886);
nor UO_1267 (O_1267,N_14832,N_14926);
or UO_1268 (O_1268,N_14935,N_14951);
and UO_1269 (O_1269,N_14832,N_14897);
nor UO_1270 (O_1270,N_14818,N_14872);
or UO_1271 (O_1271,N_14919,N_14920);
or UO_1272 (O_1272,N_14995,N_14901);
xnor UO_1273 (O_1273,N_14993,N_14921);
nand UO_1274 (O_1274,N_14808,N_14904);
and UO_1275 (O_1275,N_14892,N_14970);
xor UO_1276 (O_1276,N_14892,N_14886);
xnor UO_1277 (O_1277,N_14873,N_14842);
xor UO_1278 (O_1278,N_14917,N_14934);
and UO_1279 (O_1279,N_14853,N_14872);
nand UO_1280 (O_1280,N_14828,N_14831);
or UO_1281 (O_1281,N_14963,N_14913);
xnor UO_1282 (O_1282,N_14840,N_14939);
or UO_1283 (O_1283,N_14945,N_14849);
and UO_1284 (O_1284,N_14805,N_14882);
nor UO_1285 (O_1285,N_14906,N_14862);
nand UO_1286 (O_1286,N_14937,N_14961);
xnor UO_1287 (O_1287,N_14906,N_14823);
xnor UO_1288 (O_1288,N_14897,N_14827);
xor UO_1289 (O_1289,N_14963,N_14846);
xnor UO_1290 (O_1290,N_14824,N_14880);
and UO_1291 (O_1291,N_14879,N_14895);
or UO_1292 (O_1292,N_14926,N_14957);
nand UO_1293 (O_1293,N_14973,N_14914);
nor UO_1294 (O_1294,N_14852,N_14836);
nor UO_1295 (O_1295,N_14997,N_14993);
nand UO_1296 (O_1296,N_14903,N_14975);
nand UO_1297 (O_1297,N_14825,N_14845);
nor UO_1298 (O_1298,N_14979,N_14897);
nand UO_1299 (O_1299,N_14807,N_14872);
xnor UO_1300 (O_1300,N_14926,N_14865);
nand UO_1301 (O_1301,N_14908,N_14801);
xor UO_1302 (O_1302,N_14985,N_14871);
nand UO_1303 (O_1303,N_14883,N_14805);
and UO_1304 (O_1304,N_14922,N_14888);
or UO_1305 (O_1305,N_14812,N_14901);
nor UO_1306 (O_1306,N_14950,N_14973);
xnor UO_1307 (O_1307,N_14980,N_14984);
xor UO_1308 (O_1308,N_14937,N_14990);
nor UO_1309 (O_1309,N_14942,N_14916);
nand UO_1310 (O_1310,N_14969,N_14981);
or UO_1311 (O_1311,N_14838,N_14868);
nand UO_1312 (O_1312,N_14800,N_14908);
or UO_1313 (O_1313,N_14999,N_14873);
nand UO_1314 (O_1314,N_14868,N_14872);
nand UO_1315 (O_1315,N_14898,N_14976);
or UO_1316 (O_1316,N_14869,N_14810);
xnor UO_1317 (O_1317,N_14839,N_14990);
nand UO_1318 (O_1318,N_14915,N_14809);
nor UO_1319 (O_1319,N_14960,N_14944);
and UO_1320 (O_1320,N_14925,N_14906);
nand UO_1321 (O_1321,N_14908,N_14952);
nand UO_1322 (O_1322,N_14836,N_14993);
and UO_1323 (O_1323,N_14887,N_14879);
nor UO_1324 (O_1324,N_14981,N_14998);
nand UO_1325 (O_1325,N_14935,N_14941);
or UO_1326 (O_1326,N_14920,N_14869);
or UO_1327 (O_1327,N_14944,N_14889);
or UO_1328 (O_1328,N_14832,N_14805);
or UO_1329 (O_1329,N_14888,N_14849);
nand UO_1330 (O_1330,N_14891,N_14920);
or UO_1331 (O_1331,N_14877,N_14992);
nor UO_1332 (O_1332,N_14867,N_14865);
xor UO_1333 (O_1333,N_14862,N_14814);
xnor UO_1334 (O_1334,N_14982,N_14918);
xnor UO_1335 (O_1335,N_14899,N_14924);
or UO_1336 (O_1336,N_14902,N_14903);
nor UO_1337 (O_1337,N_14804,N_14994);
or UO_1338 (O_1338,N_14891,N_14974);
and UO_1339 (O_1339,N_14885,N_14952);
nor UO_1340 (O_1340,N_14823,N_14862);
or UO_1341 (O_1341,N_14835,N_14865);
nor UO_1342 (O_1342,N_14965,N_14818);
nand UO_1343 (O_1343,N_14899,N_14910);
or UO_1344 (O_1344,N_14855,N_14834);
nor UO_1345 (O_1345,N_14810,N_14906);
xnor UO_1346 (O_1346,N_14861,N_14986);
nor UO_1347 (O_1347,N_14803,N_14887);
and UO_1348 (O_1348,N_14837,N_14876);
nand UO_1349 (O_1349,N_14815,N_14934);
xnor UO_1350 (O_1350,N_14916,N_14979);
xor UO_1351 (O_1351,N_14946,N_14973);
nand UO_1352 (O_1352,N_14963,N_14865);
nand UO_1353 (O_1353,N_14919,N_14926);
xor UO_1354 (O_1354,N_14960,N_14894);
and UO_1355 (O_1355,N_14952,N_14911);
nand UO_1356 (O_1356,N_14844,N_14849);
and UO_1357 (O_1357,N_14866,N_14977);
xor UO_1358 (O_1358,N_14850,N_14985);
xnor UO_1359 (O_1359,N_14805,N_14917);
and UO_1360 (O_1360,N_14823,N_14969);
nand UO_1361 (O_1361,N_14880,N_14816);
or UO_1362 (O_1362,N_14847,N_14906);
xor UO_1363 (O_1363,N_14837,N_14838);
xnor UO_1364 (O_1364,N_14823,N_14981);
or UO_1365 (O_1365,N_14887,N_14864);
xnor UO_1366 (O_1366,N_14961,N_14935);
nand UO_1367 (O_1367,N_14926,N_14955);
or UO_1368 (O_1368,N_14805,N_14959);
xor UO_1369 (O_1369,N_14970,N_14851);
nand UO_1370 (O_1370,N_14805,N_14942);
nor UO_1371 (O_1371,N_14945,N_14951);
nand UO_1372 (O_1372,N_14969,N_14880);
nor UO_1373 (O_1373,N_14926,N_14900);
or UO_1374 (O_1374,N_14848,N_14819);
nor UO_1375 (O_1375,N_14853,N_14939);
or UO_1376 (O_1376,N_14987,N_14951);
xor UO_1377 (O_1377,N_14911,N_14979);
nor UO_1378 (O_1378,N_14843,N_14875);
and UO_1379 (O_1379,N_14824,N_14915);
or UO_1380 (O_1380,N_14879,N_14958);
or UO_1381 (O_1381,N_14842,N_14986);
xor UO_1382 (O_1382,N_14823,N_14971);
nor UO_1383 (O_1383,N_14912,N_14822);
or UO_1384 (O_1384,N_14989,N_14970);
and UO_1385 (O_1385,N_14852,N_14953);
nand UO_1386 (O_1386,N_14842,N_14884);
or UO_1387 (O_1387,N_14928,N_14910);
xor UO_1388 (O_1388,N_14973,N_14923);
or UO_1389 (O_1389,N_14918,N_14900);
and UO_1390 (O_1390,N_14975,N_14878);
and UO_1391 (O_1391,N_14987,N_14858);
or UO_1392 (O_1392,N_14925,N_14951);
or UO_1393 (O_1393,N_14801,N_14919);
xnor UO_1394 (O_1394,N_14889,N_14920);
and UO_1395 (O_1395,N_14800,N_14932);
nand UO_1396 (O_1396,N_14825,N_14841);
or UO_1397 (O_1397,N_14911,N_14972);
nor UO_1398 (O_1398,N_14908,N_14824);
nand UO_1399 (O_1399,N_14874,N_14939);
nor UO_1400 (O_1400,N_14989,N_14928);
and UO_1401 (O_1401,N_14936,N_14903);
nand UO_1402 (O_1402,N_14925,N_14972);
nand UO_1403 (O_1403,N_14900,N_14915);
nor UO_1404 (O_1404,N_14996,N_14898);
nand UO_1405 (O_1405,N_14996,N_14975);
and UO_1406 (O_1406,N_14881,N_14829);
xnor UO_1407 (O_1407,N_14924,N_14842);
xnor UO_1408 (O_1408,N_14952,N_14901);
nor UO_1409 (O_1409,N_14831,N_14848);
or UO_1410 (O_1410,N_14925,N_14952);
xor UO_1411 (O_1411,N_14906,N_14950);
or UO_1412 (O_1412,N_14952,N_14965);
or UO_1413 (O_1413,N_14842,N_14840);
nor UO_1414 (O_1414,N_14931,N_14923);
nor UO_1415 (O_1415,N_14913,N_14985);
and UO_1416 (O_1416,N_14932,N_14878);
xor UO_1417 (O_1417,N_14983,N_14824);
xnor UO_1418 (O_1418,N_14934,N_14836);
or UO_1419 (O_1419,N_14860,N_14855);
or UO_1420 (O_1420,N_14844,N_14824);
nand UO_1421 (O_1421,N_14852,N_14859);
nand UO_1422 (O_1422,N_14869,N_14908);
or UO_1423 (O_1423,N_14894,N_14955);
nor UO_1424 (O_1424,N_14990,N_14816);
or UO_1425 (O_1425,N_14911,N_14865);
and UO_1426 (O_1426,N_14897,N_14944);
and UO_1427 (O_1427,N_14971,N_14831);
nor UO_1428 (O_1428,N_14971,N_14946);
nor UO_1429 (O_1429,N_14951,N_14853);
nor UO_1430 (O_1430,N_14812,N_14833);
nor UO_1431 (O_1431,N_14992,N_14811);
nor UO_1432 (O_1432,N_14971,N_14879);
xnor UO_1433 (O_1433,N_14984,N_14919);
xnor UO_1434 (O_1434,N_14864,N_14865);
and UO_1435 (O_1435,N_14936,N_14825);
nor UO_1436 (O_1436,N_14967,N_14842);
or UO_1437 (O_1437,N_14821,N_14974);
xnor UO_1438 (O_1438,N_14833,N_14818);
or UO_1439 (O_1439,N_14867,N_14972);
nor UO_1440 (O_1440,N_14950,N_14866);
or UO_1441 (O_1441,N_14870,N_14858);
nor UO_1442 (O_1442,N_14907,N_14942);
nor UO_1443 (O_1443,N_14922,N_14874);
nand UO_1444 (O_1444,N_14918,N_14830);
xor UO_1445 (O_1445,N_14854,N_14933);
nand UO_1446 (O_1446,N_14959,N_14855);
xnor UO_1447 (O_1447,N_14896,N_14931);
and UO_1448 (O_1448,N_14832,N_14822);
nand UO_1449 (O_1449,N_14862,N_14819);
and UO_1450 (O_1450,N_14851,N_14827);
nor UO_1451 (O_1451,N_14875,N_14836);
nand UO_1452 (O_1452,N_14820,N_14975);
and UO_1453 (O_1453,N_14894,N_14873);
nor UO_1454 (O_1454,N_14973,N_14856);
or UO_1455 (O_1455,N_14943,N_14920);
and UO_1456 (O_1456,N_14961,N_14830);
nand UO_1457 (O_1457,N_14886,N_14819);
or UO_1458 (O_1458,N_14884,N_14817);
nor UO_1459 (O_1459,N_14954,N_14909);
and UO_1460 (O_1460,N_14835,N_14867);
and UO_1461 (O_1461,N_14878,N_14947);
nor UO_1462 (O_1462,N_14904,N_14813);
and UO_1463 (O_1463,N_14906,N_14804);
nor UO_1464 (O_1464,N_14818,N_14870);
xnor UO_1465 (O_1465,N_14922,N_14995);
or UO_1466 (O_1466,N_14920,N_14947);
nor UO_1467 (O_1467,N_14802,N_14888);
and UO_1468 (O_1468,N_14946,N_14911);
nor UO_1469 (O_1469,N_14950,N_14818);
xor UO_1470 (O_1470,N_14840,N_14897);
and UO_1471 (O_1471,N_14997,N_14911);
xnor UO_1472 (O_1472,N_14838,N_14930);
or UO_1473 (O_1473,N_14880,N_14861);
nand UO_1474 (O_1474,N_14895,N_14965);
or UO_1475 (O_1475,N_14879,N_14869);
and UO_1476 (O_1476,N_14871,N_14949);
xnor UO_1477 (O_1477,N_14989,N_14860);
or UO_1478 (O_1478,N_14822,N_14894);
xnor UO_1479 (O_1479,N_14859,N_14893);
and UO_1480 (O_1480,N_14824,N_14891);
xnor UO_1481 (O_1481,N_14947,N_14949);
nand UO_1482 (O_1482,N_14998,N_14943);
xnor UO_1483 (O_1483,N_14844,N_14992);
nor UO_1484 (O_1484,N_14890,N_14945);
nand UO_1485 (O_1485,N_14904,N_14845);
nand UO_1486 (O_1486,N_14815,N_14892);
nor UO_1487 (O_1487,N_14859,N_14921);
xor UO_1488 (O_1488,N_14876,N_14897);
nand UO_1489 (O_1489,N_14889,N_14949);
nand UO_1490 (O_1490,N_14808,N_14822);
or UO_1491 (O_1491,N_14954,N_14988);
xnor UO_1492 (O_1492,N_14854,N_14905);
nor UO_1493 (O_1493,N_14905,N_14893);
xor UO_1494 (O_1494,N_14863,N_14975);
nand UO_1495 (O_1495,N_14971,N_14803);
nor UO_1496 (O_1496,N_14931,N_14856);
nand UO_1497 (O_1497,N_14924,N_14907);
or UO_1498 (O_1498,N_14864,N_14863);
or UO_1499 (O_1499,N_14989,N_14867);
and UO_1500 (O_1500,N_14982,N_14829);
nor UO_1501 (O_1501,N_14963,N_14872);
nand UO_1502 (O_1502,N_14979,N_14902);
and UO_1503 (O_1503,N_14951,N_14863);
or UO_1504 (O_1504,N_14914,N_14935);
and UO_1505 (O_1505,N_14839,N_14911);
or UO_1506 (O_1506,N_14800,N_14966);
and UO_1507 (O_1507,N_14915,N_14876);
nor UO_1508 (O_1508,N_14844,N_14897);
and UO_1509 (O_1509,N_14856,N_14975);
or UO_1510 (O_1510,N_14950,N_14802);
and UO_1511 (O_1511,N_14871,N_14983);
nor UO_1512 (O_1512,N_14823,N_14953);
or UO_1513 (O_1513,N_14847,N_14882);
and UO_1514 (O_1514,N_14861,N_14942);
nor UO_1515 (O_1515,N_14913,N_14826);
nand UO_1516 (O_1516,N_14832,N_14932);
nor UO_1517 (O_1517,N_14812,N_14873);
nand UO_1518 (O_1518,N_14987,N_14882);
xnor UO_1519 (O_1519,N_14977,N_14806);
xor UO_1520 (O_1520,N_14810,N_14983);
nor UO_1521 (O_1521,N_14826,N_14801);
or UO_1522 (O_1522,N_14842,N_14809);
or UO_1523 (O_1523,N_14832,N_14803);
nor UO_1524 (O_1524,N_14817,N_14968);
and UO_1525 (O_1525,N_14985,N_14900);
or UO_1526 (O_1526,N_14859,N_14960);
nand UO_1527 (O_1527,N_14950,N_14826);
xor UO_1528 (O_1528,N_14991,N_14803);
and UO_1529 (O_1529,N_14873,N_14956);
xor UO_1530 (O_1530,N_14892,N_14966);
or UO_1531 (O_1531,N_14817,N_14860);
or UO_1532 (O_1532,N_14817,N_14999);
xor UO_1533 (O_1533,N_14963,N_14908);
nand UO_1534 (O_1534,N_14836,N_14903);
or UO_1535 (O_1535,N_14801,N_14895);
nand UO_1536 (O_1536,N_14865,N_14937);
nand UO_1537 (O_1537,N_14821,N_14918);
or UO_1538 (O_1538,N_14914,N_14998);
xnor UO_1539 (O_1539,N_14899,N_14994);
nor UO_1540 (O_1540,N_14859,N_14957);
or UO_1541 (O_1541,N_14997,N_14803);
nand UO_1542 (O_1542,N_14838,N_14865);
or UO_1543 (O_1543,N_14921,N_14874);
or UO_1544 (O_1544,N_14832,N_14887);
nor UO_1545 (O_1545,N_14889,N_14992);
nor UO_1546 (O_1546,N_14986,N_14956);
nand UO_1547 (O_1547,N_14961,N_14878);
nor UO_1548 (O_1548,N_14880,N_14817);
xor UO_1549 (O_1549,N_14956,N_14869);
nor UO_1550 (O_1550,N_14950,N_14873);
nor UO_1551 (O_1551,N_14974,N_14952);
nor UO_1552 (O_1552,N_14956,N_14925);
nand UO_1553 (O_1553,N_14829,N_14987);
or UO_1554 (O_1554,N_14804,N_14932);
nand UO_1555 (O_1555,N_14826,N_14908);
and UO_1556 (O_1556,N_14816,N_14846);
nor UO_1557 (O_1557,N_14922,N_14945);
xor UO_1558 (O_1558,N_14911,N_14910);
xnor UO_1559 (O_1559,N_14955,N_14984);
and UO_1560 (O_1560,N_14897,N_14881);
xor UO_1561 (O_1561,N_14863,N_14815);
nand UO_1562 (O_1562,N_14842,N_14832);
and UO_1563 (O_1563,N_14943,N_14839);
and UO_1564 (O_1564,N_14830,N_14972);
and UO_1565 (O_1565,N_14972,N_14815);
and UO_1566 (O_1566,N_14962,N_14809);
nor UO_1567 (O_1567,N_14935,N_14892);
nand UO_1568 (O_1568,N_14869,N_14878);
nor UO_1569 (O_1569,N_14810,N_14902);
nand UO_1570 (O_1570,N_14972,N_14939);
or UO_1571 (O_1571,N_14801,N_14836);
nor UO_1572 (O_1572,N_14963,N_14942);
or UO_1573 (O_1573,N_14981,N_14984);
xnor UO_1574 (O_1574,N_14806,N_14981);
xnor UO_1575 (O_1575,N_14950,N_14927);
and UO_1576 (O_1576,N_14985,N_14828);
or UO_1577 (O_1577,N_14882,N_14972);
and UO_1578 (O_1578,N_14859,N_14905);
xnor UO_1579 (O_1579,N_14874,N_14952);
or UO_1580 (O_1580,N_14957,N_14984);
or UO_1581 (O_1581,N_14902,N_14879);
xor UO_1582 (O_1582,N_14802,N_14932);
nand UO_1583 (O_1583,N_14806,N_14947);
nor UO_1584 (O_1584,N_14939,N_14896);
xor UO_1585 (O_1585,N_14894,N_14844);
and UO_1586 (O_1586,N_14890,N_14866);
xor UO_1587 (O_1587,N_14975,N_14872);
xnor UO_1588 (O_1588,N_14843,N_14844);
and UO_1589 (O_1589,N_14898,N_14828);
xor UO_1590 (O_1590,N_14955,N_14954);
or UO_1591 (O_1591,N_14932,N_14958);
nand UO_1592 (O_1592,N_14913,N_14832);
nand UO_1593 (O_1593,N_14896,N_14822);
or UO_1594 (O_1594,N_14989,N_14950);
nor UO_1595 (O_1595,N_14958,N_14869);
or UO_1596 (O_1596,N_14923,N_14834);
nor UO_1597 (O_1597,N_14827,N_14800);
and UO_1598 (O_1598,N_14908,N_14873);
and UO_1599 (O_1599,N_14803,N_14867);
nor UO_1600 (O_1600,N_14878,N_14979);
xor UO_1601 (O_1601,N_14916,N_14893);
xnor UO_1602 (O_1602,N_14819,N_14861);
or UO_1603 (O_1603,N_14857,N_14986);
or UO_1604 (O_1604,N_14833,N_14838);
nor UO_1605 (O_1605,N_14940,N_14820);
nor UO_1606 (O_1606,N_14827,N_14870);
nor UO_1607 (O_1607,N_14825,N_14945);
nand UO_1608 (O_1608,N_14808,N_14948);
nor UO_1609 (O_1609,N_14821,N_14991);
nor UO_1610 (O_1610,N_14811,N_14934);
nand UO_1611 (O_1611,N_14813,N_14972);
and UO_1612 (O_1612,N_14853,N_14842);
nor UO_1613 (O_1613,N_14818,N_14846);
or UO_1614 (O_1614,N_14873,N_14846);
xor UO_1615 (O_1615,N_14912,N_14849);
or UO_1616 (O_1616,N_14956,N_14890);
or UO_1617 (O_1617,N_14928,N_14902);
and UO_1618 (O_1618,N_14871,N_14818);
xnor UO_1619 (O_1619,N_14951,N_14808);
nand UO_1620 (O_1620,N_14914,N_14863);
and UO_1621 (O_1621,N_14983,N_14899);
and UO_1622 (O_1622,N_14907,N_14947);
or UO_1623 (O_1623,N_14940,N_14896);
nor UO_1624 (O_1624,N_14876,N_14984);
xor UO_1625 (O_1625,N_14808,N_14843);
nor UO_1626 (O_1626,N_14988,N_14994);
xnor UO_1627 (O_1627,N_14896,N_14968);
xor UO_1628 (O_1628,N_14850,N_14971);
xnor UO_1629 (O_1629,N_14812,N_14933);
nand UO_1630 (O_1630,N_14910,N_14885);
and UO_1631 (O_1631,N_14905,N_14886);
or UO_1632 (O_1632,N_14989,N_14939);
nor UO_1633 (O_1633,N_14820,N_14819);
nor UO_1634 (O_1634,N_14839,N_14963);
or UO_1635 (O_1635,N_14962,N_14946);
or UO_1636 (O_1636,N_14881,N_14870);
nand UO_1637 (O_1637,N_14949,N_14972);
xnor UO_1638 (O_1638,N_14865,N_14829);
xor UO_1639 (O_1639,N_14801,N_14898);
nand UO_1640 (O_1640,N_14969,N_14939);
and UO_1641 (O_1641,N_14911,N_14969);
xnor UO_1642 (O_1642,N_14819,N_14817);
xnor UO_1643 (O_1643,N_14984,N_14838);
nand UO_1644 (O_1644,N_14828,N_14871);
nor UO_1645 (O_1645,N_14991,N_14919);
and UO_1646 (O_1646,N_14849,N_14808);
or UO_1647 (O_1647,N_14829,N_14917);
nand UO_1648 (O_1648,N_14849,N_14958);
xnor UO_1649 (O_1649,N_14999,N_14993);
and UO_1650 (O_1650,N_14828,N_14810);
or UO_1651 (O_1651,N_14908,N_14819);
nand UO_1652 (O_1652,N_14943,N_14851);
nand UO_1653 (O_1653,N_14852,N_14944);
nor UO_1654 (O_1654,N_14814,N_14923);
nor UO_1655 (O_1655,N_14977,N_14819);
or UO_1656 (O_1656,N_14850,N_14965);
nand UO_1657 (O_1657,N_14856,N_14821);
nor UO_1658 (O_1658,N_14826,N_14953);
nor UO_1659 (O_1659,N_14931,N_14954);
and UO_1660 (O_1660,N_14815,N_14964);
and UO_1661 (O_1661,N_14905,N_14863);
xnor UO_1662 (O_1662,N_14871,N_14864);
nor UO_1663 (O_1663,N_14839,N_14894);
and UO_1664 (O_1664,N_14874,N_14857);
nor UO_1665 (O_1665,N_14969,N_14822);
and UO_1666 (O_1666,N_14887,N_14982);
and UO_1667 (O_1667,N_14807,N_14819);
and UO_1668 (O_1668,N_14949,N_14984);
nand UO_1669 (O_1669,N_14911,N_14989);
nand UO_1670 (O_1670,N_14999,N_14821);
nand UO_1671 (O_1671,N_14982,N_14942);
nor UO_1672 (O_1672,N_14848,N_14910);
and UO_1673 (O_1673,N_14856,N_14854);
nor UO_1674 (O_1674,N_14876,N_14870);
and UO_1675 (O_1675,N_14856,N_14877);
xor UO_1676 (O_1676,N_14802,N_14922);
xor UO_1677 (O_1677,N_14984,N_14960);
nor UO_1678 (O_1678,N_14831,N_14918);
nand UO_1679 (O_1679,N_14912,N_14954);
and UO_1680 (O_1680,N_14803,N_14912);
nor UO_1681 (O_1681,N_14849,N_14821);
or UO_1682 (O_1682,N_14815,N_14913);
nand UO_1683 (O_1683,N_14959,N_14934);
and UO_1684 (O_1684,N_14957,N_14812);
xnor UO_1685 (O_1685,N_14844,N_14959);
xnor UO_1686 (O_1686,N_14835,N_14881);
nor UO_1687 (O_1687,N_14996,N_14812);
and UO_1688 (O_1688,N_14981,N_14975);
or UO_1689 (O_1689,N_14851,N_14926);
nor UO_1690 (O_1690,N_14982,N_14836);
or UO_1691 (O_1691,N_14940,N_14902);
nor UO_1692 (O_1692,N_14885,N_14929);
nor UO_1693 (O_1693,N_14978,N_14921);
nand UO_1694 (O_1694,N_14802,N_14821);
nand UO_1695 (O_1695,N_14972,N_14889);
nand UO_1696 (O_1696,N_14873,N_14929);
nor UO_1697 (O_1697,N_14806,N_14807);
nand UO_1698 (O_1698,N_14843,N_14877);
xor UO_1699 (O_1699,N_14978,N_14842);
and UO_1700 (O_1700,N_14893,N_14923);
nand UO_1701 (O_1701,N_14850,N_14918);
nor UO_1702 (O_1702,N_14902,N_14917);
xor UO_1703 (O_1703,N_14910,N_14922);
nand UO_1704 (O_1704,N_14866,N_14886);
and UO_1705 (O_1705,N_14904,N_14920);
nor UO_1706 (O_1706,N_14804,N_14949);
nor UO_1707 (O_1707,N_14847,N_14848);
nand UO_1708 (O_1708,N_14960,N_14858);
or UO_1709 (O_1709,N_14906,N_14958);
nand UO_1710 (O_1710,N_14849,N_14933);
and UO_1711 (O_1711,N_14861,N_14992);
and UO_1712 (O_1712,N_14952,N_14859);
and UO_1713 (O_1713,N_14921,N_14832);
or UO_1714 (O_1714,N_14856,N_14956);
nand UO_1715 (O_1715,N_14902,N_14865);
nor UO_1716 (O_1716,N_14825,N_14980);
nand UO_1717 (O_1717,N_14809,N_14901);
nand UO_1718 (O_1718,N_14840,N_14928);
nor UO_1719 (O_1719,N_14868,N_14810);
nor UO_1720 (O_1720,N_14835,N_14843);
nor UO_1721 (O_1721,N_14860,N_14849);
nand UO_1722 (O_1722,N_14985,N_14979);
nand UO_1723 (O_1723,N_14918,N_14985);
or UO_1724 (O_1724,N_14957,N_14980);
nor UO_1725 (O_1725,N_14840,N_14944);
or UO_1726 (O_1726,N_14895,N_14957);
xor UO_1727 (O_1727,N_14992,N_14936);
or UO_1728 (O_1728,N_14906,N_14841);
or UO_1729 (O_1729,N_14920,N_14983);
nor UO_1730 (O_1730,N_14817,N_14842);
nand UO_1731 (O_1731,N_14948,N_14817);
nand UO_1732 (O_1732,N_14941,N_14984);
and UO_1733 (O_1733,N_14988,N_14965);
nand UO_1734 (O_1734,N_14833,N_14945);
or UO_1735 (O_1735,N_14940,N_14868);
nand UO_1736 (O_1736,N_14883,N_14916);
and UO_1737 (O_1737,N_14821,N_14854);
xnor UO_1738 (O_1738,N_14960,N_14831);
and UO_1739 (O_1739,N_14977,N_14868);
xor UO_1740 (O_1740,N_14931,N_14979);
and UO_1741 (O_1741,N_14923,N_14858);
and UO_1742 (O_1742,N_14863,N_14930);
nand UO_1743 (O_1743,N_14908,N_14836);
or UO_1744 (O_1744,N_14930,N_14974);
xor UO_1745 (O_1745,N_14973,N_14909);
xor UO_1746 (O_1746,N_14896,N_14959);
xnor UO_1747 (O_1747,N_14922,N_14846);
or UO_1748 (O_1748,N_14884,N_14973);
nand UO_1749 (O_1749,N_14965,N_14817);
and UO_1750 (O_1750,N_14841,N_14804);
nor UO_1751 (O_1751,N_14921,N_14934);
xor UO_1752 (O_1752,N_14859,N_14907);
nor UO_1753 (O_1753,N_14813,N_14878);
and UO_1754 (O_1754,N_14857,N_14957);
nor UO_1755 (O_1755,N_14851,N_14962);
nor UO_1756 (O_1756,N_14892,N_14923);
nor UO_1757 (O_1757,N_14821,N_14835);
or UO_1758 (O_1758,N_14852,N_14952);
nor UO_1759 (O_1759,N_14950,N_14964);
nor UO_1760 (O_1760,N_14956,N_14858);
and UO_1761 (O_1761,N_14816,N_14916);
or UO_1762 (O_1762,N_14880,N_14933);
or UO_1763 (O_1763,N_14869,N_14809);
nand UO_1764 (O_1764,N_14896,N_14997);
xnor UO_1765 (O_1765,N_14985,N_14814);
nor UO_1766 (O_1766,N_14903,N_14999);
and UO_1767 (O_1767,N_14985,N_14835);
or UO_1768 (O_1768,N_14876,N_14958);
and UO_1769 (O_1769,N_14918,N_14971);
and UO_1770 (O_1770,N_14859,N_14959);
nand UO_1771 (O_1771,N_14816,N_14984);
xor UO_1772 (O_1772,N_14843,N_14904);
nor UO_1773 (O_1773,N_14934,N_14899);
xor UO_1774 (O_1774,N_14840,N_14800);
nand UO_1775 (O_1775,N_14835,N_14853);
or UO_1776 (O_1776,N_14934,N_14864);
or UO_1777 (O_1777,N_14816,N_14857);
nor UO_1778 (O_1778,N_14822,N_14903);
or UO_1779 (O_1779,N_14939,N_14833);
or UO_1780 (O_1780,N_14808,N_14810);
nand UO_1781 (O_1781,N_14850,N_14994);
xnor UO_1782 (O_1782,N_14975,N_14869);
and UO_1783 (O_1783,N_14932,N_14910);
and UO_1784 (O_1784,N_14824,N_14927);
or UO_1785 (O_1785,N_14888,N_14889);
nand UO_1786 (O_1786,N_14887,N_14944);
or UO_1787 (O_1787,N_14834,N_14848);
and UO_1788 (O_1788,N_14843,N_14821);
or UO_1789 (O_1789,N_14900,N_14821);
xor UO_1790 (O_1790,N_14901,N_14916);
nor UO_1791 (O_1791,N_14909,N_14990);
or UO_1792 (O_1792,N_14840,N_14893);
and UO_1793 (O_1793,N_14881,N_14979);
and UO_1794 (O_1794,N_14924,N_14943);
and UO_1795 (O_1795,N_14959,N_14898);
xor UO_1796 (O_1796,N_14824,N_14851);
xnor UO_1797 (O_1797,N_14905,N_14976);
and UO_1798 (O_1798,N_14857,N_14888);
or UO_1799 (O_1799,N_14976,N_14869);
nand UO_1800 (O_1800,N_14877,N_14935);
xnor UO_1801 (O_1801,N_14849,N_14930);
and UO_1802 (O_1802,N_14989,N_14992);
or UO_1803 (O_1803,N_14958,N_14872);
and UO_1804 (O_1804,N_14977,N_14933);
nand UO_1805 (O_1805,N_14869,N_14968);
nand UO_1806 (O_1806,N_14949,N_14816);
and UO_1807 (O_1807,N_14891,N_14846);
or UO_1808 (O_1808,N_14853,N_14804);
and UO_1809 (O_1809,N_14837,N_14981);
and UO_1810 (O_1810,N_14851,N_14949);
or UO_1811 (O_1811,N_14938,N_14823);
xor UO_1812 (O_1812,N_14851,N_14842);
and UO_1813 (O_1813,N_14801,N_14934);
and UO_1814 (O_1814,N_14941,N_14936);
nand UO_1815 (O_1815,N_14884,N_14880);
and UO_1816 (O_1816,N_14800,N_14977);
or UO_1817 (O_1817,N_14926,N_14899);
xnor UO_1818 (O_1818,N_14859,N_14930);
and UO_1819 (O_1819,N_14898,N_14848);
or UO_1820 (O_1820,N_14867,N_14973);
nand UO_1821 (O_1821,N_14907,N_14979);
nand UO_1822 (O_1822,N_14931,N_14857);
and UO_1823 (O_1823,N_14912,N_14844);
xnor UO_1824 (O_1824,N_14947,N_14913);
nor UO_1825 (O_1825,N_14970,N_14819);
nor UO_1826 (O_1826,N_14825,N_14907);
nor UO_1827 (O_1827,N_14995,N_14903);
and UO_1828 (O_1828,N_14905,N_14919);
nor UO_1829 (O_1829,N_14974,N_14940);
xor UO_1830 (O_1830,N_14984,N_14865);
and UO_1831 (O_1831,N_14938,N_14928);
or UO_1832 (O_1832,N_14985,N_14862);
and UO_1833 (O_1833,N_14871,N_14946);
nor UO_1834 (O_1834,N_14950,N_14998);
nand UO_1835 (O_1835,N_14814,N_14935);
nand UO_1836 (O_1836,N_14878,N_14861);
or UO_1837 (O_1837,N_14812,N_14943);
xor UO_1838 (O_1838,N_14849,N_14843);
xnor UO_1839 (O_1839,N_14821,N_14959);
or UO_1840 (O_1840,N_14944,N_14838);
nand UO_1841 (O_1841,N_14928,N_14898);
nand UO_1842 (O_1842,N_14897,N_14885);
nand UO_1843 (O_1843,N_14918,N_14922);
nor UO_1844 (O_1844,N_14985,N_14843);
or UO_1845 (O_1845,N_14822,N_14824);
nand UO_1846 (O_1846,N_14885,N_14896);
or UO_1847 (O_1847,N_14905,N_14803);
nand UO_1848 (O_1848,N_14943,N_14984);
xnor UO_1849 (O_1849,N_14898,N_14889);
xor UO_1850 (O_1850,N_14952,N_14897);
or UO_1851 (O_1851,N_14848,N_14830);
nand UO_1852 (O_1852,N_14825,N_14943);
or UO_1853 (O_1853,N_14841,N_14992);
nor UO_1854 (O_1854,N_14953,N_14812);
nand UO_1855 (O_1855,N_14953,N_14851);
nand UO_1856 (O_1856,N_14967,N_14866);
nor UO_1857 (O_1857,N_14978,N_14809);
and UO_1858 (O_1858,N_14889,N_14975);
nor UO_1859 (O_1859,N_14852,N_14964);
xor UO_1860 (O_1860,N_14933,N_14824);
nand UO_1861 (O_1861,N_14905,N_14867);
and UO_1862 (O_1862,N_14848,N_14976);
xnor UO_1863 (O_1863,N_14935,N_14888);
nor UO_1864 (O_1864,N_14836,N_14861);
nor UO_1865 (O_1865,N_14880,N_14826);
and UO_1866 (O_1866,N_14983,N_14894);
or UO_1867 (O_1867,N_14896,N_14888);
nor UO_1868 (O_1868,N_14941,N_14970);
or UO_1869 (O_1869,N_14826,N_14849);
nand UO_1870 (O_1870,N_14895,N_14882);
xor UO_1871 (O_1871,N_14985,N_14848);
xnor UO_1872 (O_1872,N_14864,N_14828);
xnor UO_1873 (O_1873,N_14836,N_14962);
nor UO_1874 (O_1874,N_14914,N_14877);
nor UO_1875 (O_1875,N_14898,N_14979);
xor UO_1876 (O_1876,N_14913,N_14921);
nand UO_1877 (O_1877,N_14864,N_14931);
xnor UO_1878 (O_1878,N_14988,N_14818);
or UO_1879 (O_1879,N_14937,N_14880);
and UO_1880 (O_1880,N_14899,N_14891);
nand UO_1881 (O_1881,N_14972,N_14890);
and UO_1882 (O_1882,N_14966,N_14849);
xor UO_1883 (O_1883,N_14848,N_14989);
or UO_1884 (O_1884,N_14900,N_14960);
or UO_1885 (O_1885,N_14924,N_14998);
and UO_1886 (O_1886,N_14855,N_14836);
nor UO_1887 (O_1887,N_14896,N_14870);
and UO_1888 (O_1888,N_14990,N_14838);
and UO_1889 (O_1889,N_14915,N_14875);
xor UO_1890 (O_1890,N_14824,N_14905);
or UO_1891 (O_1891,N_14872,N_14921);
nor UO_1892 (O_1892,N_14891,N_14936);
nand UO_1893 (O_1893,N_14995,N_14933);
and UO_1894 (O_1894,N_14924,N_14933);
nand UO_1895 (O_1895,N_14842,N_14812);
nor UO_1896 (O_1896,N_14936,N_14914);
xor UO_1897 (O_1897,N_14880,N_14926);
nor UO_1898 (O_1898,N_14947,N_14894);
nand UO_1899 (O_1899,N_14925,N_14859);
nor UO_1900 (O_1900,N_14829,N_14975);
or UO_1901 (O_1901,N_14850,N_14847);
or UO_1902 (O_1902,N_14835,N_14863);
or UO_1903 (O_1903,N_14850,N_14879);
nand UO_1904 (O_1904,N_14928,N_14994);
or UO_1905 (O_1905,N_14873,N_14917);
xor UO_1906 (O_1906,N_14935,N_14867);
nor UO_1907 (O_1907,N_14833,N_14968);
nand UO_1908 (O_1908,N_14969,N_14948);
or UO_1909 (O_1909,N_14859,N_14839);
nand UO_1910 (O_1910,N_14972,N_14822);
nor UO_1911 (O_1911,N_14816,N_14811);
nand UO_1912 (O_1912,N_14841,N_14996);
or UO_1913 (O_1913,N_14941,N_14928);
nor UO_1914 (O_1914,N_14909,N_14865);
or UO_1915 (O_1915,N_14908,N_14885);
nor UO_1916 (O_1916,N_14815,N_14951);
or UO_1917 (O_1917,N_14932,N_14838);
and UO_1918 (O_1918,N_14852,N_14896);
and UO_1919 (O_1919,N_14815,N_14950);
and UO_1920 (O_1920,N_14857,N_14871);
nand UO_1921 (O_1921,N_14806,N_14820);
or UO_1922 (O_1922,N_14812,N_14913);
or UO_1923 (O_1923,N_14866,N_14988);
and UO_1924 (O_1924,N_14844,N_14899);
nand UO_1925 (O_1925,N_14804,N_14893);
nor UO_1926 (O_1926,N_14969,N_14886);
nand UO_1927 (O_1927,N_14948,N_14954);
xnor UO_1928 (O_1928,N_14804,N_14993);
and UO_1929 (O_1929,N_14948,N_14961);
and UO_1930 (O_1930,N_14842,N_14950);
xor UO_1931 (O_1931,N_14916,N_14888);
nor UO_1932 (O_1932,N_14996,N_14809);
xnor UO_1933 (O_1933,N_14849,N_14898);
nand UO_1934 (O_1934,N_14896,N_14882);
xnor UO_1935 (O_1935,N_14891,N_14809);
or UO_1936 (O_1936,N_14926,N_14843);
xor UO_1937 (O_1937,N_14800,N_14991);
or UO_1938 (O_1938,N_14992,N_14931);
nand UO_1939 (O_1939,N_14902,N_14873);
nand UO_1940 (O_1940,N_14875,N_14820);
xor UO_1941 (O_1941,N_14974,N_14968);
xor UO_1942 (O_1942,N_14881,N_14805);
and UO_1943 (O_1943,N_14939,N_14827);
and UO_1944 (O_1944,N_14975,N_14906);
nor UO_1945 (O_1945,N_14826,N_14983);
nor UO_1946 (O_1946,N_14936,N_14975);
or UO_1947 (O_1947,N_14894,N_14829);
nand UO_1948 (O_1948,N_14931,N_14800);
nor UO_1949 (O_1949,N_14968,N_14809);
nand UO_1950 (O_1950,N_14928,N_14803);
xnor UO_1951 (O_1951,N_14959,N_14804);
and UO_1952 (O_1952,N_14922,N_14912);
nor UO_1953 (O_1953,N_14957,N_14953);
nand UO_1954 (O_1954,N_14954,N_14830);
nor UO_1955 (O_1955,N_14870,N_14999);
xor UO_1956 (O_1956,N_14850,N_14906);
or UO_1957 (O_1957,N_14803,N_14929);
and UO_1958 (O_1958,N_14853,N_14882);
nand UO_1959 (O_1959,N_14931,N_14819);
nand UO_1960 (O_1960,N_14971,N_14941);
and UO_1961 (O_1961,N_14815,N_14908);
nand UO_1962 (O_1962,N_14995,N_14821);
xnor UO_1963 (O_1963,N_14878,N_14931);
or UO_1964 (O_1964,N_14956,N_14928);
nor UO_1965 (O_1965,N_14875,N_14924);
or UO_1966 (O_1966,N_14816,N_14998);
xnor UO_1967 (O_1967,N_14985,N_14869);
nand UO_1968 (O_1968,N_14858,N_14976);
nand UO_1969 (O_1969,N_14850,N_14917);
and UO_1970 (O_1970,N_14811,N_14914);
and UO_1971 (O_1971,N_14875,N_14966);
nor UO_1972 (O_1972,N_14824,N_14812);
xor UO_1973 (O_1973,N_14943,N_14838);
nor UO_1974 (O_1974,N_14934,N_14888);
or UO_1975 (O_1975,N_14883,N_14858);
or UO_1976 (O_1976,N_14839,N_14977);
nand UO_1977 (O_1977,N_14884,N_14846);
or UO_1978 (O_1978,N_14839,N_14953);
nand UO_1979 (O_1979,N_14950,N_14926);
or UO_1980 (O_1980,N_14924,N_14945);
nand UO_1981 (O_1981,N_14945,N_14806);
nor UO_1982 (O_1982,N_14837,N_14940);
nor UO_1983 (O_1983,N_14986,N_14962);
xor UO_1984 (O_1984,N_14804,N_14901);
nor UO_1985 (O_1985,N_14997,N_14832);
and UO_1986 (O_1986,N_14820,N_14895);
nor UO_1987 (O_1987,N_14869,N_14972);
nor UO_1988 (O_1988,N_14857,N_14890);
xnor UO_1989 (O_1989,N_14839,N_14986);
nor UO_1990 (O_1990,N_14894,N_14826);
nor UO_1991 (O_1991,N_14903,N_14939);
and UO_1992 (O_1992,N_14986,N_14843);
or UO_1993 (O_1993,N_14884,N_14974);
nand UO_1994 (O_1994,N_14842,N_14961);
xor UO_1995 (O_1995,N_14830,N_14952);
and UO_1996 (O_1996,N_14904,N_14897);
xor UO_1997 (O_1997,N_14952,N_14845);
nand UO_1998 (O_1998,N_14904,N_14952);
and UO_1999 (O_1999,N_14957,N_14831);
endmodule