module basic_750_5000_1000_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_96,In_444);
xnor U1 (N_1,In_655,In_59);
or U2 (N_2,In_698,In_659);
xor U3 (N_3,In_195,In_592);
nand U4 (N_4,In_161,In_368);
xnor U5 (N_5,In_653,In_610);
nand U6 (N_6,In_572,In_372);
or U7 (N_7,In_640,In_329);
nand U8 (N_8,In_309,In_646);
nor U9 (N_9,In_304,In_109);
or U10 (N_10,In_259,In_31);
and U11 (N_11,In_136,In_39);
and U12 (N_12,In_94,In_322);
or U13 (N_13,In_582,In_686);
nor U14 (N_14,In_101,In_250);
nand U15 (N_15,In_164,In_268);
nand U16 (N_16,In_615,In_605);
or U17 (N_17,In_564,In_670);
nand U18 (N_18,In_117,In_201);
xnor U19 (N_19,In_194,In_350);
or U20 (N_20,In_104,In_599);
nand U21 (N_21,In_383,In_699);
nand U22 (N_22,In_489,In_251);
xor U23 (N_23,In_513,In_86);
and U24 (N_24,In_330,In_139);
or U25 (N_25,In_666,In_531);
nor U26 (N_26,In_651,In_622);
nand U27 (N_27,In_38,In_0);
or U28 (N_28,In_275,In_456);
and U29 (N_29,In_281,In_256);
nand U30 (N_30,In_393,In_714);
or U31 (N_31,In_517,In_518);
nor U32 (N_32,In_515,In_709);
and U33 (N_33,In_265,In_108);
or U34 (N_34,In_432,In_665);
nand U35 (N_35,In_574,In_362);
xor U36 (N_36,In_213,In_124);
or U37 (N_37,In_723,In_143);
or U38 (N_38,In_371,In_676);
and U39 (N_39,In_591,In_70);
xor U40 (N_40,In_335,In_370);
xnor U41 (N_41,In_618,In_697);
nand U42 (N_42,In_21,In_742);
or U43 (N_43,In_80,In_211);
nand U44 (N_44,In_293,In_332);
or U45 (N_45,In_272,In_155);
xnor U46 (N_46,In_50,In_392);
or U47 (N_47,In_118,In_289);
or U48 (N_48,In_707,In_431);
nand U49 (N_49,In_713,In_316);
nand U50 (N_50,In_246,In_604);
nor U51 (N_51,In_342,In_214);
nand U52 (N_52,In_637,In_9);
or U53 (N_53,In_299,In_29);
nor U54 (N_54,In_89,In_354);
xnor U55 (N_55,In_650,In_282);
xor U56 (N_56,In_166,In_380);
xnor U57 (N_57,In_427,In_516);
and U58 (N_58,In_398,In_730);
xnor U59 (N_59,In_310,In_84);
xnor U60 (N_60,In_349,In_638);
and U61 (N_61,In_486,In_46);
or U62 (N_62,In_381,In_588);
and U63 (N_63,In_173,In_336);
and U64 (N_64,In_583,In_216);
or U65 (N_65,In_594,In_656);
and U66 (N_66,In_99,In_401);
or U67 (N_67,In_684,In_154);
nor U68 (N_68,In_276,In_673);
and U69 (N_69,In_125,In_77);
nor U70 (N_70,In_478,In_505);
nand U71 (N_71,In_128,In_508);
or U72 (N_72,In_327,In_253);
and U73 (N_73,In_185,In_127);
and U74 (N_74,In_577,In_473);
nand U75 (N_75,In_247,In_437);
nor U76 (N_76,In_641,In_262);
nand U77 (N_77,In_123,In_140);
and U78 (N_78,In_150,In_306);
nor U79 (N_79,In_187,In_132);
nor U80 (N_80,In_345,In_716);
nor U81 (N_81,In_667,In_603);
nor U82 (N_82,In_25,In_3);
nand U83 (N_83,In_727,In_578);
or U84 (N_84,In_511,In_79);
or U85 (N_85,In_720,In_303);
nand U86 (N_86,In_643,In_28);
or U87 (N_87,In_729,In_191);
nor U88 (N_88,In_151,In_204);
nand U89 (N_89,In_521,In_743);
xor U90 (N_90,In_722,In_545);
and U91 (N_91,In_365,In_43);
xnor U92 (N_92,In_543,In_134);
nor U93 (N_93,In_55,In_7);
and U94 (N_94,In_424,In_333);
nor U95 (N_95,In_560,In_584);
nand U96 (N_96,In_47,In_248);
or U97 (N_97,In_343,In_319);
nor U98 (N_98,In_174,In_644);
nand U99 (N_99,In_170,In_355);
xor U100 (N_100,In_26,In_103);
and U101 (N_101,In_748,In_307);
nand U102 (N_102,In_664,In_575);
or U103 (N_103,In_446,N_3);
nand U104 (N_104,In_146,In_744);
nand U105 (N_105,In_606,N_69);
xor U106 (N_106,In_657,In_189);
or U107 (N_107,In_220,In_110);
and U108 (N_108,In_274,In_325);
and U109 (N_109,In_224,In_404);
xnor U110 (N_110,In_179,In_454);
nor U111 (N_111,In_130,In_376);
nand U112 (N_112,In_559,In_106);
and U113 (N_113,N_85,In_739);
xor U114 (N_114,In_426,In_529);
xnor U115 (N_115,N_33,In_193);
nor U116 (N_116,N_89,In_416);
nor U117 (N_117,In_704,In_37);
xnor U118 (N_118,In_514,In_557);
or U119 (N_119,In_694,In_595);
nand U120 (N_120,In_76,In_300);
nor U121 (N_121,In_361,In_4);
xor U122 (N_122,N_1,N_50);
and U123 (N_123,In_226,In_159);
xnor U124 (N_124,N_64,In_339);
xnor U125 (N_125,In_10,In_176);
and U126 (N_126,N_32,In_425);
nor U127 (N_127,In_600,In_409);
and U128 (N_128,In_620,N_67);
or U129 (N_129,In_535,In_662);
xor U130 (N_130,In_227,In_242);
xor U131 (N_131,In_597,In_477);
and U132 (N_132,N_35,In_51);
nor U133 (N_133,In_135,In_741);
and U134 (N_134,In_196,In_200);
nand U135 (N_135,In_612,N_22);
or U136 (N_136,In_617,In_54);
and U137 (N_137,N_72,In_616);
nor U138 (N_138,In_255,In_504);
or U139 (N_139,N_82,In_702);
nand U140 (N_140,N_58,N_13);
and U141 (N_141,In_573,In_467);
and U142 (N_142,In_296,N_55);
xor U143 (N_143,In_126,In_749);
and U144 (N_144,In_232,In_692);
xor U145 (N_145,In_453,N_93);
or U146 (N_146,N_90,N_2);
xnor U147 (N_147,In_510,In_369);
and U148 (N_148,In_62,In_88);
or U149 (N_149,In_405,In_602);
and U150 (N_150,In_225,In_280);
xor U151 (N_151,In_311,In_223);
or U152 (N_152,In_169,In_415);
or U153 (N_153,In_447,In_593);
nor U154 (N_154,In_399,In_206);
xnor U155 (N_155,In_131,In_679);
nor U156 (N_156,In_721,In_484);
xor U157 (N_157,In_495,In_210);
or U158 (N_158,In_114,N_29);
and U159 (N_159,In_279,In_480);
nor U160 (N_160,In_178,In_147);
xor U161 (N_161,In_229,In_555);
nand U162 (N_162,In_121,In_563);
nor U163 (N_163,In_526,In_388);
nand U164 (N_164,In_56,In_61);
or U165 (N_165,In_540,N_5);
nor U166 (N_166,In_683,In_737);
nand U167 (N_167,N_95,N_21);
or U168 (N_168,In_724,In_156);
nor U169 (N_169,In_693,In_261);
or U170 (N_170,In_718,N_74);
nand U171 (N_171,In_423,In_298);
nand U172 (N_172,In_462,In_435);
nand U173 (N_173,In_465,N_15);
nand U174 (N_174,In_44,In_351);
xnor U175 (N_175,In_358,In_421);
or U176 (N_176,In_534,In_337);
nor U177 (N_177,In_690,In_119);
or U178 (N_178,N_6,In_522);
or U179 (N_179,In_550,In_115);
xnor U180 (N_180,In_341,In_158);
or U181 (N_181,In_418,N_59);
nand U182 (N_182,In_202,In_496);
xor U183 (N_183,N_96,In_288);
nor U184 (N_184,In_53,N_79);
nor U185 (N_185,In_252,In_429);
or U186 (N_186,In_182,In_263);
nor U187 (N_187,In_218,In_314);
nand U188 (N_188,In_162,In_685);
nand U189 (N_189,N_19,In_579);
and U190 (N_190,In_344,In_317);
or U191 (N_191,N_94,In_19);
nand U192 (N_192,In_661,In_553);
nand U193 (N_193,In_257,N_63);
and U194 (N_194,In_634,N_54);
xnor U195 (N_195,N_99,In_241);
nor U196 (N_196,In_363,N_36);
nand U197 (N_197,In_738,In_377);
nor U198 (N_198,N_88,In_561);
nand U199 (N_199,In_41,In_340);
or U200 (N_200,In_209,N_156);
nor U201 (N_201,In_687,In_623);
nand U202 (N_202,N_151,N_147);
nor U203 (N_203,In_611,In_285);
and U204 (N_204,In_523,In_601);
or U205 (N_205,In_481,In_621);
or U206 (N_206,In_541,N_117);
nor U207 (N_207,In_221,N_150);
or U208 (N_208,N_119,In_414);
nand U209 (N_209,N_145,In_493);
and U210 (N_210,In_375,In_558);
and U211 (N_211,N_191,In_566);
xnor U212 (N_212,N_62,In_649);
nand U213 (N_213,In_458,In_323);
xor U214 (N_214,In_576,N_73);
nand U215 (N_215,N_34,In_17);
or U216 (N_216,In_491,In_474);
or U217 (N_217,In_501,In_706);
nor U218 (N_218,N_17,In_30);
and U219 (N_219,In_144,In_113);
nor U220 (N_220,N_71,N_27);
nor U221 (N_221,In_449,In_149);
xor U222 (N_222,In_745,In_15);
nand U223 (N_223,In_569,In_287);
xor U224 (N_224,In_348,In_5);
and U225 (N_225,N_52,In_273);
and U226 (N_226,In_494,N_126);
or U227 (N_227,N_47,In_387);
xnor U228 (N_228,In_530,In_525);
or U229 (N_229,In_292,In_471);
nand U230 (N_230,N_24,In_466);
and U231 (N_231,In_439,In_452);
nor U232 (N_232,In_18,In_509);
nand U233 (N_233,In_177,In_461);
or U234 (N_234,In_502,In_445);
nor U235 (N_235,In_11,In_645);
nor U236 (N_236,In_45,In_22);
or U237 (N_237,In_313,In_36);
nand U238 (N_238,In_234,In_556);
or U239 (N_239,N_49,In_290);
and U240 (N_240,In_442,In_192);
nand U241 (N_241,In_608,In_688);
or U242 (N_242,In_485,In_283);
nand U243 (N_243,N_157,In_712);
nor U244 (N_244,In_152,In_199);
xor U245 (N_245,In_674,N_190);
and U246 (N_246,N_115,N_51);
or U247 (N_247,N_83,N_178);
or U248 (N_248,In_717,In_407);
nor U249 (N_249,N_109,In_705);
nor U250 (N_250,In_347,In_675);
nand U251 (N_251,N_8,In_65);
nand U252 (N_252,In_448,In_98);
nand U253 (N_253,N_187,In_14);
or U254 (N_254,N_175,In_73);
nand U255 (N_255,In_165,N_101);
or U256 (N_256,In_105,In_180);
or U257 (N_257,In_613,N_77);
nand U258 (N_258,In_72,In_506);
or U259 (N_259,In_527,In_270);
and U260 (N_260,In_16,N_38);
or U261 (N_261,In_367,N_7);
xor U262 (N_262,In_297,N_118);
xnor U263 (N_263,In_436,In_689);
and U264 (N_264,In_122,In_428);
nand U265 (N_265,In_291,In_116);
or U266 (N_266,In_237,N_184);
or U267 (N_267,In_228,In_512);
and U268 (N_268,N_105,N_172);
xnor U269 (N_269,In_548,In_57);
nand U270 (N_270,In_324,In_52);
xor U271 (N_271,In_490,In_32);
xor U272 (N_272,In_410,N_68);
nand U273 (N_273,In_732,In_747);
nand U274 (N_274,In_395,In_81);
nor U275 (N_275,In_654,In_107);
xor U276 (N_276,In_148,In_635);
nor U277 (N_277,In_532,N_131);
nor U278 (N_278,In_389,In_631);
and U279 (N_279,In_48,In_172);
nand U280 (N_280,In_492,N_152);
or U281 (N_281,In_364,In_519);
xnor U282 (N_282,In_546,In_138);
and U283 (N_283,N_170,In_205);
and U284 (N_284,In_78,N_194);
and U285 (N_285,In_391,In_668);
and U286 (N_286,N_199,In_451);
or U287 (N_287,In_691,N_142);
nor U288 (N_288,In_642,N_41);
or U289 (N_289,In_598,In_459);
and U290 (N_290,N_169,N_174);
nand U291 (N_291,N_140,In_190);
and U292 (N_292,In_207,N_165);
or U293 (N_293,N_25,N_197);
xor U294 (N_294,In_483,In_286);
nor U295 (N_295,In_500,In_567);
or U296 (N_296,In_648,In_671);
nor U297 (N_297,In_547,In_85);
nand U298 (N_298,In_681,In_479);
or U299 (N_299,In_538,In_625);
nor U300 (N_300,In_353,In_639);
xor U301 (N_301,N_297,N_205);
and U302 (N_302,In_396,N_220);
and U303 (N_303,In_295,N_159);
nor U304 (N_304,In_528,In_168);
or U305 (N_305,In_82,In_633);
nand U306 (N_306,N_291,In_69);
or U307 (N_307,N_149,In_6);
xnor U308 (N_308,N_243,In_696);
and U309 (N_309,In_91,In_27);
nor U310 (N_310,In_33,In_142);
xor U311 (N_311,In_64,N_75);
or U312 (N_312,In_590,In_422);
and U313 (N_313,In_312,N_137);
xnor U314 (N_314,In_596,N_251);
nand U315 (N_315,In_507,In_302);
nor U316 (N_316,N_86,N_12);
nand U317 (N_317,N_133,N_211);
xnor U318 (N_318,N_70,N_136);
or U319 (N_319,N_244,In_320);
nand U320 (N_320,In_740,N_273);
and U321 (N_321,In_34,N_295);
or U322 (N_322,In_629,N_222);
or U323 (N_323,In_384,In_586);
xnor U324 (N_324,In_520,In_258);
and U325 (N_325,N_164,In_544);
nand U326 (N_326,In_678,N_293);
or U327 (N_327,In_562,In_475);
nor U328 (N_328,In_95,N_264);
nand U329 (N_329,N_188,In_539);
and U330 (N_330,In_20,In_609);
nand U331 (N_331,In_284,In_470);
or U332 (N_332,In_542,In_163);
and U333 (N_333,In_267,N_183);
nor U334 (N_334,In_412,In_408);
nand U335 (N_335,N_252,In_708);
nand U336 (N_336,In_400,N_277);
or U337 (N_337,In_331,In_269);
nand U338 (N_338,N_114,N_221);
nand U339 (N_339,N_250,N_110);
nor U340 (N_340,N_223,In_93);
xor U341 (N_341,In_266,In_663);
nor U342 (N_342,In_239,In_403);
nor U343 (N_343,N_176,In_360);
and U344 (N_344,N_299,In_497);
nor U345 (N_345,In_554,In_321);
or U346 (N_346,N_177,N_37);
or U347 (N_347,N_229,In_12);
and U348 (N_348,N_40,In_188);
xnor U349 (N_349,In_397,N_241);
nand U350 (N_350,N_160,N_14);
xor U351 (N_351,N_10,In_183);
xnor U352 (N_352,In_587,N_285);
nand U353 (N_353,In_24,N_228);
nand U354 (N_354,In_90,N_60);
nand U355 (N_355,In_733,N_216);
nand U356 (N_356,In_102,N_39);
xnor U357 (N_357,In_167,N_97);
xnor U358 (N_358,N_130,N_100);
nand U359 (N_359,N_143,In_695);
and U360 (N_360,In_570,N_76);
xnor U361 (N_361,In_672,In_301);
nand U362 (N_362,In_40,N_255);
xor U363 (N_363,In_464,In_243);
and U364 (N_364,N_45,In_476);
or U365 (N_365,In_413,N_181);
nand U366 (N_366,N_78,N_168);
nand U367 (N_367,N_209,In_208);
or U368 (N_368,In_133,N_43);
or U369 (N_369,In_580,In_682);
nor U370 (N_370,N_290,N_265);
xnor U371 (N_371,N_166,In_334);
or U372 (N_372,N_270,N_20);
nand U373 (N_373,In_420,N_230);
or U374 (N_374,N_107,In_565);
nand U375 (N_375,In_157,N_203);
xnor U376 (N_376,In_619,N_148);
or U377 (N_377,N_44,N_233);
xor U378 (N_378,N_284,In_215);
nand U379 (N_379,In_66,N_261);
nor U380 (N_380,N_0,N_196);
xnor U381 (N_381,In_378,N_127);
and U382 (N_382,In_245,In_472);
xor U383 (N_383,N_298,N_245);
xnor U384 (N_384,In_411,In_254);
and U385 (N_385,In_524,N_11);
and U386 (N_386,N_289,In_87);
nor U387 (N_387,In_92,N_260);
nand U388 (N_388,In_549,N_281);
and U389 (N_389,N_218,In_100);
nand U390 (N_390,N_212,In_315);
and U391 (N_391,In_735,N_53);
or U392 (N_392,N_238,In_503);
nand U393 (N_393,In_628,In_1);
nor U394 (N_394,In_129,N_206);
xnor U395 (N_395,In_203,N_288);
nor U396 (N_396,In_438,N_154);
xnor U397 (N_397,In_441,In_374);
and U398 (N_398,In_719,In_328);
xor U399 (N_399,In_746,N_57);
and U400 (N_400,N_31,N_65);
xor U401 (N_401,N_207,N_9);
or U402 (N_402,N_268,N_302);
nand U403 (N_403,N_314,In_726);
or U404 (N_404,N_87,N_227);
nand U405 (N_405,N_198,N_388);
or U406 (N_406,N_329,In_457);
or U407 (N_407,N_278,N_310);
nor U408 (N_408,N_201,N_210);
or U409 (N_409,In_482,N_316);
nor U410 (N_410,In_552,N_121);
xnor U411 (N_411,N_326,N_353);
or U412 (N_412,In_294,In_240);
nor U413 (N_413,N_276,In_137);
xnor U414 (N_414,N_320,N_269);
and U415 (N_415,N_4,In_352);
and U416 (N_416,In_731,N_340);
nor U417 (N_417,N_236,In_305);
or U418 (N_418,N_249,In_184);
nor U419 (N_419,N_279,In_233);
nor U420 (N_420,N_327,In_463);
nand U421 (N_421,N_129,N_371);
nor U422 (N_422,N_347,N_373);
nor U423 (N_423,In_60,N_263);
nor U424 (N_424,N_385,In_181);
or U425 (N_425,In_487,In_624);
and U426 (N_426,N_372,In_589);
and U427 (N_427,In_145,N_381);
nand U428 (N_428,In_63,N_18);
and U429 (N_429,N_204,N_397);
nor U430 (N_430,In_198,N_23);
and U431 (N_431,In_68,N_56);
nor U432 (N_432,In_498,N_376);
nand U433 (N_433,N_259,N_274);
xnor U434 (N_434,N_173,N_306);
or U435 (N_435,N_189,N_239);
or U436 (N_436,In_468,In_715);
or U437 (N_437,N_319,N_305);
nor U438 (N_438,In_571,N_167);
nand U439 (N_439,N_186,In_366);
and U440 (N_440,In_359,N_363);
or U441 (N_441,N_98,N_337);
and U442 (N_442,N_124,N_358);
nor U443 (N_443,In_551,N_308);
nor U444 (N_444,In_212,In_734);
or U445 (N_445,In_585,In_677);
nand U446 (N_446,N_345,In_278);
nand U447 (N_447,In_175,N_339);
xor U448 (N_448,In_402,In_443);
xor U449 (N_449,N_360,N_392);
and U450 (N_450,N_362,N_309);
nand U451 (N_451,In_680,In_230);
or U452 (N_452,N_283,In_499);
nand U453 (N_453,N_179,N_365);
nor U454 (N_454,In_607,N_355);
nand U455 (N_455,In_308,N_272);
and U456 (N_456,N_224,N_61);
xor U457 (N_457,In_244,In_222);
xor U458 (N_458,N_158,N_342);
nand U459 (N_459,N_366,N_301);
or U460 (N_460,N_346,N_359);
or U461 (N_461,N_113,N_348);
or U462 (N_462,N_102,In_736);
nand U463 (N_463,N_247,N_161);
or U464 (N_464,N_374,In_23);
xor U465 (N_465,In_235,N_399);
nor U466 (N_466,N_344,In_217);
nor U467 (N_467,N_394,N_379);
or U468 (N_468,In_160,N_248);
nor U469 (N_469,N_208,N_328);
nand U470 (N_470,N_391,N_390);
xor U471 (N_471,In_271,In_630);
or U472 (N_472,N_300,N_334);
nor U473 (N_473,In_669,N_296);
nand U474 (N_474,In_74,N_120);
nor U475 (N_475,N_387,In_260);
nor U476 (N_476,N_123,In_249);
or U477 (N_477,N_304,In_186);
and U478 (N_478,In_373,In_701);
nand U479 (N_479,In_469,In_700);
xnor U480 (N_480,N_370,N_317);
nor U481 (N_481,In_632,N_341);
or U482 (N_482,N_106,N_349);
nand U483 (N_483,N_215,N_253);
and U484 (N_484,N_144,N_343);
nand U485 (N_485,N_280,N_84);
nand U486 (N_486,In_430,N_315);
xor U487 (N_487,In_417,In_346);
nand U488 (N_488,N_398,In_433);
xor U489 (N_489,In_49,N_313);
or U490 (N_490,N_232,In_710);
nor U491 (N_491,In_390,N_377);
and U492 (N_492,In_385,N_384);
and U493 (N_493,N_219,N_330);
nand U494 (N_494,N_271,N_323);
xor U495 (N_495,N_389,N_146);
and U496 (N_496,In_326,N_294);
xnor U497 (N_497,N_16,In_197);
nand U498 (N_498,In_357,N_262);
and U499 (N_499,In_636,N_258);
nor U500 (N_500,N_322,N_66);
and U501 (N_501,In_338,N_481);
nand U502 (N_502,N_350,N_457);
xor U503 (N_503,In_627,N_292);
nor U504 (N_504,In_111,N_240);
nor U505 (N_505,N_420,N_336);
xnor U506 (N_506,N_80,N_482);
xor U507 (N_507,N_335,In_141);
or U508 (N_508,N_138,In_318);
xor U509 (N_509,N_408,In_13);
nor U510 (N_510,In_75,N_367);
or U511 (N_511,N_498,In_382);
or U512 (N_512,In_406,In_450);
xnor U513 (N_513,N_111,N_386);
or U514 (N_514,N_477,In_386);
nand U515 (N_515,N_266,N_437);
and U516 (N_516,N_242,N_333);
and U517 (N_517,N_202,N_473);
and U518 (N_518,N_476,In_455);
and U519 (N_519,N_368,N_321);
nor U520 (N_520,N_338,N_369);
nand U521 (N_521,N_405,In_35);
nor U522 (N_522,In_440,N_450);
nor U523 (N_523,N_487,N_485);
or U524 (N_524,N_332,N_122);
nor U525 (N_525,N_419,In_58);
and U526 (N_526,N_382,N_471);
xor U527 (N_527,In_728,N_441);
nand U528 (N_528,N_467,N_162);
nand U529 (N_529,N_423,N_234);
and U530 (N_530,N_286,N_312);
or U531 (N_531,In_626,N_424);
nor U532 (N_532,In_277,N_445);
and U533 (N_533,N_492,N_403);
nand U534 (N_534,N_185,N_451);
nand U535 (N_535,N_378,N_182);
xor U536 (N_536,N_303,N_478);
nor U537 (N_537,N_429,In_171);
and U538 (N_538,N_422,N_354);
xnor U539 (N_539,In_8,In_356);
or U540 (N_540,N_488,N_410);
xnor U541 (N_541,N_400,N_417);
xnor U542 (N_542,N_103,N_416);
and U543 (N_543,N_491,N_46);
nand U544 (N_544,In_71,N_108);
xor U545 (N_545,N_396,N_395);
nor U546 (N_546,N_447,N_472);
or U547 (N_547,N_427,In_703);
xnor U548 (N_548,N_494,In_97);
nand U549 (N_549,In_660,N_225);
nand U550 (N_550,N_455,In_647);
or U551 (N_551,N_104,N_383);
nand U552 (N_552,N_128,N_446);
nand U553 (N_553,N_325,N_463);
nand U554 (N_554,In_238,N_267);
or U555 (N_555,N_461,N_195);
xnor U556 (N_556,In_568,N_42);
nand U557 (N_557,In_652,N_351);
nor U558 (N_558,N_428,In_112);
nand U559 (N_559,N_483,N_421);
nor U560 (N_560,N_434,N_307);
and U561 (N_561,N_406,In_236);
and U562 (N_562,N_438,N_432);
and U563 (N_563,N_480,N_356);
nor U564 (N_564,In_711,N_246);
or U565 (N_565,In_67,N_499);
nand U566 (N_566,N_217,N_444);
nor U567 (N_567,N_415,N_214);
nor U568 (N_568,N_401,N_407);
xor U569 (N_569,N_490,N_496);
or U570 (N_570,N_213,N_484);
nor U571 (N_571,In_231,In_536);
xor U572 (N_572,N_466,N_393);
nor U573 (N_573,N_171,N_364);
nor U574 (N_574,In_614,N_440);
xnor U575 (N_575,N_155,N_470);
nand U576 (N_576,N_453,N_331);
or U577 (N_577,N_91,In_153);
nand U578 (N_578,N_26,N_28);
nand U579 (N_579,N_442,N_235);
nor U580 (N_580,N_464,N_116);
or U581 (N_581,N_112,N_237);
and U582 (N_582,In_537,In_264);
nand U583 (N_583,N_380,In_42);
or U584 (N_584,N_493,N_436);
or U585 (N_585,In_120,N_448);
nor U586 (N_586,N_192,N_409);
xor U587 (N_587,N_486,N_254);
nor U588 (N_588,N_352,N_460);
nor U589 (N_589,In_533,N_200);
and U590 (N_590,N_231,N_431);
xor U591 (N_591,N_92,In_394);
nand U592 (N_592,N_361,N_282);
xnor U593 (N_593,N_357,N_414);
xnor U594 (N_594,N_139,N_452);
nor U595 (N_595,In_581,In_219);
and U596 (N_596,N_430,N_443);
nand U597 (N_597,In_725,In_83);
nor U598 (N_598,N_411,N_454);
and U599 (N_599,N_449,In_419);
nor U600 (N_600,N_574,N_531);
and U601 (N_601,N_582,N_536);
or U602 (N_602,N_551,N_565);
nand U603 (N_603,N_543,N_527);
nand U604 (N_604,N_489,In_434);
xnor U605 (N_605,N_509,N_404);
xor U606 (N_606,N_311,N_30);
nand U607 (N_607,N_587,N_81);
xnor U608 (N_608,N_557,N_180);
nor U609 (N_609,N_465,N_193);
nor U610 (N_610,N_458,N_584);
nand U611 (N_611,N_596,N_501);
and U612 (N_612,N_497,N_530);
xnor U613 (N_613,N_598,N_514);
xor U614 (N_614,N_583,N_418);
and U615 (N_615,N_541,N_537);
xnor U616 (N_616,N_581,N_570);
xnor U617 (N_617,N_456,In_2);
nand U618 (N_618,N_132,N_586);
nand U619 (N_619,N_577,N_426);
nor U620 (N_620,N_545,In_658);
xor U621 (N_621,N_375,N_535);
nand U622 (N_622,N_564,N_469);
nand U623 (N_623,N_529,N_544);
nor U624 (N_624,N_516,N_568);
and U625 (N_625,N_562,N_589);
nor U626 (N_626,N_546,N_226);
and U627 (N_627,N_513,N_502);
nor U628 (N_628,N_507,N_573);
or U629 (N_629,N_519,N_558);
xor U630 (N_630,N_578,N_538);
nor U631 (N_631,N_534,N_561);
xnor U632 (N_632,N_528,N_125);
nand U633 (N_633,In_488,N_505);
nor U634 (N_634,N_591,N_402);
or U635 (N_635,N_504,N_542);
and U636 (N_636,N_522,N_433);
and U637 (N_637,N_495,N_135);
nor U638 (N_638,N_517,N_318);
nor U639 (N_639,N_518,N_163);
nand U640 (N_640,N_512,N_588);
nand U641 (N_641,N_503,N_566);
nor U642 (N_642,N_547,N_552);
or U643 (N_643,N_468,N_287);
and U644 (N_644,N_569,N_462);
and U645 (N_645,N_257,N_475);
xnor U646 (N_646,N_520,N_555);
xnor U647 (N_647,N_153,N_576);
xor U648 (N_648,N_525,N_593);
xnor U649 (N_649,N_590,In_460);
nor U650 (N_650,N_539,N_533);
and U651 (N_651,N_549,N_592);
or U652 (N_652,In_379,N_585);
and U653 (N_653,N_567,N_256);
xnor U654 (N_654,N_413,N_508);
nand U655 (N_655,N_579,N_559);
and U656 (N_656,N_439,N_515);
and U657 (N_657,N_134,N_506);
xnor U658 (N_658,N_599,N_553);
nand U659 (N_659,N_575,N_523);
and U660 (N_660,N_510,N_141);
and U661 (N_661,N_435,N_532);
or U662 (N_662,N_324,N_554);
or U663 (N_663,N_556,N_540);
and U664 (N_664,N_595,N_425);
xnor U665 (N_665,N_474,N_412);
and U666 (N_666,N_459,N_524);
xor U667 (N_667,N_563,N_580);
xor U668 (N_668,N_572,N_594);
or U669 (N_669,N_48,N_597);
nor U670 (N_670,N_479,N_571);
nand U671 (N_671,N_550,N_526);
and U672 (N_672,N_548,N_560);
nor U673 (N_673,N_521,N_500);
nor U674 (N_674,N_275,N_511);
nand U675 (N_675,N_462,N_535);
xor U676 (N_676,N_532,N_81);
nand U677 (N_677,N_597,N_537);
and U678 (N_678,N_588,N_501);
or U679 (N_679,N_595,N_505);
nand U680 (N_680,N_30,N_507);
xor U681 (N_681,N_479,N_520);
nor U682 (N_682,N_597,N_575);
nor U683 (N_683,N_226,N_554);
or U684 (N_684,N_599,N_425);
and U685 (N_685,N_549,N_580);
and U686 (N_686,N_287,N_567);
nand U687 (N_687,N_542,N_134);
nand U688 (N_688,N_518,In_460);
xnor U689 (N_689,N_439,N_561);
xnor U690 (N_690,N_596,N_570);
xnor U691 (N_691,N_564,N_132);
xor U692 (N_692,N_571,N_468);
xor U693 (N_693,N_563,N_459);
nor U694 (N_694,N_531,N_497);
or U695 (N_695,N_501,N_599);
nor U696 (N_696,N_529,N_586);
or U697 (N_697,In_488,N_141);
xnor U698 (N_698,N_553,N_507);
nand U699 (N_699,N_599,N_535);
or U700 (N_700,N_624,N_668);
and U701 (N_701,N_618,N_637);
xor U702 (N_702,N_654,N_653);
nand U703 (N_703,N_687,N_684);
nor U704 (N_704,N_673,N_667);
xor U705 (N_705,N_699,N_671);
xor U706 (N_706,N_609,N_632);
or U707 (N_707,N_614,N_688);
nand U708 (N_708,N_613,N_666);
nor U709 (N_709,N_607,N_651);
and U710 (N_710,N_694,N_693);
nor U711 (N_711,N_600,N_625);
or U712 (N_712,N_674,N_626);
nand U713 (N_713,N_663,N_675);
nand U714 (N_714,N_658,N_647);
nand U715 (N_715,N_603,N_644);
nor U716 (N_716,N_605,N_616);
xnor U717 (N_717,N_682,N_611);
nand U718 (N_718,N_652,N_606);
xnor U719 (N_719,N_617,N_610);
nand U720 (N_720,N_638,N_623);
xor U721 (N_721,N_696,N_665);
nand U722 (N_722,N_620,N_612);
nand U723 (N_723,N_669,N_659);
nor U724 (N_724,N_698,N_628);
nand U725 (N_725,N_629,N_630);
nand U726 (N_726,N_622,N_641);
nor U727 (N_727,N_642,N_608);
xor U728 (N_728,N_615,N_692);
xnor U729 (N_729,N_672,N_686);
nor U730 (N_730,N_627,N_639);
nand U731 (N_731,N_661,N_660);
and U732 (N_732,N_646,N_601);
and U733 (N_733,N_636,N_604);
nor U734 (N_734,N_640,N_635);
nand U735 (N_735,N_650,N_655);
nand U736 (N_736,N_679,N_697);
nor U737 (N_737,N_649,N_695);
or U738 (N_738,N_621,N_670);
nor U739 (N_739,N_645,N_676);
nand U740 (N_740,N_680,N_631);
or U741 (N_741,N_690,N_648);
xor U742 (N_742,N_634,N_691);
nor U743 (N_743,N_619,N_685);
or U744 (N_744,N_657,N_677);
nand U745 (N_745,N_689,N_662);
nand U746 (N_746,N_683,N_678);
or U747 (N_747,N_681,N_664);
and U748 (N_748,N_633,N_602);
nand U749 (N_749,N_656,N_643);
xnor U750 (N_750,N_653,N_604);
and U751 (N_751,N_694,N_656);
nor U752 (N_752,N_651,N_685);
nand U753 (N_753,N_658,N_657);
and U754 (N_754,N_622,N_660);
nand U755 (N_755,N_699,N_690);
nand U756 (N_756,N_658,N_640);
xnor U757 (N_757,N_667,N_652);
xor U758 (N_758,N_685,N_652);
or U759 (N_759,N_635,N_678);
and U760 (N_760,N_694,N_687);
or U761 (N_761,N_681,N_619);
xor U762 (N_762,N_691,N_612);
or U763 (N_763,N_621,N_623);
nor U764 (N_764,N_654,N_642);
and U765 (N_765,N_613,N_640);
nor U766 (N_766,N_637,N_673);
xnor U767 (N_767,N_642,N_618);
or U768 (N_768,N_666,N_667);
and U769 (N_769,N_635,N_634);
xnor U770 (N_770,N_669,N_671);
nand U771 (N_771,N_683,N_699);
xor U772 (N_772,N_625,N_640);
xnor U773 (N_773,N_660,N_633);
or U774 (N_774,N_678,N_605);
xor U775 (N_775,N_653,N_634);
xor U776 (N_776,N_626,N_634);
and U777 (N_777,N_646,N_683);
xnor U778 (N_778,N_666,N_692);
or U779 (N_779,N_642,N_643);
nor U780 (N_780,N_610,N_698);
xor U781 (N_781,N_688,N_605);
or U782 (N_782,N_679,N_611);
and U783 (N_783,N_668,N_623);
or U784 (N_784,N_643,N_617);
and U785 (N_785,N_630,N_648);
or U786 (N_786,N_632,N_655);
xnor U787 (N_787,N_665,N_644);
xor U788 (N_788,N_631,N_673);
xnor U789 (N_789,N_605,N_640);
or U790 (N_790,N_617,N_675);
or U791 (N_791,N_655,N_681);
and U792 (N_792,N_670,N_615);
and U793 (N_793,N_679,N_606);
xor U794 (N_794,N_694,N_671);
or U795 (N_795,N_652,N_624);
nor U796 (N_796,N_674,N_618);
or U797 (N_797,N_627,N_615);
nand U798 (N_798,N_685,N_635);
nor U799 (N_799,N_627,N_676);
xor U800 (N_800,N_727,N_737);
xor U801 (N_801,N_762,N_763);
or U802 (N_802,N_768,N_709);
nand U803 (N_803,N_793,N_720);
xor U804 (N_804,N_767,N_743);
xnor U805 (N_805,N_723,N_745);
and U806 (N_806,N_794,N_717);
and U807 (N_807,N_738,N_719);
and U808 (N_808,N_755,N_790);
nor U809 (N_809,N_778,N_729);
nor U810 (N_810,N_740,N_787);
or U811 (N_811,N_775,N_779);
xor U812 (N_812,N_749,N_735);
nand U813 (N_813,N_707,N_782);
nand U814 (N_814,N_726,N_744);
nor U815 (N_815,N_747,N_785);
or U816 (N_816,N_757,N_780);
nor U817 (N_817,N_784,N_716);
or U818 (N_818,N_711,N_789);
nor U819 (N_819,N_713,N_730);
or U820 (N_820,N_774,N_725);
nor U821 (N_821,N_764,N_792);
nand U822 (N_822,N_786,N_753);
nor U823 (N_823,N_751,N_760);
xor U824 (N_824,N_776,N_773);
nor U825 (N_825,N_731,N_708);
nor U826 (N_826,N_791,N_777);
xnor U827 (N_827,N_718,N_756);
or U828 (N_828,N_736,N_722);
and U829 (N_829,N_703,N_712);
and U830 (N_830,N_758,N_734);
xnor U831 (N_831,N_795,N_781);
xnor U832 (N_832,N_799,N_701);
nor U833 (N_833,N_752,N_797);
nor U834 (N_834,N_705,N_728);
xor U835 (N_835,N_715,N_704);
xor U836 (N_836,N_742,N_761);
xnor U837 (N_837,N_721,N_770);
nor U838 (N_838,N_714,N_765);
or U839 (N_839,N_771,N_733);
nand U840 (N_840,N_710,N_702);
and U841 (N_841,N_732,N_700);
nor U842 (N_842,N_766,N_739);
or U843 (N_843,N_788,N_748);
nand U844 (N_844,N_754,N_759);
or U845 (N_845,N_741,N_798);
nand U846 (N_846,N_750,N_783);
nor U847 (N_847,N_724,N_796);
xor U848 (N_848,N_769,N_772);
nor U849 (N_849,N_706,N_746);
xor U850 (N_850,N_739,N_744);
nand U851 (N_851,N_792,N_725);
nor U852 (N_852,N_759,N_707);
xor U853 (N_853,N_748,N_759);
or U854 (N_854,N_780,N_775);
nand U855 (N_855,N_788,N_789);
nor U856 (N_856,N_797,N_784);
and U857 (N_857,N_739,N_700);
nand U858 (N_858,N_740,N_723);
nor U859 (N_859,N_755,N_763);
nor U860 (N_860,N_725,N_766);
and U861 (N_861,N_712,N_777);
and U862 (N_862,N_705,N_776);
nor U863 (N_863,N_737,N_723);
and U864 (N_864,N_717,N_705);
xor U865 (N_865,N_773,N_775);
and U866 (N_866,N_740,N_783);
xor U867 (N_867,N_725,N_740);
or U868 (N_868,N_795,N_785);
nand U869 (N_869,N_783,N_763);
nand U870 (N_870,N_706,N_789);
nor U871 (N_871,N_793,N_764);
or U872 (N_872,N_759,N_722);
or U873 (N_873,N_700,N_764);
and U874 (N_874,N_781,N_798);
xnor U875 (N_875,N_734,N_701);
and U876 (N_876,N_791,N_708);
and U877 (N_877,N_720,N_715);
and U878 (N_878,N_726,N_708);
xor U879 (N_879,N_709,N_704);
or U880 (N_880,N_743,N_797);
and U881 (N_881,N_732,N_701);
xor U882 (N_882,N_761,N_752);
or U883 (N_883,N_746,N_712);
xor U884 (N_884,N_751,N_769);
or U885 (N_885,N_734,N_775);
xor U886 (N_886,N_758,N_771);
nand U887 (N_887,N_724,N_788);
nor U888 (N_888,N_759,N_736);
nor U889 (N_889,N_702,N_714);
nor U890 (N_890,N_737,N_732);
and U891 (N_891,N_765,N_790);
nor U892 (N_892,N_754,N_777);
xor U893 (N_893,N_701,N_710);
nand U894 (N_894,N_773,N_779);
nand U895 (N_895,N_776,N_788);
or U896 (N_896,N_755,N_789);
or U897 (N_897,N_701,N_748);
nor U898 (N_898,N_733,N_734);
xnor U899 (N_899,N_713,N_790);
xor U900 (N_900,N_880,N_838);
nor U901 (N_901,N_887,N_889);
xnor U902 (N_902,N_897,N_803);
nand U903 (N_903,N_869,N_845);
and U904 (N_904,N_823,N_854);
or U905 (N_905,N_834,N_878);
nor U906 (N_906,N_873,N_892);
nand U907 (N_907,N_886,N_847);
nand U908 (N_908,N_885,N_837);
nor U909 (N_909,N_839,N_804);
and U910 (N_910,N_816,N_835);
or U911 (N_911,N_875,N_810);
xor U912 (N_912,N_884,N_852);
and U913 (N_913,N_891,N_822);
nor U914 (N_914,N_824,N_801);
nor U915 (N_915,N_846,N_865);
or U916 (N_916,N_841,N_836);
nor U917 (N_917,N_861,N_876);
xnor U918 (N_918,N_871,N_853);
and U919 (N_919,N_855,N_868);
xor U920 (N_920,N_879,N_849);
and U921 (N_921,N_820,N_800);
and U922 (N_922,N_833,N_888);
nand U923 (N_923,N_893,N_856);
or U924 (N_924,N_831,N_867);
or U925 (N_925,N_842,N_883);
xor U926 (N_926,N_840,N_830);
nand U927 (N_927,N_811,N_848);
nor U928 (N_928,N_877,N_894);
xnor U929 (N_929,N_806,N_826);
xnor U930 (N_930,N_857,N_890);
or U931 (N_931,N_815,N_870);
or U932 (N_932,N_812,N_828);
or U933 (N_933,N_863,N_898);
xor U934 (N_934,N_896,N_808);
nand U935 (N_935,N_858,N_862);
nor U936 (N_936,N_850,N_805);
nor U937 (N_937,N_860,N_807);
nor U938 (N_938,N_813,N_899);
and U939 (N_939,N_881,N_819);
nand U940 (N_940,N_814,N_872);
and U941 (N_941,N_802,N_882);
nor U942 (N_942,N_866,N_825);
nand U943 (N_943,N_809,N_832);
nor U944 (N_944,N_821,N_827);
nor U945 (N_945,N_864,N_895);
and U946 (N_946,N_859,N_874);
xnor U947 (N_947,N_829,N_818);
nor U948 (N_948,N_844,N_851);
or U949 (N_949,N_843,N_817);
and U950 (N_950,N_869,N_883);
or U951 (N_951,N_800,N_860);
or U952 (N_952,N_873,N_837);
nor U953 (N_953,N_844,N_864);
nor U954 (N_954,N_811,N_858);
nor U955 (N_955,N_897,N_863);
nor U956 (N_956,N_822,N_885);
and U957 (N_957,N_861,N_893);
or U958 (N_958,N_816,N_851);
or U959 (N_959,N_843,N_873);
xor U960 (N_960,N_844,N_898);
nor U961 (N_961,N_834,N_811);
nand U962 (N_962,N_854,N_828);
xor U963 (N_963,N_817,N_884);
nand U964 (N_964,N_822,N_843);
nor U965 (N_965,N_881,N_869);
or U966 (N_966,N_890,N_838);
nand U967 (N_967,N_812,N_810);
xor U968 (N_968,N_899,N_833);
and U969 (N_969,N_822,N_816);
and U970 (N_970,N_831,N_800);
nor U971 (N_971,N_814,N_845);
or U972 (N_972,N_867,N_830);
nand U973 (N_973,N_886,N_858);
and U974 (N_974,N_821,N_866);
xnor U975 (N_975,N_808,N_826);
nand U976 (N_976,N_887,N_842);
or U977 (N_977,N_806,N_885);
and U978 (N_978,N_838,N_809);
xnor U979 (N_979,N_858,N_850);
and U980 (N_980,N_868,N_853);
nor U981 (N_981,N_817,N_872);
xor U982 (N_982,N_813,N_850);
and U983 (N_983,N_875,N_871);
or U984 (N_984,N_824,N_873);
or U985 (N_985,N_834,N_839);
nor U986 (N_986,N_828,N_805);
or U987 (N_987,N_872,N_822);
nand U988 (N_988,N_841,N_855);
and U989 (N_989,N_894,N_819);
or U990 (N_990,N_829,N_887);
nor U991 (N_991,N_833,N_854);
nor U992 (N_992,N_864,N_889);
xnor U993 (N_993,N_837,N_877);
and U994 (N_994,N_879,N_869);
xnor U995 (N_995,N_859,N_817);
xnor U996 (N_996,N_861,N_888);
nor U997 (N_997,N_825,N_850);
and U998 (N_998,N_892,N_883);
xnor U999 (N_999,N_841,N_816);
and U1000 (N_1000,N_977,N_957);
or U1001 (N_1001,N_994,N_928);
nand U1002 (N_1002,N_904,N_914);
xnor U1003 (N_1003,N_921,N_954);
xnor U1004 (N_1004,N_970,N_980);
nand U1005 (N_1005,N_925,N_965);
or U1006 (N_1006,N_968,N_915);
or U1007 (N_1007,N_963,N_975);
nor U1008 (N_1008,N_910,N_976);
or U1009 (N_1009,N_930,N_929);
or U1010 (N_1010,N_916,N_958);
nor U1011 (N_1011,N_985,N_993);
xor U1012 (N_1012,N_919,N_999);
xor U1013 (N_1013,N_991,N_966);
and U1014 (N_1014,N_920,N_982);
or U1015 (N_1015,N_992,N_949);
nor U1016 (N_1016,N_947,N_946);
nand U1017 (N_1017,N_937,N_981);
nand U1018 (N_1018,N_997,N_911);
nand U1019 (N_1019,N_940,N_951);
and U1020 (N_1020,N_955,N_990);
nor U1021 (N_1021,N_979,N_901);
nor U1022 (N_1022,N_972,N_969);
xor U1023 (N_1023,N_909,N_987);
nor U1024 (N_1024,N_971,N_917);
xor U1025 (N_1025,N_944,N_922);
nand U1026 (N_1026,N_907,N_996);
nor U1027 (N_1027,N_945,N_903);
or U1028 (N_1028,N_936,N_933);
or U1029 (N_1029,N_995,N_927);
xor U1030 (N_1030,N_932,N_902);
xnor U1031 (N_1031,N_923,N_918);
nand U1032 (N_1032,N_988,N_934);
or U1033 (N_1033,N_984,N_964);
or U1034 (N_1034,N_939,N_908);
xor U1035 (N_1035,N_989,N_941);
or U1036 (N_1036,N_900,N_926);
xnor U1037 (N_1037,N_931,N_953);
xnor U1038 (N_1038,N_924,N_986);
nor U1039 (N_1039,N_978,N_906);
nand U1040 (N_1040,N_913,N_998);
xnor U1041 (N_1041,N_938,N_942);
xnor U1042 (N_1042,N_974,N_961);
nor U1043 (N_1043,N_956,N_973);
xor U1044 (N_1044,N_943,N_935);
xor U1045 (N_1045,N_905,N_952);
and U1046 (N_1046,N_983,N_950);
and U1047 (N_1047,N_959,N_962);
or U1048 (N_1048,N_960,N_912);
and U1049 (N_1049,N_948,N_967);
nor U1050 (N_1050,N_940,N_930);
and U1051 (N_1051,N_912,N_949);
nor U1052 (N_1052,N_967,N_901);
or U1053 (N_1053,N_947,N_974);
nand U1054 (N_1054,N_989,N_924);
nand U1055 (N_1055,N_903,N_909);
nor U1056 (N_1056,N_907,N_989);
or U1057 (N_1057,N_932,N_964);
nor U1058 (N_1058,N_985,N_995);
nand U1059 (N_1059,N_987,N_922);
or U1060 (N_1060,N_989,N_975);
or U1061 (N_1061,N_904,N_929);
nand U1062 (N_1062,N_997,N_928);
and U1063 (N_1063,N_966,N_906);
xnor U1064 (N_1064,N_983,N_968);
or U1065 (N_1065,N_922,N_951);
xnor U1066 (N_1066,N_908,N_986);
nor U1067 (N_1067,N_966,N_932);
xnor U1068 (N_1068,N_982,N_909);
and U1069 (N_1069,N_977,N_933);
xor U1070 (N_1070,N_902,N_922);
nand U1071 (N_1071,N_922,N_901);
nor U1072 (N_1072,N_974,N_906);
xor U1073 (N_1073,N_963,N_971);
nand U1074 (N_1074,N_913,N_934);
nand U1075 (N_1075,N_954,N_989);
or U1076 (N_1076,N_998,N_912);
nor U1077 (N_1077,N_980,N_908);
or U1078 (N_1078,N_942,N_928);
xnor U1079 (N_1079,N_975,N_956);
and U1080 (N_1080,N_981,N_965);
nand U1081 (N_1081,N_915,N_974);
and U1082 (N_1082,N_948,N_989);
or U1083 (N_1083,N_917,N_989);
nor U1084 (N_1084,N_999,N_959);
or U1085 (N_1085,N_922,N_945);
and U1086 (N_1086,N_910,N_925);
or U1087 (N_1087,N_991,N_925);
or U1088 (N_1088,N_991,N_990);
xnor U1089 (N_1089,N_917,N_943);
or U1090 (N_1090,N_981,N_901);
nand U1091 (N_1091,N_979,N_958);
or U1092 (N_1092,N_959,N_921);
nor U1093 (N_1093,N_916,N_920);
or U1094 (N_1094,N_903,N_990);
nand U1095 (N_1095,N_926,N_935);
and U1096 (N_1096,N_977,N_904);
nand U1097 (N_1097,N_920,N_980);
or U1098 (N_1098,N_943,N_996);
or U1099 (N_1099,N_948,N_947);
or U1100 (N_1100,N_1021,N_1075);
nor U1101 (N_1101,N_1022,N_1082);
or U1102 (N_1102,N_1097,N_1061);
nand U1103 (N_1103,N_1028,N_1092);
xnor U1104 (N_1104,N_1025,N_1006);
or U1105 (N_1105,N_1089,N_1066);
or U1106 (N_1106,N_1064,N_1001);
nor U1107 (N_1107,N_1019,N_1005);
xor U1108 (N_1108,N_1096,N_1033);
or U1109 (N_1109,N_1091,N_1030);
nor U1110 (N_1110,N_1026,N_1036);
nand U1111 (N_1111,N_1054,N_1002);
or U1112 (N_1112,N_1045,N_1043);
nand U1113 (N_1113,N_1050,N_1098);
and U1114 (N_1114,N_1038,N_1051);
xor U1115 (N_1115,N_1067,N_1027);
nand U1116 (N_1116,N_1053,N_1017);
or U1117 (N_1117,N_1073,N_1081);
and U1118 (N_1118,N_1049,N_1069);
xnor U1119 (N_1119,N_1085,N_1056);
or U1120 (N_1120,N_1088,N_1057);
and U1121 (N_1121,N_1046,N_1065);
and U1122 (N_1122,N_1087,N_1035);
or U1123 (N_1123,N_1007,N_1093);
nor U1124 (N_1124,N_1090,N_1048);
or U1125 (N_1125,N_1011,N_1000);
or U1126 (N_1126,N_1059,N_1074);
or U1127 (N_1127,N_1068,N_1037);
nand U1128 (N_1128,N_1063,N_1095);
or U1129 (N_1129,N_1047,N_1080);
nand U1130 (N_1130,N_1083,N_1055);
and U1131 (N_1131,N_1052,N_1084);
nor U1132 (N_1132,N_1023,N_1044);
or U1133 (N_1133,N_1013,N_1072);
nor U1134 (N_1134,N_1016,N_1010);
nand U1135 (N_1135,N_1009,N_1071);
nand U1136 (N_1136,N_1078,N_1014);
nand U1137 (N_1137,N_1004,N_1041);
nor U1138 (N_1138,N_1042,N_1012);
and U1139 (N_1139,N_1099,N_1060);
xor U1140 (N_1140,N_1029,N_1070);
nor U1141 (N_1141,N_1040,N_1018);
xnor U1142 (N_1142,N_1015,N_1020);
xnor U1143 (N_1143,N_1039,N_1079);
xnor U1144 (N_1144,N_1077,N_1058);
and U1145 (N_1145,N_1003,N_1034);
or U1146 (N_1146,N_1094,N_1062);
or U1147 (N_1147,N_1032,N_1031);
or U1148 (N_1148,N_1008,N_1024);
xnor U1149 (N_1149,N_1086,N_1076);
or U1150 (N_1150,N_1005,N_1083);
and U1151 (N_1151,N_1094,N_1011);
and U1152 (N_1152,N_1084,N_1068);
nand U1153 (N_1153,N_1097,N_1057);
nor U1154 (N_1154,N_1041,N_1050);
and U1155 (N_1155,N_1051,N_1065);
or U1156 (N_1156,N_1005,N_1074);
xor U1157 (N_1157,N_1088,N_1074);
nor U1158 (N_1158,N_1050,N_1068);
nand U1159 (N_1159,N_1005,N_1095);
xor U1160 (N_1160,N_1053,N_1019);
xor U1161 (N_1161,N_1084,N_1072);
and U1162 (N_1162,N_1006,N_1044);
and U1163 (N_1163,N_1050,N_1066);
and U1164 (N_1164,N_1081,N_1024);
and U1165 (N_1165,N_1071,N_1012);
nor U1166 (N_1166,N_1060,N_1027);
and U1167 (N_1167,N_1049,N_1076);
nand U1168 (N_1168,N_1017,N_1026);
or U1169 (N_1169,N_1099,N_1098);
and U1170 (N_1170,N_1041,N_1033);
nor U1171 (N_1171,N_1035,N_1053);
nor U1172 (N_1172,N_1086,N_1055);
nand U1173 (N_1173,N_1077,N_1059);
nor U1174 (N_1174,N_1018,N_1006);
or U1175 (N_1175,N_1075,N_1037);
nand U1176 (N_1176,N_1041,N_1017);
nand U1177 (N_1177,N_1008,N_1079);
or U1178 (N_1178,N_1013,N_1014);
nor U1179 (N_1179,N_1094,N_1079);
or U1180 (N_1180,N_1072,N_1095);
nand U1181 (N_1181,N_1010,N_1008);
or U1182 (N_1182,N_1064,N_1073);
xnor U1183 (N_1183,N_1041,N_1053);
nand U1184 (N_1184,N_1050,N_1058);
nor U1185 (N_1185,N_1098,N_1096);
or U1186 (N_1186,N_1003,N_1064);
nand U1187 (N_1187,N_1095,N_1031);
nand U1188 (N_1188,N_1069,N_1048);
xor U1189 (N_1189,N_1039,N_1001);
or U1190 (N_1190,N_1065,N_1061);
xor U1191 (N_1191,N_1005,N_1012);
xor U1192 (N_1192,N_1011,N_1022);
and U1193 (N_1193,N_1098,N_1066);
nand U1194 (N_1194,N_1005,N_1009);
or U1195 (N_1195,N_1050,N_1053);
and U1196 (N_1196,N_1048,N_1009);
xor U1197 (N_1197,N_1027,N_1077);
xnor U1198 (N_1198,N_1087,N_1059);
and U1199 (N_1199,N_1004,N_1023);
nor U1200 (N_1200,N_1195,N_1173);
nor U1201 (N_1201,N_1186,N_1174);
and U1202 (N_1202,N_1177,N_1199);
nand U1203 (N_1203,N_1168,N_1158);
xor U1204 (N_1204,N_1103,N_1191);
or U1205 (N_1205,N_1197,N_1104);
and U1206 (N_1206,N_1156,N_1119);
nand U1207 (N_1207,N_1135,N_1127);
nor U1208 (N_1208,N_1175,N_1171);
nor U1209 (N_1209,N_1159,N_1110);
and U1210 (N_1210,N_1117,N_1193);
and U1211 (N_1211,N_1140,N_1149);
xnor U1212 (N_1212,N_1137,N_1147);
nor U1213 (N_1213,N_1116,N_1170);
or U1214 (N_1214,N_1157,N_1162);
nor U1215 (N_1215,N_1196,N_1112);
and U1216 (N_1216,N_1153,N_1144);
xor U1217 (N_1217,N_1107,N_1181);
nand U1218 (N_1218,N_1188,N_1176);
xnor U1219 (N_1219,N_1120,N_1145);
nand U1220 (N_1220,N_1151,N_1154);
nand U1221 (N_1221,N_1169,N_1136);
and U1222 (N_1222,N_1152,N_1106);
nand U1223 (N_1223,N_1124,N_1185);
nand U1224 (N_1224,N_1161,N_1148);
xnor U1225 (N_1225,N_1190,N_1184);
and U1226 (N_1226,N_1132,N_1101);
or U1227 (N_1227,N_1160,N_1183);
and U1228 (N_1228,N_1138,N_1142);
and U1229 (N_1229,N_1122,N_1133);
nand U1230 (N_1230,N_1114,N_1146);
nand U1231 (N_1231,N_1102,N_1130);
and U1232 (N_1232,N_1198,N_1121);
and U1233 (N_1233,N_1123,N_1194);
and U1234 (N_1234,N_1111,N_1166);
xor U1235 (N_1235,N_1143,N_1192);
nor U1236 (N_1236,N_1167,N_1178);
nor U1237 (N_1237,N_1164,N_1150);
or U1238 (N_1238,N_1165,N_1129);
or U1239 (N_1239,N_1125,N_1100);
and U1240 (N_1240,N_1113,N_1115);
nor U1241 (N_1241,N_1118,N_1105);
and U1242 (N_1242,N_1134,N_1126);
nand U1243 (N_1243,N_1182,N_1187);
nor U1244 (N_1244,N_1180,N_1172);
and U1245 (N_1245,N_1163,N_1179);
or U1246 (N_1246,N_1131,N_1139);
nand U1247 (N_1247,N_1128,N_1155);
and U1248 (N_1248,N_1141,N_1109);
nor U1249 (N_1249,N_1189,N_1108);
nor U1250 (N_1250,N_1160,N_1182);
xnor U1251 (N_1251,N_1133,N_1140);
nand U1252 (N_1252,N_1169,N_1143);
nand U1253 (N_1253,N_1121,N_1199);
nor U1254 (N_1254,N_1152,N_1127);
or U1255 (N_1255,N_1123,N_1122);
nand U1256 (N_1256,N_1170,N_1167);
xnor U1257 (N_1257,N_1160,N_1171);
nand U1258 (N_1258,N_1119,N_1189);
nor U1259 (N_1259,N_1183,N_1152);
or U1260 (N_1260,N_1181,N_1179);
or U1261 (N_1261,N_1149,N_1117);
xnor U1262 (N_1262,N_1124,N_1180);
and U1263 (N_1263,N_1164,N_1119);
xnor U1264 (N_1264,N_1176,N_1192);
nand U1265 (N_1265,N_1193,N_1178);
and U1266 (N_1266,N_1122,N_1186);
nor U1267 (N_1267,N_1162,N_1109);
or U1268 (N_1268,N_1173,N_1150);
or U1269 (N_1269,N_1117,N_1104);
nor U1270 (N_1270,N_1185,N_1171);
nand U1271 (N_1271,N_1198,N_1190);
nor U1272 (N_1272,N_1144,N_1188);
and U1273 (N_1273,N_1135,N_1143);
nand U1274 (N_1274,N_1140,N_1185);
or U1275 (N_1275,N_1176,N_1103);
nand U1276 (N_1276,N_1155,N_1124);
and U1277 (N_1277,N_1107,N_1116);
and U1278 (N_1278,N_1177,N_1108);
nand U1279 (N_1279,N_1190,N_1149);
xnor U1280 (N_1280,N_1105,N_1177);
xnor U1281 (N_1281,N_1196,N_1142);
xor U1282 (N_1282,N_1150,N_1194);
or U1283 (N_1283,N_1114,N_1163);
and U1284 (N_1284,N_1140,N_1127);
and U1285 (N_1285,N_1192,N_1149);
and U1286 (N_1286,N_1174,N_1183);
and U1287 (N_1287,N_1166,N_1159);
nor U1288 (N_1288,N_1185,N_1127);
or U1289 (N_1289,N_1126,N_1117);
nor U1290 (N_1290,N_1153,N_1152);
or U1291 (N_1291,N_1193,N_1132);
or U1292 (N_1292,N_1196,N_1117);
xnor U1293 (N_1293,N_1186,N_1170);
or U1294 (N_1294,N_1184,N_1147);
xnor U1295 (N_1295,N_1153,N_1166);
nand U1296 (N_1296,N_1129,N_1101);
xor U1297 (N_1297,N_1198,N_1154);
and U1298 (N_1298,N_1181,N_1126);
nor U1299 (N_1299,N_1185,N_1113);
or U1300 (N_1300,N_1265,N_1257);
or U1301 (N_1301,N_1250,N_1206);
nand U1302 (N_1302,N_1251,N_1211);
or U1303 (N_1303,N_1231,N_1220);
or U1304 (N_1304,N_1207,N_1237);
and U1305 (N_1305,N_1223,N_1281);
and U1306 (N_1306,N_1238,N_1201);
or U1307 (N_1307,N_1298,N_1268);
or U1308 (N_1308,N_1283,N_1299);
xor U1309 (N_1309,N_1233,N_1285);
or U1310 (N_1310,N_1278,N_1284);
and U1311 (N_1311,N_1255,N_1282);
xor U1312 (N_1312,N_1294,N_1262);
xor U1313 (N_1313,N_1240,N_1208);
or U1314 (N_1314,N_1204,N_1297);
and U1315 (N_1315,N_1225,N_1270);
and U1316 (N_1316,N_1256,N_1286);
or U1317 (N_1317,N_1295,N_1280);
and U1318 (N_1318,N_1269,N_1246);
nand U1319 (N_1319,N_1212,N_1224);
xor U1320 (N_1320,N_1229,N_1239);
nor U1321 (N_1321,N_1273,N_1218);
nand U1322 (N_1322,N_1234,N_1252);
nor U1323 (N_1323,N_1275,N_1259);
or U1324 (N_1324,N_1221,N_1279);
or U1325 (N_1325,N_1244,N_1222);
or U1326 (N_1326,N_1203,N_1202);
nand U1327 (N_1327,N_1287,N_1243);
or U1328 (N_1328,N_1236,N_1277);
or U1329 (N_1329,N_1216,N_1291);
and U1330 (N_1330,N_1272,N_1263);
and U1331 (N_1331,N_1249,N_1253);
or U1332 (N_1332,N_1266,N_1245);
nand U1333 (N_1333,N_1289,N_1267);
nand U1334 (N_1334,N_1290,N_1274);
and U1335 (N_1335,N_1247,N_1213);
xor U1336 (N_1336,N_1219,N_1230);
nand U1337 (N_1337,N_1288,N_1210);
nand U1338 (N_1338,N_1217,N_1232);
nand U1339 (N_1339,N_1264,N_1292);
and U1340 (N_1340,N_1258,N_1293);
nor U1341 (N_1341,N_1235,N_1200);
and U1342 (N_1342,N_1227,N_1209);
and U1343 (N_1343,N_1260,N_1215);
xnor U1344 (N_1344,N_1241,N_1254);
xor U1345 (N_1345,N_1271,N_1276);
xor U1346 (N_1346,N_1242,N_1205);
nor U1347 (N_1347,N_1296,N_1261);
xor U1348 (N_1348,N_1228,N_1214);
xnor U1349 (N_1349,N_1248,N_1226);
nor U1350 (N_1350,N_1238,N_1273);
xnor U1351 (N_1351,N_1239,N_1212);
or U1352 (N_1352,N_1255,N_1278);
xnor U1353 (N_1353,N_1223,N_1274);
and U1354 (N_1354,N_1220,N_1249);
nor U1355 (N_1355,N_1282,N_1206);
nand U1356 (N_1356,N_1274,N_1269);
and U1357 (N_1357,N_1240,N_1260);
nor U1358 (N_1358,N_1257,N_1276);
nand U1359 (N_1359,N_1223,N_1285);
nand U1360 (N_1360,N_1256,N_1269);
or U1361 (N_1361,N_1215,N_1219);
nand U1362 (N_1362,N_1208,N_1242);
and U1363 (N_1363,N_1259,N_1226);
nand U1364 (N_1364,N_1251,N_1225);
nand U1365 (N_1365,N_1264,N_1285);
nand U1366 (N_1366,N_1259,N_1216);
nor U1367 (N_1367,N_1257,N_1253);
xnor U1368 (N_1368,N_1257,N_1228);
nor U1369 (N_1369,N_1258,N_1225);
or U1370 (N_1370,N_1248,N_1228);
nand U1371 (N_1371,N_1268,N_1205);
and U1372 (N_1372,N_1281,N_1237);
xor U1373 (N_1373,N_1248,N_1217);
xor U1374 (N_1374,N_1247,N_1239);
or U1375 (N_1375,N_1214,N_1239);
nor U1376 (N_1376,N_1295,N_1291);
nor U1377 (N_1377,N_1283,N_1291);
xor U1378 (N_1378,N_1211,N_1212);
nor U1379 (N_1379,N_1222,N_1213);
or U1380 (N_1380,N_1248,N_1297);
or U1381 (N_1381,N_1291,N_1253);
nand U1382 (N_1382,N_1271,N_1208);
xnor U1383 (N_1383,N_1281,N_1228);
xnor U1384 (N_1384,N_1221,N_1227);
or U1385 (N_1385,N_1274,N_1237);
or U1386 (N_1386,N_1211,N_1258);
and U1387 (N_1387,N_1209,N_1234);
xnor U1388 (N_1388,N_1245,N_1272);
or U1389 (N_1389,N_1298,N_1239);
xnor U1390 (N_1390,N_1248,N_1271);
nand U1391 (N_1391,N_1240,N_1217);
xnor U1392 (N_1392,N_1230,N_1251);
or U1393 (N_1393,N_1265,N_1284);
xnor U1394 (N_1394,N_1212,N_1264);
xnor U1395 (N_1395,N_1219,N_1284);
nor U1396 (N_1396,N_1236,N_1276);
xor U1397 (N_1397,N_1223,N_1211);
or U1398 (N_1398,N_1221,N_1237);
and U1399 (N_1399,N_1258,N_1252);
nor U1400 (N_1400,N_1329,N_1360);
and U1401 (N_1401,N_1343,N_1386);
nand U1402 (N_1402,N_1350,N_1325);
xor U1403 (N_1403,N_1346,N_1374);
nand U1404 (N_1404,N_1376,N_1341);
and U1405 (N_1405,N_1378,N_1314);
nand U1406 (N_1406,N_1368,N_1308);
or U1407 (N_1407,N_1327,N_1385);
and U1408 (N_1408,N_1348,N_1377);
xor U1409 (N_1409,N_1317,N_1387);
or U1410 (N_1410,N_1357,N_1372);
nor U1411 (N_1411,N_1352,N_1354);
xnor U1412 (N_1412,N_1393,N_1331);
and U1413 (N_1413,N_1303,N_1340);
xnor U1414 (N_1414,N_1306,N_1337);
nand U1415 (N_1415,N_1388,N_1307);
and U1416 (N_1416,N_1355,N_1363);
nand U1417 (N_1417,N_1390,N_1389);
nor U1418 (N_1418,N_1370,N_1358);
and U1419 (N_1419,N_1328,N_1342);
xnor U1420 (N_1420,N_1312,N_1304);
or U1421 (N_1421,N_1361,N_1396);
or U1422 (N_1422,N_1364,N_1332);
nand U1423 (N_1423,N_1399,N_1375);
and U1424 (N_1424,N_1394,N_1300);
nand U1425 (N_1425,N_1339,N_1359);
nand U1426 (N_1426,N_1353,N_1310);
xor U1427 (N_1427,N_1391,N_1336);
xnor U1428 (N_1428,N_1397,N_1323);
nand U1429 (N_1429,N_1302,N_1335);
and U1430 (N_1430,N_1369,N_1320);
and U1431 (N_1431,N_1345,N_1380);
xnor U1432 (N_1432,N_1382,N_1324);
nor U1433 (N_1433,N_1395,N_1373);
and U1434 (N_1434,N_1321,N_1305);
or U1435 (N_1435,N_1381,N_1367);
nor U1436 (N_1436,N_1383,N_1356);
nor U1437 (N_1437,N_1333,N_1315);
or U1438 (N_1438,N_1371,N_1366);
nand U1439 (N_1439,N_1379,N_1398);
and U1440 (N_1440,N_1351,N_1392);
nor U1441 (N_1441,N_1301,N_1318);
nor U1442 (N_1442,N_1311,N_1322);
or U1443 (N_1443,N_1309,N_1384);
or U1444 (N_1444,N_1347,N_1334);
and U1445 (N_1445,N_1316,N_1344);
nand U1446 (N_1446,N_1349,N_1313);
nand U1447 (N_1447,N_1319,N_1362);
and U1448 (N_1448,N_1338,N_1326);
nor U1449 (N_1449,N_1330,N_1365);
nor U1450 (N_1450,N_1370,N_1390);
nor U1451 (N_1451,N_1355,N_1395);
or U1452 (N_1452,N_1334,N_1352);
nand U1453 (N_1453,N_1353,N_1368);
nor U1454 (N_1454,N_1343,N_1361);
nor U1455 (N_1455,N_1313,N_1321);
nand U1456 (N_1456,N_1317,N_1361);
and U1457 (N_1457,N_1370,N_1393);
xor U1458 (N_1458,N_1305,N_1374);
xnor U1459 (N_1459,N_1357,N_1348);
and U1460 (N_1460,N_1374,N_1353);
nor U1461 (N_1461,N_1382,N_1360);
nand U1462 (N_1462,N_1392,N_1324);
nor U1463 (N_1463,N_1307,N_1373);
and U1464 (N_1464,N_1322,N_1366);
and U1465 (N_1465,N_1395,N_1307);
or U1466 (N_1466,N_1305,N_1306);
xnor U1467 (N_1467,N_1320,N_1382);
nor U1468 (N_1468,N_1354,N_1346);
nor U1469 (N_1469,N_1307,N_1326);
nor U1470 (N_1470,N_1335,N_1308);
nand U1471 (N_1471,N_1333,N_1387);
xnor U1472 (N_1472,N_1332,N_1341);
nand U1473 (N_1473,N_1351,N_1336);
nand U1474 (N_1474,N_1395,N_1372);
and U1475 (N_1475,N_1394,N_1374);
or U1476 (N_1476,N_1351,N_1374);
nand U1477 (N_1477,N_1347,N_1377);
xor U1478 (N_1478,N_1368,N_1331);
and U1479 (N_1479,N_1308,N_1323);
or U1480 (N_1480,N_1386,N_1384);
xnor U1481 (N_1481,N_1361,N_1349);
nand U1482 (N_1482,N_1331,N_1310);
nor U1483 (N_1483,N_1367,N_1365);
and U1484 (N_1484,N_1360,N_1385);
xor U1485 (N_1485,N_1337,N_1376);
and U1486 (N_1486,N_1397,N_1316);
nand U1487 (N_1487,N_1339,N_1360);
xor U1488 (N_1488,N_1306,N_1387);
or U1489 (N_1489,N_1376,N_1386);
nor U1490 (N_1490,N_1370,N_1339);
or U1491 (N_1491,N_1372,N_1315);
nor U1492 (N_1492,N_1321,N_1353);
nand U1493 (N_1493,N_1304,N_1369);
and U1494 (N_1494,N_1323,N_1371);
nor U1495 (N_1495,N_1336,N_1373);
nor U1496 (N_1496,N_1306,N_1340);
or U1497 (N_1497,N_1311,N_1349);
nand U1498 (N_1498,N_1374,N_1362);
nor U1499 (N_1499,N_1365,N_1325);
nor U1500 (N_1500,N_1458,N_1461);
xnor U1501 (N_1501,N_1456,N_1472);
and U1502 (N_1502,N_1451,N_1422);
nand U1503 (N_1503,N_1408,N_1490);
xor U1504 (N_1504,N_1444,N_1435);
or U1505 (N_1505,N_1404,N_1427);
nor U1506 (N_1506,N_1480,N_1432);
xnor U1507 (N_1507,N_1453,N_1497);
or U1508 (N_1508,N_1447,N_1406);
and U1509 (N_1509,N_1449,N_1403);
or U1510 (N_1510,N_1411,N_1448);
or U1511 (N_1511,N_1452,N_1487);
and U1512 (N_1512,N_1423,N_1426);
and U1513 (N_1513,N_1481,N_1437);
xnor U1514 (N_1514,N_1474,N_1442);
nor U1515 (N_1515,N_1428,N_1499);
or U1516 (N_1516,N_1464,N_1455);
and U1517 (N_1517,N_1469,N_1483);
nand U1518 (N_1518,N_1482,N_1417);
and U1519 (N_1519,N_1496,N_1471);
xor U1520 (N_1520,N_1475,N_1429);
nor U1521 (N_1521,N_1488,N_1477);
or U1522 (N_1522,N_1454,N_1409);
xor U1523 (N_1523,N_1410,N_1414);
nor U1524 (N_1524,N_1478,N_1465);
and U1525 (N_1525,N_1457,N_1418);
and U1526 (N_1526,N_1425,N_1419);
or U1527 (N_1527,N_1459,N_1443);
xnor U1528 (N_1528,N_1462,N_1493);
xnor U1529 (N_1529,N_1441,N_1420);
xor U1530 (N_1530,N_1486,N_1494);
nor U1531 (N_1531,N_1433,N_1401);
xor U1532 (N_1532,N_1424,N_1491);
xnor U1533 (N_1533,N_1415,N_1402);
or U1534 (N_1534,N_1498,N_1484);
xor U1535 (N_1535,N_1416,N_1492);
xor U1536 (N_1536,N_1430,N_1405);
and U1537 (N_1537,N_1445,N_1413);
and U1538 (N_1538,N_1438,N_1468);
nand U1539 (N_1539,N_1489,N_1421);
xor U1540 (N_1540,N_1470,N_1407);
nand U1541 (N_1541,N_1450,N_1485);
xnor U1542 (N_1542,N_1467,N_1412);
xnor U1543 (N_1543,N_1479,N_1440);
nor U1544 (N_1544,N_1460,N_1400);
and U1545 (N_1545,N_1436,N_1463);
xor U1546 (N_1546,N_1446,N_1431);
nor U1547 (N_1547,N_1495,N_1476);
xnor U1548 (N_1548,N_1439,N_1434);
xnor U1549 (N_1549,N_1466,N_1473);
or U1550 (N_1550,N_1454,N_1466);
xnor U1551 (N_1551,N_1410,N_1422);
nor U1552 (N_1552,N_1487,N_1443);
and U1553 (N_1553,N_1449,N_1423);
and U1554 (N_1554,N_1490,N_1456);
and U1555 (N_1555,N_1461,N_1407);
xnor U1556 (N_1556,N_1422,N_1460);
xnor U1557 (N_1557,N_1440,N_1487);
and U1558 (N_1558,N_1425,N_1400);
and U1559 (N_1559,N_1447,N_1409);
nand U1560 (N_1560,N_1407,N_1439);
nor U1561 (N_1561,N_1407,N_1486);
xnor U1562 (N_1562,N_1402,N_1414);
nor U1563 (N_1563,N_1406,N_1475);
and U1564 (N_1564,N_1440,N_1414);
xnor U1565 (N_1565,N_1422,N_1465);
and U1566 (N_1566,N_1466,N_1448);
xor U1567 (N_1567,N_1477,N_1419);
nand U1568 (N_1568,N_1492,N_1461);
or U1569 (N_1569,N_1448,N_1489);
xnor U1570 (N_1570,N_1460,N_1435);
nor U1571 (N_1571,N_1451,N_1497);
nor U1572 (N_1572,N_1406,N_1456);
nor U1573 (N_1573,N_1417,N_1476);
nand U1574 (N_1574,N_1437,N_1442);
or U1575 (N_1575,N_1403,N_1454);
nand U1576 (N_1576,N_1466,N_1404);
xnor U1577 (N_1577,N_1439,N_1452);
nand U1578 (N_1578,N_1406,N_1412);
nand U1579 (N_1579,N_1471,N_1413);
xor U1580 (N_1580,N_1411,N_1461);
or U1581 (N_1581,N_1448,N_1433);
nor U1582 (N_1582,N_1434,N_1484);
xor U1583 (N_1583,N_1408,N_1409);
and U1584 (N_1584,N_1457,N_1411);
nand U1585 (N_1585,N_1416,N_1423);
and U1586 (N_1586,N_1447,N_1474);
and U1587 (N_1587,N_1433,N_1457);
xor U1588 (N_1588,N_1471,N_1438);
nand U1589 (N_1589,N_1443,N_1494);
nor U1590 (N_1590,N_1423,N_1427);
xor U1591 (N_1591,N_1440,N_1464);
or U1592 (N_1592,N_1421,N_1450);
or U1593 (N_1593,N_1484,N_1464);
nand U1594 (N_1594,N_1467,N_1494);
xnor U1595 (N_1595,N_1434,N_1488);
nor U1596 (N_1596,N_1456,N_1429);
and U1597 (N_1597,N_1420,N_1450);
and U1598 (N_1598,N_1455,N_1412);
nor U1599 (N_1599,N_1450,N_1484);
or U1600 (N_1600,N_1591,N_1529);
or U1601 (N_1601,N_1565,N_1512);
nand U1602 (N_1602,N_1570,N_1545);
nor U1603 (N_1603,N_1509,N_1586);
nor U1604 (N_1604,N_1500,N_1501);
nand U1605 (N_1605,N_1513,N_1550);
nor U1606 (N_1606,N_1525,N_1514);
nor U1607 (N_1607,N_1560,N_1527);
xnor U1608 (N_1608,N_1541,N_1578);
nand U1609 (N_1609,N_1543,N_1532);
xnor U1610 (N_1610,N_1519,N_1597);
xor U1611 (N_1611,N_1576,N_1535);
or U1612 (N_1612,N_1548,N_1510);
and U1613 (N_1613,N_1568,N_1575);
nand U1614 (N_1614,N_1506,N_1544);
xor U1615 (N_1615,N_1562,N_1572);
xor U1616 (N_1616,N_1505,N_1542);
xor U1617 (N_1617,N_1558,N_1502);
nand U1618 (N_1618,N_1553,N_1537);
xor U1619 (N_1619,N_1573,N_1508);
or U1620 (N_1620,N_1540,N_1567);
nor U1621 (N_1621,N_1574,N_1523);
nor U1622 (N_1622,N_1546,N_1584);
or U1623 (N_1623,N_1539,N_1592);
nand U1624 (N_1624,N_1557,N_1590);
nand U1625 (N_1625,N_1595,N_1561);
nand U1626 (N_1626,N_1504,N_1522);
and U1627 (N_1627,N_1533,N_1507);
nor U1628 (N_1628,N_1520,N_1528);
and U1629 (N_1629,N_1538,N_1593);
nor U1630 (N_1630,N_1551,N_1554);
nor U1631 (N_1631,N_1577,N_1549);
and U1632 (N_1632,N_1555,N_1511);
and U1633 (N_1633,N_1582,N_1599);
or U1634 (N_1634,N_1598,N_1559);
nor U1635 (N_1635,N_1534,N_1581);
or U1636 (N_1636,N_1571,N_1563);
and U1637 (N_1637,N_1564,N_1580);
nand U1638 (N_1638,N_1596,N_1588);
nand U1639 (N_1639,N_1517,N_1526);
and U1640 (N_1640,N_1585,N_1530);
xnor U1641 (N_1641,N_1589,N_1515);
or U1642 (N_1642,N_1594,N_1583);
or U1643 (N_1643,N_1516,N_1587);
nor U1644 (N_1644,N_1547,N_1579);
nand U1645 (N_1645,N_1566,N_1552);
xnor U1646 (N_1646,N_1521,N_1524);
nor U1647 (N_1647,N_1536,N_1531);
xnor U1648 (N_1648,N_1518,N_1503);
or U1649 (N_1649,N_1569,N_1556);
nand U1650 (N_1650,N_1520,N_1500);
xor U1651 (N_1651,N_1586,N_1533);
nor U1652 (N_1652,N_1543,N_1566);
or U1653 (N_1653,N_1551,N_1581);
nand U1654 (N_1654,N_1585,N_1511);
or U1655 (N_1655,N_1539,N_1548);
nand U1656 (N_1656,N_1541,N_1573);
nor U1657 (N_1657,N_1567,N_1500);
nor U1658 (N_1658,N_1514,N_1570);
xnor U1659 (N_1659,N_1517,N_1558);
nand U1660 (N_1660,N_1539,N_1513);
nor U1661 (N_1661,N_1591,N_1561);
or U1662 (N_1662,N_1549,N_1587);
and U1663 (N_1663,N_1531,N_1591);
nor U1664 (N_1664,N_1526,N_1565);
nand U1665 (N_1665,N_1561,N_1549);
nand U1666 (N_1666,N_1512,N_1504);
or U1667 (N_1667,N_1515,N_1505);
nor U1668 (N_1668,N_1587,N_1514);
nand U1669 (N_1669,N_1599,N_1588);
xor U1670 (N_1670,N_1536,N_1571);
or U1671 (N_1671,N_1502,N_1509);
nor U1672 (N_1672,N_1535,N_1545);
xor U1673 (N_1673,N_1519,N_1531);
nand U1674 (N_1674,N_1597,N_1595);
nand U1675 (N_1675,N_1554,N_1593);
nor U1676 (N_1676,N_1553,N_1509);
and U1677 (N_1677,N_1580,N_1570);
nor U1678 (N_1678,N_1532,N_1593);
or U1679 (N_1679,N_1549,N_1517);
and U1680 (N_1680,N_1501,N_1551);
or U1681 (N_1681,N_1538,N_1548);
xor U1682 (N_1682,N_1570,N_1556);
and U1683 (N_1683,N_1537,N_1548);
and U1684 (N_1684,N_1584,N_1540);
nor U1685 (N_1685,N_1580,N_1535);
xnor U1686 (N_1686,N_1593,N_1587);
nand U1687 (N_1687,N_1531,N_1565);
nor U1688 (N_1688,N_1544,N_1591);
and U1689 (N_1689,N_1576,N_1514);
nand U1690 (N_1690,N_1569,N_1573);
and U1691 (N_1691,N_1516,N_1572);
nand U1692 (N_1692,N_1578,N_1521);
xnor U1693 (N_1693,N_1544,N_1555);
or U1694 (N_1694,N_1503,N_1522);
and U1695 (N_1695,N_1558,N_1545);
xnor U1696 (N_1696,N_1530,N_1590);
or U1697 (N_1697,N_1506,N_1599);
and U1698 (N_1698,N_1528,N_1534);
nand U1699 (N_1699,N_1575,N_1551);
nand U1700 (N_1700,N_1613,N_1680);
nand U1701 (N_1701,N_1618,N_1619);
nand U1702 (N_1702,N_1651,N_1653);
nor U1703 (N_1703,N_1686,N_1617);
nand U1704 (N_1704,N_1666,N_1667);
and U1705 (N_1705,N_1673,N_1658);
or U1706 (N_1706,N_1638,N_1699);
nor U1707 (N_1707,N_1688,N_1691);
and U1708 (N_1708,N_1676,N_1631);
nand U1709 (N_1709,N_1641,N_1662);
xnor U1710 (N_1710,N_1642,N_1636);
nor U1711 (N_1711,N_1648,N_1603);
xnor U1712 (N_1712,N_1620,N_1633);
and U1713 (N_1713,N_1668,N_1678);
xor U1714 (N_1714,N_1623,N_1692);
and U1715 (N_1715,N_1696,N_1624);
and U1716 (N_1716,N_1665,N_1632);
nand U1717 (N_1717,N_1654,N_1644);
and U1718 (N_1718,N_1616,N_1602);
xnor U1719 (N_1719,N_1647,N_1645);
or U1720 (N_1720,N_1611,N_1625);
xor U1721 (N_1721,N_1697,N_1682);
xnor U1722 (N_1722,N_1612,N_1601);
xnor U1723 (N_1723,N_1640,N_1639);
or U1724 (N_1724,N_1669,N_1609);
nand U1725 (N_1725,N_1693,N_1637);
and U1726 (N_1726,N_1626,N_1670);
nand U1727 (N_1727,N_1674,N_1677);
nor U1728 (N_1728,N_1659,N_1661);
nor U1729 (N_1729,N_1656,N_1605);
xor U1730 (N_1730,N_1675,N_1671);
xor U1731 (N_1731,N_1629,N_1650);
nor U1732 (N_1732,N_1681,N_1679);
nand U1733 (N_1733,N_1690,N_1695);
nand U1734 (N_1734,N_1687,N_1663);
xor U1735 (N_1735,N_1614,N_1622);
nand U1736 (N_1736,N_1635,N_1600);
xnor U1737 (N_1737,N_1606,N_1672);
or U1738 (N_1738,N_1652,N_1615);
nand U1739 (N_1739,N_1610,N_1604);
xor U1740 (N_1740,N_1649,N_1684);
nor U1741 (N_1741,N_1634,N_1657);
or U1742 (N_1742,N_1628,N_1655);
and U1743 (N_1743,N_1607,N_1630);
nor U1744 (N_1744,N_1698,N_1646);
xor U1745 (N_1745,N_1685,N_1643);
nor U1746 (N_1746,N_1608,N_1683);
or U1747 (N_1747,N_1689,N_1694);
nand U1748 (N_1748,N_1660,N_1627);
nand U1749 (N_1749,N_1664,N_1621);
nor U1750 (N_1750,N_1626,N_1654);
and U1751 (N_1751,N_1678,N_1620);
and U1752 (N_1752,N_1610,N_1669);
nand U1753 (N_1753,N_1698,N_1669);
nor U1754 (N_1754,N_1645,N_1634);
or U1755 (N_1755,N_1616,N_1666);
xnor U1756 (N_1756,N_1619,N_1614);
and U1757 (N_1757,N_1680,N_1644);
nand U1758 (N_1758,N_1643,N_1673);
nor U1759 (N_1759,N_1697,N_1618);
or U1760 (N_1760,N_1638,N_1610);
nand U1761 (N_1761,N_1669,N_1614);
xor U1762 (N_1762,N_1684,N_1645);
and U1763 (N_1763,N_1663,N_1678);
xor U1764 (N_1764,N_1609,N_1631);
nand U1765 (N_1765,N_1658,N_1684);
xor U1766 (N_1766,N_1683,N_1673);
nand U1767 (N_1767,N_1623,N_1631);
or U1768 (N_1768,N_1694,N_1623);
and U1769 (N_1769,N_1664,N_1653);
xnor U1770 (N_1770,N_1652,N_1639);
and U1771 (N_1771,N_1665,N_1675);
nand U1772 (N_1772,N_1640,N_1694);
xor U1773 (N_1773,N_1635,N_1610);
nor U1774 (N_1774,N_1686,N_1692);
nor U1775 (N_1775,N_1684,N_1602);
nor U1776 (N_1776,N_1618,N_1603);
and U1777 (N_1777,N_1699,N_1628);
and U1778 (N_1778,N_1693,N_1692);
xor U1779 (N_1779,N_1651,N_1678);
and U1780 (N_1780,N_1619,N_1661);
nand U1781 (N_1781,N_1629,N_1648);
nor U1782 (N_1782,N_1623,N_1607);
and U1783 (N_1783,N_1689,N_1646);
xnor U1784 (N_1784,N_1659,N_1611);
xor U1785 (N_1785,N_1625,N_1676);
xor U1786 (N_1786,N_1657,N_1617);
nand U1787 (N_1787,N_1653,N_1683);
nand U1788 (N_1788,N_1605,N_1640);
xor U1789 (N_1789,N_1614,N_1665);
and U1790 (N_1790,N_1640,N_1632);
and U1791 (N_1791,N_1638,N_1666);
nand U1792 (N_1792,N_1615,N_1626);
nand U1793 (N_1793,N_1648,N_1652);
nand U1794 (N_1794,N_1613,N_1689);
nor U1795 (N_1795,N_1690,N_1642);
and U1796 (N_1796,N_1615,N_1620);
nor U1797 (N_1797,N_1676,N_1623);
nand U1798 (N_1798,N_1657,N_1638);
or U1799 (N_1799,N_1606,N_1677);
xor U1800 (N_1800,N_1761,N_1719);
nor U1801 (N_1801,N_1742,N_1735);
nand U1802 (N_1802,N_1740,N_1751);
and U1803 (N_1803,N_1705,N_1759);
or U1804 (N_1804,N_1711,N_1792);
xnor U1805 (N_1805,N_1793,N_1782);
xor U1806 (N_1806,N_1791,N_1772);
nand U1807 (N_1807,N_1773,N_1790);
nor U1808 (N_1808,N_1744,N_1766);
nand U1809 (N_1809,N_1700,N_1727);
and U1810 (N_1810,N_1722,N_1778);
and U1811 (N_1811,N_1750,N_1713);
xor U1812 (N_1812,N_1752,N_1777);
and U1813 (N_1813,N_1756,N_1754);
nor U1814 (N_1814,N_1734,N_1786);
or U1815 (N_1815,N_1731,N_1724);
and U1816 (N_1816,N_1758,N_1765);
nand U1817 (N_1817,N_1769,N_1798);
nor U1818 (N_1818,N_1764,N_1714);
or U1819 (N_1819,N_1774,N_1755);
or U1820 (N_1820,N_1703,N_1785);
and U1821 (N_1821,N_1712,N_1797);
nand U1822 (N_1822,N_1741,N_1723);
nor U1823 (N_1823,N_1736,N_1757);
xnor U1824 (N_1824,N_1707,N_1732);
or U1825 (N_1825,N_1737,N_1763);
nand U1826 (N_1826,N_1789,N_1771);
nand U1827 (N_1827,N_1781,N_1708);
or U1828 (N_1828,N_1783,N_1702);
xnor U1829 (N_1829,N_1746,N_1720);
xor U1830 (N_1830,N_1775,N_1787);
xor U1831 (N_1831,N_1776,N_1770);
nor U1832 (N_1832,N_1706,N_1717);
nand U1833 (N_1833,N_1784,N_1704);
and U1834 (N_1834,N_1718,N_1795);
and U1835 (N_1835,N_1794,N_1730);
nor U1836 (N_1836,N_1749,N_1738);
nand U1837 (N_1837,N_1780,N_1726);
nand U1838 (N_1838,N_1745,N_1743);
and U1839 (N_1839,N_1739,N_1733);
nor U1840 (N_1840,N_1779,N_1716);
and U1841 (N_1841,N_1725,N_1796);
nor U1842 (N_1842,N_1721,N_1710);
nand U1843 (N_1843,N_1753,N_1709);
nand U1844 (N_1844,N_1762,N_1768);
xnor U1845 (N_1845,N_1747,N_1728);
xnor U1846 (N_1846,N_1715,N_1767);
xnor U1847 (N_1847,N_1729,N_1748);
and U1848 (N_1848,N_1788,N_1701);
and U1849 (N_1849,N_1799,N_1760);
or U1850 (N_1850,N_1714,N_1777);
or U1851 (N_1851,N_1786,N_1785);
nand U1852 (N_1852,N_1707,N_1791);
nor U1853 (N_1853,N_1759,N_1761);
and U1854 (N_1854,N_1772,N_1739);
and U1855 (N_1855,N_1726,N_1773);
xor U1856 (N_1856,N_1760,N_1748);
or U1857 (N_1857,N_1715,N_1738);
nor U1858 (N_1858,N_1757,N_1777);
nand U1859 (N_1859,N_1798,N_1748);
or U1860 (N_1860,N_1798,N_1799);
or U1861 (N_1861,N_1755,N_1788);
and U1862 (N_1862,N_1796,N_1707);
nand U1863 (N_1863,N_1713,N_1777);
nor U1864 (N_1864,N_1736,N_1791);
nand U1865 (N_1865,N_1757,N_1768);
nand U1866 (N_1866,N_1727,N_1711);
or U1867 (N_1867,N_1757,N_1759);
nand U1868 (N_1868,N_1764,N_1750);
and U1869 (N_1869,N_1765,N_1723);
or U1870 (N_1870,N_1753,N_1703);
xnor U1871 (N_1871,N_1717,N_1720);
and U1872 (N_1872,N_1744,N_1764);
nand U1873 (N_1873,N_1740,N_1738);
and U1874 (N_1874,N_1786,N_1772);
and U1875 (N_1875,N_1781,N_1773);
nor U1876 (N_1876,N_1760,N_1738);
nand U1877 (N_1877,N_1753,N_1799);
nor U1878 (N_1878,N_1730,N_1782);
or U1879 (N_1879,N_1791,N_1728);
nor U1880 (N_1880,N_1722,N_1717);
nor U1881 (N_1881,N_1751,N_1756);
nor U1882 (N_1882,N_1778,N_1779);
nor U1883 (N_1883,N_1775,N_1748);
nor U1884 (N_1884,N_1773,N_1711);
nor U1885 (N_1885,N_1724,N_1730);
xnor U1886 (N_1886,N_1749,N_1758);
and U1887 (N_1887,N_1745,N_1742);
and U1888 (N_1888,N_1780,N_1735);
nor U1889 (N_1889,N_1766,N_1794);
nor U1890 (N_1890,N_1726,N_1772);
and U1891 (N_1891,N_1760,N_1767);
and U1892 (N_1892,N_1747,N_1704);
nor U1893 (N_1893,N_1773,N_1737);
xor U1894 (N_1894,N_1731,N_1717);
and U1895 (N_1895,N_1711,N_1736);
nor U1896 (N_1896,N_1731,N_1795);
and U1897 (N_1897,N_1705,N_1750);
and U1898 (N_1898,N_1799,N_1723);
or U1899 (N_1899,N_1756,N_1777);
nor U1900 (N_1900,N_1856,N_1818);
nand U1901 (N_1901,N_1814,N_1822);
xor U1902 (N_1902,N_1870,N_1817);
and U1903 (N_1903,N_1809,N_1805);
and U1904 (N_1904,N_1865,N_1857);
and U1905 (N_1905,N_1868,N_1815);
xor U1906 (N_1906,N_1811,N_1881);
xnor U1907 (N_1907,N_1861,N_1821);
and U1908 (N_1908,N_1883,N_1826);
nor U1909 (N_1909,N_1819,N_1871);
and U1910 (N_1910,N_1807,N_1879);
nor U1911 (N_1911,N_1812,N_1849);
xnor U1912 (N_1912,N_1810,N_1802);
nor U1913 (N_1913,N_1829,N_1867);
or U1914 (N_1914,N_1846,N_1823);
and U1915 (N_1915,N_1882,N_1893);
xnor U1916 (N_1916,N_1813,N_1897);
nand U1917 (N_1917,N_1840,N_1875);
or U1918 (N_1918,N_1877,N_1852);
and U1919 (N_1919,N_1833,N_1848);
xor U1920 (N_1920,N_1844,N_1837);
nor U1921 (N_1921,N_1873,N_1864);
xor U1922 (N_1922,N_1816,N_1851);
and U1923 (N_1923,N_1894,N_1860);
nor U1924 (N_1924,N_1859,N_1843);
and U1925 (N_1925,N_1841,N_1891);
and U1926 (N_1926,N_1880,N_1838);
xnor U1927 (N_1927,N_1804,N_1831);
nand U1928 (N_1928,N_1863,N_1827);
and U1929 (N_1929,N_1801,N_1820);
and U1930 (N_1930,N_1853,N_1806);
nor U1931 (N_1931,N_1854,N_1892);
xnor U1932 (N_1932,N_1872,N_1836);
xnor U1933 (N_1933,N_1886,N_1896);
and U1934 (N_1934,N_1862,N_1899);
or U1935 (N_1935,N_1839,N_1898);
nand U1936 (N_1936,N_1869,N_1858);
nor U1937 (N_1937,N_1825,N_1885);
and U1938 (N_1938,N_1824,N_1884);
or U1939 (N_1939,N_1889,N_1832);
and U1940 (N_1940,N_1850,N_1887);
nand U1941 (N_1941,N_1842,N_1834);
and U1942 (N_1942,N_1847,N_1878);
and U1943 (N_1943,N_1895,N_1888);
nand U1944 (N_1944,N_1800,N_1855);
nand U1945 (N_1945,N_1830,N_1803);
and U1946 (N_1946,N_1835,N_1845);
nand U1947 (N_1947,N_1876,N_1874);
and U1948 (N_1948,N_1866,N_1808);
xnor U1949 (N_1949,N_1828,N_1890);
nor U1950 (N_1950,N_1841,N_1854);
or U1951 (N_1951,N_1807,N_1891);
xor U1952 (N_1952,N_1888,N_1870);
nor U1953 (N_1953,N_1881,N_1803);
nand U1954 (N_1954,N_1829,N_1849);
nor U1955 (N_1955,N_1855,N_1867);
nand U1956 (N_1956,N_1836,N_1802);
and U1957 (N_1957,N_1881,N_1800);
nand U1958 (N_1958,N_1842,N_1887);
xnor U1959 (N_1959,N_1895,N_1870);
xor U1960 (N_1960,N_1836,N_1896);
xor U1961 (N_1961,N_1829,N_1820);
and U1962 (N_1962,N_1845,N_1890);
nand U1963 (N_1963,N_1832,N_1831);
nor U1964 (N_1964,N_1805,N_1807);
and U1965 (N_1965,N_1849,N_1886);
and U1966 (N_1966,N_1830,N_1859);
xor U1967 (N_1967,N_1888,N_1811);
xor U1968 (N_1968,N_1818,N_1844);
nor U1969 (N_1969,N_1853,N_1820);
nor U1970 (N_1970,N_1848,N_1805);
and U1971 (N_1971,N_1861,N_1876);
or U1972 (N_1972,N_1894,N_1893);
xor U1973 (N_1973,N_1848,N_1874);
xnor U1974 (N_1974,N_1859,N_1833);
nand U1975 (N_1975,N_1873,N_1874);
and U1976 (N_1976,N_1888,N_1813);
or U1977 (N_1977,N_1854,N_1844);
nor U1978 (N_1978,N_1808,N_1834);
and U1979 (N_1979,N_1879,N_1875);
and U1980 (N_1980,N_1824,N_1857);
xnor U1981 (N_1981,N_1802,N_1884);
nor U1982 (N_1982,N_1805,N_1852);
and U1983 (N_1983,N_1806,N_1883);
or U1984 (N_1984,N_1891,N_1833);
nor U1985 (N_1985,N_1865,N_1810);
or U1986 (N_1986,N_1889,N_1883);
or U1987 (N_1987,N_1868,N_1861);
nor U1988 (N_1988,N_1899,N_1878);
and U1989 (N_1989,N_1878,N_1883);
nand U1990 (N_1990,N_1846,N_1870);
or U1991 (N_1991,N_1800,N_1806);
or U1992 (N_1992,N_1896,N_1847);
nand U1993 (N_1993,N_1822,N_1866);
xor U1994 (N_1994,N_1875,N_1805);
or U1995 (N_1995,N_1808,N_1842);
nor U1996 (N_1996,N_1863,N_1884);
nand U1997 (N_1997,N_1844,N_1857);
nor U1998 (N_1998,N_1819,N_1815);
and U1999 (N_1999,N_1827,N_1885);
or U2000 (N_2000,N_1958,N_1935);
xnor U2001 (N_2001,N_1955,N_1906);
xnor U2002 (N_2002,N_1933,N_1917);
and U2003 (N_2003,N_1912,N_1913);
xor U2004 (N_2004,N_1972,N_1963);
or U2005 (N_2005,N_1992,N_1932);
nand U2006 (N_2006,N_1937,N_1981);
or U2007 (N_2007,N_1915,N_1965);
and U2008 (N_2008,N_1985,N_1929);
or U2009 (N_2009,N_1959,N_1986);
xnor U2010 (N_2010,N_1901,N_1982);
and U2011 (N_2011,N_1920,N_1909);
and U2012 (N_2012,N_1941,N_1988);
and U2013 (N_2013,N_1956,N_1940);
nor U2014 (N_2014,N_1926,N_1989);
or U2015 (N_2015,N_1990,N_1987);
nand U2016 (N_2016,N_1942,N_1925);
or U2017 (N_2017,N_1922,N_1934);
nand U2018 (N_2018,N_1924,N_1961);
xor U2019 (N_2019,N_1954,N_1908);
nand U2020 (N_2020,N_1951,N_1991);
nand U2021 (N_2021,N_1976,N_1931);
nand U2022 (N_2022,N_1952,N_1948);
nor U2023 (N_2023,N_1977,N_1984);
nor U2024 (N_2024,N_1918,N_1968);
xnor U2025 (N_2025,N_1923,N_1994);
xor U2026 (N_2026,N_1997,N_1953);
nand U2027 (N_2027,N_1964,N_1936);
nand U2028 (N_2028,N_1914,N_1962);
or U2029 (N_2029,N_1993,N_1974);
xor U2030 (N_2030,N_1911,N_1995);
nor U2031 (N_2031,N_1980,N_1966);
nor U2032 (N_2032,N_1904,N_1947);
nor U2033 (N_2033,N_1967,N_1996);
or U2034 (N_2034,N_1949,N_1916);
and U2035 (N_2035,N_1939,N_1910);
and U2036 (N_2036,N_1999,N_1900);
nor U2037 (N_2037,N_1902,N_1957);
nand U2038 (N_2038,N_1905,N_1944);
xor U2039 (N_2039,N_1978,N_1921);
and U2040 (N_2040,N_1973,N_1950);
nand U2041 (N_2041,N_1945,N_1907);
xor U2042 (N_2042,N_1938,N_1930);
xor U2043 (N_2043,N_1998,N_1970);
nand U2044 (N_2044,N_1919,N_1927);
nor U2045 (N_2045,N_1979,N_1943);
nand U2046 (N_2046,N_1946,N_1971);
nand U2047 (N_2047,N_1975,N_1903);
nor U2048 (N_2048,N_1960,N_1969);
xnor U2049 (N_2049,N_1928,N_1983);
and U2050 (N_2050,N_1903,N_1995);
nor U2051 (N_2051,N_1930,N_1903);
or U2052 (N_2052,N_1903,N_1920);
and U2053 (N_2053,N_1919,N_1942);
and U2054 (N_2054,N_1933,N_1930);
nand U2055 (N_2055,N_1901,N_1973);
xor U2056 (N_2056,N_1956,N_1955);
or U2057 (N_2057,N_1986,N_1932);
or U2058 (N_2058,N_1902,N_1909);
and U2059 (N_2059,N_1992,N_1907);
and U2060 (N_2060,N_1913,N_1958);
xnor U2061 (N_2061,N_1960,N_1983);
nor U2062 (N_2062,N_1963,N_1956);
nor U2063 (N_2063,N_1960,N_1924);
or U2064 (N_2064,N_1919,N_1967);
xnor U2065 (N_2065,N_1924,N_1995);
nor U2066 (N_2066,N_1951,N_1961);
nand U2067 (N_2067,N_1947,N_1907);
or U2068 (N_2068,N_1904,N_1934);
xor U2069 (N_2069,N_1950,N_1974);
xor U2070 (N_2070,N_1948,N_1977);
nand U2071 (N_2071,N_1994,N_1949);
nand U2072 (N_2072,N_1981,N_1904);
and U2073 (N_2073,N_1934,N_1900);
or U2074 (N_2074,N_1901,N_1996);
nand U2075 (N_2075,N_1941,N_1921);
nor U2076 (N_2076,N_1966,N_1906);
nand U2077 (N_2077,N_1999,N_1959);
nor U2078 (N_2078,N_1999,N_1906);
xor U2079 (N_2079,N_1990,N_1959);
or U2080 (N_2080,N_1917,N_1984);
and U2081 (N_2081,N_1900,N_1943);
or U2082 (N_2082,N_1988,N_1993);
xnor U2083 (N_2083,N_1977,N_1962);
nor U2084 (N_2084,N_1948,N_1938);
and U2085 (N_2085,N_1970,N_1995);
xnor U2086 (N_2086,N_1937,N_1931);
and U2087 (N_2087,N_1933,N_1964);
xor U2088 (N_2088,N_1939,N_1905);
and U2089 (N_2089,N_1962,N_1937);
nor U2090 (N_2090,N_1933,N_1918);
or U2091 (N_2091,N_1967,N_1907);
nor U2092 (N_2092,N_1984,N_1924);
nand U2093 (N_2093,N_1974,N_1921);
or U2094 (N_2094,N_1933,N_1971);
or U2095 (N_2095,N_1966,N_1969);
and U2096 (N_2096,N_1931,N_1947);
and U2097 (N_2097,N_1992,N_1906);
or U2098 (N_2098,N_1930,N_1972);
nor U2099 (N_2099,N_1945,N_1970);
nand U2100 (N_2100,N_2045,N_2075);
and U2101 (N_2101,N_2013,N_2064);
or U2102 (N_2102,N_2037,N_2073);
xor U2103 (N_2103,N_2007,N_2067);
or U2104 (N_2104,N_2049,N_2061);
or U2105 (N_2105,N_2068,N_2089);
xnor U2106 (N_2106,N_2058,N_2093);
and U2107 (N_2107,N_2081,N_2095);
and U2108 (N_2108,N_2001,N_2020);
nand U2109 (N_2109,N_2078,N_2040);
xor U2110 (N_2110,N_2033,N_2015);
nor U2111 (N_2111,N_2031,N_2042);
or U2112 (N_2112,N_2071,N_2080);
xnor U2113 (N_2113,N_2006,N_2070);
and U2114 (N_2114,N_2084,N_2027);
xnor U2115 (N_2115,N_2021,N_2003);
xor U2116 (N_2116,N_2050,N_2085);
or U2117 (N_2117,N_2030,N_2072);
nor U2118 (N_2118,N_2029,N_2094);
and U2119 (N_2119,N_2014,N_2032);
nand U2120 (N_2120,N_2017,N_2018);
xor U2121 (N_2121,N_2057,N_2048);
nor U2122 (N_2122,N_2056,N_2090);
and U2123 (N_2123,N_2009,N_2099);
nor U2124 (N_2124,N_2028,N_2054);
or U2125 (N_2125,N_2098,N_2034);
and U2126 (N_2126,N_2087,N_2059);
xor U2127 (N_2127,N_2062,N_2038);
xor U2128 (N_2128,N_2026,N_2019);
xor U2129 (N_2129,N_2063,N_2023);
or U2130 (N_2130,N_2004,N_2083);
or U2131 (N_2131,N_2036,N_2043);
nand U2132 (N_2132,N_2055,N_2076);
or U2133 (N_2133,N_2079,N_2091);
nor U2134 (N_2134,N_2082,N_2052);
or U2135 (N_2135,N_2065,N_2088);
nor U2136 (N_2136,N_2066,N_2086);
nor U2137 (N_2137,N_2025,N_2016);
nand U2138 (N_2138,N_2008,N_2022);
nor U2139 (N_2139,N_2053,N_2005);
nand U2140 (N_2140,N_2060,N_2092);
xnor U2141 (N_2141,N_2035,N_2044);
nor U2142 (N_2142,N_2002,N_2024);
nand U2143 (N_2143,N_2000,N_2097);
xor U2144 (N_2144,N_2047,N_2077);
and U2145 (N_2145,N_2069,N_2074);
or U2146 (N_2146,N_2039,N_2046);
or U2147 (N_2147,N_2051,N_2096);
nor U2148 (N_2148,N_2011,N_2041);
xnor U2149 (N_2149,N_2010,N_2012);
xor U2150 (N_2150,N_2010,N_2053);
xor U2151 (N_2151,N_2083,N_2090);
nand U2152 (N_2152,N_2040,N_2024);
or U2153 (N_2153,N_2058,N_2014);
xnor U2154 (N_2154,N_2073,N_2005);
nor U2155 (N_2155,N_2016,N_2058);
xnor U2156 (N_2156,N_2017,N_2060);
and U2157 (N_2157,N_2001,N_2071);
nand U2158 (N_2158,N_2037,N_2044);
and U2159 (N_2159,N_2064,N_2073);
nor U2160 (N_2160,N_2039,N_2052);
and U2161 (N_2161,N_2021,N_2067);
nand U2162 (N_2162,N_2061,N_2047);
xor U2163 (N_2163,N_2029,N_2097);
nor U2164 (N_2164,N_2087,N_2045);
or U2165 (N_2165,N_2001,N_2050);
or U2166 (N_2166,N_2039,N_2009);
xor U2167 (N_2167,N_2085,N_2086);
nor U2168 (N_2168,N_2017,N_2055);
xnor U2169 (N_2169,N_2033,N_2025);
and U2170 (N_2170,N_2059,N_2072);
xnor U2171 (N_2171,N_2097,N_2008);
and U2172 (N_2172,N_2007,N_2048);
nand U2173 (N_2173,N_2076,N_2017);
nor U2174 (N_2174,N_2087,N_2077);
nor U2175 (N_2175,N_2046,N_2050);
nor U2176 (N_2176,N_2093,N_2000);
xor U2177 (N_2177,N_2054,N_2007);
and U2178 (N_2178,N_2069,N_2053);
or U2179 (N_2179,N_2030,N_2044);
xor U2180 (N_2180,N_2045,N_2082);
nand U2181 (N_2181,N_2083,N_2011);
nor U2182 (N_2182,N_2095,N_2000);
xor U2183 (N_2183,N_2039,N_2038);
nor U2184 (N_2184,N_2072,N_2078);
or U2185 (N_2185,N_2099,N_2021);
nand U2186 (N_2186,N_2054,N_2037);
xor U2187 (N_2187,N_2016,N_2023);
nor U2188 (N_2188,N_2058,N_2035);
nor U2189 (N_2189,N_2065,N_2024);
nor U2190 (N_2190,N_2079,N_2010);
nand U2191 (N_2191,N_2021,N_2053);
and U2192 (N_2192,N_2060,N_2009);
nand U2193 (N_2193,N_2027,N_2070);
nor U2194 (N_2194,N_2023,N_2052);
nand U2195 (N_2195,N_2086,N_2018);
nand U2196 (N_2196,N_2093,N_2069);
nor U2197 (N_2197,N_2028,N_2016);
nand U2198 (N_2198,N_2040,N_2044);
or U2199 (N_2199,N_2056,N_2099);
nor U2200 (N_2200,N_2146,N_2114);
xnor U2201 (N_2201,N_2148,N_2183);
xor U2202 (N_2202,N_2136,N_2160);
nor U2203 (N_2203,N_2102,N_2119);
or U2204 (N_2204,N_2120,N_2111);
nor U2205 (N_2205,N_2110,N_2199);
or U2206 (N_2206,N_2181,N_2132);
xnor U2207 (N_2207,N_2154,N_2109);
and U2208 (N_2208,N_2152,N_2122);
nand U2209 (N_2209,N_2150,N_2108);
nand U2210 (N_2210,N_2194,N_2179);
nand U2211 (N_2211,N_2123,N_2128);
or U2212 (N_2212,N_2176,N_2187);
xnor U2213 (N_2213,N_2127,N_2185);
and U2214 (N_2214,N_2157,N_2158);
nor U2215 (N_2215,N_2144,N_2163);
nand U2216 (N_2216,N_2198,N_2118);
nand U2217 (N_2217,N_2197,N_2103);
xnor U2218 (N_2218,N_2180,N_2143);
xor U2219 (N_2219,N_2107,N_2161);
or U2220 (N_2220,N_2147,N_2193);
nand U2221 (N_2221,N_2162,N_2168);
xnor U2222 (N_2222,N_2124,N_2177);
or U2223 (N_2223,N_2137,N_2184);
or U2224 (N_2224,N_2159,N_2182);
xor U2225 (N_2225,N_2116,N_2133);
xnor U2226 (N_2226,N_2167,N_2173);
or U2227 (N_2227,N_2174,N_2131);
or U2228 (N_2228,N_2126,N_2153);
nand U2229 (N_2229,N_2141,N_2105);
nor U2230 (N_2230,N_2169,N_2186);
nor U2231 (N_2231,N_2113,N_2189);
or U2232 (N_2232,N_2166,N_2188);
nand U2233 (N_2233,N_2145,N_2170);
and U2234 (N_2234,N_2156,N_2106);
and U2235 (N_2235,N_2142,N_2195);
nand U2236 (N_2236,N_2138,N_2100);
nor U2237 (N_2237,N_2121,N_2178);
xor U2238 (N_2238,N_2165,N_2151);
nor U2239 (N_2239,N_2125,N_2172);
xnor U2240 (N_2240,N_2101,N_2135);
nand U2241 (N_2241,N_2190,N_2191);
nand U2242 (N_2242,N_2164,N_2155);
and U2243 (N_2243,N_2112,N_2134);
and U2244 (N_2244,N_2175,N_2192);
or U2245 (N_2245,N_2129,N_2196);
or U2246 (N_2246,N_2140,N_2117);
and U2247 (N_2247,N_2171,N_2130);
nand U2248 (N_2248,N_2104,N_2115);
xor U2249 (N_2249,N_2139,N_2149);
and U2250 (N_2250,N_2107,N_2180);
xor U2251 (N_2251,N_2156,N_2189);
xnor U2252 (N_2252,N_2143,N_2106);
or U2253 (N_2253,N_2110,N_2151);
xor U2254 (N_2254,N_2190,N_2150);
and U2255 (N_2255,N_2146,N_2141);
nor U2256 (N_2256,N_2152,N_2151);
and U2257 (N_2257,N_2150,N_2136);
nor U2258 (N_2258,N_2153,N_2194);
or U2259 (N_2259,N_2184,N_2197);
or U2260 (N_2260,N_2141,N_2190);
xnor U2261 (N_2261,N_2186,N_2122);
and U2262 (N_2262,N_2165,N_2130);
and U2263 (N_2263,N_2167,N_2147);
and U2264 (N_2264,N_2171,N_2112);
nor U2265 (N_2265,N_2192,N_2134);
or U2266 (N_2266,N_2100,N_2144);
nand U2267 (N_2267,N_2113,N_2127);
or U2268 (N_2268,N_2144,N_2103);
xor U2269 (N_2269,N_2158,N_2189);
and U2270 (N_2270,N_2189,N_2172);
nand U2271 (N_2271,N_2181,N_2155);
and U2272 (N_2272,N_2173,N_2130);
nand U2273 (N_2273,N_2150,N_2157);
nor U2274 (N_2274,N_2126,N_2169);
nand U2275 (N_2275,N_2106,N_2190);
nand U2276 (N_2276,N_2198,N_2144);
xnor U2277 (N_2277,N_2106,N_2113);
or U2278 (N_2278,N_2119,N_2133);
nor U2279 (N_2279,N_2155,N_2157);
or U2280 (N_2280,N_2196,N_2134);
nand U2281 (N_2281,N_2124,N_2195);
xnor U2282 (N_2282,N_2115,N_2137);
and U2283 (N_2283,N_2168,N_2179);
and U2284 (N_2284,N_2103,N_2157);
nand U2285 (N_2285,N_2182,N_2160);
or U2286 (N_2286,N_2125,N_2160);
and U2287 (N_2287,N_2105,N_2166);
nor U2288 (N_2288,N_2163,N_2107);
nand U2289 (N_2289,N_2152,N_2108);
xor U2290 (N_2290,N_2109,N_2105);
and U2291 (N_2291,N_2161,N_2177);
and U2292 (N_2292,N_2122,N_2135);
nor U2293 (N_2293,N_2154,N_2178);
and U2294 (N_2294,N_2185,N_2137);
or U2295 (N_2295,N_2154,N_2181);
nor U2296 (N_2296,N_2166,N_2136);
xnor U2297 (N_2297,N_2168,N_2155);
nand U2298 (N_2298,N_2105,N_2138);
nand U2299 (N_2299,N_2171,N_2151);
or U2300 (N_2300,N_2280,N_2224);
nand U2301 (N_2301,N_2238,N_2248);
nand U2302 (N_2302,N_2254,N_2214);
or U2303 (N_2303,N_2282,N_2265);
xor U2304 (N_2304,N_2237,N_2220);
or U2305 (N_2305,N_2236,N_2294);
or U2306 (N_2306,N_2273,N_2219);
nor U2307 (N_2307,N_2247,N_2267);
xor U2308 (N_2308,N_2204,N_2284);
and U2309 (N_2309,N_2277,N_2289);
and U2310 (N_2310,N_2274,N_2250);
nand U2311 (N_2311,N_2230,N_2240);
and U2312 (N_2312,N_2263,N_2291);
nor U2313 (N_2313,N_2246,N_2212);
and U2314 (N_2314,N_2245,N_2286);
nor U2315 (N_2315,N_2234,N_2207);
nor U2316 (N_2316,N_2253,N_2241);
or U2317 (N_2317,N_2221,N_2292);
xnor U2318 (N_2318,N_2270,N_2257);
xnor U2319 (N_2319,N_2295,N_2217);
or U2320 (N_2320,N_2258,N_2215);
nor U2321 (N_2321,N_2256,N_2251);
nand U2322 (N_2322,N_2229,N_2210);
nor U2323 (N_2323,N_2208,N_2239);
and U2324 (N_2324,N_2264,N_2203);
nor U2325 (N_2325,N_2225,N_2211);
and U2326 (N_2326,N_2278,N_2202);
and U2327 (N_2327,N_2233,N_2269);
or U2328 (N_2328,N_2223,N_2228);
and U2329 (N_2329,N_2260,N_2288);
and U2330 (N_2330,N_2209,N_2252);
xnor U2331 (N_2331,N_2205,N_2262);
and U2332 (N_2332,N_2206,N_2299);
and U2333 (N_2333,N_2243,N_2242);
or U2334 (N_2334,N_2296,N_2244);
xor U2335 (N_2335,N_2290,N_2297);
and U2336 (N_2336,N_2283,N_2268);
nor U2337 (N_2337,N_2271,N_2285);
nand U2338 (N_2338,N_2226,N_2218);
nor U2339 (N_2339,N_2279,N_2213);
and U2340 (N_2340,N_2222,N_2287);
nand U2341 (N_2341,N_2255,N_2293);
nand U2342 (N_2342,N_2232,N_2227);
or U2343 (N_2343,N_2231,N_2266);
or U2344 (N_2344,N_2281,N_2275);
xnor U2345 (N_2345,N_2249,N_2259);
or U2346 (N_2346,N_2272,N_2298);
nand U2347 (N_2347,N_2216,N_2200);
nand U2348 (N_2348,N_2261,N_2235);
nor U2349 (N_2349,N_2276,N_2201);
xor U2350 (N_2350,N_2276,N_2266);
nor U2351 (N_2351,N_2241,N_2272);
or U2352 (N_2352,N_2238,N_2268);
nand U2353 (N_2353,N_2219,N_2253);
xnor U2354 (N_2354,N_2247,N_2256);
nor U2355 (N_2355,N_2204,N_2298);
nand U2356 (N_2356,N_2255,N_2263);
nand U2357 (N_2357,N_2264,N_2241);
or U2358 (N_2358,N_2212,N_2269);
nand U2359 (N_2359,N_2294,N_2220);
nand U2360 (N_2360,N_2280,N_2211);
nor U2361 (N_2361,N_2262,N_2257);
nand U2362 (N_2362,N_2278,N_2237);
xor U2363 (N_2363,N_2260,N_2267);
xnor U2364 (N_2364,N_2287,N_2218);
or U2365 (N_2365,N_2215,N_2217);
and U2366 (N_2366,N_2207,N_2265);
or U2367 (N_2367,N_2201,N_2256);
nor U2368 (N_2368,N_2273,N_2294);
nand U2369 (N_2369,N_2214,N_2259);
nand U2370 (N_2370,N_2288,N_2217);
nand U2371 (N_2371,N_2222,N_2290);
nand U2372 (N_2372,N_2248,N_2269);
nor U2373 (N_2373,N_2295,N_2207);
nor U2374 (N_2374,N_2213,N_2294);
nor U2375 (N_2375,N_2296,N_2205);
nor U2376 (N_2376,N_2257,N_2286);
or U2377 (N_2377,N_2256,N_2235);
and U2378 (N_2378,N_2295,N_2208);
xor U2379 (N_2379,N_2256,N_2252);
or U2380 (N_2380,N_2280,N_2239);
nand U2381 (N_2381,N_2212,N_2287);
and U2382 (N_2382,N_2232,N_2202);
nor U2383 (N_2383,N_2266,N_2240);
and U2384 (N_2384,N_2207,N_2214);
nand U2385 (N_2385,N_2200,N_2204);
nor U2386 (N_2386,N_2205,N_2283);
nor U2387 (N_2387,N_2216,N_2298);
nand U2388 (N_2388,N_2273,N_2292);
nor U2389 (N_2389,N_2229,N_2268);
nor U2390 (N_2390,N_2269,N_2299);
nor U2391 (N_2391,N_2222,N_2201);
or U2392 (N_2392,N_2213,N_2295);
or U2393 (N_2393,N_2263,N_2268);
nor U2394 (N_2394,N_2211,N_2266);
nor U2395 (N_2395,N_2231,N_2203);
or U2396 (N_2396,N_2226,N_2262);
nor U2397 (N_2397,N_2253,N_2290);
xnor U2398 (N_2398,N_2202,N_2240);
nand U2399 (N_2399,N_2299,N_2268);
or U2400 (N_2400,N_2332,N_2362);
nand U2401 (N_2401,N_2380,N_2316);
nand U2402 (N_2402,N_2357,N_2300);
and U2403 (N_2403,N_2349,N_2322);
and U2404 (N_2404,N_2345,N_2306);
and U2405 (N_2405,N_2374,N_2305);
xnor U2406 (N_2406,N_2388,N_2303);
nand U2407 (N_2407,N_2314,N_2343);
and U2408 (N_2408,N_2378,N_2354);
xor U2409 (N_2409,N_2346,N_2321);
and U2410 (N_2410,N_2341,N_2326);
nand U2411 (N_2411,N_2336,N_2318);
xnor U2412 (N_2412,N_2340,N_2348);
and U2413 (N_2413,N_2361,N_2344);
nor U2414 (N_2414,N_2391,N_2363);
or U2415 (N_2415,N_2395,N_2373);
xnor U2416 (N_2416,N_2350,N_2379);
or U2417 (N_2417,N_2317,N_2372);
nor U2418 (N_2418,N_2311,N_2360);
nand U2419 (N_2419,N_2337,N_2319);
xnor U2420 (N_2420,N_2397,N_2366);
or U2421 (N_2421,N_2392,N_2365);
and U2422 (N_2422,N_2308,N_2399);
and U2423 (N_2423,N_2393,N_2371);
and U2424 (N_2424,N_2382,N_2310);
and U2425 (N_2425,N_2359,N_2304);
nand U2426 (N_2426,N_2339,N_2367);
nand U2427 (N_2427,N_2369,N_2313);
and U2428 (N_2428,N_2355,N_2375);
or U2429 (N_2429,N_2301,N_2368);
nand U2430 (N_2430,N_2383,N_2328);
and U2431 (N_2431,N_2335,N_2386);
or U2432 (N_2432,N_2323,N_2370);
and U2433 (N_2433,N_2320,N_2396);
xnor U2434 (N_2434,N_2342,N_2356);
and U2435 (N_2435,N_2390,N_2327);
nand U2436 (N_2436,N_2376,N_2331);
or U2437 (N_2437,N_2387,N_2351);
and U2438 (N_2438,N_2307,N_2352);
nand U2439 (N_2439,N_2324,N_2325);
nor U2440 (N_2440,N_2312,N_2377);
xnor U2441 (N_2441,N_2347,N_2334);
xor U2442 (N_2442,N_2330,N_2364);
nand U2443 (N_2443,N_2338,N_2329);
xor U2444 (N_2444,N_2385,N_2353);
nor U2445 (N_2445,N_2302,N_2384);
or U2446 (N_2446,N_2394,N_2315);
xnor U2447 (N_2447,N_2389,N_2398);
nand U2448 (N_2448,N_2309,N_2333);
and U2449 (N_2449,N_2358,N_2381);
and U2450 (N_2450,N_2350,N_2338);
or U2451 (N_2451,N_2316,N_2393);
nor U2452 (N_2452,N_2315,N_2392);
nor U2453 (N_2453,N_2368,N_2337);
xor U2454 (N_2454,N_2306,N_2355);
nand U2455 (N_2455,N_2383,N_2323);
xnor U2456 (N_2456,N_2334,N_2314);
or U2457 (N_2457,N_2371,N_2326);
and U2458 (N_2458,N_2328,N_2325);
and U2459 (N_2459,N_2317,N_2345);
or U2460 (N_2460,N_2324,N_2389);
or U2461 (N_2461,N_2310,N_2383);
xor U2462 (N_2462,N_2303,N_2306);
and U2463 (N_2463,N_2351,N_2388);
nor U2464 (N_2464,N_2300,N_2382);
nor U2465 (N_2465,N_2332,N_2311);
xor U2466 (N_2466,N_2360,N_2387);
xnor U2467 (N_2467,N_2350,N_2342);
or U2468 (N_2468,N_2338,N_2303);
or U2469 (N_2469,N_2363,N_2347);
or U2470 (N_2470,N_2345,N_2396);
nor U2471 (N_2471,N_2388,N_2394);
nor U2472 (N_2472,N_2300,N_2378);
nor U2473 (N_2473,N_2389,N_2305);
or U2474 (N_2474,N_2372,N_2392);
nand U2475 (N_2475,N_2342,N_2396);
nor U2476 (N_2476,N_2399,N_2334);
nand U2477 (N_2477,N_2373,N_2322);
nor U2478 (N_2478,N_2353,N_2352);
or U2479 (N_2479,N_2303,N_2370);
nor U2480 (N_2480,N_2345,N_2302);
nand U2481 (N_2481,N_2340,N_2347);
xor U2482 (N_2482,N_2386,N_2333);
and U2483 (N_2483,N_2335,N_2382);
xnor U2484 (N_2484,N_2371,N_2346);
xor U2485 (N_2485,N_2366,N_2359);
nor U2486 (N_2486,N_2326,N_2348);
xnor U2487 (N_2487,N_2302,N_2337);
nand U2488 (N_2488,N_2350,N_2388);
nor U2489 (N_2489,N_2376,N_2389);
nor U2490 (N_2490,N_2386,N_2301);
xor U2491 (N_2491,N_2313,N_2356);
and U2492 (N_2492,N_2387,N_2383);
and U2493 (N_2493,N_2381,N_2304);
and U2494 (N_2494,N_2322,N_2383);
nand U2495 (N_2495,N_2305,N_2341);
nand U2496 (N_2496,N_2339,N_2309);
and U2497 (N_2497,N_2387,N_2373);
xnor U2498 (N_2498,N_2328,N_2399);
nand U2499 (N_2499,N_2319,N_2380);
or U2500 (N_2500,N_2414,N_2481);
xor U2501 (N_2501,N_2401,N_2432);
xnor U2502 (N_2502,N_2400,N_2462);
and U2503 (N_2503,N_2422,N_2425);
nand U2504 (N_2504,N_2452,N_2460);
or U2505 (N_2505,N_2486,N_2467);
nor U2506 (N_2506,N_2413,N_2411);
or U2507 (N_2507,N_2433,N_2497);
or U2508 (N_2508,N_2419,N_2488);
nor U2509 (N_2509,N_2439,N_2441);
and U2510 (N_2510,N_2475,N_2404);
and U2511 (N_2511,N_2494,N_2447);
nand U2512 (N_2512,N_2436,N_2476);
and U2513 (N_2513,N_2457,N_2429);
or U2514 (N_2514,N_2456,N_2435);
and U2515 (N_2515,N_2465,N_2468);
nor U2516 (N_2516,N_2498,N_2412);
or U2517 (N_2517,N_2461,N_2445);
and U2518 (N_2518,N_2440,N_2430);
or U2519 (N_2519,N_2417,N_2485);
xnor U2520 (N_2520,N_2471,N_2454);
nor U2521 (N_2521,N_2470,N_2491);
nor U2522 (N_2522,N_2428,N_2442);
nand U2523 (N_2523,N_2406,N_2431);
or U2524 (N_2524,N_2496,N_2463);
nand U2525 (N_2525,N_2480,N_2420);
xor U2526 (N_2526,N_2408,N_2455);
xnor U2527 (N_2527,N_2444,N_2472);
and U2528 (N_2528,N_2489,N_2492);
nand U2529 (N_2529,N_2479,N_2451);
nor U2530 (N_2530,N_2466,N_2459);
and U2531 (N_2531,N_2448,N_2409);
and U2532 (N_2532,N_2482,N_2410);
nand U2533 (N_2533,N_2478,N_2446);
xor U2534 (N_2534,N_2499,N_2449);
nor U2535 (N_2535,N_2473,N_2483);
or U2536 (N_2536,N_2423,N_2416);
and U2537 (N_2537,N_2427,N_2484);
nor U2538 (N_2538,N_2458,N_2495);
and U2539 (N_2539,N_2418,N_2405);
or U2540 (N_2540,N_2450,N_2487);
or U2541 (N_2541,N_2426,N_2415);
xor U2542 (N_2542,N_2490,N_2403);
xnor U2543 (N_2543,N_2421,N_2443);
xor U2544 (N_2544,N_2477,N_2469);
or U2545 (N_2545,N_2474,N_2493);
nand U2546 (N_2546,N_2464,N_2438);
xnor U2547 (N_2547,N_2402,N_2453);
nor U2548 (N_2548,N_2424,N_2437);
or U2549 (N_2549,N_2407,N_2434);
nand U2550 (N_2550,N_2491,N_2409);
xnor U2551 (N_2551,N_2467,N_2477);
and U2552 (N_2552,N_2425,N_2491);
nand U2553 (N_2553,N_2497,N_2491);
xor U2554 (N_2554,N_2404,N_2416);
nand U2555 (N_2555,N_2498,N_2474);
and U2556 (N_2556,N_2450,N_2414);
nor U2557 (N_2557,N_2440,N_2497);
nand U2558 (N_2558,N_2448,N_2467);
xnor U2559 (N_2559,N_2451,N_2421);
nor U2560 (N_2560,N_2438,N_2437);
xnor U2561 (N_2561,N_2426,N_2459);
nand U2562 (N_2562,N_2466,N_2464);
and U2563 (N_2563,N_2400,N_2403);
nor U2564 (N_2564,N_2473,N_2451);
xor U2565 (N_2565,N_2409,N_2404);
or U2566 (N_2566,N_2426,N_2485);
and U2567 (N_2567,N_2480,N_2443);
nand U2568 (N_2568,N_2461,N_2404);
or U2569 (N_2569,N_2424,N_2479);
xnor U2570 (N_2570,N_2451,N_2438);
and U2571 (N_2571,N_2473,N_2452);
nand U2572 (N_2572,N_2429,N_2430);
or U2573 (N_2573,N_2431,N_2457);
nand U2574 (N_2574,N_2407,N_2403);
nor U2575 (N_2575,N_2404,N_2496);
nand U2576 (N_2576,N_2400,N_2460);
nor U2577 (N_2577,N_2487,N_2429);
nor U2578 (N_2578,N_2437,N_2420);
nand U2579 (N_2579,N_2414,N_2482);
and U2580 (N_2580,N_2478,N_2449);
nor U2581 (N_2581,N_2406,N_2463);
and U2582 (N_2582,N_2460,N_2431);
and U2583 (N_2583,N_2404,N_2497);
and U2584 (N_2584,N_2442,N_2468);
and U2585 (N_2585,N_2443,N_2466);
xnor U2586 (N_2586,N_2480,N_2436);
xnor U2587 (N_2587,N_2412,N_2453);
nor U2588 (N_2588,N_2434,N_2427);
or U2589 (N_2589,N_2437,N_2497);
xnor U2590 (N_2590,N_2490,N_2460);
nor U2591 (N_2591,N_2407,N_2417);
or U2592 (N_2592,N_2492,N_2479);
nand U2593 (N_2593,N_2401,N_2454);
nor U2594 (N_2594,N_2407,N_2484);
xor U2595 (N_2595,N_2439,N_2493);
xnor U2596 (N_2596,N_2440,N_2482);
or U2597 (N_2597,N_2471,N_2487);
nand U2598 (N_2598,N_2419,N_2436);
or U2599 (N_2599,N_2465,N_2490);
or U2600 (N_2600,N_2509,N_2514);
and U2601 (N_2601,N_2508,N_2519);
nor U2602 (N_2602,N_2595,N_2586);
and U2603 (N_2603,N_2572,N_2510);
nand U2604 (N_2604,N_2597,N_2526);
xnor U2605 (N_2605,N_2583,N_2505);
or U2606 (N_2606,N_2532,N_2520);
nor U2607 (N_2607,N_2546,N_2535);
nand U2608 (N_2608,N_2548,N_2525);
and U2609 (N_2609,N_2554,N_2584);
or U2610 (N_2610,N_2538,N_2581);
nand U2611 (N_2611,N_2580,N_2573);
nor U2612 (N_2612,N_2585,N_2558);
nor U2613 (N_2613,N_2515,N_2575);
nor U2614 (N_2614,N_2506,N_2523);
or U2615 (N_2615,N_2588,N_2528);
xor U2616 (N_2616,N_2522,N_2593);
nor U2617 (N_2617,N_2543,N_2534);
xor U2618 (N_2618,N_2552,N_2539);
nand U2619 (N_2619,N_2599,N_2545);
nand U2620 (N_2620,N_2570,N_2507);
or U2621 (N_2621,N_2587,N_2596);
nand U2622 (N_2622,N_2578,N_2521);
and U2623 (N_2623,N_2555,N_2549);
and U2624 (N_2624,N_2574,N_2536);
nor U2625 (N_2625,N_2542,N_2531);
nor U2626 (N_2626,N_2561,N_2568);
nor U2627 (N_2627,N_2513,N_2512);
nor U2628 (N_2628,N_2517,N_2563);
and U2629 (N_2629,N_2566,N_2500);
or U2630 (N_2630,N_2503,N_2551);
and U2631 (N_2631,N_2553,N_2592);
xor U2632 (N_2632,N_2565,N_2590);
nor U2633 (N_2633,N_2511,N_2559);
nor U2634 (N_2634,N_2537,N_2529);
xor U2635 (N_2635,N_2589,N_2560);
and U2636 (N_2636,N_2550,N_2557);
nor U2637 (N_2637,N_2567,N_2530);
or U2638 (N_2638,N_2576,N_2540);
or U2639 (N_2639,N_2591,N_2582);
nor U2640 (N_2640,N_2541,N_2562);
xor U2641 (N_2641,N_2564,N_2544);
or U2642 (N_2642,N_2518,N_2556);
nand U2643 (N_2643,N_2579,N_2527);
nor U2644 (N_2644,N_2502,N_2577);
nand U2645 (N_2645,N_2504,N_2524);
nor U2646 (N_2646,N_2594,N_2569);
and U2647 (N_2647,N_2501,N_2516);
or U2648 (N_2648,N_2533,N_2598);
and U2649 (N_2649,N_2547,N_2571);
or U2650 (N_2650,N_2533,N_2538);
nand U2651 (N_2651,N_2549,N_2570);
or U2652 (N_2652,N_2545,N_2588);
nand U2653 (N_2653,N_2518,N_2520);
nand U2654 (N_2654,N_2589,N_2577);
and U2655 (N_2655,N_2551,N_2525);
nand U2656 (N_2656,N_2556,N_2570);
and U2657 (N_2657,N_2543,N_2520);
and U2658 (N_2658,N_2504,N_2521);
or U2659 (N_2659,N_2598,N_2541);
and U2660 (N_2660,N_2590,N_2550);
and U2661 (N_2661,N_2541,N_2568);
nor U2662 (N_2662,N_2525,N_2540);
xnor U2663 (N_2663,N_2512,N_2569);
nand U2664 (N_2664,N_2538,N_2559);
or U2665 (N_2665,N_2590,N_2547);
or U2666 (N_2666,N_2529,N_2564);
and U2667 (N_2667,N_2566,N_2531);
xnor U2668 (N_2668,N_2527,N_2548);
or U2669 (N_2669,N_2593,N_2536);
xor U2670 (N_2670,N_2587,N_2544);
or U2671 (N_2671,N_2527,N_2561);
and U2672 (N_2672,N_2591,N_2506);
nor U2673 (N_2673,N_2558,N_2555);
nand U2674 (N_2674,N_2547,N_2554);
or U2675 (N_2675,N_2540,N_2554);
nand U2676 (N_2676,N_2580,N_2566);
or U2677 (N_2677,N_2593,N_2543);
nor U2678 (N_2678,N_2570,N_2581);
or U2679 (N_2679,N_2505,N_2551);
or U2680 (N_2680,N_2538,N_2517);
xnor U2681 (N_2681,N_2549,N_2578);
xnor U2682 (N_2682,N_2550,N_2583);
xnor U2683 (N_2683,N_2556,N_2598);
xnor U2684 (N_2684,N_2589,N_2535);
or U2685 (N_2685,N_2592,N_2535);
xnor U2686 (N_2686,N_2597,N_2544);
xnor U2687 (N_2687,N_2517,N_2509);
or U2688 (N_2688,N_2514,N_2528);
xor U2689 (N_2689,N_2511,N_2584);
nand U2690 (N_2690,N_2579,N_2512);
or U2691 (N_2691,N_2567,N_2525);
xor U2692 (N_2692,N_2519,N_2520);
or U2693 (N_2693,N_2596,N_2557);
nand U2694 (N_2694,N_2583,N_2508);
xor U2695 (N_2695,N_2562,N_2515);
xor U2696 (N_2696,N_2579,N_2591);
nor U2697 (N_2697,N_2589,N_2595);
nor U2698 (N_2698,N_2552,N_2523);
xnor U2699 (N_2699,N_2535,N_2574);
nor U2700 (N_2700,N_2695,N_2686);
and U2701 (N_2701,N_2629,N_2641);
nand U2702 (N_2702,N_2650,N_2682);
nor U2703 (N_2703,N_2662,N_2609);
and U2704 (N_2704,N_2617,N_2669);
or U2705 (N_2705,N_2676,N_2653);
or U2706 (N_2706,N_2615,N_2656);
xnor U2707 (N_2707,N_2652,N_2612);
xor U2708 (N_2708,N_2628,N_2605);
and U2709 (N_2709,N_2680,N_2657);
or U2710 (N_2710,N_2688,N_2647);
xor U2711 (N_2711,N_2636,N_2670);
or U2712 (N_2712,N_2614,N_2633);
and U2713 (N_2713,N_2603,N_2608);
xor U2714 (N_2714,N_2602,N_2619);
xnor U2715 (N_2715,N_2623,N_2634);
nand U2716 (N_2716,N_2681,N_2699);
nor U2717 (N_2717,N_2661,N_2626);
xnor U2718 (N_2718,N_2646,N_2601);
and U2719 (N_2719,N_2672,N_2625);
and U2720 (N_2720,N_2687,N_2689);
nor U2721 (N_2721,N_2697,N_2654);
nor U2722 (N_2722,N_2698,N_2671);
nor U2723 (N_2723,N_2620,N_2643);
nand U2724 (N_2724,N_2673,N_2692);
or U2725 (N_2725,N_2691,N_2637);
nor U2726 (N_2726,N_2616,N_2666);
or U2727 (N_2727,N_2678,N_2649);
nand U2728 (N_2728,N_2684,N_2611);
nand U2729 (N_2729,N_2663,N_2607);
xor U2730 (N_2730,N_2606,N_2694);
xor U2731 (N_2731,N_2675,N_2664);
or U2732 (N_2732,N_2604,N_2642);
nor U2733 (N_2733,N_2645,N_2613);
nor U2734 (N_2734,N_2674,N_2696);
nor U2735 (N_2735,N_2667,N_2632);
xnor U2736 (N_2736,N_2639,N_2618);
nand U2737 (N_2737,N_2693,N_2651);
or U2738 (N_2738,N_2631,N_2679);
nand U2739 (N_2739,N_2638,N_2610);
nor U2740 (N_2740,N_2630,N_2624);
nand U2741 (N_2741,N_2655,N_2690);
or U2742 (N_2742,N_2627,N_2668);
nor U2743 (N_2743,N_2648,N_2659);
or U2744 (N_2744,N_2660,N_2644);
and U2745 (N_2745,N_2640,N_2677);
nor U2746 (N_2746,N_2658,N_2665);
and U2747 (N_2747,N_2685,N_2621);
nand U2748 (N_2748,N_2600,N_2635);
xor U2749 (N_2749,N_2683,N_2622);
nand U2750 (N_2750,N_2613,N_2656);
xnor U2751 (N_2751,N_2668,N_2614);
nand U2752 (N_2752,N_2633,N_2652);
and U2753 (N_2753,N_2692,N_2624);
and U2754 (N_2754,N_2600,N_2646);
xnor U2755 (N_2755,N_2683,N_2682);
and U2756 (N_2756,N_2687,N_2645);
nand U2757 (N_2757,N_2600,N_2605);
or U2758 (N_2758,N_2630,N_2663);
or U2759 (N_2759,N_2612,N_2679);
nand U2760 (N_2760,N_2610,N_2670);
nand U2761 (N_2761,N_2630,N_2645);
nand U2762 (N_2762,N_2660,N_2642);
xor U2763 (N_2763,N_2648,N_2650);
nand U2764 (N_2764,N_2613,N_2673);
and U2765 (N_2765,N_2698,N_2682);
or U2766 (N_2766,N_2662,N_2637);
nor U2767 (N_2767,N_2659,N_2680);
nand U2768 (N_2768,N_2619,N_2601);
nand U2769 (N_2769,N_2647,N_2619);
xor U2770 (N_2770,N_2692,N_2621);
xor U2771 (N_2771,N_2692,N_2634);
nor U2772 (N_2772,N_2654,N_2604);
nand U2773 (N_2773,N_2631,N_2669);
or U2774 (N_2774,N_2668,N_2617);
or U2775 (N_2775,N_2633,N_2673);
xnor U2776 (N_2776,N_2619,N_2692);
nor U2777 (N_2777,N_2618,N_2679);
xor U2778 (N_2778,N_2673,N_2688);
or U2779 (N_2779,N_2604,N_2632);
or U2780 (N_2780,N_2635,N_2659);
xor U2781 (N_2781,N_2663,N_2670);
and U2782 (N_2782,N_2696,N_2660);
nor U2783 (N_2783,N_2608,N_2620);
nand U2784 (N_2784,N_2622,N_2635);
nand U2785 (N_2785,N_2602,N_2665);
nand U2786 (N_2786,N_2666,N_2684);
nor U2787 (N_2787,N_2642,N_2628);
nand U2788 (N_2788,N_2675,N_2671);
xor U2789 (N_2789,N_2606,N_2632);
xor U2790 (N_2790,N_2640,N_2646);
xor U2791 (N_2791,N_2689,N_2609);
xnor U2792 (N_2792,N_2645,N_2664);
or U2793 (N_2793,N_2605,N_2607);
and U2794 (N_2794,N_2651,N_2619);
nand U2795 (N_2795,N_2613,N_2604);
or U2796 (N_2796,N_2615,N_2624);
nand U2797 (N_2797,N_2604,N_2602);
and U2798 (N_2798,N_2659,N_2643);
and U2799 (N_2799,N_2607,N_2646);
and U2800 (N_2800,N_2751,N_2730);
and U2801 (N_2801,N_2759,N_2763);
and U2802 (N_2802,N_2717,N_2772);
xor U2803 (N_2803,N_2733,N_2761);
or U2804 (N_2804,N_2754,N_2740);
or U2805 (N_2805,N_2705,N_2743);
nand U2806 (N_2806,N_2799,N_2735);
xnor U2807 (N_2807,N_2755,N_2715);
nor U2808 (N_2808,N_2798,N_2778);
xnor U2809 (N_2809,N_2702,N_2727);
or U2810 (N_2810,N_2708,N_2757);
nand U2811 (N_2811,N_2721,N_2775);
nor U2812 (N_2812,N_2732,N_2787);
nor U2813 (N_2813,N_2704,N_2771);
nor U2814 (N_2814,N_2790,N_2764);
nor U2815 (N_2815,N_2710,N_2776);
and U2816 (N_2816,N_2747,N_2700);
xor U2817 (N_2817,N_2737,N_2725);
nor U2818 (N_2818,N_2783,N_2788);
xor U2819 (N_2819,N_2709,N_2774);
nor U2820 (N_2820,N_2749,N_2716);
and U2821 (N_2821,N_2742,N_2728);
xnor U2822 (N_2822,N_2765,N_2729);
and U2823 (N_2823,N_2784,N_2760);
xnor U2824 (N_2824,N_2770,N_2748);
or U2825 (N_2825,N_2745,N_2756);
nor U2826 (N_2826,N_2794,N_2780);
or U2827 (N_2827,N_2722,N_2738);
nor U2828 (N_2828,N_2785,N_2723);
nand U2829 (N_2829,N_2758,N_2762);
and U2830 (N_2830,N_2718,N_2719);
and U2831 (N_2831,N_2731,N_2773);
xnor U2832 (N_2832,N_2782,N_2712);
xnor U2833 (N_2833,N_2766,N_2786);
nor U2834 (N_2834,N_2750,N_2720);
nor U2835 (N_2835,N_2789,N_2713);
and U2836 (N_2836,N_2781,N_2752);
xor U2837 (N_2837,N_2726,N_2707);
and U2838 (N_2838,N_2777,N_2724);
and U2839 (N_2839,N_2741,N_2746);
nand U2840 (N_2840,N_2744,N_2736);
and U2841 (N_2841,N_2793,N_2792);
and U2842 (N_2842,N_2768,N_2795);
xor U2843 (N_2843,N_2769,N_2703);
nor U2844 (N_2844,N_2753,N_2734);
and U2845 (N_2845,N_2767,N_2714);
nor U2846 (N_2846,N_2796,N_2706);
xnor U2847 (N_2847,N_2711,N_2739);
nand U2848 (N_2848,N_2779,N_2797);
or U2849 (N_2849,N_2701,N_2791);
nor U2850 (N_2850,N_2761,N_2787);
or U2851 (N_2851,N_2799,N_2746);
and U2852 (N_2852,N_2732,N_2768);
nand U2853 (N_2853,N_2755,N_2766);
nand U2854 (N_2854,N_2741,N_2775);
nand U2855 (N_2855,N_2745,N_2760);
and U2856 (N_2856,N_2726,N_2716);
xnor U2857 (N_2857,N_2720,N_2709);
xor U2858 (N_2858,N_2761,N_2755);
and U2859 (N_2859,N_2724,N_2716);
xor U2860 (N_2860,N_2784,N_2799);
and U2861 (N_2861,N_2705,N_2777);
and U2862 (N_2862,N_2799,N_2754);
or U2863 (N_2863,N_2799,N_2792);
nand U2864 (N_2864,N_2737,N_2782);
and U2865 (N_2865,N_2731,N_2758);
nor U2866 (N_2866,N_2733,N_2714);
xor U2867 (N_2867,N_2733,N_2794);
nand U2868 (N_2868,N_2768,N_2764);
nor U2869 (N_2869,N_2790,N_2785);
nor U2870 (N_2870,N_2784,N_2713);
and U2871 (N_2871,N_2735,N_2782);
nor U2872 (N_2872,N_2765,N_2723);
nor U2873 (N_2873,N_2795,N_2798);
xnor U2874 (N_2874,N_2732,N_2790);
xnor U2875 (N_2875,N_2724,N_2758);
or U2876 (N_2876,N_2747,N_2752);
and U2877 (N_2877,N_2711,N_2707);
or U2878 (N_2878,N_2735,N_2741);
nor U2879 (N_2879,N_2798,N_2750);
or U2880 (N_2880,N_2729,N_2728);
nand U2881 (N_2881,N_2757,N_2735);
nor U2882 (N_2882,N_2731,N_2781);
or U2883 (N_2883,N_2786,N_2749);
xnor U2884 (N_2884,N_2775,N_2720);
nand U2885 (N_2885,N_2717,N_2704);
xor U2886 (N_2886,N_2763,N_2740);
nand U2887 (N_2887,N_2713,N_2744);
and U2888 (N_2888,N_2791,N_2744);
nand U2889 (N_2889,N_2757,N_2772);
nor U2890 (N_2890,N_2799,N_2727);
and U2891 (N_2891,N_2787,N_2745);
xor U2892 (N_2892,N_2780,N_2748);
xnor U2893 (N_2893,N_2737,N_2773);
nor U2894 (N_2894,N_2743,N_2703);
nand U2895 (N_2895,N_2729,N_2788);
nor U2896 (N_2896,N_2701,N_2783);
or U2897 (N_2897,N_2701,N_2751);
nand U2898 (N_2898,N_2726,N_2741);
and U2899 (N_2899,N_2750,N_2742);
or U2900 (N_2900,N_2897,N_2815);
or U2901 (N_2901,N_2870,N_2805);
nor U2902 (N_2902,N_2842,N_2871);
nor U2903 (N_2903,N_2879,N_2819);
xnor U2904 (N_2904,N_2854,N_2835);
nor U2905 (N_2905,N_2881,N_2896);
nor U2906 (N_2906,N_2851,N_2872);
xor U2907 (N_2907,N_2804,N_2814);
nand U2908 (N_2908,N_2806,N_2843);
and U2909 (N_2909,N_2803,N_2811);
and U2910 (N_2910,N_2876,N_2863);
nand U2911 (N_2911,N_2891,N_2883);
and U2912 (N_2912,N_2867,N_2848);
and U2913 (N_2913,N_2887,N_2825);
nor U2914 (N_2914,N_2846,N_2834);
xor U2915 (N_2915,N_2895,N_2894);
and U2916 (N_2916,N_2885,N_2841);
and U2917 (N_2917,N_2807,N_2844);
nand U2918 (N_2918,N_2830,N_2817);
or U2919 (N_2919,N_2852,N_2833);
or U2920 (N_2920,N_2874,N_2882);
and U2921 (N_2921,N_2828,N_2838);
and U2922 (N_2922,N_2808,N_2816);
and U2923 (N_2923,N_2898,N_2827);
and U2924 (N_2924,N_2801,N_2878);
or U2925 (N_2925,N_2875,N_2864);
nor U2926 (N_2926,N_2866,N_2831);
and U2927 (N_2927,N_2893,N_2818);
or U2928 (N_2928,N_2809,N_2839);
xor U2929 (N_2929,N_2822,N_2892);
or U2930 (N_2930,N_2860,N_2889);
or U2931 (N_2931,N_2853,N_2812);
and U2932 (N_2932,N_2884,N_2861);
xnor U2933 (N_2933,N_2832,N_2890);
nand U2934 (N_2934,N_2836,N_2823);
xnor U2935 (N_2935,N_2855,N_2847);
or U2936 (N_2936,N_2869,N_2824);
nand U2937 (N_2937,N_2877,N_2840);
and U2938 (N_2938,N_2826,N_2845);
or U2939 (N_2939,N_2813,N_2821);
nand U2940 (N_2940,N_2829,N_2865);
xor U2941 (N_2941,N_2859,N_2873);
xnor U2942 (N_2942,N_2800,N_2850);
or U2943 (N_2943,N_2899,N_2886);
nor U2944 (N_2944,N_2880,N_2857);
nor U2945 (N_2945,N_2849,N_2856);
nor U2946 (N_2946,N_2810,N_2868);
nand U2947 (N_2947,N_2820,N_2888);
or U2948 (N_2948,N_2802,N_2837);
and U2949 (N_2949,N_2862,N_2858);
nor U2950 (N_2950,N_2849,N_2807);
nor U2951 (N_2951,N_2802,N_2882);
xor U2952 (N_2952,N_2829,N_2882);
nand U2953 (N_2953,N_2896,N_2876);
xnor U2954 (N_2954,N_2840,N_2825);
or U2955 (N_2955,N_2827,N_2884);
and U2956 (N_2956,N_2866,N_2833);
nor U2957 (N_2957,N_2883,N_2845);
or U2958 (N_2958,N_2896,N_2882);
nand U2959 (N_2959,N_2809,N_2834);
and U2960 (N_2960,N_2852,N_2894);
or U2961 (N_2961,N_2857,N_2861);
xnor U2962 (N_2962,N_2839,N_2820);
xor U2963 (N_2963,N_2897,N_2837);
xor U2964 (N_2964,N_2875,N_2894);
xnor U2965 (N_2965,N_2837,N_2824);
or U2966 (N_2966,N_2815,N_2837);
nand U2967 (N_2967,N_2843,N_2884);
xnor U2968 (N_2968,N_2841,N_2820);
nand U2969 (N_2969,N_2867,N_2892);
or U2970 (N_2970,N_2877,N_2891);
nor U2971 (N_2971,N_2829,N_2817);
xor U2972 (N_2972,N_2871,N_2883);
nor U2973 (N_2973,N_2890,N_2887);
and U2974 (N_2974,N_2849,N_2865);
or U2975 (N_2975,N_2834,N_2873);
nand U2976 (N_2976,N_2897,N_2805);
xnor U2977 (N_2977,N_2806,N_2873);
and U2978 (N_2978,N_2878,N_2822);
and U2979 (N_2979,N_2803,N_2849);
or U2980 (N_2980,N_2882,N_2897);
xnor U2981 (N_2981,N_2897,N_2860);
nand U2982 (N_2982,N_2829,N_2870);
or U2983 (N_2983,N_2895,N_2866);
xnor U2984 (N_2984,N_2891,N_2874);
or U2985 (N_2985,N_2877,N_2801);
nand U2986 (N_2986,N_2856,N_2838);
nor U2987 (N_2987,N_2810,N_2871);
and U2988 (N_2988,N_2836,N_2808);
nand U2989 (N_2989,N_2866,N_2868);
nor U2990 (N_2990,N_2874,N_2822);
and U2991 (N_2991,N_2889,N_2886);
xnor U2992 (N_2992,N_2860,N_2835);
nand U2993 (N_2993,N_2897,N_2838);
nand U2994 (N_2994,N_2852,N_2859);
or U2995 (N_2995,N_2840,N_2881);
nor U2996 (N_2996,N_2833,N_2814);
nand U2997 (N_2997,N_2834,N_2822);
nor U2998 (N_2998,N_2806,N_2831);
nand U2999 (N_2999,N_2899,N_2885);
and U3000 (N_3000,N_2914,N_2919);
and U3001 (N_3001,N_2955,N_2944);
and U3002 (N_3002,N_2931,N_2990);
or U3003 (N_3003,N_2941,N_2996);
nand U3004 (N_3004,N_2908,N_2976);
nand U3005 (N_3005,N_2937,N_2983);
nand U3006 (N_3006,N_2917,N_2992);
and U3007 (N_3007,N_2991,N_2902);
xor U3008 (N_3008,N_2966,N_2918);
or U3009 (N_3009,N_2995,N_2960);
xnor U3010 (N_3010,N_2988,N_2994);
nand U3011 (N_3011,N_2910,N_2925);
and U3012 (N_3012,N_2943,N_2926);
or U3013 (N_3013,N_2948,N_2975);
and U3014 (N_3014,N_2978,N_2911);
nand U3015 (N_3015,N_2924,N_2971);
xor U3016 (N_3016,N_2989,N_2905);
nor U3017 (N_3017,N_2950,N_2952);
and U3018 (N_3018,N_2979,N_2939);
xor U3019 (N_3019,N_2933,N_2974);
or U3020 (N_3020,N_2956,N_2915);
and U3021 (N_3021,N_2981,N_2945);
nor U3022 (N_3022,N_2977,N_2935);
xor U3023 (N_3023,N_2965,N_2970);
and U3024 (N_3024,N_2984,N_2936);
nand U3025 (N_3025,N_2982,N_2942);
nand U3026 (N_3026,N_2958,N_2972);
nor U3027 (N_3027,N_2929,N_2932);
or U3028 (N_3028,N_2923,N_2928);
or U3029 (N_3029,N_2946,N_2985);
and U3030 (N_3030,N_2969,N_2934);
or U3031 (N_3031,N_2987,N_2909);
xnor U3032 (N_3032,N_2903,N_2980);
or U3033 (N_3033,N_2951,N_2913);
or U3034 (N_3034,N_2959,N_2973);
nand U3035 (N_3035,N_2940,N_2998);
xnor U3036 (N_3036,N_2986,N_2901);
xor U3037 (N_3037,N_2947,N_2968);
nand U3038 (N_3038,N_2904,N_2900);
or U3039 (N_3039,N_2967,N_2916);
nand U3040 (N_3040,N_2962,N_2927);
xor U3041 (N_3041,N_2961,N_2993);
nand U3042 (N_3042,N_2938,N_2920);
and U3043 (N_3043,N_2957,N_2954);
nor U3044 (N_3044,N_2997,N_2999);
nand U3045 (N_3045,N_2906,N_2907);
nand U3046 (N_3046,N_2912,N_2953);
or U3047 (N_3047,N_2930,N_2964);
xor U3048 (N_3048,N_2921,N_2963);
nand U3049 (N_3049,N_2922,N_2949);
nand U3050 (N_3050,N_2989,N_2998);
and U3051 (N_3051,N_2941,N_2940);
or U3052 (N_3052,N_2987,N_2907);
xor U3053 (N_3053,N_2941,N_2958);
xor U3054 (N_3054,N_2961,N_2982);
and U3055 (N_3055,N_2922,N_2996);
nand U3056 (N_3056,N_2989,N_2997);
or U3057 (N_3057,N_2968,N_2953);
or U3058 (N_3058,N_2934,N_2996);
or U3059 (N_3059,N_2995,N_2905);
and U3060 (N_3060,N_2932,N_2942);
nor U3061 (N_3061,N_2929,N_2941);
xnor U3062 (N_3062,N_2905,N_2996);
xor U3063 (N_3063,N_2945,N_2955);
nor U3064 (N_3064,N_2996,N_2947);
or U3065 (N_3065,N_2980,N_2983);
or U3066 (N_3066,N_2995,N_2997);
and U3067 (N_3067,N_2959,N_2967);
or U3068 (N_3068,N_2973,N_2976);
nand U3069 (N_3069,N_2984,N_2993);
and U3070 (N_3070,N_2924,N_2956);
xnor U3071 (N_3071,N_2977,N_2937);
nand U3072 (N_3072,N_2937,N_2942);
and U3073 (N_3073,N_2972,N_2917);
or U3074 (N_3074,N_2983,N_2914);
nand U3075 (N_3075,N_2908,N_2951);
nand U3076 (N_3076,N_2946,N_2925);
or U3077 (N_3077,N_2942,N_2916);
and U3078 (N_3078,N_2966,N_2985);
xnor U3079 (N_3079,N_2975,N_2910);
nand U3080 (N_3080,N_2925,N_2957);
or U3081 (N_3081,N_2916,N_2985);
xnor U3082 (N_3082,N_2966,N_2916);
nand U3083 (N_3083,N_2923,N_2963);
or U3084 (N_3084,N_2956,N_2946);
nand U3085 (N_3085,N_2984,N_2918);
or U3086 (N_3086,N_2931,N_2922);
nor U3087 (N_3087,N_2938,N_2969);
and U3088 (N_3088,N_2980,N_2954);
xor U3089 (N_3089,N_2943,N_2934);
or U3090 (N_3090,N_2917,N_2911);
nand U3091 (N_3091,N_2968,N_2981);
and U3092 (N_3092,N_2992,N_2957);
nand U3093 (N_3093,N_2992,N_2924);
or U3094 (N_3094,N_2945,N_2948);
or U3095 (N_3095,N_2993,N_2998);
nand U3096 (N_3096,N_2951,N_2933);
xor U3097 (N_3097,N_2909,N_2919);
or U3098 (N_3098,N_2913,N_2966);
nor U3099 (N_3099,N_2958,N_2902);
and U3100 (N_3100,N_3004,N_3037);
nand U3101 (N_3101,N_3003,N_3094);
and U3102 (N_3102,N_3029,N_3049);
or U3103 (N_3103,N_3020,N_3001);
or U3104 (N_3104,N_3018,N_3015);
or U3105 (N_3105,N_3013,N_3023);
nand U3106 (N_3106,N_3071,N_3022);
or U3107 (N_3107,N_3079,N_3010);
nand U3108 (N_3108,N_3093,N_3057);
and U3109 (N_3109,N_3025,N_3055);
xor U3110 (N_3110,N_3048,N_3008);
nand U3111 (N_3111,N_3090,N_3081);
nand U3112 (N_3112,N_3042,N_3092);
xor U3113 (N_3113,N_3097,N_3085);
nand U3114 (N_3114,N_3051,N_3016);
xor U3115 (N_3115,N_3095,N_3083);
or U3116 (N_3116,N_3011,N_3005);
nor U3117 (N_3117,N_3087,N_3059);
xnor U3118 (N_3118,N_3098,N_3047);
nand U3119 (N_3119,N_3084,N_3044);
nor U3120 (N_3120,N_3034,N_3086);
and U3121 (N_3121,N_3056,N_3021);
nor U3122 (N_3122,N_3074,N_3028);
nor U3123 (N_3123,N_3075,N_3041);
nor U3124 (N_3124,N_3007,N_3082);
xnor U3125 (N_3125,N_3054,N_3027);
or U3126 (N_3126,N_3006,N_3096);
and U3127 (N_3127,N_3072,N_3060);
or U3128 (N_3128,N_3063,N_3050);
nand U3129 (N_3129,N_3067,N_3080);
nand U3130 (N_3130,N_3058,N_3032);
xor U3131 (N_3131,N_3066,N_3045);
nand U3132 (N_3132,N_3019,N_3052);
and U3133 (N_3133,N_3065,N_3062);
nand U3134 (N_3134,N_3069,N_3039);
nand U3135 (N_3135,N_3024,N_3064);
xnor U3136 (N_3136,N_3017,N_3043);
nand U3137 (N_3137,N_3070,N_3026);
nand U3138 (N_3138,N_3076,N_3012);
nor U3139 (N_3139,N_3046,N_3014);
and U3140 (N_3140,N_3030,N_3068);
xnor U3141 (N_3141,N_3073,N_3033);
and U3142 (N_3142,N_3035,N_3036);
nor U3143 (N_3143,N_3002,N_3089);
or U3144 (N_3144,N_3009,N_3088);
nor U3145 (N_3145,N_3038,N_3053);
nand U3146 (N_3146,N_3040,N_3099);
and U3147 (N_3147,N_3031,N_3077);
or U3148 (N_3148,N_3000,N_3091);
or U3149 (N_3149,N_3061,N_3078);
xnor U3150 (N_3150,N_3080,N_3094);
and U3151 (N_3151,N_3098,N_3082);
and U3152 (N_3152,N_3028,N_3000);
or U3153 (N_3153,N_3034,N_3045);
or U3154 (N_3154,N_3043,N_3026);
nor U3155 (N_3155,N_3057,N_3064);
and U3156 (N_3156,N_3096,N_3097);
or U3157 (N_3157,N_3032,N_3060);
nand U3158 (N_3158,N_3052,N_3028);
and U3159 (N_3159,N_3098,N_3076);
and U3160 (N_3160,N_3004,N_3057);
and U3161 (N_3161,N_3027,N_3036);
or U3162 (N_3162,N_3097,N_3019);
and U3163 (N_3163,N_3055,N_3005);
xor U3164 (N_3164,N_3039,N_3029);
and U3165 (N_3165,N_3025,N_3078);
xor U3166 (N_3166,N_3013,N_3015);
nand U3167 (N_3167,N_3082,N_3054);
nand U3168 (N_3168,N_3089,N_3086);
xnor U3169 (N_3169,N_3030,N_3037);
nand U3170 (N_3170,N_3068,N_3050);
nor U3171 (N_3171,N_3027,N_3032);
nor U3172 (N_3172,N_3085,N_3019);
nand U3173 (N_3173,N_3022,N_3030);
xor U3174 (N_3174,N_3020,N_3089);
nand U3175 (N_3175,N_3099,N_3096);
and U3176 (N_3176,N_3043,N_3022);
or U3177 (N_3177,N_3033,N_3065);
or U3178 (N_3178,N_3057,N_3028);
or U3179 (N_3179,N_3069,N_3027);
xnor U3180 (N_3180,N_3082,N_3066);
or U3181 (N_3181,N_3044,N_3043);
xor U3182 (N_3182,N_3063,N_3029);
nand U3183 (N_3183,N_3076,N_3069);
nor U3184 (N_3184,N_3077,N_3083);
nand U3185 (N_3185,N_3079,N_3055);
nor U3186 (N_3186,N_3011,N_3088);
nand U3187 (N_3187,N_3025,N_3064);
or U3188 (N_3188,N_3009,N_3069);
nand U3189 (N_3189,N_3034,N_3017);
and U3190 (N_3190,N_3004,N_3020);
and U3191 (N_3191,N_3016,N_3034);
nand U3192 (N_3192,N_3042,N_3004);
or U3193 (N_3193,N_3042,N_3028);
and U3194 (N_3194,N_3094,N_3067);
nand U3195 (N_3195,N_3066,N_3098);
nor U3196 (N_3196,N_3073,N_3020);
xor U3197 (N_3197,N_3019,N_3065);
nand U3198 (N_3198,N_3030,N_3032);
nand U3199 (N_3199,N_3093,N_3063);
xnor U3200 (N_3200,N_3129,N_3107);
xnor U3201 (N_3201,N_3190,N_3176);
or U3202 (N_3202,N_3116,N_3177);
xnor U3203 (N_3203,N_3148,N_3130);
nand U3204 (N_3204,N_3159,N_3134);
nand U3205 (N_3205,N_3150,N_3167);
nor U3206 (N_3206,N_3185,N_3135);
or U3207 (N_3207,N_3115,N_3164);
or U3208 (N_3208,N_3152,N_3181);
or U3209 (N_3209,N_3153,N_3145);
nor U3210 (N_3210,N_3121,N_3192);
nor U3211 (N_3211,N_3187,N_3126);
or U3212 (N_3212,N_3199,N_3131);
nor U3213 (N_3213,N_3162,N_3172);
nand U3214 (N_3214,N_3178,N_3195);
and U3215 (N_3215,N_3113,N_3171);
nand U3216 (N_3216,N_3109,N_3143);
nor U3217 (N_3217,N_3197,N_3166);
nor U3218 (N_3218,N_3139,N_3161);
and U3219 (N_3219,N_3111,N_3157);
nand U3220 (N_3220,N_3102,N_3198);
nor U3221 (N_3221,N_3169,N_3124);
and U3222 (N_3222,N_3158,N_3184);
and U3223 (N_3223,N_3179,N_3173);
or U3224 (N_3224,N_3141,N_3182);
or U3225 (N_3225,N_3138,N_3120);
xor U3226 (N_3226,N_3137,N_3183);
and U3227 (N_3227,N_3106,N_3105);
nand U3228 (N_3228,N_3142,N_3165);
nor U3229 (N_3229,N_3119,N_3117);
nor U3230 (N_3230,N_3175,N_3156);
xor U3231 (N_3231,N_3191,N_3140);
xor U3232 (N_3232,N_3104,N_3101);
xnor U3233 (N_3233,N_3194,N_3133);
xnor U3234 (N_3234,N_3163,N_3151);
and U3235 (N_3235,N_3189,N_3193);
nor U3236 (N_3236,N_3122,N_3144);
nor U3237 (N_3237,N_3149,N_3160);
and U3238 (N_3238,N_3174,N_3100);
nand U3239 (N_3239,N_3188,N_3168);
nand U3240 (N_3240,N_3125,N_3127);
or U3241 (N_3241,N_3155,N_3146);
xnor U3242 (N_3242,N_3114,N_3186);
or U3243 (N_3243,N_3103,N_3180);
nand U3244 (N_3244,N_3123,N_3196);
and U3245 (N_3245,N_3118,N_3108);
nand U3246 (N_3246,N_3110,N_3170);
and U3247 (N_3247,N_3128,N_3136);
or U3248 (N_3248,N_3112,N_3154);
and U3249 (N_3249,N_3147,N_3132);
or U3250 (N_3250,N_3162,N_3176);
nor U3251 (N_3251,N_3193,N_3179);
nor U3252 (N_3252,N_3167,N_3114);
nor U3253 (N_3253,N_3113,N_3105);
xor U3254 (N_3254,N_3139,N_3143);
and U3255 (N_3255,N_3194,N_3122);
nand U3256 (N_3256,N_3121,N_3138);
or U3257 (N_3257,N_3144,N_3179);
xnor U3258 (N_3258,N_3191,N_3179);
xnor U3259 (N_3259,N_3175,N_3180);
or U3260 (N_3260,N_3135,N_3194);
or U3261 (N_3261,N_3178,N_3169);
nand U3262 (N_3262,N_3178,N_3112);
xnor U3263 (N_3263,N_3196,N_3151);
and U3264 (N_3264,N_3115,N_3162);
xnor U3265 (N_3265,N_3172,N_3189);
or U3266 (N_3266,N_3179,N_3123);
nand U3267 (N_3267,N_3163,N_3149);
xnor U3268 (N_3268,N_3131,N_3158);
xnor U3269 (N_3269,N_3199,N_3111);
and U3270 (N_3270,N_3187,N_3136);
nor U3271 (N_3271,N_3106,N_3187);
xor U3272 (N_3272,N_3104,N_3135);
and U3273 (N_3273,N_3123,N_3194);
nand U3274 (N_3274,N_3146,N_3132);
or U3275 (N_3275,N_3159,N_3116);
nor U3276 (N_3276,N_3135,N_3112);
nor U3277 (N_3277,N_3148,N_3108);
or U3278 (N_3278,N_3182,N_3117);
or U3279 (N_3279,N_3179,N_3176);
nor U3280 (N_3280,N_3154,N_3130);
or U3281 (N_3281,N_3199,N_3118);
nor U3282 (N_3282,N_3131,N_3152);
nand U3283 (N_3283,N_3149,N_3151);
nor U3284 (N_3284,N_3172,N_3177);
nor U3285 (N_3285,N_3141,N_3164);
or U3286 (N_3286,N_3133,N_3113);
nand U3287 (N_3287,N_3144,N_3145);
nor U3288 (N_3288,N_3131,N_3198);
nand U3289 (N_3289,N_3118,N_3181);
xor U3290 (N_3290,N_3161,N_3183);
nor U3291 (N_3291,N_3129,N_3191);
and U3292 (N_3292,N_3193,N_3129);
xor U3293 (N_3293,N_3142,N_3146);
nand U3294 (N_3294,N_3168,N_3120);
nor U3295 (N_3295,N_3139,N_3149);
nor U3296 (N_3296,N_3132,N_3157);
xor U3297 (N_3297,N_3174,N_3134);
or U3298 (N_3298,N_3145,N_3122);
xor U3299 (N_3299,N_3110,N_3168);
nor U3300 (N_3300,N_3248,N_3249);
and U3301 (N_3301,N_3205,N_3219);
nor U3302 (N_3302,N_3212,N_3262);
and U3303 (N_3303,N_3220,N_3290);
xnor U3304 (N_3304,N_3261,N_3218);
or U3305 (N_3305,N_3228,N_3260);
xor U3306 (N_3306,N_3286,N_3253);
xor U3307 (N_3307,N_3276,N_3241);
nand U3308 (N_3308,N_3272,N_3294);
or U3309 (N_3309,N_3265,N_3250);
xor U3310 (N_3310,N_3298,N_3270);
and U3311 (N_3311,N_3239,N_3217);
nand U3312 (N_3312,N_3285,N_3213);
or U3313 (N_3313,N_3224,N_3207);
xnor U3314 (N_3314,N_3278,N_3259);
nor U3315 (N_3315,N_3245,N_3223);
nand U3316 (N_3316,N_3266,N_3226);
or U3317 (N_3317,N_3283,N_3273);
nand U3318 (N_3318,N_3268,N_3281);
nand U3319 (N_3319,N_3274,N_3234);
or U3320 (N_3320,N_3222,N_3277);
nor U3321 (N_3321,N_3208,N_3255);
and U3322 (N_3322,N_3257,N_3288);
xor U3323 (N_3323,N_3269,N_3236);
xnor U3324 (N_3324,N_3242,N_3204);
xnor U3325 (N_3325,N_3247,N_3292);
nor U3326 (N_3326,N_3252,N_3221);
nor U3327 (N_3327,N_3280,N_3206);
and U3328 (N_3328,N_3256,N_3264);
nand U3329 (N_3329,N_3232,N_3214);
nor U3330 (N_3330,N_3231,N_3287);
or U3331 (N_3331,N_3258,N_3295);
and U3332 (N_3332,N_3238,N_3297);
and U3333 (N_3333,N_3279,N_3209);
xnor U3334 (N_3334,N_3200,N_3230);
nand U3335 (N_3335,N_3251,N_3293);
or U3336 (N_3336,N_3240,N_3267);
nand U3337 (N_3337,N_3210,N_3233);
and U3338 (N_3338,N_3201,N_3237);
nand U3339 (N_3339,N_3263,N_3211);
xor U3340 (N_3340,N_3284,N_3202);
xnor U3341 (N_3341,N_3229,N_3244);
nand U3342 (N_3342,N_3216,N_3235);
xor U3343 (N_3343,N_3243,N_3275);
nand U3344 (N_3344,N_3271,N_3227);
nand U3345 (N_3345,N_3203,N_3296);
or U3346 (N_3346,N_3289,N_3225);
nor U3347 (N_3347,N_3299,N_3254);
xnor U3348 (N_3348,N_3282,N_3246);
xor U3349 (N_3349,N_3215,N_3291);
and U3350 (N_3350,N_3258,N_3297);
xnor U3351 (N_3351,N_3277,N_3224);
or U3352 (N_3352,N_3264,N_3217);
and U3353 (N_3353,N_3203,N_3211);
nor U3354 (N_3354,N_3203,N_3227);
or U3355 (N_3355,N_3231,N_3292);
and U3356 (N_3356,N_3238,N_3209);
and U3357 (N_3357,N_3224,N_3246);
xor U3358 (N_3358,N_3275,N_3260);
nor U3359 (N_3359,N_3219,N_3221);
nor U3360 (N_3360,N_3213,N_3264);
or U3361 (N_3361,N_3222,N_3238);
or U3362 (N_3362,N_3234,N_3292);
xnor U3363 (N_3363,N_3252,N_3261);
nor U3364 (N_3364,N_3288,N_3202);
nor U3365 (N_3365,N_3248,N_3255);
nand U3366 (N_3366,N_3225,N_3292);
nor U3367 (N_3367,N_3293,N_3210);
and U3368 (N_3368,N_3289,N_3235);
nand U3369 (N_3369,N_3238,N_3284);
xnor U3370 (N_3370,N_3263,N_3293);
or U3371 (N_3371,N_3277,N_3250);
nor U3372 (N_3372,N_3223,N_3259);
nor U3373 (N_3373,N_3284,N_3206);
nand U3374 (N_3374,N_3253,N_3250);
or U3375 (N_3375,N_3289,N_3236);
or U3376 (N_3376,N_3221,N_3291);
and U3377 (N_3377,N_3295,N_3202);
nand U3378 (N_3378,N_3277,N_3262);
xnor U3379 (N_3379,N_3285,N_3242);
and U3380 (N_3380,N_3293,N_3228);
and U3381 (N_3381,N_3276,N_3232);
nand U3382 (N_3382,N_3242,N_3216);
nand U3383 (N_3383,N_3240,N_3257);
nor U3384 (N_3384,N_3298,N_3242);
xnor U3385 (N_3385,N_3238,N_3248);
or U3386 (N_3386,N_3217,N_3284);
nor U3387 (N_3387,N_3210,N_3264);
nand U3388 (N_3388,N_3253,N_3275);
nand U3389 (N_3389,N_3200,N_3240);
nor U3390 (N_3390,N_3241,N_3250);
nor U3391 (N_3391,N_3225,N_3242);
or U3392 (N_3392,N_3288,N_3205);
and U3393 (N_3393,N_3249,N_3253);
and U3394 (N_3394,N_3269,N_3297);
xor U3395 (N_3395,N_3289,N_3255);
or U3396 (N_3396,N_3240,N_3232);
and U3397 (N_3397,N_3274,N_3264);
nand U3398 (N_3398,N_3260,N_3269);
or U3399 (N_3399,N_3246,N_3248);
and U3400 (N_3400,N_3334,N_3343);
xnor U3401 (N_3401,N_3392,N_3331);
nand U3402 (N_3402,N_3371,N_3303);
xor U3403 (N_3403,N_3338,N_3341);
or U3404 (N_3404,N_3370,N_3358);
nor U3405 (N_3405,N_3380,N_3352);
nor U3406 (N_3406,N_3368,N_3376);
xnor U3407 (N_3407,N_3357,N_3348);
and U3408 (N_3408,N_3329,N_3372);
or U3409 (N_3409,N_3311,N_3325);
xor U3410 (N_3410,N_3328,N_3353);
xor U3411 (N_3411,N_3318,N_3345);
and U3412 (N_3412,N_3387,N_3342);
or U3413 (N_3413,N_3332,N_3366);
and U3414 (N_3414,N_3308,N_3374);
or U3415 (N_3415,N_3326,N_3309);
and U3416 (N_3416,N_3373,N_3322);
xnor U3417 (N_3417,N_3384,N_3363);
nand U3418 (N_3418,N_3347,N_3360);
and U3419 (N_3419,N_3354,N_3385);
or U3420 (N_3420,N_3333,N_3365);
xor U3421 (N_3421,N_3382,N_3351);
xor U3422 (N_3422,N_3302,N_3317);
or U3423 (N_3423,N_3324,N_3316);
nand U3424 (N_3424,N_3340,N_3301);
or U3425 (N_3425,N_3398,N_3327);
xnor U3426 (N_3426,N_3336,N_3391);
and U3427 (N_3427,N_3397,N_3355);
nor U3428 (N_3428,N_3349,N_3344);
or U3429 (N_3429,N_3396,N_3362);
nand U3430 (N_3430,N_3381,N_3304);
or U3431 (N_3431,N_3364,N_3350);
nand U3432 (N_3432,N_3300,N_3389);
and U3433 (N_3433,N_3367,N_3395);
and U3434 (N_3434,N_3359,N_3323);
and U3435 (N_3435,N_3388,N_3306);
xnor U3436 (N_3436,N_3399,N_3369);
or U3437 (N_3437,N_3337,N_3313);
or U3438 (N_3438,N_3335,N_3320);
and U3439 (N_3439,N_3375,N_3393);
nor U3440 (N_3440,N_3330,N_3390);
xnor U3441 (N_3441,N_3394,N_3310);
and U3442 (N_3442,N_3307,N_3361);
or U3443 (N_3443,N_3315,N_3386);
and U3444 (N_3444,N_3319,N_3356);
and U3445 (N_3445,N_3305,N_3339);
nand U3446 (N_3446,N_3321,N_3379);
nor U3447 (N_3447,N_3383,N_3314);
nor U3448 (N_3448,N_3378,N_3346);
nor U3449 (N_3449,N_3312,N_3377);
and U3450 (N_3450,N_3379,N_3358);
or U3451 (N_3451,N_3303,N_3366);
and U3452 (N_3452,N_3361,N_3341);
nand U3453 (N_3453,N_3336,N_3397);
nand U3454 (N_3454,N_3390,N_3324);
and U3455 (N_3455,N_3381,N_3324);
nor U3456 (N_3456,N_3333,N_3371);
or U3457 (N_3457,N_3388,N_3309);
or U3458 (N_3458,N_3332,N_3311);
and U3459 (N_3459,N_3361,N_3351);
and U3460 (N_3460,N_3355,N_3395);
and U3461 (N_3461,N_3394,N_3309);
or U3462 (N_3462,N_3367,N_3342);
nand U3463 (N_3463,N_3335,N_3337);
nor U3464 (N_3464,N_3326,N_3313);
or U3465 (N_3465,N_3399,N_3364);
nand U3466 (N_3466,N_3301,N_3334);
xor U3467 (N_3467,N_3397,N_3315);
nand U3468 (N_3468,N_3338,N_3382);
or U3469 (N_3469,N_3356,N_3382);
nor U3470 (N_3470,N_3333,N_3330);
nor U3471 (N_3471,N_3340,N_3360);
or U3472 (N_3472,N_3353,N_3321);
xnor U3473 (N_3473,N_3351,N_3379);
nand U3474 (N_3474,N_3377,N_3324);
and U3475 (N_3475,N_3341,N_3311);
and U3476 (N_3476,N_3324,N_3334);
nand U3477 (N_3477,N_3317,N_3378);
or U3478 (N_3478,N_3346,N_3371);
nand U3479 (N_3479,N_3358,N_3399);
xnor U3480 (N_3480,N_3346,N_3362);
nand U3481 (N_3481,N_3354,N_3328);
and U3482 (N_3482,N_3375,N_3358);
nand U3483 (N_3483,N_3336,N_3321);
nor U3484 (N_3484,N_3312,N_3325);
nand U3485 (N_3485,N_3323,N_3373);
xnor U3486 (N_3486,N_3346,N_3317);
and U3487 (N_3487,N_3324,N_3387);
xor U3488 (N_3488,N_3331,N_3342);
or U3489 (N_3489,N_3351,N_3347);
and U3490 (N_3490,N_3366,N_3370);
and U3491 (N_3491,N_3359,N_3388);
or U3492 (N_3492,N_3368,N_3395);
or U3493 (N_3493,N_3399,N_3336);
nand U3494 (N_3494,N_3391,N_3308);
xnor U3495 (N_3495,N_3398,N_3390);
nor U3496 (N_3496,N_3310,N_3354);
and U3497 (N_3497,N_3378,N_3380);
nor U3498 (N_3498,N_3339,N_3382);
nand U3499 (N_3499,N_3379,N_3378);
or U3500 (N_3500,N_3468,N_3400);
xor U3501 (N_3501,N_3498,N_3408);
and U3502 (N_3502,N_3457,N_3492);
xor U3503 (N_3503,N_3433,N_3421);
or U3504 (N_3504,N_3440,N_3409);
and U3505 (N_3505,N_3414,N_3489);
and U3506 (N_3506,N_3424,N_3485);
nand U3507 (N_3507,N_3472,N_3434);
nand U3508 (N_3508,N_3451,N_3436);
and U3509 (N_3509,N_3464,N_3448);
nor U3510 (N_3510,N_3419,N_3403);
nand U3511 (N_3511,N_3474,N_3449);
and U3512 (N_3512,N_3453,N_3402);
or U3513 (N_3513,N_3450,N_3423);
or U3514 (N_3514,N_3454,N_3428);
nor U3515 (N_3515,N_3435,N_3469);
or U3516 (N_3516,N_3482,N_3405);
nand U3517 (N_3517,N_3456,N_3486);
xor U3518 (N_3518,N_3415,N_3430);
nand U3519 (N_3519,N_3404,N_3459);
nand U3520 (N_3520,N_3446,N_3426);
xnor U3521 (N_3521,N_3470,N_3483);
xnor U3522 (N_3522,N_3427,N_3493);
nand U3523 (N_3523,N_3425,N_3491);
or U3524 (N_3524,N_3438,N_3475);
xor U3525 (N_3525,N_3447,N_3477);
nor U3526 (N_3526,N_3478,N_3429);
nand U3527 (N_3527,N_3439,N_3437);
nor U3528 (N_3528,N_3413,N_3467);
nand U3529 (N_3529,N_3466,N_3444);
nand U3530 (N_3530,N_3499,N_3443);
or U3531 (N_3531,N_3417,N_3490);
nand U3532 (N_3532,N_3445,N_3494);
or U3533 (N_3533,N_3442,N_3488);
and U3534 (N_3534,N_3431,N_3497);
nor U3535 (N_3535,N_3411,N_3432);
nand U3536 (N_3536,N_3471,N_3458);
and U3537 (N_3537,N_3496,N_3418);
or U3538 (N_3538,N_3420,N_3412);
xor U3539 (N_3539,N_3473,N_3407);
or U3540 (N_3540,N_3460,N_3416);
nand U3541 (N_3541,N_3479,N_3476);
xnor U3542 (N_3542,N_3481,N_3487);
nand U3543 (N_3543,N_3452,N_3455);
or U3544 (N_3544,N_3463,N_3441);
nor U3545 (N_3545,N_3480,N_3462);
and U3546 (N_3546,N_3406,N_3465);
xor U3547 (N_3547,N_3422,N_3484);
and U3548 (N_3548,N_3495,N_3401);
and U3549 (N_3549,N_3410,N_3461);
xor U3550 (N_3550,N_3445,N_3433);
xor U3551 (N_3551,N_3477,N_3436);
nand U3552 (N_3552,N_3430,N_3471);
xnor U3553 (N_3553,N_3489,N_3458);
xnor U3554 (N_3554,N_3408,N_3429);
nor U3555 (N_3555,N_3423,N_3457);
nor U3556 (N_3556,N_3464,N_3456);
and U3557 (N_3557,N_3424,N_3489);
and U3558 (N_3558,N_3454,N_3493);
xnor U3559 (N_3559,N_3411,N_3422);
or U3560 (N_3560,N_3483,N_3486);
xnor U3561 (N_3561,N_3412,N_3437);
nand U3562 (N_3562,N_3462,N_3475);
and U3563 (N_3563,N_3469,N_3455);
or U3564 (N_3564,N_3494,N_3405);
nor U3565 (N_3565,N_3439,N_3433);
or U3566 (N_3566,N_3486,N_3409);
and U3567 (N_3567,N_3406,N_3462);
or U3568 (N_3568,N_3487,N_3456);
nand U3569 (N_3569,N_3494,N_3427);
or U3570 (N_3570,N_3450,N_3498);
or U3571 (N_3571,N_3440,N_3490);
nand U3572 (N_3572,N_3467,N_3452);
and U3573 (N_3573,N_3491,N_3448);
and U3574 (N_3574,N_3438,N_3432);
nand U3575 (N_3575,N_3421,N_3402);
nor U3576 (N_3576,N_3421,N_3417);
xor U3577 (N_3577,N_3496,N_3482);
nor U3578 (N_3578,N_3476,N_3411);
xor U3579 (N_3579,N_3427,N_3432);
nor U3580 (N_3580,N_3480,N_3430);
xnor U3581 (N_3581,N_3414,N_3419);
and U3582 (N_3582,N_3478,N_3459);
nor U3583 (N_3583,N_3494,N_3470);
nor U3584 (N_3584,N_3439,N_3454);
xor U3585 (N_3585,N_3415,N_3477);
or U3586 (N_3586,N_3415,N_3470);
xnor U3587 (N_3587,N_3487,N_3435);
and U3588 (N_3588,N_3436,N_3487);
nor U3589 (N_3589,N_3453,N_3416);
and U3590 (N_3590,N_3458,N_3413);
and U3591 (N_3591,N_3413,N_3469);
and U3592 (N_3592,N_3418,N_3465);
nor U3593 (N_3593,N_3400,N_3411);
and U3594 (N_3594,N_3404,N_3485);
and U3595 (N_3595,N_3477,N_3480);
nor U3596 (N_3596,N_3457,N_3479);
xor U3597 (N_3597,N_3430,N_3458);
xor U3598 (N_3598,N_3419,N_3496);
and U3599 (N_3599,N_3492,N_3444);
or U3600 (N_3600,N_3568,N_3590);
and U3601 (N_3601,N_3553,N_3529);
or U3602 (N_3602,N_3560,N_3559);
nor U3603 (N_3603,N_3526,N_3569);
and U3604 (N_3604,N_3510,N_3574);
xor U3605 (N_3605,N_3594,N_3506);
or U3606 (N_3606,N_3592,N_3501);
and U3607 (N_3607,N_3538,N_3585);
or U3608 (N_3608,N_3583,N_3502);
nand U3609 (N_3609,N_3561,N_3579);
nand U3610 (N_3610,N_3557,N_3528);
or U3611 (N_3611,N_3537,N_3581);
and U3612 (N_3612,N_3500,N_3556);
or U3613 (N_3613,N_3575,N_3512);
and U3614 (N_3614,N_3563,N_3566);
xnor U3615 (N_3615,N_3535,N_3588);
nand U3616 (N_3616,N_3562,N_3518);
or U3617 (N_3617,N_3533,N_3513);
nand U3618 (N_3618,N_3520,N_3564);
nand U3619 (N_3619,N_3525,N_3571);
nor U3620 (N_3620,N_3573,N_3546);
xor U3621 (N_3621,N_3584,N_3554);
and U3622 (N_3622,N_3555,N_3534);
nand U3623 (N_3623,N_3565,N_3552);
xnor U3624 (N_3624,N_3595,N_3541);
and U3625 (N_3625,N_3547,N_3543);
and U3626 (N_3626,N_3540,N_3527);
or U3627 (N_3627,N_3567,N_3530);
or U3628 (N_3628,N_3515,N_3548);
and U3629 (N_3629,N_3545,N_3522);
nand U3630 (N_3630,N_3516,N_3558);
or U3631 (N_3631,N_3532,N_3536);
nor U3632 (N_3632,N_3578,N_3591);
nor U3633 (N_3633,N_3531,N_3596);
and U3634 (N_3634,N_3586,N_3544);
nor U3635 (N_3635,N_3508,N_3509);
and U3636 (N_3636,N_3505,N_3549);
or U3637 (N_3637,N_3503,N_3519);
and U3638 (N_3638,N_3580,N_3514);
and U3639 (N_3639,N_3523,N_3570);
and U3640 (N_3640,N_3517,N_3598);
and U3641 (N_3641,N_3593,N_3504);
and U3642 (N_3642,N_3524,N_3511);
nand U3643 (N_3643,N_3582,N_3576);
and U3644 (N_3644,N_3597,N_3587);
or U3645 (N_3645,N_3550,N_3507);
or U3646 (N_3646,N_3577,N_3521);
xnor U3647 (N_3647,N_3589,N_3539);
nor U3648 (N_3648,N_3599,N_3551);
nor U3649 (N_3649,N_3572,N_3542);
or U3650 (N_3650,N_3566,N_3540);
nand U3651 (N_3651,N_3545,N_3588);
and U3652 (N_3652,N_3590,N_3575);
nor U3653 (N_3653,N_3584,N_3576);
nor U3654 (N_3654,N_3500,N_3561);
xnor U3655 (N_3655,N_3528,N_3508);
xnor U3656 (N_3656,N_3558,N_3571);
xnor U3657 (N_3657,N_3532,N_3597);
or U3658 (N_3658,N_3557,N_3540);
nor U3659 (N_3659,N_3510,N_3560);
or U3660 (N_3660,N_3512,N_3508);
nand U3661 (N_3661,N_3519,N_3505);
and U3662 (N_3662,N_3541,N_3506);
and U3663 (N_3663,N_3509,N_3536);
xor U3664 (N_3664,N_3594,N_3556);
and U3665 (N_3665,N_3582,N_3512);
or U3666 (N_3666,N_3564,N_3540);
nor U3667 (N_3667,N_3530,N_3584);
nor U3668 (N_3668,N_3593,N_3514);
nand U3669 (N_3669,N_3525,N_3543);
nand U3670 (N_3670,N_3530,N_3524);
and U3671 (N_3671,N_3516,N_3559);
or U3672 (N_3672,N_3519,N_3526);
and U3673 (N_3673,N_3586,N_3582);
and U3674 (N_3674,N_3533,N_3558);
and U3675 (N_3675,N_3580,N_3539);
nand U3676 (N_3676,N_3536,N_3538);
xor U3677 (N_3677,N_3571,N_3538);
nand U3678 (N_3678,N_3509,N_3576);
nand U3679 (N_3679,N_3530,N_3571);
xnor U3680 (N_3680,N_3518,N_3567);
or U3681 (N_3681,N_3572,N_3588);
and U3682 (N_3682,N_3582,N_3506);
nand U3683 (N_3683,N_3559,N_3542);
nand U3684 (N_3684,N_3562,N_3539);
nand U3685 (N_3685,N_3573,N_3552);
and U3686 (N_3686,N_3574,N_3584);
nor U3687 (N_3687,N_3537,N_3501);
nor U3688 (N_3688,N_3567,N_3509);
or U3689 (N_3689,N_3596,N_3504);
nand U3690 (N_3690,N_3577,N_3571);
xor U3691 (N_3691,N_3533,N_3502);
nor U3692 (N_3692,N_3512,N_3520);
nand U3693 (N_3693,N_3544,N_3500);
nor U3694 (N_3694,N_3561,N_3571);
and U3695 (N_3695,N_3524,N_3590);
or U3696 (N_3696,N_3516,N_3511);
nand U3697 (N_3697,N_3514,N_3520);
xor U3698 (N_3698,N_3581,N_3586);
nor U3699 (N_3699,N_3562,N_3558);
nor U3700 (N_3700,N_3694,N_3671);
or U3701 (N_3701,N_3676,N_3628);
nand U3702 (N_3702,N_3607,N_3673);
or U3703 (N_3703,N_3654,N_3661);
xnor U3704 (N_3704,N_3687,N_3655);
and U3705 (N_3705,N_3615,N_3613);
nor U3706 (N_3706,N_3681,N_3636);
and U3707 (N_3707,N_3685,N_3651);
nor U3708 (N_3708,N_3619,N_3639);
nor U3709 (N_3709,N_3674,N_3689);
nor U3710 (N_3710,N_3611,N_3646);
nor U3711 (N_3711,N_3677,N_3643);
xor U3712 (N_3712,N_3668,N_3605);
xor U3713 (N_3713,N_3645,N_3641);
nand U3714 (N_3714,N_3672,N_3663);
nand U3715 (N_3715,N_3631,N_3610);
xor U3716 (N_3716,N_3601,N_3640);
xor U3717 (N_3717,N_3644,N_3632);
nand U3718 (N_3718,N_3683,N_3647);
xor U3719 (N_3719,N_3626,N_3684);
xor U3720 (N_3720,N_3692,N_3603);
xnor U3721 (N_3721,N_3696,N_3670);
nand U3722 (N_3722,N_3667,N_3648);
nand U3723 (N_3723,N_3693,N_3690);
nor U3724 (N_3724,N_3642,N_3635);
nor U3725 (N_3725,N_3633,N_3669);
nor U3726 (N_3726,N_3618,N_3627);
nor U3727 (N_3727,N_3698,N_3609);
nor U3728 (N_3728,N_3662,N_3617);
nand U3729 (N_3729,N_3675,N_3659);
nor U3730 (N_3730,N_3604,N_3602);
nor U3731 (N_3731,N_3620,N_3630);
xnor U3732 (N_3732,N_3680,N_3634);
xnor U3733 (N_3733,N_3614,N_3688);
xnor U3734 (N_3734,N_3697,N_3678);
xor U3735 (N_3735,N_3652,N_3699);
nand U3736 (N_3736,N_3649,N_3629);
and U3737 (N_3737,N_3657,N_3600);
or U3738 (N_3738,N_3612,N_3665);
nor U3739 (N_3739,N_3606,N_3625);
and U3740 (N_3740,N_3622,N_3691);
and U3741 (N_3741,N_3679,N_3637);
nor U3742 (N_3742,N_3686,N_3653);
nor U3743 (N_3743,N_3695,N_3666);
nor U3744 (N_3744,N_3616,N_3650);
xor U3745 (N_3745,N_3621,N_3682);
nand U3746 (N_3746,N_3664,N_3624);
and U3747 (N_3747,N_3658,N_3660);
xnor U3748 (N_3748,N_3608,N_3623);
nor U3749 (N_3749,N_3656,N_3638);
nand U3750 (N_3750,N_3690,N_3686);
xor U3751 (N_3751,N_3678,N_3688);
and U3752 (N_3752,N_3646,N_3609);
and U3753 (N_3753,N_3652,N_3666);
nand U3754 (N_3754,N_3661,N_3675);
nor U3755 (N_3755,N_3602,N_3667);
and U3756 (N_3756,N_3621,N_3604);
xor U3757 (N_3757,N_3644,N_3619);
nor U3758 (N_3758,N_3626,N_3622);
xnor U3759 (N_3759,N_3632,N_3650);
or U3760 (N_3760,N_3653,N_3671);
nand U3761 (N_3761,N_3622,N_3674);
or U3762 (N_3762,N_3614,N_3684);
nor U3763 (N_3763,N_3600,N_3635);
and U3764 (N_3764,N_3637,N_3646);
nor U3765 (N_3765,N_3689,N_3627);
xnor U3766 (N_3766,N_3622,N_3644);
or U3767 (N_3767,N_3608,N_3643);
and U3768 (N_3768,N_3695,N_3649);
nor U3769 (N_3769,N_3622,N_3665);
and U3770 (N_3770,N_3645,N_3636);
xnor U3771 (N_3771,N_3615,N_3658);
xnor U3772 (N_3772,N_3603,N_3684);
xnor U3773 (N_3773,N_3631,N_3680);
and U3774 (N_3774,N_3621,N_3653);
and U3775 (N_3775,N_3668,N_3691);
nor U3776 (N_3776,N_3655,N_3683);
and U3777 (N_3777,N_3654,N_3672);
and U3778 (N_3778,N_3693,N_3611);
and U3779 (N_3779,N_3621,N_3633);
nor U3780 (N_3780,N_3620,N_3644);
xnor U3781 (N_3781,N_3698,N_3668);
nor U3782 (N_3782,N_3652,N_3600);
xnor U3783 (N_3783,N_3648,N_3651);
nand U3784 (N_3784,N_3666,N_3645);
nand U3785 (N_3785,N_3662,N_3642);
nand U3786 (N_3786,N_3631,N_3632);
xor U3787 (N_3787,N_3637,N_3611);
nor U3788 (N_3788,N_3650,N_3601);
nor U3789 (N_3789,N_3677,N_3642);
or U3790 (N_3790,N_3600,N_3625);
nor U3791 (N_3791,N_3625,N_3660);
nor U3792 (N_3792,N_3641,N_3629);
nand U3793 (N_3793,N_3685,N_3690);
nor U3794 (N_3794,N_3600,N_3631);
xor U3795 (N_3795,N_3690,N_3689);
nor U3796 (N_3796,N_3659,N_3613);
nor U3797 (N_3797,N_3616,N_3623);
nand U3798 (N_3798,N_3611,N_3617);
and U3799 (N_3799,N_3602,N_3612);
and U3800 (N_3800,N_3762,N_3714);
and U3801 (N_3801,N_3733,N_3797);
xnor U3802 (N_3802,N_3771,N_3786);
and U3803 (N_3803,N_3787,N_3779);
xor U3804 (N_3804,N_3773,N_3725);
nand U3805 (N_3805,N_3750,N_3777);
nand U3806 (N_3806,N_3778,N_3723);
xor U3807 (N_3807,N_3713,N_3781);
and U3808 (N_3808,N_3728,N_3768);
and U3809 (N_3809,N_3716,N_3755);
xor U3810 (N_3810,N_3794,N_3754);
or U3811 (N_3811,N_3718,N_3737);
or U3812 (N_3812,N_3784,N_3705);
nand U3813 (N_3813,N_3747,N_3709);
and U3814 (N_3814,N_3701,N_3711);
or U3815 (N_3815,N_3706,N_3772);
and U3816 (N_3816,N_3799,N_3795);
xnor U3817 (N_3817,N_3782,N_3769);
nand U3818 (N_3818,N_3788,N_3746);
xor U3819 (N_3819,N_3798,N_3757);
or U3820 (N_3820,N_3745,N_3702);
nor U3821 (N_3821,N_3722,N_3761);
xnor U3822 (N_3822,N_3790,N_3738);
nor U3823 (N_3823,N_3708,N_3776);
and U3824 (N_3824,N_3748,N_3796);
xnor U3825 (N_3825,N_3707,N_3780);
nor U3826 (N_3826,N_3726,N_3720);
nand U3827 (N_3827,N_3793,N_3749);
nor U3828 (N_3828,N_3710,N_3730);
or U3829 (N_3829,N_3700,N_3727);
xnor U3830 (N_3830,N_3765,N_3717);
nor U3831 (N_3831,N_3766,N_3715);
or U3832 (N_3832,N_3736,N_3752);
and U3833 (N_3833,N_3734,N_3763);
or U3834 (N_3834,N_3742,N_3744);
or U3835 (N_3835,N_3751,N_3719);
xor U3836 (N_3836,N_3785,N_3764);
nor U3837 (N_3837,N_3724,N_3792);
nand U3838 (N_3838,N_3756,N_3703);
xor U3839 (N_3839,N_3741,N_3775);
nor U3840 (N_3840,N_3729,N_3791);
or U3841 (N_3841,N_3739,N_3770);
nor U3842 (N_3842,N_3767,N_3732);
nand U3843 (N_3843,N_3758,N_3760);
xor U3844 (N_3844,N_3740,N_3704);
nand U3845 (N_3845,N_3759,N_3731);
and U3846 (N_3846,N_3753,N_3743);
xnor U3847 (N_3847,N_3774,N_3789);
or U3848 (N_3848,N_3721,N_3735);
nand U3849 (N_3849,N_3783,N_3712);
and U3850 (N_3850,N_3701,N_3786);
nand U3851 (N_3851,N_3721,N_3786);
or U3852 (N_3852,N_3797,N_3722);
and U3853 (N_3853,N_3743,N_3778);
and U3854 (N_3854,N_3768,N_3729);
or U3855 (N_3855,N_3785,N_3771);
or U3856 (N_3856,N_3786,N_3774);
nor U3857 (N_3857,N_3741,N_3782);
nand U3858 (N_3858,N_3726,N_3735);
or U3859 (N_3859,N_3757,N_3774);
nor U3860 (N_3860,N_3781,N_3706);
or U3861 (N_3861,N_3722,N_3759);
or U3862 (N_3862,N_3767,N_3766);
nor U3863 (N_3863,N_3735,N_3702);
xor U3864 (N_3864,N_3744,N_3771);
nand U3865 (N_3865,N_3705,N_3767);
and U3866 (N_3866,N_3708,N_3793);
and U3867 (N_3867,N_3799,N_3769);
and U3868 (N_3868,N_3765,N_3703);
nand U3869 (N_3869,N_3798,N_3712);
or U3870 (N_3870,N_3766,N_3798);
nand U3871 (N_3871,N_3784,N_3725);
and U3872 (N_3872,N_3781,N_3724);
xnor U3873 (N_3873,N_3767,N_3789);
nand U3874 (N_3874,N_3766,N_3737);
and U3875 (N_3875,N_3714,N_3774);
and U3876 (N_3876,N_3788,N_3742);
nand U3877 (N_3877,N_3727,N_3788);
xor U3878 (N_3878,N_3799,N_3741);
and U3879 (N_3879,N_3736,N_3791);
xor U3880 (N_3880,N_3736,N_3794);
xor U3881 (N_3881,N_3789,N_3749);
nand U3882 (N_3882,N_3722,N_3795);
nand U3883 (N_3883,N_3751,N_3736);
or U3884 (N_3884,N_3767,N_3758);
nand U3885 (N_3885,N_3777,N_3771);
and U3886 (N_3886,N_3773,N_3768);
and U3887 (N_3887,N_3734,N_3748);
and U3888 (N_3888,N_3737,N_3781);
xor U3889 (N_3889,N_3716,N_3770);
or U3890 (N_3890,N_3725,N_3778);
xor U3891 (N_3891,N_3780,N_3729);
xor U3892 (N_3892,N_3706,N_3713);
and U3893 (N_3893,N_3752,N_3773);
nor U3894 (N_3894,N_3764,N_3753);
nor U3895 (N_3895,N_3795,N_3784);
and U3896 (N_3896,N_3739,N_3718);
nor U3897 (N_3897,N_3753,N_3744);
nand U3898 (N_3898,N_3741,N_3781);
nand U3899 (N_3899,N_3753,N_3720);
or U3900 (N_3900,N_3846,N_3889);
and U3901 (N_3901,N_3823,N_3826);
nor U3902 (N_3902,N_3875,N_3837);
nand U3903 (N_3903,N_3842,N_3880);
nand U3904 (N_3904,N_3829,N_3862);
nor U3905 (N_3905,N_3854,N_3899);
and U3906 (N_3906,N_3845,N_3805);
nor U3907 (N_3907,N_3873,N_3856);
or U3908 (N_3908,N_3897,N_3841);
nand U3909 (N_3909,N_3881,N_3809);
and U3910 (N_3910,N_3840,N_3872);
nand U3911 (N_3911,N_3863,N_3825);
nand U3912 (N_3912,N_3808,N_3814);
nand U3913 (N_3913,N_3839,N_3869);
nand U3914 (N_3914,N_3815,N_3851);
nand U3915 (N_3915,N_3857,N_3894);
nand U3916 (N_3916,N_3813,N_3865);
or U3917 (N_3917,N_3828,N_3818);
or U3918 (N_3918,N_3852,N_3895);
and U3919 (N_3919,N_3870,N_3855);
nand U3920 (N_3920,N_3896,N_3801);
and U3921 (N_3921,N_3876,N_3866);
xnor U3922 (N_3922,N_3860,N_3830);
xnor U3923 (N_3923,N_3804,N_3827);
or U3924 (N_3924,N_3891,N_3848);
or U3925 (N_3925,N_3893,N_3832);
and U3926 (N_3926,N_3835,N_3802);
xor U3927 (N_3927,N_3824,N_3838);
xor U3928 (N_3928,N_3864,N_3820);
or U3929 (N_3929,N_3859,N_3887);
xor U3930 (N_3930,N_3885,N_3877);
and U3931 (N_3931,N_3850,N_3834);
nand U3932 (N_3932,N_3831,N_3874);
nand U3933 (N_3933,N_3858,N_3811);
nor U3934 (N_3934,N_3879,N_3817);
or U3935 (N_3935,N_3812,N_3822);
and U3936 (N_3936,N_3833,N_3884);
nand U3937 (N_3937,N_3847,N_3871);
and U3938 (N_3938,N_3810,N_3867);
nand U3939 (N_3939,N_3836,N_3844);
nor U3940 (N_3940,N_3821,N_3886);
nor U3941 (N_3941,N_3861,N_3888);
nor U3942 (N_3942,N_3890,N_3807);
nand U3943 (N_3943,N_3800,N_3853);
nand U3944 (N_3944,N_3878,N_3898);
nand U3945 (N_3945,N_3868,N_3819);
xnor U3946 (N_3946,N_3803,N_3816);
or U3947 (N_3947,N_3843,N_3882);
nor U3948 (N_3948,N_3892,N_3806);
and U3949 (N_3949,N_3883,N_3849);
nor U3950 (N_3950,N_3842,N_3835);
and U3951 (N_3951,N_3848,N_3874);
xnor U3952 (N_3952,N_3850,N_3862);
nand U3953 (N_3953,N_3807,N_3880);
and U3954 (N_3954,N_3890,N_3872);
nor U3955 (N_3955,N_3864,N_3821);
or U3956 (N_3956,N_3822,N_3846);
or U3957 (N_3957,N_3899,N_3814);
nand U3958 (N_3958,N_3899,N_3896);
nand U3959 (N_3959,N_3875,N_3865);
nand U3960 (N_3960,N_3824,N_3873);
or U3961 (N_3961,N_3833,N_3888);
nand U3962 (N_3962,N_3858,N_3833);
and U3963 (N_3963,N_3859,N_3813);
nand U3964 (N_3964,N_3817,N_3858);
and U3965 (N_3965,N_3834,N_3842);
or U3966 (N_3966,N_3818,N_3821);
or U3967 (N_3967,N_3886,N_3882);
and U3968 (N_3968,N_3889,N_3894);
or U3969 (N_3969,N_3818,N_3825);
xor U3970 (N_3970,N_3840,N_3878);
or U3971 (N_3971,N_3851,N_3808);
or U3972 (N_3972,N_3843,N_3885);
nor U3973 (N_3973,N_3848,N_3802);
xor U3974 (N_3974,N_3875,N_3854);
nand U3975 (N_3975,N_3829,N_3825);
nand U3976 (N_3976,N_3887,N_3883);
or U3977 (N_3977,N_3851,N_3826);
nor U3978 (N_3978,N_3841,N_3801);
xnor U3979 (N_3979,N_3822,N_3826);
and U3980 (N_3980,N_3839,N_3854);
nand U3981 (N_3981,N_3810,N_3804);
nand U3982 (N_3982,N_3840,N_3818);
xnor U3983 (N_3983,N_3802,N_3826);
or U3984 (N_3984,N_3843,N_3896);
and U3985 (N_3985,N_3860,N_3841);
nand U3986 (N_3986,N_3857,N_3815);
nor U3987 (N_3987,N_3882,N_3821);
nor U3988 (N_3988,N_3811,N_3812);
nor U3989 (N_3989,N_3838,N_3852);
and U3990 (N_3990,N_3851,N_3854);
or U3991 (N_3991,N_3870,N_3892);
nor U3992 (N_3992,N_3852,N_3800);
xnor U3993 (N_3993,N_3889,N_3845);
nand U3994 (N_3994,N_3816,N_3897);
xnor U3995 (N_3995,N_3825,N_3831);
xor U3996 (N_3996,N_3856,N_3876);
and U3997 (N_3997,N_3836,N_3853);
nor U3998 (N_3998,N_3864,N_3858);
nor U3999 (N_3999,N_3878,N_3856);
nand U4000 (N_4000,N_3900,N_3963);
nand U4001 (N_4001,N_3970,N_3935);
nand U4002 (N_4002,N_3955,N_3967);
xor U4003 (N_4003,N_3979,N_3916);
xor U4004 (N_4004,N_3998,N_3927);
nor U4005 (N_4005,N_3990,N_3992);
nor U4006 (N_4006,N_3971,N_3912);
nand U4007 (N_4007,N_3949,N_3987);
xnor U4008 (N_4008,N_3968,N_3903);
nand U4009 (N_4009,N_3993,N_3953);
nand U4010 (N_4010,N_3928,N_3997);
xor U4011 (N_4011,N_3984,N_3961);
and U4012 (N_4012,N_3924,N_3937);
xnor U4013 (N_4013,N_3918,N_3904);
and U4014 (N_4014,N_3948,N_3950);
xnor U4015 (N_4015,N_3983,N_3995);
nor U4016 (N_4016,N_3914,N_3908);
xor U4017 (N_4017,N_3945,N_3939);
nor U4018 (N_4018,N_3958,N_3905);
nor U4019 (N_4019,N_3994,N_3952);
and U4020 (N_4020,N_3956,N_3943);
nand U4021 (N_4021,N_3969,N_3941);
xor U4022 (N_4022,N_3986,N_3921);
and U4023 (N_4023,N_3960,N_3981);
xnor U4024 (N_4024,N_3965,N_3902);
or U4025 (N_4025,N_3944,N_3996);
xor U4026 (N_4026,N_3988,N_3947);
xor U4027 (N_4027,N_3982,N_3913);
nand U4028 (N_4028,N_3917,N_3951);
nand U4029 (N_4029,N_3932,N_3959);
and U4030 (N_4030,N_3980,N_3938);
and U4031 (N_4031,N_3972,N_3942);
and U4032 (N_4032,N_3966,N_3925);
nand U4033 (N_4033,N_3930,N_3975);
nor U4034 (N_4034,N_3906,N_3929);
xor U4035 (N_4035,N_3919,N_3985);
or U4036 (N_4036,N_3991,N_3926);
xor U4037 (N_4037,N_3931,N_3957);
nand U4038 (N_4038,N_3933,N_3920);
xnor U4039 (N_4039,N_3911,N_3954);
and U4040 (N_4040,N_3946,N_3962);
or U4041 (N_4041,N_3973,N_3909);
or U4042 (N_4042,N_3989,N_3907);
nand U4043 (N_4043,N_3976,N_3974);
nor U4044 (N_4044,N_3934,N_3999);
nand U4045 (N_4045,N_3964,N_3936);
xor U4046 (N_4046,N_3910,N_3922);
or U4047 (N_4047,N_3923,N_3978);
nand U4048 (N_4048,N_3940,N_3915);
nand U4049 (N_4049,N_3901,N_3977);
xnor U4050 (N_4050,N_3960,N_3988);
nor U4051 (N_4051,N_3907,N_3944);
or U4052 (N_4052,N_3970,N_3960);
xnor U4053 (N_4053,N_3947,N_3977);
nor U4054 (N_4054,N_3901,N_3907);
nor U4055 (N_4055,N_3933,N_3942);
nand U4056 (N_4056,N_3907,N_3949);
xnor U4057 (N_4057,N_3919,N_3934);
and U4058 (N_4058,N_3984,N_3968);
xor U4059 (N_4059,N_3941,N_3915);
nor U4060 (N_4060,N_3980,N_3988);
and U4061 (N_4061,N_3910,N_3926);
and U4062 (N_4062,N_3966,N_3924);
nand U4063 (N_4063,N_3923,N_3980);
nor U4064 (N_4064,N_3917,N_3939);
nor U4065 (N_4065,N_3986,N_3979);
nor U4066 (N_4066,N_3908,N_3928);
nor U4067 (N_4067,N_3994,N_3932);
and U4068 (N_4068,N_3920,N_3963);
or U4069 (N_4069,N_3991,N_3982);
xor U4070 (N_4070,N_3968,N_3944);
nand U4071 (N_4071,N_3968,N_3912);
xnor U4072 (N_4072,N_3964,N_3961);
xor U4073 (N_4073,N_3952,N_3907);
nand U4074 (N_4074,N_3974,N_3996);
nand U4075 (N_4075,N_3952,N_3927);
nor U4076 (N_4076,N_3935,N_3933);
nor U4077 (N_4077,N_3971,N_3939);
xnor U4078 (N_4078,N_3908,N_3972);
or U4079 (N_4079,N_3930,N_3921);
xnor U4080 (N_4080,N_3989,N_3955);
nand U4081 (N_4081,N_3970,N_3979);
or U4082 (N_4082,N_3994,N_3943);
and U4083 (N_4083,N_3941,N_3903);
and U4084 (N_4084,N_3959,N_3958);
xor U4085 (N_4085,N_3946,N_3975);
nand U4086 (N_4086,N_3932,N_3969);
or U4087 (N_4087,N_3983,N_3999);
and U4088 (N_4088,N_3945,N_3926);
or U4089 (N_4089,N_3995,N_3925);
nor U4090 (N_4090,N_3976,N_3956);
nor U4091 (N_4091,N_3931,N_3932);
or U4092 (N_4092,N_3997,N_3998);
nor U4093 (N_4093,N_3943,N_3972);
nor U4094 (N_4094,N_3986,N_3953);
nand U4095 (N_4095,N_3978,N_3907);
nor U4096 (N_4096,N_3920,N_3916);
and U4097 (N_4097,N_3990,N_3956);
nand U4098 (N_4098,N_3927,N_3987);
nor U4099 (N_4099,N_3972,N_3978);
and U4100 (N_4100,N_4049,N_4017);
nor U4101 (N_4101,N_4004,N_4053);
nand U4102 (N_4102,N_4058,N_4016);
xor U4103 (N_4103,N_4061,N_4085);
or U4104 (N_4104,N_4025,N_4042);
nand U4105 (N_4105,N_4092,N_4034);
nand U4106 (N_4106,N_4005,N_4048);
nor U4107 (N_4107,N_4037,N_4050);
nor U4108 (N_4108,N_4008,N_4014);
nand U4109 (N_4109,N_4038,N_4010);
nand U4110 (N_4110,N_4075,N_4015);
xor U4111 (N_4111,N_4044,N_4072);
xor U4112 (N_4112,N_4094,N_4097);
nand U4113 (N_4113,N_4003,N_4023);
or U4114 (N_4114,N_4096,N_4082);
xnor U4115 (N_4115,N_4059,N_4027);
nor U4116 (N_4116,N_4039,N_4099);
or U4117 (N_4117,N_4046,N_4036);
nand U4118 (N_4118,N_4095,N_4056);
or U4119 (N_4119,N_4089,N_4011);
nand U4120 (N_4120,N_4024,N_4071);
nor U4121 (N_4121,N_4043,N_4000);
nand U4122 (N_4122,N_4081,N_4063);
xor U4123 (N_4123,N_4078,N_4076);
and U4124 (N_4124,N_4084,N_4021);
xnor U4125 (N_4125,N_4031,N_4077);
nor U4126 (N_4126,N_4060,N_4088);
nor U4127 (N_4127,N_4013,N_4057);
and U4128 (N_4128,N_4029,N_4098);
nor U4129 (N_4129,N_4086,N_4041);
nor U4130 (N_4130,N_4035,N_4090);
nor U4131 (N_4131,N_4070,N_4074);
or U4132 (N_4132,N_4066,N_4064);
nand U4133 (N_4133,N_4093,N_4067);
xnor U4134 (N_4134,N_4001,N_4083);
and U4135 (N_4135,N_4002,N_4055);
and U4136 (N_4136,N_4012,N_4026);
nand U4137 (N_4137,N_4052,N_4032);
xnor U4138 (N_4138,N_4079,N_4006);
xor U4139 (N_4139,N_4065,N_4087);
nand U4140 (N_4140,N_4009,N_4091);
nand U4141 (N_4141,N_4045,N_4080);
nor U4142 (N_4142,N_4007,N_4028);
nor U4143 (N_4143,N_4062,N_4030);
and U4144 (N_4144,N_4040,N_4073);
and U4145 (N_4145,N_4047,N_4068);
xnor U4146 (N_4146,N_4069,N_4019);
nor U4147 (N_4147,N_4022,N_4051);
xnor U4148 (N_4148,N_4020,N_4033);
nor U4149 (N_4149,N_4018,N_4054);
nor U4150 (N_4150,N_4057,N_4030);
and U4151 (N_4151,N_4022,N_4088);
nand U4152 (N_4152,N_4094,N_4037);
nand U4153 (N_4153,N_4078,N_4095);
xnor U4154 (N_4154,N_4070,N_4075);
xor U4155 (N_4155,N_4039,N_4057);
and U4156 (N_4156,N_4035,N_4083);
or U4157 (N_4157,N_4049,N_4057);
and U4158 (N_4158,N_4065,N_4009);
nor U4159 (N_4159,N_4077,N_4011);
or U4160 (N_4160,N_4069,N_4060);
nor U4161 (N_4161,N_4099,N_4010);
and U4162 (N_4162,N_4076,N_4077);
and U4163 (N_4163,N_4024,N_4012);
xor U4164 (N_4164,N_4037,N_4075);
and U4165 (N_4165,N_4025,N_4019);
xor U4166 (N_4166,N_4093,N_4052);
nor U4167 (N_4167,N_4043,N_4039);
and U4168 (N_4168,N_4090,N_4060);
or U4169 (N_4169,N_4099,N_4041);
nor U4170 (N_4170,N_4034,N_4008);
xor U4171 (N_4171,N_4010,N_4072);
or U4172 (N_4172,N_4004,N_4079);
nand U4173 (N_4173,N_4021,N_4069);
and U4174 (N_4174,N_4070,N_4015);
xor U4175 (N_4175,N_4065,N_4091);
or U4176 (N_4176,N_4007,N_4004);
xor U4177 (N_4177,N_4051,N_4094);
nor U4178 (N_4178,N_4098,N_4010);
nand U4179 (N_4179,N_4057,N_4040);
nor U4180 (N_4180,N_4039,N_4031);
and U4181 (N_4181,N_4018,N_4056);
xor U4182 (N_4182,N_4090,N_4025);
nand U4183 (N_4183,N_4076,N_4064);
nand U4184 (N_4184,N_4029,N_4085);
nor U4185 (N_4185,N_4066,N_4098);
and U4186 (N_4186,N_4014,N_4079);
nor U4187 (N_4187,N_4034,N_4007);
nand U4188 (N_4188,N_4057,N_4095);
or U4189 (N_4189,N_4094,N_4010);
nand U4190 (N_4190,N_4078,N_4054);
xor U4191 (N_4191,N_4059,N_4025);
nor U4192 (N_4192,N_4003,N_4071);
and U4193 (N_4193,N_4037,N_4068);
nand U4194 (N_4194,N_4076,N_4061);
nand U4195 (N_4195,N_4062,N_4025);
and U4196 (N_4196,N_4044,N_4016);
or U4197 (N_4197,N_4071,N_4088);
and U4198 (N_4198,N_4019,N_4008);
and U4199 (N_4199,N_4009,N_4049);
xnor U4200 (N_4200,N_4100,N_4111);
or U4201 (N_4201,N_4183,N_4156);
nor U4202 (N_4202,N_4113,N_4178);
xor U4203 (N_4203,N_4146,N_4166);
xnor U4204 (N_4204,N_4180,N_4137);
xnor U4205 (N_4205,N_4124,N_4196);
nand U4206 (N_4206,N_4109,N_4186);
nand U4207 (N_4207,N_4167,N_4134);
nand U4208 (N_4208,N_4139,N_4135);
or U4209 (N_4209,N_4132,N_4157);
or U4210 (N_4210,N_4129,N_4116);
nor U4211 (N_4211,N_4120,N_4171);
and U4212 (N_4212,N_4150,N_4189);
xor U4213 (N_4213,N_4114,N_4187);
xor U4214 (N_4214,N_4182,N_4142);
nand U4215 (N_4215,N_4194,N_4147);
and U4216 (N_4216,N_4172,N_4105);
nand U4217 (N_4217,N_4122,N_4136);
nor U4218 (N_4218,N_4127,N_4123);
nor U4219 (N_4219,N_4153,N_4121);
or U4220 (N_4220,N_4162,N_4191);
and U4221 (N_4221,N_4101,N_4154);
xor U4222 (N_4222,N_4141,N_4179);
xnor U4223 (N_4223,N_4148,N_4174);
xor U4224 (N_4224,N_4128,N_4192);
nor U4225 (N_4225,N_4133,N_4130);
or U4226 (N_4226,N_4149,N_4199);
nand U4227 (N_4227,N_4138,N_4158);
and U4228 (N_4228,N_4119,N_4185);
nand U4229 (N_4229,N_4131,N_4125);
nand U4230 (N_4230,N_4106,N_4144);
nor U4231 (N_4231,N_4195,N_4181);
nand U4232 (N_4232,N_4159,N_4126);
xnor U4233 (N_4233,N_4173,N_4163);
nand U4234 (N_4234,N_4103,N_4161);
nor U4235 (N_4235,N_4104,N_4112);
xnor U4236 (N_4236,N_4169,N_4152);
or U4237 (N_4237,N_4175,N_4108);
or U4238 (N_4238,N_4176,N_4110);
nor U4239 (N_4239,N_4165,N_4188);
or U4240 (N_4240,N_4168,N_4118);
and U4241 (N_4241,N_4198,N_4145);
or U4242 (N_4242,N_4193,N_4155);
nor U4243 (N_4243,N_4184,N_4151);
nor U4244 (N_4244,N_4164,N_4170);
nor U4245 (N_4245,N_4177,N_4197);
or U4246 (N_4246,N_4102,N_4117);
xnor U4247 (N_4247,N_4143,N_4115);
nor U4248 (N_4248,N_4160,N_4140);
nor U4249 (N_4249,N_4107,N_4190);
or U4250 (N_4250,N_4155,N_4180);
or U4251 (N_4251,N_4199,N_4116);
nor U4252 (N_4252,N_4193,N_4132);
nor U4253 (N_4253,N_4148,N_4157);
nand U4254 (N_4254,N_4154,N_4140);
or U4255 (N_4255,N_4182,N_4146);
and U4256 (N_4256,N_4135,N_4132);
xor U4257 (N_4257,N_4178,N_4126);
and U4258 (N_4258,N_4175,N_4144);
and U4259 (N_4259,N_4178,N_4132);
or U4260 (N_4260,N_4150,N_4105);
nand U4261 (N_4261,N_4165,N_4117);
nor U4262 (N_4262,N_4181,N_4170);
and U4263 (N_4263,N_4111,N_4129);
and U4264 (N_4264,N_4105,N_4155);
or U4265 (N_4265,N_4134,N_4152);
or U4266 (N_4266,N_4198,N_4192);
or U4267 (N_4267,N_4122,N_4175);
xor U4268 (N_4268,N_4157,N_4188);
and U4269 (N_4269,N_4176,N_4138);
xor U4270 (N_4270,N_4187,N_4169);
xnor U4271 (N_4271,N_4114,N_4115);
or U4272 (N_4272,N_4146,N_4199);
and U4273 (N_4273,N_4126,N_4137);
and U4274 (N_4274,N_4176,N_4115);
nand U4275 (N_4275,N_4127,N_4115);
nand U4276 (N_4276,N_4171,N_4150);
nor U4277 (N_4277,N_4103,N_4134);
xor U4278 (N_4278,N_4167,N_4172);
nor U4279 (N_4279,N_4196,N_4125);
and U4280 (N_4280,N_4195,N_4103);
nand U4281 (N_4281,N_4110,N_4114);
nor U4282 (N_4282,N_4155,N_4157);
nand U4283 (N_4283,N_4172,N_4176);
nor U4284 (N_4284,N_4110,N_4198);
nor U4285 (N_4285,N_4139,N_4146);
or U4286 (N_4286,N_4126,N_4183);
nor U4287 (N_4287,N_4102,N_4184);
xor U4288 (N_4288,N_4195,N_4173);
nand U4289 (N_4289,N_4169,N_4166);
and U4290 (N_4290,N_4106,N_4170);
xor U4291 (N_4291,N_4186,N_4139);
xnor U4292 (N_4292,N_4156,N_4117);
xnor U4293 (N_4293,N_4146,N_4151);
or U4294 (N_4294,N_4168,N_4169);
xor U4295 (N_4295,N_4146,N_4130);
or U4296 (N_4296,N_4169,N_4131);
or U4297 (N_4297,N_4173,N_4133);
and U4298 (N_4298,N_4198,N_4138);
nor U4299 (N_4299,N_4148,N_4133);
or U4300 (N_4300,N_4214,N_4238);
and U4301 (N_4301,N_4261,N_4218);
nand U4302 (N_4302,N_4241,N_4230);
and U4303 (N_4303,N_4232,N_4296);
xnor U4304 (N_4304,N_4297,N_4226);
xor U4305 (N_4305,N_4250,N_4248);
or U4306 (N_4306,N_4253,N_4270);
and U4307 (N_4307,N_4206,N_4245);
nor U4308 (N_4308,N_4260,N_4262);
nand U4309 (N_4309,N_4224,N_4235);
nor U4310 (N_4310,N_4294,N_4280);
and U4311 (N_4311,N_4283,N_4279);
xnor U4312 (N_4312,N_4292,N_4263);
nor U4313 (N_4313,N_4220,N_4289);
and U4314 (N_4314,N_4287,N_4210);
xnor U4315 (N_4315,N_4255,N_4272);
xnor U4316 (N_4316,N_4200,N_4237);
and U4317 (N_4317,N_4221,N_4205);
xnor U4318 (N_4318,N_4229,N_4222);
nand U4319 (N_4319,N_4265,N_4201);
and U4320 (N_4320,N_4251,N_4290);
or U4321 (N_4321,N_4268,N_4285);
nor U4322 (N_4322,N_4247,N_4249);
and U4323 (N_4323,N_4213,N_4225);
nor U4324 (N_4324,N_4239,N_4208);
xor U4325 (N_4325,N_4273,N_4286);
nand U4326 (N_4326,N_4298,N_4291);
nor U4327 (N_4327,N_4257,N_4254);
nand U4328 (N_4328,N_4234,N_4227);
xor U4329 (N_4329,N_4211,N_4275);
xor U4330 (N_4330,N_4278,N_4259);
nor U4331 (N_4331,N_4240,N_4203);
xnor U4332 (N_4332,N_4209,N_4244);
or U4333 (N_4333,N_4276,N_4284);
xor U4334 (N_4334,N_4264,N_4223);
nor U4335 (N_4335,N_4267,N_4246);
or U4336 (N_4336,N_4299,N_4231);
or U4337 (N_4337,N_4271,N_4233);
nand U4338 (N_4338,N_4281,N_4288);
xnor U4339 (N_4339,N_4269,N_4219);
nand U4340 (N_4340,N_4277,N_4258);
xnor U4341 (N_4341,N_4217,N_4207);
and U4342 (N_4342,N_4243,N_4274);
nand U4343 (N_4343,N_4242,N_4216);
and U4344 (N_4344,N_4282,N_4204);
or U4345 (N_4345,N_4228,N_4252);
and U4346 (N_4346,N_4202,N_4266);
or U4347 (N_4347,N_4236,N_4293);
and U4348 (N_4348,N_4295,N_4215);
and U4349 (N_4349,N_4212,N_4256);
xor U4350 (N_4350,N_4207,N_4293);
xnor U4351 (N_4351,N_4256,N_4259);
and U4352 (N_4352,N_4255,N_4214);
or U4353 (N_4353,N_4227,N_4275);
or U4354 (N_4354,N_4206,N_4257);
xnor U4355 (N_4355,N_4213,N_4270);
nor U4356 (N_4356,N_4248,N_4253);
or U4357 (N_4357,N_4275,N_4201);
nor U4358 (N_4358,N_4269,N_4298);
nor U4359 (N_4359,N_4260,N_4254);
nand U4360 (N_4360,N_4247,N_4239);
xnor U4361 (N_4361,N_4221,N_4216);
or U4362 (N_4362,N_4211,N_4231);
or U4363 (N_4363,N_4283,N_4284);
nand U4364 (N_4364,N_4254,N_4216);
or U4365 (N_4365,N_4204,N_4213);
and U4366 (N_4366,N_4213,N_4281);
and U4367 (N_4367,N_4287,N_4258);
or U4368 (N_4368,N_4245,N_4269);
nand U4369 (N_4369,N_4227,N_4219);
nand U4370 (N_4370,N_4230,N_4208);
nand U4371 (N_4371,N_4204,N_4228);
xnor U4372 (N_4372,N_4249,N_4293);
nand U4373 (N_4373,N_4244,N_4242);
nor U4374 (N_4374,N_4238,N_4288);
nor U4375 (N_4375,N_4269,N_4251);
nand U4376 (N_4376,N_4280,N_4276);
nand U4377 (N_4377,N_4274,N_4240);
or U4378 (N_4378,N_4287,N_4247);
nor U4379 (N_4379,N_4289,N_4273);
and U4380 (N_4380,N_4208,N_4295);
or U4381 (N_4381,N_4287,N_4286);
or U4382 (N_4382,N_4290,N_4293);
nor U4383 (N_4383,N_4229,N_4285);
xor U4384 (N_4384,N_4277,N_4267);
nand U4385 (N_4385,N_4271,N_4273);
or U4386 (N_4386,N_4292,N_4237);
xnor U4387 (N_4387,N_4229,N_4246);
nand U4388 (N_4388,N_4253,N_4233);
xnor U4389 (N_4389,N_4217,N_4234);
and U4390 (N_4390,N_4293,N_4211);
xor U4391 (N_4391,N_4279,N_4213);
or U4392 (N_4392,N_4257,N_4222);
nor U4393 (N_4393,N_4268,N_4279);
nand U4394 (N_4394,N_4200,N_4233);
or U4395 (N_4395,N_4240,N_4221);
or U4396 (N_4396,N_4271,N_4249);
xnor U4397 (N_4397,N_4274,N_4232);
nor U4398 (N_4398,N_4282,N_4258);
nand U4399 (N_4399,N_4255,N_4200);
nor U4400 (N_4400,N_4344,N_4356);
nor U4401 (N_4401,N_4300,N_4398);
xnor U4402 (N_4402,N_4330,N_4351);
nor U4403 (N_4403,N_4369,N_4381);
and U4404 (N_4404,N_4342,N_4331);
nand U4405 (N_4405,N_4317,N_4375);
xnor U4406 (N_4406,N_4347,N_4348);
xnor U4407 (N_4407,N_4307,N_4388);
xor U4408 (N_4408,N_4350,N_4380);
xor U4409 (N_4409,N_4349,N_4314);
nor U4410 (N_4410,N_4385,N_4316);
and U4411 (N_4411,N_4305,N_4357);
nand U4412 (N_4412,N_4333,N_4318);
and U4413 (N_4413,N_4336,N_4361);
xor U4414 (N_4414,N_4335,N_4309);
or U4415 (N_4415,N_4395,N_4358);
nor U4416 (N_4416,N_4332,N_4327);
and U4417 (N_4417,N_4387,N_4377);
nor U4418 (N_4418,N_4338,N_4399);
and U4419 (N_4419,N_4319,N_4306);
nor U4420 (N_4420,N_4322,N_4312);
nor U4421 (N_4421,N_4325,N_4382);
and U4422 (N_4422,N_4311,N_4374);
or U4423 (N_4423,N_4334,N_4362);
nor U4424 (N_4424,N_4301,N_4313);
xnor U4425 (N_4425,N_4364,N_4368);
nor U4426 (N_4426,N_4339,N_4355);
or U4427 (N_4427,N_4366,N_4376);
and U4428 (N_4428,N_4341,N_4384);
nor U4429 (N_4429,N_4326,N_4337);
and U4430 (N_4430,N_4359,N_4304);
or U4431 (N_4431,N_4393,N_4320);
nor U4432 (N_4432,N_4352,N_4363);
xnor U4433 (N_4433,N_4371,N_4310);
nor U4434 (N_4434,N_4340,N_4343);
and U4435 (N_4435,N_4346,N_4386);
xnor U4436 (N_4436,N_4365,N_4345);
xor U4437 (N_4437,N_4373,N_4303);
nand U4438 (N_4438,N_4367,N_4390);
or U4439 (N_4439,N_4383,N_4328);
nor U4440 (N_4440,N_4379,N_4324);
or U4441 (N_4441,N_4360,N_4315);
nand U4442 (N_4442,N_4392,N_4378);
nor U4443 (N_4443,N_4321,N_4329);
xnor U4444 (N_4444,N_4394,N_4391);
or U4445 (N_4445,N_4372,N_4308);
or U4446 (N_4446,N_4354,N_4323);
nor U4447 (N_4447,N_4353,N_4397);
nor U4448 (N_4448,N_4302,N_4370);
or U4449 (N_4449,N_4396,N_4389);
nor U4450 (N_4450,N_4356,N_4323);
xor U4451 (N_4451,N_4325,N_4307);
nor U4452 (N_4452,N_4394,N_4312);
or U4453 (N_4453,N_4328,N_4346);
nand U4454 (N_4454,N_4306,N_4335);
or U4455 (N_4455,N_4353,N_4321);
nand U4456 (N_4456,N_4349,N_4344);
nor U4457 (N_4457,N_4324,N_4363);
or U4458 (N_4458,N_4312,N_4307);
and U4459 (N_4459,N_4310,N_4354);
and U4460 (N_4460,N_4339,N_4321);
nor U4461 (N_4461,N_4334,N_4361);
and U4462 (N_4462,N_4313,N_4338);
nor U4463 (N_4463,N_4304,N_4329);
and U4464 (N_4464,N_4313,N_4305);
and U4465 (N_4465,N_4346,N_4303);
xor U4466 (N_4466,N_4350,N_4301);
nor U4467 (N_4467,N_4388,N_4346);
nand U4468 (N_4468,N_4393,N_4357);
nor U4469 (N_4469,N_4356,N_4396);
xnor U4470 (N_4470,N_4361,N_4321);
or U4471 (N_4471,N_4378,N_4371);
or U4472 (N_4472,N_4306,N_4379);
xor U4473 (N_4473,N_4389,N_4301);
nand U4474 (N_4474,N_4360,N_4386);
xor U4475 (N_4475,N_4303,N_4326);
nor U4476 (N_4476,N_4375,N_4321);
and U4477 (N_4477,N_4332,N_4354);
or U4478 (N_4478,N_4320,N_4384);
or U4479 (N_4479,N_4326,N_4312);
or U4480 (N_4480,N_4359,N_4306);
xnor U4481 (N_4481,N_4388,N_4383);
nor U4482 (N_4482,N_4354,N_4338);
xor U4483 (N_4483,N_4371,N_4363);
xnor U4484 (N_4484,N_4384,N_4304);
xnor U4485 (N_4485,N_4300,N_4307);
or U4486 (N_4486,N_4309,N_4307);
nor U4487 (N_4487,N_4382,N_4346);
nor U4488 (N_4488,N_4345,N_4315);
nand U4489 (N_4489,N_4352,N_4348);
and U4490 (N_4490,N_4380,N_4382);
or U4491 (N_4491,N_4376,N_4354);
nand U4492 (N_4492,N_4334,N_4370);
or U4493 (N_4493,N_4350,N_4341);
or U4494 (N_4494,N_4393,N_4315);
xor U4495 (N_4495,N_4309,N_4337);
or U4496 (N_4496,N_4366,N_4367);
xor U4497 (N_4497,N_4392,N_4307);
nand U4498 (N_4498,N_4312,N_4366);
nor U4499 (N_4499,N_4342,N_4373);
nor U4500 (N_4500,N_4487,N_4478);
or U4501 (N_4501,N_4423,N_4435);
xor U4502 (N_4502,N_4426,N_4410);
and U4503 (N_4503,N_4469,N_4477);
and U4504 (N_4504,N_4405,N_4489);
xor U4505 (N_4505,N_4453,N_4488);
nor U4506 (N_4506,N_4436,N_4474);
and U4507 (N_4507,N_4444,N_4430);
nand U4508 (N_4508,N_4463,N_4497);
nor U4509 (N_4509,N_4422,N_4437);
nand U4510 (N_4510,N_4481,N_4493);
xnor U4511 (N_4511,N_4445,N_4466);
nand U4512 (N_4512,N_4417,N_4450);
xnor U4513 (N_4513,N_4428,N_4461);
nand U4514 (N_4514,N_4448,N_4494);
and U4515 (N_4515,N_4452,N_4484);
nor U4516 (N_4516,N_4457,N_4498);
and U4517 (N_4517,N_4479,N_4414);
xnor U4518 (N_4518,N_4467,N_4432);
nand U4519 (N_4519,N_4472,N_4447);
nor U4520 (N_4520,N_4455,N_4458);
nand U4521 (N_4521,N_4429,N_4480);
xnor U4522 (N_4522,N_4442,N_4411);
nor U4523 (N_4523,N_4473,N_4486);
nor U4524 (N_4524,N_4454,N_4434);
and U4525 (N_4525,N_4439,N_4418);
xor U4526 (N_4526,N_4406,N_4483);
nor U4527 (N_4527,N_4409,N_4460);
xor U4528 (N_4528,N_4496,N_4403);
xor U4529 (N_4529,N_4499,N_4420);
nor U4530 (N_4530,N_4456,N_4441);
nand U4531 (N_4531,N_4443,N_4425);
nand U4532 (N_4532,N_4475,N_4438);
xor U4533 (N_4533,N_4464,N_4476);
nand U4534 (N_4534,N_4412,N_4491);
or U4535 (N_4535,N_4440,N_4431);
and U4536 (N_4536,N_4449,N_4495);
nand U4537 (N_4537,N_4451,N_4402);
nor U4538 (N_4538,N_4482,N_4421);
and U4539 (N_4539,N_4427,N_4433);
nor U4540 (N_4540,N_4415,N_4492);
xor U4541 (N_4541,N_4485,N_4400);
or U4542 (N_4542,N_4468,N_4471);
nor U4543 (N_4543,N_4416,N_4459);
or U4544 (N_4544,N_4419,N_4408);
nor U4545 (N_4545,N_4446,N_4470);
nor U4546 (N_4546,N_4465,N_4407);
nor U4547 (N_4547,N_4490,N_4404);
nor U4548 (N_4548,N_4424,N_4462);
xnor U4549 (N_4549,N_4401,N_4413);
xor U4550 (N_4550,N_4425,N_4499);
xor U4551 (N_4551,N_4428,N_4475);
or U4552 (N_4552,N_4458,N_4448);
and U4553 (N_4553,N_4485,N_4473);
nand U4554 (N_4554,N_4475,N_4424);
or U4555 (N_4555,N_4403,N_4498);
nor U4556 (N_4556,N_4481,N_4448);
and U4557 (N_4557,N_4432,N_4457);
and U4558 (N_4558,N_4495,N_4428);
nand U4559 (N_4559,N_4404,N_4408);
xnor U4560 (N_4560,N_4486,N_4490);
nor U4561 (N_4561,N_4415,N_4439);
xnor U4562 (N_4562,N_4493,N_4421);
xnor U4563 (N_4563,N_4482,N_4445);
xor U4564 (N_4564,N_4402,N_4484);
or U4565 (N_4565,N_4406,N_4447);
xor U4566 (N_4566,N_4437,N_4412);
xnor U4567 (N_4567,N_4485,N_4484);
xnor U4568 (N_4568,N_4466,N_4426);
nand U4569 (N_4569,N_4451,N_4406);
nor U4570 (N_4570,N_4487,N_4461);
xnor U4571 (N_4571,N_4404,N_4467);
xor U4572 (N_4572,N_4498,N_4428);
or U4573 (N_4573,N_4423,N_4449);
or U4574 (N_4574,N_4417,N_4473);
nand U4575 (N_4575,N_4482,N_4402);
xor U4576 (N_4576,N_4482,N_4424);
nor U4577 (N_4577,N_4466,N_4402);
nand U4578 (N_4578,N_4499,N_4438);
nor U4579 (N_4579,N_4465,N_4468);
xor U4580 (N_4580,N_4401,N_4443);
xor U4581 (N_4581,N_4446,N_4460);
or U4582 (N_4582,N_4436,N_4400);
nor U4583 (N_4583,N_4456,N_4485);
nand U4584 (N_4584,N_4496,N_4444);
or U4585 (N_4585,N_4499,N_4440);
and U4586 (N_4586,N_4443,N_4470);
nor U4587 (N_4587,N_4465,N_4410);
and U4588 (N_4588,N_4409,N_4453);
nand U4589 (N_4589,N_4449,N_4483);
nand U4590 (N_4590,N_4467,N_4465);
nand U4591 (N_4591,N_4491,N_4464);
xor U4592 (N_4592,N_4443,N_4486);
or U4593 (N_4593,N_4408,N_4485);
xnor U4594 (N_4594,N_4466,N_4487);
nor U4595 (N_4595,N_4417,N_4433);
nor U4596 (N_4596,N_4474,N_4496);
nor U4597 (N_4597,N_4400,N_4462);
and U4598 (N_4598,N_4415,N_4471);
and U4599 (N_4599,N_4482,N_4438);
nor U4600 (N_4600,N_4585,N_4559);
xnor U4601 (N_4601,N_4535,N_4562);
and U4602 (N_4602,N_4555,N_4567);
nor U4603 (N_4603,N_4557,N_4542);
nand U4604 (N_4604,N_4524,N_4545);
xor U4605 (N_4605,N_4563,N_4552);
or U4606 (N_4606,N_4577,N_4515);
xor U4607 (N_4607,N_4532,N_4592);
xnor U4608 (N_4608,N_4588,N_4553);
or U4609 (N_4609,N_4572,N_4501);
nor U4610 (N_4610,N_4531,N_4514);
nor U4611 (N_4611,N_4580,N_4503);
nor U4612 (N_4612,N_4573,N_4546);
xor U4613 (N_4613,N_4596,N_4564);
and U4614 (N_4614,N_4508,N_4561);
and U4615 (N_4615,N_4587,N_4541);
xor U4616 (N_4616,N_4500,N_4569);
and U4617 (N_4617,N_4519,N_4551);
or U4618 (N_4618,N_4560,N_4583);
and U4619 (N_4619,N_4533,N_4518);
nor U4620 (N_4620,N_4591,N_4548);
and U4621 (N_4621,N_4554,N_4568);
or U4622 (N_4622,N_4538,N_4575);
xnor U4623 (N_4623,N_4547,N_4550);
and U4624 (N_4624,N_4565,N_4570);
or U4625 (N_4625,N_4534,N_4504);
nor U4626 (N_4626,N_4566,N_4543);
nor U4627 (N_4627,N_4544,N_4558);
nor U4628 (N_4628,N_4556,N_4597);
or U4629 (N_4629,N_4511,N_4513);
nor U4630 (N_4630,N_4516,N_4574);
nor U4631 (N_4631,N_4576,N_4578);
and U4632 (N_4632,N_4595,N_4594);
and U4633 (N_4633,N_4536,N_4598);
nand U4634 (N_4634,N_4507,N_4528);
nand U4635 (N_4635,N_4582,N_4510);
xnor U4636 (N_4636,N_4521,N_4527);
and U4637 (N_4637,N_4593,N_4581);
nand U4638 (N_4638,N_4539,N_4517);
and U4639 (N_4639,N_4505,N_4549);
nor U4640 (N_4640,N_4590,N_4530);
xor U4641 (N_4641,N_4525,N_4540);
and U4642 (N_4642,N_4512,N_4509);
and U4643 (N_4643,N_4522,N_4571);
xnor U4644 (N_4644,N_4537,N_4506);
and U4645 (N_4645,N_4586,N_4589);
nand U4646 (N_4646,N_4584,N_4529);
or U4647 (N_4647,N_4599,N_4502);
and U4648 (N_4648,N_4520,N_4579);
xor U4649 (N_4649,N_4526,N_4523);
nor U4650 (N_4650,N_4542,N_4527);
or U4651 (N_4651,N_4568,N_4557);
nand U4652 (N_4652,N_4573,N_4506);
or U4653 (N_4653,N_4588,N_4508);
or U4654 (N_4654,N_4559,N_4523);
nor U4655 (N_4655,N_4520,N_4545);
and U4656 (N_4656,N_4523,N_4582);
or U4657 (N_4657,N_4520,N_4539);
xnor U4658 (N_4658,N_4568,N_4595);
nor U4659 (N_4659,N_4561,N_4578);
xnor U4660 (N_4660,N_4570,N_4594);
or U4661 (N_4661,N_4538,N_4555);
nand U4662 (N_4662,N_4560,N_4575);
and U4663 (N_4663,N_4523,N_4583);
xnor U4664 (N_4664,N_4592,N_4584);
and U4665 (N_4665,N_4535,N_4509);
and U4666 (N_4666,N_4530,N_4569);
nor U4667 (N_4667,N_4559,N_4543);
nand U4668 (N_4668,N_4593,N_4513);
and U4669 (N_4669,N_4525,N_4595);
and U4670 (N_4670,N_4515,N_4580);
nand U4671 (N_4671,N_4576,N_4551);
xnor U4672 (N_4672,N_4593,N_4516);
nand U4673 (N_4673,N_4552,N_4590);
and U4674 (N_4674,N_4552,N_4594);
nor U4675 (N_4675,N_4592,N_4597);
nor U4676 (N_4676,N_4513,N_4509);
nand U4677 (N_4677,N_4555,N_4588);
xor U4678 (N_4678,N_4533,N_4543);
and U4679 (N_4679,N_4541,N_4524);
and U4680 (N_4680,N_4517,N_4548);
and U4681 (N_4681,N_4532,N_4572);
and U4682 (N_4682,N_4591,N_4599);
and U4683 (N_4683,N_4540,N_4510);
and U4684 (N_4684,N_4579,N_4557);
or U4685 (N_4685,N_4519,N_4567);
nor U4686 (N_4686,N_4540,N_4587);
nor U4687 (N_4687,N_4533,N_4575);
and U4688 (N_4688,N_4520,N_4581);
xor U4689 (N_4689,N_4597,N_4542);
and U4690 (N_4690,N_4532,N_4598);
or U4691 (N_4691,N_4580,N_4595);
nand U4692 (N_4692,N_4500,N_4564);
and U4693 (N_4693,N_4553,N_4516);
nand U4694 (N_4694,N_4562,N_4565);
xor U4695 (N_4695,N_4576,N_4567);
nor U4696 (N_4696,N_4584,N_4547);
nand U4697 (N_4697,N_4538,N_4520);
xor U4698 (N_4698,N_4584,N_4515);
nor U4699 (N_4699,N_4572,N_4521);
nor U4700 (N_4700,N_4641,N_4610);
nand U4701 (N_4701,N_4653,N_4600);
and U4702 (N_4702,N_4646,N_4695);
nand U4703 (N_4703,N_4636,N_4661);
nand U4704 (N_4704,N_4656,N_4671);
xnor U4705 (N_4705,N_4662,N_4659);
nand U4706 (N_4706,N_4611,N_4660);
nor U4707 (N_4707,N_4657,N_4678);
nor U4708 (N_4708,N_4687,N_4670);
nand U4709 (N_4709,N_4673,N_4621);
xnor U4710 (N_4710,N_4626,N_4627);
and U4711 (N_4711,N_4633,N_4614);
xnor U4712 (N_4712,N_4651,N_4680);
nor U4713 (N_4713,N_4652,N_4639);
nor U4714 (N_4714,N_4619,N_4612);
nand U4715 (N_4715,N_4604,N_4649);
nand U4716 (N_4716,N_4689,N_4609);
xnor U4717 (N_4717,N_4686,N_4668);
xor U4718 (N_4718,N_4632,N_4683);
and U4719 (N_4719,N_4630,N_4643);
xor U4720 (N_4720,N_4628,N_4629);
or U4721 (N_4721,N_4665,N_4675);
nand U4722 (N_4722,N_4688,N_4637);
and U4723 (N_4723,N_4624,N_4605);
nor U4724 (N_4724,N_4658,N_4677);
or U4725 (N_4725,N_4622,N_4645);
xor U4726 (N_4726,N_4634,N_4664);
nor U4727 (N_4727,N_4691,N_4638);
xnor U4728 (N_4728,N_4607,N_4617);
nand U4729 (N_4729,N_4603,N_4699);
or U4730 (N_4730,N_4631,N_4679);
and U4731 (N_4731,N_4696,N_4642);
nor U4732 (N_4732,N_4601,N_4644);
nand U4733 (N_4733,N_4625,N_4674);
xnor U4734 (N_4734,N_4602,N_4681);
xnor U4735 (N_4735,N_4615,N_4672);
nand U4736 (N_4736,N_4684,N_4613);
and U4737 (N_4737,N_4694,N_4667);
nor U4738 (N_4738,N_4640,N_4697);
and U4739 (N_4739,N_4693,N_4616);
xor U4740 (N_4740,N_4650,N_4655);
nor U4741 (N_4741,N_4654,N_4685);
or U4742 (N_4742,N_4682,N_4690);
xor U4743 (N_4743,N_4676,N_4606);
or U4744 (N_4744,N_4663,N_4648);
and U4745 (N_4745,N_4647,N_4666);
or U4746 (N_4746,N_4635,N_4623);
xor U4747 (N_4747,N_4618,N_4692);
nor U4748 (N_4748,N_4608,N_4669);
nor U4749 (N_4749,N_4698,N_4620);
xnor U4750 (N_4750,N_4689,N_4688);
and U4751 (N_4751,N_4690,N_4656);
or U4752 (N_4752,N_4643,N_4621);
and U4753 (N_4753,N_4652,N_4615);
or U4754 (N_4754,N_4674,N_4648);
nand U4755 (N_4755,N_4647,N_4675);
nand U4756 (N_4756,N_4692,N_4634);
and U4757 (N_4757,N_4639,N_4620);
xnor U4758 (N_4758,N_4682,N_4612);
nand U4759 (N_4759,N_4674,N_4685);
nand U4760 (N_4760,N_4621,N_4609);
nand U4761 (N_4761,N_4619,N_4693);
nand U4762 (N_4762,N_4692,N_4667);
and U4763 (N_4763,N_4619,N_4641);
and U4764 (N_4764,N_4696,N_4670);
and U4765 (N_4765,N_4667,N_4638);
nand U4766 (N_4766,N_4694,N_4683);
and U4767 (N_4767,N_4643,N_4667);
and U4768 (N_4768,N_4629,N_4676);
and U4769 (N_4769,N_4694,N_4626);
or U4770 (N_4770,N_4615,N_4608);
nand U4771 (N_4771,N_4619,N_4668);
xor U4772 (N_4772,N_4601,N_4647);
nor U4773 (N_4773,N_4618,N_4666);
nor U4774 (N_4774,N_4673,N_4640);
nand U4775 (N_4775,N_4676,N_4609);
xnor U4776 (N_4776,N_4699,N_4601);
and U4777 (N_4777,N_4659,N_4620);
nand U4778 (N_4778,N_4620,N_4615);
xnor U4779 (N_4779,N_4653,N_4664);
and U4780 (N_4780,N_4616,N_4620);
nand U4781 (N_4781,N_4670,N_4681);
nor U4782 (N_4782,N_4684,N_4672);
nor U4783 (N_4783,N_4663,N_4639);
or U4784 (N_4784,N_4625,N_4637);
and U4785 (N_4785,N_4649,N_4647);
xnor U4786 (N_4786,N_4614,N_4678);
and U4787 (N_4787,N_4697,N_4681);
xor U4788 (N_4788,N_4693,N_4629);
xnor U4789 (N_4789,N_4621,N_4615);
and U4790 (N_4790,N_4630,N_4612);
or U4791 (N_4791,N_4650,N_4682);
or U4792 (N_4792,N_4617,N_4600);
and U4793 (N_4793,N_4642,N_4674);
xor U4794 (N_4794,N_4675,N_4679);
or U4795 (N_4795,N_4696,N_4690);
nor U4796 (N_4796,N_4617,N_4671);
and U4797 (N_4797,N_4634,N_4655);
nand U4798 (N_4798,N_4610,N_4682);
and U4799 (N_4799,N_4687,N_4652);
and U4800 (N_4800,N_4758,N_4701);
or U4801 (N_4801,N_4763,N_4743);
or U4802 (N_4802,N_4742,N_4767);
nor U4803 (N_4803,N_4707,N_4728);
nor U4804 (N_4804,N_4761,N_4791);
nand U4805 (N_4805,N_4721,N_4770);
or U4806 (N_4806,N_4760,N_4797);
nor U4807 (N_4807,N_4712,N_4768);
xor U4808 (N_4808,N_4739,N_4792);
or U4809 (N_4809,N_4772,N_4740);
and U4810 (N_4810,N_4724,N_4723);
or U4811 (N_4811,N_4700,N_4780);
or U4812 (N_4812,N_4789,N_4717);
and U4813 (N_4813,N_4727,N_4720);
nor U4814 (N_4814,N_4746,N_4798);
and U4815 (N_4815,N_4719,N_4702);
and U4816 (N_4816,N_4783,N_4790);
and U4817 (N_4817,N_4710,N_4730);
nor U4818 (N_4818,N_4750,N_4796);
and U4819 (N_4819,N_4786,N_4753);
nor U4820 (N_4820,N_4714,N_4765);
xnor U4821 (N_4821,N_4713,N_4747);
nor U4822 (N_4822,N_4788,N_4734);
nand U4823 (N_4823,N_4776,N_4775);
and U4824 (N_4824,N_4781,N_4784);
or U4825 (N_4825,N_4715,N_4745);
xnor U4826 (N_4826,N_4762,N_4722);
xnor U4827 (N_4827,N_4754,N_4779);
and U4828 (N_4828,N_4774,N_4733);
or U4829 (N_4829,N_4771,N_4757);
nand U4830 (N_4830,N_4737,N_4773);
xor U4831 (N_4831,N_4705,N_4759);
nor U4832 (N_4832,N_4729,N_4778);
nor U4833 (N_4833,N_4764,N_4785);
or U4834 (N_4834,N_4795,N_4755);
nand U4835 (N_4835,N_4794,N_4703);
nor U4836 (N_4836,N_4738,N_4748);
nor U4837 (N_4837,N_4766,N_4752);
nand U4838 (N_4838,N_4732,N_4741);
or U4839 (N_4839,N_4777,N_4708);
nand U4840 (N_4840,N_4782,N_4718);
nand U4841 (N_4841,N_4725,N_4709);
and U4842 (N_4842,N_4711,N_4736);
or U4843 (N_4843,N_4716,N_4706);
nand U4844 (N_4844,N_4799,N_4731);
nor U4845 (N_4845,N_4744,N_4749);
and U4846 (N_4846,N_4726,N_4793);
nand U4847 (N_4847,N_4704,N_4735);
or U4848 (N_4848,N_4756,N_4769);
or U4849 (N_4849,N_4787,N_4751);
or U4850 (N_4850,N_4762,N_4774);
nor U4851 (N_4851,N_4771,N_4725);
and U4852 (N_4852,N_4708,N_4747);
nor U4853 (N_4853,N_4783,N_4742);
and U4854 (N_4854,N_4753,N_4775);
xor U4855 (N_4855,N_4792,N_4756);
or U4856 (N_4856,N_4744,N_4706);
nor U4857 (N_4857,N_4754,N_4718);
nand U4858 (N_4858,N_4747,N_4779);
or U4859 (N_4859,N_4705,N_4746);
nor U4860 (N_4860,N_4773,N_4772);
and U4861 (N_4861,N_4752,N_4796);
nand U4862 (N_4862,N_4700,N_4797);
or U4863 (N_4863,N_4788,N_4756);
xnor U4864 (N_4864,N_4754,N_4794);
nor U4865 (N_4865,N_4770,N_4752);
or U4866 (N_4866,N_4745,N_4742);
and U4867 (N_4867,N_4788,N_4740);
or U4868 (N_4868,N_4778,N_4775);
and U4869 (N_4869,N_4774,N_4738);
and U4870 (N_4870,N_4758,N_4745);
nor U4871 (N_4871,N_4765,N_4719);
nand U4872 (N_4872,N_4790,N_4753);
xnor U4873 (N_4873,N_4727,N_4763);
nand U4874 (N_4874,N_4739,N_4745);
and U4875 (N_4875,N_4710,N_4796);
or U4876 (N_4876,N_4728,N_4788);
nand U4877 (N_4877,N_4731,N_4715);
nor U4878 (N_4878,N_4757,N_4768);
xor U4879 (N_4879,N_4718,N_4715);
nor U4880 (N_4880,N_4781,N_4739);
nor U4881 (N_4881,N_4758,N_4715);
xor U4882 (N_4882,N_4700,N_4776);
nor U4883 (N_4883,N_4742,N_4702);
xor U4884 (N_4884,N_4721,N_4784);
nor U4885 (N_4885,N_4759,N_4707);
nor U4886 (N_4886,N_4769,N_4752);
nor U4887 (N_4887,N_4731,N_4764);
or U4888 (N_4888,N_4705,N_4725);
or U4889 (N_4889,N_4745,N_4751);
xor U4890 (N_4890,N_4763,N_4715);
nand U4891 (N_4891,N_4772,N_4792);
and U4892 (N_4892,N_4744,N_4797);
or U4893 (N_4893,N_4779,N_4700);
or U4894 (N_4894,N_4711,N_4715);
nand U4895 (N_4895,N_4782,N_4726);
nor U4896 (N_4896,N_4722,N_4720);
and U4897 (N_4897,N_4748,N_4721);
or U4898 (N_4898,N_4740,N_4731);
and U4899 (N_4899,N_4797,N_4747);
or U4900 (N_4900,N_4888,N_4830);
nor U4901 (N_4901,N_4841,N_4881);
or U4902 (N_4902,N_4880,N_4860);
nor U4903 (N_4903,N_4826,N_4805);
xor U4904 (N_4904,N_4889,N_4853);
xor U4905 (N_4905,N_4802,N_4856);
xnor U4906 (N_4906,N_4834,N_4819);
or U4907 (N_4907,N_4811,N_4894);
nor U4908 (N_4908,N_4837,N_4831);
and U4909 (N_4909,N_4852,N_4833);
and U4910 (N_4910,N_4896,N_4846);
and U4911 (N_4911,N_4818,N_4840);
xnor U4912 (N_4912,N_4800,N_4828);
or U4913 (N_4913,N_4870,N_4832);
or U4914 (N_4914,N_4887,N_4882);
nand U4915 (N_4915,N_4845,N_4847);
xnor U4916 (N_4916,N_4807,N_4886);
xor U4917 (N_4917,N_4810,N_4850);
or U4918 (N_4918,N_4806,N_4835);
xor U4919 (N_4919,N_4890,N_4849);
nand U4920 (N_4920,N_4895,N_4893);
or U4921 (N_4921,N_4864,N_4885);
and U4922 (N_4922,N_4876,N_4865);
nand U4923 (N_4923,N_4843,N_4822);
or U4924 (N_4924,N_4804,N_4812);
or U4925 (N_4925,N_4883,N_4862);
nor U4926 (N_4926,N_4855,N_4874);
or U4927 (N_4927,N_4857,N_4884);
xnor U4928 (N_4928,N_4866,N_4813);
or U4929 (N_4929,N_4801,N_4838);
nor U4930 (N_4930,N_4877,N_4829);
nor U4931 (N_4931,N_4809,N_4827);
xnor U4932 (N_4932,N_4858,N_4899);
nor U4933 (N_4933,N_4823,N_4898);
and U4934 (N_4934,N_4839,N_4825);
xor U4935 (N_4935,N_4821,N_4875);
nand U4936 (N_4936,N_4872,N_4861);
xor U4937 (N_4937,N_4863,N_4816);
nor U4938 (N_4938,N_4867,N_4868);
nor U4939 (N_4939,N_4854,N_4844);
xnor U4940 (N_4940,N_4808,N_4873);
nand U4941 (N_4941,N_4836,N_4803);
nand U4942 (N_4942,N_4891,N_4842);
nor U4943 (N_4943,N_4815,N_4871);
or U4944 (N_4944,N_4859,N_4869);
xnor U4945 (N_4945,N_4824,N_4851);
and U4946 (N_4946,N_4878,N_4848);
and U4947 (N_4947,N_4892,N_4814);
nor U4948 (N_4948,N_4897,N_4879);
xnor U4949 (N_4949,N_4820,N_4817);
or U4950 (N_4950,N_4853,N_4860);
xor U4951 (N_4951,N_4895,N_4863);
nand U4952 (N_4952,N_4899,N_4842);
xor U4953 (N_4953,N_4819,N_4810);
and U4954 (N_4954,N_4837,N_4836);
nand U4955 (N_4955,N_4804,N_4860);
and U4956 (N_4956,N_4843,N_4816);
nand U4957 (N_4957,N_4848,N_4872);
and U4958 (N_4958,N_4805,N_4870);
and U4959 (N_4959,N_4827,N_4857);
and U4960 (N_4960,N_4814,N_4856);
xnor U4961 (N_4961,N_4820,N_4891);
nand U4962 (N_4962,N_4830,N_4849);
and U4963 (N_4963,N_4874,N_4830);
and U4964 (N_4964,N_4847,N_4801);
xor U4965 (N_4965,N_4835,N_4801);
nand U4966 (N_4966,N_4872,N_4880);
or U4967 (N_4967,N_4879,N_4810);
nand U4968 (N_4968,N_4896,N_4816);
xor U4969 (N_4969,N_4872,N_4877);
nand U4970 (N_4970,N_4800,N_4827);
and U4971 (N_4971,N_4868,N_4815);
or U4972 (N_4972,N_4867,N_4807);
xnor U4973 (N_4973,N_4809,N_4858);
xnor U4974 (N_4974,N_4805,N_4812);
xor U4975 (N_4975,N_4812,N_4800);
or U4976 (N_4976,N_4885,N_4888);
xnor U4977 (N_4977,N_4894,N_4821);
nand U4978 (N_4978,N_4890,N_4822);
nor U4979 (N_4979,N_4809,N_4886);
or U4980 (N_4980,N_4865,N_4850);
or U4981 (N_4981,N_4847,N_4815);
nand U4982 (N_4982,N_4815,N_4897);
nor U4983 (N_4983,N_4806,N_4897);
nand U4984 (N_4984,N_4854,N_4866);
and U4985 (N_4985,N_4806,N_4847);
or U4986 (N_4986,N_4850,N_4802);
or U4987 (N_4987,N_4869,N_4843);
and U4988 (N_4988,N_4854,N_4800);
nand U4989 (N_4989,N_4891,N_4808);
xor U4990 (N_4990,N_4836,N_4857);
nand U4991 (N_4991,N_4853,N_4871);
nand U4992 (N_4992,N_4845,N_4870);
nand U4993 (N_4993,N_4881,N_4896);
xor U4994 (N_4994,N_4865,N_4836);
and U4995 (N_4995,N_4802,N_4846);
and U4996 (N_4996,N_4890,N_4854);
and U4997 (N_4997,N_4875,N_4893);
nand U4998 (N_4998,N_4848,N_4840);
nand U4999 (N_4999,N_4870,N_4868);
or UO_0 (O_0,N_4963,N_4925);
xor UO_1 (O_1,N_4979,N_4975);
nand UO_2 (O_2,N_4910,N_4926);
nor UO_3 (O_3,N_4957,N_4944);
nor UO_4 (O_4,N_4901,N_4972);
xor UO_5 (O_5,N_4968,N_4900);
or UO_6 (O_6,N_4948,N_4919);
xor UO_7 (O_7,N_4971,N_4933);
xor UO_8 (O_8,N_4916,N_4902);
nand UO_9 (O_9,N_4946,N_4922);
and UO_10 (O_10,N_4929,N_4997);
nand UO_11 (O_11,N_4907,N_4905);
and UO_12 (O_12,N_4993,N_4962);
and UO_13 (O_13,N_4986,N_4985);
nor UO_14 (O_14,N_4953,N_4969);
or UO_15 (O_15,N_4956,N_4999);
nand UO_16 (O_16,N_4937,N_4915);
or UO_17 (O_17,N_4981,N_4918);
nor UO_18 (O_18,N_4960,N_4932);
or UO_19 (O_19,N_4994,N_4941);
or UO_20 (O_20,N_4920,N_4978);
or UO_21 (O_21,N_4906,N_4992);
or UO_22 (O_22,N_4936,N_4908);
or UO_23 (O_23,N_4996,N_4909);
xor UO_24 (O_24,N_4943,N_4984);
xor UO_25 (O_25,N_4983,N_4942);
nor UO_26 (O_26,N_4961,N_4923);
xor UO_27 (O_27,N_4967,N_4955);
nor UO_28 (O_28,N_4970,N_4940);
nor UO_29 (O_29,N_4982,N_4974);
and UO_30 (O_30,N_4917,N_4949);
xnor UO_31 (O_31,N_4966,N_4976);
or UO_32 (O_32,N_4995,N_4980);
and UO_33 (O_33,N_4931,N_4991);
xor UO_34 (O_34,N_4938,N_4945);
and UO_35 (O_35,N_4930,N_4947);
and UO_36 (O_36,N_4973,N_4988);
xnor UO_37 (O_37,N_4987,N_4952);
or UO_38 (O_38,N_4911,N_4913);
and UO_39 (O_39,N_4935,N_4965);
or UO_40 (O_40,N_4964,N_4921);
and UO_41 (O_41,N_4912,N_4934);
nor UO_42 (O_42,N_4924,N_4950);
xnor UO_43 (O_43,N_4998,N_4954);
and UO_44 (O_44,N_4990,N_4989);
nor UO_45 (O_45,N_4914,N_4927);
and UO_46 (O_46,N_4959,N_4951);
xor UO_47 (O_47,N_4977,N_4939);
nor UO_48 (O_48,N_4904,N_4903);
and UO_49 (O_49,N_4958,N_4928);
nand UO_50 (O_50,N_4987,N_4944);
nand UO_51 (O_51,N_4906,N_4974);
nor UO_52 (O_52,N_4957,N_4931);
nor UO_53 (O_53,N_4986,N_4919);
nor UO_54 (O_54,N_4990,N_4930);
nand UO_55 (O_55,N_4930,N_4924);
nand UO_56 (O_56,N_4900,N_4919);
or UO_57 (O_57,N_4917,N_4946);
and UO_58 (O_58,N_4934,N_4916);
xnor UO_59 (O_59,N_4984,N_4990);
xnor UO_60 (O_60,N_4950,N_4943);
xnor UO_61 (O_61,N_4903,N_4939);
xnor UO_62 (O_62,N_4980,N_4908);
or UO_63 (O_63,N_4980,N_4978);
or UO_64 (O_64,N_4938,N_4988);
nand UO_65 (O_65,N_4906,N_4958);
or UO_66 (O_66,N_4936,N_4972);
nor UO_67 (O_67,N_4991,N_4975);
or UO_68 (O_68,N_4997,N_4970);
and UO_69 (O_69,N_4904,N_4934);
nand UO_70 (O_70,N_4980,N_4981);
nor UO_71 (O_71,N_4947,N_4979);
and UO_72 (O_72,N_4973,N_4915);
or UO_73 (O_73,N_4983,N_4925);
nor UO_74 (O_74,N_4992,N_4981);
nor UO_75 (O_75,N_4905,N_4923);
nor UO_76 (O_76,N_4900,N_4986);
xor UO_77 (O_77,N_4939,N_4991);
and UO_78 (O_78,N_4961,N_4941);
nor UO_79 (O_79,N_4907,N_4977);
or UO_80 (O_80,N_4986,N_4944);
or UO_81 (O_81,N_4949,N_4945);
nand UO_82 (O_82,N_4961,N_4927);
and UO_83 (O_83,N_4900,N_4947);
or UO_84 (O_84,N_4990,N_4945);
and UO_85 (O_85,N_4912,N_4977);
xor UO_86 (O_86,N_4967,N_4998);
and UO_87 (O_87,N_4957,N_4932);
xor UO_88 (O_88,N_4984,N_4955);
xnor UO_89 (O_89,N_4946,N_4918);
xor UO_90 (O_90,N_4942,N_4939);
nor UO_91 (O_91,N_4996,N_4907);
or UO_92 (O_92,N_4978,N_4915);
nor UO_93 (O_93,N_4965,N_4971);
nor UO_94 (O_94,N_4901,N_4976);
nand UO_95 (O_95,N_4918,N_4949);
xor UO_96 (O_96,N_4992,N_4978);
nor UO_97 (O_97,N_4947,N_4964);
and UO_98 (O_98,N_4930,N_4996);
nor UO_99 (O_99,N_4938,N_4968);
and UO_100 (O_100,N_4908,N_4967);
and UO_101 (O_101,N_4940,N_4912);
nand UO_102 (O_102,N_4953,N_4947);
nor UO_103 (O_103,N_4921,N_4992);
or UO_104 (O_104,N_4960,N_4968);
nand UO_105 (O_105,N_4972,N_4963);
nor UO_106 (O_106,N_4940,N_4954);
xor UO_107 (O_107,N_4924,N_4971);
or UO_108 (O_108,N_4966,N_4943);
nor UO_109 (O_109,N_4937,N_4924);
and UO_110 (O_110,N_4943,N_4915);
and UO_111 (O_111,N_4935,N_4944);
xnor UO_112 (O_112,N_4951,N_4917);
nor UO_113 (O_113,N_4939,N_4911);
xor UO_114 (O_114,N_4984,N_4923);
xnor UO_115 (O_115,N_4984,N_4989);
or UO_116 (O_116,N_4945,N_4911);
nor UO_117 (O_117,N_4980,N_4900);
nor UO_118 (O_118,N_4941,N_4901);
or UO_119 (O_119,N_4990,N_4906);
or UO_120 (O_120,N_4912,N_4948);
and UO_121 (O_121,N_4976,N_4917);
xor UO_122 (O_122,N_4900,N_4954);
nor UO_123 (O_123,N_4907,N_4934);
or UO_124 (O_124,N_4994,N_4923);
or UO_125 (O_125,N_4922,N_4967);
and UO_126 (O_126,N_4938,N_4924);
or UO_127 (O_127,N_4909,N_4949);
and UO_128 (O_128,N_4998,N_4950);
or UO_129 (O_129,N_4974,N_4934);
or UO_130 (O_130,N_4997,N_4954);
nand UO_131 (O_131,N_4981,N_4970);
or UO_132 (O_132,N_4906,N_4946);
nand UO_133 (O_133,N_4918,N_4968);
nor UO_134 (O_134,N_4982,N_4931);
xnor UO_135 (O_135,N_4923,N_4922);
nor UO_136 (O_136,N_4946,N_4979);
or UO_137 (O_137,N_4999,N_4957);
xor UO_138 (O_138,N_4900,N_4982);
xor UO_139 (O_139,N_4984,N_4968);
nand UO_140 (O_140,N_4990,N_4947);
xor UO_141 (O_141,N_4938,N_4970);
nor UO_142 (O_142,N_4940,N_4918);
or UO_143 (O_143,N_4904,N_4912);
nand UO_144 (O_144,N_4982,N_4976);
and UO_145 (O_145,N_4922,N_4953);
xor UO_146 (O_146,N_4970,N_4952);
nor UO_147 (O_147,N_4984,N_4927);
and UO_148 (O_148,N_4914,N_4981);
and UO_149 (O_149,N_4985,N_4987);
nand UO_150 (O_150,N_4984,N_4946);
nand UO_151 (O_151,N_4936,N_4938);
or UO_152 (O_152,N_4999,N_4909);
nor UO_153 (O_153,N_4994,N_4938);
xnor UO_154 (O_154,N_4917,N_4929);
nor UO_155 (O_155,N_4991,N_4914);
nor UO_156 (O_156,N_4943,N_4977);
nor UO_157 (O_157,N_4960,N_4955);
nand UO_158 (O_158,N_4976,N_4977);
xnor UO_159 (O_159,N_4969,N_4911);
xnor UO_160 (O_160,N_4913,N_4910);
or UO_161 (O_161,N_4947,N_4941);
xnor UO_162 (O_162,N_4931,N_4932);
xnor UO_163 (O_163,N_4938,N_4984);
and UO_164 (O_164,N_4904,N_4933);
xnor UO_165 (O_165,N_4993,N_4932);
nand UO_166 (O_166,N_4940,N_4962);
nand UO_167 (O_167,N_4958,N_4949);
and UO_168 (O_168,N_4942,N_4934);
nor UO_169 (O_169,N_4989,N_4934);
or UO_170 (O_170,N_4983,N_4917);
nor UO_171 (O_171,N_4952,N_4918);
or UO_172 (O_172,N_4961,N_4968);
or UO_173 (O_173,N_4973,N_4999);
or UO_174 (O_174,N_4914,N_4992);
nand UO_175 (O_175,N_4934,N_4957);
xnor UO_176 (O_176,N_4965,N_4961);
nor UO_177 (O_177,N_4966,N_4995);
or UO_178 (O_178,N_4918,N_4972);
or UO_179 (O_179,N_4970,N_4954);
and UO_180 (O_180,N_4905,N_4903);
nor UO_181 (O_181,N_4976,N_4967);
xnor UO_182 (O_182,N_4943,N_4906);
xnor UO_183 (O_183,N_4994,N_4986);
and UO_184 (O_184,N_4911,N_4964);
nor UO_185 (O_185,N_4909,N_4901);
xor UO_186 (O_186,N_4929,N_4975);
nor UO_187 (O_187,N_4953,N_4934);
nor UO_188 (O_188,N_4901,N_4989);
or UO_189 (O_189,N_4990,N_4959);
and UO_190 (O_190,N_4975,N_4941);
or UO_191 (O_191,N_4903,N_4900);
xor UO_192 (O_192,N_4968,N_4989);
nor UO_193 (O_193,N_4983,N_4921);
xor UO_194 (O_194,N_4901,N_4902);
and UO_195 (O_195,N_4900,N_4952);
nand UO_196 (O_196,N_4991,N_4974);
and UO_197 (O_197,N_4959,N_4919);
or UO_198 (O_198,N_4933,N_4925);
xor UO_199 (O_199,N_4976,N_4954);
and UO_200 (O_200,N_4979,N_4993);
and UO_201 (O_201,N_4921,N_4931);
and UO_202 (O_202,N_4948,N_4970);
nand UO_203 (O_203,N_4913,N_4970);
xor UO_204 (O_204,N_4997,N_4916);
nand UO_205 (O_205,N_4935,N_4940);
and UO_206 (O_206,N_4959,N_4991);
nor UO_207 (O_207,N_4950,N_4908);
or UO_208 (O_208,N_4967,N_4905);
or UO_209 (O_209,N_4971,N_4934);
nor UO_210 (O_210,N_4918,N_4998);
xnor UO_211 (O_211,N_4913,N_4946);
nand UO_212 (O_212,N_4996,N_4932);
nand UO_213 (O_213,N_4965,N_4921);
nand UO_214 (O_214,N_4900,N_4936);
nand UO_215 (O_215,N_4992,N_4982);
xor UO_216 (O_216,N_4950,N_4956);
nand UO_217 (O_217,N_4943,N_4911);
or UO_218 (O_218,N_4956,N_4935);
xor UO_219 (O_219,N_4982,N_4927);
nor UO_220 (O_220,N_4920,N_4926);
nor UO_221 (O_221,N_4903,N_4920);
nand UO_222 (O_222,N_4980,N_4929);
or UO_223 (O_223,N_4925,N_4996);
nor UO_224 (O_224,N_4973,N_4971);
nand UO_225 (O_225,N_4907,N_4954);
nor UO_226 (O_226,N_4995,N_4978);
nor UO_227 (O_227,N_4997,N_4906);
nand UO_228 (O_228,N_4991,N_4993);
nand UO_229 (O_229,N_4985,N_4950);
nor UO_230 (O_230,N_4952,N_4988);
nand UO_231 (O_231,N_4960,N_4926);
or UO_232 (O_232,N_4943,N_4916);
and UO_233 (O_233,N_4905,N_4904);
nand UO_234 (O_234,N_4928,N_4932);
xnor UO_235 (O_235,N_4930,N_4955);
nor UO_236 (O_236,N_4935,N_4987);
and UO_237 (O_237,N_4901,N_4981);
xor UO_238 (O_238,N_4971,N_4993);
nor UO_239 (O_239,N_4986,N_4968);
and UO_240 (O_240,N_4920,N_4907);
and UO_241 (O_241,N_4962,N_4942);
or UO_242 (O_242,N_4928,N_4934);
and UO_243 (O_243,N_4941,N_4938);
and UO_244 (O_244,N_4954,N_4932);
and UO_245 (O_245,N_4986,N_4972);
nor UO_246 (O_246,N_4952,N_4966);
nand UO_247 (O_247,N_4993,N_4955);
nor UO_248 (O_248,N_4934,N_4925);
xnor UO_249 (O_249,N_4925,N_4952);
or UO_250 (O_250,N_4992,N_4913);
or UO_251 (O_251,N_4922,N_4949);
or UO_252 (O_252,N_4954,N_4981);
nor UO_253 (O_253,N_4998,N_4944);
nor UO_254 (O_254,N_4907,N_4975);
xnor UO_255 (O_255,N_4957,N_4913);
nor UO_256 (O_256,N_4906,N_4918);
xnor UO_257 (O_257,N_4919,N_4930);
xor UO_258 (O_258,N_4933,N_4915);
nand UO_259 (O_259,N_4911,N_4938);
nand UO_260 (O_260,N_4905,N_4968);
and UO_261 (O_261,N_4911,N_4984);
or UO_262 (O_262,N_4961,N_4910);
nor UO_263 (O_263,N_4976,N_4918);
or UO_264 (O_264,N_4926,N_4930);
or UO_265 (O_265,N_4938,N_4959);
or UO_266 (O_266,N_4919,N_4979);
xnor UO_267 (O_267,N_4924,N_4928);
nor UO_268 (O_268,N_4916,N_4948);
nor UO_269 (O_269,N_4906,N_4962);
nor UO_270 (O_270,N_4959,N_4929);
or UO_271 (O_271,N_4995,N_4901);
nand UO_272 (O_272,N_4951,N_4941);
nor UO_273 (O_273,N_4929,N_4984);
nor UO_274 (O_274,N_4981,N_4969);
nand UO_275 (O_275,N_4996,N_4973);
and UO_276 (O_276,N_4908,N_4957);
nor UO_277 (O_277,N_4941,N_4904);
and UO_278 (O_278,N_4943,N_4976);
or UO_279 (O_279,N_4978,N_4902);
nor UO_280 (O_280,N_4920,N_4996);
nand UO_281 (O_281,N_4965,N_4925);
nor UO_282 (O_282,N_4928,N_4972);
nor UO_283 (O_283,N_4918,N_4987);
xnor UO_284 (O_284,N_4967,N_4965);
or UO_285 (O_285,N_4997,N_4919);
xor UO_286 (O_286,N_4936,N_4907);
and UO_287 (O_287,N_4925,N_4917);
nor UO_288 (O_288,N_4972,N_4994);
and UO_289 (O_289,N_4940,N_4972);
nand UO_290 (O_290,N_4918,N_4994);
xnor UO_291 (O_291,N_4963,N_4994);
xor UO_292 (O_292,N_4986,N_4973);
nor UO_293 (O_293,N_4937,N_4996);
and UO_294 (O_294,N_4943,N_4931);
and UO_295 (O_295,N_4970,N_4960);
xnor UO_296 (O_296,N_4989,N_4900);
nand UO_297 (O_297,N_4967,N_4979);
nor UO_298 (O_298,N_4976,N_4933);
and UO_299 (O_299,N_4905,N_4978);
and UO_300 (O_300,N_4977,N_4930);
nor UO_301 (O_301,N_4933,N_4962);
nand UO_302 (O_302,N_4993,N_4966);
nor UO_303 (O_303,N_4944,N_4955);
nand UO_304 (O_304,N_4981,N_4962);
xnor UO_305 (O_305,N_4951,N_4956);
nand UO_306 (O_306,N_4948,N_4987);
xnor UO_307 (O_307,N_4979,N_4931);
nor UO_308 (O_308,N_4964,N_4994);
and UO_309 (O_309,N_4927,N_4995);
nor UO_310 (O_310,N_4974,N_4966);
xor UO_311 (O_311,N_4935,N_4967);
nor UO_312 (O_312,N_4983,N_4944);
nor UO_313 (O_313,N_4963,N_4965);
or UO_314 (O_314,N_4942,N_4955);
and UO_315 (O_315,N_4957,N_4922);
nand UO_316 (O_316,N_4948,N_4930);
or UO_317 (O_317,N_4941,N_4942);
nand UO_318 (O_318,N_4911,N_4994);
nand UO_319 (O_319,N_4986,N_4961);
nand UO_320 (O_320,N_4918,N_4932);
or UO_321 (O_321,N_4964,N_4903);
nand UO_322 (O_322,N_4925,N_4987);
nor UO_323 (O_323,N_4991,N_4902);
xnor UO_324 (O_324,N_4982,N_4930);
nor UO_325 (O_325,N_4985,N_4930);
nor UO_326 (O_326,N_4945,N_4953);
xnor UO_327 (O_327,N_4934,N_4983);
nand UO_328 (O_328,N_4998,N_4942);
xor UO_329 (O_329,N_4967,N_4910);
xnor UO_330 (O_330,N_4908,N_4917);
xor UO_331 (O_331,N_4911,N_4927);
or UO_332 (O_332,N_4900,N_4934);
nand UO_333 (O_333,N_4954,N_4968);
xnor UO_334 (O_334,N_4956,N_4985);
nor UO_335 (O_335,N_4983,N_4959);
and UO_336 (O_336,N_4971,N_4979);
xor UO_337 (O_337,N_4968,N_4939);
nand UO_338 (O_338,N_4960,N_4949);
or UO_339 (O_339,N_4942,N_4967);
nor UO_340 (O_340,N_4911,N_4904);
or UO_341 (O_341,N_4970,N_4955);
xnor UO_342 (O_342,N_4940,N_4989);
xnor UO_343 (O_343,N_4959,N_4981);
nand UO_344 (O_344,N_4967,N_4927);
xnor UO_345 (O_345,N_4973,N_4966);
or UO_346 (O_346,N_4985,N_4954);
nand UO_347 (O_347,N_4948,N_4932);
xnor UO_348 (O_348,N_4993,N_4985);
or UO_349 (O_349,N_4919,N_4982);
and UO_350 (O_350,N_4931,N_4904);
nor UO_351 (O_351,N_4916,N_4949);
or UO_352 (O_352,N_4956,N_4960);
nand UO_353 (O_353,N_4987,N_4923);
xor UO_354 (O_354,N_4986,N_4999);
nand UO_355 (O_355,N_4903,N_4930);
nor UO_356 (O_356,N_4904,N_4917);
nand UO_357 (O_357,N_4907,N_4997);
or UO_358 (O_358,N_4983,N_4915);
nor UO_359 (O_359,N_4918,N_4956);
nand UO_360 (O_360,N_4935,N_4943);
nor UO_361 (O_361,N_4991,N_4948);
xor UO_362 (O_362,N_4920,N_4969);
xor UO_363 (O_363,N_4910,N_4986);
nor UO_364 (O_364,N_4972,N_4915);
or UO_365 (O_365,N_4909,N_4956);
xnor UO_366 (O_366,N_4904,N_4952);
xnor UO_367 (O_367,N_4992,N_4933);
nor UO_368 (O_368,N_4956,N_4961);
xnor UO_369 (O_369,N_4903,N_4912);
and UO_370 (O_370,N_4987,N_4900);
and UO_371 (O_371,N_4988,N_4978);
and UO_372 (O_372,N_4939,N_4910);
nor UO_373 (O_373,N_4924,N_4909);
nor UO_374 (O_374,N_4907,N_4952);
nor UO_375 (O_375,N_4968,N_4946);
nor UO_376 (O_376,N_4984,N_4922);
nand UO_377 (O_377,N_4947,N_4970);
or UO_378 (O_378,N_4922,N_4952);
nor UO_379 (O_379,N_4959,N_4995);
xor UO_380 (O_380,N_4985,N_4996);
and UO_381 (O_381,N_4989,N_4994);
and UO_382 (O_382,N_4987,N_4937);
nand UO_383 (O_383,N_4977,N_4935);
xor UO_384 (O_384,N_4929,N_4924);
nand UO_385 (O_385,N_4941,N_4933);
and UO_386 (O_386,N_4911,N_4961);
xnor UO_387 (O_387,N_4940,N_4941);
or UO_388 (O_388,N_4918,N_4988);
nand UO_389 (O_389,N_4919,N_4908);
and UO_390 (O_390,N_4989,N_4952);
nor UO_391 (O_391,N_4944,N_4925);
and UO_392 (O_392,N_4996,N_4965);
nor UO_393 (O_393,N_4982,N_4935);
nor UO_394 (O_394,N_4963,N_4983);
or UO_395 (O_395,N_4902,N_4938);
and UO_396 (O_396,N_4926,N_4914);
nor UO_397 (O_397,N_4934,N_4999);
nor UO_398 (O_398,N_4916,N_4914);
xor UO_399 (O_399,N_4910,N_4902);
xor UO_400 (O_400,N_4905,N_4987);
or UO_401 (O_401,N_4954,N_4919);
or UO_402 (O_402,N_4953,N_4913);
nor UO_403 (O_403,N_4933,N_4994);
and UO_404 (O_404,N_4980,N_4982);
or UO_405 (O_405,N_4947,N_4913);
nand UO_406 (O_406,N_4994,N_4993);
or UO_407 (O_407,N_4907,N_4958);
nor UO_408 (O_408,N_4934,N_4920);
or UO_409 (O_409,N_4988,N_4990);
xor UO_410 (O_410,N_4970,N_4974);
nand UO_411 (O_411,N_4948,N_4909);
xnor UO_412 (O_412,N_4935,N_4972);
xor UO_413 (O_413,N_4939,N_4948);
or UO_414 (O_414,N_4936,N_4906);
xnor UO_415 (O_415,N_4974,N_4986);
or UO_416 (O_416,N_4933,N_4921);
xnor UO_417 (O_417,N_4907,N_4942);
and UO_418 (O_418,N_4959,N_4977);
and UO_419 (O_419,N_4995,N_4924);
xor UO_420 (O_420,N_4909,N_4926);
and UO_421 (O_421,N_4903,N_4911);
xnor UO_422 (O_422,N_4978,N_4908);
nor UO_423 (O_423,N_4964,N_4943);
xor UO_424 (O_424,N_4918,N_4904);
nor UO_425 (O_425,N_4979,N_4908);
nand UO_426 (O_426,N_4973,N_4983);
xnor UO_427 (O_427,N_4987,N_4988);
nor UO_428 (O_428,N_4960,N_4921);
and UO_429 (O_429,N_4991,N_4919);
xor UO_430 (O_430,N_4970,N_4965);
xnor UO_431 (O_431,N_4986,N_4959);
xor UO_432 (O_432,N_4977,N_4968);
xnor UO_433 (O_433,N_4955,N_4961);
nand UO_434 (O_434,N_4993,N_4914);
nand UO_435 (O_435,N_4993,N_4902);
nand UO_436 (O_436,N_4998,N_4929);
xor UO_437 (O_437,N_4969,N_4967);
xor UO_438 (O_438,N_4981,N_4966);
or UO_439 (O_439,N_4981,N_4921);
nand UO_440 (O_440,N_4984,N_4925);
nor UO_441 (O_441,N_4954,N_4916);
and UO_442 (O_442,N_4952,N_4999);
nor UO_443 (O_443,N_4972,N_4976);
or UO_444 (O_444,N_4979,N_4995);
or UO_445 (O_445,N_4938,N_4956);
xor UO_446 (O_446,N_4943,N_4920);
and UO_447 (O_447,N_4979,N_4936);
nand UO_448 (O_448,N_4929,N_4919);
xnor UO_449 (O_449,N_4911,N_4954);
or UO_450 (O_450,N_4976,N_4944);
nor UO_451 (O_451,N_4955,N_4968);
and UO_452 (O_452,N_4930,N_4986);
or UO_453 (O_453,N_4916,N_4913);
nand UO_454 (O_454,N_4999,N_4958);
nor UO_455 (O_455,N_4930,N_4945);
and UO_456 (O_456,N_4993,N_4916);
nor UO_457 (O_457,N_4945,N_4933);
or UO_458 (O_458,N_4949,N_4993);
xor UO_459 (O_459,N_4907,N_4944);
nor UO_460 (O_460,N_4931,N_4902);
or UO_461 (O_461,N_4911,N_4942);
nor UO_462 (O_462,N_4920,N_4991);
nor UO_463 (O_463,N_4992,N_4973);
or UO_464 (O_464,N_4986,N_4903);
or UO_465 (O_465,N_4950,N_4909);
nand UO_466 (O_466,N_4990,N_4917);
nor UO_467 (O_467,N_4985,N_4952);
nor UO_468 (O_468,N_4960,N_4913);
nor UO_469 (O_469,N_4934,N_4940);
and UO_470 (O_470,N_4955,N_4917);
xnor UO_471 (O_471,N_4990,N_4969);
xnor UO_472 (O_472,N_4932,N_4966);
and UO_473 (O_473,N_4925,N_4966);
or UO_474 (O_474,N_4912,N_4925);
nor UO_475 (O_475,N_4902,N_4955);
or UO_476 (O_476,N_4903,N_4955);
and UO_477 (O_477,N_4990,N_4964);
or UO_478 (O_478,N_4972,N_4947);
and UO_479 (O_479,N_4940,N_4946);
nand UO_480 (O_480,N_4964,N_4908);
nor UO_481 (O_481,N_4937,N_4976);
nand UO_482 (O_482,N_4911,N_4906);
nor UO_483 (O_483,N_4932,N_4921);
or UO_484 (O_484,N_4974,N_4981);
or UO_485 (O_485,N_4956,N_4983);
or UO_486 (O_486,N_4989,N_4967);
and UO_487 (O_487,N_4959,N_4910);
nor UO_488 (O_488,N_4932,N_4920);
nor UO_489 (O_489,N_4981,N_4994);
or UO_490 (O_490,N_4943,N_4960);
nor UO_491 (O_491,N_4921,N_4923);
nor UO_492 (O_492,N_4915,N_4952);
and UO_493 (O_493,N_4931,N_4970);
xnor UO_494 (O_494,N_4962,N_4932);
and UO_495 (O_495,N_4939,N_4958);
nand UO_496 (O_496,N_4972,N_4970);
nor UO_497 (O_497,N_4954,N_4920);
xor UO_498 (O_498,N_4920,N_4974);
or UO_499 (O_499,N_4947,N_4956);
nand UO_500 (O_500,N_4932,N_4933);
xnor UO_501 (O_501,N_4923,N_4963);
and UO_502 (O_502,N_4987,N_4974);
and UO_503 (O_503,N_4977,N_4948);
and UO_504 (O_504,N_4920,N_4983);
xor UO_505 (O_505,N_4916,N_4922);
and UO_506 (O_506,N_4902,N_4959);
or UO_507 (O_507,N_4942,N_4986);
nor UO_508 (O_508,N_4912,N_4974);
and UO_509 (O_509,N_4936,N_4921);
nand UO_510 (O_510,N_4959,N_4944);
xor UO_511 (O_511,N_4988,N_4991);
or UO_512 (O_512,N_4997,N_4974);
xor UO_513 (O_513,N_4969,N_4994);
nor UO_514 (O_514,N_4947,N_4926);
and UO_515 (O_515,N_4960,N_4999);
nand UO_516 (O_516,N_4938,N_4954);
and UO_517 (O_517,N_4980,N_4937);
or UO_518 (O_518,N_4986,N_4907);
xor UO_519 (O_519,N_4957,N_4985);
and UO_520 (O_520,N_4940,N_4977);
nor UO_521 (O_521,N_4927,N_4920);
xor UO_522 (O_522,N_4989,N_4925);
and UO_523 (O_523,N_4999,N_4938);
and UO_524 (O_524,N_4930,N_4952);
xnor UO_525 (O_525,N_4917,N_4963);
and UO_526 (O_526,N_4950,N_4964);
xor UO_527 (O_527,N_4966,N_4939);
xor UO_528 (O_528,N_4978,N_4972);
xor UO_529 (O_529,N_4976,N_4948);
nor UO_530 (O_530,N_4980,N_4933);
nand UO_531 (O_531,N_4933,N_4975);
and UO_532 (O_532,N_4943,N_4937);
and UO_533 (O_533,N_4991,N_4943);
nor UO_534 (O_534,N_4911,N_4973);
nor UO_535 (O_535,N_4991,N_4986);
xnor UO_536 (O_536,N_4958,N_4951);
and UO_537 (O_537,N_4980,N_4924);
nand UO_538 (O_538,N_4911,N_4976);
xnor UO_539 (O_539,N_4945,N_4951);
xor UO_540 (O_540,N_4994,N_4952);
and UO_541 (O_541,N_4912,N_4915);
nor UO_542 (O_542,N_4922,N_4973);
xor UO_543 (O_543,N_4903,N_4932);
and UO_544 (O_544,N_4989,N_4930);
xnor UO_545 (O_545,N_4922,N_4986);
xnor UO_546 (O_546,N_4922,N_4963);
and UO_547 (O_547,N_4986,N_4917);
or UO_548 (O_548,N_4998,N_4985);
and UO_549 (O_549,N_4981,N_4908);
nor UO_550 (O_550,N_4940,N_4913);
and UO_551 (O_551,N_4957,N_4986);
and UO_552 (O_552,N_4920,N_4979);
xnor UO_553 (O_553,N_4981,N_4934);
nand UO_554 (O_554,N_4913,N_4988);
nand UO_555 (O_555,N_4932,N_4989);
xor UO_556 (O_556,N_4920,N_4922);
or UO_557 (O_557,N_4990,N_4925);
and UO_558 (O_558,N_4997,N_4939);
and UO_559 (O_559,N_4974,N_4916);
nand UO_560 (O_560,N_4906,N_4989);
xor UO_561 (O_561,N_4947,N_4923);
nor UO_562 (O_562,N_4948,N_4904);
nor UO_563 (O_563,N_4996,N_4963);
nor UO_564 (O_564,N_4918,N_4933);
xor UO_565 (O_565,N_4960,N_4939);
and UO_566 (O_566,N_4930,N_4957);
nand UO_567 (O_567,N_4923,N_4918);
and UO_568 (O_568,N_4954,N_4939);
nor UO_569 (O_569,N_4953,N_4908);
nand UO_570 (O_570,N_4965,N_4977);
and UO_571 (O_571,N_4986,N_4965);
or UO_572 (O_572,N_4935,N_4918);
nand UO_573 (O_573,N_4900,N_4956);
nor UO_574 (O_574,N_4923,N_4983);
or UO_575 (O_575,N_4911,N_4949);
or UO_576 (O_576,N_4975,N_4969);
and UO_577 (O_577,N_4942,N_4987);
nor UO_578 (O_578,N_4929,N_4914);
and UO_579 (O_579,N_4921,N_4968);
or UO_580 (O_580,N_4921,N_4961);
and UO_581 (O_581,N_4946,N_4988);
or UO_582 (O_582,N_4977,N_4915);
nand UO_583 (O_583,N_4975,N_4902);
nand UO_584 (O_584,N_4984,N_4917);
and UO_585 (O_585,N_4964,N_4918);
xor UO_586 (O_586,N_4980,N_4961);
nor UO_587 (O_587,N_4923,N_4915);
xnor UO_588 (O_588,N_4909,N_4961);
nand UO_589 (O_589,N_4932,N_4904);
or UO_590 (O_590,N_4944,N_4991);
and UO_591 (O_591,N_4926,N_4997);
nor UO_592 (O_592,N_4964,N_4978);
nor UO_593 (O_593,N_4926,N_4950);
nand UO_594 (O_594,N_4946,N_4971);
and UO_595 (O_595,N_4939,N_4932);
nand UO_596 (O_596,N_4992,N_4924);
or UO_597 (O_597,N_4973,N_4978);
xnor UO_598 (O_598,N_4910,N_4951);
xor UO_599 (O_599,N_4955,N_4922);
xnor UO_600 (O_600,N_4966,N_4988);
nor UO_601 (O_601,N_4994,N_4902);
nor UO_602 (O_602,N_4907,N_4983);
nand UO_603 (O_603,N_4944,N_4970);
xnor UO_604 (O_604,N_4908,N_4992);
or UO_605 (O_605,N_4938,N_4972);
nor UO_606 (O_606,N_4971,N_4955);
xor UO_607 (O_607,N_4986,N_4993);
xor UO_608 (O_608,N_4949,N_4978);
or UO_609 (O_609,N_4955,N_4988);
and UO_610 (O_610,N_4910,N_4932);
nor UO_611 (O_611,N_4939,N_4947);
and UO_612 (O_612,N_4985,N_4926);
or UO_613 (O_613,N_4955,N_4997);
nor UO_614 (O_614,N_4988,N_4940);
nand UO_615 (O_615,N_4912,N_4980);
and UO_616 (O_616,N_4934,N_4914);
xnor UO_617 (O_617,N_4900,N_4912);
and UO_618 (O_618,N_4923,N_4920);
nor UO_619 (O_619,N_4956,N_4962);
or UO_620 (O_620,N_4979,N_4945);
or UO_621 (O_621,N_4912,N_4930);
nor UO_622 (O_622,N_4914,N_4940);
xnor UO_623 (O_623,N_4911,N_4947);
nand UO_624 (O_624,N_4998,N_4987);
and UO_625 (O_625,N_4939,N_4994);
and UO_626 (O_626,N_4914,N_4977);
nand UO_627 (O_627,N_4952,N_4959);
nor UO_628 (O_628,N_4910,N_4954);
and UO_629 (O_629,N_4989,N_4920);
nand UO_630 (O_630,N_4923,N_4912);
or UO_631 (O_631,N_4937,N_4959);
xnor UO_632 (O_632,N_4936,N_4954);
xor UO_633 (O_633,N_4926,N_4956);
and UO_634 (O_634,N_4937,N_4932);
nand UO_635 (O_635,N_4967,N_4926);
nor UO_636 (O_636,N_4942,N_4930);
nor UO_637 (O_637,N_4999,N_4974);
xor UO_638 (O_638,N_4990,N_4905);
xnor UO_639 (O_639,N_4949,N_4937);
and UO_640 (O_640,N_4926,N_4932);
and UO_641 (O_641,N_4974,N_4958);
or UO_642 (O_642,N_4938,N_4910);
and UO_643 (O_643,N_4966,N_4970);
nand UO_644 (O_644,N_4984,N_4998);
nor UO_645 (O_645,N_4961,N_4993);
and UO_646 (O_646,N_4938,N_4939);
nand UO_647 (O_647,N_4973,N_4923);
xor UO_648 (O_648,N_4998,N_4988);
nor UO_649 (O_649,N_4944,N_4930);
xor UO_650 (O_650,N_4957,N_4912);
and UO_651 (O_651,N_4908,N_4922);
nand UO_652 (O_652,N_4981,N_4904);
xnor UO_653 (O_653,N_4915,N_4935);
or UO_654 (O_654,N_4927,N_4942);
xnor UO_655 (O_655,N_4976,N_4942);
or UO_656 (O_656,N_4960,N_4919);
and UO_657 (O_657,N_4910,N_4997);
and UO_658 (O_658,N_4933,N_4949);
and UO_659 (O_659,N_4958,N_4918);
or UO_660 (O_660,N_4932,N_4984);
xor UO_661 (O_661,N_4934,N_4956);
nor UO_662 (O_662,N_4948,N_4989);
nor UO_663 (O_663,N_4966,N_4937);
nor UO_664 (O_664,N_4989,N_4959);
and UO_665 (O_665,N_4996,N_4938);
xnor UO_666 (O_666,N_4928,N_4973);
and UO_667 (O_667,N_4919,N_4990);
and UO_668 (O_668,N_4904,N_4979);
nand UO_669 (O_669,N_4953,N_4938);
nand UO_670 (O_670,N_4951,N_4978);
nor UO_671 (O_671,N_4931,N_4941);
nand UO_672 (O_672,N_4993,N_4921);
xnor UO_673 (O_673,N_4929,N_4996);
or UO_674 (O_674,N_4990,N_4981);
and UO_675 (O_675,N_4910,N_4923);
and UO_676 (O_676,N_4993,N_4977);
or UO_677 (O_677,N_4943,N_4954);
and UO_678 (O_678,N_4969,N_4961);
nand UO_679 (O_679,N_4937,N_4911);
or UO_680 (O_680,N_4925,N_4937);
nand UO_681 (O_681,N_4904,N_4916);
and UO_682 (O_682,N_4977,N_4947);
nand UO_683 (O_683,N_4951,N_4953);
nor UO_684 (O_684,N_4985,N_4955);
or UO_685 (O_685,N_4945,N_4916);
nor UO_686 (O_686,N_4968,N_4904);
nor UO_687 (O_687,N_4996,N_4914);
and UO_688 (O_688,N_4997,N_4953);
xnor UO_689 (O_689,N_4920,N_4965);
or UO_690 (O_690,N_4999,N_4968);
and UO_691 (O_691,N_4993,N_4948);
or UO_692 (O_692,N_4960,N_4909);
or UO_693 (O_693,N_4932,N_4965);
and UO_694 (O_694,N_4915,N_4925);
or UO_695 (O_695,N_4981,N_4935);
and UO_696 (O_696,N_4917,N_4945);
xnor UO_697 (O_697,N_4974,N_4984);
xnor UO_698 (O_698,N_4938,N_4915);
nand UO_699 (O_699,N_4966,N_4909);
or UO_700 (O_700,N_4909,N_4945);
and UO_701 (O_701,N_4956,N_4948);
xor UO_702 (O_702,N_4962,N_4926);
nor UO_703 (O_703,N_4945,N_4929);
and UO_704 (O_704,N_4903,N_4997);
xor UO_705 (O_705,N_4952,N_4962);
or UO_706 (O_706,N_4905,N_4994);
or UO_707 (O_707,N_4999,N_4920);
nor UO_708 (O_708,N_4952,N_4929);
nand UO_709 (O_709,N_4947,N_4993);
nand UO_710 (O_710,N_4988,N_4976);
or UO_711 (O_711,N_4958,N_4961);
nand UO_712 (O_712,N_4969,N_4933);
nand UO_713 (O_713,N_4924,N_4943);
xnor UO_714 (O_714,N_4955,N_4934);
and UO_715 (O_715,N_4936,N_4965);
nor UO_716 (O_716,N_4924,N_4981);
nor UO_717 (O_717,N_4973,N_4930);
and UO_718 (O_718,N_4996,N_4950);
or UO_719 (O_719,N_4970,N_4978);
nor UO_720 (O_720,N_4973,N_4937);
or UO_721 (O_721,N_4996,N_4934);
xnor UO_722 (O_722,N_4900,N_4902);
or UO_723 (O_723,N_4904,N_4965);
xnor UO_724 (O_724,N_4948,N_4998);
nand UO_725 (O_725,N_4952,N_4935);
xor UO_726 (O_726,N_4912,N_4991);
or UO_727 (O_727,N_4937,N_4990);
or UO_728 (O_728,N_4905,N_4947);
nor UO_729 (O_729,N_4941,N_4906);
nand UO_730 (O_730,N_4992,N_4910);
nor UO_731 (O_731,N_4934,N_4941);
and UO_732 (O_732,N_4942,N_4902);
nand UO_733 (O_733,N_4999,N_4996);
nor UO_734 (O_734,N_4960,N_4975);
nor UO_735 (O_735,N_4989,N_4950);
nand UO_736 (O_736,N_4959,N_4997);
or UO_737 (O_737,N_4902,N_4986);
nor UO_738 (O_738,N_4963,N_4936);
xnor UO_739 (O_739,N_4956,N_4939);
or UO_740 (O_740,N_4973,N_4940);
nand UO_741 (O_741,N_4985,N_4979);
nor UO_742 (O_742,N_4923,N_4909);
xnor UO_743 (O_743,N_4939,N_4959);
or UO_744 (O_744,N_4982,N_4969);
and UO_745 (O_745,N_4921,N_4956);
or UO_746 (O_746,N_4937,N_4951);
nand UO_747 (O_747,N_4924,N_4977);
nor UO_748 (O_748,N_4941,N_4912);
nor UO_749 (O_749,N_4900,N_4957);
or UO_750 (O_750,N_4939,N_4934);
or UO_751 (O_751,N_4939,N_4983);
xnor UO_752 (O_752,N_4983,N_4949);
and UO_753 (O_753,N_4904,N_4921);
and UO_754 (O_754,N_4982,N_4954);
and UO_755 (O_755,N_4925,N_4980);
or UO_756 (O_756,N_4976,N_4921);
or UO_757 (O_757,N_4993,N_4926);
and UO_758 (O_758,N_4961,N_4957);
nand UO_759 (O_759,N_4947,N_4916);
or UO_760 (O_760,N_4901,N_4966);
xor UO_761 (O_761,N_4971,N_4989);
or UO_762 (O_762,N_4992,N_4994);
nor UO_763 (O_763,N_4997,N_4990);
xor UO_764 (O_764,N_4967,N_4953);
or UO_765 (O_765,N_4918,N_4944);
and UO_766 (O_766,N_4920,N_4987);
or UO_767 (O_767,N_4951,N_4968);
xnor UO_768 (O_768,N_4905,N_4912);
xor UO_769 (O_769,N_4904,N_4927);
nor UO_770 (O_770,N_4950,N_4983);
nand UO_771 (O_771,N_4939,N_4975);
and UO_772 (O_772,N_4984,N_4967);
or UO_773 (O_773,N_4915,N_4945);
nand UO_774 (O_774,N_4948,N_4920);
nor UO_775 (O_775,N_4939,N_4935);
and UO_776 (O_776,N_4946,N_4923);
nor UO_777 (O_777,N_4997,N_4982);
xor UO_778 (O_778,N_4918,N_4925);
or UO_779 (O_779,N_4969,N_4931);
and UO_780 (O_780,N_4917,N_4969);
or UO_781 (O_781,N_4942,N_4952);
nor UO_782 (O_782,N_4977,N_4966);
nor UO_783 (O_783,N_4992,N_4925);
or UO_784 (O_784,N_4927,N_4976);
nor UO_785 (O_785,N_4915,N_4928);
and UO_786 (O_786,N_4947,N_4992);
xnor UO_787 (O_787,N_4943,N_4972);
nand UO_788 (O_788,N_4930,N_4909);
nand UO_789 (O_789,N_4962,N_4968);
or UO_790 (O_790,N_4995,N_4910);
nand UO_791 (O_791,N_4905,N_4965);
nand UO_792 (O_792,N_4949,N_4979);
nor UO_793 (O_793,N_4911,N_4965);
xnor UO_794 (O_794,N_4913,N_4905);
xnor UO_795 (O_795,N_4909,N_4997);
or UO_796 (O_796,N_4916,N_4996);
nor UO_797 (O_797,N_4958,N_4990);
nor UO_798 (O_798,N_4936,N_4950);
or UO_799 (O_799,N_4959,N_4915);
or UO_800 (O_800,N_4957,N_4964);
and UO_801 (O_801,N_4903,N_4913);
and UO_802 (O_802,N_4976,N_4928);
nor UO_803 (O_803,N_4989,N_4987);
or UO_804 (O_804,N_4923,N_4996);
nand UO_805 (O_805,N_4969,N_4910);
or UO_806 (O_806,N_4915,N_4998);
nand UO_807 (O_807,N_4983,N_4902);
and UO_808 (O_808,N_4921,N_4967);
nor UO_809 (O_809,N_4967,N_4959);
or UO_810 (O_810,N_4927,N_4988);
nor UO_811 (O_811,N_4951,N_4952);
xnor UO_812 (O_812,N_4972,N_4964);
xor UO_813 (O_813,N_4907,N_4962);
xnor UO_814 (O_814,N_4915,N_4951);
nor UO_815 (O_815,N_4970,N_4996);
nand UO_816 (O_816,N_4910,N_4940);
or UO_817 (O_817,N_4931,N_4986);
nor UO_818 (O_818,N_4991,N_4999);
xnor UO_819 (O_819,N_4998,N_4916);
xnor UO_820 (O_820,N_4943,N_4993);
nor UO_821 (O_821,N_4918,N_4950);
xnor UO_822 (O_822,N_4953,N_4995);
nor UO_823 (O_823,N_4971,N_4936);
xor UO_824 (O_824,N_4962,N_4916);
nor UO_825 (O_825,N_4989,N_4988);
or UO_826 (O_826,N_4991,N_4909);
nor UO_827 (O_827,N_4960,N_4908);
and UO_828 (O_828,N_4937,N_4917);
xnor UO_829 (O_829,N_4942,N_4994);
nor UO_830 (O_830,N_4984,N_4947);
and UO_831 (O_831,N_4979,N_4916);
and UO_832 (O_832,N_4939,N_4999);
xor UO_833 (O_833,N_4943,N_4929);
nor UO_834 (O_834,N_4975,N_4913);
nand UO_835 (O_835,N_4926,N_4943);
nor UO_836 (O_836,N_4977,N_4984);
or UO_837 (O_837,N_4995,N_4938);
nor UO_838 (O_838,N_4986,N_4988);
or UO_839 (O_839,N_4985,N_4923);
and UO_840 (O_840,N_4911,N_4946);
nand UO_841 (O_841,N_4971,N_4905);
and UO_842 (O_842,N_4970,N_4943);
nor UO_843 (O_843,N_4996,N_4995);
or UO_844 (O_844,N_4930,N_4962);
nand UO_845 (O_845,N_4938,N_4973);
or UO_846 (O_846,N_4941,N_4908);
nor UO_847 (O_847,N_4941,N_4943);
nand UO_848 (O_848,N_4935,N_4923);
nor UO_849 (O_849,N_4955,N_4920);
and UO_850 (O_850,N_4946,N_4975);
nand UO_851 (O_851,N_4989,N_4969);
and UO_852 (O_852,N_4930,N_4916);
or UO_853 (O_853,N_4963,N_4956);
and UO_854 (O_854,N_4973,N_4982);
nand UO_855 (O_855,N_4936,N_4992);
and UO_856 (O_856,N_4940,N_4907);
or UO_857 (O_857,N_4972,N_4953);
xnor UO_858 (O_858,N_4939,N_4913);
nand UO_859 (O_859,N_4977,N_4974);
nor UO_860 (O_860,N_4977,N_4978);
or UO_861 (O_861,N_4916,N_4968);
or UO_862 (O_862,N_4954,N_4905);
or UO_863 (O_863,N_4936,N_4912);
nor UO_864 (O_864,N_4987,N_4931);
and UO_865 (O_865,N_4914,N_4966);
or UO_866 (O_866,N_4969,N_4995);
xnor UO_867 (O_867,N_4974,N_4988);
nor UO_868 (O_868,N_4901,N_4958);
or UO_869 (O_869,N_4944,N_4939);
nand UO_870 (O_870,N_4963,N_4955);
nor UO_871 (O_871,N_4935,N_4905);
or UO_872 (O_872,N_4988,N_4916);
nand UO_873 (O_873,N_4977,N_4941);
nand UO_874 (O_874,N_4989,N_4998);
and UO_875 (O_875,N_4997,N_4985);
xor UO_876 (O_876,N_4978,N_4901);
or UO_877 (O_877,N_4980,N_4955);
nand UO_878 (O_878,N_4920,N_4935);
xnor UO_879 (O_879,N_4962,N_4925);
nand UO_880 (O_880,N_4901,N_4913);
and UO_881 (O_881,N_4939,N_4936);
nand UO_882 (O_882,N_4936,N_4983);
nor UO_883 (O_883,N_4945,N_4940);
xor UO_884 (O_884,N_4924,N_4960);
nand UO_885 (O_885,N_4937,N_4919);
nand UO_886 (O_886,N_4985,N_4922);
and UO_887 (O_887,N_4956,N_4936);
or UO_888 (O_888,N_4982,N_4949);
and UO_889 (O_889,N_4941,N_4959);
and UO_890 (O_890,N_4928,N_4941);
nand UO_891 (O_891,N_4990,N_4949);
xor UO_892 (O_892,N_4939,N_4984);
nand UO_893 (O_893,N_4950,N_4920);
nor UO_894 (O_894,N_4917,N_4994);
nor UO_895 (O_895,N_4984,N_4975);
and UO_896 (O_896,N_4978,N_4914);
and UO_897 (O_897,N_4920,N_4933);
nand UO_898 (O_898,N_4980,N_4950);
nand UO_899 (O_899,N_4960,N_4979);
or UO_900 (O_900,N_4994,N_4995);
or UO_901 (O_901,N_4936,N_4915);
nand UO_902 (O_902,N_4922,N_4942);
and UO_903 (O_903,N_4935,N_4938);
nand UO_904 (O_904,N_4977,N_4999);
and UO_905 (O_905,N_4953,N_4948);
nand UO_906 (O_906,N_4968,N_4944);
xnor UO_907 (O_907,N_4932,N_4925);
nand UO_908 (O_908,N_4965,N_4943);
xor UO_909 (O_909,N_4990,N_4901);
or UO_910 (O_910,N_4913,N_4986);
and UO_911 (O_911,N_4916,N_4941);
xor UO_912 (O_912,N_4955,N_4989);
xor UO_913 (O_913,N_4977,N_4931);
nor UO_914 (O_914,N_4954,N_4956);
xor UO_915 (O_915,N_4936,N_4916);
or UO_916 (O_916,N_4934,N_4970);
nand UO_917 (O_917,N_4968,N_4917);
xor UO_918 (O_918,N_4974,N_4917);
and UO_919 (O_919,N_4990,N_4918);
nor UO_920 (O_920,N_4998,N_4990);
nand UO_921 (O_921,N_4928,N_4978);
nand UO_922 (O_922,N_4988,N_4931);
nor UO_923 (O_923,N_4956,N_4929);
xnor UO_924 (O_924,N_4928,N_4906);
and UO_925 (O_925,N_4927,N_4952);
or UO_926 (O_926,N_4922,N_4944);
xnor UO_927 (O_927,N_4992,N_4948);
nor UO_928 (O_928,N_4952,N_4965);
and UO_929 (O_929,N_4917,N_4940);
or UO_930 (O_930,N_4924,N_4932);
and UO_931 (O_931,N_4985,N_4937);
xnor UO_932 (O_932,N_4942,N_4946);
nand UO_933 (O_933,N_4925,N_4947);
xnor UO_934 (O_934,N_4979,N_4955);
and UO_935 (O_935,N_4986,N_4987);
or UO_936 (O_936,N_4970,N_4922);
nor UO_937 (O_937,N_4982,N_4984);
or UO_938 (O_938,N_4985,N_4978);
and UO_939 (O_939,N_4948,N_4908);
nand UO_940 (O_940,N_4920,N_4963);
and UO_941 (O_941,N_4947,N_4928);
or UO_942 (O_942,N_4901,N_4985);
nand UO_943 (O_943,N_4956,N_4923);
nand UO_944 (O_944,N_4980,N_4965);
nand UO_945 (O_945,N_4931,N_4965);
xor UO_946 (O_946,N_4986,N_4995);
nor UO_947 (O_947,N_4951,N_4967);
or UO_948 (O_948,N_4921,N_4902);
and UO_949 (O_949,N_4941,N_4949);
nor UO_950 (O_950,N_4922,N_4983);
and UO_951 (O_951,N_4987,N_4956);
or UO_952 (O_952,N_4975,N_4931);
or UO_953 (O_953,N_4957,N_4907);
nand UO_954 (O_954,N_4998,N_4946);
and UO_955 (O_955,N_4964,N_4987);
or UO_956 (O_956,N_4921,N_4905);
xnor UO_957 (O_957,N_4992,N_4904);
nand UO_958 (O_958,N_4975,N_4964);
nand UO_959 (O_959,N_4945,N_4994);
and UO_960 (O_960,N_4946,N_4973);
nor UO_961 (O_961,N_4929,N_4961);
or UO_962 (O_962,N_4997,N_4934);
xor UO_963 (O_963,N_4974,N_4923);
or UO_964 (O_964,N_4933,N_4979);
nor UO_965 (O_965,N_4953,N_4962);
nor UO_966 (O_966,N_4982,N_4958);
and UO_967 (O_967,N_4998,N_4981);
or UO_968 (O_968,N_4998,N_4917);
xor UO_969 (O_969,N_4953,N_4955);
nor UO_970 (O_970,N_4908,N_4916);
and UO_971 (O_971,N_4952,N_4973);
and UO_972 (O_972,N_4934,N_4929);
or UO_973 (O_973,N_4905,N_4963);
and UO_974 (O_974,N_4961,N_4974);
nand UO_975 (O_975,N_4976,N_4965);
nor UO_976 (O_976,N_4961,N_4942);
xor UO_977 (O_977,N_4933,N_4990);
or UO_978 (O_978,N_4903,N_4924);
nand UO_979 (O_979,N_4979,N_4962);
xnor UO_980 (O_980,N_4994,N_4914);
and UO_981 (O_981,N_4949,N_4912);
nor UO_982 (O_982,N_4920,N_4929);
nand UO_983 (O_983,N_4938,N_4967);
nor UO_984 (O_984,N_4925,N_4914);
nand UO_985 (O_985,N_4970,N_4962);
and UO_986 (O_986,N_4992,N_4967);
xnor UO_987 (O_987,N_4904,N_4966);
and UO_988 (O_988,N_4974,N_4945);
nor UO_989 (O_989,N_4959,N_4926);
nor UO_990 (O_990,N_4956,N_4996);
or UO_991 (O_991,N_4982,N_4910);
nand UO_992 (O_992,N_4914,N_4945);
nor UO_993 (O_993,N_4902,N_4964);
nand UO_994 (O_994,N_4983,N_4971);
nor UO_995 (O_995,N_4913,N_4934);
nor UO_996 (O_996,N_4959,N_4908);
or UO_997 (O_997,N_4959,N_4942);
or UO_998 (O_998,N_4903,N_4946);
xor UO_999 (O_999,N_4941,N_4953);
endmodule