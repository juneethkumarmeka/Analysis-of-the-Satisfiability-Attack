module basic_500_3000_500_3_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_350,In_250);
nand U1 (N_1,In_473,In_283);
nand U2 (N_2,In_342,In_437);
nor U3 (N_3,In_388,In_67);
and U4 (N_4,In_228,In_58);
nor U5 (N_5,In_259,In_212);
nor U6 (N_6,In_30,In_293);
and U7 (N_7,In_211,In_2);
or U8 (N_8,In_97,In_475);
and U9 (N_9,In_296,In_420);
nand U10 (N_10,In_221,In_76);
or U11 (N_11,In_9,In_251);
and U12 (N_12,In_80,In_155);
nor U13 (N_13,In_143,In_215);
nor U14 (N_14,In_268,In_75);
or U15 (N_15,In_219,In_282);
xnor U16 (N_16,In_375,In_112);
and U17 (N_17,In_148,In_305);
nand U18 (N_18,In_216,In_156);
nand U19 (N_19,In_175,In_429);
or U20 (N_20,In_40,In_416);
or U21 (N_21,In_37,In_399);
or U22 (N_22,In_363,In_263);
and U23 (N_23,In_418,In_207);
nand U24 (N_24,In_131,In_371);
and U25 (N_25,In_455,In_186);
or U26 (N_26,In_33,In_272);
nor U27 (N_27,In_482,In_379);
nand U28 (N_28,In_391,In_410);
nand U29 (N_29,In_73,In_306);
and U30 (N_30,In_334,In_213);
nor U31 (N_31,In_43,In_88);
and U32 (N_32,In_494,In_360);
nor U33 (N_33,In_61,In_466);
and U34 (N_34,In_394,In_280);
nand U35 (N_35,In_49,In_159);
or U36 (N_36,In_173,In_140);
nor U37 (N_37,In_498,In_191);
and U38 (N_38,In_8,In_493);
nor U39 (N_39,In_474,In_315);
nor U40 (N_40,In_258,In_65);
and U41 (N_41,In_181,In_165);
and U42 (N_42,In_29,In_101);
and U43 (N_43,In_337,In_68);
and U44 (N_44,In_446,In_415);
or U45 (N_45,In_166,In_271);
and U46 (N_46,In_374,In_190);
nor U47 (N_47,In_402,In_430);
and U48 (N_48,In_380,In_208);
nand U49 (N_49,In_260,In_93);
nand U50 (N_50,In_161,In_352);
nor U51 (N_51,In_254,In_425);
or U52 (N_52,In_96,In_64);
nor U53 (N_53,In_123,In_324);
or U54 (N_54,In_274,In_486);
nor U55 (N_55,In_206,In_104);
nand U56 (N_56,In_339,In_257);
nor U57 (N_57,In_318,In_434);
nand U58 (N_58,In_92,In_397);
nor U59 (N_59,In_309,In_365);
nor U60 (N_60,In_362,In_433);
and U61 (N_61,In_39,In_330);
nor U62 (N_62,In_338,In_264);
nor U63 (N_63,In_193,In_141);
or U64 (N_64,In_133,In_162);
nor U65 (N_65,In_55,In_361);
nand U66 (N_66,In_115,In_202);
or U67 (N_67,In_203,In_421);
nand U68 (N_68,In_12,In_21);
or U69 (N_69,In_78,In_103);
or U70 (N_70,In_378,In_79);
nand U71 (N_71,In_403,In_303);
nor U72 (N_72,In_1,In_479);
nor U73 (N_73,In_273,In_354);
nor U74 (N_74,In_428,In_495);
or U75 (N_75,In_441,In_89);
or U76 (N_76,In_470,In_16);
or U77 (N_77,In_314,In_146);
or U78 (N_78,In_333,In_460);
or U79 (N_79,In_99,In_328);
nor U80 (N_80,In_347,In_6);
and U81 (N_81,In_329,In_147);
nand U82 (N_82,In_356,In_438);
nand U83 (N_83,In_126,In_246);
nand U84 (N_84,In_138,In_381);
xnor U85 (N_85,In_270,In_50);
nor U86 (N_86,In_46,In_366);
xor U87 (N_87,In_467,In_152);
and U88 (N_88,In_239,In_226);
nor U89 (N_89,In_195,In_277);
or U90 (N_90,In_163,In_431);
nand U91 (N_91,In_368,In_436);
nand U92 (N_92,In_139,In_462);
nand U93 (N_93,In_426,In_313);
or U94 (N_94,In_13,In_154);
xor U95 (N_95,In_192,In_201);
nand U96 (N_96,In_320,In_308);
nand U97 (N_97,In_449,In_35);
nand U98 (N_98,In_18,In_160);
and U99 (N_99,In_164,In_122);
nor U100 (N_100,In_84,In_340);
and U101 (N_101,In_177,In_188);
and U102 (N_102,In_405,In_174);
nand U103 (N_103,In_278,In_15);
nand U104 (N_104,In_336,In_102);
nor U105 (N_105,In_71,In_419);
nand U106 (N_106,In_236,In_265);
nor U107 (N_107,In_396,In_376);
and U108 (N_108,In_204,In_243);
and U109 (N_109,In_456,In_233);
or U110 (N_110,In_294,In_52);
or U111 (N_111,In_59,In_86);
nand U112 (N_112,In_241,In_407);
or U113 (N_113,In_34,In_158);
or U114 (N_114,In_244,In_497);
nand U115 (N_115,In_288,In_325);
xnor U116 (N_116,In_414,In_432);
nor U117 (N_117,In_284,In_448);
nor U118 (N_118,In_121,In_304);
or U119 (N_119,In_232,In_105);
or U120 (N_120,In_25,In_279);
and U121 (N_121,In_180,In_222);
or U122 (N_122,In_491,In_44);
nor U123 (N_123,In_41,In_27);
nand U124 (N_124,In_286,In_287);
nand U125 (N_125,In_297,In_157);
nor U126 (N_126,In_401,In_469);
nor U127 (N_127,In_36,In_344);
or U128 (N_128,In_178,In_38);
nand U129 (N_129,In_345,In_220);
or U130 (N_130,In_24,In_0);
or U131 (N_131,In_171,In_323);
nor U132 (N_132,In_468,In_179);
nand U133 (N_133,In_307,In_47);
nor U134 (N_134,In_217,In_377);
and U135 (N_135,In_487,In_302);
nor U136 (N_136,In_31,In_463);
nor U137 (N_137,In_404,In_214);
and U138 (N_138,In_176,In_245);
nand U139 (N_139,In_83,In_189);
nand U140 (N_140,In_234,In_316);
nor U141 (N_141,In_477,In_488);
or U142 (N_142,In_382,In_137);
and U143 (N_143,In_94,In_172);
nor U144 (N_144,In_348,In_230);
or U145 (N_145,In_247,In_332);
or U146 (N_146,In_117,In_132);
nor U147 (N_147,In_10,In_136);
or U148 (N_148,In_372,In_276);
nand U149 (N_149,In_184,In_224);
and U150 (N_150,In_484,In_128);
nand U151 (N_151,In_134,In_406);
or U152 (N_152,In_3,In_261);
or U153 (N_153,In_398,In_107);
or U154 (N_154,In_390,In_341);
and U155 (N_155,In_223,In_125);
or U156 (N_156,In_472,In_321);
or U157 (N_157,In_235,In_269);
nor U158 (N_158,In_292,In_311);
and U159 (N_159,In_322,In_77);
and U160 (N_160,In_343,In_11);
and U161 (N_161,In_295,In_422);
nor U162 (N_162,In_48,In_225);
and U163 (N_163,In_481,In_256);
and U164 (N_164,In_490,In_227);
nand U165 (N_165,In_119,In_262);
or U166 (N_166,In_28,In_442);
or U167 (N_167,In_301,In_127);
or U168 (N_168,In_182,In_300);
nand U169 (N_169,In_54,In_349);
or U170 (N_170,In_478,In_317);
and U171 (N_171,In_400,In_389);
nor U172 (N_172,In_267,In_253);
xor U173 (N_173,In_185,In_395);
and U174 (N_174,In_82,In_298);
and U175 (N_175,In_106,In_110);
and U176 (N_176,In_22,In_445);
nor U177 (N_177,In_145,In_450);
and U178 (N_178,In_238,In_205);
nor U179 (N_179,In_423,In_57);
nor U180 (N_180,In_95,In_5);
or U181 (N_181,In_26,In_447);
nand U182 (N_182,In_335,In_369);
xnor U183 (N_183,In_7,In_385);
nor U184 (N_184,In_461,In_499);
and U185 (N_185,In_116,In_364);
and U186 (N_186,In_496,In_454);
nor U187 (N_187,In_231,In_74);
nor U188 (N_188,In_413,In_383);
nor U189 (N_189,In_109,In_209);
nor U190 (N_190,In_87,In_151);
and U191 (N_191,In_62,In_476);
nand U192 (N_192,In_480,In_142);
nor U193 (N_193,In_60,In_319);
or U194 (N_194,In_124,In_457);
or U195 (N_195,In_440,In_153);
nand U196 (N_196,In_199,In_310);
nand U197 (N_197,In_483,In_444);
or U198 (N_198,In_45,In_144);
nor U199 (N_199,In_453,In_100);
nand U200 (N_200,In_130,In_19);
and U201 (N_201,In_69,In_285);
nor U202 (N_202,In_489,In_4);
nand U203 (N_203,In_427,In_240);
xnor U204 (N_204,In_70,In_194);
and U205 (N_205,In_443,In_187);
and U206 (N_206,In_168,In_120);
nand U207 (N_207,In_51,In_56);
or U208 (N_208,In_459,In_464);
or U209 (N_209,In_290,In_417);
and U210 (N_210,In_358,In_108);
or U211 (N_211,In_218,In_424);
or U212 (N_212,In_242,In_266);
nand U213 (N_213,In_118,In_465);
or U214 (N_214,In_357,In_312);
and U215 (N_215,In_412,In_275);
and U216 (N_216,In_66,In_169);
and U217 (N_217,In_252,In_435);
or U218 (N_218,In_85,In_197);
and U219 (N_219,In_370,In_327);
nand U220 (N_220,In_458,In_485);
nand U221 (N_221,In_359,In_20);
and U222 (N_222,In_90,In_113);
nor U223 (N_223,In_299,In_196);
nand U224 (N_224,In_281,In_392);
nand U225 (N_225,In_411,In_439);
and U226 (N_226,In_408,In_170);
nor U227 (N_227,In_167,In_237);
and U228 (N_228,In_210,In_387);
or U229 (N_229,In_72,In_373);
nand U230 (N_230,In_53,In_150);
nand U231 (N_231,In_98,In_91);
nor U232 (N_232,In_81,In_331);
or U233 (N_233,In_346,In_289);
nand U234 (N_234,In_384,In_386);
nand U235 (N_235,In_14,In_248);
and U236 (N_236,In_129,In_351);
nor U237 (N_237,In_326,In_393);
and U238 (N_238,In_452,In_114);
nand U239 (N_239,In_32,In_409);
xnor U240 (N_240,In_17,In_42);
nor U241 (N_241,In_291,In_229);
or U242 (N_242,In_198,In_471);
nand U243 (N_243,In_23,In_200);
and U244 (N_244,In_353,In_249);
nor U245 (N_245,In_135,In_355);
and U246 (N_246,In_111,In_367);
nor U247 (N_247,In_451,In_183);
or U248 (N_248,In_492,In_63);
nand U249 (N_249,In_255,In_149);
or U250 (N_250,In_374,In_22);
nor U251 (N_251,In_241,In_417);
nand U252 (N_252,In_364,In_458);
xnor U253 (N_253,In_260,In_178);
nand U254 (N_254,In_388,In_495);
or U255 (N_255,In_328,In_173);
nor U256 (N_256,In_291,In_347);
nand U257 (N_257,In_474,In_230);
nand U258 (N_258,In_31,In_277);
and U259 (N_259,In_443,In_409);
and U260 (N_260,In_448,In_463);
and U261 (N_261,In_249,In_383);
nand U262 (N_262,In_486,In_131);
nor U263 (N_263,In_97,In_434);
xnor U264 (N_264,In_201,In_127);
or U265 (N_265,In_237,In_21);
nand U266 (N_266,In_417,In_448);
or U267 (N_267,In_307,In_133);
nand U268 (N_268,In_214,In_144);
nand U269 (N_269,In_368,In_231);
xnor U270 (N_270,In_91,In_7);
nand U271 (N_271,In_251,In_29);
or U272 (N_272,In_483,In_376);
nor U273 (N_273,In_227,In_331);
nor U274 (N_274,In_193,In_445);
and U275 (N_275,In_272,In_269);
or U276 (N_276,In_129,In_204);
nand U277 (N_277,In_180,In_209);
or U278 (N_278,In_253,In_31);
nor U279 (N_279,In_201,In_68);
or U280 (N_280,In_149,In_475);
nor U281 (N_281,In_293,In_291);
and U282 (N_282,In_342,In_288);
nand U283 (N_283,In_289,In_422);
or U284 (N_284,In_310,In_346);
nor U285 (N_285,In_13,In_29);
or U286 (N_286,In_187,In_299);
nor U287 (N_287,In_482,In_30);
nor U288 (N_288,In_34,In_146);
or U289 (N_289,In_89,In_234);
and U290 (N_290,In_297,In_190);
and U291 (N_291,In_179,In_277);
or U292 (N_292,In_360,In_392);
nand U293 (N_293,In_238,In_474);
nor U294 (N_294,In_279,In_256);
nand U295 (N_295,In_196,In_38);
nor U296 (N_296,In_344,In_429);
xor U297 (N_297,In_459,In_181);
or U298 (N_298,In_438,In_347);
or U299 (N_299,In_471,In_14);
and U300 (N_300,In_448,In_207);
nand U301 (N_301,In_377,In_375);
and U302 (N_302,In_161,In_494);
nand U303 (N_303,In_353,In_243);
nand U304 (N_304,In_336,In_386);
nand U305 (N_305,In_468,In_109);
nor U306 (N_306,In_448,In_243);
nor U307 (N_307,In_202,In_188);
nor U308 (N_308,In_405,In_289);
and U309 (N_309,In_358,In_279);
and U310 (N_310,In_47,In_77);
or U311 (N_311,In_375,In_36);
or U312 (N_312,In_443,In_71);
and U313 (N_313,In_177,In_28);
or U314 (N_314,In_396,In_162);
nand U315 (N_315,In_63,In_268);
nor U316 (N_316,In_387,In_131);
or U317 (N_317,In_323,In_27);
nor U318 (N_318,In_442,In_64);
or U319 (N_319,In_329,In_430);
and U320 (N_320,In_472,In_53);
nor U321 (N_321,In_452,In_403);
and U322 (N_322,In_453,In_440);
and U323 (N_323,In_323,In_314);
xor U324 (N_324,In_153,In_117);
nand U325 (N_325,In_198,In_432);
nand U326 (N_326,In_12,In_0);
nor U327 (N_327,In_378,In_271);
nor U328 (N_328,In_176,In_388);
and U329 (N_329,In_380,In_386);
and U330 (N_330,In_298,In_273);
or U331 (N_331,In_191,In_367);
nor U332 (N_332,In_67,In_92);
nand U333 (N_333,In_242,In_371);
or U334 (N_334,In_496,In_18);
nor U335 (N_335,In_126,In_108);
and U336 (N_336,In_295,In_380);
or U337 (N_337,In_314,In_390);
nor U338 (N_338,In_182,In_380);
nand U339 (N_339,In_348,In_28);
nand U340 (N_340,In_173,In_339);
or U341 (N_341,In_113,In_413);
nor U342 (N_342,In_72,In_289);
or U343 (N_343,In_94,In_456);
and U344 (N_344,In_301,In_62);
nor U345 (N_345,In_123,In_74);
or U346 (N_346,In_248,In_400);
or U347 (N_347,In_183,In_186);
nand U348 (N_348,In_233,In_484);
and U349 (N_349,In_479,In_442);
and U350 (N_350,In_376,In_454);
nor U351 (N_351,In_410,In_474);
nand U352 (N_352,In_182,In_378);
or U353 (N_353,In_94,In_206);
nor U354 (N_354,In_167,In_305);
and U355 (N_355,In_304,In_169);
nand U356 (N_356,In_459,In_204);
or U357 (N_357,In_199,In_85);
or U358 (N_358,In_261,In_36);
nor U359 (N_359,In_273,In_406);
nor U360 (N_360,In_301,In_448);
or U361 (N_361,In_489,In_48);
nand U362 (N_362,In_17,In_389);
or U363 (N_363,In_493,In_398);
nand U364 (N_364,In_462,In_255);
and U365 (N_365,In_403,In_30);
and U366 (N_366,In_244,In_113);
or U367 (N_367,In_487,In_125);
nor U368 (N_368,In_52,In_115);
nor U369 (N_369,In_227,In_34);
and U370 (N_370,In_122,In_286);
nand U371 (N_371,In_60,In_96);
nor U372 (N_372,In_22,In_406);
xor U373 (N_373,In_100,In_45);
and U374 (N_374,In_389,In_336);
nor U375 (N_375,In_358,In_390);
and U376 (N_376,In_396,In_332);
or U377 (N_377,In_323,In_282);
nand U378 (N_378,In_479,In_191);
and U379 (N_379,In_94,In_394);
and U380 (N_380,In_357,In_421);
and U381 (N_381,In_388,In_151);
and U382 (N_382,In_259,In_230);
or U383 (N_383,In_73,In_262);
nand U384 (N_384,In_357,In_347);
and U385 (N_385,In_290,In_186);
nor U386 (N_386,In_282,In_313);
and U387 (N_387,In_342,In_28);
xor U388 (N_388,In_328,In_25);
nor U389 (N_389,In_384,In_289);
nor U390 (N_390,In_400,In_161);
nor U391 (N_391,In_105,In_249);
and U392 (N_392,In_70,In_258);
nor U393 (N_393,In_151,In_113);
nand U394 (N_394,In_204,In_211);
and U395 (N_395,In_493,In_445);
and U396 (N_396,In_144,In_160);
or U397 (N_397,In_69,In_282);
or U398 (N_398,In_44,In_43);
nand U399 (N_399,In_278,In_103);
nand U400 (N_400,In_45,In_300);
or U401 (N_401,In_94,In_414);
nor U402 (N_402,In_64,In_180);
and U403 (N_403,In_388,In_380);
and U404 (N_404,In_420,In_95);
nand U405 (N_405,In_118,In_394);
or U406 (N_406,In_43,In_0);
nand U407 (N_407,In_212,In_3);
or U408 (N_408,In_158,In_441);
and U409 (N_409,In_488,In_71);
xnor U410 (N_410,In_495,In_249);
or U411 (N_411,In_144,In_391);
and U412 (N_412,In_475,In_334);
nand U413 (N_413,In_457,In_348);
nand U414 (N_414,In_194,In_104);
xor U415 (N_415,In_311,In_207);
nor U416 (N_416,In_409,In_46);
and U417 (N_417,In_423,In_229);
nor U418 (N_418,In_297,In_46);
or U419 (N_419,In_7,In_254);
nand U420 (N_420,In_453,In_318);
or U421 (N_421,In_198,In_30);
nor U422 (N_422,In_30,In_71);
nor U423 (N_423,In_93,In_204);
and U424 (N_424,In_244,In_458);
nand U425 (N_425,In_462,In_358);
nor U426 (N_426,In_367,In_436);
nand U427 (N_427,In_204,In_177);
nor U428 (N_428,In_254,In_400);
or U429 (N_429,In_17,In_407);
nor U430 (N_430,In_213,In_88);
and U431 (N_431,In_132,In_203);
nor U432 (N_432,In_239,In_499);
nand U433 (N_433,In_217,In_438);
nor U434 (N_434,In_14,In_469);
nor U435 (N_435,In_100,In_245);
or U436 (N_436,In_454,In_261);
nand U437 (N_437,In_367,In_269);
and U438 (N_438,In_338,In_376);
nand U439 (N_439,In_399,In_58);
and U440 (N_440,In_279,In_430);
or U441 (N_441,In_52,In_332);
or U442 (N_442,In_367,In_278);
or U443 (N_443,In_221,In_26);
or U444 (N_444,In_198,In_448);
nand U445 (N_445,In_154,In_254);
or U446 (N_446,In_415,In_183);
or U447 (N_447,In_481,In_56);
or U448 (N_448,In_80,In_246);
nor U449 (N_449,In_401,In_457);
nor U450 (N_450,In_208,In_303);
nand U451 (N_451,In_50,In_448);
nand U452 (N_452,In_146,In_479);
nand U453 (N_453,In_282,In_199);
nor U454 (N_454,In_202,In_172);
nor U455 (N_455,In_193,In_414);
and U456 (N_456,In_123,In_141);
nand U457 (N_457,In_302,In_243);
and U458 (N_458,In_35,In_313);
or U459 (N_459,In_119,In_308);
nor U460 (N_460,In_154,In_336);
and U461 (N_461,In_211,In_223);
and U462 (N_462,In_275,In_147);
nand U463 (N_463,In_441,In_276);
and U464 (N_464,In_371,In_123);
nor U465 (N_465,In_496,In_169);
nand U466 (N_466,In_347,In_340);
or U467 (N_467,In_109,In_336);
and U468 (N_468,In_305,In_394);
nor U469 (N_469,In_133,In_85);
nand U470 (N_470,In_176,In_37);
or U471 (N_471,In_63,In_466);
and U472 (N_472,In_488,In_28);
nand U473 (N_473,In_17,In_40);
nor U474 (N_474,In_394,In_397);
nand U475 (N_475,In_278,In_169);
and U476 (N_476,In_278,In_157);
and U477 (N_477,In_217,In_238);
nand U478 (N_478,In_325,In_287);
or U479 (N_479,In_461,In_474);
and U480 (N_480,In_297,In_478);
or U481 (N_481,In_228,In_22);
and U482 (N_482,In_300,In_200);
nand U483 (N_483,In_408,In_57);
nor U484 (N_484,In_462,In_443);
and U485 (N_485,In_343,In_302);
nor U486 (N_486,In_264,In_403);
nand U487 (N_487,In_13,In_403);
nand U488 (N_488,In_247,In_44);
nor U489 (N_489,In_376,In_448);
and U490 (N_490,In_88,In_62);
nand U491 (N_491,In_45,In_352);
and U492 (N_492,In_233,In_375);
nor U493 (N_493,In_264,In_129);
xnor U494 (N_494,In_310,In_151);
or U495 (N_495,In_307,In_66);
or U496 (N_496,In_336,In_173);
and U497 (N_497,In_439,In_90);
and U498 (N_498,In_428,In_382);
nor U499 (N_499,In_204,In_286);
or U500 (N_500,In_260,In_374);
nor U501 (N_501,In_12,In_407);
nand U502 (N_502,In_433,In_223);
and U503 (N_503,In_444,In_339);
or U504 (N_504,In_2,In_293);
nand U505 (N_505,In_330,In_490);
or U506 (N_506,In_50,In_142);
or U507 (N_507,In_186,In_70);
nand U508 (N_508,In_398,In_490);
nand U509 (N_509,In_456,In_115);
xor U510 (N_510,In_184,In_421);
or U511 (N_511,In_92,In_120);
or U512 (N_512,In_435,In_368);
nand U513 (N_513,In_281,In_261);
and U514 (N_514,In_140,In_71);
nor U515 (N_515,In_447,In_125);
nor U516 (N_516,In_127,In_481);
nand U517 (N_517,In_59,In_380);
nand U518 (N_518,In_225,In_101);
or U519 (N_519,In_142,In_438);
nor U520 (N_520,In_485,In_402);
nand U521 (N_521,In_397,In_378);
or U522 (N_522,In_498,In_227);
nand U523 (N_523,In_230,In_189);
and U524 (N_524,In_46,In_261);
and U525 (N_525,In_464,In_63);
and U526 (N_526,In_189,In_4);
or U527 (N_527,In_400,In_92);
nor U528 (N_528,In_439,In_220);
nor U529 (N_529,In_359,In_365);
nor U530 (N_530,In_262,In_3);
and U531 (N_531,In_74,In_394);
or U532 (N_532,In_416,In_348);
nand U533 (N_533,In_314,In_243);
or U534 (N_534,In_313,In_190);
and U535 (N_535,In_82,In_31);
and U536 (N_536,In_134,In_178);
and U537 (N_537,In_22,In_326);
nor U538 (N_538,In_99,In_305);
and U539 (N_539,In_337,In_10);
nand U540 (N_540,In_411,In_384);
nand U541 (N_541,In_222,In_388);
nor U542 (N_542,In_478,In_409);
nor U543 (N_543,In_238,In_142);
nand U544 (N_544,In_436,In_386);
or U545 (N_545,In_237,In_4);
or U546 (N_546,In_253,In_76);
nand U547 (N_547,In_80,In_471);
and U548 (N_548,In_435,In_384);
or U549 (N_549,In_168,In_109);
nand U550 (N_550,In_106,In_427);
and U551 (N_551,In_159,In_150);
or U552 (N_552,In_251,In_321);
nor U553 (N_553,In_369,In_30);
and U554 (N_554,In_261,In_323);
or U555 (N_555,In_365,In_40);
nand U556 (N_556,In_128,In_372);
or U557 (N_557,In_9,In_495);
nand U558 (N_558,In_92,In_387);
and U559 (N_559,In_448,In_195);
and U560 (N_560,In_302,In_494);
nor U561 (N_561,In_268,In_208);
and U562 (N_562,In_448,In_350);
or U563 (N_563,In_316,In_272);
or U564 (N_564,In_437,In_117);
and U565 (N_565,In_91,In_430);
nand U566 (N_566,In_496,In_139);
nand U567 (N_567,In_54,In_192);
and U568 (N_568,In_247,In_197);
nor U569 (N_569,In_105,In_208);
nand U570 (N_570,In_413,In_341);
and U571 (N_571,In_280,In_125);
nor U572 (N_572,In_419,In_217);
nor U573 (N_573,In_207,In_180);
and U574 (N_574,In_313,In_119);
nand U575 (N_575,In_295,In_341);
nor U576 (N_576,In_421,In_23);
or U577 (N_577,In_429,In_28);
or U578 (N_578,In_410,In_200);
and U579 (N_579,In_231,In_146);
nor U580 (N_580,In_140,In_468);
nand U581 (N_581,In_381,In_62);
or U582 (N_582,In_291,In_183);
xnor U583 (N_583,In_70,In_332);
nand U584 (N_584,In_466,In_234);
and U585 (N_585,In_323,In_457);
and U586 (N_586,In_351,In_416);
and U587 (N_587,In_222,In_26);
and U588 (N_588,In_26,In_7);
and U589 (N_589,In_162,In_305);
nor U590 (N_590,In_317,In_322);
nand U591 (N_591,In_187,In_457);
or U592 (N_592,In_24,In_346);
or U593 (N_593,In_222,In_177);
and U594 (N_594,In_153,In_488);
and U595 (N_595,In_279,In_40);
nand U596 (N_596,In_338,In_13);
nor U597 (N_597,In_156,In_174);
or U598 (N_598,In_293,In_187);
nor U599 (N_599,In_447,In_185);
or U600 (N_600,In_390,In_115);
nand U601 (N_601,In_270,In_147);
or U602 (N_602,In_236,In_427);
nand U603 (N_603,In_263,In_441);
or U604 (N_604,In_282,In_96);
nor U605 (N_605,In_332,In_474);
nor U606 (N_606,In_312,In_121);
and U607 (N_607,In_7,In_78);
and U608 (N_608,In_197,In_318);
and U609 (N_609,In_4,In_386);
nor U610 (N_610,In_63,In_284);
and U611 (N_611,In_234,In_37);
nor U612 (N_612,In_380,In_184);
or U613 (N_613,In_480,In_219);
or U614 (N_614,In_280,In_441);
or U615 (N_615,In_303,In_61);
and U616 (N_616,In_61,In_329);
and U617 (N_617,In_272,In_220);
nor U618 (N_618,In_212,In_12);
or U619 (N_619,In_83,In_227);
nand U620 (N_620,In_213,In_225);
nand U621 (N_621,In_314,In_410);
nor U622 (N_622,In_99,In_442);
or U623 (N_623,In_19,In_203);
and U624 (N_624,In_238,In_371);
nand U625 (N_625,In_47,In_359);
or U626 (N_626,In_193,In_327);
and U627 (N_627,In_101,In_199);
or U628 (N_628,In_60,In_179);
or U629 (N_629,In_355,In_109);
xnor U630 (N_630,In_420,In_351);
nand U631 (N_631,In_347,In_256);
and U632 (N_632,In_485,In_460);
or U633 (N_633,In_51,In_60);
nand U634 (N_634,In_397,In_139);
nor U635 (N_635,In_280,In_268);
or U636 (N_636,In_406,In_265);
nor U637 (N_637,In_207,In_140);
nor U638 (N_638,In_47,In_173);
nor U639 (N_639,In_35,In_47);
nor U640 (N_640,In_487,In_389);
nand U641 (N_641,In_148,In_96);
nand U642 (N_642,In_36,In_398);
nand U643 (N_643,In_477,In_24);
and U644 (N_644,In_270,In_37);
and U645 (N_645,In_412,In_334);
and U646 (N_646,In_247,In_155);
or U647 (N_647,In_495,In_397);
nand U648 (N_648,In_462,In_470);
and U649 (N_649,In_285,In_92);
nor U650 (N_650,In_450,In_8);
and U651 (N_651,In_320,In_225);
nand U652 (N_652,In_243,In_41);
xor U653 (N_653,In_69,In_257);
and U654 (N_654,In_127,In_314);
and U655 (N_655,In_16,In_220);
nand U656 (N_656,In_380,In_382);
and U657 (N_657,In_376,In_288);
nor U658 (N_658,In_89,In_250);
nand U659 (N_659,In_118,In_7);
or U660 (N_660,In_108,In_351);
or U661 (N_661,In_93,In_289);
or U662 (N_662,In_459,In_412);
nor U663 (N_663,In_429,In_413);
and U664 (N_664,In_419,In_98);
and U665 (N_665,In_199,In_196);
nor U666 (N_666,In_160,In_417);
nand U667 (N_667,In_6,In_349);
nor U668 (N_668,In_247,In_458);
or U669 (N_669,In_369,In_404);
nor U670 (N_670,In_495,In_105);
nand U671 (N_671,In_111,In_65);
and U672 (N_672,In_378,In_53);
and U673 (N_673,In_466,In_426);
or U674 (N_674,In_444,In_385);
or U675 (N_675,In_477,In_358);
or U676 (N_676,In_77,In_305);
and U677 (N_677,In_241,In_203);
nor U678 (N_678,In_210,In_42);
or U679 (N_679,In_84,In_407);
or U680 (N_680,In_447,In_223);
or U681 (N_681,In_216,In_13);
nand U682 (N_682,In_148,In_491);
or U683 (N_683,In_166,In_132);
or U684 (N_684,In_137,In_56);
nor U685 (N_685,In_332,In_153);
or U686 (N_686,In_103,In_350);
nor U687 (N_687,In_63,In_440);
and U688 (N_688,In_4,In_438);
nand U689 (N_689,In_35,In_330);
nor U690 (N_690,In_118,In_410);
and U691 (N_691,In_372,In_227);
xor U692 (N_692,In_192,In_93);
nor U693 (N_693,In_298,In_141);
and U694 (N_694,In_485,In_21);
nand U695 (N_695,In_146,In_42);
nor U696 (N_696,In_177,In_243);
nor U697 (N_697,In_60,In_141);
and U698 (N_698,In_421,In_294);
and U699 (N_699,In_54,In_94);
or U700 (N_700,In_53,In_380);
and U701 (N_701,In_64,In_258);
nand U702 (N_702,In_153,In_387);
and U703 (N_703,In_245,In_111);
nand U704 (N_704,In_210,In_245);
nand U705 (N_705,In_327,In_26);
and U706 (N_706,In_496,In_142);
nor U707 (N_707,In_223,In_92);
nor U708 (N_708,In_107,In_79);
or U709 (N_709,In_61,In_352);
nor U710 (N_710,In_104,In_70);
nor U711 (N_711,In_34,In_336);
nand U712 (N_712,In_244,In_34);
nor U713 (N_713,In_70,In_445);
nor U714 (N_714,In_457,In_11);
or U715 (N_715,In_79,In_101);
nor U716 (N_716,In_124,In_496);
nor U717 (N_717,In_268,In_380);
nand U718 (N_718,In_300,In_320);
xnor U719 (N_719,In_436,In_179);
and U720 (N_720,In_100,In_414);
nand U721 (N_721,In_173,In_164);
or U722 (N_722,In_143,In_391);
nand U723 (N_723,In_310,In_144);
nand U724 (N_724,In_79,In_396);
xnor U725 (N_725,In_173,In_357);
nand U726 (N_726,In_89,In_39);
or U727 (N_727,In_354,In_85);
or U728 (N_728,In_347,In_103);
or U729 (N_729,In_261,In_359);
or U730 (N_730,In_395,In_260);
nor U731 (N_731,In_201,In_308);
or U732 (N_732,In_311,In_379);
and U733 (N_733,In_218,In_223);
nand U734 (N_734,In_305,In_135);
or U735 (N_735,In_411,In_359);
or U736 (N_736,In_485,In_408);
nand U737 (N_737,In_407,In_347);
or U738 (N_738,In_397,In_0);
and U739 (N_739,In_421,In_454);
nand U740 (N_740,In_437,In_47);
nor U741 (N_741,In_385,In_302);
nor U742 (N_742,In_324,In_290);
nand U743 (N_743,In_464,In_11);
xnor U744 (N_744,In_467,In_158);
xnor U745 (N_745,In_145,In_335);
or U746 (N_746,In_91,In_177);
or U747 (N_747,In_375,In_37);
xnor U748 (N_748,In_348,In_53);
or U749 (N_749,In_369,In_201);
and U750 (N_750,In_235,In_219);
nand U751 (N_751,In_240,In_25);
nor U752 (N_752,In_321,In_170);
nor U753 (N_753,In_146,In_117);
xnor U754 (N_754,In_354,In_319);
xor U755 (N_755,In_475,In_281);
nand U756 (N_756,In_172,In_445);
xor U757 (N_757,In_215,In_282);
nand U758 (N_758,In_229,In_50);
nor U759 (N_759,In_83,In_219);
and U760 (N_760,In_249,In_344);
nand U761 (N_761,In_43,In_491);
or U762 (N_762,In_58,In_156);
nor U763 (N_763,In_137,In_163);
nor U764 (N_764,In_285,In_463);
nand U765 (N_765,In_278,In_201);
or U766 (N_766,In_358,In_57);
nor U767 (N_767,In_224,In_480);
and U768 (N_768,In_305,In_390);
nand U769 (N_769,In_128,In_457);
and U770 (N_770,In_24,In_204);
and U771 (N_771,In_45,In_325);
nor U772 (N_772,In_137,In_446);
nand U773 (N_773,In_212,In_316);
or U774 (N_774,In_95,In_57);
nor U775 (N_775,In_263,In_325);
nor U776 (N_776,In_240,In_208);
nor U777 (N_777,In_346,In_194);
and U778 (N_778,In_78,In_391);
nor U779 (N_779,In_471,In_51);
and U780 (N_780,In_463,In_429);
xor U781 (N_781,In_263,In_419);
nand U782 (N_782,In_348,In_221);
or U783 (N_783,In_205,In_455);
or U784 (N_784,In_154,In_391);
nand U785 (N_785,In_323,In_189);
or U786 (N_786,In_103,In_484);
and U787 (N_787,In_1,In_2);
and U788 (N_788,In_282,In_150);
nor U789 (N_789,In_143,In_496);
and U790 (N_790,In_275,In_78);
nand U791 (N_791,In_159,In_182);
nand U792 (N_792,In_245,In_308);
or U793 (N_793,In_307,In_140);
nor U794 (N_794,In_87,In_166);
nand U795 (N_795,In_150,In_271);
nand U796 (N_796,In_493,In_170);
or U797 (N_797,In_426,In_102);
xnor U798 (N_798,In_363,In_442);
xor U799 (N_799,In_323,In_96);
and U800 (N_800,In_91,In_363);
or U801 (N_801,In_69,In_318);
or U802 (N_802,In_312,In_326);
nand U803 (N_803,In_225,In_365);
xor U804 (N_804,In_108,In_245);
nor U805 (N_805,In_95,In_279);
nor U806 (N_806,In_370,In_387);
nor U807 (N_807,In_466,In_92);
nand U808 (N_808,In_45,In_286);
and U809 (N_809,In_479,In_325);
and U810 (N_810,In_332,In_93);
xor U811 (N_811,In_115,In_257);
nor U812 (N_812,In_176,In_54);
and U813 (N_813,In_0,In_463);
nor U814 (N_814,In_404,In_465);
and U815 (N_815,In_431,In_174);
and U816 (N_816,In_388,In_420);
nor U817 (N_817,In_110,In_252);
and U818 (N_818,In_334,In_93);
nor U819 (N_819,In_396,In_210);
and U820 (N_820,In_19,In_354);
or U821 (N_821,In_417,In_355);
or U822 (N_822,In_83,In_121);
nand U823 (N_823,In_321,In_380);
and U824 (N_824,In_145,In_64);
nor U825 (N_825,In_170,In_264);
nor U826 (N_826,In_10,In_429);
or U827 (N_827,In_184,In_409);
or U828 (N_828,In_131,In_319);
nand U829 (N_829,In_407,In_450);
or U830 (N_830,In_427,In_241);
or U831 (N_831,In_103,In_21);
or U832 (N_832,In_393,In_230);
nand U833 (N_833,In_467,In_154);
nor U834 (N_834,In_441,In_103);
or U835 (N_835,In_423,In_273);
nand U836 (N_836,In_12,In_493);
nor U837 (N_837,In_174,In_158);
nor U838 (N_838,In_96,In_58);
or U839 (N_839,In_347,In_140);
nor U840 (N_840,In_455,In_216);
nand U841 (N_841,In_40,In_196);
or U842 (N_842,In_195,In_59);
nand U843 (N_843,In_394,In_53);
and U844 (N_844,In_403,In_221);
or U845 (N_845,In_475,In_39);
nand U846 (N_846,In_410,In_498);
and U847 (N_847,In_481,In_363);
nor U848 (N_848,In_202,In_298);
nand U849 (N_849,In_254,In_103);
and U850 (N_850,In_458,In_121);
nor U851 (N_851,In_446,In_283);
xnor U852 (N_852,In_327,In_450);
nand U853 (N_853,In_252,In_185);
and U854 (N_854,In_137,In_34);
and U855 (N_855,In_423,In_123);
or U856 (N_856,In_224,In_153);
or U857 (N_857,In_6,In_204);
nand U858 (N_858,In_186,In_338);
or U859 (N_859,In_84,In_222);
or U860 (N_860,In_60,In_21);
nand U861 (N_861,In_423,In_96);
and U862 (N_862,In_47,In_372);
nor U863 (N_863,In_88,In_450);
or U864 (N_864,In_156,In_42);
and U865 (N_865,In_491,In_263);
xor U866 (N_866,In_280,In_495);
and U867 (N_867,In_396,In_170);
nand U868 (N_868,In_331,In_335);
and U869 (N_869,In_364,In_491);
or U870 (N_870,In_136,In_338);
nand U871 (N_871,In_394,In_422);
or U872 (N_872,In_420,In_201);
nor U873 (N_873,In_72,In_123);
or U874 (N_874,In_229,In_100);
and U875 (N_875,In_210,In_160);
nor U876 (N_876,In_365,In_103);
nor U877 (N_877,In_482,In_320);
or U878 (N_878,In_411,In_366);
nand U879 (N_879,In_403,In_256);
nor U880 (N_880,In_380,In_320);
and U881 (N_881,In_298,In_392);
nand U882 (N_882,In_357,In_195);
nor U883 (N_883,In_255,In_422);
or U884 (N_884,In_455,In_217);
xor U885 (N_885,In_162,In_315);
or U886 (N_886,In_181,In_385);
and U887 (N_887,In_83,In_311);
nor U888 (N_888,In_429,In_274);
or U889 (N_889,In_299,In_15);
nand U890 (N_890,In_257,In_204);
and U891 (N_891,In_59,In_302);
nand U892 (N_892,In_14,In_69);
xor U893 (N_893,In_474,In_411);
and U894 (N_894,In_226,In_109);
or U895 (N_895,In_120,In_345);
nor U896 (N_896,In_188,In_331);
nand U897 (N_897,In_279,In_55);
and U898 (N_898,In_294,In_341);
nor U899 (N_899,In_494,In_348);
nand U900 (N_900,In_274,In_352);
nand U901 (N_901,In_153,In_238);
nor U902 (N_902,In_141,In_34);
xor U903 (N_903,In_41,In_136);
or U904 (N_904,In_135,In_395);
nand U905 (N_905,In_350,In_108);
nor U906 (N_906,In_25,In_155);
nor U907 (N_907,In_14,In_252);
nand U908 (N_908,In_333,In_456);
and U909 (N_909,In_263,In_291);
or U910 (N_910,In_482,In_439);
nor U911 (N_911,In_62,In_352);
and U912 (N_912,In_229,In_405);
nor U913 (N_913,In_122,In_188);
nor U914 (N_914,In_442,In_68);
nor U915 (N_915,In_143,In_277);
nor U916 (N_916,In_111,In_306);
nor U917 (N_917,In_220,In_190);
nor U918 (N_918,In_247,In_215);
nor U919 (N_919,In_344,In_274);
or U920 (N_920,In_359,In_192);
nor U921 (N_921,In_363,In_482);
or U922 (N_922,In_498,In_154);
nor U923 (N_923,In_229,In_208);
and U924 (N_924,In_304,In_453);
and U925 (N_925,In_30,In_443);
or U926 (N_926,In_250,In_139);
or U927 (N_927,In_263,In_197);
nand U928 (N_928,In_451,In_195);
or U929 (N_929,In_281,In_122);
and U930 (N_930,In_468,In_430);
or U931 (N_931,In_209,In_410);
nand U932 (N_932,In_267,In_90);
and U933 (N_933,In_387,In_165);
or U934 (N_934,In_224,In_457);
or U935 (N_935,In_44,In_321);
nor U936 (N_936,In_360,In_224);
nor U937 (N_937,In_64,In_38);
nand U938 (N_938,In_299,In_443);
nand U939 (N_939,In_434,In_201);
and U940 (N_940,In_169,In_456);
nor U941 (N_941,In_286,In_264);
nor U942 (N_942,In_373,In_57);
or U943 (N_943,In_222,In_361);
nor U944 (N_944,In_86,In_309);
or U945 (N_945,In_299,In_161);
and U946 (N_946,In_297,In_22);
and U947 (N_947,In_75,In_222);
and U948 (N_948,In_434,In_116);
nand U949 (N_949,In_271,In_199);
nand U950 (N_950,In_53,In_267);
or U951 (N_951,In_326,In_123);
nand U952 (N_952,In_193,In_482);
and U953 (N_953,In_359,In_78);
and U954 (N_954,In_421,In_190);
or U955 (N_955,In_225,In_181);
nand U956 (N_956,In_496,In_413);
nor U957 (N_957,In_419,In_167);
nand U958 (N_958,In_59,In_58);
nand U959 (N_959,In_458,In_109);
nand U960 (N_960,In_23,In_86);
nor U961 (N_961,In_136,In_438);
or U962 (N_962,In_425,In_76);
or U963 (N_963,In_203,In_331);
or U964 (N_964,In_325,In_320);
and U965 (N_965,In_493,In_468);
or U966 (N_966,In_206,In_240);
and U967 (N_967,In_80,In_477);
nor U968 (N_968,In_270,In_379);
or U969 (N_969,In_294,In_270);
nand U970 (N_970,In_53,In_411);
nand U971 (N_971,In_308,In_408);
or U972 (N_972,In_37,In_72);
nand U973 (N_973,In_136,In_286);
and U974 (N_974,In_40,In_427);
and U975 (N_975,In_393,In_235);
or U976 (N_976,In_9,In_258);
nand U977 (N_977,In_121,In_305);
or U978 (N_978,In_275,In_416);
and U979 (N_979,In_182,In_109);
nor U980 (N_980,In_197,In_252);
nand U981 (N_981,In_36,In_409);
nor U982 (N_982,In_327,In_270);
and U983 (N_983,In_182,In_27);
or U984 (N_984,In_476,In_373);
and U985 (N_985,In_240,In_384);
nand U986 (N_986,In_35,In_181);
and U987 (N_987,In_92,In_350);
nand U988 (N_988,In_94,In_98);
or U989 (N_989,In_244,In_182);
and U990 (N_990,In_5,In_470);
or U991 (N_991,In_128,In_274);
or U992 (N_992,In_341,In_126);
nand U993 (N_993,In_413,In_111);
and U994 (N_994,In_35,In_300);
and U995 (N_995,In_196,In_424);
nand U996 (N_996,In_238,In_430);
nor U997 (N_997,In_265,In_304);
or U998 (N_998,In_141,In_228);
and U999 (N_999,In_236,In_52);
or U1000 (N_1000,N_846,N_519);
nor U1001 (N_1001,N_243,N_408);
and U1002 (N_1002,N_432,N_495);
nor U1003 (N_1003,N_740,N_518);
or U1004 (N_1004,N_636,N_264);
nand U1005 (N_1005,N_657,N_553);
nor U1006 (N_1006,N_650,N_308);
xnor U1007 (N_1007,N_952,N_763);
or U1008 (N_1008,N_725,N_119);
or U1009 (N_1009,N_444,N_560);
nand U1010 (N_1010,N_602,N_307);
and U1011 (N_1011,N_460,N_809);
or U1012 (N_1012,N_780,N_434);
and U1013 (N_1013,N_411,N_224);
or U1014 (N_1014,N_765,N_153);
or U1015 (N_1015,N_915,N_821);
or U1016 (N_1016,N_754,N_72);
nor U1017 (N_1017,N_849,N_394);
nor U1018 (N_1018,N_808,N_668);
nor U1019 (N_1019,N_59,N_700);
xnor U1020 (N_1020,N_175,N_615);
nor U1021 (N_1021,N_859,N_940);
and U1022 (N_1022,N_907,N_572);
nand U1023 (N_1023,N_274,N_909);
nor U1024 (N_1024,N_240,N_222);
nor U1025 (N_1025,N_208,N_608);
or U1026 (N_1026,N_166,N_866);
and U1027 (N_1027,N_894,N_82);
and U1028 (N_1028,N_68,N_674);
and U1029 (N_1029,N_450,N_750);
nand U1030 (N_1030,N_397,N_664);
nand U1031 (N_1031,N_491,N_928);
and U1032 (N_1032,N_498,N_488);
or U1033 (N_1033,N_832,N_283);
nor U1034 (N_1034,N_351,N_246);
or U1035 (N_1035,N_178,N_600);
nand U1036 (N_1036,N_922,N_764);
or U1037 (N_1037,N_338,N_681);
or U1038 (N_1038,N_298,N_417);
and U1039 (N_1039,N_36,N_237);
nor U1040 (N_1040,N_862,N_94);
nand U1041 (N_1041,N_269,N_516);
or U1042 (N_1042,N_704,N_624);
or U1043 (N_1043,N_333,N_261);
nor U1044 (N_1044,N_113,N_289);
nand U1045 (N_1045,N_115,N_556);
nand U1046 (N_1046,N_1,N_935);
nand U1047 (N_1047,N_638,N_379);
or U1048 (N_1048,N_996,N_21);
nand U1049 (N_1049,N_100,N_597);
or U1050 (N_1050,N_86,N_167);
nor U1051 (N_1051,N_235,N_229);
nand U1052 (N_1052,N_402,N_496);
nand U1053 (N_1053,N_447,N_574);
and U1054 (N_1054,N_457,N_469);
nand U1055 (N_1055,N_471,N_304);
nor U1056 (N_1056,N_232,N_67);
nor U1057 (N_1057,N_456,N_771);
nor U1058 (N_1058,N_876,N_651);
or U1059 (N_1059,N_212,N_554);
xor U1060 (N_1060,N_284,N_843);
and U1061 (N_1061,N_248,N_79);
nor U1062 (N_1062,N_288,N_489);
nor U1063 (N_1063,N_135,N_173);
or U1064 (N_1064,N_58,N_218);
nand U1065 (N_1065,N_938,N_33);
nor U1066 (N_1066,N_181,N_238);
or U1067 (N_1067,N_661,N_586);
nand U1068 (N_1068,N_815,N_873);
and U1069 (N_1069,N_576,N_155);
nand U1070 (N_1070,N_392,N_623);
nand U1071 (N_1071,N_705,N_901);
or U1072 (N_1072,N_864,N_943);
or U1073 (N_1073,N_699,N_850);
and U1074 (N_1074,N_865,N_634);
nand U1075 (N_1075,N_893,N_227);
nand U1076 (N_1076,N_202,N_92);
and U1077 (N_1077,N_327,N_453);
or U1078 (N_1078,N_716,N_570);
nor U1079 (N_1079,N_415,N_340);
nand U1080 (N_1080,N_861,N_287);
nor U1081 (N_1081,N_326,N_622);
and U1082 (N_1082,N_975,N_695);
nor U1083 (N_1083,N_344,N_937);
and U1084 (N_1084,N_449,N_913);
nor U1085 (N_1085,N_116,N_39);
nand U1086 (N_1086,N_689,N_256);
nor U1087 (N_1087,N_69,N_799);
or U1088 (N_1088,N_215,N_603);
nor U1089 (N_1089,N_31,N_561);
nand U1090 (N_1090,N_347,N_573);
or U1091 (N_1091,N_803,N_370);
nand U1092 (N_1092,N_384,N_688);
and U1093 (N_1093,N_52,N_881);
nand U1094 (N_1094,N_512,N_328);
or U1095 (N_1095,N_663,N_900);
nor U1096 (N_1096,N_34,N_852);
nor U1097 (N_1097,N_366,N_2);
and U1098 (N_1098,N_748,N_766);
nand U1099 (N_1099,N_321,N_376);
nor U1100 (N_1100,N_840,N_823);
nor U1101 (N_1101,N_65,N_300);
nor U1102 (N_1102,N_487,N_522);
and U1103 (N_1103,N_25,N_436);
nor U1104 (N_1104,N_422,N_412);
xnor U1105 (N_1105,N_168,N_12);
nor U1106 (N_1106,N_867,N_587);
or U1107 (N_1107,N_182,N_233);
nor U1108 (N_1108,N_761,N_680);
nor U1109 (N_1109,N_474,N_929);
or U1110 (N_1110,N_584,N_589);
or U1111 (N_1111,N_446,N_293);
and U1112 (N_1112,N_606,N_851);
or U1113 (N_1113,N_738,N_197);
nand U1114 (N_1114,N_787,N_57);
or U1115 (N_1115,N_118,N_784);
and U1116 (N_1116,N_410,N_981);
and U1117 (N_1117,N_942,N_545);
and U1118 (N_1118,N_965,N_102);
or U1119 (N_1119,N_953,N_160);
nor U1120 (N_1120,N_962,N_713);
or U1121 (N_1121,N_280,N_869);
and U1122 (N_1122,N_140,N_426);
and U1123 (N_1123,N_797,N_656);
xnor U1124 (N_1124,N_993,N_42);
nor U1125 (N_1125,N_386,N_985);
and U1126 (N_1126,N_789,N_563);
nor U1127 (N_1127,N_322,N_466);
nand U1128 (N_1128,N_180,N_895);
or U1129 (N_1129,N_273,N_336);
and U1130 (N_1130,N_473,N_236);
or U1131 (N_1131,N_54,N_106);
or U1132 (N_1132,N_593,N_908);
nor U1133 (N_1133,N_997,N_87);
and U1134 (N_1134,N_348,N_970);
nand U1135 (N_1135,N_101,N_921);
or U1136 (N_1136,N_37,N_147);
and U1137 (N_1137,N_27,N_226);
and U1138 (N_1138,N_632,N_254);
nor U1139 (N_1139,N_192,N_275);
nand U1140 (N_1140,N_369,N_477);
nor U1141 (N_1141,N_501,N_999);
and U1142 (N_1142,N_626,N_209);
nand U1143 (N_1143,N_188,N_198);
nor U1144 (N_1144,N_22,N_837);
nand U1145 (N_1145,N_196,N_958);
and U1146 (N_1146,N_398,N_744);
or U1147 (N_1147,N_125,N_992);
or U1148 (N_1148,N_978,N_637);
nor U1149 (N_1149,N_64,N_737);
and U1150 (N_1150,N_319,N_159);
nand U1151 (N_1151,N_162,N_241);
or U1152 (N_1152,N_442,N_482);
and U1153 (N_1153,N_80,N_391);
and U1154 (N_1154,N_524,N_10);
nand U1155 (N_1155,N_774,N_559);
nor U1156 (N_1156,N_15,N_4);
and U1157 (N_1157,N_550,N_874);
and U1158 (N_1158,N_85,N_355);
nor U1159 (N_1159,N_372,N_189);
nor U1160 (N_1160,N_891,N_431);
nand U1161 (N_1161,N_219,N_99);
or U1162 (N_1162,N_790,N_914);
nor U1163 (N_1163,N_123,N_295);
nand U1164 (N_1164,N_174,N_423);
nor U1165 (N_1165,N_380,N_131);
and U1166 (N_1166,N_715,N_834);
nor U1167 (N_1167,N_898,N_373);
nand U1168 (N_1168,N_918,N_381);
or U1169 (N_1169,N_210,N_506);
or U1170 (N_1170,N_360,N_647);
nand U1171 (N_1171,N_510,N_731);
and U1172 (N_1172,N_536,N_49);
nor U1173 (N_1173,N_30,N_217);
and U1174 (N_1174,N_714,N_8);
nor U1175 (N_1175,N_521,N_961);
or U1176 (N_1176,N_762,N_11);
nand U1177 (N_1177,N_537,N_598);
xor U1178 (N_1178,N_591,N_503);
nor U1179 (N_1179,N_389,N_788);
nand U1180 (N_1180,N_826,N_368);
or U1181 (N_1181,N_3,N_403);
nand U1182 (N_1182,N_919,N_204);
or U1183 (N_1183,N_730,N_927);
and U1184 (N_1184,N_126,N_438);
or U1185 (N_1185,N_378,N_323);
nand U1186 (N_1186,N_706,N_9);
and U1187 (N_1187,N_547,N_991);
or U1188 (N_1188,N_562,N_467);
or U1189 (N_1189,N_16,N_583);
or U1190 (N_1190,N_614,N_708);
xor U1191 (N_1191,N_599,N_461);
nand U1192 (N_1192,N_811,N_805);
nand U1193 (N_1193,N_183,N_980);
nor U1194 (N_1194,N_47,N_6);
or U1195 (N_1195,N_694,N_413);
or U1196 (N_1196,N_427,N_430);
nand U1197 (N_1197,N_455,N_483);
and U1198 (N_1198,N_653,N_546);
nand U1199 (N_1199,N_393,N_697);
or U1200 (N_1200,N_205,N_356);
nand U1201 (N_1201,N_542,N_76);
nor U1202 (N_1202,N_200,N_783);
or U1203 (N_1203,N_353,N_282);
and U1204 (N_1204,N_569,N_267);
and U1205 (N_1205,N_858,N_833);
or U1206 (N_1206,N_676,N_649);
and U1207 (N_1207,N_769,N_549);
nor U1208 (N_1208,N_409,N_244);
nor U1209 (N_1209,N_310,N_646);
or U1210 (N_1210,N_825,N_625);
nor U1211 (N_1211,N_829,N_499);
and U1212 (N_1212,N_374,N_459);
and U1213 (N_1213,N_964,N_818);
nand U1214 (N_1214,N_605,N_151);
or U1215 (N_1215,N_48,N_214);
and U1216 (N_1216,N_145,N_74);
nand U1217 (N_1217,N_0,N_617);
and U1218 (N_1218,N_231,N_324);
nor U1219 (N_1219,N_485,N_946);
or U1220 (N_1220,N_306,N_643);
or U1221 (N_1221,N_984,N_303);
nor U1222 (N_1222,N_702,N_296);
or U1223 (N_1223,N_136,N_828);
nor U1224 (N_1224,N_581,N_130);
nand U1225 (N_1225,N_252,N_741);
or U1226 (N_1226,N_627,N_749);
or U1227 (N_1227,N_251,N_419);
nor U1228 (N_1228,N_523,N_358);
and U1229 (N_1229,N_95,N_899);
and U1230 (N_1230,N_601,N_870);
and U1231 (N_1231,N_290,N_590);
nand U1232 (N_1232,N_880,N_77);
or U1233 (N_1233,N_314,N_673);
nand U1234 (N_1234,N_170,N_19);
or U1235 (N_1235,N_971,N_81);
and U1236 (N_1236,N_493,N_317);
nor U1237 (N_1237,N_262,N_242);
nor U1238 (N_1238,N_635,N_791);
or U1239 (N_1239,N_558,N_195);
and U1240 (N_1240,N_539,N_332);
xor U1241 (N_1241,N_448,N_968);
or U1242 (N_1242,N_257,N_966);
nand U1243 (N_1243,N_936,N_350);
and U1244 (N_1244,N_732,N_352);
and U1245 (N_1245,N_110,N_944);
and U1246 (N_1246,N_451,N_365);
nand U1247 (N_1247,N_916,N_278);
and U1248 (N_1248,N_223,N_396);
or U1249 (N_1249,N_759,N_247);
or U1250 (N_1250,N_728,N_13);
nand U1251 (N_1251,N_988,N_190);
or U1252 (N_1252,N_810,N_470);
or U1253 (N_1253,N_472,N_50);
and U1254 (N_1254,N_594,N_777);
nand U1255 (N_1255,N_817,N_579);
nand U1256 (N_1256,N_806,N_390);
or U1257 (N_1257,N_973,N_112);
nand U1258 (N_1258,N_107,N_756);
nor U1259 (N_1259,N_860,N_529);
nand U1260 (N_1260,N_7,N_475);
nor U1261 (N_1261,N_954,N_185);
nand U1262 (N_1262,N_41,N_266);
or U1263 (N_1263,N_781,N_729);
or U1264 (N_1264,N_193,N_727);
and U1265 (N_1265,N_611,N_575);
nand U1266 (N_1266,N_747,N_671);
nand U1267 (N_1267,N_685,N_526);
and U1268 (N_1268,N_724,N_629);
nor U1269 (N_1269,N_525,N_709);
and U1270 (N_1270,N_710,N_320);
nor U1271 (N_1271,N_565,N_270);
and U1272 (N_1272,N_755,N_230);
or U1273 (N_1273,N_819,N_464);
or U1274 (N_1274,N_479,N_429);
nor U1275 (N_1275,N_630,N_211);
or U1276 (N_1276,N_620,N_665);
or U1277 (N_1277,N_703,N_201);
nor U1278 (N_1278,N_62,N_122);
nand U1279 (N_1279,N_105,N_903);
and U1280 (N_1280,N_842,N_800);
and U1281 (N_1281,N_655,N_281);
and U1282 (N_1282,N_543,N_845);
and U1283 (N_1283,N_5,N_585);
or U1284 (N_1284,N_88,N_707);
or U1285 (N_1285,N_97,N_930);
nand U1286 (N_1286,N_844,N_712);
and U1287 (N_1287,N_607,N_399);
nand U1288 (N_1288,N_103,N_772);
and U1289 (N_1289,N_640,N_920);
nor U1290 (N_1290,N_207,N_794);
or U1291 (N_1291,N_20,N_141);
and U1292 (N_1292,N_154,N_481);
and U1293 (N_1293,N_316,N_443);
nor U1294 (N_1294,N_802,N_70);
or U1295 (N_1295,N_268,N_588);
nand U1296 (N_1296,N_385,N_568);
xor U1297 (N_1297,N_362,N_854);
or U1298 (N_1298,N_566,N_187);
nand U1299 (N_1299,N_249,N_150);
nor U1300 (N_1300,N_63,N_437);
and U1301 (N_1301,N_677,N_445);
and U1302 (N_1302,N_172,N_824);
or U1303 (N_1303,N_633,N_28);
nand U1304 (N_1304,N_814,N_142);
and U1305 (N_1305,N_779,N_877);
or U1306 (N_1306,N_425,N_302);
or U1307 (N_1307,N_986,N_511);
nand U1308 (N_1308,N_691,N_14);
nor U1309 (N_1309,N_294,N_675);
or U1310 (N_1310,N_186,N_149);
and U1311 (N_1311,N_478,N_923);
nor U1312 (N_1312,N_619,N_813);
or U1313 (N_1313,N_698,N_171);
and U1314 (N_1314,N_114,N_692);
nor U1315 (N_1315,N_311,N_129);
nor U1316 (N_1316,N_158,N_841);
or U1317 (N_1317,N_330,N_830);
nand U1318 (N_1318,N_902,N_341);
nor U1319 (N_1319,N_795,N_742);
nand U1320 (N_1320,N_441,N_642);
or U1321 (N_1321,N_305,N_505);
or U1322 (N_1322,N_299,N_371);
and U1323 (N_1323,N_335,N_216);
nand U1324 (N_1324,N_276,N_904);
and U1325 (N_1325,N_648,N_367);
or U1326 (N_1326,N_260,N_990);
or U1327 (N_1327,N_345,N_947);
nor U1328 (N_1328,N_253,N_773);
nand U1329 (N_1329,N_956,N_959);
and U1330 (N_1330,N_83,N_812);
nor U1331 (N_1331,N_279,N_465);
nand U1332 (N_1332,N_743,N_977);
and U1333 (N_1333,N_517,N_361);
nor U1334 (N_1334,N_234,N_339);
and U1335 (N_1335,N_124,N_592);
and U1336 (N_1336,N_343,N_654);
nor U1337 (N_1337,N_73,N_334);
or U1338 (N_1338,N_882,N_363);
or U1339 (N_1339,N_428,N_169);
nor U1340 (N_1340,N_911,N_857);
or U1341 (N_1341,N_683,N_711);
and U1342 (N_1342,N_796,N_871);
nand U1343 (N_1343,N_492,N_272);
or U1344 (N_1344,N_931,N_838);
nor U1345 (N_1345,N_520,N_509);
nand U1346 (N_1346,N_312,N_721);
or U1347 (N_1347,N_17,N_906);
or U1348 (N_1348,N_515,N_133);
or U1349 (N_1349,N_604,N_382);
nand U1350 (N_1350,N_872,N_435);
and U1351 (N_1351,N_687,N_404);
or U1352 (N_1352,N_60,N_255);
or U1353 (N_1353,N_258,N_46);
nand U1354 (N_1354,N_701,N_177);
nor U1355 (N_1355,N_645,N_785);
nand U1356 (N_1356,N_421,N_497);
or U1357 (N_1357,N_801,N_476);
and U1358 (N_1358,N_152,N_945);
or U1359 (N_1359,N_78,N_291);
nor U1360 (N_1360,N_134,N_40);
nor U1361 (N_1361,N_760,N_24);
or U1362 (N_1362,N_318,N_164);
or U1363 (N_1363,N_400,N_315);
and U1364 (N_1364,N_782,N_108);
nor U1365 (N_1365,N_420,N_357);
or U1366 (N_1366,N_804,N_631);
or U1367 (N_1367,N_395,N_121);
xor U1368 (N_1368,N_84,N_979);
or U1369 (N_1369,N_199,N_61);
nand U1370 (N_1370,N_504,N_416);
nand U1371 (N_1371,N_179,N_96);
nand U1372 (N_1372,N_191,N_679);
or U1373 (N_1373,N_669,N_406);
nand U1374 (N_1374,N_486,N_337);
nand U1375 (N_1375,N_342,N_452);
nor U1376 (N_1376,N_736,N_822);
or U1377 (N_1377,N_758,N_723);
or U1378 (N_1378,N_331,N_245);
or U1379 (N_1379,N_165,N_745);
nand U1380 (N_1380,N_955,N_735);
nor U1381 (N_1381,N_949,N_890);
or U1382 (N_1382,N_746,N_271);
or U1383 (N_1383,N_387,N_53);
nand U1384 (N_1384,N_535,N_690);
nor U1385 (N_1385,N_93,N_527);
nand U1386 (N_1386,N_856,N_836);
and U1387 (N_1387,N_91,N_879);
and U1388 (N_1388,N_847,N_109);
nor U1389 (N_1389,N_578,N_939);
and U1390 (N_1390,N_839,N_56);
and U1391 (N_1391,N_577,N_816);
nand U1392 (N_1392,N_888,N_567);
or U1393 (N_1393,N_51,N_484);
or U1394 (N_1394,N_286,N_621);
nand U1395 (N_1395,N_994,N_983);
nand U1396 (N_1396,N_644,N_827);
or U1397 (N_1397,N_490,N_544);
or U1398 (N_1398,N_552,N_309);
nor U1399 (N_1399,N_184,N_739);
xor U1400 (N_1400,N_684,N_250);
or U1401 (N_1401,N_807,N_995);
nand U1402 (N_1402,N_752,N_424);
nor U1403 (N_1403,N_375,N_127);
nor U1404 (N_1404,N_146,N_221);
or U1405 (N_1405,N_662,N_555);
and U1406 (N_1406,N_383,N_462);
or U1407 (N_1407,N_138,N_767);
or U1408 (N_1408,N_329,N_98);
and U1409 (N_1409,N_494,N_228);
nor U1410 (N_1410,N_757,N_407);
or U1411 (N_1411,N_530,N_557);
nand U1412 (N_1412,N_660,N_719);
and U1413 (N_1413,N_144,N_696);
nand U1414 (N_1414,N_855,N_848);
or U1415 (N_1415,N_682,N_941);
nor U1416 (N_1416,N_957,N_433);
or U1417 (N_1417,N_540,N_932);
xor U1418 (N_1418,N_71,N_770);
nand U1419 (N_1419,N_718,N_458);
nor U1420 (N_1420,N_66,N_292);
nand U1421 (N_1421,N_439,N_974);
nor U1422 (N_1422,N_658,N_18);
or U1423 (N_1423,N_143,N_117);
and U1424 (N_1424,N_157,N_910);
and U1425 (N_1425,N_925,N_831);
and U1426 (N_1426,N_89,N_502);
nand U1427 (N_1427,N_533,N_26);
or U1428 (N_1428,N_969,N_868);
nor U1429 (N_1429,N_889,N_951);
and U1430 (N_1430,N_693,N_377);
and U1431 (N_1431,N_998,N_551);
nand U1432 (N_1432,N_354,N_285);
nand U1433 (N_1433,N_43,N_595);
and U1434 (N_1434,N_641,N_414);
nand U1435 (N_1435,N_686,N_775);
nor U1436 (N_1436,N_161,N_440);
nand U1437 (N_1437,N_878,N_912);
or U1438 (N_1438,N_44,N_297);
or U1439 (N_1439,N_513,N_618);
and U1440 (N_1440,N_156,N_531);
or U1441 (N_1441,N_564,N_726);
and U1442 (N_1442,N_853,N_753);
nor U1443 (N_1443,N_778,N_480);
or U1444 (N_1444,N_38,N_596);
nand U1445 (N_1445,N_950,N_672);
nor U1446 (N_1446,N_885,N_960);
nand U1447 (N_1447,N_733,N_137);
or U1448 (N_1448,N_265,N_734);
nor U1449 (N_1449,N_532,N_548);
and U1450 (N_1450,N_917,N_768);
nand U1451 (N_1451,N_132,N_933);
or U1452 (N_1452,N_325,N_32);
or U1453 (N_1453,N_239,N_792);
and U1454 (N_1454,N_659,N_666);
nor U1455 (N_1455,N_616,N_793);
nor U1456 (N_1456,N_454,N_786);
or U1457 (N_1457,N_987,N_163);
and U1458 (N_1458,N_90,N_405);
or U1459 (N_1459,N_628,N_982);
and U1460 (N_1460,N_905,N_364);
nor U1461 (N_1461,N_508,N_887);
or U1462 (N_1462,N_963,N_301);
nand U1463 (N_1463,N_976,N_875);
nand U1464 (N_1464,N_111,N_948);
nand U1465 (N_1465,N_538,N_139);
nand U1466 (N_1466,N_798,N_776);
and U1467 (N_1467,N_259,N_213);
nand U1468 (N_1468,N_401,N_206);
nor U1469 (N_1469,N_967,N_897);
nor U1470 (N_1470,N_717,N_104);
and U1471 (N_1471,N_883,N_580);
nand U1472 (N_1472,N_388,N_896);
nand U1473 (N_1473,N_176,N_652);
nand U1474 (N_1474,N_120,N_720);
or U1475 (N_1475,N_751,N_934);
and U1476 (N_1476,N_612,N_468);
and U1477 (N_1477,N_835,N_55);
nor U1478 (N_1478,N_514,N_972);
xor U1479 (N_1479,N_884,N_892);
and U1480 (N_1480,N_75,N_678);
and U1481 (N_1481,N_528,N_639);
or U1482 (N_1482,N_610,N_541);
nor U1483 (N_1483,N_194,N_507);
nand U1484 (N_1484,N_609,N_263);
and U1485 (N_1485,N_722,N_23);
and U1486 (N_1486,N_989,N_500);
nand U1487 (N_1487,N_820,N_277);
or U1488 (N_1488,N_148,N_220);
or U1489 (N_1489,N_346,N_926);
nand U1490 (N_1490,N_313,N_667);
nor U1491 (N_1491,N_463,N_924);
nand U1492 (N_1492,N_45,N_571);
nand U1493 (N_1493,N_225,N_35);
nor U1494 (N_1494,N_670,N_349);
and U1495 (N_1495,N_359,N_863);
nor U1496 (N_1496,N_613,N_128);
nand U1497 (N_1497,N_203,N_534);
and U1498 (N_1498,N_886,N_418);
or U1499 (N_1499,N_582,N_29);
or U1500 (N_1500,N_741,N_523);
or U1501 (N_1501,N_73,N_6);
or U1502 (N_1502,N_589,N_451);
nor U1503 (N_1503,N_725,N_152);
nor U1504 (N_1504,N_923,N_888);
nor U1505 (N_1505,N_749,N_974);
nand U1506 (N_1506,N_504,N_395);
or U1507 (N_1507,N_537,N_871);
xnor U1508 (N_1508,N_591,N_869);
nand U1509 (N_1509,N_199,N_306);
and U1510 (N_1510,N_158,N_665);
or U1511 (N_1511,N_852,N_780);
and U1512 (N_1512,N_668,N_640);
and U1513 (N_1513,N_258,N_11);
or U1514 (N_1514,N_388,N_532);
nand U1515 (N_1515,N_619,N_507);
or U1516 (N_1516,N_647,N_346);
nor U1517 (N_1517,N_163,N_524);
nor U1518 (N_1518,N_415,N_577);
and U1519 (N_1519,N_536,N_866);
nand U1520 (N_1520,N_978,N_475);
nor U1521 (N_1521,N_352,N_102);
and U1522 (N_1522,N_260,N_488);
or U1523 (N_1523,N_752,N_276);
nand U1524 (N_1524,N_272,N_619);
nor U1525 (N_1525,N_80,N_14);
or U1526 (N_1526,N_419,N_955);
and U1527 (N_1527,N_937,N_857);
or U1528 (N_1528,N_843,N_86);
xnor U1529 (N_1529,N_343,N_775);
and U1530 (N_1530,N_509,N_59);
nor U1531 (N_1531,N_768,N_746);
nand U1532 (N_1532,N_529,N_617);
and U1533 (N_1533,N_156,N_573);
and U1534 (N_1534,N_954,N_179);
and U1535 (N_1535,N_848,N_866);
or U1536 (N_1536,N_693,N_689);
and U1537 (N_1537,N_983,N_39);
or U1538 (N_1538,N_959,N_500);
xnor U1539 (N_1539,N_293,N_442);
and U1540 (N_1540,N_581,N_758);
or U1541 (N_1541,N_893,N_470);
nand U1542 (N_1542,N_437,N_141);
nor U1543 (N_1543,N_566,N_536);
or U1544 (N_1544,N_960,N_110);
xor U1545 (N_1545,N_746,N_5);
or U1546 (N_1546,N_517,N_245);
or U1547 (N_1547,N_628,N_480);
or U1548 (N_1548,N_663,N_285);
and U1549 (N_1549,N_96,N_703);
nor U1550 (N_1550,N_226,N_28);
or U1551 (N_1551,N_417,N_318);
and U1552 (N_1552,N_309,N_432);
nor U1553 (N_1553,N_61,N_64);
nor U1554 (N_1554,N_78,N_674);
nor U1555 (N_1555,N_399,N_843);
and U1556 (N_1556,N_623,N_400);
nand U1557 (N_1557,N_895,N_707);
or U1558 (N_1558,N_863,N_337);
or U1559 (N_1559,N_957,N_891);
or U1560 (N_1560,N_350,N_700);
and U1561 (N_1561,N_427,N_466);
or U1562 (N_1562,N_835,N_554);
and U1563 (N_1563,N_202,N_817);
and U1564 (N_1564,N_263,N_840);
nor U1565 (N_1565,N_50,N_378);
nand U1566 (N_1566,N_422,N_753);
and U1567 (N_1567,N_695,N_270);
and U1568 (N_1568,N_356,N_846);
or U1569 (N_1569,N_852,N_3);
or U1570 (N_1570,N_518,N_617);
nor U1571 (N_1571,N_944,N_192);
xor U1572 (N_1572,N_449,N_930);
nor U1573 (N_1573,N_391,N_279);
nand U1574 (N_1574,N_333,N_820);
or U1575 (N_1575,N_785,N_348);
nor U1576 (N_1576,N_424,N_971);
and U1577 (N_1577,N_866,N_140);
nand U1578 (N_1578,N_239,N_946);
xnor U1579 (N_1579,N_131,N_626);
nand U1580 (N_1580,N_489,N_997);
and U1581 (N_1581,N_288,N_791);
and U1582 (N_1582,N_517,N_301);
or U1583 (N_1583,N_797,N_8);
or U1584 (N_1584,N_369,N_152);
and U1585 (N_1585,N_74,N_719);
nor U1586 (N_1586,N_55,N_810);
nand U1587 (N_1587,N_814,N_309);
nand U1588 (N_1588,N_700,N_470);
xor U1589 (N_1589,N_156,N_273);
nand U1590 (N_1590,N_180,N_875);
nor U1591 (N_1591,N_652,N_211);
or U1592 (N_1592,N_394,N_257);
or U1593 (N_1593,N_541,N_505);
and U1594 (N_1594,N_165,N_161);
and U1595 (N_1595,N_593,N_487);
nor U1596 (N_1596,N_148,N_932);
xnor U1597 (N_1597,N_972,N_741);
or U1598 (N_1598,N_28,N_483);
nand U1599 (N_1599,N_428,N_528);
or U1600 (N_1600,N_482,N_517);
nand U1601 (N_1601,N_680,N_492);
nand U1602 (N_1602,N_406,N_315);
and U1603 (N_1603,N_302,N_669);
and U1604 (N_1604,N_813,N_337);
and U1605 (N_1605,N_10,N_189);
or U1606 (N_1606,N_406,N_15);
and U1607 (N_1607,N_318,N_764);
nand U1608 (N_1608,N_926,N_272);
and U1609 (N_1609,N_667,N_786);
nand U1610 (N_1610,N_923,N_806);
nand U1611 (N_1611,N_936,N_112);
nand U1612 (N_1612,N_613,N_860);
nor U1613 (N_1613,N_820,N_790);
nor U1614 (N_1614,N_662,N_719);
nand U1615 (N_1615,N_148,N_399);
nor U1616 (N_1616,N_687,N_342);
or U1617 (N_1617,N_535,N_443);
and U1618 (N_1618,N_575,N_205);
and U1619 (N_1619,N_217,N_571);
nand U1620 (N_1620,N_592,N_193);
nand U1621 (N_1621,N_899,N_491);
nor U1622 (N_1622,N_477,N_501);
nand U1623 (N_1623,N_691,N_424);
and U1624 (N_1624,N_915,N_132);
and U1625 (N_1625,N_90,N_672);
nand U1626 (N_1626,N_833,N_726);
nand U1627 (N_1627,N_598,N_827);
nor U1628 (N_1628,N_635,N_330);
nor U1629 (N_1629,N_334,N_107);
nor U1630 (N_1630,N_255,N_843);
nor U1631 (N_1631,N_728,N_766);
nor U1632 (N_1632,N_440,N_339);
xor U1633 (N_1633,N_382,N_678);
or U1634 (N_1634,N_216,N_186);
or U1635 (N_1635,N_954,N_257);
nor U1636 (N_1636,N_992,N_419);
nand U1637 (N_1637,N_120,N_905);
nand U1638 (N_1638,N_89,N_683);
nor U1639 (N_1639,N_260,N_10);
and U1640 (N_1640,N_655,N_652);
or U1641 (N_1641,N_316,N_37);
nand U1642 (N_1642,N_783,N_418);
nand U1643 (N_1643,N_916,N_303);
and U1644 (N_1644,N_942,N_289);
xnor U1645 (N_1645,N_71,N_451);
nor U1646 (N_1646,N_545,N_319);
xnor U1647 (N_1647,N_360,N_731);
nor U1648 (N_1648,N_992,N_61);
or U1649 (N_1649,N_307,N_733);
nand U1650 (N_1650,N_461,N_160);
xor U1651 (N_1651,N_781,N_132);
and U1652 (N_1652,N_660,N_446);
nor U1653 (N_1653,N_884,N_43);
nor U1654 (N_1654,N_848,N_530);
or U1655 (N_1655,N_801,N_739);
or U1656 (N_1656,N_433,N_924);
nor U1657 (N_1657,N_137,N_926);
nand U1658 (N_1658,N_505,N_439);
nand U1659 (N_1659,N_556,N_671);
or U1660 (N_1660,N_330,N_275);
and U1661 (N_1661,N_137,N_772);
and U1662 (N_1662,N_471,N_641);
or U1663 (N_1663,N_960,N_482);
nand U1664 (N_1664,N_202,N_285);
nand U1665 (N_1665,N_322,N_744);
or U1666 (N_1666,N_690,N_818);
nand U1667 (N_1667,N_593,N_827);
nand U1668 (N_1668,N_794,N_711);
nand U1669 (N_1669,N_236,N_643);
or U1670 (N_1670,N_956,N_591);
nand U1671 (N_1671,N_965,N_220);
or U1672 (N_1672,N_681,N_795);
nor U1673 (N_1673,N_134,N_637);
nor U1674 (N_1674,N_132,N_788);
nor U1675 (N_1675,N_845,N_287);
xnor U1676 (N_1676,N_95,N_642);
nor U1677 (N_1677,N_426,N_544);
and U1678 (N_1678,N_432,N_81);
nand U1679 (N_1679,N_232,N_377);
nor U1680 (N_1680,N_53,N_282);
nand U1681 (N_1681,N_620,N_900);
and U1682 (N_1682,N_232,N_902);
and U1683 (N_1683,N_672,N_810);
and U1684 (N_1684,N_589,N_262);
nor U1685 (N_1685,N_553,N_962);
nor U1686 (N_1686,N_209,N_729);
or U1687 (N_1687,N_818,N_742);
nand U1688 (N_1688,N_961,N_191);
nand U1689 (N_1689,N_870,N_87);
nand U1690 (N_1690,N_844,N_155);
and U1691 (N_1691,N_169,N_528);
xor U1692 (N_1692,N_655,N_430);
nor U1693 (N_1693,N_202,N_279);
nand U1694 (N_1694,N_747,N_211);
nor U1695 (N_1695,N_922,N_6);
and U1696 (N_1696,N_160,N_958);
or U1697 (N_1697,N_496,N_893);
nor U1698 (N_1698,N_390,N_631);
nand U1699 (N_1699,N_525,N_46);
nor U1700 (N_1700,N_520,N_515);
and U1701 (N_1701,N_576,N_239);
nand U1702 (N_1702,N_426,N_920);
nand U1703 (N_1703,N_922,N_548);
or U1704 (N_1704,N_526,N_232);
and U1705 (N_1705,N_521,N_121);
nor U1706 (N_1706,N_176,N_418);
nand U1707 (N_1707,N_384,N_721);
and U1708 (N_1708,N_193,N_139);
or U1709 (N_1709,N_387,N_487);
nand U1710 (N_1710,N_544,N_806);
or U1711 (N_1711,N_409,N_638);
and U1712 (N_1712,N_722,N_929);
or U1713 (N_1713,N_783,N_275);
nor U1714 (N_1714,N_632,N_613);
nand U1715 (N_1715,N_172,N_957);
nor U1716 (N_1716,N_213,N_130);
and U1717 (N_1717,N_879,N_137);
or U1718 (N_1718,N_199,N_445);
or U1719 (N_1719,N_957,N_780);
xnor U1720 (N_1720,N_84,N_874);
or U1721 (N_1721,N_708,N_878);
and U1722 (N_1722,N_193,N_953);
nand U1723 (N_1723,N_247,N_508);
and U1724 (N_1724,N_85,N_947);
and U1725 (N_1725,N_143,N_876);
nor U1726 (N_1726,N_472,N_640);
nor U1727 (N_1727,N_324,N_696);
and U1728 (N_1728,N_17,N_534);
and U1729 (N_1729,N_614,N_36);
nor U1730 (N_1730,N_790,N_870);
nand U1731 (N_1731,N_948,N_941);
nor U1732 (N_1732,N_317,N_374);
nor U1733 (N_1733,N_660,N_595);
xnor U1734 (N_1734,N_506,N_903);
nand U1735 (N_1735,N_249,N_279);
nand U1736 (N_1736,N_867,N_967);
nand U1737 (N_1737,N_53,N_679);
or U1738 (N_1738,N_81,N_651);
or U1739 (N_1739,N_27,N_384);
nand U1740 (N_1740,N_280,N_311);
and U1741 (N_1741,N_734,N_202);
nand U1742 (N_1742,N_492,N_662);
nand U1743 (N_1743,N_41,N_368);
and U1744 (N_1744,N_765,N_362);
or U1745 (N_1745,N_498,N_955);
nor U1746 (N_1746,N_517,N_533);
and U1747 (N_1747,N_606,N_487);
and U1748 (N_1748,N_332,N_458);
nor U1749 (N_1749,N_402,N_611);
nor U1750 (N_1750,N_99,N_677);
nand U1751 (N_1751,N_953,N_382);
nor U1752 (N_1752,N_13,N_746);
nor U1753 (N_1753,N_549,N_595);
nand U1754 (N_1754,N_103,N_166);
and U1755 (N_1755,N_194,N_605);
or U1756 (N_1756,N_6,N_144);
nor U1757 (N_1757,N_553,N_885);
nor U1758 (N_1758,N_554,N_257);
and U1759 (N_1759,N_626,N_163);
nand U1760 (N_1760,N_961,N_840);
or U1761 (N_1761,N_756,N_766);
or U1762 (N_1762,N_669,N_156);
nor U1763 (N_1763,N_393,N_600);
nand U1764 (N_1764,N_716,N_5);
or U1765 (N_1765,N_552,N_64);
nor U1766 (N_1766,N_0,N_234);
and U1767 (N_1767,N_271,N_778);
nor U1768 (N_1768,N_363,N_97);
nor U1769 (N_1769,N_524,N_125);
or U1770 (N_1770,N_518,N_236);
nand U1771 (N_1771,N_551,N_701);
nor U1772 (N_1772,N_278,N_633);
or U1773 (N_1773,N_721,N_413);
and U1774 (N_1774,N_277,N_518);
and U1775 (N_1775,N_123,N_477);
and U1776 (N_1776,N_754,N_204);
or U1777 (N_1777,N_982,N_843);
nand U1778 (N_1778,N_147,N_678);
and U1779 (N_1779,N_27,N_321);
xor U1780 (N_1780,N_144,N_877);
and U1781 (N_1781,N_273,N_947);
nand U1782 (N_1782,N_908,N_688);
nor U1783 (N_1783,N_602,N_758);
nor U1784 (N_1784,N_895,N_87);
nor U1785 (N_1785,N_738,N_785);
and U1786 (N_1786,N_459,N_807);
nor U1787 (N_1787,N_351,N_65);
nand U1788 (N_1788,N_481,N_479);
nor U1789 (N_1789,N_745,N_109);
nor U1790 (N_1790,N_436,N_330);
nand U1791 (N_1791,N_573,N_222);
nor U1792 (N_1792,N_797,N_587);
or U1793 (N_1793,N_694,N_447);
nand U1794 (N_1794,N_732,N_258);
nor U1795 (N_1795,N_700,N_177);
or U1796 (N_1796,N_190,N_576);
and U1797 (N_1797,N_929,N_210);
nand U1798 (N_1798,N_620,N_414);
or U1799 (N_1799,N_672,N_839);
nand U1800 (N_1800,N_2,N_295);
nand U1801 (N_1801,N_53,N_640);
or U1802 (N_1802,N_726,N_477);
and U1803 (N_1803,N_506,N_298);
or U1804 (N_1804,N_621,N_561);
or U1805 (N_1805,N_208,N_744);
nor U1806 (N_1806,N_594,N_676);
and U1807 (N_1807,N_293,N_490);
nor U1808 (N_1808,N_896,N_125);
nand U1809 (N_1809,N_606,N_650);
nand U1810 (N_1810,N_883,N_390);
nand U1811 (N_1811,N_322,N_774);
nor U1812 (N_1812,N_307,N_893);
or U1813 (N_1813,N_509,N_713);
nand U1814 (N_1814,N_81,N_982);
or U1815 (N_1815,N_584,N_39);
nand U1816 (N_1816,N_409,N_84);
and U1817 (N_1817,N_588,N_427);
nand U1818 (N_1818,N_920,N_780);
or U1819 (N_1819,N_414,N_553);
nor U1820 (N_1820,N_601,N_842);
nand U1821 (N_1821,N_866,N_379);
nand U1822 (N_1822,N_826,N_440);
nand U1823 (N_1823,N_261,N_352);
and U1824 (N_1824,N_820,N_634);
nand U1825 (N_1825,N_710,N_722);
or U1826 (N_1826,N_612,N_277);
nor U1827 (N_1827,N_115,N_405);
nand U1828 (N_1828,N_836,N_455);
or U1829 (N_1829,N_374,N_554);
or U1830 (N_1830,N_460,N_652);
nor U1831 (N_1831,N_593,N_288);
and U1832 (N_1832,N_988,N_368);
and U1833 (N_1833,N_941,N_694);
or U1834 (N_1834,N_521,N_970);
and U1835 (N_1835,N_91,N_115);
nand U1836 (N_1836,N_207,N_625);
nor U1837 (N_1837,N_165,N_544);
nand U1838 (N_1838,N_337,N_816);
nand U1839 (N_1839,N_32,N_35);
nand U1840 (N_1840,N_241,N_810);
and U1841 (N_1841,N_688,N_718);
nor U1842 (N_1842,N_138,N_925);
or U1843 (N_1843,N_775,N_145);
and U1844 (N_1844,N_871,N_798);
and U1845 (N_1845,N_251,N_337);
nor U1846 (N_1846,N_723,N_300);
or U1847 (N_1847,N_964,N_406);
nor U1848 (N_1848,N_396,N_80);
nor U1849 (N_1849,N_707,N_643);
and U1850 (N_1850,N_28,N_454);
and U1851 (N_1851,N_19,N_726);
or U1852 (N_1852,N_707,N_457);
or U1853 (N_1853,N_89,N_946);
nand U1854 (N_1854,N_447,N_314);
nand U1855 (N_1855,N_594,N_754);
xor U1856 (N_1856,N_162,N_128);
nor U1857 (N_1857,N_33,N_893);
and U1858 (N_1858,N_40,N_737);
and U1859 (N_1859,N_870,N_899);
and U1860 (N_1860,N_182,N_663);
nor U1861 (N_1861,N_702,N_135);
and U1862 (N_1862,N_503,N_538);
nor U1863 (N_1863,N_422,N_886);
nand U1864 (N_1864,N_727,N_611);
or U1865 (N_1865,N_632,N_934);
or U1866 (N_1866,N_861,N_769);
or U1867 (N_1867,N_51,N_713);
nor U1868 (N_1868,N_39,N_609);
and U1869 (N_1869,N_242,N_527);
nand U1870 (N_1870,N_736,N_748);
or U1871 (N_1871,N_722,N_188);
nand U1872 (N_1872,N_488,N_761);
or U1873 (N_1873,N_801,N_802);
and U1874 (N_1874,N_90,N_219);
or U1875 (N_1875,N_998,N_990);
and U1876 (N_1876,N_535,N_965);
nor U1877 (N_1877,N_642,N_264);
nand U1878 (N_1878,N_699,N_953);
nor U1879 (N_1879,N_344,N_665);
or U1880 (N_1880,N_338,N_317);
or U1881 (N_1881,N_358,N_13);
nand U1882 (N_1882,N_837,N_337);
or U1883 (N_1883,N_804,N_344);
nand U1884 (N_1884,N_445,N_463);
or U1885 (N_1885,N_315,N_895);
or U1886 (N_1886,N_581,N_485);
and U1887 (N_1887,N_511,N_212);
nand U1888 (N_1888,N_846,N_647);
or U1889 (N_1889,N_101,N_439);
or U1890 (N_1890,N_460,N_457);
or U1891 (N_1891,N_918,N_386);
and U1892 (N_1892,N_486,N_364);
nand U1893 (N_1893,N_456,N_491);
or U1894 (N_1894,N_717,N_193);
nor U1895 (N_1895,N_69,N_808);
and U1896 (N_1896,N_332,N_693);
nand U1897 (N_1897,N_141,N_95);
nor U1898 (N_1898,N_501,N_18);
nor U1899 (N_1899,N_591,N_231);
nor U1900 (N_1900,N_350,N_402);
and U1901 (N_1901,N_660,N_659);
nor U1902 (N_1902,N_483,N_276);
xnor U1903 (N_1903,N_252,N_817);
nand U1904 (N_1904,N_777,N_758);
and U1905 (N_1905,N_837,N_967);
or U1906 (N_1906,N_760,N_874);
and U1907 (N_1907,N_978,N_544);
and U1908 (N_1908,N_237,N_223);
and U1909 (N_1909,N_212,N_79);
or U1910 (N_1910,N_730,N_216);
or U1911 (N_1911,N_248,N_866);
or U1912 (N_1912,N_123,N_393);
nor U1913 (N_1913,N_952,N_796);
nor U1914 (N_1914,N_842,N_504);
and U1915 (N_1915,N_499,N_201);
nand U1916 (N_1916,N_555,N_114);
xnor U1917 (N_1917,N_157,N_988);
and U1918 (N_1918,N_784,N_605);
nand U1919 (N_1919,N_773,N_705);
nand U1920 (N_1920,N_901,N_130);
and U1921 (N_1921,N_49,N_11);
and U1922 (N_1922,N_31,N_889);
or U1923 (N_1923,N_195,N_855);
or U1924 (N_1924,N_764,N_942);
or U1925 (N_1925,N_245,N_448);
nand U1926 (N_1926,N_760,N_154);
and U1927 (N_1927,N_695,N_15);
nand U1928 (N_1928,N_917,N_358);
nor U1929 (N_1929,N_649,N_789);
nand U1930 (N_1930,N_395,N_792);
and U1931 (N_1931,N_287,N_983);
xnor U1932 (N_1932,N_57,N_42);
or U1933 (N_1933,N_393,N_541);
and U1934 (N_1934,N_735,N_227);
or U1935 (N_1935,N_382,N_118);
or U1936 (N_1936,N_950,N_124);
nor U1937 (N_1937,N_916,N_206);
nor U1938 (N_1938,N_550,N_561);
or U1939 (N_1939,N_542,N_195);
nand U1940 (N_1940,N_325,N_387);
nor U1941 (N_1941,N_425,N_638);
or U1942 (N_1942,N_188,N_68);
or U1943 (N_1943,N_3,N_793);
and U1944 (N_1944,N_359,N_279);
nor U1945 (N_1945,N_509,N_545);
nor U1946 (N_1946,N_472,N_741);
nand U1947 (N_1947,N_999,N_24);
or U1948 (N_1948,N_506,N_263);
and U1949 (N_1949,N_908,N_807);
and U1950 (N_1950,N_228,N_112);
and U1951 (N_1951,N_252,N_507);
or U1952 (N_1952,N_559,N_372);
and U1953 (N_1953,N_757,N_188);
nand U1954 (N_1954,N_326,N_783);
or U1955 (N_1955,N_326,N_609);
and U1956 (N_1956,N_547,N_236);
nor U1957 (N_1957,N_721,N_306);
nor U1958 (N_1958,N_80,N_388);
or U1959 (N_1959,N_463,N_914);
or U1960 (N_1960,N_300,N_919);
and U1961 (N_1961,N_512,N_409);
nor U1962 (N_1962,N_57,N_869);
or U1963 (N_1963,N_401,N_563);
or U1964 (N_1964,N_187,N_973);
or U1965 (N_1965,N_183,N_989);
and U1966 (N_1966,N_152,N_919);
and U1967 (N_1967,N_449,N_74);
or U1968 (N_1968,N_88,N_315);
nand U1969 (N_1969,N_673,N_486);
and U1970 (N_1970,N_639,N_875);
nor U1971 (N_1971,N_572,N_640);
and U1972 (N_1972,N_332,N_649);
nor U1973 (N_1973,N_649,N_848);
or U1974 (N_1974,N_383,N_836);
xnor U1975 (N_1975,N_965,N_661);
or U1976 (N_1976,N_138,N_237);
nand U1977 (N_1977,N_454,N_798);
or U1978 (N_1978,N_301,N_721);
and U1979 (N_1979,N_94,N_536);
nor U1980 (N_1980,N_468,N_402);
or U1981 (N_1981,N_432,N_112);
or U1982 (N_1982,N_254,N_389);
nor U1983 (N_1983,N_930,N_694);
nand U1984 (N_1984,N_356,N_605);
and U1985 (N_1985,N_454,N_220);
or U1986 (N_1986,N_502,N_404);
nor U1987 (N_1987,N_633,N_730);
nand U1988 (N_1988,N_114,N_288);
nor U1989 (N_1989,N_933,N_575);
and U1990 (N_1990,N_948,N_614);
or U1991 (N_1991,N_813,N_893);
nand U1992 (N_1992,N_290,N_166);
nor U1993 (N_1993,N_185,N_538);
or U1994 (N_1994,N_555,N_607);
and U1995 (N_1995,N_243,N_56);
nand U1996 (N_1996,N_162,N_662);
and U1997 (N_1997,N_626,N_958);
or U1998 (N_1998,N_113,N_332);
or U1999 (N_1999,N_669,N_415);
and U2000 (N_2000,N_1307,N_1534);
nor U2001 (N_2001,N_1229,N_1440);
nand U2002 (N_2002,N_1470,N_1488);
or U2003 (N_2003,N_1504,N_1801);
nor U2004 (N_2004,N_1429,N_1035);
nand U2005 (N_2005,N_1660,N_1262);
nor U2006 (N_2006,N_1879,N_1602);
nor U2007 (N_2007,N_1665,N_1690);
and U2008 (N_2008,N_1528,N_1086);
nand U2009 (N_2009,N_1006,N_1479);
or U2010 (N_2010,N_1437,N_1640);
nor U2011 (N_2011,N_1755,N_1386);
nor U2012 (N_2012,N_1216,N_1512);
or U2013 (N_2013,N_1092,N_1682);
nor U2014 (N_2014,N_1716,N_1244);
nor U2015 (N_2015,N_1638,N_1826);
nand U2016 (N_2016,N_1093,N_1431);
nand U2017 (N_2017,N_1727,N_1586);
and U2018 (N_2018,N_1592,N_1471);
nand U2019 (N_2019,N_1017,N_1940);
xor U2020 (N_2020,N_1966,N_1570);
nor U2021 (N_2021,N_1717,N_1062);
nor U2022 (N_2022,N_1579,N_1725);
or U2023 (N_2023,N_1162,N_1938);
nor U2024 (N_2024,N_1712,N_1274);
nand U2025 (N_2025,N_1719,N_1650);
nand U2026 (N_2026,N_1078,N_1347);
or U2027 (N_2027,N_1907,N_1654);
nand U2028 (N_2028,N_1365,N_1409);
or U2029 (N_2029,N_1530,N_1259);
nor U2030 (N_2030,N_1079,N_1831);
and U2031 (N_2031,N_1893,N_1948);
nor U2032 (N_2032,N_1781,N_1340);
nor U2033 (N_2033,N_1549,N_1069);
and U2034 (N_2034,N_1761,N_1758);
and U2035 (N_2035,N_1770,N_1258);
and U2036 (N_2036,N_1949,N_1523);
nand U2037 (N_2037,N_1203,N_1361);
or U2038 (N_2038,N_1656,N_1873);
nor U2039 (N_2039,N_1862,N_1852);
and U2040 (N_2040,N_1005,N_1388);
nand U2041 (N_2041,N_1942,N_1188);
nand U2042 (N_2042,N_1978,N_1498);
nand U2043 (N_2043,N_1950,N_1765);
and U2044 (N_2044,N_1449,N_1676);
or U2045 (N_2045,N_1526,N_1000);
and U2046 (N_2046,N_1769,N_1222);
and U2047 (N_2047,N_1446,N_1641);
or U2048 (N_2048,N_1915,N_1473);
and U2049 (N_2049,N_1497,N_1689);
or U2050 (N_2050,N_1700,N_1010);
xnor U2051 (N_2051,N_1568,N_1125);
nor U2052 (N_2052,N_1351,N_1320);
and U2053 (N_2053,N_1809,N_1913);
nor U2054 (N_2054,N_1159,N_1445);
xnor U2055 (N_2055,N_1402,N_1970);
nand U2056 (N_2056,N_1548,N_1668);
nor U2057 (N_2057,N_1545,N_1969);
and U2058 (N_2058,N_1444,N_1757);
and U2059 (N_2059,N_1461,N_1465);
nand U2060 (N_2060,N_1042,N_1711);
and U2061 (N_2061,N_1778,N_1101);
nor U2062 (N_2062,N_1945,N_1722);
and U2063 (N_2063,N_1897,N_1655);
nor U2064 (N_2064,N_1904,N_1301);
nand U2065 (N_2065,N_1776,N_1968);
nor U2066 (N_2066,N_1242,N_1118);
xnor U2067 (N_2067,N_1923,N_1191);
nand U2068 (N_2068,N_1344,N_1580);
nor U2069 (N_2069,N_1956,N_1173);
nand U2070 (N_2070,N_1922,N_1363);
or U2071 (N_2071,N_1859,N_1611);
nand U2072 (N_2072,N_1605,N_1463);
nor U2073 (N_2073,N_1318,N_1898);
and U2074 (N_2074,N_1051,N_1232);
xor U2075 (N_2075,N_1517,N_1126);
or U2076 (N_2076,N_1315,N_1477);
nor U2077 (N_2077,N_1759,N_1306);
nand U2078 (N_2078,N_1516,N_1934);
or U2079 (N_2079,N_1235,N_1043);
nor U2080 (N_2080,N_1960,N_1877);
nand U2081 (N_2081,N_1348,N_1182);
and U2082 (N_2082,N_1730,N_1028);
and U2083 (N_2083,N_1167,N_1190);
nor U2084 (N_2084,N_1397,N_1398);
and U2085 (N_2085,N_1275,N_1659);
nor U2086 (N_2086,N_1202,N_1925);
and U2087 (N_2087,N_1147,N_1379);
xor U2088 (N_2088,N_1239,N_1982);
and U2089 (N_2089,N_1436,N_1736);
or U2090 (N_2090,N_1603,N_1697);
nand U2091 (N_2091,N_1657,N_1642);
nor U2092 (N_2092,N_1869,N_1354);
xnor U2093 (N_2093,N_1481,N_1854);
nand U2094 (N_2094,N_1120,N_1296);
nor U2095 (N_2095,N_1482,N_1377);
or U2096 (N_2096,N_1735,N_1292);
or U2097 (N_2097,N_1175,N_1737);
or U2098 (N_2098,N_1334,N_1376);
and U2099 (N_2099,N_1688,N_1228);
and U2100 (N_2100,N_1316,N_1583);
or U2101 (N_2101,N_1090,N_1492);
or U2102 (N_2102,N_1508,N_1663);
or U2103 (N_2103,N_1888,N_1382);
or U2104 (N_2104,N_1231,N_1550);
nand U2105 (N_2105,N_1076,N_1073);
or U2106 (N_2106,N_1667,N_1658);
and U2107 (N_2107,N_1480,N_1752);
or U2108 (N_2108,N_1196,N_1872);
or U2109 (N_2109,N_1068,N_1527);
nor U2110 (N_2110,N_1369,N_1355);
nand U2111 (N_2111,N_1706,N_1693);
and U2112 (N_2112,N_1815,N_1691);
nand U2113 (N_2113,N_1082,N_1217);
nor U2114 (N_2114,N_1339,N_1977);
or U2115 (N_2115,N_1738,N_1142);
nor U2116 (N_2116,N_1600,N_1958);
and U2117 (N_2117,N_1598,N_1824);
nand U2118 (N_2118,N_1720,N_1786);
or U2119 (N_2119,N_1687,N_1303);
or U2120 (N_2120,N_1614,N_1390);
xor U2121 (N_2121,N_1562,N_1053);
nand U2122 (N_2122,N_1260,N_1763);
and U2123 (N_2123,N_1176,N_1694);
nand U2124 (N_2124,N_1885,N_1476);
or U2125 (N_2125,N_1410,N_1561);
nand U2126 (N_2126,N_1353,N_1279);
nand U2127 (N_2127,N_1785,N_1345);
nor U2128 (N_2128,N_1400,N_1556);
nor U2129 (N_2129,N_1679,N_1782);
nor U2130 (N_2130,N_1109,N_1161);
nand U2131 (N_2131,N_1812,N_1403);
or U2132 (N_2132,N_1462,N_1341);
nor U2133 (N_2133,N_1247,N_1324);
nor U2134 (N_2134,N_1633,N_1245);
and U2135 (N_2135,N_1936,N_1077);
nand U2136 (N_2136,N_1312,N_1485);
nor U2137 (N_2137,N_1146,N_1140);
nand U2138 (N_2138,N_1004,N_1417);
or U2139 (N_2139,N_1947,N_1343);
nor U2140 (N_2140,N_1074,N_1141);
or U2141 (N_2141,N_1362,N_1513);
nor U2142 (N_2142,N_1129,N_1529);
nand U2143 (N_2143,N_1645,N_1851);
and U2144 (N_2144,N_1566,N_1571);
or U2145 (N_2145,N_1021,N_1286);
nor U2146 (N_2146,N_1180,N_1623);
nand U2147 (N_2147,N_1048,N_1984);
and U2148 (N_2148,N_1935,N_1853);
and U2149 (N_2149,N_1384,N_1186);
nor U2150 (N_2150,N_1002,N_1880);
nand U2151 (N_2151,N_1747,N_1046);
nand U2152 (N_2152,N_1317,N_1993);
and U2153 (N_2153,N_1091,N_1961);
or U2154 (N_2154,N_1111,N_1165);
and U2155 (N_2155,N_1096,N_1237);
xnor U2156 (N_2156,N_1024,N_1174);
nand U2157 (N_2157,N_1756,N_1308);
nand U2158 (N_2158,N_1675,N_1768);
nor U2159 (N_2159,N_1849,N_1543);
and U2160 (N_2160,N_1421,N_1336);
nand U2161 (N_2161,N_1559,N_1327);
or U2162 (N_2162,N_1472,N_1536);
nand U2163 (N_2163,N_1293,N_1025);
nor U2164 (N_2164,N_1774,N_1882);
nand U2165 (N_2165,N_1932,N_1300);
and U2166 (N_2166,N_1484,N_1749);
nand U2167 (N_2167,N_1066,N_1843);
nor U2168 (N_2168,N_1825,N_1926);
or U2169 (N_2169,N_1425,N_1796);
and U2170 (N_2170,N_1531,N_1589);
nor U2171 (N_2171,N_1451,N_1015);
and U2172 (N_2172,N_1772,N_1804);
and U2173 (N_2173,N_1263,N_1597);
or U2174 (N_2174,N_1820,N_1364);
and U2175 (N_2175,N_1486,N_1503);
or U2176 (N_2176,N_1442,N_1154);
nor U2177 (N_2177,N_1405,N_1617);
nand U2178 (N_2178,N_1204,N_1314);
and U2179 (N_2179,N_1927,N_1407);
nor U2180 (N_2180,N_1569,N_1621);
nor U2181 (N_2181,N_1903,N_1194);
and U2182 (N_2182,N_1268,N_1418);
nor U2183 (N_2183,N_1835,N_1065);
nor U2184 (N_2184,N_1828,N_1878);
nand U2185 (N_2185,N_1813,N_1610);
nor U2186 (N_2186,N_1489,N_1917);
and U2187 (N_2187,N_1726,N_1766);
or U2188 (N_2188,N_1883,N_1537);
and U2189 (N_2189,N_1585,N_1653);
or U2190 (N_2190,N_1322,N_1951);
nor U2191 (N_2191,N_1514,N_1220);
or U2192 (N_2192,N_1064,N_1703);
and U2193 (N_2193,N_1789,N_1171);
nand U2194 (N_2194,N_1153,N_1001);
or U2195 (N_2195,N_1563,N_1587);
or U2196 (N_2196,N_1817,N_1670);
or U2197 (N_2197,N_1088,N_1810);
nor U2198 (N_2198,N_1187,N_1325);
and U2199 (N_2199,N_1211,N_1535);
nand U2200 (N_2200,N_1920,N_1057);
xnor U2201 (N_2201,N_1494,N_1764);
and U2202 (N_2202,N_1075,N_1741);
nand U2203 (N_2203,N_1681,N_1166);
and U2204 (N_2204,N_1609,N_1867);
nor U2205 (N_2205,N_1150,N_1169);
nand U2206 (N_2206,N_1210,N_1834);
nor U2207 (N_2207,N_1930,N_1013);
and U2208 (N_2208,N_1071,N_1988);
xnor U2209 (N_2209,N_1085,N_1201);
nor U2210 (N_2210,N_1252,N_1366);
and U2211 (N_2211,N_1249,N_1019);
or U2212 (N_2212,N_1792,N_1282);
or U2213 (N_2213,N_1295,N_1328);
nor U2214 (N_2214,N_1814,N_1375);
or U2215 (N_2215,N_1775,N_1123);
nor U2216 (N_2216,N_1372,N_1469);
nor U2217 (N_2217,N_1790,N_1290);
or U2218 (N_2218,N_1806,N_1246);
nor U2219 (N_2219,N_1291,N_1520);
nor U2220 (N_2220,N_1370,N_1900);
nor U2221 (N_2221,N_1627,N_1330);
nor U2222 (N_2222,N_1373,N_1499);
and U2223 (N_2223,N_1198,N_1404);
nand U2224 (N_2224,N_1047,N_1464);
nor U2225 (N_2225,N_1857,N_1729);
and U2226 (N_2226,N_1261,N_1845);
or U2227 (N_2227,N_1981,N_1428);
xor U2228 (N_2228,N_1127,N_1116);
or U2229 (N_2229,N_1063,N_1624);
and U2230 (N_2230,N_1505,N_1713);
nand U2231 (N_2231,N_1594,N_1954);
or U2232 (N_2232,N_1215,N_1992);
and U2233 (N_2233,N_1224,N_1193);
nand U2234 (N_2234,N_1619,N_1858);
nor U2235 (N_2235,N_1933,N_1420);
xor U2236 (N_2236,N_1467,N_1164);
or U2237 (N_2237,N_1266,N_1276);
nor U2238 (N_2238,N_1281,N_1784);
or U2239 (N_2239,N_1698,N_1884);
nor U2240 (N_2240,N_1762,N_1524);
nand U2241 (N_2241,N_1137,N_1299);
nand U2242 (N_2242,N_1124,N_1952);
or U2243 (N_2243,N_1034,N_1385);
nand U2244 (N_2244,N_1582,N_1692);
nor U2245 (N_2245,N_1648,N_1780);
nand U2246 (N_2246,N_1329,N_1115);
nand U2247 (N_2247,N_1117,N_1226);
nand U2248 (N_2248,N_1728,N_1604);
and U2249 (N_2249,N_1636,N_1413);
or U2250 (N_2250,N_1056,N_1967);
or U2251 (N_2251,N_1510,N_1731);
and U2252 (N_2252,N_1448,N_1906);
and U2253 (N_2253,N_1715,N_1267);
nand U2254 (N_2254,N_1432,N_1718);
and U2255 (N_2255,N_1595,N_1827);
or U2256 (N_2256,N_1836,N_1995);
nand U2257 (N_2257,N_1319,N_1613);
nor U2258 (N_2258,N_1760,N_1918);
and U2259 (N_2259,N_1646,N_1661);
and U2260 (N_2260,N_1225,N_1238);
or U2261 (N_2261,N_1230,N_1509);
nand U2262 (N_2262,N_1389,N_1170);
nand U2263 (N_2263,N_1861,N_1639);
nand U2264 (N_2264,N_1380,N_1278);
or U2265 (N_2265,N_1601,N_1138);
nor U2266 (N_2266,N_1212,N_1045);
nor U2267 (N_2267,N_1634,N_1447);
nor U2268 (N_2268,N_1061,N_1576);
nor U2269 (N_2269,N_1547,N_1136);
nand U2270 (N_2270,N_1108,N_1538);
nand U2271 (N_2271,N_1145,N_1119);
nand U2272 (N_2272,N_1644,N_1651);
nor U2273 (N_2273,N_1012,N_1501);
or U2274 (N_2274,N_1975,N_1822);
or U2275 (N_2275,N_1352,N_1856);
nor U2276 (N_2276,N_1026,N_1483);
nand U2277 (N_2277,N_1060,N_1829);
or U2278 (N_2278,N_1899,N_1475);
nor U2279 (N_2279,N_1236,N_1632);
or U2280 (N_2280,N_1953,N_1864);
or U2281 (N_2281,N_1020,N_1921);
and U2282 (N_2282,N_1909,N_1438);
nand U2283 (N_2283,N_1052,N_1748);
nand U2284 (N_2284,N_1423,N_1998);
and U2285 (N_2285,N_1837,N_1037);
nor U2286 (N_2286,N_1257,N_1374);
and U2287 (N_2287,N_1072,N_1155);
and U2288 (N_2288,N_1087,N_1014);
nor U2289 (N_2289,N_1011,N_1038);
nor U2290 (N_2290,N_1144,N_1100);
nand U2291 (N_2291,N_1132,N_1099);
nand U2292 (N_2292,N_1795,N_1183);
nor U2293 (N_2293,N_1331,N_1359);
and U2294 (N_2294,N_1205,N_1098);
or U2295 (N_2295,N_1590,N_1886);
nand U2296 (N_2296,N_1185,N_1452);
and U2297 (N_2297,N_1050,N_1674);
nor U2298 (N_2298,N_1989,N_1647);
nor U2299 (N_2299,N_1532,N_1192);
or U2300 (N_2300,N_1112,N_1049);
or U2301 (N_2301,N_1607,N_1067);
or U2302 (N_2302,N_1030,N_1889);
and U2303 (N_2303,N_1914,N_1294);
and U2304 (N_2304,N_1671,N_1393);
nand U2305 (N_2305,N_1626,N_1771);
nand U2306 (N_2306,N_1114,N_1288);
and U2307 (N_2307,N_1608,N_1102);
and U2308 (N_2308,N_1468,N_1036);
xnor U2309 (N_2309,N_1816,N_1459);
or U2310 (N_2310,N_1433,N_1416);
nand U2311 (N_2311,N_1350,N_1957);
nand U2312 (N_2312,N_1892,N_1788);
and U2313 (N_2313,N_1008,N_1901);
and U2314 (N_2314,N_1539,N_1846);
nor U2315 (N_2315,N_1911,N_1678);
nand U2316 (N_2316,N_1223,N_1751);
and U2317 (N_2317,N_1832,N_1773);
or U2318 (N_2318,N_1250,N_1199);
and U2319 (N_2319,N_1996,N_1016);
or U2320 (N_2320,N_1151,N_1573);
nor U2321 (N_2321,N_1551,N_1284);
nor U2322 (N_2322,N_1213,N_1148);
and U2323 (N_2323,N_1669,N_1553);
and U2324 (N_2324,N_1896,N_1860);
or U2325 (N_2325,N_1179,N_1387);
nand U2326 (N_2326,N_1924,N_1441);
nor U2327 (N_2327,N_1818,N_1696);
nor U2328 (N_2328,N_1044,N_1971);
or U2329 (N_2329,N_1955,N_1839);
or U2330 (N_2330,N_1985,N_1283);
or U2331 (N_2331,N_1723,N_1980);
or U2332 (N_2332,N_1027,N_1411);
or U2333 (N_2333,N_1285,N_1221);
xnor U2334 (N_2334,N_1596,N_1652);
and U2335 (N_2335,N_1163,N_1705);
nand U2336 (N_2336,N_1401,N_1708);
and U2337 (N_2337,N_1040,N_1890);
and U2338 (N_2338,N_1577,N_1875);
or U2339 (N_2339,N_1139,N_1280);
nor U2340 (N_2340,N_1360,N_1206);
nand U2341 (N_2341,N_1160,N_1131);
or U2342 (N_2342,N_1219,N_1113);
and U2343 (N_2343,N_1699,N_1800);
and U2344 (N_2344,N_1855,N_1743);
nand U2345 (N_2345,N_1256,N_1335);
nor U2346 (N_2346,N_1628,N_1309);
and U2347 (N_2347,N_1939,N_1630);
nor U2348 (N_2348,N_1039,N_1134);
or U2349 (N_2349,N_1152,N_1787);
nor U2350 (N_2350,N_1218,N_1253);
or U2351 (N_2351,N_1805,N_1833);
or U2352 (N_2352,N_1097,N_1168);
nor U2353 (N_2353,N_1214,N_1519);
or U2354 (N_2354,N_1631,N_1578);
nor U2355 (N_2355,N_1346,N_1332);
nand U2356 (N_2356,N_1635,N_1083);
xnor U2357 (N_2357,N_1866,N_1754);
nand U2358 (N_2358,N_1629,N_1838);
nand U2359 (N_2359,N_1394,N_1511);
nor U2360 (N_2360,N_1745,N_1902);
nand U2361 (N_2361,N_1991,N_1599);
and U2362 (N_2362,N_1337,N_1615);
and U2363 (N_2363,N_1287,N_1426);
nor U2364 (N_2364,N_1986,N_1891);
and U2365 (N_2365,N_1121,N_1894);
or U2366 (N_2366,N_1910,N_1392);
nor U2367 (N_2367,N_1189,N_1022);
or U2368 (N_2368,N_1031,N_1518);
nor U2369 (N_2369,N_1620,N_1546);
nor U2370 (N_2370,N_1540,N_1181);
nand U2371 (N_2371,N_1094,N_1739);
and U2372 (N_2372,N_1349,N_1973);
or U2373 (N_2373,N_1574,N_1271);
nand U2374 (N_2374,N_1172,N_1686);
nand U2375 (N_2375,N_1821,N_1265);
or U2376 (N_2376,N_1310,N_1059);
and U2377 (N_2377,N_1702,N_1430);
nand U2378 (N_2378,N_1707,N_1564);
nand U2379 (N_2379,N_1807,N_1870);
nor U2380 (N_2380,N_1055,N_1106);
or U2381 (N_2381,N_1740,N_1422);
nand U2382 (N_2382,N_1302,N_1378);
or U2383 (N_2383,N_1871,N_1311);
nor U2384 (N_2384,N_1704,N_1128);
nor U2385 (N_2385,N_1721,N_1248);
or U2386 (N_2386,N_1474,N_1500);
nand U2387 (N_2387,N_1797,N_1750);
nand U2388 (N_2388,N_1666,N_1495);
and U2389 (N_2389,N_1803,N_1777);
or U2390 (N_2390,N_1943,N_1009);
and U2391 (N_2391,N_1876,N_1156);
and U2392 (N_2392,N_1522,N_1070);
and U2393 (N_2393,N_1999,N_1233);
or U2394 (N_2394,N_1356,N_1673);
or U2395 (N_2395,N_1637,N_1408);
or U2396 (N_2396,N_1798,N_1542);
or U2397 (N_2397,N_1478,N_1701);
or U2398 (N_2398,N_1558,N_1555);
or U2399 (N_2399,N_1625,N_1456);
nand U2400 (N_2400,N_1412,N_1427);
nand U2401 (N_2401,N_1841,N_1865);
and U2402 (N_2402,N_1868,N_1819);
and U2403 (N_2403,N_1983,N_1714);
nor U2404 (N_2404,N_1808,N_1184);
xor U2405 (N_2405,N_1919,N_1506);
and U2406 (N_2406,N_1916,N_1502);
and U2407 (N_2407,N_1227,N_1272);
and U2408 (N_2408,N_1089,N_1107);
and U2409 (N_2409,N_1593,N_1779);
nand U2410 (N_2410,N_1466,N_1618);
and U2411 (N_2411,N_1251,N_1453);
and U2412 (N_2412,N_1965,N_1994);
nor U2413 (N_2413,N_1054,N_1080);
or U2414 (N_2414,N_1929,N_1643);
and U2415 (N_2415,N_1460,N_1612);
and U2416 (N_2416,N_1490,N_1326);
or U2417 (N_2417,N_1842,N_1616);
nor U2418 (N_2418,N_1240,N_1912);
nor U2419 (N_2419,N_1987,N_1525);
nand U2420 (N_2420,N_1895,N_1304);
nand U2421 (N_2421,N_1685,N_1990);
or U2422 (N_2422,N_1560,N_1439);
and U2423 (N_2423,N_1584,N_1964);
nor U2424 (N_2424,N_1143,N_1371);
nand U2425 (N_2425,N_1081,N_1588);
nor U2426 (N_2426,N_1533,N_1130);
nand U2427 (N_2427,N_1208,N_1793);
nand U2428 (N_2428,N_1567,N_1084);
nor U2429 (N_2429,N_1496,N_1434);
or U2430 (N_2430,N_1783,N_1333);
or U2431 (N_2431,N_1794,N_1976);
nand U2432 (N_2432,N_1840,N_1207);
or U2433 (N_2433,N_1032,N_1269);
or U2434 (N_2434,N_1158,N_1414);
or U2435 (N_2435,N_1887,N_1135);
xnor U2436 (N_2436,N_1799,N_1368);
or U2437 (N_2437,N_1305,N_1338);
and U2438 (N_2438,N_1767,N_1110);
and U2439 (N_2439,N_1830,N_1881);
or U2440 (N_2440,N_1018,N_1342);
or U2441 (N_2441,N_1255,N_1680);
nand U2442 (N_2442,N_1450,N_1104);
nor U2443 (N_2443,N_1243,N_1734);
nor U2444 (N_2444,N_1406,N_1095);
nor U2445 (N_2445,N_1905,N_1742);
or U2446 (N_2446,N_1554,N_1358);
nand U2447 (N_2447,N_1541,N_1023);
nor U2448 (N_2448,N_1298,N_1908);
xor U2449 (N_2449,N_1321,N_1487);
and U2450 (N_2450,N_1732,N_1695);
or U2451 (N_2451,N_1277,N_1844);
and U2452 (N_2452,N_1591,N_1455);
nor U2453 (N_2453,N_1963,N_1848);
or U2454 (N_2454,N_1724,N_1937);
nor U2455 (N_2455,N_1744,N_1493);
or U2456 (N_2456,N_1133,N_1289);
nand U2457 (N_2457,N_1946,N_1007);
or U2458 (N_2458,N_1003,N_1200);
nor U2459 (N_2459,N_1058,N_1974);
nor U2460 (N_2460,N_1381,N_1383);
nor U2461 (N_2461,N_1122,N_1041);
nor U2462 (N_2462,N_1649,N_1391);
nor U2463 (N_2463,N_1850,N_1823);
nor U2464 (N_2464,N_1419,N_1273);
or U2465 (N_2465,N_1234,N_1515);
nand U2466 (N_2466,N_1457,N_1997);
or U2467 (N_2467,N_1270,N_1454);
and U2468 (N_2468,N_1662,N_1149);
or U2469 (N_2469,N_1622,N_1572);
nor U2470 (N_2470,N_1415,N_1847);
nor U2471 (N_2471,N_1399,N_1684);
and U2472 (N_2472,N_1195,N_1029);
nor U2473 (N_2473,N_1357,N_1177);
nor U2474 (N_2474,N_1753,N_1395);
nor U2475 (N_2475,N_1979,N_1552);
and U2476 (N_2476,N_1791,N_1209);
nor U2477 (N_2477,N_1491,N_1435);
nor U2478 (N_2478,N_1557,N_1241);
nand U2479 (N_2479,N_1944,N_1105);
nor U2480 (N_2480,N_1931,N_1521);
nor U2481 (N_2481,N_1606,N_1507);
or U2482 (N_2482,N_1581,N_1683);
nand U2483 (N_2483,N_1677,N_1178);
or U2484 (N_2484,N_1443,N_1733);
nor U2485 (N_2485,N_1033,N_1941);
nor U2486 (N_2486,N_1254,N_1575);
nor U2487 (N_2487,N_1424,N_1709);
or U2488 (N_2488,N_1972,N_1458);
nor U2489 (N_2489,N_1313,N_1746);
nand U2490 (N_2490,N_1157,N_1802);
or U2491 (N_2491,N_1544,N_1264);
or U2492 (N_2492,N_1565,N_1297);
or U2493 (N_2493,N_1962,N_1811);
nand U2494 (N_2494,N_1874,N_1710);
nor U2495 (N_2495,N_1863,N_1197);
or U2496 (N_2496,N_1928,N_1103);
nor U2497 (N_2497,N_1323,N_1664);
nor U2498 (N_2498,N_1959,N_1367);
and U2499 (N_2499,N_1672,N_1396);
nor U2500 (N_2500,N_1434,N_1060);
nand U2501 (N_2501,N_1617,N_1590);
nor U2502 (N_2502,N_1570,N_1403);
nand U2503 (N_2503,N_1896,N_1622);
and U2504 (N_2504,N_1585,N_1364);
or U2505 (N_2505,N_1959,N_1932);
nand U2506 (N_2506,N_1836,N_1258);
and U2507 (N_2507,N_1584,N_1431);
or U2508 (N_2508,N_1851,N_1937);
and U2509 (N_2509,N_1632,N_1652);
nor U2510 (N_2510,N_1458,N_1991);
nor U2511 (N_2511,N_1995,N_1065);
or U2512 (N_2512,N_1354,N_1023);
nand U2513 (N_2513,N_1756,N_1641);
or U2514 (N_2514,N_1262,N_1347);
xor U2515 (N_2515,N_1187,N_1414);
nand U2516 (N_2516,N_1249,N_1200);
nand U2517 (N_2517,N_1824,N_1958);
or U2518 (N_2518,N_1922,N_1114);
and U2519 (N_2519,N_1278,N_1790);
or U2520 (N_2520,N_1004,N_1864);
or U2521 (N_2521,N_1026,N_1724);
and U2522 (N_2522,N_1682,N_1510);
xnor U2523 (N_2523,N_1737,N_1631);
and U2524 (N_2524,N_1267,N_1409);
and U2525 (N_2525,N_1405,N_1813);
nand U2526 (N_2526,N_1214,N_1774);
nor U2527 (N_2527,N_1333,N_1564);
or U2528 (N_2528,N_1538,N_1641);
nor U2529 (N_2529,N_1462,N_1983);
nand U2530 (N_2530,N_1014,N_1852);
or U2531 (N_2531,N_1997,N_1093);
nor U2532 (N_2532,N_1309,N_1780);
nor U2533 (N_2533,N_1246,N_1247);
or U2534 (N_2534,N_1724,N_1854);
and U2535 (N_2535,N_1710,N_1576);
nand U2536 (N_2536,N_1125,N_1592);
nor U2537 (N_2537,N_1155,N_1606);
nor U2538 (N_2538,N_1705,N_1539);
or U2539 (N_2539,N_1955,N_1912);
nand U2540 (N_2540,N_1816,N_1920);
and U2541 (N_2541,N_1209,N_1222);
or U2542 (N_2542,N_1843,N_1358);
nand U2543 (N_2543,N_1483,N_1183);
nand U2544 (N_2544,N_1421,N_1919);
or U2545 (N_2545,N_1640,N_1479);
nand U2546 (N_2546,N_1445,N_1935);
nand U2547 (N_2547,N_1887,N_1806);
nand U2548 (N_2548,N_1738,N_1982);
nor U2549 (N_2549,N_1490,N_1799);
nor U2550 (N_2550,N_1451,N_1516);
or U2551 (N_2551,N_1841,N_1623);
and U2552 (N_2552,N_1491,N_1742);
or U2553 (N_2553,N_1541,N_1555);
and U2554 (N_2554,N_1822,N_1083);
nor U2555 (N_2555,N_1710,N_1929);
and U2556 (N_2556,N_1049,N_1345);
and U2557 (N_2557,N_1778,N_1398);
xnor U2558 (N_2558,N_1201,N_1133);
nand U2559 (N_2559,N_1967,N_1096);
and U2560 (N_2560,N_1531,N_1681);
or U2561 (N_2561,N_1438,N_1682);
and U2562 (N_2562,N_1649,N_1137);
nand U2563 (N_2563,N_1538,N_1704);
and U2564 (N_2564,N_1632,N_1464);
nand U2565 (N_2565,N_1886,N_1209);
nand U2566 (N_2566,N_1347,N_1936);
nor U2567 (N_2567,N_1663,N_1630);
nor U2568 (N_2568,N_1735,N_1381);
or U2569 (N_2569,N_1145,N_1365);
nand U2570 (N_2570,N_1967,N_1900);
or U2571 (N_2571,N_1886,N_1913);
nor U2572 (N_2572,N_1482,N_1100);
nand U2573 (N_2573,N_1835,N_1428);
and U2574 (N_2574,N_1861,N_1357);
xnor U2575 (N_2575,N_1703,N_1060);
xnor U2576 (N_2576,N_1101,N_1087);
nand U2577 (N_2577,N_1113,N_1664);
nand U2578 (N_2578,N_1580,N_1264);
and U2579 (N_2579,N_1864,N_1752);
or U2580 (N_2580,N_1181,N_1869);
or U2581 (N_2581,N_1678,N_1422);
nor U2582 (N_2582,N_1089,N_1786);
nor U2583 (N_2583,N_1131,N_1271);
nor U2584 (N_2584,N_1691,N_1999);
and U2585 (N_2585,N_1784,N_1047);
or U2586 (N_2586,N_1177,N_1073);
nor U2587 (N_2587,N_1119,N_1847);
and U2588 (N_2588,N_1792,N_1755);
and U2589 (N_2589,N_1317,N_1338);
and U2590 (N_2590,N_1065,N_1460);
and U2591 (N_2591,N_1432,N_1006);
nand U2592 (N_2592,N_1135,N_1326);
nor U2593 (N_2593,N_1095,N_1727);
nor U2594 (N_2594,N_1708,N_1778);
and U2595 (N_2595,N_1285,N_1578);
nor U2596 (N_2596,N_1088,N_1279);
or U2597 (N_2597,N_1904,N_1256);
nor U2598 (N_2598,N_1642,N_1394);
nor U2599 (N_2599,N_1011,N_1623);
or U2600 (N_2600,N_1958,N_1261);
and U2601 (N_2601,N_1865,N_1106);
nor U2602 (N_2602,N_1469,N_1213);
nor U2603 (N_2603,N_1782,N_1943);
nand U2604 (N_2604,N_1703,N_1776);
nand U2605 (N_2605,N_1224,N_1700);
nand U2606 (N_2606,N_1710,N_1186);
and U2607 (N_2607,N_1954,N_1537);
nand U2608 (N_2608,N_1120,N_1730);
nand U2609 (N_2609,N_1411,N_1178);
and U2610 (N_2610,N_1197,N_1206);
and U2611 (N_2611,N_1267,N_1637);
nand U2612 (N_2612,N_1861,N_1386);
nand U2613 (N_2613,N_1792,N_1138);
nand U2614 (N_2614,N_1100,N_1188);
xor U2615 (N_2615,N_1428,N_1423);
or U2616 (N_2616,N_1719,N_1513);
nand U2617 (N_2617,N_1604,N_1175);
nor U2618 (N_2618,N_1920,N_1327);
and U2619 (N_2619,N_1472,N_1953);
and U2620 (N_2620,N_1479,N_1650);
or U2621 (N_2621,N_1750,N_1027);
and U2622 (N_2622,N_1002,N_1761);
nand U2623 (N_2623,N_1563,N_1851);
nor U2624 (N_2624,N_1063,N_1354);
nor U2625 (N_2625,N_1022,N_1828);
nand U2626 (N_2626,N_1179,N_1025);
nand U2627 (N_2627,N_1082,N_1013);
nand U2628 (N_2628,N_1531,N_1405);
and U2629 (N_2629,N_1168,N_1751);
or U2630 (N_2630,N_1065,N_1543);
or U2631 (N_2631,N_1231,N_1988);
nand U2632 (N_2632,N_1043,N_1388);
or U2633 (N_2633,N_1198,N_1541);
nand U2634 (N_2634,N_1386,N_1812);
and U2635 (N_2635,N_1915,N_1625);
and U2636 (N_2636,N_1812,N_1301);
and U2637 (N_2637,N_1386,N_1781);
nand U2638 (N_2638,N_1526,N_1021);
xor U2639 (N_2639,N_1493,N_1481);
nand U2640 (N_2640,N_1828,N_1767);
nand U2641 (N_2641,N_1338,N_1064);
nor U2642 (N_2642,N_1505,N_1091);
nand U2643 (N_2643,N_1553,N_1656);
nand U2644 (N_2644,N_1581,N_1511);
nand U2645 (N_2645,N_1204,N_1139);
or U2646 (N_2646,N_1769,N_1553);
and U2647 (N_2647,N_1958,N_1537);
nand U2648 (N_2648,N_1637,N_1596);
or U2649 (N_2649,N_1589,N_1043);
and U2650 (N_2650,N_1831,N_1415);
or U2651 (N_2651,N_1788,N_1364);
nor U2652 (N_2652,N_1391,N_1688);
or U2653 (N_2653,N_1854,N_1156);
or U2654 (N_2654,N_1202,N_1636);
nand U2655 (N_2655,N_1883,N_1025);
and U2656 (N_2656,N_1587,N_1800);
nand U2657 (N_2657,N_1438,N_1579);
nand U2658 (N_2658,N_1439,N_1901);
nand U2659 (N_2659,N_1381,N_1515);
and U2660 (N_2660,N_1560,N_1659);
nor U2661 (N_2661,N_1399,N_1012);
nor U2662 (N_2662,N_1353,N_1419);
nor U2663 (N_2663,N_1318,N_1664);
nand U2664 (N_2664,N_1698,N_1415);
and U2665 (N_2665,N_1279,N_1412);
nor U2666 (N_2666,N_1049,N_1260);
or U2667 (N_2667,N_1610,N_1799);
or U2668 (N_2668,N_1977,N_1655);
or U2669 (N_2669,N_1628,N_1654);
and U2670 (N_2670,N_1424,N_1122);
or U2671 (N_2671,N_1050,N_1478);
nand U2672 (N_2672,N_1245,N_1932);
xor U2673 (N_2673,N_1806,N_1539);
and U2674 (N_2674,N_1297,N_1732);
or U2675 (N_2675,N_1362,N_1478);
nor U2676 (N_2676,N_1196,N_1476);
nor U2677 (N_2677,N_1494,N_1347);
nor U2678 (N_2678,N_1941,N_1403);
nor U2679 (N_2679,N_1067,N_1967);
nand U2680 (N_2680,N_1614,N_1335);
and U2681 (N_2681,N_1055,N_1843);
nor U2682 (N_2682,N_1832,N_1290);
and U2683 (N_2683,N_1353,N_1948);
or U2684 (N_2684,N_1689,N_1680);
nor U2685 (N_2685,N_1277,N_1382);
nor U2686 (N_2686,N_1525,N_1876);
and U2687 (N_2687,N_1393,N_1689);
xnor U2688 (N_2688,N_1091,N_1886);
or U2689 (N_2689,N_1266,N_1663);
nand U2690 (N_2690,N_1995,N_1223);
and U2691 (N_2691,N_1949,N_1692);
or U2692 (N_2692,N_1482,N_1585);
or U2693 (N_2693,N_1434,N_1346);
or U2694 (N_2694,N_1721,N_1709);
nor U2695 (N_2695,N_1681,N_1904);
or U2696 (N_2696,N_1475,N_1609);
or U2697 (N_2697,N_1171,N_1487);
or U2698 (N_2698,N_1737,N_1255);
or U2699 (N_2699,N_1092,N_1586);
nor U2700 (N_2700,N_1483,N_1050);
or U2701 (N_2701,N_1504,N_1149);
nor U2702 (N_2702,N_1974,N_1964);
nor U2703 (N_2703,N_1844,N_1656);
and U2704 (N_2704,N_1388,N_1926);
or U2705 (N_2705,N_1679,N_1523);
nor U2706 (N_2706,N_1466,N_1965);
nand U2707 (N_2707,N_1148,N_1549);
and U2708 (N_2708,N_1511,N_1687);
nand U2709 (N_2709,N_1814,N_1383);
and U2710 (N_2710,N_1482,N_1610);
nor U2711 (N_2711,N_1998,N_1529);
nor U2712 (N_2712,N_1159,N_1440);
or U2713 (N_2713,N_1246,N_1092);
and U2714 (N_2714,N_1843,N_1252);
and U2715 (N_2715,N_1964,N_1987);
and U2716 (N_2716,N_1600,N_1637);
and U2717 (N_2717,N_1670,N_1332);
nand U2718 (N_2718,N_1422,N_1895);
nor U2719 (N_2719,N_1565,N_1367);
and U2720 (N_2720,N_1746,N_1473);
nand U2721 (N_2721,N_1611,N_1111);
or U2722 (N_2722,N_1952,N_1965);
nand U2723 (N_2723,N_1836,N_1937);
nand U2724 (N_2724,N_1281,N_1548);
or U2725 (N_2725,N_1815,N_1576);
nand U2726 (N_2726,N_1898,N_1212);
or U2727 (N_2727,N_1289,N_1225);
xnor U2728 (N_2728,N_1461,N_1116);
xnor U2729 (N_2729,N_1809,N_1872);
and U2730 (N_2730,N_1630,N_1026);
xor U2731 (N_2731,N_1633,N_1777);
or U2732 (N_2732,N_1344,N_1741);
or U2733 (N_2733,N_1476,N_1824);
and U2734 (N_2734,N_1867,N_1245);
nand U2735 (N_2735,N_1073,N_1133);
xor U2736 (N_2736,N_1297,N_1137);
nor U2737 (N_2737,N_1741,N_1638);
nor U2738 (N_2738,N_1822,N_1824);
and U2739 (N_2739,N_1501,N_1630);
or U2740 (N_2740,N_1171,N_1194);
and U2741 (N_2741,N_1833,N_1957);
or U2742 (N_2742,N_1825,N_1079);
or U2743 (N_2743,N_1650,N_1287);
nor U2744 (N_2744,N_1440,N_1413);
nor U2745 (N_2745,N_1679,N_1231);
or U2746 (N_2746,N_1235,N_1736);
nand U2747 (N_2747,N_1890,N_1658);
xor U2748 (N_2748,N_1029,N_1792);
nand U2749 (N_2749,N_1093,N_1529);
or U2750 (N_2750,N_1555,N_1389);
nand U2751 (N_2751,N_1080,N_1471);
and U2752 (N_2752,N_1127,N_1088);
and U2753 (N_2753,N_1437,N_1001);
nand U2754 (N_2754,N_1003,N_1730);
or U2755 (N_2755,N_1695,N_1529);
nand U2756 (N_2756,N_1749,N_1756);
nand U2757 (N_2757,N_1426,N_1139);
and U2758 (N_2758,N_1330,N_1664);
xnor U2759 (N_2759,N_1503,N_1670);
and U2760 (N_2760,N_1832,N_1769);
nand U2761 (N_2761,N_1159,N_1774);
or U2762 (N_2762,N_1120,N_1578);
nand U2763 (N_2763,N_1556,N_1428);
and U2764 (N_2764,N_1955,N_1220);
nand U2765 (N_2765,N_1093,N_1460);
and U2766 (N_2766,N_1762,N_1552);
nor U2767 (N_2767,N_1194,N_1516);
nand U2768 (N_2768,N_1234,N_1473);
or U2769 (N_2769,N_1141,N_1179);
nand U2770 (N_2770,N_1572,N_1385);
and U2771 (N_2771,N_1724,N_1755);
nand U2772 (N_2772,N_1567,N_1403);
and U2773 (N_2773,N_1154,N_1568);
nor U2774 (N_2774,N_1768,N_1500);
nor U2775 (N_2775,N_1934,N_1867);
nand U2776 (N_2776,N_1684,N_1808);
nand U2777 (N_2777,N_1266,N_1451);
nor U2778 (N_2778,N_1035,N_1181);
and U2779 (N_2779,N_1505,N_1630);
nor U2780 (N_2780,N_1793,N_1460);
xnor U2781 (N_2781,N_1822,N_1037);
and U2782 (N_2782,N_1687,N_1780);
nand U2783 (N_2783,N_1897,N_1333);
nand U2784 (N_2784,N_1823,N_1489);
and U2785 (N_2785,N_1964,N_1668);
or U2786 (N_2786,N_1778,N_1285);
or U2787 (N_2787,N_1066,N_1145);
or U2788 (N_2788,N_1766,N_1042);
nor U2789 (N_2789,N_1824,N_1612);
nor U2790 (N_2790,N_1617,N_1787);
nor U2791 (N_2791,N_1017,N_1133);
or U2792 (N_2792,N_1070,N_1512);
nor U2793 (N_2793,N_1903,N_1040);
nor U2794 (N_2794,N_1789,N_1844);
nand U2795 (N_2795,N_1126,N_1791);
or U2796 (N_2796,N_1753,N_1217);
or U2797 (N_2797,N_1753,N_1102);
xor U2798 (N_2798,N_1992,N_1460);
or U2799 (N_2799,N_1631,N_1715);
nand U2800 (N_2800,N_1118,N_1218);
and U2801 (N_2801,N_1652,N_1528);
or U2802 (N_2802,N_1990,N_1274);
or U2803 (N_2803,N_1967,N_1954);
nor U2804 (N_2804,N_1036,N_1248);
nand U2805 (N_2805,N_1111,N_1141);
and U2806 (N_2806,N_1693,N_1729);
or U2807 (N_2807,N_1608,N_1261);
nand U2808 (N_2808,N_1118,N_1400);
nor U2809 (N_2809,N_1879,N_1752);
and U2810 (N_2810,N_1993,N_1306);
nand U2811 (N_2811,N_1904,N_1760);
nor U2812 (N_2812,N_1808,N_1502);
nand U2813 (N_2813,N_1595,N_1741);
nand U2814 (N_2814,N_1134,N_1789);
and U2815 (N_2815,N_1755,N_1199);
nor U2816 (N_2816,N_1854,N_1378);
nand U2817 (N_2817,N_1205,N_1314);
nand U2818 (N_2818,N_1591,N_1644);
and U2819 (N_2819,N_1276,N_1731);
or U2820 (N_2820,N_1831,N_1410);
or U2821 (N_2821,N_1150,N_1875);
and U2822 (N_2822,N_1019,N_1250);
nor U2823 (N_2823,N_1852,N_1851);
and U2824 (N_2824,N_1809,N_1758);
or U2825 (N_2825,N_1741,N_1951);
nand U2826 (N_2826,N_1129,N_1420);
nand U2827 (N_2827,N_1159,N_1025);
nand U2828 (N_2828,N_1073,N_1213);
xnor U2829 (N_2829,N_1826,N_1957);
nor U2830 (N_2830,N_1629,N_1653);
nor U2831 (N_2831,N_1213,N_1804);
nand U2832 (N_2832,N_1754,N_1187);
and U2833 (N_2833,N_1724,N_1801);
or U2834 (N_2834,N_1199,N_1923);
or U2835 (N_2835,N_1901,N_1461);
or U2836 (N_2836,N_1808,N_1313);
nand U2837 (N_2837,N_1032,N_1858);
and U2838 (N_2838,N_1056,N_1208);
or U2839 (N_2839,N_1382,N_1441);
or U2840 (N_2840,N_1446,N_1139);
or U2841 (N_2841,N_1171,N_1296);
nand U2842 (N_2842,N_1647,N_1461);
nand U2843 (N_2843,N_1120,N_1379);
nand U2844 (N_2844,N_1240,N_1244);
nand U2845 (N_2845,N_1119,N_1943);
nor U2846 (N_2846,N_1876,N_1113);
or U2847 (N_2847,N_1513,N_1633);
or U2848 (N_2848,N_1341,N_1311);
and U2849 (N_2849,N_1539,N_1026);
and U2850 (N_2850,N_1885,N_1706);
or U2851 (N_2851,N_1912,N_1053);
or U2852 (N_2852,N_1973,N_1398);
nor U2853 (N_2853,N_1278,N_1877);
nand U2854 (N_2854,N_1962,N_1502);
nor U2855 (N_2855,N_1106,N_1581);
or U2856 (N_2856,N_1533,N_1148);
or U2857 (N_2857,N_1885,N_1894);
and U2858 (N_2858,N_1759,N_1045);
nor U2859 (N_2859,N_1442,N_1257);
nand U2860 (N_2860,N_1154,N_1908);
nor U2861 (N_2861,N_1108,N_1532);
nand U2862 (N_2862,N_1839,N_1089);
or U2863 (N_2863,N_1102,N_1570);
and U2864 (N_2864,N_1923,N_1670);
nor U2865 (N_2865,N_1606,N_1814);
nand U2866 (N_2866,N_1403,N_1528);
or U2867 (N_2867,N_1601,N_1458);
nand U2868 (N_2868,N_1145,N_1433);
nor U2869 (N_2869,N_1395,N_1942);
and U2870 (N_2870,N_1861,N_1889);
and U2871 (N_2871,N_1767,N_1479);
and U2872 (N_2872,N_1527,N_1979);
nand U2873 (N_2873,N_1627,N_1780);
and U2874 (N_2874,N_1022,N_1978);
and U2875 (N_2875,N_1624,N_1293);
and U2876 (N_2876,N_1799,N_1550);
xor U2877 (N_2877,N_1654,N_1428);
nor U2878 (N_2878,N_1661,N_1711);
nor U2879 (N_2879,N_1539,N_1661);
or U2880 (N_2880,N_1463,N_1550);
nand U2881 (N_2881,N_1984,N_1459);
or U2882 (N_2882,N_1592,N_1904);
nor U2883 (N_2883,N_1172,N_1394);
and U2884 (N_2884,N_1021,N_1188);
nand U2885 (N_2885,N_1869,N_1562);
or U2886 (N_2886,N_1508,N_1360);
and U2887 (N_2887,N_1476,N_1224);
nand U2888 (N_2888,N_1227,N_1453);
nand U2889 (N_2889,N_1630,N_1112);
nor U2890 (N_2890,N_1174,N_1926);
and U2891 (N_2891,N_1531,N_1445);
and U2892 (N_2892,N_1118,N_1998);
nand U2893 (N_2893,N_1456,N_1889);
nor U2894 (N_2894,N_1162,N_1920);
and U2895 (N_2895,N_1417,N_1947);
nand U2896 (N_2896,N_1170,N_1503);
nand U2897 (N_2897,N_1955,N_1350);
nand U2898 (N_2898,N_1313,N_1185);
nand U2899 (N_2899,N_1802,N_1868);
or U2900 (N_2900,N_1955,N_1688);
or U2901 (N_2901,N_1931,N_1309);
and U2902 (N_2902,N_1750,N_1339);
and U2903 (N_2903,N_1704,N_1915);
or U2904 (N_2904,N_1002,N_1416);
nor U2905 (N_2905,N_1831,N_1173);
or U2906 (N_2906,N_1544,N_1439);
nand U2907 (N_2907,N_1871,N_1284);
nand U2908 (N_2908,N_1349,N_1762);
or U2909 (N_2909,N_1136,N_1139);
or U2910 (N_2910,N_1886,N_1672);
and U2911 (N_2911,N_1529,N_1766);
nand U2912 (N_2912,N_1478,N_1509);
or U2913 (N_2913,N_1466,N_1422);
nor U2914 (N_2914,N_1122,N_1021);
nand U2915 (N_2915,N_1278,N_1699);
nand U2916 (N_2916,N_1415,N_1109);
nor U2917 (N_2917,N_1607,N_1755);
or U2918 (N_2918,N_1845,N_1674);
or U2919 (N_2919,N_1788,N_1685);
or U2920 (N_2920,N_1326,N_1042);
nand U2921 (N_2921,N_1002,N_1140);
nand U2922 (N_2922,N_1771,N_1101);
and U2923 (N_2923,N_1323,N_1716);
and U2924 (N_2924,N_1109,N_1130);
and U2925 (N_2925,N_1512,N_1355);
or U2926 (N_2926,N_1546,N_1634);
nand U2927 (N_2927,N_1672,N_1729);
and U2928 (N_2928,N_1323,N_1264);
and U2929 (N_2929,N_1890,N_1206);
and U2930 (N_2930,N_1800,N_1458);
nor U2931 (N_2931,N_1968,N_1401);
or U2932 (N_2932,N_1015,N_1112);
or U2933 (N_2933,N_1990,N_1397);
nor U2934 (N_2934,N_1788,N_1737);
nand U2935 (N_2935,N_1903,N_1750);
nand U2936 (N_2936,N_1529,N_1440);
xor U2937 (N_2937,N_1826,N_1265);
or U2938 (N_2938,N_1254,N_1217);
or U2939 (N_2939,N_1462,N_1232);
and U2940 (N_2940,N_1530,N_1441);
or U2941 (N_2941,N_1528,N_1010);
and U2942 (N_2942,N_1528,N_1573);
nand U2943 (N_2943,N_1657,N_1857);
nor U2944 (N_2944,N_1945,N_1581);
or U2945 (N_2945,N_1623,N_1417);
or U2946 (N_2946,N_1463,N_1841);
nand U2947 (N_2947,N_1523,N_1007);
and U2948 (N_2948,N_1456,N_1795);
or U2949 (N_2949,N_1051,N_1135);
and U2950 (N_2950,N_1535,N_1682);
or U2951 (N_2951,N_1941,N_1427);
or U2952 (N_2952,N_1470,N_1030);
or U2953 (N_2953,N_1272,N_1304);
and U2954 (N_2954,N_1873,N_1983);
nor U2955 (N_2955,N_1669,N_1978);
nor U2956 (N_2956,N_1199,N_1482);
nand U2957 (N_2957,N_1089,N_1368);
and U2958 (N_2958,N_1327,N_1070);
and U2959 (N_2959,N_1036,N_1412);
nor U2960 (N_2960,N_1033,N_1864);
or U2961 (N_2961,N_1732,N_1019);
or U2962 (N_2962,N_1961,N_1607);
or U2963 (N_2963,N_1201,N_1137);
and U2964 (N_2964,N_1485,N_1112);
nor U2965 (N_2965,N_1659,N_1021);
nand U2966 (N_2966,N_1010,N_1956);
and U2967 (N_2967,N_1732,N_1100);
and U2968 (N_2968,N_1315,N_1273);
or U2969 (N_2969,N_1330,N_1181);
or U2970 (N_2970,N_1411,N_1774);
or U2971 (N_2971,N_1199,N_1776);
and U2972 (N_2972,N_1022,N_1723);
nand U2973 (N_2973,N_1681,N_1522);
and U2974 (N_2974,N_1982,N_1956);
nand U2975 (N_2975,N_1195,N_1762);
nor U2976 (N_2976,N_1672,N_1430);
nor U2977 (N_2977,N_1676,N_1111);
and U2978 (N_2978,N_1112,N_1957);
or U2979 (N_2979,N_1612,N_1453);
or U2980 (N_2980,N_1098,N_1365);
and U2981 (N_2981,N_1257,N_1971);
and U2982 (N_2982,N_1264,N_1901);
and U2983 (N_2983,N_1148,N_1721);
or U2984 (N_2984,N_1397,N_1278);
nor U2985 (N_2985,N_1041,N_1691);
or U2986 (N_2986,N_1833,N_1229);
or U2987 (N_2987,N_1533,N_1575);
or U2988 (N_2988,N_1140,N_1694);
and U2989 (N_2989,N_1419,N_1929);
and U2990 (N_2990,N_1308,N_1953);
or U2991 (N_2991,N_1806,N_1984);
nand U2992 (N_2992,N_1502,N_1125);
and U2993 (N_2993,N_1107,N_1312);
nor U2994 (N_2994,N_1365,N_1678);
nor U2995 (N_2995,N_1933,N_1764);
or U2996 (N_2996,N_1796,N_1633);
and U2997 (N_2997,N_1014,N_1215);
or U2998 (N_2998,N_1437,N_1615);
nand U2999 (N_2999,N_1806,N_1534);
and UO_0 (O_0,N_2137,N_2681);
nor UO_1 (O_1,N_2676,N_2506);
nor UO_2 (O_2,N_2135,N_2818);
nand UO_3 (O_3,N_2330,N_2193);
nor UO_4 (O_4,N_2656,N_2958);
or UO_5 (O_5,N_2232,N_2071);
nand UO_6 (O_6,N_2194,N_2192);
nand UO_7 (O_7,N_2225,N_2337);
nor UO_8 (O_8,N_2566,N_2738);
nor UO_9 (O_9,N_2186,N_2074);
and UO_10 (O_10,N_2978,N_2085);
nand UO_11 (O_11,N_2065,N_2590);
xnor UO_12 (O_12,N_2298,N_2254);
nor UO_13 (O_13,N_2576,N_2423);
or UO_14 (O_14,N_2712,N_2018);
or UO_15 (O_15,N_2104,N_2737);
or UO_16 (O_16,N_2495,N_2341);
or UO_17 (O_17,N_2468,N_2498);
and UO_18 (O_18,N_2526,N_2094);
nor UO_19 (O_19,N_2106,N_2770);
nand UO_20 (O_20,N_2392,N_2711);
nor UO_21 (O_21,N_2642,N_2872);
and UO_22 (O_22,N_2101,N_2521);
nand UO_23 (O_23,N_2155,N_2285);
nor UO_24 (O_24,N_2683,N_2374);
nand UO_25 (O_25,N_2952,N_2512);
nor UO_26 (O_26,N_2722,N_2785);
and UO_27 (O_27,N_2097,N_2114);
nor UO_28 (O_28,N_2763,N_2025);
and UO_29 (O_29,N_2125,N_2587);
nand UO_30 (O_30,N_2052,N_2427);
nor UO_31 (O_31,N_2593,N_2312);
and UO_32 (O_32,N_2405,N_2203);
nand UO_33 (O_33,N_2629,N_2791);
nand UO_34 (O_34,N_2489,N_2633);
or UO_35 (O_35,N_2527,N_2202);
or UO_36 (O_36,N_2724,N_2670);
and UO_37 (O_37,N_2229,N_2607);
nor UO_38 (O_38,N_2242,N_2180);
and UO_39 (O_39,N_2934,N_2517);
nand UO_40 (O_40,N_2462,N_2914);
nor UO_41 (O_41,N_2831,N_2128);
or UO_42 (O_42,N_2212,N_2231);
xnor UO_43 (O_43,N_2136,N_2664);
and UO_44 (O_44,N_2451,N_2222);
nor UO_45 (O_45,N_2523,N_2956);
nand UO_46 (O_46,N_2378,N_2399);
and UO_47 (O_47,N_2145,N_2649);
or UO_48 (O_48,N_2033,N_2695);
nand UO_49 (O_49,N_2532,N_2460);
nand UO_50 (O_50,N_2141,N_2430);
nor UO_51 (O_51,N_2111,N_2256);
xor UO_52 (O_52,N_2009,N_2979);
nand UO_53 (O_53,N_2339,N_2448);
or UO_54 (O_54,N_2588,N_2385);
and UO_55 (O_55,N_2048,N_2159);
nand UO_56 (O_56,N_2343,N_2581);
nand UO_57 (O_57,N_2240,N_2515);
and UO_58 (O_58,N_2239,N_2019);
and UO_59 (O_59,N_2181,N_2665);
nor UO_60 (O_60,N_2214,N_2003);
or UO_61 (O_61,N_2975,N_2334);
nand UO_62 (O_62,N_2046,N_2945);
or UO_63 (O_63,N_2736,N_2432);
nand UO_64 (O_64,N_2062,N_2210);
or UO_65 (O_65,N_2568,N_2098);
nor UO_66 (O_66,N_2936,N_2319);
nand UO_67 (O_67,N_2497,N_2929);
nand UO_68 (O_68,N_2821,N_2290);
nand UO_69 (O_69,N_2361,N_2227);
or UO_70 (O_70,N_2802,N_2316);
nand UO_71 (O_71,N_2200,N_2351);
or UO_72 (O_72,N_2959,N_2579);
and UO_73 (O_73,N_2093,N_2038);
nor UO_74 (O_74,N_2031,N_2260);
nor UO_75 (O_75,N_2733,N_2209);
and UO_76 (O_76,N_2977,N_2863);
nor UO_77 (O_77,N_2262,N_2322);
or UO_78 (O_78,N_2966,N_2331);
or UO_79 (O_79,N_2798,N_2981);
and UO_80 (O_80,N_2621,N_2589);
and UO_81 (O_81,N_2586,N_2610);
nor UO_82 (O_82,N_2414,N_2400);
or UO_83 (O_83,N_2110,N_2190);
and UO_84 (O_84,N_2205,N_2546);
nor UO_85 (O_85,N_2467,N_2769);
or UO_86 (O_86,N_2648,N_2848);
and UO_87 (O_87,N_2404,N_2620);
and UO_88 (O_88,N_2483,N_2698);
nor UO_89 (O_89,N_2756,N_2974);
nor UO_90 (O_90,N_2236,N_2369);
nand UO_91 (O_91,N_2021,N_2650);
and UO_92 (O_92,N_2069,N_2353);
nand UO_93 (O_93,N_2707,N_2365);
xor UO_94 (O_94,N_2571,N_2187);
and UO_95 (O_95,N_2117,N_2286);
and UO_96 (O_96,N_2504,N_2158);
and UO_97 (O_97,N_2324,N_2268);
and UO_98 (O_98,N_2016,N_2655);
or UO_99 (O_99,N_2360,N_2790);
or UO_100 (O_100,N_2816,N_2538);
nand UO_101 (O_101,N_2051,N_2058);
and UO_102 (O_102,N_2191,N_2425);
nor UO_103 (O_103,N_2255,N_2464);
nand UO_104 (O_104,N_2728,N_2803);
nand UO_105 (O_105,N_2600,N_2854);
nand UO_106 (O_106,N_2643,N_2787);
nand UO_107 (O_107,N_2927,N_2134);
and UO_108 (O_108,N_2456,N_2053);
and UO_109 (O_109,N_2109,N_2118);
xor UO_110 (O_110,N_2049,N_2596);
or UO_111 (O_111,N_2431,N_2948);
and UO_112 (O_112,N_2772,N_2985);
and UO_113 (O_113,N_2257,N_2674);
or UO_114 (O_114,N_2663,N_2710);
or UO_115 (O_115,N_2921,N_2638);
or UO_116 (O_116,N_2799,N_2562);
or UO_117 (O_117,N_2296,N_2627);
nand UO_118 (O_118,N_2548,N_2153);
nor UO_119 (O_119,N_2869,N_2394);
nor UO_120 (O_120,N_2716,N_2315);
and UO_121 (O_121,N_2631,N_2154);
or UO_122 (O_122,N_2107,N_2905);
nand UO_123 (O_123,N_2529,N_2366);
or UO_124 (O_124,N_2918,N_2499);
or UO_125 (O_125,N_2199,N_2513);
nand UO_126 (O_126,N_2303,N_2639);
nand UO_127 (O_127,N_2265,N_2352);
nand UO_128 (O_128,N_2359,N_2358);
nand UO_129 (O_129,N_2563,N_2878);
nor UO_130 (O_130,N_2595,N_2332);
nand UO_131 (O_131,N_2955,N_2026);
nand UO_132 (O_132,N_2865,N_2278);
and UO_133 (O_133,N_2604,N_2856);
and UO_134 (O_134,N_2625,N_2687);
xor UO_135 (O_135,N_2133,N_2689);
and UO_136 (O_136,N_2029,N_2349);
nand UO_137 (O_137,N_2694,N_2731);
or UO_138 (O_138,N_2807,N_2441);
and UO_139 (O_139,N_2237,N_2357);
nor UO_140 (O_140,N_2690,N_2808);
or UO_141 (O_141,N_2218,N_2273);
nor UO_142 (O_142,N_2761,N_2552);
xnor UO_143 (O_143,N_2091,N_2701);
nand UO_144 (O_144,N_2006,N_2647);
and UO_145 (O_145,N_2165,N_2535);
or UO_146 (O_146,N_2252,N_2473);
and UO_147 (O_147,N_2061,N_2164);
or UO_148 (O_148,N_2868,N_2894);
or UO_149 (O_149,N_2904,N_2614);
nand UO_150 (O_150,N_2853,N_2264);
and UO_151 (O_151,N_2304,N_2082);
and UO_152 (O_152,N_2188,N_2602);
xnor UO_153 (O_153,N_2245,N_2951);
xnor UO_154 (O_154,N_2024,N_2911);
nand UO_155 (O_155,N_2603,N_2491);
xnor UO_156 (O_156,N_2741,N_2962);
and UO_157 (O_157,N_2308,N_2395);
or UO_158 (O_158,N_2823,N_2553);
and UO_159 (O_159,N_2470,N_2105);
nor UO_160 (O_160,N_2015,N_2980);
nor UO_161 (O_161,N_2348,N_2855);
nand UO_162 (O_162,N_2534,N_2204);
nand UO_163 (O_163,N_2801,N_2100);
and UO_164 (O_164,N_2311,N_2993);
nand UO_165 (O_165,N_2703,N_2176);
nand UO_166 (O_166,N_2510,N_2524);
and UO_167 (O_167,N_2465,N_2671);
or UO_168 (O_168,N_2350,N_2411);
xnor UO_169 (O_169,N_2035,N_2652);
nor UO_170 (O_170,N_2897,N_2679);
nor UO_171 (O_171,N_2857,N_2909);
nand UO_172 (O_172,N_2879,N_2577);
nor UO_173 (O_173,N_2615,N_2088);
nor UO_174 (O_174,N_2640,N_2384);
nor UO_175 (O_175,N_2752,N_2197);
and UO_176 (O_176,N_2055,N_2208);
xnor UO_177 (O_177,N_2436,N_2090);
nand UO_178 (O_178,N_2368,N_2965);
or UO_179 (O_179,N_2266,N_2333);
and UO_180 (O_180,N_2380,N_2813);
nand UO_181 (O_181,N_2480,N_2221);
nor UO_182 (O_182,N_2444,N_2281);
or UO_183 (O_183,N_2377,N_2001);
nor UO_184 (O_184,N_2140,N_2887);
or UO_185 (O_185,N_2833,N_2626);
and UO_186 (O_186,N_2129,N_2166);
nand UO_187 (O_187,N_2259,N_2344);
or UO_188 (O_188,N_2036,N_2463);
nor UO_189 (O_189,N_2811,N_2834);
nor UO_190 (O_190,N_2277,N_2042);
nor UO_191 (O_191,N_2836,N_2215);
and UO_192 (O_192,N_2528,N_2178);
xnor UO_193 (O_193,N_2820,N_2922);
or UO_194 (O_194,N_2745,N_2250);
nor UO_195 (O_195,N_2623,N_2138);
nand UO_196 (O_196,N_2500,N_2556);
and UO_197 (O_197,N_2906,N_2835);
nand UO_198 (O_198,N_2119,N_2075);
nor UO_199 (O_199,N_2949,N_2641);
xor UO_200 (O_200,N_2244,N_2605);
or UO_201 (O_201,N_2781,N_2383);
nor UO_202 (O_202,N_2850,N_2270);
nand UO_203 (O_203,N_2447,N_2433);
nand UO_204 (O_204,N_2597,N_2880);
nand UO_205 (O_205,N_2907,N_2081);
or UO_206 (O_206,N_2540,N_2459);
nor UO_207 (O_207,N_2492,N_2327);
nor UO_208 (O_208,N_2990,N_2709);
nor UO_209 (O_209,N_2825,N_2890);
xor UO_210 (O_210,N_2828,N_2788);
nor UO_211 (O_211,N_2410,N_2829);
nor UO_212 (O_212,N_2372,N_2446);
nand UO_213 (O_213,N_2452,N_2940);
or UO_214 (O_214,N_2219,N_2428);
nor UO_215 (O_215,N_2066,N_2345);
nor UO_216 (O_216,N_2485,N_2832);
nor UO_217 (O_217,N_2809,N_2735);
or UO_218 (O_218,N_2415,N_2937);
or UO_219 (O_219,N_2987,N_2892);
or UO_220 (O_220,N_2908,N_2654);
nand UO_221 (O_221,N_2582,N_2401);
nor UO_222 (O_222,N_2971,N_2935);
and UO_223 (O_223,N_2010,N_2957);
nor UO_224 (O_224,N_2750,N_2926);
and UO_225 (O_225,N_2037,N_2874);
nand UO_226 (O_226,N_2618,N_2749);
nor UO_227 (O_227,N_2005,N_2995);
nor UO_228 (O_228,N_2142,N_2336);
nor UO_229 (O_229,N_2913,N_2784);
and UO_230 (O_230,N_2122,N_2680);
or UO_231 (O_231,N_2915,N_2347);
nor UO_232 (O_232,N_2338,N_2841);
and UO_233 (O_233,N_2613,N_2354);
nor UO_234 (O_234,N_2891,N_2078);
or UO_235 (O_235,N_2877,N_2849);
or UO_236 (O_236,N_2175,N_2697);
and UO_237 (O_237,N_2783,N_2509);
and UO_238 (O_238,N_2184,N_2757);
and UO_239 (O_239,N_2771,N_2403);
or UO_240 (O_240,N_2216,N_2466);
nor UO_241 (O_241,N_2050,N_2173);
nand UO_242 (O_242,N_2541,N_2557);
nand UO_243 (O_243,N_2007,N_2148);
or UO_244 (O_244,N_2653,N_2246);
and UO_245 (O_245,N_2634,N_2668);
nor UO_246 (O_246,N_2660,N_2022);
and UO_247 (O_247,N_2764,N_2840);
and UO_248 (O_248,N_2407,N_2476);
nor UO_249 (O_249,N_2207,N_2773);
or UO_250 (O_250,N_2041,N_2000);
and UO_251 (O_251,N_2691,N_2282);
nor UO_252 (O_252,N_2012,N_2941);
and UO_253 (O_253,N_2726,N_2651);
nor UO_254 (O_254,N_2559,N_2008);
or UO_255 (O_255,N_2560,N_2233);
nor UO_256 (O_256,N_2249,N_2885);
and UO_257 (O_257,N_2686,N_2531);
and UO_258 (O_258,N_2973,N_2481);
nor UO_259 (O_259,N_2040,N_2964);
or UO_260 (O_260,N_2706,N_2174);
or UO_261 (O_261,N_2434,N_2858);
nand UO_262 (O_262,N_2299,N_2606);
or UO_263 (O_263,N_2822,N_2371);
nor UO_264 (O_264,N_2472,N_2326);
or UO_265 (O_265,N_2954,N_2744);
nand UO_266 (O_266,N_2873,N_2393);
and UO_267 (O_267,N_2083,N_2886);
nor UO_268 (O_268,N_2211,N_2947);
and UO_269 (O_269,N_2039,N_2149);
nor UO_270 (O_270,N_2126,N_2599);
nand UO_271 (O_271,N_2253,N_2759);
nand UO_272 (O_272,N_2309,N_2542);
xnor UO_273 (O_273,N_2646,N_2429);
and UO_274 (O_274,N_2131,N_2121);
nor UO_275 (O_275,N_2213,N_2340);
nand UO_276 (O_276,N_2346,N_2002);
or UO_277 (O_277,N_2147,N_2944);
or UO_278 (O_278,N_2310,N_2056);
or UO_279 (O_279,N_2778,N_2043);
or UO_280 (O_280,N_2505,N_2496);
or UO_281 (O_281,N_2682,N_2398);
nand UO_282 (O_282,N_2223,N_2087);
and UO_283 (O_283,N_2748,N_2774);
nor UO_284 (O_284,N_2846,N_2437);
and UO_285 (O_285,N_2960,N_2765);
or UO_286 (O_286,N_2684,N_2457);
nor UO_287 (O_287,N_2795,N_2930);
and UO_288 (O_288,N_2901,N_2899);
nor UO_289 (O_289,N_2068,N_2157);
and UO_290 (O_290,N_2426,N_2617);
and UO_291 (O_291,N_2842,N_2072);
and UO_292 (O_292,N_2389,N_2747);
and UO_293 (O_293,N_2079,N_2185);
nand UO_294 (O_294,N_2705,N_2775);
and UO_295 (O_295,N_2814,N_2720);
nor UO_296 (O_296,N_2673,N_2171);
nor UO_297 (O_297,N_2102,N_2287);
or UO_298 (O_298,N_2696,N_2408);
nor UO_299 (O_299,N_2659,N_2819);
and UO_300 (O_300,N_2279,N_2030);
nor UO_301 (O_301,N_2804,N_2946);
nand UO_302 (O_302,N_2516,N_2362);
and UO_303 (O_303,N_2983,N_2969);
nand UO_304 (O_304,N_2047,N_2989);
nor UO_305 (O_305,N_2230,N_2440);
and UO_306 (O_306,N_2866,N_2297);
or UO_307 (O_307,N_2723,N_2363);
nor UO_308 (O_308,N_2932,N_2045);
or UO_309 (O_309,N_2306,N_2555);
or UO_310 (O_310,N_2396,N_2511);
or UO_311 (O_311,N_2044,N_2013);
or UO_312 (O_312,N_2730,N_2554);
nor UO_313 (O_313,N_2616,N_2902);
and UO_314 (O_314,N_2851,N_2439);
or UO_315 (O_315,N_2537,N_2567);
and UO_316 (O_316,N_2972,N_2089);
nor UO_317 (O_317,N_2386,N_2424);
and UO_318 (O_318,N_2817,N_2170);
and UO_319 (O_319,N_2514,N_2875);
or UO_320 (O_320,N_2261,N_2220);
or UO_321 (O_321,N_2997,N_2718);
and UO_322 (O_322,N_2275,N_2307);
or UO_323 (O_323,N_2291,N_2120);
nor UO_324 (O_324,N_2786,N_2217);
nand UO_325 (O_325,N_2637,N_2238);
and UO_326 (O_326,N_2084,N_2961);
or UO_327 (O_327,N_2067,N_2898);
or UO_328 (O_328,N_2561,N_2151);
nand UO_329 (O_329,N_2421,N_2318);
nand UO_330 (O_330,N_2234,N_2017);
nand UO_331 (O_331,N_2494,N_2370);
or UO_332 (O_332,N_2413,N_2475);
nand UO_333 (O_333,N_2267,N_2520);
and UO_334 (O_334,N_2924,N_2584);
and UO_335 (O_335,N_2477,N_2367);
or UO_336 (O_336,N_2438,N_2645);
nand UO_337 (O_337,N_2881,N_2487);
nor UO_338 (O_338,N_2753,N_2984);
and UO_339 (O_339,N_2806,N_2533);
nor UO_340 (O_340,N_2417,N_2488);
or UO_341 (O_341,N_2177,N_2702);
or UO_342 (O_342,N_2076,N_2796);
nand UO_343 (O_343,N_2355,N_2635);
or UO_344 (O_344,N_2580,N_2172);
nor UO_345 (O_345,N_2550,N_2493);
and UO_346 (O_346,N_2740,N_2843);
nand UO_347 (O_347,N_2910,N_2800);
or UO_348 (O_348,N_2592,N_2143);
xor UO_349 (O_349,N_2864,N_2382);
or UO_350 (O_350,N_2391,N_2416);
nor UO_351 (O_351,N_2073,N_2920);
and UO_352 (O_352,N_2996,N_2057);
or UO_353 (O_353,N_2601,N_2574);
and UO_354 (O_354,N_2195,N_2675);
nor UO_355 (O_355,N_2127,N_2742);
and UO_356 (O_356,N_2402,N_2471);
or UO_357 (O_357,N_2096,N_2323);
xor UO_358 (O_358,N_2667,N_2305);
nor UO_359 (O_359,N_2876,N_2992);
and UO_360 (O_360,N_2182,N_2445);
and UO_361 (O_361,N_2685,N_2179);
nor UO_362 (O_362,N_2302,N_2274);
nand UO_363 (O_363,N_2789,N_2630);
or UO_364 (O_364,N_2435,N_2280);
nand UO_365 (O_365,N_2294,N_2912);
nor UO_366 (O_366,N_2168,N_2688);
and UO_367 (O_367,N_2183,N_2976);
or UO_368 (O_368,N_2794,N_2525);
nor UO_369 (O_369,N_2612,N_2070);
nor UO_370 (O_370,N_2004,N_2867);
and UO_371 (O_371,N_2609,N_2241);
nand UO_372 (O_372,N_2314,N_2486);
nor UO_373 (O_373,N_2717,N_2064);
or UO_374 (O_374,N_2490,N_2708);
xor UO_375 (O_375,N_2461,N_2518);
xor UO_376 (O_376,N_2263,N_2719);
and UO_377 (O_377,N_2713,N_2086);
nand UO_378 (O_378,N_2160,N_2206);
nand UO_379 (O_379,N_2953,N_2228);
nor UO_380 (O_380,N_2727,N_2999);
or UO_381 (O_381,N_2545,N_2011);
and UO_382 (O_382,N_2732,N_2276);
and UO_383 (O_383,N_2739,N_2569);
or UO_384 (O_384,N_2196,N_2888);
nand UO_385 (O_385,N_2201,N_2845);
nor UO_386 (O_386,N_2988,N_2130);
and UO_387 (O_387,N_2839,N_2077);
and UO_388 (O_388,N_2636,N_2862);
and UO_389 (O_389,N_2743,N_2116);
or UO_390 (O_390,N_2916,N_2776);
nor UO_391 (O_391,N_2099,N_2295);
nand UO_392 (O_392,N_2700,N_2812);
nand UO_393 (O_393,N_2247,N_2933);
or UO_394 (O_394,N_2390,N_2805);
and UO_395 (O_395,N_2611,N_2450);
nand UO_396 (O_396,N_2939,N_2132);
nor UO_397 (O_397,N_2226,N_2883);
and UO_398 (O_398,N_2375,N_2925);
or UO_399 (O_399,N_2474,N_2054);
xnor UO_400 (O_400,N_2321,N_2028);
or UO_401 (O_401,N_2288,N_2289);
nor UO_402 (O_402,N_2669,N_2284);
nand UO_403 (O_403,N_2032,N_2942);
nand UO_404 (O_404,N_2469,N_2169);
nor UO_405 (O_405,N_2547,N_2189);
and UO_406 (O_406,N_2662,N_2292);
and UO_407 (O_407,N_2419,N_2558);
nand UO_408 (O_408,N_2248,N_2837);
and UO_409 (O_409,N_2591,N_2115);
and UO_410 (O_410,N_2139,N_2672);
or UO_411 (O_411,N_2815,N_2144);
xnor UO_412 (O_412,N_2658,N_2508);
or UO_413 (O_413,N_2824,N_2388);
and UO_414 (O_414,N_2725,N_2454);
and UO_415 (O_415,N_2420,N_2931);
or UO_416 (O_416,N_2826,N_2092);
nand UO_417 (O_417,N_2329,N_2146);
nor UO_418 (O_418,N_2755,N_2746);
or UO_419 (O_419,N_2994,N_2644);
nand UO_420 (O_420,N_2950,N_2986);
nand UO_421 (O_421,N_2301,N_2624);
or UO_422 (O_422,N_2585,N_2928);
nand UO_423 (O_423,N_2060,N_2564);
nor UO_424 (O_424,N_2870,N_2455);
and UO_425 (O_425,N_2838,N_2758);
and UO_426 (O_426,N_2243,N_2766);
nor UO_427 (O_427,N_2397,N_2572);
and UO_428 (O_428,N_2777,N_2573);
nor UO_429 (O_429,N_2721,N_2967);
nand UO_430 (O_430,N_2103,N_2608);
nor UO_431 (O_431,N_2714,N_2861);
or UO_432 (O_432,N_2543,N_2530);
xnor UO_433 (O_433,N_2412,N_2300);
and UO_434 (O_434,N_2484,N_2896);
nor UO_435 (O_435,N_2859,N_2998);
nand UO_436 (O_436,N_2482,N_2917);
nor UO_437 (O_437,N_2123,N_2903);
and UO_438 (O_438,N_2762,N_2991);
and UO_439 (O_439,N_2479,N_2751);
nor UO_440 (O_440,N_2968,N_2882);
and UO_441 (O_441,N_2871,N_2381);
nor UO_442 (O_442,N_2923,N_2293);
nor UO_443 (O_443,N_2113,N_2622);
nand UO_444 (O_444,N_2779,N_2023);
or UO_445 (O_445,N_2729,N_2224);
xor UO_446 (O_446,N_2442,N_2628);
nor UO_447 (O_447,N_2919,N_2889);
nand UO_448 (O_448,N_2379,N_2376);
nand UO_449 (O_449,N_2693,N_2269);
or UO_450 (O_450,N_2578,N_2124);
nor UO_451 (O_451,N_2666,N_2251);
nand UO_452 (O_452,N_2313,N_2830);
and UO_453 (O_453,N_2373,N_2320);
or UO_454 (O_454,N_2943,N_2443);
nor UO_455 (O_455,N_2059,N_2063);
or UO_456 (O_456,N_2768,N_2895);
nand UO_457 (O_457,N_2760,N_2317);
nor UO_458 (O_458,N_2792,N_2519);
nand UO_459 (O_459,N_2565,N_2271);
or UO_460 (O_460,N_2342,N_2478);
nor UO_461 (O_461,N_2235,N_2827);
nor UO_462 (O_462,N_2409,N_2551);
nand UO_463 (O_463,N_2156,N_2797);
and UO_464 (O_464,N_2162,N_2982);
and UO_465 (O_465,N_2938,N_2356);
nor UO_466 (O_466,N_2406,N_2014);
nor UO_467 (O_467,N_2844,N_2860);
or UO_468 (O_468,N_2893,N_2678);
or UO_469 (O_469,N_2422,N_2034);
nand UO_470 (O_470,N_2598,N_2198);
and UO_471 (O_471,N_2328,N_2364);
nor UO_472 (O_472,N_2549,N_2112);
xnor UO_473 (O_473,N_2501,N_2449);
nor UO_474 (O_474,N_2418,N_2900);
nand UO_475 (O_475,N_2522,N_2734);
and UO_476 (O_476,N_2583,N_2152);
nor UO_477 (O_477,N_2767,N_2325);
nand UO_478 (O_478,N_2335,N_2458);
nand UO_479 (O_479,N_2810,N_2027);
and UO_480 (O_480,N_2507,N_2163);
and UO_481 (O_481,N_2661,N_2632);
nor UO_482 (O_482,N_2847,N_2780);
and UO_483 (O_483,N_2536,N_2272);
and UO_484 (O_484,N_2704,N_2150);
or UO_485 (O_485,N_2970,N_2108);
or UO_486 (O_486,N_2619,N_2095);
or UO_487 (O_487,N_2539,N_2594);
and UO_488 (O_488,N_2258,N_2793);
and UO_489 (O_489,N_2167,N_2754);
and UO_490 (O_490,N_2544,N_2453);
nor UO_491 (O_491,N_2570,N_2692);
and UO_492 (O_492,N_2782,N_2699);
or UO_493 (O_493,N_2283,N_2080);
nand UO_494 (O_494,N_2657,N_2020);
or UO_495 (O_495,N_2884,N_2715);
nand UO_496 (O_496,N_2963,N_2852);
nor UO_497 (O_497,N_2161,N_2503);
xor UO_498 (O_498,N_2502,N_2677);
or UO_499 (O_499,N_2387,N_2575);
endmodule