module basic_500_3000_500_30_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_76,In_424);
or U1 (N_1,In_311,In_490);
nor U2 (N_2,In_419,In_427);
nand U3 (N_3,In_360,In_149);
or U4 (N_4,In_469,In_11);
nand U5 (N_5,In_335,In_162);
or U6 (N_6,In_24,In_275);
and U7 (N_7,In_414,In_60);
nor U8 (N_8,In_470,In_382);
xor U9 (N_9,In_242,In_172);
nand U10 (N_10,In_446,In_114);
nand U11 (N_11,In_347,In_411);
nand U12 (N_12,In_219,In_160);
xnor U13 (N_13,In_0,In_227);
or U14 (N_14,In_453,In_357);
nand U15 (N_15,In_75,In_237);
nand U16 (N_16,In_494,In_302);
nor U17 (N_17,In_452,In_273);
nor U18 (N_18,In_83,In_5);
and U19 (N_19,In_240,In_89);
xor U20 (N_20,In_66,In_194);
xor U21 (N_21,In_464,In_27);
nand U22 (N_22,In_284,In_256);
nand U23 (N_23,In_210,In_129);
xnor U24 (N_24,In_203,In_271);
and U25 (N_25,In_291,In_313);
and U26 (N_26,In_229,In_165);
nand U27 (N_27,In_393,In_394);
or U28 (N_28,In_163,In_383);
and U29 (N_29,In_95,In_14);
and U30 (N_30,In_475,In_22);
nor U31 (N_31,In_224,In_127);
or U32 (N_32,In_178,In_488);
nand U33 (N_33,In_23,In_111);
or U34 (N_34,In_140,In_230);
and U35 (N_35,In_344,In_78);
or U36 (N_36,In_496,In_159);
nand U37 (N_37,In_251,In_212);
nand U38 (N_38,In_186,In_417);
xnor U39 (N_39,In_4,In_118);
or U40 (N_40,In_231,In_450);
or U41 (N_41,In_290,In_216);
nand U42 (N_42,In_415,In_269);
nand U43 (N_43,In_405,In_312);
nor U44 (N_44,In_410,In_143);
xor U45 (N_45,In_443,In_9);
or U46 (N_46,In_45,In_305);
and U47 (N_47,In_130,In_385);
and U48 (N_48,In_119,In_479);
or U49 (N_49,In_396,In_377);
or U50 (N_50,In_117,In_183);
or U51 (N_51,In_218,In_461);
nor U52 (N_52,In_297,In_367);
and U53 (N_53,In_98,In_106);
or U54 (N_54,In_154,In_155);
and U55 (N_55,In_131,In_472);
xor U56 (N_56,In_59,In_190);
and U57 (N_57,In_128,In_21);
xor U58 (N_58,In_348,In_486);
nand U59 (N_59,In_198,In_199);
nand U60 (N_60,In_37,In_316);
xor U61 (N_61,In_380,In_105);
or U62 (N_62,In_18,In_327);
xor U63 (N_63,In_116,In_173);
or U64 (N_64,In_495,In_91);
nor U65 (N_65,In_293,In_179);
or U66 (N_66,In_425,In_402);
or U67 (N_67,In_152,In_191);
or U68 (N_68,In_192,In_341);
nor U69 (N_69,In_120,In_399);
xor U70 (N_70,In_362,In_221);
nand U71 (N_71,In_478,In_90);
nand U72 (N_72,In_384,In_351);
nand U73 (N_73,In_448,In_77);
xnor U74 (N_74,In_349,In_168);
nand U75 (N_75,In_426,In_28);
and U76 (N_76,In_79,In_233);
and U77 (N_77,In_338,In_94);
xor U78 (N_78,In_434,In_126);
xor U79 (N_79,In_325,In_264);
nor U80 (N_80,In_492,In_298);
xor U81 (N_81,In_54,In_304);
nand U82 (N_82,In_222,In_200);
nand U83 (N_83,In_93,In_65);
or U84 (N_84,In_401,In_47);
and U85 (N_85,In_343,In_436);
or U86 (N_86,In_39,In_403);
xor U87 (N_87,In_438,In_247);
nor U88 (N_88,In_70,In_205);
and U89 (N_89,In_96,In_404);
xor U90 (N_90,In_202,In_281);
nor U91 (N_91,In_13,In_487);
or U92 (N_92,In_225,In_337);
nor U93 (N_93,In_36,In_87);
xor U94 (N_94,In_62,In_71);
and U95 (N_95,In_40,In_258);
nand U96 (N_96,In_462,In_369);
nand U97 (N_97,In_339,In_318);
xnor U98 (N_98,In_181,In_439);
xor U99 (N_99,In_390,In_484);
or U100 (N_100,In_352,In_241);
and U101 (N_101,In_49,N_86);
xnor U102 (N_102,In_454,In_182);
xnor U103 (N_103,In_364,In_68);
and U104 (N_104,N_96,In_286);
and U105 (N_105,N_41,In_215);
or U106 (N_106,In_169,In_374);
or U107 (N_107,In_303,N_13);
xor U108 (N_108,In_197,N_34);
nor U109 (N_109,In_358,In_322);
xor U110 (N_110,In_250,N_82);
xnor U111 (N_111,In_135,N_11);
or U112 (N_112,In_317,In_30);
or U113 (N_113,N_65,N_62);
nor U114 (N_114,In_157,In_416);
or U115 (N_115,In_228,In_57);
xor U116 (N_116,In_370,In_456);
and U117 (N_117,In_180,N_51);
xnor U118 (N_118,In_223,In_429);
nand U119 (N_119,N_98,In_171);
or U120 (N_120,N_44,N_3);
and U121 (N_121,N_30,In_74);
and U122 (N_122,N_57,In_244);
xor U123 (N_123,N_63,N_89);
nor U124 (N_124,N_12,N_88);
and U125 (N_125,In_321,N_71);
nand U126 (N_126,N_74,N_72);
nor U127 (N_127,In_102,In_308);
nor U128 (N_128,In_451,In_391);
or U129 (N_129,N_59,In_42);
and U130 (N_130,In_468,In_234);
and U131 (N_131,In_356,In_243);
or U132 (N_132,In_283,In_29);
nor U133 (N_133,N_97,In_177);
nand U134 (N_134,N_33,N_7);
nor U135 (N_135,In_56,In_55);
xnor U136 (N_136,In_207,In_17);
and U137 (N_137,N_16,In_259);
nor U138 (N_138,In_373,N_67);
and U139 (N_139,In_33,In_278);
xor U140 (N_140,In_381,In_420);
nor U141 (N_141,In_334,In_458);
nor U142 (N_142,In_144,In_35);
or U143 (N_143,N_38,N_81);
xor U144 (N_144,In_142,In_148);
nand U145 (N_145,In_175,N_76);
or U146 (N_146,In_331,In_248);
or U147 (N_147,In_289,In_31);
or U148 (N_148,In_387,In_145);
and U149 (N_149,In_326,N_46);
and U150 (N_150,N_42,In_307);
and U151 (N_151,N_55,In_406);
nand U152 (N_152,In_254,In_236);
nand U153 (N_153,In_255,In_34);
nand U154 (N_154,In_32,In_133);
and U155 (N_155,In_473,N_36);
xor U156 (N_156,In_12,In_466);
or U157 (N_157,In_187,In_433);
and U158 (N_158,In_196,In_151);
or U159 (N_159,In_397,In_108);
xor U160 (N_160,In_103,In_459);
nand U161 (N_161,N_73,In_166);
and U162 (N_162,In_156,In_265);
or U163 (N_163,N_94,N_90);
and U164 (N_164,In_146,In_430);
and U165 (N_165,In_449,N_84);
and U166 (N_166,In_354,In_463);
nor U167 (N_167,In_252,In_16);
or U168 (N_168,N_39,In_25);
or U169 (N_169,In_353,In_440);
xor U170 (N_170,In_355,In_340);
nor U171 (N_171,In_262,In_73);
and U172 (N_172,N_8,In_235);
and U173 (N_173,In_44,In_306);
xor U174 (N_174,N_40,N_31);
nand U175 (N_175,In_209,In_121);
or U176 (N_176,In_1,In_92);
nor U177 (N_177,In_287,In_88);
xnor U178 (N_178,In_141,In_272);
or U179 (N_179,In_99,In_6);
and U180 (N_180,In_167,In_445);
xnor U181 (N_181,In_476,N_10);
nor U182 (N_182,In_310,N_32);
or U183 (N_183,In_153,In_371);
and U184 (N_184,In_109,N_20);
and U185 (N_185,In_239,N_95);
nor U186 (N_186,N_99,In_20);
nor U187 (N_187,N_70,In_112);
or U188 (N_188,N_37,In_441);
nor U189 (N_189,In_296,In_184);
and U190 (N_190,In_493,In_43);
nor U191 (N_191,N_21,In_46);
xor U192 (N_192,N_83,N_1);
nor U193 (N_193,In_471,In_418);
nand U194 (N_194,In_261,In_211);
or U195 (N_195,In_10,In_407);
nand U196 (N_196,In_137,In_260);
nand U197 (N_197,In_80,In_138);
nand U198 (N_198,N_2,In_53);
nor U199 (N_199,In_101,N_75);
and U200 (N_200,N_17,N_102);
nor U201 (N_201,N_157,N_132);
or U202 (N_202,In_193,N_181);
or U203 (N_203,In_115,In_195);
xor U204 (N_204,In_400,In_104);
and U205 (N_205,In_455,N_186);
xor U206 (N_206,In_41,In_412);
and U207 (N_207,N_196,N_4);
nor U208 (N_208,N_66,In_253);
or U209 (N_209,N_110,In_319);
nand U210 (N_210,N_78,In_408);
nor U211 (N_211,In_378,In_274);
nand U212 (N_212,In_489,In_123);
nand U213 (N_213,In_499,N_144);
nand U214 (N_214,N_154,N_187);
nand U215 (N_215,In_365,N_147);
and U216 (N_216,In_97,N_149);
nor U217 (N_217,N_61,N_195);
nor U218 (N_218,In_368,N_199);
xor U219 (N_219,In_366,In_482);
xnor U220 (N_220,In_288,N_191);
xnor U221 (N_221,In_238,In_132);
nand U222 (N_222,N_52,In_189);
and U223 (N_223,N_182,N_140);
nor U224 (N_224,N_174,In_363);
and U225 (N_225,N_160,In_388);
nand U226 (N_226,N_108,In_164);
nand U227 (N_227,In_280,In_295);
nor U228 (N_228,N_192,In_245);
nor U229 (N_229,N_197,N_134);
and U230 (N_230,In_389,N_115);
nand U231 (N_231,N_93,In_226);
or U232 (N_232,N_167,In_292);
xnor U233 (N_233,N_0,N_179);
and U234 (N_234,N_100,N_129);
nor U235 (N_235,N_54,In_134);
xor U236 (N_236,N_188,In_332);
or U237 (N_237,In_375,N_79);
and U238 (N_238,N_194,In_386);
and U239 (N_239,In_213,In_435);
and U240 (N_240,N_164,N_47);
and U241 (N_241,N_23,In_257);
and U242 (N_242,In_315,In_413);
nor U243 (N_243,In_72,In_320);
nand U244 (N_244,In_158,In_447);
and U245 (N_245,N_104,In_147);
nand U246 (N_246,N_178,In_263);
nor U247 (N_247,In_246,N_171);
and U248 (N_248,N_114,N_198);
or U249 (N_249,In_421,In_483);
xor U250 (N_250,N_126,N_5);
xnor U251 (N_251,In_110,In_485);
nor U252 (N_252,N_105,N_29);
nand U253 (N_253,In_81,In_2);
or U254 (N_254,In_345,N_14);
nor U255 (N_255,N_60,N_177);
or U256 (N_256,In_270,In_67);
nor U257 (N_257,N_18,In_329);
nor U258 (N_258,N_68,In_437);
xnor U259 (N_259,N_49,N_172);
or U260 (N_260,N_64,N_124);
xnor U261 (N_261,N_35,In_314);
nor U262 (N_262,N_92,In_266);
nor U263 (N_263,N_27,In_174);
xnor U264 (N_264,In_185,In_48);
nor U265 (N_265,N_103,N_183);
nand U266 (N_266,In_8,N_80);
nand U267 (N_267,N_113,In_38);
nand U268 (N_268,N_176,In_107);
nor U269 (N_269,N_123,N_142);
nand U270 (N_270,N_162,In_15);
nand U271 (N_271,In_277,N_153);
nor U272 (N_272,In_64,In_491);
nand U273 (N_273,In_376,N_155);
nor U274 (N_274,In_50,N_148);
nand U275 (N_275,In_58,In_279);
or U276 (N_276,In_176,N_184);
nor U277 (N_277,N_158,In_268);
nor U278 (N_278,N_85,N_136);
nand U279 (N_279,In_220,N_141);
nor U280 (N_280,N_137,N_125);
nor U281 (N_281,In_432,N_48);
or U282 (N_282,N_22,N_166);
and U283 (N_283,In_398,N_190);
xor U284 (N_284,N_91,N_117);
xnor U285 (N_285,N_116,In_409);
nor U286 (N_286,N_69,In_299);
and U287 (N_287,In_150,In_444);
nand U288 (N_288,N_28,N_109);
or U289 (N_289,In_324,N_107);
nand U290 (N_290,In_3,In_267);
and U291 (N_291,In_361,N_152);
nor U292 (N_292,In_113,In_392);
or U293 (N_293,N_161,N_159);
xor U294 (N_294,N_56,In_100);
or U295 (N_295,In_481,In_201);
and U296 (N_296,N_50,In_457);
xor U297 (N_297,In_498,N_151);
and U298 (N_298,N_19,In_423);
xnor U299 (N_299,In_69,N_156);
xor U300 (N_300,N_290,N_211);
or U301 (N_301,N_276,N_270);
and U302 (N_302,N_227,N_246);
xor U303 (N_303,In_460,N_228);
nor U304 (N_304,N_231,N_168);
or U305 (N_305,N_264,In_125);
nand U306 (N_306,In_395,In_82);
nand U307 (N_307,In_333,N_224);
nand U308 (N_308,N_220,N_234);
xnor U309 (N_309,N_232,In_336);
nor U310 (N_310,N_121,N_118);
nor U311 (N_311,N_201,N_283);
xor U312 (N_312,N_245,N_298);
nand U313 (N_313,N_222,N_278);
and U314 (N_314,In_465,N_260);
xnor U315 (N_315,N_271,N_281);
nor U316 (N_316,N_130,N_254);
nand U317 (N_317,N_219,In_7);
xnor U318 (N_318,N_131,N_252);
nand U319 (N_319,N_204,In_276);
or U320 (N_320,N_253,N_170);
or U321 (N_321,N_133,In_428);
nand U322 (N_322,N_128,N_119);
and U323 (N_323,N_262,N_120);
nand U324 (N_324,N_25,N_214);
or U325 (N_325,N_203,In_282);
nand U326 (N_326,In_330,N_239);
or U327 (N_327,In_309,N_274);
xor U328 (N_328,N_297,N_206);
nor U329 (N_329,In_208,N_217);
nor U330 (N_330,N_277,N_266);
and U331 (N_331,N_291,In_350);
xor U332 (N_332,In_477,In_52);
nand U333 (N_333,N_235,N_242);
nor U334 (N_334,In_26,N_233);
or U335 (N_335,N_175,N_288);
nand U336 (N_336,N_226,In_474);
or U337 (N_337,N_282,In_61);
and U338 (N_338,N_241,N_200);
xnor U339 (N_339,In_342,N_205);
or U340 (N_340,In_431,N_207);
and U341 (N_341,N_173,N_24);
xnor U342 (N_342,N_169,N_58);
and U343 (N_343,N_138,N_279);
nand U344 (N_344,In_214,N_45);
or U345 (N_345,N_261,N_257);
nand U346 (N_346,N_77,In_442);
and U347 (N_347,N_87,N_240);
xor U348 (N_348,N_244,N_202);
xnor U349 (N_349,In_122,N_285);
or U350 (N_350,In_86,N_43);
or U351 (N_351,N_284,In_249);
xor U352 (N_352,In_328,In_63);
or U353 (N_353,In_467,N_185);
and U354 (N_354,N_236,In_217);
nand U355 (N_355,In_372,In_301);
nand U356 (N_356,N_213,In_85);
nor U357 (N_357,N_106,In_232);
or U358 (N_358,N_15,N_286);
or U359 (N_359,N_295,N_269);
or U360 (N_360,N_243,N_299);
xnor U361 (N_361,N_216,In_188);
nor U362 (N_362,In_124,N_293);
nand U363 (N_363,In_285,N_250);
and U364 (N_364,N_145,N_122);
and U365 (N_365,In_84,N_189);
nor U366 (N_366,In_51,N_135);
nor U367 (N_367,N_165,N_209);
and U368 (N_368,N_53,N_238);
xor U369 (N_369,N_146,N_127);
or U370 (N_370,N_280,N_215);
nor U371 (N_371,In_206,N_193);
or U372 (N_372,N_229,In_346);
and U373 (N_373,N_111,N_139);
or U374 (N_374,N_237,N_112);
nand U375 (N_375,N_223,In_161);
xnor U376 (N_376,In_480,N_210);
and U377 (N_377,N_230,N_258);
xnor U378 (N_378,N_248,In_422);
xor U379 (N_379,In_359,In_136);
and U380 (N_380,N_26,N_256);
xnor U381 (N_381,In_300,In_170);
nor U382 (N_382,N_263,N_180);
nand U383 (N_383,N_292,N_273);
and U384 (N_384,N_6,N_294);
and U385 (N_385,In_204,N_268);
nor U386 (N_386,N_259,In_497);
and U387 (N_387,N_163,N_101);
xnor U388 (N_388,N_296,N_212);
nand U389 (N_389,In_139,In_379);
nor U390 (N_390,N_150,N_143);
nor U391 (N_391,N_221,In_19);
xnor U392 (N_392,N_225,N_251);
nor U393 (N_393,In_323,N_272);
nand U394 (N_394,N_9,N_208);
and U395 (N_395,N_255,N_287);
and U396 (N_396,N_289,N_249);
or U397 (N_397,In_294,N_267);
or U398 (N_398,N_275,N_265);
xor U399 (N_399,N_218,N_247);
nand U400 (N_400,N_331,N_383);
or U401 (N_401,N_392,N_346);
nand U402 (N_402,N_355,N_399);
and U403 (N_403,N_338,N_328);
nand U404 (N_404,N_345,N_381);
xor U405 (N_405,N_359,N_390);
and U406 (N_406,N_318,N_382);
or U407 (N_407,N_301,N_315);
nor U408 (N_408,N_327,N_317);
nor U409 (N_409,N_394,N_370);
nand U410 (N_410,N_324,N_393);
nor U411 (N_411,N_341,N_351);
or U412 (N_412,N_352,N_363);
and U413 (N_413,N_316,N_364);
xnor U414 (N_414,N_313,N_333);
nor U415 (N_415,N_362,N_342);
and U416 (N_416,N_358,N_320);
nand U417 (N_417,N_369,N_360);
xor U418 (N_418,N_374,N_300);
xor U419 (N_419,N_373,N_319);
or U420 (N_420,N_309,N_388);
and U421 (N_421,N_326,N_302);
xor U422 (N_422,N_308,N_347);
xnor U423 (N_423,N_391,N_305);
nand U424 (N_424,N_310,N_397);
nand U425 (N_425,N_376,N_385);
nor U426 (N_426,N_343,N_365);
or U427 (N_427,N_387,N_372);
or U428 (N_428,N_337,N_306);
or U429 (N_429,N_330,N_350);
and U430 (N_430,N_340,N_356);
nand U431 (N_431,N_377,N_334);
and U432 (N_432,N_384,N_339);
and U433 (N_433,N_395,N_398);
or U434 (N_434,N_322,N_314);
and U435 (N_435,N_379,N_312);
xnor U436 (N_436,N_329,N_323);
nand U437 (N_437,N_349,N_307);
or U438 (N_438,N_311,N_357);
nand U439 (N_439,N_361,N_321);
nand U440 (N_440,N_371,N_335);
nor U441 (N_441,N_366,N_353);
and U442 (N_442,N_367,N_336);
nand U443 (N_443,N_386,N_375);
or U444 (N_444,N_378,N_354);
and U445 (N_445,N_348,N_380);
nand U446 (N_446,N_368,N_325);
xor U447 (N_447,N_332,N_396);
nand U448 (N_448,N_304,N_389);
and U449 (N_449,N_303,N_344);
nor U450 (N_450,N_328,N_388);
nand U451 (N_451,N_307,N_317);
or U452 (N_452,N_315,N_383);
nand U453 (N_453,N_331,N_387);
and U454 (N_454,N_317,N_325);
xor U455 (N_455,N_396,N_353);
nor U456 (N_456,N_303,N_366);
nor U457 (N_457,N_300,N_358);
nand U458 (N_458,N_352,N_316);
and U459 (N_459,N_315,N_311);
xor U460 (N_460,N_375,N_301);
nor U461 (N_461,N_374,N_317);
nor U462 (N_462,N_326,N_327);
xor U463 (N_463,N_342,N_303);
and U464 (N_464,N_324,N_360);
nand U465 (N_465,N_362,N_373);
or U466 (N_466,N_324,N_361);
or U467 (N_467,N_368,N_340);
nor U468 (N_468,N_390,N_312);
xor U469 (N_469,N_361,N_330);
nor U470 (N_470,N_342,N_361);
nor U471 (N_471,N_322,N_374);
nor U472 (N_472,N_364,N_351);
xnor U473 (N_473,N_384,N_300);
nand U474 (N_474,N_344,N_394);
or U475 (N_475,N_350,N_313);
nand U476 (N_476,N_320,N_354);
and U477 (N_477,N_368,N_351);
and U478 (N_478,N_379,N_307);
or U479 (N_479,N_345,N_377);
or U480 (N_480,N_323,N_372);
nor U481 (N_481,N_396,N_395);
xor U482 (N_482,N_347,N_354);
xnor U483 (N_483,N_335,N_357);
nor U484 (N_484,N_349,N_386);
xor U485 (N_485,N_350,N_329);
xnor U486 (N_486,N_398,N_359);
xor U487 (N_487,N_396,N_376);
xor U488 (N_488,N_346,N_339);
xor U489 (N_489,N_387,N_347);
and U490 (N_490,N_316,N_394);
xor U491 (N_491,N_308,N_358);
nor U492 (N_492,N_306,N_311);
or U493 (N_493,N_358,N_382);
nor U494 (N_494,N_364,N_319);
or U495 (N_495,N_370,N_343);
nand U496 (N_496,N_376,N_386);
nand U497 (N_497,N_343,N_395);
nand U498 (N_498,N_353,N_367);
and U499 (N_499,N_352,N_382);
and U500 (N_500,N_444,N_475);
nor U501 (N_501,N_409,N_465);
nor U502 (N_502,N_470,N_499);
nand U503 (N_503,N_414,N_464);
xnor U504 (N_504,N_481,N_495);
and U505 (N_505,N_426,N_491);
and U506 (N_506,N_431,N_445);
nand U507 (N_507,N_419,N_441);
or U508 (N_508,N_484,N_483);
and U509 (N_509,N_497,N_466);
xnor U510 (N_510,N_478,N_402);
xnor U511 (N_511,N_450,N_489);
or U512 (N_512,N_451,N_418);
or U513 (N_513,N_458,N_428);
and U514 (N_514,N_435,N_420);
nand U515 (N_515,N_437,N_463);
and U516 (N_516,N_448,N_460);
xnor U517 (N_517,N_468,N_410);
nor U518 (N_518,N_439,N_477);
and U519 (N_519,N_492,N_446);
xor U520 (N_520,N_442,N_443);
or U521 (N_521,N_433,N_494);
nor U522 (N_522,N_440,N_421);
and U523 (N_523,N_413,N_403);
and U524 (N_524,N_488,N_411);
and U525 (N_525,N_429,N_438);
nor U526 (N_526,N_476,N_436);
and U527 (N_527,N_498,N_425);
or U528 (N_528,N_469,N_467);
nor U529 (N_529,N_493,N_496);
xnor U530 (N_530,N_473,N_406);
or U531 (N_531,N_407,N_482);
nand U532 (N_532,N_412,N_423);
and U533 (N_533,N_462,N_480);
or U534 (N_534,N_454,N_486);
or U535 (N_535,N_422,N_408);
and U536 (N_536,N_455,N_490);
or U537 (N_537,N_456,N_417);
nor U538 (N_538,N_452,N_453);
nand U539 (N_539,N_449,N_400);
nor U540 (N_540,N_401,N_474);
or U541 (N_541,N_424,N_430);
or U542 (N_542,N_432,N_472);
or U543 (N_543,N_415,N_485);
nand U544 (N_544,N_457,N_416);
nand U545 (N_545,N_459,N_461);
xnor U546 (N_546,N_404,N_405);
and U547 (N_547,N_479,N_471);
and U548 (N_548,N_427,N_487);
xnor U549 (N_549,N_434,N_447);
and U550 (N_550,N_406,N_400);
xor U551 (N_551,N_447,N_406);
nor U552 (N_552,N_447,N_438);
nor U553 (N_553,N_423,N_413);
nor U554 (N_554,N_472,N_448);
xnor U555 (N_555,N_497,N_459);
nor U556 (N_556,N_475,N_471);
nand U557 (N_557,N_447,N_491);
nand U558 (N_558,N_489,N_491);
xor U559 (N_559,N_420,N_428);
and U560 (N_560,N_432,N_404);
or U561 (N_561,N_410,N_401);
xnor U562 (N_562,N_475,N_485);
nor U563 (N_563,N_444,N_422);
nand U564 (N_564,N_455,N_431);
and U565 (N_565,N_459,N_430);
and U566 (N_566,N_433,N_474);
and U567 (N_567,N_484,N_401);
or U568 (N_568,N_408,N_410);
nor U569 (N_569,N_468,N_466);
xnor U570 (N_570,N_484,N_430);
or U571 (N_571,N_415,N_491);
or U572 (N_572,N_415,N_458);
nand U573 (N_573,N_440,N_493);
xnor U574 (N_574,N_425,N_485);
xor U575 (N_575,N_450,N_402);
and U576 (N_576,N_477,N_420);
nor U577 (N_577,N_422,N_470);
xnor U578 (N_578,N_419,N_433);
nand U579 (N_579,N_477,N_402);
xor U580 (N_580,N_420,N_451);
xor U581 (N_581,N_464,N_413);
nand U582 (N_582,N_493,N_420);
or U583 (N_583,N_414,N_426);
and U584 (N_584,N_454,N_463);
nor U585 (N_585,N_439,N_444);
nor U586 (N_586,N_454,N_421);
nor U587 (N_587,N_421,N_431);
or U588 (N_588,N_456,N_465);
xnor U589 (N_589,N_431,N_413);
nor U590 (N_590,N_483,N_417);
or U591 (N_591,N_429,N_406);
xor U592 (N_592,N_470,N_485);
or U593 (N_593,N_474,N_415);
nor U594 (N_594,N_421,N_484);
or U595 (N_595,N_487,N_475);
nor U596 (N_596,N_478,N_457);
or U597 (N_597,N_439,N_413);
and U598 (N_598,N_411,N_457);
and U599 (N_599,N_484,N_443);
and U600 (N_600,N_552,N_598);
and U601 (N_601,N_550,N_597);
or U602 (N_602,N_518,N_587);
nand U603 (N_603,N_585,N_522);
and U604 (N_604,N_508,N_529);
and U605 (N_605,N_599,N_576);
nand U606 (N_606,N_525,N_504);
or U607 (N_607,N_543,N_548);
nor U608 (N_608,N_530,N_590);
or U609 (N_609,N_563,N_596);
nand U610 (N_610,N_592,N_568);
nand U611 (N_611,N_521,N_527);
and U612 (N_612,N_577,N_559);
and U613 (N_613,N_594,N_534);
or U614 (N_614,N_578,N_512);
or U615 (N_615,N_581,N_560);
nand U616 (N_616,N_555,N_588);
and U617 (N_617,N_566,N_516);
xnor U618 (N_618,N_574,N_547);
nand U619 (N_619,N_557,N_584);
and U620 (N_620,N_505,N_583);
or U621 (N_621,N_517,N_519);
or U622 (N_622,N_523,N_501);
nand U623 (N_623,N_520,N_573);
or U624 (N_624,N_593,N_500);
nor U625 (N_625,N_513,N_591);
and U626 (N_626,N_515,N_514);
nor U627 (N_627,N_589,N_532);
or U628 (N_628,N_542,N_503);
and U629 (N_629,N_561,N_540);
xor U630 (N_630,N_536,N_579);
and U631 (N_631,N_537,N_507);
xor U632 (N_632,N_549,N_580);
xnor U633 (N_633,N_531,N_528);
nand U634 (N_634,N_526,N_553);
nand U635 (N_635,N_586,N_575);
and U636 (N_636,N_541,N_506);
nand U637 (N_637,N_546,N_545);
and U638 (N_638,N_565,N_511);
nand U639 (N_639,N_571,N_533);
xnor U640 (N_640,N_510,N_509);
nand U641 (N_641,N_595,N_539);
nor U642 (N_642,N_572,N_564);
or U643 (N_643,N_502,N_538);
and U644 (N_644,N_524,N_551);
xnor U645 (N_645,N_582,N_535);
xnor U646 (N_646,N_558,N_569);
xor U647 (N_647,N_567,N_544);
nor U648 (N_648,N_556,N_562);
or U649 (N_649,N_554,N_570);
xnor U650 (N_650,N_514,N_501);
or U651 (N_651,N_505,N_591);
or U652 (N_652,N_527,N_516);
and U653 (N_653,N_541,N_535);
or U654 (N_654,N_591,N_560);
nand U655 (N_655,N_567,N_553);
xor U656 (N_656,N_516,N_590);
xor U657 (N_657,N_593,N_547);
nand U658 (N_658,N_535,N_593);
and U659 (N_659,N_515,N_556);
xor U660 (N_660,N_549,N_525);
or U661 (N_661,N_526,N_522);
nand U662 (N_662,N_599,N_553);
and U663 (N_663,N_526,N_550);
nand U664 (N_664,N_518,N_582);
xor U665 (N_665,N_506,N_569);
nor U666 (N_666,N_529,N_528);
and U667 (N_667,N_520,N_591);
and U668 (N_668,N_552,N_584);
and U669 (N_669,N_569,N_518);
xnor U670 (N_670,N_528,N_579);
and U671 (N_671,N_531,N_522);
nand U672 (N_672,N_547,N_533);
nand U673 (N_673,N_583,N_596);
or U674 (N_674,N_507,N_533);
nor U675 (N_675,N_539,N_514);
or U676 (N_676,N_543,N_500);
and U677 (N_677,N_517,N_576);
xnor U678 (N_678,N_502,N_507);
xor U679 (N_679,N_545,N_527);
xor U680 (N_680,N_536,N_506);
and U681 (N_681,N_504,N_518);
and U682 (N_682,N_538,N_587);
nor U683 (N_683,N_581,N_512);
xor U684 (N_684,N_581,N_515);
nor U685 (N_685,N_507,N_578);
nor U686 (N_686,N_527,N_526);
nor U687 (N_687,N_501,N_513);
nand U688 (N_688,N_594,N_537);
xnor U689 (N_689,N_536,N_523);
or U690 (N_690,N_585,N_513);
and U691 (N_691,N_566,N_535);
or U692 (N_692,N_533,N_589);
or U693 (N_693,N_552,N_578);
nor U694 (N_694,N_524,N_538);
nor U695 (N_695,N_526,N_518);
nor U696 (N_696,N_533,N_569);
nand U697 (N_697,N_566,N_521);
xor U698 (N_698,N_542,N_500);
and U699 (N_699,N_541,N_555);
or U700 (N_700,N_695,N_652);
or U701 (N_701,N_624,N_689);
and U702 (N_702,N_602,N_667);
and U703 (N_703,N_638,N_601);
nor U704 (N_704,N_678,N_635);
nor U705 (N_705,N_661,N_639);
nor U706 (N_706,N_653,N_604);
xnor U707 (N_707,N_693,N_671);
nand U708 (N_708,N_609,N_644);
nand U709 (N_709,N_658,N_686);
nor U710 (N_710,N_647,N_657);
nor U711 (N_711,N_632,N_676);
nand U712 (N_712,N_649,N_614);
xor U713 (N_713,N_674,N_626);
and U714 (N_714,N_672,N_688);
and U715 (N_715,N_692,N_616);
or U716 (N_716,N_675,N_603);
or U717 (N_717,N_643,N_600);
nand U718 (N_718,N_659,N_613);
nand U719 (N_719,N_669,N_683);
xnor U720 (N_720,N_610,N_621);
nor U721 (N_721,N_642,N_654);
nor U722 (N_722,N_650,N_637);
or U723 (N_723,N_681,N_611);
and U724 (N_724,N_631,N_690);
xnor U725 (N_725,N_617,N_655);
nor U726 (N_726,N_646,N_677);
or U727 (N_727,N_687,N_696);
or U728 (N_728,N_622,N_664);
or U729 (N_729,N_606,N_685);
nor U730 (N_730,N_679,N_615);
xor U731 (N_731,N_684,N_682);
xor U732 (N_732,N_627,N_618);
and U733 (N_733,N_668,N_697);
nand U734 (N_734,N_680,N_633);
nor U735 (N_735,N_619,N_629);
nor U736 (N_736,N_612,N_648);
nor U737 (N_737,N_651,N_634);
xnor U738 (N_738,N_641,N_694);
nand U739 (N_739,N_623,N_636);
xnor U740 (N_740,N_673,N_620);
or U741 (N_741,N_663,N_699);
nand U742 (N_742,N_662,N_665);
or U743 (N_743,N_656,N_608);
xnor U744 (N_744,N_698,N_607);
and U745 (N_745,N_660,N_691);
xnor U746 (N_746,N_628,N_630);
nand U747 (N_747,N_645,N_666);
xnor U748 (N_748,N_640,N_625);
xnor U749 (N_749,N_670,N_605);
and U750 (N_750,N_654,N_645);
xor U751 (N_751,N_609,N_682);
xnor U752 (N_752,N_694,N_639);
or U753 (N_753,N_624,N_684);
xor U754 (N_754,N_646,N_629);
or U755 (N_755,N_621,N_617);
or U756 (N_756,N_629,N_637);
and U757 (N_757,N_697,N_661);
and U758 (N_758,N_661,N_641);
nor U759 (N_759,N_622,N_679);
nand U760 (N_760,N_662,N_673);
xor U761 (N_761,N_609,N_634);
or U762 (N_762,N_625,N_658);
nor U763 (N_763,N_653,N_666);
nand U764 (N_764,N_612,N_610);
and U765 (N_765,N_675,N_669);
and U766 (N_766,N_601,N_633);
and U767 (N_767,N_643,N_687);
nor U768 (N_768,N_683,N_605);
xor U769 (N_769,N_641,N_674);
nand U770 (N_770,N_604,N_640);
xnor U771 (N_771,N_677,N_609);
or U772 (N_772,N_688,N_608);
or U773 (N_773,N_665,N_679);
or U774 (N_774,N_653,N_677);
and U775 (N_775,N_662,N_645);
xnor U776 (N_776,N_620,N_626);
nand U777 (N_777,N_646,N_609);
nand U778 (N_778,N_682,N_656);
nor U779 (N_779,N_628,N_671);
nand U780 (N_780,N_681,N_639);
nand U781 (N_781,N_673,N_643);
nand U782 (N_782,N_600,N_686);
or U783 (N_783,N_620,N_608);
nor U784 (N_784,N_643,N_661);
xnor U785 (N_785,N_670,N_691);
nand U786 (N_786,N_611,N_651);
and U787 (N_787,N_685,N_609);
and U788 (N_788,N_692,N_667);
nor U789 (N_789,N_697,N_623);
and U790 (N_790,N_665,N_696);
and U791 (N_791,N_675,N_607);
nand U792 (N_792,N_698,N_650);
and U793 (N_793,N_621,N_616);
nand U794 (N_794,N_650,N_636);
and U795 (N_795,N_621,N_696);
nand U796 (N_796,N_613,N_631);
or U797 (N_797,N_671,N_616);
xnor U798 (N_798,N_627,N_695);
or U799 (N_799,N_653,N_698);
or U800 (N_800,N_785,N_763);
and U801 (N_801,N_744,N_720);
nor U802 (N_802,N_746,N_731);
xnor U803 (N_803,N_703,N_737);
xor U804 (N_804,N_711,N_791);
nor U805 (N_805,N_733,N_762);
nand U806 (N_806,N_768,N_755);
nor U807 (N_807,N_714,N_753);
or U808 (N_808,N_759,N_715);
or U809 (N_809,N_776,N_705);
nor U810 (N_810,N_794,N_738);
xor U811 (N_811,N_792,N_741);
or U812 (N_812,N_745,N_771);
xnor U813 (N_813,N_749,N_770);
nor U814 (N_814,N_765,N_751);
nor U815 (N_815,N_787,N_707);
and U816 (N_816,N_708,N_793);
or U817 (N_817,N_717,N_784);
nor U818 (N_818,N_724,N_712);
xor U819 (N_819,N_783,N_760);
xor U820 (N_820,N_713,N_701);
xor U821 (N_821,N_774,N_723);
nor U822 (N_822,N_706,N_775);
xnor U823 (N_823,N_778,N_748);
nand U824 (N_824,N_782,N_797);
and U825 (N_825,N_798,N_750);
or U826 (N_826,N_747,N_735);
or U827 (N_827,N_700,N_734);
nand U828 (N_828,N_726,N_722);
nor U829 (N_829,N_739,N_752);
or U830 (N_830,N_718,N_728);
nor U831 (N_831,N_725,N_757);
or U832 (N_832,N_799,N_742);
nand U833 (N_833,N_796,N_780);
xor U834 (N_834,N_777,N_743);
or U835 (N_835,N_761,N_789);
nand U836 (N_836,N_766,N_781);
xnor U837 (N_837,N_754,N_758);
nand U838 (N_838,N_736,N_756);
or U839 (N_839,N_767,N_704);
nand U840 (N_840,N_719,N_740);
xnor U841 (N_841,N_773,N_772);
nor U842 (N_842,N_702,N_795);
xor U843 (N_843,N_730,N_779);
or U844 (N_844,N_790,N_710);
and U845 (N_845,N_721,N_709);
nand U846 (N_846,N_716,N_729);
or U847 (N_847,N_732,N_764);
nand U848 (N_848,N_769,N_727);
xnor U849 (N_849,N_788,N_786);
nor U850 (N_850,N_718,N_724);
nor U851 (N_851,N_725,N_722);
xnor U852 (N_852,N_794,N_716);
nand U853 (N_853,N_767,N_733);
and U854 (N_854,N_764,N_738);
and U855 (N_855,N_777,N_739);
xnor U856 (N_856,N_728,N_751);
nor U857 (N_857,N_759,N_702);
xor U858 (N_858,N_711,N_734);
nor U859 (N_859,N_762,N_753);
and U860 (N_860,N_779,N_788);
xor U861 (N_861,N_723,N_722);
nor U862 (N_862,N_719,N_795);
nor U863 (N_863,N_799,N_775);
xnor U864 (N_864,N_742,N_730);
nand U865 (N_865,N_783,N_796);
or U866 (N_866,N_796,N_739);
xor U867 (N_867,N_782,N_746);
nand U868 (N_868,N_744,N_762);
xor U869 (N_869,N_798,N_756);
xor U870 (N_870,N_741,N_763);
xnor U871 (N_871,N_795,N_708);
nor U872 (N_872,N_730,N_768);
nor U873 (N_873,N_722,N_715);
and U874 (N_874,N_739,N_756);
nor U875 (N_875,N_749,N_731);
xor U876 (N_876,N_752,N_775);
nand U877 (N_877,N_791,N_795);
nor U878 (N_878,N_736,N_781);
nand U879 (N_879,N_729,N_786);
nand U880 (N_880,N_710,N_796);
nand U881 (N_881,N_776,N_758);
xor U882 (N_882,N_700,N_761);
nor U883 (N_883,N_723,N_729);
and U884 (N_884,N_742,N_772);
nor U885 (N_885,N_705,N_790);
or U886 (N_886,N_737,N_710);
or U887 (N_887,N_743,N_750);
nor U888 (N_888,N_728,N_715);
nor U889 (N_889,N_757,N_780);
or U890 (N_890,N_725,N_783);
or U891 (N_891,N_733,N_701);
and U892 (N_892,N_716,N_777);
nand U893 (N_893,N_710,N_789);
and U894 (N_894,N_702,N_717);
nand U895 (N_895,N_791,N_744);
or U896 (N_896,N_765,N_789);
nand U897 (N_897,N_794,N_745);
nand U898 (N_898,N_725,N_714);
nand U899 (N_899,N_726,N_774);
nor U900 (N_900,N_856,N_809);
or U901 (N_901,N_816,N_847);
and U902 (N_902,N_884,N_890);
and U903 (N_903,N_898,N_849);
nor U904 (N_904,N_808,N_881);
nor U905 (N_905,N_801,N_807);
xnor U906 (N_906,N_851,N_872);
xnor U907 (N_907,N_818,N_826);
xnor U908 (N_908,N_854,N_817);
and U909 (N_909,N_824,N_877);
nand U910 (N_910,N_861,N_855);
nor U911 (N_911,N_837,N_870);
and U912 (N_912,N_839,N_843);
nor U913 (N_913,N_848,N_806);
nor U914 (N_914,N_862,N_814);
and U915 (N_915,N_878,N_800);
or U916 (N_916,N_876,N_857);
or U917 (N_917,N_812,N_873);
xnor U918 (N_918,N_838,N_874);
xnor U919 (N_919,N_805,N_882);
nand U920 (N_920,N_832,N_819);
xor U921 (N_921,N_892,N_835);
nor U922 (N_922,N_827,N_825);
nand U923 (N_923,N_820,N_811);
or U924 (N_924,N_871,N_864);
nand U925 (N_925,N_893,N_803);
or U926 (N_926,N_859,N_845);
nor U927 (N_927,N_858,N_863);
nor U928 (N_928,N_888,N_886);
nor U929 (N_929,N_831,N_852);
nand U930 (N_930,N_828,N_869);
xnor U931 (N_931,N_887,N_815);
xnor U932 (N_932,N_810,N_899);
nor U933 (N_933,N_875,N_885);
or U934 (N_934,N_842,N_834);
or U935 (N_935,N_866,N_844);
xor U936 (N_936,N_830,N_891);
or U937 (N_937,N_889,N_813);
xor U938 (N_938,N_853,N_865);
or U939 (N_939,N_846,N_821);
nand U940 (N_940,N_836,N_804);
xor U941 (N_941,N_895,N_879);
or U942 (N_942,N_850,N_896);
nor U943 (N_943,N_822,N_860);
or U944 (N_944,N_841,N_894);
or U945 (N_945,N_880,N_829);
nand U946 (N_946,N_897,N_867);
xor U947 (N_947,N_883,N_840);
nor U948 (N_948,N_823,N_802);
nor U949 (N_949,N_868,N_833);
and U950 (N_950,N_806,N_864);
nand U951 (N_951,N_866,N_855);
nand U952 (N_952,N_811,N_877);
xnor U953 (N_953,N_856,N_843);
xnor U954 (N_954,N_893,N_820);
or U955 (N_955,N_870,N_882);
xor U956 (N_956,N_817,N_835);
and U957 (N_957,N_882,N_848);
and U958 (N_958,N_852,N_850);
nand U959 (N_959,N_825,N_833);
nand U960 (N_960,N_882,N_844);
xnor U961 (N_961,N_857,N_816);
and U962 (N_962,N_849,N_868);
xnor U963 (N_963,N_839,N_826);
or U964 (N_964,N_872,N_876);
or U965 (N_965,N_861,N_890);
nor U966 (N_966,N_807,N_859);
and U967 (N_967,N_842,N_809);
and U968 (N_968,N_871,N_805);
nor U969 (N_969,N_895,N_830);
xor U970 (N_970,N_833,N_814);
nand U971 (N_971,N_873,N_854);
or U972 (N_972,N_815,N_838);
nand U973 (N_973,N_834,N_861);
xor U974 (N_974,N_844,N_809);
xor U975 (N_975,N_875,N_810);
and U976 (N_976,N_830,N_820);
nor U977 (N_977,N_843,N_858);
nor U978 (N_978,N_849,N_825);
xor U979 (N_979,N_846,N_892);
nor U980 (N_980,N_864,N_856);
and U981 (N_981,N_851,N_864);
nand U982 (N_982,N_880,N_821);
nand U983 (N_983,N_833,N_818);
nand U984 (N_984,N_876,N_800);
and U985 (N_985,N_893,N_810);
xor U986 (N_986,N_832,N_833);
or U987 (N_987,N_830,N_826);
nor U988 (N_988,N_835,N_877);
xnor U989 (N_989,N_857,N_831);
and U990 (N_990,N_846,N_886);
nand U991 (N_991,N_897,N_840);
or U992 (N_992,N_858,N_880);
xor U993 (N_993,N_833,N_895);
xnor U994 (N_994,N_808,N_883);
nand U995 (N_995,N_817,N_862);
xor U996 (N_996,N_861,N_841);
xor U997 (N_997,N_821,N_865);
nor U998 (N_998,N_853,N_877);
xnor U999 (N_999,N_822,N_883);
nor U1000 (N_1000,N_942,N_949);
nand U1001 (N_1001,N_947,N_944);
xnor U1002 (N_1002,N_982,N_918);
nor U1003 (N_1003,N_912,N_986);
xor U1004 (N_1004,N_921,N_935);
nand U1005 (N_1005,N_934,N_915);
or U1006 (N_1006,N_997,N_961);
xnor U1007 (N_1007,N_966,N_930);
nand U1008 (N_1008,N_979,N_992);
or U1009 (N_1009,N_953,N_938);
and U1010 (N_1010,N_985,N_907);
nand U1011 (N_1011,N_922,N_945);
nand U1012 (N_1012,N_959,N_906);
nor U1013 (N_1013,N_983,N_990);
and U1014 (N_1014,N_940,N_927);
nand U1015 (N_1015,N_937,N_969);
or U1016 (N_1016,N_984,N_914);
nand U1017 (N_1017,N_933,N_963);
or U1018 (N_1018,N_943,N_941);
nand U1019 (N_1019,N_996,N_994);
and U1020 (N_1020,N_957,N_999);
xnor U1021 (N_1021,N_950,N_951);
xnor U1022 (N_1022,N_916,N_978);
and U1023 (N_1023,N_967,N_926);
nor U1024 (N_1024,N_901,N_974);
nand U1025 (N_1025,N_975,N_929);
or U1026 (N_1026,N_923,N_952);
and U1027 (N_1027,N_968,N_920);
or U1028 (N_1028,N_905,N_970);
and U1029 (N_1029,N_928,N_991);
xnor U1030 (N_1030,N_932,N_977);
xor U1031 (N_1031,N_989,N_993);
and U1032 (N_1032,N_946,N_954);
xor U1033 (N_1033,N_980,N_972);
nand U1034 (N_1034,N_962,N_903);
and U1035 (N_1035,N_900,N_925);
and U1036 (N_1036,N_987,N_960);
or U1037 (N_1037,N_936,N_917);
nand U1038 (N_1038,N_904,N_998);
nand U1039 (N_1039,N_908,N_948);
nand U1040 (N_1040,N_973,N_965);
nand U1041 (N_1041,N_971,N_988);
and U1042 (N_1042,N_976,N_955);
and U1043 (N_1043,N_910,N_958);
and U1044 (N_1044,N_964,N_919);
nand U1045 (N_1045,N_913,N_931);
xor U1046 (N_1046,N_911,N_981);
and U1047 (N_1047,N_902,N_995);
nand U1048 (N_1048,N_924,N_956);
or U1049 (N_1049,N_939,N_909);
or U1050 (N_1050,N_972,N_958);
xnor U1051 (N_1051,N_939,N_991);
or U1052 (N_1052,N_950,N_946);
and U1053 (N_1053,N_972,N_915);
nor U1054 (N_1054,N_940,N_956);
or U1055 (N_1055,N_941,N_918);
nor U1056 (N_1056,N_944,N_909);
xnor U1057 (N_1057,N_935,N_942);
xor U1058 (N_1058,N_919,N_931);
or U1059 (N_1059,N_920,N_948);
nor U1060 (N_1060,N_992,N_912);
and U1061 (N_1061,N_969,N_974);
nand U1062 (N_1062,N_917,N_983);
xnor U1063 (N_1063,N_978,N_971);
xor U1064 (N_1064,N_967,N_902);
xnor U1065 (N_1065,N_983,N_967);
xor U1066 (N_1066,N_942,N_909);
and U1067 (N_1067,N_942,N_981);
xor U1068 (N_1068,N_922,N_996);
or U1069 (N_1069,N_917,N_951);
or U1070 (N_1070,N_938,N_945);
nand U1071 (N_1071,N_929,N_946);
and U1072 (N_1072,N_913,N_929);
and U1073 (N_1073,N_926,N_925);
nand U1074 (N_1074,N_907,N_902);
and U1075 (N_1075,N_932,N_962);
or U1076 (N_1076,N_907,N_960);
xnor U1077 (N_1077,N_929,N_901);
nand U1078 (N_1078,N_938,N_985);
or U1079 (N_1079,N_951,N_984);
nor U1080 (N_1080,N_998,N_917);
or U1081 (N_1081,N_931,N_906);
nor U1082 (N_1082,N_900,N_993);
and U1083 (N_1083,N_976,N_990);
nand U1084 (N_1084,N_920,N_938);
and U1085 (N_1085,N_969,N_907);
or U1086 (N_1086,N_928,N_945);
nor U1087 (N_1087,N_928,N_916);
xnor U1088 (N_1088,N_930,N_955);
nand U1089 (N_1089,N_924,N_901);
or U1090 (N_1090,N_985,N_978);
nand U1091 (N_1091,N_973,N_956);
nand U1092 (N_1092,N_953,N_922);
or U1093 (N_1093,N_933,N_958);
xnor U1094 (N_1094,N_917,N_934);
and U1095 (N_1095,N_958,N_948);
nor U1096 (N_1096,N_938,N_952);
nand U1097 (N_1097,N_975,N_915);
nand U1098 (N_1098,N_926,N_984);
xor U1099 (N_1099,N_999,N_948);
and U1100 (N_1100,N_1036,N_1063);
and U1101 (N_1101,N_1024,N_1086);
nor U1102 (N_1102,N_1014,N_1060);
and U1103 (N_1103,N_1002,N_1032);
or U1104 (N_1104,N_1096,N_1039);
xor U1105 (N_1105,N_1083,N_1098);
and U1106 (N_1106,N_1010,N_1057);
nand U1107 (N_1107,N_1090,N_1028);
and U1108 (N_1108,N_1008,N_1029);
or U1109 (N_1109,N_1064,N_1033);
nand U1110 (N_1110,N_1013,N_1005);
or U1111 (N_1111,N_1052,N_1011);
nand U1112 (N_1112,N_1000,N_1088);
and U1113 (N_1113,N_1045,N_1049);
and U1114 (N_1114,N_1006,N_1001);
nor U1115 (N_1115,N_1056,N_1012);
xnor U1116 (N_1116,N_1051,N_1079);
nor U1117 (N_1117,N_1007,N_1071);
xor U1118 (N_1118,N_1054,N_1048);
nor U1119 (N_1119,N_1059,N_1018);
and U1120 (N_1120,N_1035,N_1055);
and U1121 (N_1121,N_1040,N_1093);
nand U1122 (N_1122,N_1047,N_1075);
xnor U1123 (N_1123,N_1020,N_1061);
nor U1124 (N_1124,N_1030,N_1095);
and U1125 (N_1125,N_1097,N_1034);
or U1126 (N_1126,N_1026,N_1069);
nand U1127 (N_1127,N_1091,N_1043);
or U1128 (N_1128,N_1016,N_1017);
and U1129 (N_1129,N_1094,N_1073);
or U1130 (N_1130,N_1038,N_1070);
nand U1131 (N_1131,N_1021,N_1078);
xnor U1132 (N_1132,N_1058,N_1025);
or U1133 (N_1133,N_1041,N_1009);
nor U1134 (N_1134,N_1015,N_1050);
nand U1135 (N_1135,N_1031,N_1099);
and U1136 (N_1136,N_1082,N_1072);
xnor U1137 (N_1137,N_1053,N_1074);
nor U1138 (N_1138,N_1027,N_1089);
nor U1139 (N_1139,N_1081,N_1003);
or U1140 (N_1140,N_1067,N_1080);
nor U1141 (N_1141,N_1077,N_1062);
xnor U1142 (N_1142,N_1019,N_1065);
nand U1143 (N_1143,N_1022,N_1087);
nor U1144 (N_1144,N_1076,N_1004);
xnor U1145 (N_1145,N_1042,N_1092);
or U1146 (N_1146,N_1044,N_1084);
and U1147 (N_1147,N_1085,N_1068);
and U1148 (N_1148,N_1023,N_1037);
xor U1149 (N_1149,N_1046,N_1066);
or U1150 (N_1150,N_1087,N_1053);
xnor U1151 (N_1151,N_1075,N_1025);
xor U1152 (N_1152,N_1094,N_1058);
xnor U1153 (N_1153,N_1097,N_1012);
xnor U1154 (N_1154,N_1059,N_1077);
nand U1155 (N_1155,N_1011,N_1038);
nor U1156 (N_1156,N_1026,N_1052);
xor U1157 (N_1157,N_1053,N_1050);
nor U1158 (N_1158,N_1075,N_1011);
nand U1159 (N_1159,N_1035,N_1044);
nand U1160 (N_1160,N_1099,N_1045);
and U1161 (N_1161,N_1009,N_1031);
xor U1162 (N_1162,N_1035,N_1019);
or U1163 (N_1163,N_1093,N_1087);
xor U1164 (N_1164,N_1041,N_1001);
xnor U1165 (N_1165,N_1043,N_1066);
xor U1166 (N_1166,N_1092,N_1026);
or U1167 (N_1167,N_1026,N_1047);
or U1168 (N_1168,N_1057,N_1065);
nor U1169 (N_1169,N_1025,N_1092);
or U1170 (N_1170,N_1011,N_1001);
and U1171 (N_1171,N_1043,N_1030);
and U1172 (N_1172,N_1054,N_1019);
nor U1173 (N_1173,N_1081,N_1063);
and U1174 (N_1174,N_1028,N_1052);
xor U1175 (N_1175,N_1017,N_1056);
nor U1176 (N_1176,N_1024,N_1015);
xnor U1177 (N_1177,N_1009,N_1050);
or U1178 (N_1178,N_1097,N_1047);
xnor U1179 (N_1179,N_1081,N_1057);
nand U1180 (N_1180,N_1008,N_1052);
xor U1181 (N_1181,N_1093,N_1069);
nand U1182 (N_1182,N_1095,N_1062);
xnor U1183 (N_1183,N_1060,N_1000);
nand U1184 (N_1184,N_1029,N_1091);
or U1185 (N_1185,N_1023,N_1029);
nor U1186 (N_1186,N_1084,N_1081);
nor U1187 (N_1187,N_1025,N_1091);
nor U1188 (N_1188,N_1085,N_1097);
nor U1189 (N_1189,N_1089,N_1079);
xor U1190 (N_1190,N_1018,N_1056);
or U1191 (N_1191,N_1088,N_1035);
or U1192 (N_1192,N_1057,N_1029);
nand U1193 (N_1193,N_1041,N_1099);
or U1194 (N_1194,N_1044,N_1079);
and U1195 (N_1195,N_1045,N_1066);
nand U1196 (N_1196,N_1080,N_1004);
xnor U1197 (N_1197,N_1087,N_1080);
nand U1198 (N_1198,N_1069,N_1062);
nand U1199 (N_1199,N_1016,N_1060);
nor U1200 (N_1200,N_1157,N_1116);
nand U1201 (N_1201,N_1102,N_1131);
nand U1202 (N_1202,N_1171,N_1142);
nand U1203 (N_1203,N_1156,N_1101);
or U1204 (N_1204,N_1179,N_1103);
nand U1205 (N_1205,N_1182,N_1120);
or U1206 (N_1206,N_1111,N_1114);
nand U1207 (N_1207,N_1112,N_1196);
or U1208 (N_1208,N_1115,N_1192);
nand U1209 (N_1209,N_1123,N_1110);
nor U1210 (N_1210,N_1100,N_1152);
xnor U1211 (N_1211,N_1194,N_1145);
nand U1212 (N_1212,N_1137,N_1198);
nand U1213 (N_1213,N_1189,N_1127);
nor U1214 (N_1214,N_1195,N_1176);
xnor U1215 (N_1215,N_1193,N_1148);
nor U1216 (N_1216,N_1118,N_1155);
nand U1217 (N_1217,N_1170,N_1122);
or U1218 (N_1218,N_1187,N_1175);
xnor U1219 (N_1219,N_1188,N_1138);
and U1220 (N_1220,N_1184,N_1134);
or U1221 (N_1221,N_1199,N_1154);
or U1222 (N_1222,N_1167,N_1190);
nor U1223 (N_1223,N_1132,N_1169);
and U1224 (N_1224,N_1130,N_1147);
nand U1225 (N_1225,N_1172,N_1183);
xor U1226 (N_1226,N_1160,N_1173);
and U1227 (N_1227,N_1149,N_1150);
nand U1228 (N_1228,N_1124,N_1121);
and U1229 (N_1229,N_1166,N_1136);
xor U1230 (N_1230,N_1153,N_1159);
nor U1231 (N_1231,N_1181,N_1117);
or U1232 (N_1232,N_1191,N_1178);
and U1233 (N_1233,N_1113,N_1163);
or U1234 (N_1234,N_1161,N_1126);
nand U1235 (N_1235,N_1165,N_1108);
and U1236 (N_1236,N_1139,N_1119);
or U1237 (N_1237,N_1107,N_1129);
and U1238 (N_1238,N_1162,N_1186);
nor U1239 (N_1239,N_1151,N_1164);
and U1240 (N_1240,N_1106,N_1105);
xor U1241 (N_1241,N_1180,N_1141);
xor U1242 (N_1242,N_1174,N_1177);
nor U1243 (N_1243,N_1143,N_1125);
or U1244 (N_1244,N_1133,N_1104);
and U1245 (N_1245,N_1140,N_1144);
or U1246 (N_1246,N_1185,N_1197);
nor U1247 (N_1247,N_1109,N_1158);
nor U1248 (N_1248,N_1146,N_1168);
xnor U1249 (N_1249,N_1128,N_1135);
and U1250 (N_1250,N_1112,N_1158);
or U1251 (N_1251,N_1198,N_1164);
or U1252 (N_1252,N_1185,N_1124);
and U1253 (N_1253,N_1148,N_1132);
xor U1254 (N_1254,N_1110,N_1192);
xnor U1255 (N_1255,N_1160,N_1176);
and U1256 (N_1256,N_1115,N_1117);
nor U1257 (N_1257,N_1169,N_1195);
nand U1258 (N_1258,N_1182,N_1126);
and U1259 (N_1259,N_1159,N_1141);
nor U1260 (N_1260,N_1153,N_1139);
and U1261 (N_1261,N_1105,N_1146);
nand U1262 (N_1262,N_1177,N_1124);
or U1263 (N_1263,N_1164,N_1118);
and U1264 (N_1264,N_1150,N_1138);
xor U1265 (N_1265,N_1116,N_1155);
nand U1266 (N_1266,N_1172,N_1173);
nor U1267 (N_1267,N_1127,N_1138);
nand U1268 (N_1268,N_1187,N_1118);
and U1269 (N_1269,N_1122,N_1128);
nand U1270 (N_1270,N_1147,N_1100);
nand U1271 (N_1271,N_1101,N_1166);
nor U1272 (N_1272,N_1123,N_1150);
and U1273 (N_1273,N_1179,N_1104);
xnor U1274 (N_1274,N_1169,N_1137);
nand U1275 (N_1275,N_1146,N_1175);
xnor U1276 (N_1276,N_1134,N_1194);
or U1277 (N_1277,N_1143,N_1199);
nand U1278 (N_1278,N_1101,N_1142);
and U1279 (N_1279,N_1126,N_1105);
nor U1280 (N_1280,N_1158,N_1147);
or U1281 (N_1281,N_1179,N_1177);
nand U1282 (N_1282,N_1183,N_1198);
xnor U1283 (N_1283,N_1129,N_1137);
or U1284 (N_1284,N_1110,N_1187);
nor U1285 (N_1285,N_1195,N_1115);
nor U1286 (N_1286,N_1177,N_1197);
xnor U1287 (N_1287,N_1192,N_1145);
and U1288 (N_1288,N_1155,N_1180);
nand U1289 (N_1289,N_1164,N_1105);
nand U1290 (N_1290,N_1165,N_1190);
nand U1291 (N_1291,N_1142,N_1135);
or U1292 (N_1292,N_1127,N_1100);
xnor U1293 (N_1293,N_1170,N_1185);
nand U1294 (N_1294,N_1176,N_1179);
nor U1295 (N_1295,N_1153,N_1178);
nand U1296 (N_1296,N_1141,N_1175);
nand U1297 (N_1297,N_1140,N_1181);
nor U1298 (N_1298,N_1192,N_1191);
and U1299 (N_1299,N_1128,N_1186);
nand U1300 (N_1300,N_1206,N_1298);
nor U1301 (N_1301,N_1243,N_1267);
and U1302 (N_1302,N_1226,N_1250);
xnor U1303 (N_1303,N_1284,N_1275);
or U1304 (N_1304,N_1287,N_1205);
nand U1305 (N_1305,N_1263,N_1283);
or U1306 (N_1306,N_1292,N_1214);
or U1307 (N_1307,N_1217,N_1255);
nor U1308 (N_1308,N_1269,N_1264);
nand U1309 (N_1309,N_1208,N_1215);
or U1310 (N_1310,N_1297,N_1222);
xor U1311 (N_1311,N_1220,N_1228);
xor U1312 (N_1312,N_1235,N_1246);
or U1313 (N_1313,N_1234,N_1249);
or U1314 (N_1314,N_1266,N_1259);
and U1315 (N_1315,N_1230,N_1218);
or U1316 (N_1316,N_1211,N_1242);
and U1317 (N_1317,N_1289,N_1247);
nor U1318 (N_1318,N_1207,N_1291);
nor U1319 (N_1319,N_1256,N_1252);
nand U1320 (N_1320,N_1286,N_1271);
nand U1321 (N_1321,N_1257,N_1279);
nand U1322 (N_1322,N_1210,N_1261);
nor U1323 (N_1323,N_1251,N_1212);
nand U1324 (N_1324,N_1233,N_1224);
nor U1325 (N_1325,N_1232,N_1274);
or U1326 (N_1326,N_1293,N_1202);
nand U1327 (N_1327,N_1245,N_1231);
xnor U1328 (N_1328,N_1236,N_1288);
xor U1329 (N_1329,N_1273,N_1280);
nor U1330 (N_1330,N_1201,N_1258);
nand U1331 (N_1331,N_1260,N_1270);
xnor U1332 (N_1332,N_1200,N_1248);
or U1333 (N_1333,N_1204,N_1262);
or U1334 (N_1334,N_1239,N_1296);
xor U1335 (N_1335,N_1281,N_1254);
nand U1336 (N_1336,N_1294,N_1238);
nor U1337 (N_1337,N_1216,N_1229);
or U1338 (N_1338,N_1290,N_1278);
nand U1339 (N_1339,N_1223,N_1237);
or U1340 (N_1340,N_1295,N_1265);
nand U1341 (N_1341,N_1241,N_1209);
nor U1342 (N_1342,N_1253,N_1276);
or U1343 (N_1343,N_1277,N_1221);
and U1344 (N_1344,N_1203,N_1225);
and U1345 (N_1345,N_1272,N_1213);
xnor U1346 (N_1346,N_1285,N_1282);
or U1347 (N_1347,N_1219,N_1299);
and U1348 (N_1348,N_1268,N_1244);
nand U1349 (N_1349,N_1240,N_1227);
nand U1350 (N_1350,N_1253,N_1218);
and U1351 (N_1351,N_1291,N_1227);
or U1352 (N_1352,N_1253,N_1231);
and U1353 (N_1353,N_1299,N_1251);
or U1354 (N_1354,N_1293,N_1286);
xor U1355 (N_1355,N_1217,N_1230);
and U1356 (N_1356,N_1260,N_1220);
and U1357 (N_1357,N_1213,N_1261);
nand U1358 (N_1358,N_1288,N_1219);
nor U1359 (N_1359,N_1248,N_1228);
and U1360 (N_1360,N_1297,N_1221);
and U1361 (N_1361,N_1210,N_1269);
xor U1362 (N_1362,N_1230,N_1207);
or U1363 (N_1363,N_1221,N_1245);
nand U1364 (N_1364,N_1209,N_1254);
xor U1365 (N_1365,N_1234,N_1296);
or U1366 (N_1366,N_1229,N_1281);
xnor U1367 (N_1367,N_1280,N_1275);
xnor U1368 (N_1368,N_1201,N_1251);
nor U1369 (N_1369,N_1201,N_1267);
and U1370 (N_1370,N_1241,N_1201);
or U1371 (N_1371,N_1250,N_1297);
and U1372 (N_1372,N_1232,N_1231);
xnor U1373 (N_1373,N_1244,N_1235);
nor U1374 (N_1374,N_1255,N_1235);
xnor U1375 (N_1375,N_1259,N_1232);
xnor U1376 (N_1376,N_1267,N_1264);
nor U1377 (N_1377,N_1264,N_1244);
or U1378 (N_1378,N_1293,N_1282);
nand U1379 (N_1379,N_1293,N_1266);
nand U1380 (N_1380,N_1210,N_1205);
or U1381 (N_1381,N_1275,N_1262);
or U1382 (N_1382,N_1235,N_1282);
nor U1383 (N_1383,N_1290,N_1228);
and U1384 (N_1384,N_1202,N_1269);
xor U1385 (N_1385,N_1233,N_1287);
nand U1386 (N_1386,N_1228,N_1200);
or U1387 (N_1387,N_1243,N_1289);
nor U1388 (N_1388,N_1256,N_1209);
and U1389 (N_1389,N_1297,N_1267);
and U1390 (N_1390,N_1269,N_1259);
nand U1391 (N_1391,N_1214,N_1278);
and U1392 (N_1392,N_1269,N_1214);
nor U1393 (N_1393,N_1298,N_1229);
and U1394 (N_1394,N_1205,N_1255);
xor U1395 (N_1395,N_1299,N_1267);
nor U1396 (N_1396,N_1269,N_1216);
and U1397 (N_1397,N_1251,N_1248);
nor U1398 (N_1398,N_1282,N_1264);
nand U1399 (N_1399,N_1266,N_1299);
nand U1400 (N_1400,N_1366,N_1318);
and U1401 (N_1401,N_1337,N_1320);
nand U1402 (N_1402,N_1309,N_1394);
or U1403 (N_1403,N_1356,N_1321);
or U1404 (N_1404,N_1310,N_1391);
or U1405 (N_1405,N_1326,N_1341);
or U1406 (N_1406,N_1354,N_1371);
and U1407 (N_1407,N_1399,N_1316);
nand U1408 (N_1408,N_1355,N_1330);
or U1409 (N_1409,N_1358,N_1352);
xnor U1410 (N_1410,N_1385,N_1300);
and U1411 (N_1411,N_1301,N_1389);
nor U1412 (N_1412,N_1350,N_1357);
xor U1413 (N_1413,N_1395,N_1361);
xnor U1414 (N_1414,N_1331,N_1390);
or U1415 (N_1415,N_1353,N_1377);
nor U1416 (N_1416,N_1322,N_1374);
or U1417 (N_1417,N_1376,N_1378);
or U1418 (N_1418,N_1343,N_1367);
xor U1419 (N_1419,N_1311,N_1372);
and U1420 (N_1420,N_1340,N_1347);
nor U1421 (N_1421,N_1327,N_1370);
and U1422 (N_1422,N_1303,N_1312);
or U1423 (N_1423,N_1375,N_1346);
nor U1424 (N_1424,N_1369,N_1387);
nor U1425 (N_1425,N_1332,N_1348);
nand U1426 (N_1426,N_1317,N_1319);
and U1427 (N_1427,N_1365,N_1344);
and U1428 (N_1428,N_1373,N_1313);
or U1429 (N_1429,N_1363,N_1383);
nand U1430 (N_1430,N_1392,N_1307);
nand U1431 (N_1431,N_1328,N_1384);
nand U1432 (N_1432,N_1368,N_1323);
nand U1433 (N_1433,N_1388,N_1349);
and U1434 (N_1434,N_1345,N_1315);
nor U1435 (N_1435,N_1336,N_1306);
or U1436 (N_1436,N_1379,N_1325);
xor U1437 (N_1437,N_1339,N_1302);
and U1438 (N_1438,N_1335,N_1351);
or U1439 (N_1439,N_1393,N_1381);
and U1440 (N_1440,N_1397,N_1364);
nor U1441 (N_1441,N_1396,N_1362);
nand U1442 (N_1442,N_1304,N_1338);
and U1443 (N_1443,N_1333,N_1360);
nand U1444 (N_1444,N_1329,N_1382);
or U1445 (N_1445,N_1314,N_1386);
nor U1446 (N_1446,N_1359,N_1334);
or U1447 (N_1447,N_1324,N_1305);
and U1448 (N_1448,N_1308,N_1398);
nand U1449 (N_1449,N_1342,N_1380);
nor U1450 (N_1450,N_1303,N_1364);
and U1451 (N_1451,N_1356,N_1303);
xnor U1452 (N_1452,N_1309,N_1361);
or U1453 (N_1453,N_1334,N_1313);
xnor U1454 (N_1454,N_1343,N_1399);
nor U1455 (N_1455,N_1335,N_1374);
and U1456 (N_1456,N_1311,N_1315);
nand U1457 (N_1457,N_1334,N_1386);
xor U1458 (N_1458,N_1373,N_1377);
or U1459 (N_1459,N_1389,N_1304);
nand U1460 (N_1460,N_1313,N_1304);
xnor U1461 (N_1461,N_1356,N_1392);
nor U1462 (N_1462,N_1348,N_1312);
and U1463 (N_1463,N_1345,N_1313);
nor U1464 (N_1464,N_1311,N_1380);
or U1465 (N_1465,N_1365,N_1371);
or U1466 (N_1466,N_1374,N_1365);
xnor U1467 (N_1467,N_1362,N_1367);
or U1468 (N_1468,N_1369,N_1335);
or U1469 (N_1469,N_1355,N_1332);
nand U1470 (N_1470,N_1399,N_1306);
nand U1471 (N_1471,N_1381,N_1348);
nor U1472 (N_1472,N_1388,N_1329);
xnor U1473 (N_1473,N_1368,N_1315);
xnor U1474 (N_1474,N_1345,N_1338);
and U1475 (N_1475,N_1317,N_1306);
nor U1476 (N_1476,N_1322,N_1315);
or U1477 (N_1477,N_1359,N_1365);
nor U1478 (N_1478,N_1346,N_1387);
xor U1479 (N_1479,N_1389,N_1361);
or U1480 (N_1480,N_1365,N_1369);
xnor U1481 (N_1481,N_1359,N_1384);
or U1482 (N_1482,N_1326,N_1390);
nand U1483 (N_1483,N_1338,N_1347);
and U1484 (N_1484,N_1373,N_1379);
xor U1485 (N_1485,N_1396,N_1398);
or U1486 (N_1486,N_1331,N_1347);
and U1487 (N_1487,N_1325,N_1320);
nand U1488 (N_1488,N_1395,N_1307);
and U1489 (N_1489,N_1391,N_1317);
xnor U1490 (N_1490,N_1346,N_1389);
nor U1491 (N_1491,N_1353,N_1372);
nor U1492 (N_1492,N_1363,N_1320);
or U1493 (N_1493,N_1329,N_1308);
or U1494 (N_1494,N_1394,N_1322);
xor U1495 (N_1495,N_1394,N_1374);
nor U1496 (N_1496,N_1335,N_1308);
and U1497 (N_1497,N_1359,N_1376);
or U1498 (N_1498,N_1304,N_1362);
or U1499 (N_1499,N_1353,N_1304);
nor U1500 (N_1500,N_1476,N_1457);
nor U1501 (N_1501,N_1489,N_1480);
or U1502 (N_1502,N_1483,N_1421);
nor U1503 (N_1503,N_1410,N_1435);
xnor U1504 (N_1504,N_1484,N_1487);
nor U1505 (N_1505,N_1430,N_1481);
nor U1506 (N_1506,N_1418,N_1458);
and U1507 (N_1507,N_1467,N_1447);
nor U1508 (N_1508,N_1477,N_1451);
nand U1509 (N_1509,N_1443,N_1462);
and U1510 (N_1510,N_1474,N_1422);
or U1511 (N_1511,N_1479,N_1423);
nor U1512 (N_1512,N_1468,N_1415);
xor U1513 (N_1513,N_1436,N_1411);
nor U1514 (N_1514,N_1419,N_1434);
or U1515 (N_1515,N_1472,N_1453);
and U1516 (N_1516,N_1488,N_1448);
and U1517 (N_1517,N_1405,N_1470);
or U1518 (N_1518,N_1424,N_1478);
nand U1519 (N_1519,N_1420,N_1401);
xor U1520 (N_1520,N_1409,N_1444);
nand U1521 (N_1521,N_1459,N_1417);
and U1522 (N_1522,N_1486,N_1490);
nor U1523 (N_1523,N_1456,N_1432);
xnor U1524 (N_1524,N_1455,N_1499);
nor U1525 (N_1525,N_1406,N_1441);
xor U1526 (N_1526,N_1429,N_1408);
nor U1527 (N_1527,N_1439,N_1407);
and U1528 (N_1528,N_1461,N_1498);
xnor U1529 (N_1529,N_1492,N_1445);
xor U1530 (N_1530,N_1452,N_1428);
xnor U1531 (N_1531,N_1460,N_1425);
and U1532 (N_1532,N_1475,N_1482);
or U1533 (N_1533,N_1449,N_1496);
xor U1534 (N_1534,N_1463,N_1413);
xnor U1535 (N_1535,N_1412,N_1442);
nand U1536 (N_1536,N_1433,N_1495);
or U1537 (N_1537,N_1431,N_1438);
or U1538 (N_1538,N_1473,N_1426);
and U1539 (N_1539,N_1485,N_1437);
nor U1540 (N_1540,N_1491,N_1454);
nor U1541 (N_1541,N_1427,N_1416);
or U1542 (N_1542,N_1471,N_1400);
nor U1543 (N_1543,N_1404,N_1450);
xor U1544 (N_1544,N_1440,N_1466);
and U1545 (N_1545,N_1493,N_1465);
nand U1546 (N_1546,N_1494,N_1464);
xnor U1547 (N_1547,N_1446,N_1414);
nand U1548 (N_1548,N_1402,N_1469);
or U1549 (N_1549,N_1403,N_1497);
nor U1550 (N_1550,N_1492,N_1463);
nand U1551 (N_1551,N_1498,N_1479);
and U1552 (N_1552,N_1466,N_1459);
nor U1553 (N_1553,N_1496,N_1480);
xnor U1554 (N_1554,N_1448,N_1423);
and U1555 (N_1555,N_1466,N_1494);
nand U1556 (N_1556,N_1425,N_1492);
xor U1557 (N_1557,N_1459,N_1400);
nand U1558 (N_1558,N_1467,N_1470);
or U1559 (N_1559,N_1460,N_1430);
and U1560 (N_1560,N_1492,N_1426);
and U1561 (N_1561,N_1467,N_1456);
or U1562 (N_1562,N_1443,N_1460);
xnor U1563 (N_1563,N_1428,N_1406);
or U1564 (N_1564,N_1454,N_1403);
or U1565 (N_1565,N_1459,N_1490);
xor U1566 (N_1566,N_1456,N_1452);
nor U1567 (N_1567,N_1488,N_1451);
nand U1568 (N_1568,N_1422,N_1453);
nor U1569 (N_1569,N_1429,N_1445);
nor U1570 (N_1570,N_1488,N_1443);
xor U1571 (N_1571,N_1441,N_1420);
or U1572 (N_1572,N_1428,N_1427);
and U1573 (N_1573,N_1408,N_1426);
and U1574 (N_1574,N_1429,N_1451);
xor U1575 (N_1575,N_1491,N_1487);
and U1576 (N_1576,N_1474,N_1461);
nand U1577 (N_1577,N_1458,N_1443);
xor U1578 (N_1578,N_1416,N_1429);
nand U1579 (N_1579,N_1428,N_1404);
nor U1580 (N_1580,N_1465,N_1499);
xor U1581 (N_1581,N_1484,N_1473);
and U1582 (N_1582,N_1492,N_1443);
or U1583 (N_1583,N_1412,N_1422);
xor U1584 (N_1584,N_1459,N_1452);
nand U1585 (N_1585,N_1434,N_1435);
nand U1586 (N_1586,N_1401,N_1454);
and U1587 (N_1587,N_1463,N_1414);
xnor U1588 (N_1588,N_1442,N_1494);
xnor U1589 (N_1589,N_1457,N_1446);
xnor U1590 (N_1590,N_1447,N_1456);
xnor U1591 (N_1591,N_1417,N_1494);
and U1592 (N_1592,N_1472,N_1435);
nor U1593 (N_1593,N_1441,N_1481);
nor U1594 (N_1594,N_1404,N_1433);
nand U1595 (N_1595,N_1403,N_1427);
xnor U1596 (N_1596,N_1458,N_1457);
xor U1597 (N_1597,N_1443,N_1451);
xnor U1598 (N_1598,N_1463,N_1480);
xnor U1599 (N_1599,N_1460,N_1463);
or U1600 (N_1600,N_1536,N_1524);
or U1601 (N_1601,N_1578,N_1541);
nand U1602 (N_1602,N_1511,N_1573);
or U1603 (N_1603,N_1592,N_1551);
nand U1604 (N_1604,N_1527,N_1513);
and U1605 (N_1605,N_1520,N_1572);
or U1606 (N_1606,N_1574,N_1575);
or U1607 (N_1607,N_1502,N_1518);
nor U1608 (N_1608,N_1597,N_1539);
nor U1609 (N_1609,N_1540,N_1555);
and U1610 (N_1610,N_1567,N_1598);
and U1611 (N_1611,N_1554,N_1558);
or U1612 (N_1612,N_1552,N_1534);
nor U1613 (N_1613,N_1562,N_1547);
nand U1614 (N_1614,N_1508,N_1505);
and U1615 (N_1615,N_1564,N_1589);
or U1616 (N_1616,N_1588,N_1548);
nand U1617 (N_1617,N_1537,N_1535);
nand U1618 (N_1618,N_1501,N_1563);
or U1619 (N_1619,N_1538,N_1561);
xnor U1620 (N_1620,N_1512,N_1531);
nand U1621 (N_1621,N_1569,N_1556);
nand U1622 (N_1622,N_1514,N_1521);
or U1623 (N_1623,N_1526,N_1585);
and U1624 (N_1624,N_1533,N_1580);
or U1625 (N_1625,N_1593,N_1543);
nand U1626 (N_1626,N_1532,N_1509);
or U1627 (N_1627,N_1599,N_1510);
xor U1628 (N_1628,N_1581,N_1550);
nand U1629 (N_1629,N_1528,N_1559);
nor U1630 (N_1630,N_1557,N_1586);
or U1631 (N_1631,N_1517,N_1544);
nand U1632 (N_1632,N_1570,N_1591);
nor U1633 (N_1633,N_1542,N_1568);
nand U1634 (N_1634,N_1507,N_1549);
nor U1635 (N_1635,N_1576,N_1504);
nand U1636 (N_1636,N_1500,N_1566);
or U1637 (N_1637,N_1553,N_1595);
and U1638 (N_1638,N_1560,N_1596);
nor U1639 (N_1639,N_1516,N_1582);
or U1640 (N_1640,N_1545,N_1515);
or U1641 (N_1641,N_1546,N_1590);
nand U1642 (N_1642,N_1530,N_1503);
nor U1643 (N_1643,N_1594,N_1571);
xor U1644 (N_1644,N_1579,N_1525);
nand U1645 (N_1645,N_1565,N_1577);
xor U1646 (N_1646,N_1522,N_1587);
and U1647 (N_1647,N_1519,N_1583);
xnor U1648 (N_1648,N_1584,N_1529);
and U1649 (N_1649,N_1506,N_1523);
and U1650 (N_1650,N_1589,N_1598);
nand U1651 (N_1651,N_1548,N_1505);
nor U1652 (N_1652,N_1539,N_1542);
xnor U1653 (N_1653,N_1540,N_1554);
nand U1654 (N_1654,N_1520,N_1536);
nand U1655 (N_1655,N_1533,N_1521);
and U1656 (N_1656,N_1585,N_1558);
nor U1657 (N_1657,N_1535,N_1543);
nor U1658 (N_1658,N_1577,N_1522);
xnor U1659 (N_1659,N_1589,N_1531);
xor U1660 (N_1660,N_1535,N_1585);
nand U1661 (N_1661,N_1512,N_1557);
xnor U1662 (N_1662,N_1573,N_1549);
nor U1663 (N_1663,N_1565,N_1582);
and U1664 (N_1664,N_1547,N_1544);
nor U1665 (N_1665,N_1529,N_1502);
xnor U1666 (N_1666,N_1576,N_1512);
and U1667 (N_1667,N_1513,N_1508);
nand U1668 (N_1668,N_1511,N_1564);
xnor U1669 (N_1669,N_1520,N_1579);
and U1670 (N_1670,N_1572,N_1525);
and U1671 (N_1671,N_1596,N_1572);
nor U1672 (N_1672,N_1583,N_1574);
and U1673 (N_1673,N_1567,N_1529);
nand U1674 (N_1674,N_1554,N_1589);
nor U1675 (N_1675,N_1593,N_1564);
and U1676 (N_1676,N_1578,N_1500);
and U1677 (N_1677,N_1504,N_1560);
xnor U1678 (N_1678,N_1582,N_1593);
nand U1679 (N_1679,N_1550,N_1562);
xnor U1680 (N_1680,N_1502,N_1565);
xnor U1681 (N_1681,N_1509,N_1560);
nor U1682 (N_1682,N_1529,N_1580);
or U1683 (N_1683,N_1576,N_1542);
xnor U1684 (N_1684,N_1530,N_1537);
xor U1685 (N_1685,N_1525,N_1510);
nand U1686 (N_1686,N_1541,N_1546);
nand U1687 (N_1687,N_1510,N_1598);
nor U1688 (N_1688,N_1558,N_1534);
and U1689 (N_1689,N_1544,N_1509);
nand U1690 (N_1690,N_1557,N_1567);
nand U1691 (N_1691,N_1525,N_1590);
or U1692 (N_1692,N_1511,N_1535);
nand U1693 (N_1693,N_1521,N_1587);
nor U1694 (N_1694,N_1565,N_1544);
nand U1695 (N_1695,N_1581,N_1536);
nand U1696 (N_1696,N_1556,N_1511);
and U1697 (N_1697,N_1507,N_1515);
or U1698 (N_1698,N_1589,N_1518);
xor U1699 (N_1699,N_1587,N_1534);
nor U1700 (N_1700,N_1657,N_1656);
nand U1701 (N_1701,N_1625,N_1660);
xnor U1702 (N_1702,N_1659,N_1681);
nor U1703 (N_1703,N_1665,N_1687);
and U1704 (N_1704,N_1662,N_1607);
and U1705 (N_1705,N_1667,N_1639);
nand U1706 (N_1706,N_1696,N_1683);
xnor U1707 (N_1707,N_1692,N_1644);
nor U1708 (N_1708,N_1632,N_1648);
nand U1709 (N_1709,N_1626,N_1614);
and U1710 (N_1710,N_1675,N_1610);
nor U1711 (N_1711,N_1688,N_1658);
and U1712 (N_1712,N_1690,N_1628);
nor U1713 (N_1713,N_1673,N_1602);
xor U1714 (N_1714,N_1682,N_1642);
and U1715 (N_1715,N_1651,N_1671);
nor U1716 (N_1716,N_1685,N_1645);
and U1717 (N_1717,N_1640,N_1684);
nor U1718 (N_1718,N_1679,N_1633);
and U1719 (N_1719,N_1606,N_1676);
or U1720 (N_1720,N_1641,N_1612);
xor U1721 (N_1721,N_1646,N_1624);
xor U1722 (N_1722,N_1609,N_1619);
and U1723 (N_1723,N_1617,N_1668);
nand U1724 (N_1724,N_1649,N_1647);
nand U1725 (N_1725,N_1672,N_1680);
nand U1726 (N_1726,N_1669,N_1652);
and U1727 (N_1727,N_1661,N_1627);
xnor U1728 (N_1728,N_1699,N_1697);
xor U1729 (N_1729,N_1635,N_1616);
nor U1730 (N_1730,N_1637,N_1674);
nor U1731 (N_1731,N_1663,N_1613);
nor U1732 (N_1732,N_1601,N_1608);
and U1733 (N_1733,N_1670,N_1621);
nor U1734 (N_1734,N_1664,N_1693);
nor U1735 (N_1735,N_1623,N_1677);
nor U1736 (N_1736,N_1691,N_1666);
xnor U1737 (N_1737,N_1678,N_1655);
or U1738 (N_1738,N_1694,N_1698);
xor U1739 (N_1739,N_1634,N_1603);
and U1740 (N_1740,N_1611,N_1605);
and U1741 (N_1741,N_1604,N_1654);
and U1742 (N_1742,N_1618,N_1695);
and U1743 (N_1743,N_1636,N_1629);
and U1744 (N_1744,N_1643,N_1630);
nand U1745 (N_1745,N_1622,N_1689);
and U1746 (N_1746,N_1638,N_1653);
nor U1747 (N_1747,N_1600,N_1631);
nand U1748 (N_1748,N_1686,N_1620);
xor U1749 (N_1749,N_1650,N_1615);
xor U1750 (N_1750,N_1627,N_1637);
xnor U1751 (N_1751,N_1664,N_1619);
or U1752 (N_1752,N_1699,N_1654);
or U1753 (N_1753,N_1639,N_1629);
or U1754 (N_1754,N_1676,N_1674);
nand U1755 (N_1755,N_1665,N_1623);
and U1756 (N_1756,N_1631,N_1661);
nand U1757 (N_1757,N_1635,N_1640);
nand U1758 (N_1758,N_1669,N_1658);
or U1759 (N_1759,N_1604,N_1697);
nand U1760 (N_1760,N_1613,N_1626);
nor U1761 (N_1761,N_1624,N_1696);
nand U1762 (N_1762,N_1687,N_1656);
xor U1763 (N_1763,N_1644,N_1659);
nor U1764 (N_1764,N_1674,N_1603);
nor U1765 (N_1765,N_1673,N_1669);
and U1766 (N_1766,N_1626,N_1601);
and U1767 (N_1767,N_1625,N_1612);
or U1768 (N_1768,N_1650,N_1698);
xor U1769 (N_1769,N_1650,N_1618);
nor U1770 (N_1770,N_1696,N_1688);
nor U1771 (N_1771,N_1685,N_1601);
and U1772 (N_1772,N_1629,N_1645);
and U1773 (N_1773,N_1605,N_1604);
and U1774 (N_1774,N_1616,N_1678);
nor U1775 (N_1775,N_1691,N_1601);
nor U1776 (N_1776,N_1664,N_1623);
and U1777 (N_1777,N_1641,N_1673);
and U1778 (N_1778,N_1680,N_1637);
and U1779 (N_1779,N_1624,N_1686);
and U1780 (N_1780,N_1624,N_1657);
nor U1781 (N_1781,N_1645,N_1682);
nor U1782 (N_1782,N_1659,N_1621);
xnor U1783 (N_1783,N_1665,N_1605);
and U1784 (N_1784,N_1653,N_1650);
xnor U1785 (N_1785,N_1662,N_1654);
and U1786 (N_1786,N_1644,N_1630);
and U1787 (N_1787,N_1636,N_1666);
xnor U1788 (N_1788,N_1617,N_1686);
xor U1789 (N_1789,N_1661,N_1604);
nor U1790 (N_1790,N_1605,N_1644);
xnor U1791 (N_1791,N_1659,N_1691);
or U1792 (N_1792,N_1616,N_1686);
nand U1793 (N_1793,N_1616,N_1627);
and U1794 (N_1794,N_1610,N_1617);
xor U1795 (N_1795,N_1692,N_1651);
or U1796 (N_1796,N_1629,N_1654);
nand U1797 (N_1797,N_1618,N_1660);
and U1798 (N_1798,N_1645,N_1614);
nand U1799 (N_1799,N_1600,N_1625);
nor U1800 (N_1800,N_1718,N_1728);
nor U1801 (N_1801,N_1766,N_1713);
nand U1802 (N_1802,N_1717,N_1705);
or U1803 (N_1803,N_1744,N_1759);
xor U1804 (N_1804,N_1784,N_1769);
xnor U1805 (N_1805,N_1754,N_1781);
xnor U1806 (N_1806,N_1799,N_1721);
and U1807 (N_1807,N_1730,N_1733);
and U1808 (N_1808,N_1719,N_1782);
nand U1809 (N_1809,N_1746,N_1702);
and U1810 (N_1810,N_1726,N_1793);
or U1811 (N_1811,N_1732,N_1776);
or U1812 (N_1812,N_1724,N_1780);
and U1813 (N_1813,N_1778,N_1761);
and U1814 (N_1814,N_1756,N_1758);
nor U1815 (N_1815,N_1779,N_1790);
and U1816 (N_1816,N_1723,N_1720);
and U1817 (N_1817,N_1704,N_1789);
or U1818 (N_1818,N_1787,N_1734);
or U1819 (N_1819,N_1785,N_1712);
nor U1820 (N_1820,N_1749,N_1716);
nand U1821 (N_1821,N_1792,N_1707);
nand U1822 (N_1822,N_1764,N_1755);
and U1823 (N_1823,N_1773,N_1786);
or U1824 (N_1824,N_1738,N_1763);
nor U1825 (N_1825,N_1715,N_1747);
or U1826 (N_1826,N_1736,N_1760);
or U1827 (N_1827,N_1701,N_1741);
and U1828 (N_1828,N_1714,N_1731);
xnor U1829 (N_1829,N_1703,N_1757);
nand U1830 (N_1830,N_1706,N_1752);
nor U1831 (N_1831,N_1709,N_1700);
or U1832 (N_1832,N_1751,N_1725);
nand U1833 (N_1833,N_1768,N_1767);
xor U1834 (N_1834,N_1753,N_1798);
nand U1835 (N_1835,N_1735,N_1771);
xnor U1836 (N_1836,N_1729,N_1740);
nand U1837 (N_1837,N_1770,N_1748);
and U1838 (N_1838,N_1710,N_1727);
or U1839 (N_1839,N_1708,N_1765);
nor U1840 (N_1840,N_1772,N_1745);
nor U1841 (N_1841,N_1796,N_1791);
nand U1842 (N_1842,N_1795,N_1737);
nor U1843 (N_1843,N_1739,N_1774);
or U1844 (N_1844,N_1777,N_1742);
xor U1845 (N_1845,N_1711,N_1743);
and U1846 (N_1846,N_1788,N_1783);
nor U1847 (N_1847,N_1794,N_1775);
and U1848 (N_1848,N_1762,N_1797);
nor U1849 (N_1849,N_1722,N_1750);
or U1850 (N_1850,N_1792,N_1756);
and U1851 (N_1851,N_1734,N_1779);
nand U1852 (N_1852,N_1796,N_1701);
nand U1853 (N_1853,N_1747,N_1752);
or U1854 (N_1854,N_1799,N_1778);
and U1855 (N_1855,N_1701,N_1702);
nor U1856 (N_1856,N_1767,N_1764);
nor U1857 (N_1857,N_1787,N_1793);
nand U1858 (N_1858,N_1708,N_1717);
nand U1859 (N_1859,N_1797,N_1776);
xor U1860 (N_1860,N_1785,N_1734);
and U1861 (N_1861,N_1763,N_1746);
or U1862 (N_1862,N_1717,N_1775);
nor U1863 (N_1863,N_1712,N_1756);
nand U1864 (N_1864,N_1748,N_1700);
and U1865 (N_1865,N_1777,N_1757);
xor U1866 (N_1866,N_1741,N_1778);
and U1867 (N_1867,N_1717,N_1748);
nor U1868 (N_1868,N_1799,N_1760);
nand U1869 (N_1869,N_1702,N_1713);
nand U1870 (N_1870,N_1764,N_1796);
xor U1871 (N_1871,N_1718,N_1716);
nand U1872 (N_1872,N_1752,N_1786);
and U1873 (N_1873,N_1770,N_1711);
nor U1874 (N_1874,N_1716,N_1786);
and U1875 (N_1875,N_1701,N_1715);
xnor U1876 (N_1876,N_1727,N_1722);
or U1877 (N_1877,N_1743,N_1784);
nand U1878 (N_1878,N_1747,N_1731);
nand U1879 (N_1879,N_1738,N_1742);
nor U1880 (N_1880,N_1758,N_1701);
and U1881 (N_1881,N_1789,N_1784);
xor U1882 (N_1882,N_1702,N_1794);
xnor U1883 (N_1883,N_1769,N_1766);
nor U1884 (N_1884,N_1730,N_1700);
and U1885 (N_1885,N_1706,N_1717);
or U1886 (N_1886,N_1716,N_1766);
or U1887 (N_1887,N_1724,N_1794);
nor U1888 (N_1888,N_1764,N_1766);
nand U1889 (N_1889,N_1799,N_1765);
or U1890 (N_1890,N_1719,N_1717);
nor U1891 (N_1891,N_1737,N_1721);
nor U1892 (N_1892,N_1779,N_1711);
nor U1893 (N_1893,N_1733,N_1763);
nand U1894 (N_1894,N_1797,N_1708);
and U1895 (N_1895,N_1756,N_1714);
xnor U1896 (N_1896,N_1767,N_1726);
xor U1897 (N_1897,N_1724,N_1751);
nand U1898 (N_1898,N_1726,N_1732);
nor U1899 (N_1899,N_1783,N_1711);
nand U1900 (N_1900,N_1894,N_1811);
and U1901 (N_1901,N_1816,N_1885);
nor U1902 (N_1902,N_1891,N_1876);
and U1903 (N_1903,N_1874,N_1849);
nand U1904 (N_1904,N_1820,N_1817);
xnor U1905 (N_1905,N_1837,N_1879);
nor U1906 (N_1906,N_1800,N_1802);
nor U1907 (N_1907,N_1805,N_1889);
nor U1908 (N_1908,N_1808,N_1896);
nor U1909 (N_1909,N_1856,N_1886);
nor U1910 (N_1910,N_1851,N_1826);
nand U1911 (N_1911,N_1899,N_1861);
nor U1912 (N_1912,N_1877,N_1848);
nor U1913 (N_1913,N_1884,N_1863);
nand U1914 (N_1914,N_1893,N_1853);
and U1915 (N_1915,N_1892,N_1841);
nand U1916 (N_1916,N_1806,N_1898);
and U1917 (N_1917,N_1868,N_1870);
nor U1918 (N_1918,N_1833,N_1813);
nand U1919 (N_1919,N_1840,N_1854);
nand U1920 (N_1920,N_1850,N_1895);
nor U1921 (N_1921,N_1875,N_1823);
and U1922 (N_1922,N_1821,N_1871);
or U1923 (N_1923,N_1882,N_1869);
or U1924 (N_1924,N_1838,N_1847);
or U1925 (N_1925,N_1859,N_1835);
nand U1926 (N_1926,N_1810,N_1839);
nor U1927 (N_1927,N_1887,N_1852);
or U1928 (N_1928,N_1880,N_1827);
nand U1929 (N_1929,N_1881,N_1801);
nor U1930 (N_1930,N_1807,N_1819);
or U1931 (N_1931,N_1832,N_1836);
nor U1932 (N_1932,N_1834,N_1829);
and U1933 (N_1933,N_1825,N_1814);
xnor U1934 (N_1934,N_1842,N_1866);
nand U1935 (N_1935,N_1843,N_1888);
and U1936 (N_1936,N_1864,N_1812);
and U1937 (N_1937,N_1822,N_1844);
nor U1938 (N_1938,N_1824,N_1831);
xnor U1939 (N_1939,N_1815,N_1830);
and U1940 (N_1940,N_1858,N_1860);
and U1941 (N_1941,N_1890,N_1897);
and U1942 (N_1942,N_1873,N_1883);
nand U1943 (N_1943,N_1803,N_1865);
nand U1944 (N_1944,N_1804,N_1878);
nor U1945 (N_1945,N_1867,N_1846);
and U1946 (N_1946,N_1862,N_1818);
or U1947 (N_1947,N_1828,N_1809);
nand U1948 (N_1948,N_1845,N_1872);
xor U1949 (N_1949,N_1857,N_1855);
nor U1950 (N_1950,N_1831,N_1841);
nor U1951 (N_1951,N_1862,N_1819);
nor U1952 (N_1952,N_1820,N_1832);
nor U1953 (N_1953,N_1853,N_1808);
xnor U1954 (N_1954,N_1893,N_1854);
nand U1955 (N_1955,N_1855,N_1844);
xnor U1956 (N_1956,N_1891,N_1833);
or U1957 (N_1957,N_1809,N_1860);
or U1958 (N_1958,N_1865,N_1838);
nor U1959 (N_1959,N_1868,N_1875);
or U1960 (N_1960,N_1882,N_1825);
xnor U1961 (N_1961,N_1856,N_1897);
nor U1962 (N_1962,N_1873,N_1870);
and U1963 (N_1963,N_1860,N_1800);
nand U1964 (N_1964,N_1873,N_1866);
xnor U1965 (N_1965,N_1824,N_1826);
and U1966 (N_1966,N_1873,N_1865);
xor U1967 (N_1967,N_1886,N_1888);
nor U1968 (N_1968,N_1831,N_1807);
xnor U1969 (N_1969,N_1836,N_1831);
and U1970 (N_1970,N_1880,N_1885);
xnor U1971 (N_1971,N_1890,N_1889);
or U1972 (N_1972,N_1827,N_1889);
nor U1973 (N_1973,N_1875,N_1888);
or U1974 (N_1974,N_1852,N_1811);
nor U1975 (N_1975,N_1894,N_1802);
xnor U1976 (N_1976,N_1834,N_1807);
nor U1977 (N_1977,N_1844,N_1817);
nand U1978 (N_1978,N_1826,N_1886);
nand U1979 (N_1979,N_1856,N_1891);
nor U1980 (N_1980,N_1861,N_1897);
and U1981 (N_1981,N_1840,N_1818);
nand U1982 (N_1982,N_1892,N_1812);
nor U1983 (N_1983,N_1835,N_1821);
xor U1984 (N_1984,N_1825,N_1817);
nand U1985 (N_1985,N_1871,N_1862);
or U1986 (N_1986,N_1856,N_1824);
nor U1987 (N_1987,N_1894,N_1845);
nor U1988 (N_1988,N_1802,N_1882);
nand U1989 (N_1989,N_1879,N_1876);
xnor U1990 (N_1990,N_1811,N_1843);
and U1991 (N_1991,N_1801,N_1886);
or U1992 (N_1992,N_1817,N_1860);
or U1993 (N_1993,N_1863,N_1810);
or U1994 (N_1994,N_1889,N_1851);
and U1995 (N_1995,N_1830,N_1850);
xnor U1996 (N_1996,N_1871,N_1807);
or U1997 (N_1997,N_1820,N_1870);
nand U1998 (N_1998,N_1814,N_1895);
nor U1999 (N_1999,N_1861,N_1883);
nor U2000 (N_2000,N_1950,N_1969);
nor U2001 (N_2001,N_1933,N_1949);
nand U2002 (N_2002,N_1998,N_1912);
or U2003 (N_2003,N_1945,N_1960);
or U2004 (N_2004,N_1932,N_1973);
xor U2005 (N_2005,N_1948,N_1903);
and U2006 (N_2006,N_1916,N_1935);
nand U2007 (N_2007,N_1990,N_1989);
and U2008 (N_2008,N_1909,N_1914);
nand U2009 (N_2009,N_1992,N_1936);
nand U2010 (N_2010,N_1964,N_1910);
nand U2011 (N_2011,N_1984,N_1927);
or U2012 (N_2012,N_1901,N_1962);
nand U2013 (N_2013,N_1965,N_1955);
and U2014 (N_2014,N_1941,N_1946);
nor U2015 (N_2015,N_1907,N_1956);
or U2016 (N_2016,N_1974,N_1931);
or U2017 (N_2017,N_1953,N_1900);
and U2018 (N_2018,N_1970,N_1959);
nand U2019 (N_2019,N_1966,N_1934);
nor U2020 (N_2020,N_1917,N_1938);
and U2021 (N_2021,N_1923,N_1981);
or U2022 (N_2022,N_1993,N_1921);
xnor U2023 (N_2023,N_1919,N_1928);
nand U2024 (N_2024,N_1913,N_1978);
xnor U2025 (N_2025,N_1952,N_1999);
nor U2026 (N_2026,N_1991,N_1939);
or U2027 (N_2027,N_1997,N_1926);
nor U2028 (N_2028,N_1918,N_1954);
nand U2029 (N_2029,N_1906,N_1920);
nand U2030 (N_2030,N_1977,N_1930);
or U2031 (N_2031,N_1995,N_1979);
or U2032 (N_2032,N_1937,N_1988);
or U2033 (N_2033,N_1940,N_1951);
and U2034 (N_2034,N_1986,N_1911);
xnor U2035 (N_2035,N_1976,N_1968);
or U2036 (N_2036,N_1971,N_1902);
and U2037 (N_2037,N_1915,N_1957);
nor U2038 (N_2038,N_1908,N_1904);
nor U2039 (N_2039,N_1967,N_1944);
or U2040 (N_2040,N_1947,N_1922);
nand U2041 (N_2041,N_1996,N_1985);
and U2042 (N_2042,N_1905,N_1925);
xnor U2043 (N_2043,N_1924,N_1942);
xnor U2044 (N_2044,N_1980,N_1929);
nor U2045 (N_2045,N_1982,N_1994);
nor U2046 (N_2046,N_1983,N_1975);
nor U2047 (N_2047,N_1972,N_1961);
nand U2048 (N_2048,N_1943,N_1963);
and U2049 (N_2049,N_1958,N_1987);
or U2050 (N_2050,N_1917,N_1922);
xor U2051 (N_2051,N_1941,N_1927);
nand U2052 (N_2052,N_1920,N_1925);
and U2053 (N_2053,N_1989,N_1924);
xor U2054 (N_2054,N_1911,N_1938);
and U2055 (N_2055,N_1904,N_1979);
and U2056 (N_2056,N_1926,N_1902);
or U2057 (N_2057,N_1918,N_1915);
nand U2058 (N_2058,N_1957,N_1981);
xnor U2059 (N_2059,N_1972,N_1988);
nor U2060 (N_2060,N_1907,N_1943);
xnor U2061 (N_2061,N_1992,N_1977);
nor U2062 (N_2062,N_1944,N_1997);
xnor U2063 (N_2063,N_1900,N_1943);
nor U2064 (N_2064,N_1988,N_1932);
or U2065 (N_2065,N_1957,N_1928);
and U2066 (N_2066,N_1948,N_1961);
xor U2067 (N_2067,N_1907,N_1950);
and U2068 (N_2068,N_1937,N_1933);
or U2069 (N_2069,N_1981,N_1918);
and U2070 (N_2070,N_1926,N_1962);
or U2071 (N_2071,N_1930,N_1910);
and U2072 (N_2072,N_1986,N_1948);
or U2073 (N_2073,N_1946,N_1908);
or U2074 (N_2074,N_1983,N_1962);
nor U2075 (N_2075,N_1929,N_1997);
nand U2076 (N_2076,N_1904,N_1941);
or U2077 (N_2077,N_1951,N_1945);
and U2078 (N_2078,N_1955,N_1970);
and U2079 (N_2079,N_1949,N_1920);
nor U2080 (N_2080,N_1923,N_1974);
xnor U2081 (N_2081,N_1932,N_1938);
xnor U2082 (N_2082,N_1991,N_1999);
or U2083 (N_2083,N_1989,N_1957);
nor U2084 (N_2084,N_1956,N_1982);
or U2085 (N_2085,N_1953,N_1961);
or U2086 (N_2086,N_1902,N_1938);
xnor U2087 (N_2087,N_1990,N_1950);
or U2088 (N_2088,N_1927,N_1937);
or U2089 (N_2089,N_1986,N_1964);
nand U2090 (N_2090,N_1920,N_1928);
and U2091 (N_2091,N_1972,N_1968);
nand U2092 (N_2092,N_1973,N_1950);
nor U2093 (N_2093,N_1959,N_1914);
and U2094 (N_2094,N_1959,N_1938);
nor U2095 (N_2095,N_1990,N_1902);
or U2096 (N_2096,N_1940,N_1934);
and U2097 (N_2097,N_1927,N_1981);
nand U2098 (N_2098,N_1993,N_1946);
nor U2099 (N_2099,N_1989,N_1935);
nor U2100 (N_2100,N_2017,N_2003);
and U2101 (N_2101,N_2038,N_2021);
nor U2102 (N_2102,N_2073,N_2095);
xor U2103 (N_2103,N_2001,N_2019);
or U2104 (N_2104,N_2006,N_2045);
nor U2105 (N_2105,N_2035,N_2094);
and U2106 (N_2106,N_2032,N_2076);
xnor U2107 (N_2107,N_2058,N_2025);
nand U2108 (N_2108,N_2015,N_2037);
and U2109 (N_2109,N_2084,N_2007);
nor U2110 (N_2110,N_2053,N_2010);
or U2111 (N_2111,N_2041,N_2078);
nand U2112 (N_2112,N_2044,N_2068);
and U2113 (N_2113,N_2008,N_2013);
nor U2114 (N_2114,N_2054,N_2065);
xnor U2115 (N_2115,N_2067,N_2034);
nor U2116 (N_2116,N_2082,N_2014);
nor U2117 (N_2117,N_2050,N_2009);
nand U2118 (N_2118,N_2097,N_2030);
xnor U2119 (N_2119,N_2048,N_2075);
nor U2120 (N_2120,N_2047,N_2004);
or U2121 (N_2121,N_2051,N_2022);
xor U2122 (N_2122,N_2033,N_2093);
nor U2123 (N_2123,N_2043,N_2063);
and U2124 (N_2124,N_2092,N_2029);
nand U2125 (N_2125,N_2057,N_2064);
xnor U2126 (N_2126,N_2060,N_2039);
and U2127 (N_2127,N_2049,N_2020);
xnor U2128 (N_2128,N_2083,N_2072);
nand U2129 (N_2129,N_2069,N_2012);
nor U2130 (N_2130,N_2089,N_2096);
and U2131 (N_2131,N_2016,N_2088);
nor U2132 (N_2132,N_2052,N_2055);
xnor U2133 (N_2133,N_2046,N_2024);
nor U2134 (N_2134,N_2066,N_2087);
nand U2135 (N_2135,N_2098,N_2042);
and U2136 (N_2136,N_2026,N_2040);
nand U2137 (N_2137,N_2027,N_2085);
nor U2138 (N_2138,N_2028,N_2086);
or U2139 (N_2139,N_2036,N_2071);
or U2140 (N_2140,N_2002,N_2059);
or U2141 (N_2141,N_2079,N_2090);
xor U2142 (N_2142,N_2018,N_2074);
xor U2143 (N_2143,N_2062,N_2099);
xor U2144 (N_2144,N_2080,N_2000);
xor U2145 (N_2145,N_2023,N_2091);
nor U2146 (N_2146,N_2056,N_2077);
nor U2147 (N_2147,N_2081,N_2070);
or U2148 (N_2148,N_2061,N_2031);
or U2149 (N_2149,N_2005,N_2011);
and U2150 (N_2150,N_2085,N_2030);
nor U2151 (N_2151,N_2098,N_2084);
or U2152 (N_2152,N_2084,N_2070);
or U2153 (N_2153,N_2020,N_2075);
nor U2154 (N_2154,N_2050,N_2033);
nand U2155 (N_2155,N_2023,N_2096);
and U2156 (N_2156,N_2055,N_2081);
xnor U2157 (N_2157,N_2008,N_2090);
xor U2158 (N_2158,N_2014,N_2086);
nand U2159 (N_2159,N_2048,N_2083);
xnor U2160 (N_2160,N_2083,N_2059);
xor U2161 (N_2161,N_2086,N_2083);
xor U2162 (N_2162,N_2008,N_2066);
nand U2163 (N_2163,N_2089,N_2021);
nor U2164 (N_2164,N_2086,N_2034);
nor U2165 (N_2165,N_2077,N_2012);
xnor U2166 (N_2166,N_2015,N_2042);
nand U2167 (N_2167,N_2087,N_2031);
or U2168 (N_2168,N_2073,N_2081);
and U2169 (N_2169,N_2082,N_2028);
and U2170 (N_2170,N_2030,N_2015);
and U2171 (N_2171,N_2042,N_2051);
or U2172 (N_2172,N_2059,N_2053);
nand U2173 (N_2173,N_2030,N_2009);
nor U2174 (N_2174,N_2060,N_2041);
or U2175 (N_2175,N_2045,N_2055);
or U2176 (N_2176,N_2047,N_2056);
nor U2177 (N_2177,N_2047,N_2009);
nand U2178 (N_2178,N_2007,N_2009);
xnor U2179 (N_2179,N_2014,N_2075);
or U2180 (N_2180,N_2043,N_2013);
xnor U2181 (N_2181,N_2073,N_2019);
nand U2182 (N_2182,N_2095,N_2013);
xor U2183 (N_2183,N_2005,N_2040);
or U2184 (N_2184,N_2091,N_2063);
and U2185 (N_2185,N_2007,N_2048);
xor U2186 (N_2186,N_2047,N_2057);
and U2187 (N_2187,N_2060,N_2025);
nand U2188 (N_2188,N_2038,N_2076);
and U2189 (N_2189,N_2027,N_2017);
nand U2190 (N_2190,N_2037,N_2099);
nor U2191 (N_2191,N_2080,N_2091);
xnor U2192 (N_2192,N_2024,N_2015);
nand U2193 (N_2193,N_2013,N_2087);
or U2194 (N_2194,N_2007,N_2013);
and U2195 (N_2195,N_2018,N_2040);
and U2196 (N_2196,N_2007,N_2060);
xnor U2197 (N_2197,N_2099,N_2055);
or U2198 (N_2198,N_2011,N_2039);
or U2199 (N_2199,N_2074,N_2082);
or U2200 (N_2200,N_2198,N_2162);
or U2201 (N_2201,N_2176,N_2152);
or U2202 (N_2202,N_2191,N_2135);
nor U2203 (N_2203,N_2128,N_2193);
or U2204 (N_2204,N_2169,N_2101);
nand U2205 (N_2205,N_2156,N_2130);
xor U2206 (N_2206,N_2104,N_2113);
and U2207 (N_2207,N_2129,N_2139);
xnor U2208 (N_2208,N_2151,N_2107);
nor U2209 (N_2209,N_2190,N_2106);
nand U2210 (N_2210,N_2102,N_2100);
xor U2211 (N_2211,N_2111,N_2144);
and U2212 (N_2212,N_2172,N_2182);
and U2213 (N_2213,N_2167,N_2196);
xor U2214 (N_2214,N_2122,N_2148);
or U2215 (N_2215,N_2114,N_2147);
or U2216 (N_2216,N_2165,N_2133);
or U2217 (N_2217,N_2124,N_2159);
or U2218 (N_2218,N_2185,N_2142);
nor U2219 (N_2219,N_2189,N_2163);
xor U2220 (N_2220,N_2150,N_2140);
xnor U2221 (N_2221,N_2117,N_2125);
nor U2222 (N_2222,N_2187,N_2105);
or U2223 (N_2223,N_2166,N_2146);
nor U2224 (N_2224,N_2134,N_2184);
nand U2225 (N_2225,N_2116,N_2160);
xor U2226 (N_2226,N_2158,N_2194);
or U2227 (N_2227,N_2175,N_2181);
nand U2228 (N_2228,N_2118,N_2127);
nor U2229 (N_2229,N_2164,N_2110);
or U2230 (N_2230,N_2115,N_2177);
and U2231 (N_2231,N_2137,N_2141);
nor U2232 (N_2232,N_2157,N_2171);
xor U2233 (N_2233,N_2136,N_2186);
xnor U2234 (N_2234,N_2108,N_2183);
or U2235 (N_2235,N_2112,N_2199);
nand U2236 (N_2236,N_2178,N_2131);
nand U2237 (N_2237,N_2119,N_2123);
nor U2238 (N_2238,N_2170,N_2143);
and U2239 (N_2239,N_2155,N_2132);
and U2240 (N_2240,N_2154,N_2121);
or U2241 (N_2241,N_2168,N_2188);
and U2242 (N_2242,N_2109,N_2103);
nand U2243 (N_2243,N_2195,N_2138);
or U2244 (N_2244,N_2145,N_2161);
nand U2245 (N_2245,N_2173,N_2153);
nor U2246 (N_2246,N_2126,N_2149);
and U2247 (N_2247,N_2180,N_2120);
and U2248 (N_2248,N_2179,N_2197);
and U2249 (N_2249,N_2192,N_2174);
and U2250 (N_2250,N_2160,N_2182);
xor U2251 (N_2251,N_2168,N_2103);
and U2252 (N_2252,N_2174,N_2134);
nor U2253 (N_2253,N_2146,N_2177);
nor U2254 (N_2254,N_2101,N_2115);
and U2255 (N_2255,N_2190,N_2124);
nand U2256 (N_2256,N_2190,N_2158);
nor U2257 (N_2257,N_2112,N_2197);
nand U2258 (N_2258,N_2149,N_2128);
or U2259 (N_2259,N_2155,N_2140);
xor U2260 (N_2260,N_2137,N_2145);
nor U2261 (N_2261,N_2197,N_2126);
nor U2262 (N_2262,N_2127,N_2186);
and U2263 (N_2263,N_2120,N_2188);
or U2264 (N_2264,N_2106,N_2132);
nand U2265 (N_2265,N_2196,N_2190);
and U2266 (N_2266,N_2181,N_2153);
and U2267 (N_2267,N_2182,N_2181);
or U2268 (N_2268,N_2182,N_2157);
nor U2269 (N_2269,N_2159,N_2131);
nor U2270 (N_2270,N_2101,N_2111);
xnor U2271 (N_2271,N_2135,N_2182);
nor U2272 (N_2272,N_2157,N_2183);
or U2273 (N_2273,N_2146,N_2162);
nand U2274 (N_2274,N_2183,N_2198);
or U2275 (N_2275,N_2144,N_2134);
or U2276 (N_2276,N_2154,N_2192);
xnor U2277 (N_2277,N_2161,N_2134);
and U2278 (N_2278,N_2184,N_2137);
nor U2279 (N_2279,N_2152,N_2110);
nand U2280 (N_2280,N_2129,N_2150);
nor U2281 (N_2281,N_2100,N_2174);
xnor U2282 (N_2282,N_2136,N_2160);
and U2283 (N_2283,N_2115,N_2171);
nor U2284 (N_2284,N_2167,N_2163);
xnor U2285 (N_2285,N_2128,N_2135);
and U2286 (N_2286,N_2105,N_2190);
or U2287 (N_2287,N_2108,N_2115);
and U2288 (N_2288,N_2119,N_2106);
nor U2289 (N_2289,N_2175,N_2193);
nor U2290 (N_2290,N_2162,N_2144);
xnor U2291 (N_2291,N_2114,N_2117);
or U2292 (N_2292,N_2116,N_2139);
and U2293 (N_2293,N_2142,N_2182);
xnor U2294 (N_2294,N_2118,N_2165);
and U2295 (N_2295,N_2198,N_2144);
and U2296 (N_2296,N_2113,N_2196);
nor U2297 (N_2297,N_2131,N_2101);
xor U2298 (N_2298,N_2172,N_2171);
or U2299 (N_2299,N_2116,N_2119);
nand U2300 (N_2300,N_2247,N_2275);
and U2301 (N_2301,N_2298,N_2276);
or U2302 (N_2302,N_2244,N_2237);
nor U2303 (N_2303,N_2289,N_2207);
nand U2304 (N_2304,N_2267,N_2297);
and U2305 (N_2305,N_2215,N_2211);
and U2306 (N_2306,N_2245,N_2280);
or U2307 (N_2307,N_2220,N_2252);
nand U2308 (N_2308,N_2206,N_2233);
nor U2309 (N_2309,N_2200,N_2223);
nand U2310 (N_2310,N_2264,N_2270);
xnor U2311 (N_2311,N_2261,N_2269);
or U2312 (N_2312,N_2281,N_2242);
nand U2313 (N_2313,N_2285,N_2240);
nand U2314 (N_2314,N_2271,N_2294);
nand U2315 (N_2315,N_2212,N_2255);
nand U2316 (N_2316,N_2236,N_2235);
and U2317 (N_2317,N_2202,N_2287);
nor U2318 (N_2318,N_2262,N_2263);
or U2319 (N_2319,N_2249,N_2248);
nand U2320 (N_2320,N_2213,N_2225);
nand U2321 (N_2321,N_2268,N_2241);
nand U2322 (N_2322,N_2238,N_2210);
or U2323 (N_2323,N_2282,N_2288);
or U2324 (N_2324,N_2293,N_2227);
nand U2325 (N_2325,N_2222,N_2291);
xor U2326 (N_2326,N_2219,N_2274);
xor U2327 (N_2327,N_2205,N_2278);
nand U2328 (N_2328,N_2272,N_2279);
nor U2329 (N_2329,N_2203,N_2226);
xor U2330 (N_2330,N_2254,N_2228);
nand U2331 (N_2331,N_2292,N_2218);
nand U2332 (N_2332,N_2284,N_2253);
nor U2333 (N_2333,N_2221,N_2259);
nor U2334 (N_2334,N_2296,N_2273);
or U2335 (N_2335,N_2231,N_2201);
and U2336 (N_2336,N_2290,N_2266);
nand U2337 (N_2337,N_2229,N_2230);
nand U2338 (N_2338,N_2250,N_2265);
nor U2339 (N_2339,N_2295,N_2216);
or U2340 (N_2340,N_2239,N_2257);
or U2341 (N_2341,N_2299,N_2251);
nor U2342 (N_2342,N_2232,N_2258);
xnor U2343 (N_2343,N_2243,N_2277);
xnor U2344 (N_2344,N_2286,N_2224);
or U2345 (N_2345,N_2283,N_2234);
nor U2346 (N_2346,N_2217,N_2209);
nand U2347 (N_2347,N_2246,N_2214);
xor U2348 (N_2348,N_2208,N_2256);
xor U2349 (N_2349,N_2260,N_2204);
and U2350 (N_2350,N_2268,N_2229);
nor U2351 (N_2351,N_2268,N_2223);
nand U2352 (N_2352,N_2238,N_2219);
nand U2353 (N_2353,N_2207,N_2263);
nor U2354 (N_2354,N_2216,N_2213);
nand U2355 (N_2355,N_2274,N_2273);
xor U2356 (N_2356,N_2252,N_2299);
nor U2357 (N_2357,N_2201,N_2227);
xnor U2358 (N_2358,N_2250,N_2251);
xor U2359 (N_2359,N_2202,N_2276);
nor U2360 (N_2360,N_2240,N_2256);
xnor U2361 (N_2361,N_2209,N_2279);
or U2362 (N_2362,N_2233,N_2294);
nand U2363 (N_2363,N_2282,N_2250);
nor U2364 (N_2364,N_2236,N_2209);
xnor U2365 (N_2365,N_2259,N_2231);
or U2366 (N_2366,N_2218,N_2250);
and U2367 (N_2367,N_2237,N_2226);
or U2368 (N_2368,N_2271,N_2200);
or U2369 (N_2369,N_2238,N_2243);
xnor U2370 (N_2370,N_2272,N_2277);
nor U2371 (N_2371,N_2246,N_2273);
xor U2372 (N_2372,N_2271,N_2209);
and U2373 (N_2373,N_2251,N_2229);
nor U2374 (N_2374,N_2261,N_2296);
or U2375 (N_2375,N_2210,N_2227);
and U2376 (N_2376,N_2224,N_2252);
and U2377 (N_2377,N_2271,N_2220);
nand U2378 (N_2378,N_2265,N_2216);
or U2379 (N_2379,N_2287,N_2216);
or U2380 (N_2380,N_2229,N_2235);
nor U2381 (N_2381,N_2298,N_2236);
xor U2382 (N_2382,N_2293,N_2203);
or U2383 (N_2383,N_2222,N_2221);
or U2384 (N_2384,N_2256,N_2224);
and U2385 (N_2385,N_2212,N_2249);
nand U2386 (N_2386,N_2294,N_2265);
and U2387 (N_2387,N_2231,N_2202);
or U2388 (N_2388,N_2240,N_2274);
or U2389 (N_2389,N_2214,N_2201);
xnor U2390 (N_2390,N_2239,N_2284);
nand U2391 (N_2391,N_2230,N_2245);
nand U2392 (N_2392,N_2273,N_2278);
nor U2393 (N_2393,N_2267,N_2238);
nor U2394 (N_2394,N_2264,N_2262);
nor U2395 (N_2395,N_2287,N_2225);
xnor U2396 (N_2396,N_2290,N_2282);
nor U2397 (N_2397,N_2282,N_2200);
nor U2398 (N_2398,N_2222,N_2270);
nor U2399 (N_2399,N_2203,N_2227);
nor U2400 (N_2400,N_2367,N_2397);
nor U2401 (N_2401,N_2311,N_2336);
nor U2402 (N_2402,N_2322,N_2350);
nor U2403 (N_2403,N_2357,N_2347);
or U2404 (N_2404,N_2305,N_2321);
nand U2405 (N_2405,N_2372,N_2351);
or U2406 (N_2406,N_2308,N_2395);
xnor U2407 (N_2407,N_2394,N_2314);
xnor U2408 (N_2408,N_2319,N_2380);
nor U2409 (N_2409,N_2385,N_2370);
nor U2410 (N_2410,N_2300,N_2381);
nand U2411 (N_2411,N_2360,N_2362);
nand U2412 (N_2412,N_2396,N_2334);
nand U2413 (N_2413,N_2304,N_2373);
or U2414 (N_2414,N_2375,N_2337);
or U2415 (N_2415,N_2368,N_2361);
nor U2416 (N_2416,N_2331,N_2376);
and U2417 (N_2417,N_2389,N_2384);
xnor U2418 (N_2418,N_2341,N_2315);
or U2419 (N_2419,N_2393,N_2313);
nand U2420 (N_2420,N_2316,N_2326);
or U2421 (N_2421,N_2323,N_2330);
nor U2422 (N_2422,N_2382,N_2354);
or U2423 (N_2423,N_2369,N_2349);
and U2424 (N_2424,N_2383,N_2379);
nor U2425 (N_2425,N_2339,N_2371);
nand U2426 (N_2426,N_2327,N_2387);
nand U2427 (N_2427,N_2309,N_2333);
nor U2428 (N_2428,N_2364,N_2352);
nor U2429 (N_2429,N_2358,N_2365);
xnor U2430 (N_2430,N_2391,N_2399);
and U2431 (N_2431,N_2324,N_2335);
nor U2432 (N_2432,N_2328,N_2318);
nor U2433 (N_2433,N_2338,N_2345);
xnor U2434 (N_2434,N_2359,N_2344);
or U2435 (N_2435,N_2342,N_2307);
nor U2436 (N_2436,N_2348,N_2325);
nor U2437 (N_2437,N_2329,N_2343);
nor U2438 (N_2438,N_2392,N_2356);
or U2439 (N_2439,N_2303,N_2388);
and U2440 (N_2440,N_2377,N_2390);
xnor U2441 (N_2441,N_2374,N_2366);
nor U2442 (N_2442,N_2306,N_2301);
and U2443 (N_2443,N_2332,N_2386);
nand U2444 (N_2444,N_2302,N_2312);
or U2445 (N_2445,N_2363,N_2340);
nor U2446 (N_2446,N_2355,N_2398);
or U2447 (N_2447,N_2310,N_2320);
and U2448 (N_2448,N_2353,N_2378);
and U2449 (N_2449,N_2317,N_2346);
nor U2450 (N_2450,N_2346,N_2373);
nor U2451 (N_2451,N_2365,N_2319);
nor U2452 (N_2452,N_2395,N_2321);
nor U2453 (N_2453,N_2320,N_2334);
and U2454 (N_2454,N_2342,N_2360);
or U2455 (N_2455,N_2390,N_2310);
nor U2456 (N_2456,N_2328,N_2325);
xnor U2457 (N_2457,N_2347,N_2380);
and U2458 (N_2458,N_2313,N_2314);
nand U2459 (N_2459,N_2321,N_2353);
nand U2460 (N_2460,N_2367,N_2390);
and U2461 (N_2461,N_2304,N_2346);
xor U2462 (N_2462,N_2346,N_2384);
xnor U2463 (N_2463,N_2355,N_2380);
nor U2464 (N_2464,N_2371,N_2332);
nor U2465 (N_2465,N_2308,N_2384);
nand U2466 (N_2466,N_2309,N_2328);
and U2467 (N_2467,N_2329,N_2313);
or U2468 (N_2468,N_2384,N_2366);
xor U2469 (N_2469,N_2355,N_2324);
nor U2470 (N_2470,N_2335,N_2363);
nor U2471 (N_2471,N_2365,N_2305);
nand U2472 (N_2472,N_2389,N_2387);
or U2473 (N_2473,N_2303,N_2345);
xor U2474 (N_2474,N_2305,N_2361);
nor U2475 (N_2475,N_2345,N_2346);
xnor U2476 (N_2476,N_2304,N_2329);
nand U2477 (N_2477,N_2393,N_2326);
nor U2478 (N_2478,N_2318,N_2333);
nor U2479 (N_2479,N_2310,N_2374);
nor U2480 (N_2480,N_2358,N_2337);
xor U2481 (N_2481,N_2388,N_2350);
xnor U2482 (N_2482,N_2390,N_2378);
nand U2483 (N_2483,N_2349,N_2361);
nor U2484 (N_2484,N_2378,N_2341);
xor U2485 (N_2485,N_2380,N_2307);
nor U2486 (N_2486,N_2307,N_2323);
and U2487 (N_2487,N_2368,N_2345);
and U2488 (N_2488,N_2391,N_2397);
nand U2489 (N_2489,N_2369,N_2314);
or U2490 (N_2490,N_2351,N_2305);
xnor U2491 (N_2491,N_2378,N_2309);
xor U2492 (N_2492,N_2360,N_2311);
xnor U2493 (N_2493,N_2358,N_2319);
and U2494 (N_2494,N_2370,N_2327);
xnor U2495 (N_2495,N_2325,N_2305);
and U2496 (N_2496,N_2342,N_2341);
and U2497 (N_2497,N_2373,N_2359);
xor U2498 (N_2498,N_2307,N_2339);
and U2499 (N_2499,N_2370,N_2376);
nand U2500 (N_2500,N_2452,N_2415);
xnor U2501 (N_2501,N_2467,N_2401);
nor U2502 (N_2502,N_2476,N_2498);
nand U2503 (N_2503,N_2497,N_2453);
nand U2504 (N_2504,N_2470,N_2492);
and U2505 (N_2505,N_2449,N_2432);
nor U2506 (N_2506,N_2488,N_2422);
nor U2507 (N_2507,N_2462,N_2487);
or U2508 (N_2508,N_2473,N_2483);
nand U2509 (N_2509,N_2440,N_2479);
xnor U2510 (N_2510,N_2493,N_2495);
or U2511 (N_2511,N_2446,N_2441);
and U2512 (N_2512,N_2408,N_2466);
xnor U2513 (N_2513,N_2485,N_2405);
nor U2514 (N_2514,N_2463,N_2416);
nor U2515 (N_2515,N_2469,N_2414);
or U2516 (N_2516,N_2434,N_2437);
nor U2517 (N_2517,N_2481,N_2443);
xor U2518 (N_2518,N_2410,N_2471);
nor U2519 (N_2519,N_2409,N_2477);
xnor U2520 (N_2520,N_2427,N_2404);
nand U2521 (N_2521,N_2426,N_2419);
nor U2522 (N_2522,N_2459,N_2475);
nor U2523 (N_2523,N_2445,N_2447);
xor U2524 (N_2524,N_2420,N_2455);
and U2525 (N_2525,N_2430,N_2450);
nand U2526 (N_2526,N_2451,N_2407);
xor U2527 (N_2527,N_2491,N_2474);
nand U2528 (N_2528,N_2486,N_2482);
nand U2529 (N_2529,N_2480,N_2442);
xnor U2530 (N_2530,N_2428,N_2444);
or U2531 (N_2531,N_2435,N_2423);
or U2532 (N_2532,N_2496,N_2448);
nand U2533 (N_2533,N_2402,N_2457);
nand U2534 (N_2534,N_2490,N_2439);
xnor U2535 (N_2535,N_2468,N_2484);
and U2536 (N_2536,N_2417,N_2489);
and U2537 (N_2537,N_2431,N_2460);
xor U2538 (N_2538,N_2425,N_2421);
xnor U2539 (N_2539,N_2429,N_2438);
or U2540 (N_2540,N_2403,N_2465);
nand U2541 (N_2541,N_2433,N_2494);
nor U2542 (N_2542,N_2458,N_2454);
or U2543 (N_2543,N_2400,N_2461);
nand U2544 (N_2544,N_2413,N_2478);
nand U2545 (N_2545,N_2472,N_2412);
nand U2546 (N_2546,N_2424,N_2411);
nor U2547 (N_2547,N_2436,N_2464);
nand U2548 (N_2548,N_2456,N_2418);
or U2549 (N_2549,N_2406,N_2499);
nand U2550 (N_2550,N_2451,N_2472);
nor U2551 (N_2551,N_2498,N_2496);
and U2552 (N_2552,N_2470,N_2460);
xor U2553 (N_2553,N_2490,N_2487);
nand U2554 (N_2554,N_2413,N_2498);
nand U2555 (N_2555,N_2495,N_2475);
nand U2556 (N_2556,N_2492,N_2404);
or U2557 (N_2557,N_2407,N_2494);
or U2558 (N_2558,N_2426,N_2469);
nand U2559 (N_2559,N_2415,N_2474);
nor U2560 (N_2560,N_2432,N_2403);
nand U2561 (N_2561,N_2495,N_2482);
nand U2562 (N_2562,N_2411,N_2405);
or U2563 (N_2563,N_2485,N_2426);
or U2564 (N_2564,N_2434,N_2423);
nor U2565 (N_2565,N_2458,N_2439);
nor U2566 (N_2566,N_2418,N_2446);
or U2567 (N_2567,N_2494,N_2498);
or U2568 (N_2568,N_2419,N_2463);
xnor U2569 (N_2569,N_2490,N_2451);
nand U2570 (N_2570,N_2414,N_2488);
and U2571 (N_2571,N_2498,N_2495);
or U2572 (N_2572,N_2420,N_2470);
nand U2573 (N_2573,N_2441,N_2431);
nor U2574 (N_2574,N_2492,N_2447);
or U2575 (N_2575,N_2414,N_2439);
nor U2576 (N_2576,N_2438,N_2490);
xnor U2577 (N_2577,N_2479,N_2408);
nand U2578 (N_2578,N_2449,N_2493);
xnor U2579 (N_2579,N_2477,N_2432);
nor U2580 (N_2580,N_2418,N_2496);
nor U2581 (N_2581,N_2444,N_2482);
xor U2582 (N_2582,N_2493,N_2480);
or U2583 (N_2583,N_2404,N_2441);
or U2584 (N_2584,N_2419,N_2459);
and U2585 (N_2585,N_2461,N_2464);
xor U2586 (N_2586,N_2489,N_2414);
nand U2587 (N_2587,N_2418,N_2400);
nor U2588 (N_2588,N_2400,N_2408);
xnor U2589 (N_2589,N_2416,N_2407);
nand U2590 (N_2590,N_2467,N_2406);
nand U2591 (N_2591,N_2422,N_2435);
and U2592 (N_2592,N_2472,N_2484);
xor U2593 (N_2593,N_2418,N_2489);
or U2594 (N_2594,N_2477,N_2474);
nand U2595 (N_2595,N_2457,N_2479);
and U2596 (N_2596,N_2402,N_2401);
and U2597 (N_2597,N_2452,N_2446);
or U2598 (N_2598,N_2452,N_2435);
nor U2599 (N_2599,N_2413,N_2440);
and U2600 (N_2600,N_2577,N_2588);
and U2601 (N_2601,N_2567,N_2543);
nor U2602 (N_2602,N_2598,N_2520);
nor U2603 (N_2603,N_2532,N_2591);
or U2604 (N_2604,N_2575,N_2514);
nor U2605 (N_2605,N_2590,N_2549);
nor U2606 (N_2606,N_2576,N_2522);
nand U2607 (N_2607,N_2587,N_2551);
nor U2608 (N_2608,N_2533,N_2572);
or U2609 (N_2609,N_2510,N_2560);
nor U2610 (N_2610,N_2504,N_2595);
and U2611 (N_2611,N_2557,N_2519);
nand U2612 (N_2612,N_2583,N_2553);
xnor U2613 (N_2613,N_2585,N_2597);
or U2614 (N_2614,N_2568,N_2539);
and U2615 (N_2615,N_2593,N_2582);
nor U2616 (N_2616,N_2545,N_2562);
and U2617 (N_2617,N_2594,N_2511);
nand U2618 (N_2618,N_2547,N_2515);
nand U2619 (N_2619,N_2584,N_2507);
xnor U2620 (N_2620,N_2592,N_2552);
or U2621 (N_2621,N_2525,N_2580);
nor U2622 (N_2622,N_2527,N_2581);
and U2623 (N_2623,N_2596,N_2586);
xor U2624 (N_2624,N_2500,N_2550);
nor U2625 (N_2625,N_2502,N_2546);
nand U2626 (N_2626,N_2505,N_2574);
nand U2627 (N_2627,N_2554,N_2521);
or U2628 (N_2628,N_2555,N_2542);
or U2629 (N_2629,N_2516,N_2573);
or U2630 (N_2630,N_2501,N_2536);
xnor U2631 (N_2631,N_2548,N_2517);
nand U2632 (N_2632,N_2509,N_2503);
and U2633 (N_2633,N_2579,N_2558);
xnor U2634 (N_2634,N_2563,N_2569);
xnor U2635 (N_2635,N_2566,N_2518);
nand U2636 (N_2636,N_2599,N_2508);
or U2637 (N_2637,N_2534,N_2513);
and U2638 (N_2638,N_2556,N_2565);
or U2639 (N_2639,N_2528,N_2535);
xnor U2640 (N_2640,N_2541,N_2523);
nand U2641 (N_2641,N_2561,N_2544);
and U2642 (N_2642,N_2538,N_2524);
and U2643 (N_2643,N_2529,N_2589);
or U2644 (N_2644,N_2540,N_2571);
nand U2645 (N_2645,N_2559,N_2506);
xor U2646 (N_2646,N_2526,N_2570);
and U2647 (N_2647,N_2512,N_2564);
xor U2648 (N_2648,N_2530,N_2578);
or U2649 (N_2649,N_2537,N_2531);
and U2650 (N_2650,N_2560,N_2526);
and U2651 (N_2651,N_2538,N_2575);
or U2652 (N_2652,N_2509,N_2557);
nor U2653 (N_2653,N_2552,N_2515);
xor U2654 (N_2654,N_2557,N_2548);
xor U2655 (N_2655,N_2568,N_2500);
nor U2656 (N_2656,N_2596,N_2589);
nor U2657 (N_2657,N_2517,N_2599);
nor U2658 (N_2658,N_2579,N_2516);
nor U2659 (N_2659,N_2595,N_2537);
nand U2660 (N_2660,N_2515,N_2583);
nand U2661 (N_2661,N_2514,N_2500);
and U2662 (N_2662,N_2542,N_2510);
xor U2663 (N_2663,N_2588,N_2530);
nor U2664 (N_2664,N_2519,N_2552);
or U2665 (N_2665,N_2520,N_2594);
or U2666 (N_2666,N_2574,N_2501);
or U2667 (N_2667,N_2574,N_2555);
xnor U2668 (N_2668,N_2548,N_2579);
and U2669 (N_2669,N_2598,N_2548);
nand U2670 (N_2670,N_2542,N_2504);
xor U2671 (N_2671,N_2518,N_2538);
nor U2672 (N_2672,N_2508,N_2522);
or U2673 (N_2673,N_2591,N_2575);
and U2674 (N_2674,N_2550,N_2567);
or U2675 (N_2675,N_2574,N_2541);
and U2676 (N_2676,N_2561,N_2520);
and U2677 (N_2677,N_2579,N_2502);
or U2678 (N_2678,N_2552,N_2559);
xnor U2679 (N_2679,N_2559,N_2576);
nor U2680 (N_2680,N_2578,N_2563);
nand U2681 (N_2681,N_2555,N_2528);
nor U2682 (N_2682,N_2586,N_2530);
nand U2683 (N_2683,N_2519,N_2500);
nor U2684 (N_2684,N_2586,N_2503);
nand U2685 (N_2685,N_2564,N_2521);
or U2686 (N_2686,N_2507,N_2556);
nor U2687 (N_2687,N_2549,N_2535);
nor U2688 (N_2688,N_2560,N_2581);
xor U2689 (N_2689,N_2536,N_2509);
xor U2690 (N_2690,N_2519,N_2504);
xnor U2691 (N_2691,N_2581,N_2543);
and U2692 (N_2692,N_2598,N_2596);
and U2693 (N_2693,N_2521,N_2557);
or U2694 (N_2694,N_2566,N_2545);
and U2695 (N_2695,N_2597,N_2533);
and U2696 (N_2696,N_2580,N_2592);
nor U2697 (N_2697,N_2515,N_2592);
nor U2698 (N_2698,N_2592,N_2559);
nand U2699 (N_2699,N_2595,N_2563);
and U2700 (N_2700,N_2656,N_2631);
nor U2701 (N_2701,N_2633,N_2647);
nand U2702 (N_2702,N_2675,N_2663);
xnor U2703 (N_2703,N_2667,N_2672);
nor U2704 (N_2704,N_2642,N_2628);
xnor U2705 (N_2705,N_2697,N_2621);
xnor U2706 (N_2706,N_2678,N_2687);
or U2707 (N_2707,N_2635,N_2625);
xor U2708 (N_2708,N_2618,N_2637);
and U2709 (N_2709,N_2649,N_2616);
xor U2710 (N_2710,N_2640,N_2692);
xnor U2711 (N_2711,N_2622,N_2614);
nor U2712 (N_2712,N_2693,N_2671);
and U2713 (N_2713,N_2645,N_2643);
or U2714 (N_2714,N_2666,N_2699);
nand U2715 (N_2715,N_2613,N_2677);
and U2716 (N_2716,N_2669,N_2655);
nand U2717 (N_2717,N_2652,N_2632);
nand U2718 (N_2718,N_2660,N_2641);
nor U2719 (N_2719,N_2696,N_2691);
xnor U2720 (N_2720,N_2685,N_2638);
nand U2721 (N_2721,N_2634,N_2679);
or U2722 (N_2722,N_2626,N_2617);
and U2723 (N_2723,N_2611,N_2636);
nand U2724 (N_2724,N_2620,N_2688);
nor U2725 (N_2725,N_2661,N_2607);
xor U2726 (N_2726,N_2686,N_2698);
or U2727 (N_2727,N_2690,N_2694);
and U2728 (N_2728,N_2608,N_2619);
or U2729 (N_2729,N_2629,N_2639);
and U2730 (N_2730,N_2606,N_2674);
and U2731 (N_2731,N_2654,N_2609);
xor U2732 (N_2732,N_2670,N_2601);
nand U2733 (N_2733,N_2683,N_2657);
nand U2734 (N_2734,N_2603,N_2653);
nand U2735 (N_2735,N_2650,N_2681);
nand U2736 (N_2736,N_2602,N_2610);
nand U2737 (N_2737,N_2624,N_2659);
xor U2738 (N_2738,N_2648,N_2673);
nand U2739 (N_2739,N_2662,N_2658);
nor U2740 (N_2740,N_2605,N_2600);
xnor U2741 (N_2741,N_2627,N_2604);
nand U2742 (N_2742,N_2689,N_2684);
xor U2743 (N_2743,N_2615,N_2665);
nand U2744 (N_2744,N_2680,N_2664);
nand U2745 (N_2745,N_2695,N_2676);
nor U2746 (N_2746,N_2651,N_2612);
nand U2747 (N_2747,N_2668,N_2623);
nand U2748 (N_2748,N_2630,N_2682);
nand U2749 (N_2749,N_2644,N_2646);
or U2750 (N_2750,N_2658,N_2692);
and U2751 (N_2751,N_2686,N_2618);
nor U2752 (N_2752,N_2665,N_2691);
and U2753 (N_2753,N_2691,N_2638);
nand U2754 (N_2754,N_2619,N_2637);
nand U2755 (N_2755,N_2605,N_2692);
and U2756 (N_2756,N_2671,N_2606);
or U2757 (N_2757,N_2643,N_2617);
and U2758 (N_2758,N_2643,N_2623);
nand U2759 (N_2759,N_2615,N_2673);
or U2760 (N_2760,N_2606,N_2604);
and U2761 (N_2761,N_2660,N_2667);
nand U2762 (N_2762,N_2623,N_2666);
or U2763 (N_2763,N_2655,N_2603);
nand U2764 (N_2764,N_2634,N_2611);
and U2765 (N_2765,N_2640,N_2636);
nand U2766 (N_2766,N_2612,N_2622);
nor U2767 (N_2767,N_2631,N_2688);
or U2768 (N_2768,N_2623,N_2678);
nor U2769 (N_2769,N_2633,N_2664);
nand U2770 (N_2770,N_2610,N_2629);
and U2771 (N_2771,N_2629,N_2699);
and U2772 (N_2772,N_2622,N_2603);
or U2773 (N_2773,N_2671,N_2660);
xor U2774 (N_2774,N_2671,N_2680);
nor U2775 (N_2775,N_2693,N_2675);
nand U2776 (N_2776,N_2606,N_2693);
nor U2777 (N_2777,N_2672,N_2600);
nor U2778 (N_2778,N_2689,N_2610);
xnor U2779 (N_2779,N_2612,N_2623);
or U2780 (N_2780,N_2629,N_2640);
nor U2781 (N_2781,N_2692,N_2637);
nand U2782 (N_2782,N_2692,N_2685);
nor U2783 (N_2783,N_2656,N_2600);
nand U2784 (N_2784,N_2691,N_2677);
nor U2785 (N_2785,N_2625,N_2615);
or U2786 (N_2786,N_2613,N_2668);
and U2787 (N_2787,N_2642,N_2641);
nor U2788 (N_2788,N_2660,N_2602);
xor U2789 (N_2789,N_2679,N_2645);
nand U2790 (N_2790,N_2668,N_2650);
xnor U2791 (N_2791,N_2663,N_2629);
or U2792 (N_2792,N_2631,N_2633);
or U2793 (N_2793,N_2626,N_2658);
nand U2794 (N_2794,N_2673,N_2623);
nand U2795 (N_2795,N_2688,N_2693);
nor U2796 (N_2796,N_2690,N_2699);
nand U2797 (N_2797,N_2618,N_2678);
and U2798 (N_2798,N_2632,N_2668);
nor U2799 (N_2799,N_2658,N_2668);
nor U2800 (N_2800,N_2702,N_2753);
nor U2801 (N_2801,N_2773,N_2717);
nand U2802 (N_2802,N_2729,N_2730);
xnor U2803 (N_2803,N_2779,N_2725);
and U2804 (N_2804,N_2793,N_2728);
xnor U2805 (N_2805,N_2708,N_2741);
or U2806 (N_2806,N_2710,N_2732);
or U2807 (N_2807,N_2727,N_2778);
and U2808 (N_2808,N_2722,N_2736);
and U2809 (N_2809,N_2724,N_2757);
and U2810 (N_2810,N_2719,N_2766);
nor U2811 (N_2811,N_2713,N_2734);
nand U2812 (N_2812,N_2743,N_2726);
or U2813 (N_2813,N_2745,N_2723);
and U2814 (N_2814,N_2700,N_2788);
xor U2815 (N_2815,N_2707,N_2709);
and U2816 (N_2816,N_2737,N_2777);
nand U2817 (N_2817,N_2767,N_2711);
xor U2818 (N_2818,N_2751,N_2762);
or U2819 (N_2819,N_2783,N_2786);
and U2820 (N_2820,N_2759,N_2798);
or U2821 (N_2821,N_2787,N_2774);
nor U2822 (N_2822,N_2763,N_2701);
and U2823 (N_2823,N_2771,N_2794);
and U2824 (N_2824,N_2780,N_2776);
xor U2825 (N_2825,N_2796,N_2733);
nand U2826 (N_2826,N_2756,N_2714);
xnor U2827 (N_2827,N_2797,N_2792);
nand U2828 (N_2828,N_2768,N_2772);
or U2829 (N_2829,N_2760,N_2748);
or U2830 (N_2830,N_2790,N_2781);
nand U2831 (N_2831,N_2782,N_2742);
nand U2832 (N_2832,N_2770,N_2716);
nand U2833 (N_2833,N_2795,N_2740);
nor U2834 (N_2834,N_2791,N_2705);
xor U2835 (N_2835,N_2744,N_2706);
nor U2836 (N_2836,N_2738,N_2749);
and U2837 (N_2837,N_2718,N_2703);
and U2838 (N_2838,N_2789,N_2715);
and U2839 (N_2839,N_2750,N_2704);
and U2840 (N_2840,N_2758,N_2735);
xor U2841 (N_2841,N_2761,N_2746);
and U2842 (N_2842,N_2720,N_2764);
and U2843 (N_2843,N_2712,N_2754);
nor U2844 (N_2844,N_2731,N_2765);
nor U2845 (N_2845,N_2784,N_2775);
xor U2846 (N_2846,N_2769,N_2799);
and U2847 (N_2847,N_2752,N_2755);
nand U2848 (N_2848,N_2739,N_2785);
xor U2849 (N_2849,N_2747,N_2721);
nor U2850 (N_2850,N_2704,N_2775);
and U2851 (N_2851,N_2746,N_2790);
nor U2852 (N_2852,N_2797,N_2720);
nand U2853 (N_2853,N_2787,N_2785);
nand U2854 (N_2854,N_2749,N_2722);
or U2855 (N_2855,N_2785,N_2743);
nand U2856 (N_2856,N_2746,N_2779);
and U2857 (N_2857,N_2785,N_2773);
or U2858 (N_2858,N_2738,N_2751);
and U2859 (N_2859,N_2708,N_2777);
and U2860 (N_2860,N_2729,N_2734);
xor U2861 (N_2861,N_2768,N_2751);
and U2862 (N_2862,N_2755,N_2795);
nand U2863 (N_2863,N_2783,N_2795);
or U2864 (N_2864,N_2728,N_2791);
xnor U2865 (N_2865,N_2796,N_2783);
nand U2866 (N_2866,N_2759,N_2707);
nand U2867 (N_2867,N_2771,N_2764);
xnor U2868 (N_2868,N_2764,N_2755);
and U2869 (N_2869,N_2739,N_2786);
and U2870 (N_2870,N_2762,N_2735);
xor U2871 (N_2871,N_2750,N_2723);
xnor U2872 (N_2872,N_2788,N_2770);
nor U2873 (N_2873,N_2782,N_2764);
and U2874 (N_2874,N_2741,N_2776);
or U2875 (N_2875,N_2703,N_2768);
and U2876 (N_2876,N_2739,N_2711);
and U2877 (N_2877,N_2796,N_2772);
and U2878 (N_2878,N_2747,N_2766);
nand U2879 (N_2879,N_2721,N_2756);
nor U2880 (N_2880,N_2761,N_2715);
and U2881 (N_2881,N_2748,N_2771);
nand U2882 (N_2882,N_2786,N_2759);
and U2883 (N_2883,N_2740,N_2768);
and U2884 (N_2884,N_2745,N_2703);
or U2885 (N_2885,N_2731,N_2730);
nor U2886 (N_2886,N_2765,N_2713);
or U2887 (N_2887,N_2799,N_2729);
or U2888 (N_2888,N_2767,N_2748);
and U2889 (N_2889,N_2719,N_2773);
nor U2890 (N_2890,N_2746,N_2702);
nand U2891 (N_2891,N_2776,N_2797);
or U2892 (N_2892,N_2703,N_2721);
nand U2893 (N_2893,N_2762,N_2725);
and U2894 (N_2894,N_2773,N_2734);
nor U2895 (N_2895,N_2753,N_2750);
or U2896 (N_2896,N_2727,N_2754);
xor U2897 (N_2897,N_2771,N_2723);
or U2898 (N_2898,N_2749,N_2770);
nand U2899 (N_2899,N_2794,N_2739);
xor U2900 (N_2900,N_2830,N_2837);
nor U2901 (N_2901,N_2885,N_2818);
nor U2902 (N_2902,N_2852,N_2888);
and U2903 (N_2903,N_2827,N_2803);
and U2904 (N_2904,N_2839,N_2821);
and U2905 (N_2905,N_2809,N_2810);
and U2906 (N_2906,N_2869,N_2893);
or U2907 (N_2907,N_2816,N_2833);
nor U2908 (N_2908,N_2842,N_2863);
nor U2909 (N_2909,N_2802,N_2819);
or U2910 (N_2910,N_2855,N_2861);
nand U2911 (N_2911,N_2811,N_2822);
xnor U2912 (N_2912,N_2808,N_2860);
xor U2913 (N_2913,N_2838,N_2899);
or U2914 (N_2914,N_2874,N_2826);
nand U2915 (N_2915,N_2825,N_2813);
or U2916 (N_2916,N_2870,N_2891);
nor U2917 (N_2917,N_2806,N_2881);
xnor U2918 (N_2918,N_2831,N_2864);
xnor U2919 (N_2919,N_2849,N_2854);
and U2920 (N_2920,N_2823,N_2848);
xnor U2921 (N_2921,N_2889,N_2865);
or U2922 (N_2922,N_2866,N_2843);
or U2923 (N_2923,N_2868,N_2812);
nand U2924 (N_2924,N_2815,N_2862);
or U2925 (N_2925,N_2850,N_2897);
nand U2926 (N_2926,N_2894,N_2895);
nor U2927 (N_2927,N_2857,N_2844);
nand U2928 (N_2928,N_2887,N_2876);
and U2929 (N_2929,N_2801,N_2820);
nand U2930 (N_2930,N_2834,N_2858);
or U2931 (N_2931,N_2832,N_2886);
or U2932 (N_2932,N_2845,N_2856);
nor U2933 (N_2933,N_2878,N_2883);
nor U2934 (N_2934,N_2884,N_2800);
nand U2935 (N_2935,N_2853,N_2877);
nand U2936 (N_2936,N_2841,N_2890);
or U2937 (N_2937,N_2828,N_2817);
and U2938 (N_2938,N_2882,N_2859);
nor U2939 (N_2939,N_2814,N_2880);
and U2940 (N_2940,N_2872,N_2824);
or U2941 (N_2941,N_2896,N_2873);
xor U2942 (N_2942,N_2846,N_2867);
nand U2943 (N_2943,N_2836,N_2835);
or U2944 (N_2944,N_2892,N_2898);
xor U2945 (N_2945,N_2829,N_2805);
nor U2946 (N_2946,N_2840,N_2871);
nor U2947 (N_2947,N_2851,N_2847);
or U2948 (N_2948,N_2879,N_2807);
nand U2949 (N_2949,N_2804,N_2875);
xor U2950 (N_2950,N_2822,N_2864);
nand U2951 (N_2951,N_2817,N_2805);
nor U2952 (N_2952,N_2816,N_2875);
and U2953 (N_2953,N_2866,N_2876);
xnor U2954 (N_2954,N_2880,N_2873);
xnor U2955 (N_2955,N_2843,N_2867);
xnor U2956 (N_2956,N_2859,N_2833);
or U2957 (N_2957,N_2847,N_2866);
and U2958 (N_2958,N_2814,N_2892);
and U2959 (N_2959,N_2834,N_2828);
nand U2960 (N_2960,N_2829,N_2870);
or U2961 (N_2961,N_2882,N_2833);
xor U2962 (N_2962,N_2876,N_2815);
or U2963 (N_2963,N_2863,N_2840);
xor U2964 (N_2964,N_2899,N_2802);
xnor U2965 (N_2965,N_2878,N_2831);
xnor U2966 (N_2966,N_2847,N_2819);
and U2967 (N_2967,N_2807,N_2898);
xor U2968 (N_2968,N_2895,N_2802);
nand U2969 (N_2969,N_2878,N_2876);
xnor U2970 (N_2970,N_2844,N_2843);
and U2971 (N_2971,N_2813,N_2817);
and U2972 (N_2972,N_2870,N_2855);
xnor U2973 (N_2973,N_2885,N_2867);
and U2974 (N_2974,N_2884,N_2805);
or U2975 (N_2975,N_2833,N_2854);
nor U2976 (N_2976,N_2852,N_2883);
or U2977 (N_2977,N_2838,N_2852);
or U2978 (N_2978,N_2897,N_2894);
or U2979 (N_2979,N_2843,N_2810);
or U2980 (N_2980,N_2834,N_2823);
nand U2981 (N_2981,N_2872,N_2875);
and U2982 (N_2982,N_2852,N_2895);
nor U2983 (N_2983,N_2874,N_2841);
or U2984 (N_2984,N_2898,N_2857);
nor U2985 (N_2985,N_2818,N_2884);
xor U2986 (N_2986,N_2891,N_2831);
or U2987 (N_2987,N_2891,N_2823);
or U2988 (N_2988,N_2813,N_2808);
and U2989 (N_2989,N_2894,N_2842);
nor U2990 (N_2990,N_2856,N_2876);
and U2991 (N_2991,N_2874,N_2846);
and U2992 (N_2992,N_2807,N_2858);
or U2993 (N_2993,N_2827,N_2824);
or U2994 (N_2994,N_2866,N_2883);
nor U2995 (N_2995,N_2832,N_2879);
and U2996 (N_2996,N_2842,N_2870);
or U2997 (N_2997,N_2844,N_2826);
xor U2998 (N_2998,N_2857,N_2850);
xnor U2999 (N_2999,N_2872,N_2863);
and UO_0 (O_0,N_2906,N_2981);
nand UO_1 (O_1,N_2909,N_2970);
xor UO_2 (O_2,N_2976,N_2935);
nand UO_3 (O_3,N_2927,N_2922);
xnor UO_4 (O_4,N_2924,N_2932);
or UO_5 (O_5,N_2959,N_2993);
nand UO_6 (O_6,N_2961,N_2998);
xnor UO_7 (O_7,N_2996,N_2929);
or UO_8 (O_8,N_2963,N_2964);
and UO_9 (O_9,N_2943,N_2953);
xor UO_10 (O_10,N_2958,N_2928);
nand UO_11 (O_11,N_2999,N_2977);
nand UO_12 (O_12,N_2960,N_2946);
nand UO_13 (O_13,N_2967,N_2940);
and UO_14 (O_14,N_2915,N_2901);
xor UO_15 (O_15,N_2950,N_2936);
nand UO_16 (O_16,N_2908,N_2921);
xor UO_17 (O_17,N_2937,N_2989);
nor UO_18 (O_18,N_2955,N_2947);
xnor UO_19 (O_19,N_2972,N_2916);
xnor UO_20 (O_20,N_2983,N_2978);
or UO_21 (O_21,N_2905,N_2920);
and UO_22 (O_22,N_2973,N_2945);
xnor UO_23 (O_23,N_2995,N_2980);
or UO_24 (O_24,N_2985,N_2962);
and UO_25 (O_25,N_2968,N_2931);
xor UO_26 (O_26,N_2934,N_2956);
and UO_27 (O_27,N_2965,N_2949);
nor UO_28 (O_28,N_2942,N_2994);
nand UO_29 (O_29,N_2979,N_2918);
or UO_30 (O_30,N_2914,N_2971);
or UO_31 (O_31,N_2907,N_2987);
nor UO_32 (O_32,N_2957,N_2991);
xnor UO_33 (O_33,N_2919,N_2900);
xnor UO_34 (O_34,N_2966,N_2913);
or UO_35 (O_35,N_2939,N_2982);
xor UO_36 (O_36,N_2988,N_2904);
nand UO_37 (O_37,N_2969,N_2925);
xor UO_38 (O_38,N_2954,N_2948);
nand UO_39 (O_39,N_2984,N_2903);
nand UO_40 (O_40,N_2917,N_2997);
and UO_41 (O_41,N_2952,N_2974);
or UO_42 (O_42,N_2944,N_2910);
and UO_43 (O_43,N_2923,N_2938);
nor UO_44 (O_44,N_2990,N_2926);
xor UO_45 (O_45,N_2992,N_2951);
xor UO_46 (O_46,N_2941,N_2911);
nor UO_47 (O_47,N_2930,N_2912);
nand UO_48 (O_48,N_2902,N_2975);
and UO_49 (O_49,N_2933,N_2986);
xnor UO_50 (O_50,N_2978,N_2927);
nor UO_51 (O_51,N_2920,N_2983);
nor UO_52 (O_52,N_2933,N_2907);
nand UO_53 (O_53,N_2965,N_2952);
and UO_54 (O_54,N_2943,N_2982);
or UO_55 (O_55,N_2990,N_2901);
or UO_56 (O_56,N_2904,N_2966);
nor UO_57 (O_57,N_2990,N_2975);
nor UO_58 (O_58,N_2957,N_2919);
nand UO_59 (O_59,N_2979,N_2970);
xnor UO_60 (O_60,N_2914,N_2999);
nor UO_61 (O_61,N_2908,N_2960);
or UO_62 (O_62,N_2963,N_2957);
xor UO_63 (O_63,N_2983,N_2943);
xor UO_64 (O_64,N_2970,N_2960);
nor UO_65 (O_65,N_2935,N_2946);
and UO_66 (O_66,N_2985,N_2967);
nor UO_67 (O_67,N_2995,N_2940);
xor UO_68 (O_68,N_2974,N_2929);
xnor UO_69 (O_69,N_2921,N_2958);
nand UO_70 (O_70,N_2964,N_2971);
and UO_71 (O_71,N_2988,N_2952);
nand UO_72 (O_72,N_2984,N_2982);
nand UO_73 (O_73,N_2936,N_2945);
nand UO_74 (O_74,N_2931,N_2948);
nor UO_75 (O_75,N_2902,N_2959);
or UO_76 (O_76,N_2934,N_2922);
and UO_77 (O_77,N_2945,N_2964);
xnor UO_78 (O_78,N_2985,N_2943);
or UO_79 (O_79,N_2946,N_2943);
and UO_80 (O_80,N_2930,N_2957);
nor UO_81 (O_81,N_2960,N_2937);
xor UO_82 (O_82,N_2934,N_2992);
xnor UO_83 (O_83,N_2918,N_2928);
or UO_84 (O_84,N_2986,N_2924);
nand UO_85 (O_85,N_2953,N_2977);
xor UO_86 (O_86,N_2957,N_2908);
and UO_87 (O_87,N_2987,N_2959);
and UO_88 (O_88,N_2949,N_2963);
or UO_89 (O_89,N_2958,N_2991);
nand UO_90 (O_90,N_2997,N_2914);
and UO_91 (O_91,N_2981,N_2920);
nor UO_92 (O_92,N_2943,N_2929);
xnor UO_93 (O_93,N_2950,N_2917);
nand UO_94 (O_94,N_2971,N_2907);
nand UO_95 (O_95,N_2921,N_2938);
and UO_96 (O_96,N_2965,N_2979);
and UO_97 (O_97,N_2915,N_2968);
xor UO_98 (O_98,N_2909,N_2981);
and UO_99 (O_99,N_2986,N_2952);
or UO_100 (O_100,N_2900,N_2929);
nor UO_101 (O_101,N_2929,N_2911);
or UO_102 (O_102,N_2958,N_2906);
xor UO_103 (O_103,N_2930,N_2981);
nand UO_104 (O_104,N_2974,N_2962);
and UO_105 (O_105,N_2937,N_2968);
nand UO_106 (O_106,N_2929,N_2973);
nor UO_107 (O_107,N_2977,N_2949);
nor UO_108 (O_108,N_2931,N_2925);
or UO_109 (O_109,N_2903,N_2945);
and UO_110 (O_110,N_2927,N_2966);
nor UO_111 (O_111,N_2907,N_2955);
xor UO_112 (O_112,N_2986,N_2956);
nand UO_113 (O_113,N_2924,N_2923);
or UO_114 (O_114,N_2958,N_2988);
nand UO_115 (O_115,N_2906,N_2930);
or UO_116 (O_116,N_2952,N_2932);
xnor UO_117 (O_117,N_2951,N_2968);
nand UO_118 (O_118,N_2969,N_2988);
nand UO_119 (O_119,N_2963,N_2979);
nand UO_120 (O_120,N_2961,N_2931);
and UO_121 (O_121,N_2937,N_2905);
nor UO_122 (O_122,N_2936,N_2959);
and UO_123 (O_123,N_2919,N_2929);
and UO_124 (O_124,N_2993,N_2927);
nor UO_125 (O_125,N_2948,N_2918);
or UO_126 (O_126,N_2994,N_2932);
nand UO_127 (O_127,N_2919,N_2962);
xnor UO_128 (O_128,N_2950,N_2904);
nor UO_129 (O_129,N_2944,N_2909);
xor UO_130 (O_130,N_2990,N_2972);
nand UO_131 (O_131,N_2904,N_2936);
and UO_132 (O_132,N_2938,N_2903);
xor UO_133 (O_133,N_2939,N_2994);
and UO_134 (O_134,N_2964,N_2977);
and UO_135 (O_135,N_2930,N_2979);
or UO_136 (O_136,N_2928,N_2955);
nor UO_137 (O_137,N_2922,N_2983);
nor UO_138 (O_138,N_2948,N_2990);
xnor UO_139 (O_139,N_2966,N_2952);
or UO_140 (O_140,N_2988,N_2911);
nand UO_141 (O_141,N_2970,N_2973);
nand UO_142 (O_142,N_2969,N_2983);
and UO_143 (O_143,N_2940,N_2910);
xnor UO_144 (O_144,N_2942,N_2938);
or UO_145 (O_145,N_2908,N_2976);
or UO_146 (O_146,N_2995,N_2943);
and UO_147 (O_147,N_2901,N_2933);
or UO_148 (O_148,N_2963,N_2925);
and UO_149 (O_149,N_2991,N_2990);
xnor UO_150 (O_150,N_2970,N_2951);
nand UO_151 (O_151,N_2993,N_2957);
nand UO_152 (O_152,N_2931,N_2967);
nand UO_153 (O_153,N_2931,N_2950);
nand UO_154 (O_154,N_2955,N_2926);
xor UO_155 (O_155,N_2968,N_2920);
nand UO_156 (O_156,N_2938,N_2955);
and UO_157 (O_157,N_2943,N_2991);
or UO_158 (O_158,N_2919,N_2991);
nor UO_159 (O_159,N_2935,N_2971);
xor UO_160 (O_160,N_2988,N_2917);
xnor UO_161 (O_161,N_2967,N_2998);
xnor UO_162 (O_162,N_2950,N_2903);
and UO_163 (O_163,N_2916,N_2998);
xnor UO_164 (O_164,N_2911,N_2921);
nor UO_165 (O_165,N_2961,N_2971);
and UO_166 (O_166,N_2952,N_2969);
nand UO_167 (O_167,N_2935,N_2911);
nand UO_168 (O_168,N_2932,N_2991);
nand UO_169 (O_169,N_2938,N_2915);
nor UO_170 (O_170,N_2972,N_2943);
or UO_171 (O_171,N_2940,N_2952);
nand UO_172 (O_172,N_2933,N_2956);
nand UO_173 (O_173,N_2965,N_2966);
or UO_174 (O_174,N_2935,N_2997);
nor UO_175 (O_175,N_2923,N_2997);
xnor UO_176 (O_176,N_2986,N_2928);
xnor UO_177 (O_177,N_2984,N_2910);
xor UO_178 (O_178,N_2950,N_2933);
nor UO_179 (O_179,N_2923,N_2988);
or UO_180 (O_180,N_2944,N_2902);
or UO_181 (O_181,N_2994,N_2986);
and UO_182 (O_182,N_2956,N_2932);
nand UO_183 (O_183,N_2950,N_2945);
or UO_184 (O_184,N_2944,N_2948);
and UO_185 (O_185,N_2935,N_2960);
and UO_186 (O_186,N_2938,N_2925);
nor UO_187 (O_187,N_2992,N_2937);
and UO_188 (O_188,N_2982,N_2989);
nand UO_189 (O_189,N_2964,N_2979);
xnor UO_190 (O_190,N_2974,N_2916);
nor UO_191 (O_191,N_2967,N_2964);
nand UO_192 (O_192,N_2952,N_2921);
or UO_193 (O_193,N_2982,N_2947);
nor UO_194 (O_194,N_2955,N_2991);
xnor UO_195 (O_195,N_2908,N_2922);
nor UO_196 (O_196,N_2999,N_2979);
and UO_197 (O_197,N_2905,N_2907);
and UO_198 (O_198,N_2960,N_2901);
or UO_199 (O_199,N_2987,N_2928);
nand UO_200 (O_200,N_2991,N_2980);
and UO_201 (O_201,N_2987,N_2939);
or UO_202 (O_202,N_2979,N_2977);
and UO_203 (O_203,N_2906,N_2969);
nor UO_204 (O_204,N_2919,N_2911);
xor UO_205 (O_205,N_2922,N_2954);
xnor UO_206 (O_206,N_2940,N_2917);
nand UO_207 (O_207,N_2924,N_2939);
nand UO_208 (O_208,N_2928,N_2983);
or UO_209 (O_209,N_2918,N_2932);
nand UO_210 (O_210,N_2900,N_2970);
or UO_211 (O_211,N_2957,N_2902);
and UO_212 (O_212,N_2900,N_2942);
xor UO_213 (O_213,N_2901,N_2913);
xnor UO_214 (O_214,N_2983,N_2955);
nor UO_215 (O_215,N_2990,N_2950);
nor UO_216 (O_216,N_2912,N_2913);
xnor UO_217 (O_217,N_2973,N_2933);
nor UO_218 (O_218,N_2936,N_2908);
or UO_219 (O_219,N_2998,N_2900);
and UO_220 (O_220,N_2912,N_2965);
or UO_221 (O_221,N_2913,N_2905);
nor UO_222 (O_222,N_2927,N_2912);
xor UO_223 (O_223,N_2942,N_2928);
nor UO_224 (O_224,N_2985,N_2982);
nand UO_225 (O_225,N_2965,N_2929);
and UO_226 (O_226,N_2903,N_2941);
or UO_227 (O_227,N_2925,N_2906);
or UO_228 (O_228,N_2973,N_2990);
and UO_229 (O_229,N_2926,N_2901);
nor UO_230 (O_230,N_2905,N_2931);
or UO_231 (O_231,N_2989,N_2919);
and UO_232 (O_232,N_2958,N_2999);
nor UO_233 (O_233,N_2990,N_2957);
nand UO_234 (O_234,N_2975,N_2969);
nand UO_235 (O_235,N_2941,N_2973);
and UO_236 (O_236,N_2954,N_2934);
and UO_237 (O_237,N_2934,N_2990);
nand UO_238 (O_238,N_2925,N_2979);
xor UO_239 (O_239,N_2948,N_2984);
and UO_240 (O_240,N_2940,N_2988);
and UO_241 (O_241,N_2905,N_2980);
nand UO_242 (O_242,N_2975,N_2995);
xnor UO_243 (O_243,N_2960,N_2933);
or UO_244 (O_244,N_2944,N_2979);
or UO_245 (O_245,N_2987,N_2947);
or UO_246 (O_246,N_2960,N_2953);
and UO_247 (O_247,N_2947,N_2979);
xor UO_248 (O_248,N_2940,N_2980);
nor UO_249 (O_249,N_2950,N_2930);
nand UO_250 (O_250,N_2991,N_2984);
and UO_251 (O_251,N_2987,N_2977);
xnor UO_252 (O_252,N_2905,N_2919);
and UO_253 (O_253,N_2930,N_2999);
xor UO_254 (O_254,N_2927,N_2959);
nand UO_255 (O_255,N_2920,N_2930);
nand UO_256 (O_256,N_2911,N_2940);
nor UO_257 (O_257,N_2970,N_2929);
nand UO_258 (O_258,N_2903,N_2928);
xor UO_259 (O_259,N_2980,N_2908);
nand UO_260 (O_260,N_2926,N_2931);
xor UO_261 (O_261,N_2982,N_2913);
xor UO_262 (O_262,N_2998,N_2952);
xnor UO_263 (O_263,N_2969,N_2932);
nor UO_264 (O_264,N_2900,N_2958);
and UO_265 (O_265,N_2968,N_2979);
xor UO_266 (O_266,N_2912,N_2938);
xnor UO_267 (O_267,N_2968,N_2930);
and UO_268 (O_268,N_2974,N_2988);
xnor UO_269 (O_269,N_2981,N_2975);
and UO_270 (O_270,N_2970,N_2957);
and UO_271 (O_271,N_2988,N_2903);
nor UO_272 (O_272,N_2953,N_2973);
xnor UO_273 (O_273,N_2946,N_2967);
xor UO_274 (O_274,N_2936,N_2929);
nand UO_275 (O_275,N_2947,N_2958);
xor UO_276 (O_276,N_2924,N_2974);
xor UO_277 (O_277,N_2961,N_2930);
or UO_278 (O_278,N_2939,N_2980);
nand UO_279 (O_279,N_2987,N_2961);
xnor UO_280 (O_280,N_2947,N_2940);
nor UO_281 (O_281,N_2980,N_2910);
xor UO_282 (O_282,N_2981,N_2957);
xnor UO_283 (O_283,N_2912,N_2984);
and UO_284 (O_284,N_2983,N_2919);
nor UO_285 (O_285,N_2985,N_2930);
nand UO_286 (O_286,N_2900,N_2962);
or UO_287 (O_287,N_2951,N_2991);
nor UO_288 (O_288,N_2953,N_2975);
or UO_289 (O_289,N_2927,N_2980);
xor UO_290 (O_290,N_2936,N_2917);
or UO_291 (O_291,N_2951,N_2961);
and UO_292 (O_292,N_2909,N_2976);
nor UO_293 (O_293,N_2936,N_2949);
or UO_294 (O_294,N_2909,N_2933);
nand UO_295 (O_295,N_2969,N_2900);
xor UO_296 (O_296,N_2909,N_2930);
and UO_297 (O_297,N_2978,N_2964);
or UO_298 (O_298,N_2988,N_2930);
xor UO_299 (O_299,N_2974,N_2950);
nand UO_300 (O_300,N_2930,N_2929);
nor UO_301 (O_301,N_2920,N_2964);
xor UO_302 (O_302,N_2985,N_2984);
or UO_303 (O_303,N_2913,N_2986);
xnor UO_304 (O_304,N_2924,N_2959);
or UO_305 (O_305,N_2922,N_2984);
xnor UO_306 (O_306,N_2934,N_2963);
or UO_307 (O_307,N_2930,N_2984);
nor UO_308 (O_308,N_2999,N_2943);
and UO_309 (O_309,N_2958,N_2910);
nand UO_310 (O_310,N_2944,N_2965);
and UO_311 (O_311,N_2930,N_2940);
nor UO_312 (O_312,N_2935,N_2956);
nand UO_313 (O_313,N_2941,N_2980);
and UO_314 (O_314,N_2948,N_2988);
xor UO_315 (O_315,N_2900,N_2986);
or UO_316 (O_316,N_2904,N_2929);
or UO_317 (O_317,N_2970,N_2930);
nand UO_318 (O_318,N_2972,N_2961);
or UO_319 (O_319,N_2911,N_2958);
xnor UO_320 (O_320,N_2904,N_2955);
and UO_321 (O_321,N_2985,N_2987);
nand UO_322 (O_322,N_2940,N_2981);
or UO_323 (O_323,N_2917,N_2948);
and UO_324 (O_324,N_2992,N_2980);
xor UO_325 (O_325,N_2921,N_2968);
nor UO_326 (O_326,N_2994,N_2933);
or UO_327 (O_327,N_2960,N_2999);
nand UO_328 (O_328,N_2934,N_2966);
xnor UO_329 (O_329,N_2982,N_2914);
or UO_330 (O_330,N_2965,N_2972);
nand UO_331 (O_331,N_2939,N_2908);
nand UO_332 (O_332,N_2977,N_2920);
xor UO_333 (O_333,N_2960,N_2954);
nor UO_334 (O_334,N_2953,N_2909);
nor UO_335 (O_335,N_2966,N_2996);
nor UO_336 (O_336,N_2906,N_2917);
nor UO_337 (O_337,N_2962,N_2905);
xor UO_338 (O_338,N_2956,N_2916);
nand UO_339 (O_339,N_2922,N_2973);
xnor UO_340 (O_340,N_2977,N_2973);
or UO_341 (O_341,N_2974,N_2923);
nor UO_342 (O_342,N_2986,N_2978);
xnor UO_343 (O_343,N_2911,N_2920);
and UO_344 (O_344,N_2983,N_2975);
nand UO_345 (O_345,N_2950,N_2987);
nand UO_346 (O_346,N_2957,N_2953);
xor UO_347 (O_347,N_2935,N_2951);
and UO_348 (O_348,N_2908,N_2945);
nand UO_349 (O_349,N_2978,N_2914);
and UO_350 (O_350,N_2903,N_2987);
nor UO_351 (O_351,N_2917,N_2927);
nand UO_352 (O_352,N_2963,N_2967);
xnor UO_353 (O_353,N_2984,N_2916);
xnor UO_354 (O_354,N_2926,N_2969);
nand UO_355 (O_355,N_2958,N_2998);
nand UO_356 (O_356,N_2937,N_2969);
nand UO_357 (O_357,N_2924,N_2935);
nor UO_358 (O_358,N_2976,N_2931);
or UO_359 (O_359,N_2987,N_2974);
nand UO_360 (O_360,N_2956,N_2974);
nor UO_361 (O_361,N_2907,N_2906);
nand UO_362 (O_362,N_2983,N_2997);
and UO_363 (O_363,N_2983,N_2940);
nand UO_364 (O_364,N_2980,N_2976);
nor UO_365 (O_365,N_2979,N_2924);
nand UO_366 (O_366,N_2911,N_2902);
and UO_367 (O_367,N_2956,N_2973);
nand UO_368 (O_368,N_2927,N_2953);
and UO_369 (O_369,N_2986,N_2981);
xor UO_370 (O_370,N_2998,N_2996);
xnor UO_371 (O_371,N_2997,N_2981);
and UO_372 (O_372,N_2943,N_2986);
nor UO_373 (O_373,N_2944,N_2900);
nand UO_374 (O_374,N_2914,N_2975);
or UO_375 (O_375,N_2922,N_2915);
nand UO_376 (O_376,N_2993,N_2900);
and UO_377 (O_377,N_2928,N_2927);
nand UO_378 (O_378,N_2998,N_2917);
nor UO_379 (O_379,N_2976,N_2949);
and UO_380 (O_380,N_2964,N_2952);
nand UO_381 (O_381,N_2937,N_2900);
and UO_382 (O_382,N_2972,N_2966);
nor UO_383 (O_383,N_2920,N_2902);
and UO_384 (O_384,N_2959,N_2966);
and UO_385 (O_385,N_2929,N_2984);
and UO_386 (O_386,N_2942,N_2957);
nor UO_387 (O_387,N_2987,N_2940);
and UO_388 (O_388,N_2980,N_2971);
and UO_389 (O_389,N_2926,N_2965);
xor UO_390 (O_390,N_2914,N_2921);
nor UO_391 (O_391,N_2966,N_2912);
and UO_392 (O_392,N_2977,N_2932);
nor UO_393 (O_393,N_2929,N_2992);
xnor UO_394 (O_394,N_2992,N_2989);
and UO_395 (O_395,N_2958,N_2962);
xor UO_396 (O_396,N_2980,N_2902);
and UO_397 (O_397,N_2993,N_2980);
xor UO_398 (O_398,N_2946,N_2978);
xor UO_399 (O_399,N_2902,N_2997);
xor UO_400 (O_400,N_2982,N_2901);
nor UO_401 (O_401,N_2982,N_2955);
nand UO_402 (O_402,N_2957,N_2900);
or UO_403 (O_403,N_2904,N_2993);
nor UO_404 (O_404,N_2988,N_2996);
xor UO_405 (O_405,N_2952,N_2929);
nand UO_406 (O_406,N_2994,N_2985);
nor UO_407 (O_407,N_2906,N_2936);
and UO_408 (O_408,N_2948,N_2991);
xnor UO_409 (O_409,N_2945,N_2956);
nand UO_410 (O_410,N_2958,N_2901);
or UO_411 (O_411,N_2941,N_2923);
nor UO_412 (O_412,N_2970,N_2937);
or UO_413 (O_413,N_2906,N_2964);
and UO_414 (O_414,N_2950,N_2972);
or UO_415 (O_415,N_2929,N_2941);
nor UO_416 (O_416,N_2951,N_2932);
or UO_417 (O_417,N_2912,N_2902);
xor UO_418 (O_418,N_2994,N_2968);
nand UO_419 (O_419,N_2972,N_2930);
or UO_420 (O_420,N_2921,N_2985);
or UO_421 (O_421,N_2912,N_2994);
and UO_422 (O_422,N_2986,N_2991);
and UO_423 (O_423,N_2923,N_2908);
or UO_424 (O_424,N_2936,N_2983);
and UO_425 (O_425,N_2991,N_2967);
or UO_426 (O_426,N_2997,N_2944);
xnor UO_427 (O_427,N_2968,N_2962);
nand UO_428 (O_428,N_2909,N_2937);
and UO_429 (O_429,N_2954,N_2978);
nand UO_430 (O_430,N_2953,N_2918);
xnor UO_431 (O_431,N_2957,N_2922);
nand UO_432 (O_432,N_2961,N_2989);
xnor UO_433 (O_433,N_2953,N_2952);
nand UO_434 (O_434,N_2954,N_2946);
and UO_435 (O_435,N_2950,N_2935);
or UO_436 (O_436,N_2919,N_2941);
or UO_437 (O_437,N_2993,N_2929);
xor UO_438 (O_438,N_2968,N_2972);
nor UO_439 (O_439,N_2971,N_2985);
nand UO_440 (O_440,N_2968,N_2956);
xor UO_441 (O_441,N_2995,N_2970);
xnor UO_442 (O_442,N_2965,N_2982);
nand UO_443 (O_443,N_2971,N_2981);
nand UO_444 (O_444,N_2974,N_2942);
and UO_445 (O_445,N_2995,N_2937);
nand UO_446 (O_446,N_2927,N_2906);
and UO_447 (O_447,N_2938,N_2977);
nor UO_448 (O_448,N_2931,N_2924);
nor UO_449 (O_449,N_2934,N_2939);
nand UO_450 (O_450,N_2967,N_2984);
nor UO_451 (O_451,N_2946,N_2996);
nor UO_452 (O_452,N_2956,N_2960);
nand UO_453 (O_453,N_2921,N_2931);
nand UO_454 (O_454,N_2993,N_2934);
or UO_455 (O_455,N_2926,N_2975);
or UO_456 (O_456,N_2941,N_2928);
nor UO_457 (O_457,N_2924,N_2956);
or UO_458 (O_458,N_2937,N_2911);
nand UO_459 (O_459,N_2946,N_2904);
nand UO_460 (O_460,N_2905,N_2988);
xnor UO_461 (O_461,N_2962,N_2925);
or UO_462 (O_462,N_2980,N_2948);
nand UO_463 (O_463,N_2915,N_2984);
xor UO_464 (O_464,N_2939,N_2949);
and UO_465 (O_465,N_2960,N_2932);
nand UO_466 (O_466,N_2934,N_2937);
nand UO_467 (O_467,N_2916,N_2937);
and UO_468 (O_468,N_2918,N_2994);
or UO_469 (O_469,N_2945,N_2984);
nand UO_470 (O_470,N_2980,N_2983);
or UO_471 (O_471,N_2943,N_2949);
xor UO_472 (O_472,N_2911,N_2932);
nand UO_473 (O_473,N_2983,N_2952);
and UO_474 (O_474,N_2958,N_2954);
nor UO_475 (O_475,N_2976,N_2942);
xor UO_476 (O_476,N_2930,N_2944);
and UO_477 (O_477,N_2938,N_2943);
or UO_478 (O_478,N_2961,N_2981);
and UO_479 (O_479,N_2949,N_2997);
and UO_480 (O_480,N_2947,N_2974);
or UO_481 (O_481,N_2949,N_2942);
nor UO_482 (O_482,N_2965,N_2948);
or UO_483 (O_483,N_2979,N_2956);
and UO_484 (O_484,N_2907,N_2978);
nor UO_485 (O_485,N_2935,N_2949);
and UO_486 (O_486,N_2956,N_2952);
or UO_487 (O_487,N_2942,N_2970);
or UO_488 (O_488,N_2996,N_2952);
xnor UO_489 (O_489,N_2941,N_2955);
xnor UO_490 (O_490,N_2992,N_2996);
xor UO_491 (O_491,N_2940,N_2921);
nand UO_492 (O_492,N_2923,N_2992);
xor UO_493 (O_493,N_2928,N_2963);
and UO_494 (O_494,N_2958,N_2969);
xnor UO_495 (O_495,N_2906,N_2918);
or UO_496 (O_496,N_2958,N_2907);
and UO_497 (O_497,N_2948,N_2982);
nor UO_498 (O_498,N_2908,N_2990);
and UO_499 (O_499,N_2920,N_2973);
endmodule