module basic_3000_30000_3500_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_977,In_261);
nor U1 (N_1,In_2478,In_283);
and U2 (N_2,In_982,In_1707);
and U3 (N_3,In_1546,In_1490);
or U4 (N_4,In_409,In_2832);
nor U5 (N_5,In_1523,In_1702);
nor U6 (N_6,In_399,In_625);
xnor U7 (N_7,In_1522,In_585);
nor U8 (N_8,In_2129,In_486);
nor U9 (N_9,In_1206,In_1790);
xnor U10 (N_10,In_2161,In_1765);
or U11 (N_11,In_290,In_916);
nor U12 (N_12,In_2160,In_2250);
or U13 (N_13,In_1540,In_369);
nand U14 (N_14,In_2450,In_1963);
and U15 (N_15,In_2138,In_2088);
xnor U16 (N_16,In_1257,In_1741);
xnor U17 (N_17,In_2548,In_2216);
or U18 (N_18,In_1829,In_1681);
nand U19 (N_19,In_2744,In_1222);
nand U20 (N_20,In_1167,In_1500);
xor U21 (N_21,In_1809,In_209);
nor U22 (N_22,In_147,In_696);
nor U23 (N_23,In_887,In_843);
xor U24 (N_24,In_2612,In_1125);
or U25 (N_25,In_1210,In_1375);
or U26 (N_26,In_2259,In_2654);
nor U27 (N_27,In_186,In_262);
nor U28 (N_28,In_2868,In_947);
nor U29 (N_29,In_1435,In_2435);
xor U30 (N_30,In_1282,In_763);
xnor U31 (N_31,In_1641,In_650);
nor U32 (N_32,In_2419,In_2756);
or U33 (N_33,In_1460,In_35);
and U34 (N_34,In_1288,In_2877);
or U35 (N_35,In_2409,In_1563);
and U36 (N_36,In_467,In_2580);
nor U37 (N_37,In_2067,In_2164);
xnor U38 (N_38,In_928,In_2717);
and U39 (N_39,In_116,In_79);
nand U40 (N_40,In_374,In_195);
nand U41 (N_41,In_1584,In_2150);
or U42 (N_42,In_1545,In_1729);
nand U43 (N_43,In_2010,In_2027);
nor U44 (N_44,In_1305,In_2947);
xor U45 (N_45,In_2839,In_878);
or U46 (N_46,In_2555,In_1786);
xor U47 (N_47,In_1811,In_2403);
nand U48 (N_48,In_1823,In_1204);
xor U49 (N_49,In_2030,In_905);
nor U50 (N_50,In_1935,In_232);
xnor U51 (N_51,In_1273,In_239);
nor U52 (N_52,In_2091,In_767);
and U53 (N_53,In_280,In_1801);
xor U54 (N_54,In_2809,In_1440);
xor U55 (N_55,In_226,In_407);
xor U56 (N_56,In_2917,In_2763);
nor U57 (N_57,In_2694,In_2864);
xor U58 (N_58,In_1559,In_1624);
and U59 (N_59,In_2363,In_2649);
and U60 (N_60,In_250,In_1228);
or U61 (N_61,In_2799,In_552);
xnor U62 (N_62,In_670,In_1242);
nand U63 (N_63,In_1050,In_1560);
nand U64 (N_64,In_112,In_247);
and U65 (N_65,In_1620,In_826);
and U66 (N_66,In_2514,In_939);
nor U67 (N_67,In_1386,In_2821);
nand U68 (N_68,In_1915,In_2294);
or U69 (N_69,In_2162,In_786);
and U70 (N_70,In_635,In_1984);
xor U71 (N_71,In_1936,In_532);
xnor U72 (N_72,In_2255,In_199);
and U73 (N_73,In_1571,In_353);
nand U74 (N_74,In_1143,In_1197);
and U75 (N_75,In_1045,In_748);
nor U76 (N_76,In_141,In_2385);
nand U77 (N_77,In_851,In_1528);
nor U78 (N_78,In_614,In_2080);
nand U79 (N_79,In_727,In_298);
nand U80 (N_80,In_2495,In_729);
or U81 (N_81,In_2309,In_958);
nand U82 (N_82,In_2448,In_1223);
or U83 (N_83,In_2093,In_2099);
nor U84 (N_84,In_448,In_1609);
or U85 (N_85,In_1126,In_2107);
or U86 (N_86,In_1805,In_2794);
or U87 (N_87,In_1065,In_1855);
or U88 (N_88,In_2278,In_2315);
and U89 (N_89,In_1061,In_1712);
or U90 (N_90,In_1583,In_1083);
nand U91 (N_91,In_648,In_343);
or U92 (N_92,In_674,In_379);
xor U93 (N_93,In_1055,In_1006);
xnor U94 (N_94,In_2320,In_357);
or U95 (N_95,In_2764,In_2535);
and U96 (N_96,In_811,In_151);
xnor U97 (N_97,In_1142,In_1565);
xor U98 (N_98,In_436,In_2224);
and U99 (N_99,In_2253,In_15);
or U100 (N_100,In_1152,In_2279);
nand U101 (N_101,In_1369,In_153);
nor U102 (N_102,In_2970,In_2144);
xnor U103 (N_103,In_2571,In_2222);
xor U104 (N_104,In_1578,In_1286);
nor U105 (N_105,In_556,In_251);
and U106 (N_106,In_825,In_960);
xor U107 (N_107,In_2360,In_1437);
or U108 (N_108,In_801,In_1240);
or U109 (N_109,In_800,In_2540);
xor U110 (N_110,In_452,In_198);
or U111 (N_111,In_2956,In_1037);
nor U112 (N_112,In_1180,In_1726);
xor U113 (N_113,In_672,In_1157);
xor U114 (N_114,In_2190,In_1529);
nand U115 (N_115,In_967,In_282);
xor U116 (N_116,In_1830,In_1661);
and U117 (N_117,In_527,In_2355);
xor U118 (N_118,In_2273,In_1293);
or U119 (N_119,In_230,In_2802);
and U120 (N_120,In_645,In_496);
nor U121 (N_121,In_1209,In_565);
or U122 (N_122,In_1512,In_2042);
or U123 (N_123,In_708,In_2172);
nor U124 (N_124,In_533,In_215);
and U125 (N_125,In_653,In_1821);
nand U126 (N_126,In_1260,In_2750);
or U127 (N_127,In_986,In_161);
nand U128 (N_128,In_752,In_2441);
xnor U129 (N_129,In_2038,In_589);
or U130 (N_130,In_126,In_1053);
nor U131 (N_131,In_1817,In_654);
nand U132 (N_132,In_1414,In_679);
xnor U133 (N_133,In_2520,In_2240);
or U134 (N_134,In_624,In_2773);
xnor U135 (N_135,In_2288,In_1755);
or U136 (N_136,In_2589,In_2465);
or U137 (N_137,In_480,In_2163);
nor U138 (N_138,In_2728,In_2364);
nand U139 (N_139,In_1405,In_2426);
xor U140 (N_140,In_359,In_2840);
and U141 (N_141,In_2748,In_471);
or U142 (N_142,In_1219,In_1479);
nor U143 (N_143,In_1482,In_1682);
nand U144 (N_144,In_640,In_2967);
xnor U145 (N_145,In_1237,In_951);
or U146 (N_146,In_2818,In_2658);
and U147 (N_147,In_2875,In_1903);
or U148 (N_148,In_2433,In_2083);
nand U149 (N_149,In_1417,In_737);
or U150 (N_150,In_1919,In_2766);
xor U151 (N_151,In_1954,In_1113);
xor U152 (N_152,In_1275,In_2693);
or U153 (N_153,In_1011,In_520);
and U154 (N_154,In_2578,In_1879);
xnor U155 (N_155,In_1778,In_815);
and U156 (N_156,In_693,In_979);
or U157 (N_157,In_756,In_498);
nand U158 (N_158,In_1717,In_1870);
nor U159 (N_159,In_1110,In_2343);
and U160 (N_160,In_2213,In_85);
nor U161 (N_161,In_909,In_2014);
xor U162 (N_162,In_1983,In_2114);
nand U163 (N_163,In_2289,In_1756);
xnor U164 (N_164,In_48,In_1519);
nor U165 (N_165,In_2148,In_657);
nand U166 (N_166,In_1412,In_558);
nand U167 (N_167,In_34,In_2368);
nor U168 (N_168,In_2961,In_1456);
nand U169 (N_169,In_1996,In_2638);
nand U170 (N_170,In_349,In_1473);
and U171 (N_171,In_1942,In_1934);
xnor U172 (N_172,In_2301,In_864);
xnor U173 (N_173,In_1671,In_1947);
and U174 (N_174,In_2862,In_1388);
nor U175 (N_175,In_307,In_1602);
nor U176 (N_176,In_2545,In_1542);
or U177 (N_177,In_1981,In_1406);
nand U178 (N_178,In_2721,In_2290);
nand U179 (N_179,In_1186,In_2402);
and U180 (N_180,In_465,In_2122);
and U181 (N_181,In_2192,In_188);
xor U182 (N_182,In_1310,In_736);
xor U183 (N_183,In_1953,In_1588);
nand U184 (N_184,In_722,In_263);
nor U185 (N_185,In_1069,In_1202);
xnor U186 (N_186,In_516,In_812);
nor U187 (N_187,In_959,In_2401);
xor U188 (N_188,In_747,In_181);
nor U189 (N_189,In_2601,In_1130);
nand U190 (N_190,In_2878,In_707);
and U191 (N_191,In_509,In_666);
nor U192 (N_192,In_1887,In_2912);
and U193 (N_193,In_131,In_1526);
and U194 (N_194,In_2374,In_1941);
xor U195 (N_195,In_2859,In_411);
nand U196 (N_196,In_2068,In_2445);
nand U197 (N_197,In_718,In_1909);
nor U198 (N_198,In_726,In_761);
xnor U199 (N_199,In_2782,In_972);
xnor U200 (N_200,In_2032,In_1415);
nor U201 (N_201,In_2618,In_2047);
nor U202 (N_202,In_2817,In_2632);
and U203 (N_203,In_1844,In_1754);
nand U204 (N_204,In_1154,In_749);
nor U205 (N_205,In_375,In_472);
or U206 (N_206,In_1376,In_1471);
or U207 (N_207,In_381,In_210);
and U208 (N_208,In_1396,In_566);
or U209 (N_209,In_502,In_2275);
nor U210 (N_210,In_2991,In_2988);
xor U211 (N_211,In_55,In_2989);
or U212 (N_212,In_2220,In_2106);
and U213 (N_213,In_1502,In_1556);
and U214 (N_214,In_2537,In_1047);
nand U215 (N_215,In_1908,In_867);
xnor U216 (N_216,In_2183,In_2582);
and U217 (N_217,In_462,In_1561);
and U218 (N_218,In_636,In_2843);
and U219 (N_219,In_1929,In_2890);
xnor U220 (N_220,In_2924,In_2387);
nand U221 (N_221,In_1107,In_1692);
or U222 (N_222,In_969,In_2751);
or U223 (N_223,In_2217,In_1138);
and U224 (N_224,In_1030,In_1150);
nor U225 (N_225,In_1789,In_2134);
nor U226 (N_226,In_1873,In_100);
xnor U227 (N_227,In_1899,In_577);
xnor U228 (N_228,In_1510,In_507);
nor U229 (N_229,In_863,In_1378);
nor U230 (N_230,In_2040,In_2812);
or U231 (N_231,In_965,In_1626);
or U232 (N_232,In_490,In_628);
xor U233 (N_233,In_2999,In_1135);
or U234 (N_234,In_1436,In_553);
xnor U235 (N_235,In_1991,In_2367);
nor U236 (N_236,In_1859,In_1926);
nand U237 (N_237,In_306,In_1842);
or U238 (N_238,In_2560,In_351);
xor U239 (N_239,In_1785,In_2332);
or U240 (N_240,In_1749,In_1076);
and U241 (N_241,In_2889,In_1426);
nor U242 (N_242,In_1244,In_1646);
xor U243 (N_243,In_60,In_971);
and U244 (N_244,In_1965,In_2025);
xnor U245 (N_245,In_1910,In_2130);
and U246 (N_246,In_1283,In_1858);
nand U247 (N_247,In_1553,In_1973);
nor U248 (N_248,In_605,In_597);
or U249 (N_249,In_2118,In_166);
or U250 (N_250,In_1634,In_1835);
or U251 (N_251,In_2050,In_955);
and U252 (N_252,In_2270,In_2511);
nand U253 (N_253,In_1129,In_2709);
xnor U254 (N_254,In_2602,In_2542);
xnor U255 (N_255,In_1366,In_1400);
xor U256 (N_256,In_1916,In_1458);
and U257 (N_257,In_1800,In_832);
or U258 (N_258,In_389,In_1432);
or U259 (N_259,In_260,In_2786);
and U260 (N_260,In_740,In_214);
and U261 (N_261,In_76,In_1119);
or U262 (N_262,In_1351,In_97);
nor U263 (N_263,In_1007,In_2770);
nor U264 (N_264,In_2662,In_1487);
or U265 (N_265,In_2206,In_1196);
and U266 (N_266,In_2726,In_193);
or U267 (N_267,In_160,In_187);
nand U268 (N_268,In_83,In_2795);
nand U269 (N_269,In_1589,In_2120);
nor U270 (N_270,In_1339,In_2659);
or U271 (N_271,In_2311,In_824);
and U272 (N_272,In_2642,In_2123);
and U273 (N_273,In_1716,In_601);
nand U274 (N_274,In_1813,In_331);
nand U275 (N_275,In_363,In_329);
nand U276 (N_276,In_840,In_821);
and U277 (N_277,In_2729,In_2554);
nand U278 (N_278,In_1100,In_2378);
nand U279 (N_279,In_1886,In_1428);
and U280 (N_280,In_1267,In_78);
nand U281 (N_281,In_547,In_1014);
xnor U282 (N_282,In_2396,In_1198);
or U283 (N_283,In_63,In_933);
nand U284 (N_284,In_2824,In_2981);
xnor U285 (N_285,In_537,In_2377);
nand U286 (N_286,In_772,In_517);
or U287 (N_287,In_2796,In_643);
or U288 (N_288,In_775,In_600);
and U289 (N_289,In_368,In_1884);
xor U290 (N_290,In_994,In_2267);
nand U291 (N_291,In_963,In_253);
and U292 (N_292,In_220,In_1092);
or U293 (N_293,In_272,In_2407);
xor U294 (N_294,In_1596,In_639);
xnor U295 (N_295,In_1853,In_1799);
or U296 (N_296,In_2746,In_2485);
nor U297 (N_297,In_2317,In_2372);
xnor U298 (N_298,In_1552,In_1474);
or U299 (N_299,In_1469,In_1836);
and U300 (N_300,In_102,In_134);
xor U301 (N_301,In_1291,In_105);
xor U302 (N_302,In_1136,In_2140);
xor U303 (N_303,In_1639,In_164);
xor U304 (N_304,In_2425,In_482);
nand U305 (N_305,In_1466,In_1243);
and U306 (N_306,In_2675,In_1216);
and U307 (N_307,In_1160,In_192);
and U308 (N_308,In_1203,In_1678);
and U309 (N_309,In_1342,In_1311);
nand U310 (N_310,In_2062,In_567);
nor U311 (N_311,In_2547,In_2424);
nor U312 (N_312,In_1895,In_2430);
and U313 (N_313,In_2982,In_1539);
nand U314 (N_314,In_1647,In_394);
or U315 (N_315,In_2423,In_2242);
and U316 (N_316,In_1266,In_2826);
xnor U317 (N_317,In_177,In_2575);
nor U318 (N_318,In_421,In_897);
or U319 (N_319,In_2420,In_1940);
xor U320 (N_320,In_1327,In_2249);
nand U321 (N_321,In_2447,In_2888);
or U322 (N_322,In_1253,In_884);
nand U323 (N_323,In_2020,In_2539);
or U324 (N_324,In_50,In_1489);
xnor U325 (N_325,In_1874,In_1994);
or U326 (N_326,In_333,In_1501);
xnor U327 (N_327,In_1498,In_128);
and U328 (N_328,In_2035,In_106);
and U329 (N_329,In_858,In_795);
nand U330 (N_330,In_104,In_108);
and U331 (N_331,In_2918,In_549);
xnor U332 (N_332,In_1049,In_1604);
or U333 (N_333,In_390,In_629);
xnor U334 (N_334,In_2227,In_1331);
xnor U335 (N_335,In_776,In_1068);
xnor U336 (N_336,In_719,In_2631);
or U337 (N_337,In_990,In_1075);
or U338 (N_338,In_917,In_1323);
nand U339 (N_339,In_997,In_225);
or U340 (N_340,In_618,In_723);
and U341 (N_341,In_1306,In_2735);
nor U342 (N_342,In_1147,In_446);
xnor U343 (N_343,In_2440,In_1074);
xor U344 (N_344,In_1307,In_2212);
xor U345 (N_345,In_2059,In_823);
and U346 (N_346,In_114,In_2221);
xnor U347 (N_347,In_432,In_2530);
xor U348 (N_348,In_74,In_1766);
and U349 (N_349,In_352,In_1570);
nor U350 (N_350,In_2484,In_1279);
xnor U351 (N_351,In_1285,In_857);
xor U352 (N_352,In_2958,In_291);
xor U353 (N_353,In_2084,In_2215);
xnor U354 (N_354,In_1163,In_1493);
or U355 (N_355,In_129,In_2101);
nor U356 (N_356,In_2716,In_477);
and U357 (N_357,In_1820,In_185);
nand U358 (N_358,In_1290,In_1140);
and U359 (N_359,In_293,In_1680);
xor U360 (N_360,In_2234,In_2306);
nor U361 (N_361,In_2154,In_1742);
xor U362 (N_362,In_86,In_1188);
nand U363 (N_363,In_1608,In_1041);
xnor U364 (N_364,In_1404,In_458);
nand U365 (N_365,In_2634,In_2127);
or U366 (N_366,In_551,In_2933);
or U367 (N_367,In_2146,In_852);
nor U368 (N_368,In_65,In_339);
nor U369 (N_369,In_1254,In_2738);
nor U370 (N_370,In_1826,In_1381);
nand U371 (N_371,In_721,In_396);
nand U372 (N_372,In_925,In_2997);
xor U373 (N_373,In_2948,In_2962);
xor U374 (N_374,In_607,In_2855);
or U375 (N_375,In_2318,In_1961);
nand U376 (N_376,In_1166,In_1298);
nand U377 (N_377,In_109,In_142);
nand U378 (N_378,In_1643,In_277);
and U379 (N_379,In_2976,In_2641);
nor U380 (N_380,In_483,In_1434);
xor U381 (N_381,In_57,In_2561);
and U382 (N_382,In_1452,In_1613);
nor U383 (N_383,In_2284,In_2293);
nand U384 (N_384,In_2846,In_896);
nand U385 (N_385,In_1851,In_1695);
nand U386 (N_386,In_2473,In_1063);
nand U387 (N_387,In_2277,In_2685);
and U388 (N_388,In_438,In_289);
nand U389 (N_389,In_542,In_2849);
xor U390 (N_390,In_229,In_632);
or U391 (N_391,In_2645,In_2276);
nor U392 (N_392,In_1000,In_739);
nor U393 (N_393,In_1455,In_178);
or U394 (N_394,In_2321,In_2436);
nor U395 (N_395,In_1424,In_706);
or U396 (N_396,In_1576,In_1141);
xnor U397 (N_397,In_2668,In_2995);
nor U398 (N_398,In_2008,In_2048);
xor U399 (N_399,In_1776,In_554);
and U400 (N_400,In_1457,In_746);
nand U401 (N_401,In_768,In_1499);
xnor U402 (N_402,In_588,In_2004);
xor U403 (N_403,In_315,In_2701);
and U404 (N_404,In_2239,In_2153);
xor U405 (N_405,In_2866,In_1453);
xor U406 (N_406,In_256,In_847);
nor U407 (N_407,In_1700,In_459);
nand U408 (N_408,In_1619,In_2784);
or U409 (N_409,In_941,In_575);
or U410 (N_410,In_1794,In_2103);
xnor U411 (N_411,In_1393,In_2610);
xnor U412 (N_412,In_2087,In_2196);
nand U413 (N_413,In_1753,In_1042);
xnor U414 (N_414,In_1819,In_2117);
or U415 (N_415,In_921,In_1220);
xnor U416 (N_416,In_2951,In_405);
or U417 (N_417,In_1860,In_1346);
nand U418 (N_418,In_923,In_1162);
and U419 (N_419,In_1394,In_1956);
and U420 (N_420,In_197,In_1856);
or U421 (N_421,In_698,In_699);
or U422 (N_422,In_1697,In_1322);
and U423 (N_423,In_322,In_2953);
nor U424 (N_424,In_1121,In_1410);
nand U425 (N_425,In_464,In_455);
or U426 (N_426,In_660,In_1679);
nand U427 (N_427,In_1008,In_1230);
xnor U428 (N_428,In_2456,In_2937);
nor U429 (N_429,In_1399,In_2380);
and U430 (N_430,In_2235,In_2734);
nor U431 (N_431,In_107,In_2518);
xor U432 (N_432,In_1992,In_2965);
or U433 (N_433,In_1867,In_2522);
nor U434 (N_434,In_2126,In_2813);
nand U435 (N_435,In_2412,In_1825);
nand U436 (N_436,In_19,In_1084);
nor U437 (N_437,In_441,In_1673);
nand U438 (N_438,In_2266,In_1693);
and U439 (N_439,In_17,In_257);
or U440 (N_440,In_1839,In_2427);
nor U441 (N_441,In_2597,In_2673);
xnor U442 (N_442,In_1309,In_912);
nor U443 (N_443,In_1815,In_2665);
xor U444 (N_444,In_2931,In_1738);
and U445 (N_445,In_2200,In_2712);
and U446 (N_446,In_2149,In_572);
nor U447 (N_447,In_870,In_1328);
nand U448 (N_448,In_2667,In_694);
nand U449 (N_449,In_2324,In_2028);
and U450 (N_450,In_1029,In_2979);
or U451 (N_451,In_561,In_1944);
nor U452 (N_452,In_2174,In_1224);
xnor U453 (N_453,In_1684,In_442);
and U454 (N_454,In_2244,In_420);
or U455 (N_455,In_2243,In_1928);
and U456 (N_456,In_2417,In_391);
nand U457 (N_457,In_780,In_268);
and U458 (N_458,In_1615,In_2434);
xor U459 (N_459,In_817,In_136);
xor U460 (N_460,In_265,In_2339);
and U461 (N_461,In_2467,In_2202);
and U462 (N_462,In_1215,In_2934);
nand U463 (N_463,In_23,In_2102);
and U464 (N_464,In_222,In_2651);
nand U465 (N_465,In_1390,In_73);
nor U466 (N_466,In_2198,In_1669);
nor U467 (N_467,In_1017,In_886);
or U468 (N_468,In_1979,In_1046);
xor U469 (N_469,In_2218,In_2482);
nand U470 (N_470,In_145,In_2335);
xor U471 (N_471,In_1601,In_1054);
xor U472 (N_472,In_2652,In_2558);
xor U473 (N_473,In_1767,In_81);
nor U474 (N_474,In_1494,In_2406);
nor U475 (N_475,In_410,In_2731);
and U476 (N_476,In_2463,In_233);
and U477 (N_477,In_1304,In_1880);
xor U478 (N_478,In_980,In_2108);
xnor U479 (N_479,In_1579,In_2903);
nand U480 (N_480,In_2570,In_2525);
nand U481 (N_481,In_1795,In_2489);
nand U482 (N_482,In_1866,In_2136);
xnor U483 (N_483,In_2431,In_430);
and U484 (N_484,In_492,In_1861);
or U485 (N_485,In_2262,In_685);
xor U486 (N_486,In_2919,In_1509);
and U487 (N_487,In_712,In_1127);
nor U488 (N_488,In_926,In_2492);
nor U489 (N_489,In_32,In_1106);
nor U490 (N_490,In_299,In_1637);
nor U491 (N_491,In_665,In_1666);
and U492 (N_492,In_610,In_1170);
nand U493 (N_493,In_2392,In_2837);
and U494 (N_494,In_2619,In_809);
nor U495 (N_495,In_515,In_117);
nand U496 (N_496,In_877,In_1031);
or U497 (N_497,In_1497,In_1347);
or U498 (N_498,In_45,In_279);
xor U499 (N_499,In_1231,In_2119);
nor U500 (N_500,In_397,In_755);
nand U501 (N_501,In_2847,In_709);
and U502 (N_502,In_196,In_1642);
nand U503 (N_503,In_213,In_1218);
xor U504 (N_504,In_822,In_2993);
nand U505 (N_505,In_2481,In_695);
and U506 (N_506,In_127,In_619);
or U507 (N_507,In_705,In_2704);
and U508 (N_508,In_2541,In_2787);
xor U509 (N_509,In_1320,In_713);
nor U510 (N_510,In_750,In_1051);
nand U511 (N_511,In_2927,In_541);
and U512 (N_512,In_2376,In_1688);
xnor U513 (N_513,In_560,In_2280);
and U514 (N_514,In_1312,In_1177);
or U515 (N_515,In_2066,In_174);
or U516 (N_516,In_328,In_96);
xnor U517 (N_517,In_1907,In_2024);
nand U518 (N_518,In_1341,In_2806);
or U519 (N_519,In_2798,In_1397);
nand U520 (N_520,In_29,In_2310);
and U521 (N_521,In_2531,In_0);
nand U522 (N_522,In_120,In_1448);
nor U523 (N_523,In_2326,In_2022);
or U524 (N_524,In_1344,In_1080);
and U525 (N_525,In_816,In_1664);
nor U526 (N_526,In_2347,In_1101);
or U527 (N_527,In_2044,In_935);
and U528 (N_528,In_2769,In_1883);
xor U529 (N_529,In_1611,In_1402);
or U530 (N_530,In_1207,In_2488);
or U531 (N_531,In_207,In_663);
xnor U532 (N_532,In_1403,In_595);
xor U533 (N_533,In_1833,In_702);
xnor U534 (N_534,In_434,In_992);
and U535 (N_535,In_1264,In_1952);
nand U536 (N_536,In_2745,In_2606);
or U537 (N_537,In_31,In_1099);
xor U538 (N_538,In_1768,In_2723);
xor U539 (N_539,In_899,In_1772);
xnor U540 (N_540,In_1052,In_2534);
and U541 (N_541,In_1333,In_1134);
xor U542 (N_542,In_954,In_1590);
or U543 (N_543,In_376,In_2319);
or U544 (N_544,In_1299,In_2983);
nand U545 (N_545,In_710,In_804);
nor U546 (N_546,In_2669,In_2851);
or U547 (N_547,In_297,In_2180);
or U548 (N_548,In_2232,In_58);
nor U549 (N_549,In_1889,In_1277);
or U550 (N_550,In_59,In_2105);
nand U551 (N_551,In_1164,In_525);
xor U552 (N_552,In_205,In_1597);
and U553 (N_553,In_1718,In_2480);
or U554 (N_554,In_2264,In_2604);
nand U555 (N_555,In_2305,In_2600);
xnor U556 (N_556,In_2354,In_2361);
and U557 (N_557,In_2168,In_2453);
or U558 (N_558,In_1904,In_1371);
nand U559 (N_559,In_47,In_2);
nand U560 (N_560,In_2271,In_1373);
nor U561 (N_561,In_43,In_295);
xnor U562 (N_562,In_808,In_1308);
nand U563 (N_563,In_2543,In_742);
and U564 (N_564,In_1481,In_522);
and U565 (N_565,In_123,In_902);
nor U566 (N_566,In_845,In_2886);
xnor U567 (N_567,In_534,In_2583);
or U568 (N_568,In_2922,In_2727);
and U569 (N_569,In_2767,In_2538);
nor U570 (N_570,In_336,In_678);
nor U571 (N_571,In_2132,In_231);
nor U572 (N_572,In_765,In_165);
or U573 (N_573,In_563,In_1548);
nor U574 (N_574,In_356,In_1562);
xnor U575 (N_575,In_1574,In_1221);
xnor U576 (N_576,In_1118,In_2098);
xor U577 (N_577,In_2056,In_1102);
and U578 (N_578,In_1838,In_1040);
or U579 (N_579,In_182,In_1868);
xnor U580 (N_580,In_2269,In_2792);
xor U581 (N_581,In_501,In_2331);
or U582 (N_582,In_2743,In_985);
nand U583 (N_583,In_2774,In_2998);
xnor U584 (N_584,In_661,In_2759);
or U585 (N_585,In_2852,In_2475);
and U586 (N_586,In_288,In_1969);
or U587 (N_587,In_485,In_2646);
xor U588 (N_588,In_212,In_2381);
nor U589 (N_589,In_2295,In_92);
nor U590 (N_590,In_1467,In_2089);
nand U591 (N_591,In_1775,In_898);
or U592 (N_592,In_1193,In_2238);
nand U593 (N_593,In_206,In_1200);
nand U594 (N_594,In_2788,In_403);
nand U595 (N_595,In_819,In_856);
nand U596 (N_596,In_1964,In_701);
nand U597 (N_597,In_2258,In_14);
nor U598 (N_598,In_223,In_2247);
or U599 (N_599,In_2353,In_1108);
or U600 (N_600,In_1161,N_214);
and U601 (N_601,In_2116,N_248);
nor U602 (N_602,In_568,In_1212);
nand U603 (N_603,In_1443,N_28);
nand U604 (N_604,In_2850,In_1337);
nand U605 (N_605,N_390,In_400);
nor U606 (N_606,N_407,N_186);
nor U607 (N_607,In_2464,In_2472);
xor U608 (N_608,N_165,In_1806);
nor U609 (N_609,N_182,N_552);
or U610 (N_610,In_866,In_2179);
and U611 (N_611,In_1241,N_419);
xor U612 (N_612,N_446,In_36);
xnor U613 (N_613,In_830,In_2584);
nor U614 (N_614,N_102,N_574);
nor U615 (N_615,In_194,In_264);
xor U616 (N_616,In_2771,In_1998);
and U617 (N_617,In_1841,In_2758);
xor U618 (N_618,In_18,In_1238);
or U619 (N_619,In_1518,N_23);
xor U620 (N_620,In_1740,In_1495);
or U621 (N_621,In_1010,In_2446);
nor U622 (N_622,N_358,In_895);
xor U623 (N_623,In_38,In_2041);
and U624 (N_624,N_408,N_157);
nor U625 (N_625,In_2256,N_449);
and U626 (N_626,In_2308,N_149);
nand U627 (N_627,In_1854,In_1530);
nand U628 (N_628,In_1364,In_364);
and U629 (N_629,In_861,In_2887);
xor U630 (N_630,In_2666,In_1986);
nand U631 (N_631,In_1737,In_2410);
xor U632 (N_632,N_107,In_10);
nand U633 (N_633,In_1950,N_239);
nand U634 (N_634,In_1656,In_1326);
nor U635 (N_635,In_1771,In_1703);
nand U636 (N_636,In_1175,In_1095);
nor U637 (N_637,In_1392,In_367);
and U638 (N_638,In_1822,N_267);
xnor U639 (N_639,In_2705,In_2753);
xnor U640 (N_640,In_466,N_270);
xor U641 (N_641,In_1148,In_1477);
or U642 (N_642,N_247,In_1592);
xor U643 (N_643,In_2444,In_1527);
xnor U644 (N_644,In_2272,In_1663);
or U645 (N_645,In_68,In_741);
or U646 (N_646,In_2848,In_427);
nand U647 (N_647,In_449,In_1536);
nand U648 (N_648,N_299,In_2252);
nor U649 (N_649,In_2552,In_2205);
nor U650 (N_650,N_123,In_613);
or U651 (N_651,In_2055,N_93);
nand U652 (N_652,In_524,N_453);
nor U653 (N_653,In_938,N_474);
or U654 (N_654,In_2757,In_132);
or U655 (N_655,N_264,N_370);
nor U656 (N_656,In_2690,In_1199);
xnor U657 (N_657,In_2072,In_692);
and U658 (N_658,In_155,In_386);
and U659 (N_659,In_169,In_1617);
and U660 (N_660,In_2857,In_1289);
and U661 (N_661,In_1631,In_2082);
or U662 (N_662,N_50,In_743);
or U663 (N_663,In_2230,N_126);
and U664 (N_664,In_652,In_1777);
xnor U665 (N_665,N_409,N_8);
xor U666 (N_666,In_2687,In_1922);
xnor U667 (N_667,In_848,In_1834);
nand U668 (N_668,In_1659,In_1343);
xnor U669 (N_669,In_2603,N_205);
xnor U670 (N_670,In_1002,In_2366);
xor U671 (N_671,N_582,In_2452);
nor U672 (N_672,In_2755,In_798);
and U673 (N_673,In_1213,N_535);
nand U674 (N_674,In_724,N_155);
or U675 (N_675,In_1185,In_1862);
xnor U676 (N_676,In_2896,N_98);
or U677 (N_677,In_688,N_240);
nand U678 (N_678,N_135,In_2971);
xnor U679 (N_679,In_447,In_751);
xnor U680 (N_680,In_2057,N_278);
or U681 (N_681,In_2017,In_1783);
nand U682 (N_682,In_1531,In_1653);
nand U683 (N_683,In_189,In_2382);
xor U684 (N_684,In_2874,In_2015);
nand U685 (N_685,In_834,In_1486);
nor U686 (N_686,In_2710,N_485);
xor U687 (N_687,In_1524,N_563);
or U688 (N_688,N_96,N_215);
nor U689 (N_689,In_2911,N_502);
nor U690 (N_690,N_41,N_164);
or U691 (N_691,In_1808,In_675);
nand U692 (N_692,N_385,In_2898);
and U693 (N_693,In_87,In_392);
nand U694 (N_694,In_2487,In_2429);
nand U695 (N_695,In_1111,N_325);
or U696 (N_696,In_1086,N_501);
and U697 (N_697,In_146,N_323);
nor U698 (N_698,In_2966,In_1980);
nor U699 (N_699,In_1967,In_1598);
or U700 (N_700,N_297,In_623);
nand U701 (N_701,In_115,N_290);
or U702 (N_702,In_470,In_799);
nor U703 (N_703,N_48,N_181);
xnor U704 (N_704,In_44,In_716);
xnor U705 (N_705,In_814,In_2749);
xor U706 (N_706,In_2340,In_1782);
or U707 (N_707,N_412,N_331);
and U708 (N_708,N_343,In_831);
or U709 (N_709,In_850,In_2139);
xnor U710 (N_710,In_495,In_828);
xnor U711 (N_711,In_2486,N_303);
nand U712 (N_712,In_1449,N_260);
nand U713 (N_713,N_201,In_499);
xnor U714 (N_714,N_287,In_891);
nor U715 (N_715,In_1094,In_1704);
xor U716 (N_716,In_598,In_1995);
nor U717 (N_717,In_2237,N_46);
xor U718 (N_718,In_1593,N_472);
xnor U719 (N_719,In_2636,In_2775);
nor U720 (N_720,In_1920,In_1009);
nor U721 (N_721,In_2458,In_2894);
nor U722 (N_722,In_1255,N_119);
nor U723 (N_723,In_1923,N_572);
xor U724 (N_724,In_1116,N_122);
xnor U725 (N_725,In_875,In_2663);
or U726 (N_726,In_1211,N_512);
or U727 (N_727,In_1,In_1227);
xor U728 (N_728,In_2655,In_1599);
and U729 (N_729,N_544,In_2708);
and U730 (N_730,N_140,In_1751);
and U731 (N_731,In_1724,In_56);
nor U732 (N_732,In_759,In_2173);
or U733 (N_733,In_1462,N_256);
and U734 (N_734,In_931,In_70);
and U735 (N_735,In_1594,In_2110);
nor U736 (N_736,In_176,N_86);
or U737 (N_737,N_583,In_2002);
xnor U738 (N_738,In_1516,In_1319);
nor U739 (N_739,In_855,In_1810);
nor U740 (N_740,N_450,N_371);
nor U741 (N_741,In_612,In_2231);
nand U742 (N_742,In_37,In_1492);
xnor U743 (N_743,N_337,In_1128);
nand U744 (N_744,In_3,In_69);
nor U745 (N_745,In_1674,In_673);
nand U746 (N_746,In_1654,N_142);
or U747 (N_747,N_231,In_422);
or U748 (N_748,In_2455,N_243);
xnor U749 (N_749,In_1115,In_1640);
or U750 (N_750,In_2576,In_846);
nor U751 (N_751,In_91,In_383);
and U752 (N_752,N_457,N_133);
nand U753 (N_753,In_984,In_578);
nand U754 (N_754,In_52,N_2);
or U755 (N_755,In_2245,N_352);
or U756 (N_756,In_2702,N_471);
and U757 (N_757,N_551,N_549);
nand U758 (N_758,In_249,N_425);
and U759 (N_759,In_1869,N_232);
nor U760 (N_760,In_2805,In_494);
and U761 (N_761,In_2167,N_53);
nor U762 (N_762,N_275,N_241);
nand U763 (N_763,N_249,In_493);
nor U764 (N_764,N_382,In_419);
xnor U765 (N_765,In_2815,In_1214);
nand U766 (N_766,In_423,In_1551);
and U767 (N_767,N_105,In_2608);
nand U768 (N_768,N_17,N_480);
or U769 (N_769,In_1365,In_1287);
nor U770 (N_770,In_1621,In_757);
xor U771 (N_771,N_368,In_966);
xor U772 (N_772,N_265,In_1691);
or U773 (N_773,In_2954,N_542);
and U774 (N_774,N_519,N_513);
or U775 (N_775,In_1335,In_677);
nand U776 (N_776,In_478,In_2929);
and U777 (N_777,In_1408,In_2031);
nand U778 (N_778,N_596,In_11);
nor U779 (N_779,In_1900,In_2691);
nor U780 (N_780,In_2978,In_2957);
or U781 (N_781,In_2791,In_1533);
or U782 (N_782,In_259,In_1349);
or U783 (N_783,In_2349,In_2814);
xnor U784 (N_784,In_655,In_952);
and U785 (N_785,In_2370,In_1630);
nand U786 (N_786,In_2637,N_114);
or U787 (N_787,N_555,N_137);
or U788 (N_788,N_389,In_2819);
nor U789 (N_789,In_2064,In_676);
nor U790 (N_790,N_4,In_2574);
or U791 (N_791,In_1345,N_252);
or U792 (N_792,In_2037,In_1235);
nor U793 (N_793,N_578,In_2647);
and U794 (N_794,In_2133,In_1875);
xnor U795 (N_795,In_201,In_2009);
xnor U796 (N_796,In_2208,In_2049);
nand U797 (N_797,In_2007,In_703);
or U798 (N_798,N_245,In_2474);
xnor U799 (N_799,In_649,In_2483);
xor U800 (N_800,In_488,In_111);
nor U801 (N_801,N_68,In_2437);
xnor U802 (N_802,In_2466,N_112);
and U803 (N_803,In_1169,In_1391);
xnor U804 (N_804,In_1807,In_975);
nor U805 (N_805,In_1419,In_1504);
xnor U806 (N_806,N_575,In_642);
nor U807 (N_807,N_5,In_1444);
xor U808 (N_808,In_2674,In_778);
and U809 (N_809,N_300,N_174);
nor U810 (N_810,N_379,N_286);
or U811 (N_811,In_586,In_1831);
nand U812 (N_812,In_2838,N_302);
xor U813 (N_813,In_738,In_2336);
nand U814 (N_814,In_2479,In_1261);
nand U815 (N_815,In_518,N_579);
nor U816 (N_816,In_1387,N_345);
and U817 (N_817,In_2628,In_93);
nand U818 (N_818,N_550,In_914);
and U819 (N_819,In_2737,In_2241);
nor U820 (N_820,N_349,In_1367);
or U821 (N_821,In_792,In_1912);
nor U822 (N_822,N_393,In_1350);
or U823 (N_823,In_1062,In_2207);
xnor U824 (N_824,In_1361,In_1968);
nand U825 (N_825,In_2348,In_2046);
nor U826 (N_826,In_1580,N_363);
nand U827 (N_827,In_2341,In_20);
nand U828 (N_828,In_2975,In_1066);
and U829 (N_829,In_1759,N_335);
or U830 (N_830,In_244,N_71);
xor U831 (N_831,In_1787,In_51);
xnor U832 (N_832,In_2707,In_946);
or U833 (N_833,N_196,In_627);
nor U834 (N_834,In_773,In_2350);
xor U835 (N_835,N_304,In_2713);
nand U836 (N_836,N_191,In_820);
and U837 (N_837,In_2404,N_6);
nand U838 (N_838,In_1575,In_1374);
nand U839 (N_839,N_159,N_416);
nor U840 (N_840,In_1093,In_927);
xor U841 (N_841,In_1739,In_942);
nor U842 (N_842,In_1475,In_208);
nand U843 (N_843,N_422,In_13);
nand U844 (N_844,In_2706,In_33);
nor U845 (N_845,In_2568,In_216);
xor U846 (N_846,In_2013,In_2682);
and U847 (N_847,N_79,N_455);
or U848 (N_848,In_54,In_2058);
nand U849 (N_849,In_961,N_59);
nor U850 (N_850,N_80,N_13);
xnor U851 (N_851,In_2930,In_2457);
xor U852 (N_852,In_267,In_753);
nor U853 (N_853,In_838,In_1706);
and U854 (N_854,In_2346,N_439);
nor U855 (N_855,In_1098,In_190);
nand U856 (N_856,N_198,In_957);
or U857 (N_857,In_1451,N_70);
nand U858 (N_858,In_1156,In_7);
xor U859 (N_859,In_2635,In_2203);
nand U860 (N_860,In_2777,In_1377);
and U861 (N_861,N_289,In_1694);
and U862 (N_862,N_508,In_1433);
nor U863 (N_863,In_2016,In_2005);
and U864 (N_864,N_108,In_2143);
and U865 (N_865,N_170,N_334);
nor U866 (N_866,In_1623,In_793);
or U867 (N_867,In_2670,In_1383);
nand U868 (N_868,In_468,In_1849);
xor U869 (N_869,In_2512,In_2060);
xor U870 (N_870,In_1758,In_2334);
nor U871 (N_871,In_340,In_308);
or U872 (N_872,In_2351,In_2371);
nor U873 (N_873,In_511,N_294);
xnor U874 (N_874,In_2939,In_2251);
or U875 (N_875,In_827,In_2633);
or U876 (N_876,In_2454,In_1784);
nand U877 (N_877,In_1229,In_475);
and U878 (N_878,N_558,N_136);
and U879 (N_879,In_1544,In_2940);
or U880 (N_880,N_423,In_2990);
or U881 (N_881,In_77,In_2664);
nand U882 (N_882,In_1762,N_58);
nor U883 (N_883,In_1464,In_66);
xor U884 (N_884,N_242,In_777);
xor U885 (N_885,N_106,In_2357);
and U886 (N_886,In_1179,In_2100);
or U887 (N_887,In_2556,In_1649);
xor U888 (N_888,In_347,N_479);
or U889 (N_889,In_2388,N_282);
nor U890 (N_890,N_259,In_2863);
or U891 (N_891,In_88,In_1336);
nand U892 (N_892,In_523,N_21);
xor U893 (N_893,In_2630,N_127);
nand U894 (N_894,In_2345,N_128);
nand U895 (N_895,In_2718,In_2678);
or U896 (N_896,In_286,In_445);
and U897 (N_897,N_475,In_140);
nor U898 (N_898,In_2626,In_2236);
nand U899 (N_899,In_270,In_1997);
and U900 (N_900,In_2124,In_1015);
or U901 (N_901,In_474,In_2394);
and U902 (N_902,In_910,In_700);
or U903 (N_903,In_1358,In_388);
and U904 (N_904,N_324,In_1525);
nand U905 (N_905,In_217,N_566);
xor U906 (N_906,In_543,In_684);
nand U907 (N_907,N_236,N_307);
nand U908 (N_908,N_380,N_220);
and U909 (N_909,In_1446,In_1857);
xor U910 (N_910,N_418,In_573);
xor U911 (N_911,N_541,In_732);
or U912 (N_912,In_2960,In_626);
nand U913 (N_913,N_318,In_2861);
xor U914 (N_914,N_11,In_658);
nor U915 (N_915,N_110,In_2557);
xnor U916 (N_916,In_2359,N_178);
nor U917 (N_917,In_2563,N_74);
xnor U918 (N_918,In_562,N_65);
and U919 (N_919,In_2418,N_18);
nand U920 (N_920,In_770,In_1450);
nand U921 (N_921,In_158,In_2462);
nand U922 (N_922,In_2147,In_1603);
or U923 (N_923,In_1089,In_2095);
and U924 (N_924,In_987,In_1025);
nor U925 (N_925,In_2856,In_2286);
nor U926 (N_926,N_546,In_1330);
nand U927 (N_927,In_1779,In_2779);
and U928 (N_928,N_261,N_312);
xor U929 (N_929,In_1827,N_567);
nor U930 (N_930,In_2871,In_617);
xor U931 (N_931,In_2296,In_1088);
and U932 (N_932,N_153,N_35);
nor U933 (N_933,In_686,In_1722);
and U934 (N_934,N_208,In_1357);
xor U935 (N_935,In_2656,In_1757);
or U936 (N_936,In_2155,In_1798);
or U937 (N_937,In_1003,N_520);
or U938 (N_938,N_43,In_1208);
or U939 (N_939,In_378,In_200);
and U940 (N_940,N_104,In_248);
nor U941 (N_941,In_2867,N_362);
nand U942 (N_942,In_888,N_384);
or U943 (N_943,In_2411,In_2026);
nand U944 (N_944,N_590,In_296);
nand U945 (N_945,In_1249,In_1058);
xor U946 (N_946,In_901,In_571);
and U947 (N_947,In_2926,In_294);
nand U948 (N_948,N_223,In_1297);
nor U949 (N_949,In_240,In_2092);
xnor U950 (N_950,N_253,In_1315);
xor U951 (N_951,In_769,N_111);
nor U952 (N_952,N_52,N_448);
nand U953 (N_953,In_1271,In_2551);
or U954 (N_954,In_365,In_1389);
xor U955 (N_955,N_234,In_1988);
and U956 (N_956,In_236,In_2505);
or U957 (N_957,N_154,In_1946);
nand U958 (N_958,In_2595,In_406);
and U959 (N_959,In_2302,In_1797);
and U960 (N_960,In_144,N_301);
nor U961 (N_961,In_1348,In_1773);
xnor U962 (N_962,In_2959,In_1139);
and U963 (N_963,In_574,In_2204);
xor U964 (N_964,In_500,In_2695);
xnor U965 (N_965,In_2257,In_2006);
xor U966 (N_966,In_2018,In_544);
and U967 (N_967,N_117,In_1262);
or U968 (N_968,In_2768,In_337);
xor U969 (N_969,In_2128,In_2137);
nand U970 (N_970,In_1149,In_680);
xor U971 (N_971,In_1657,In_454);
xnor U972 (N_972,In_1962,N_160);
nand U973 (N_973,In_2383,In_1605);
or U974 (N_974,N_180,N_483);
nor U975 (N_975,In_671,N_92);
nor U976 (N_976,In_504,In_2921);
and U977 (N_977,In_1097,In_211);
nor U978 (N_978,In_1752,N_592);
or U979 (N_979,In_424,In_2661);
or U980 (N_980,In_936,N_16);
xor U981 (N_981,N_426,N_585);
and U982 (N_982,N_190,In_414);
or U983 (N_983,In_2104,In_2562);
nand U984 (N_984,In_2181,In_2913);
nand U985 (N_985,In_2395,In_1993);
nand U986 (N_986,In_1582,In_631);
xnor U987 (N_987,In_1155,In_842);
nand U988 (N_988,In_2599,In_2151);
or U989 (N_989,In_2219,In_443);
and U990 (N_990,In_1747,In_555);
or U991 (N_991,In_1708,In_1480);
xor U992 (N_992,N_398,In_1517);
or U993 (N_993,N_456,In_981);
or U994 (N_994,In_2615,In_1422);
nor U995 (N_995,In_668,N_101);
nor U996 (N_996,N_199,In_1792);
nor U997 (N_997,In_1256,In_227);
or U998 (N_998,In_1848,In_481);
nand U999 (N_999,In_2389,N_293);
or U1000 (N_1000,In_2329,In_1901);
nor U1001 (N_1001,In_408,N_310);
or U1002 (N_1002,In_1958,In_803);
nor U1003 (N_1003,In_1733,In_255);
nor U1004 (N_1004,N_533,In_2607);
nand U1005 (N_1005,N_429,N_272);
and U1006 (N_1006,In_2063,In_450);
or U1007 (N_1007,N_573,In_21);
nand U1008 (N_1008,In_1190,In_2648);
nand U1009 (N_1009,In_1018,In_234);
nor U1010 (N_1010,In_149,In_1555);
xor U1011 (N_1011,N_66,In_2169);
xor U1012 (N_1012,N_328,N_490);
and U1013 (N_1013,In_1728,In_1975);
or U1014 (N_1014,In_999,In_2325);
xor U1015 (N_1015,In_871,In_2451);
nor U1016 (N_1016,In_930,N_373);
xor U1017 (N_1017,In_284,In_1711);
nand U1018 (N_1018,N_524,In_2811);
nand U1019 (N_1019,N_32,In_754);
nor U1020 (N_1020,N_64,In_2972);
and U1021 (N_1021,In_323,In_929);
nor U1022 (N_1022,In_1748,In_1918);
xor U1023 (N_1023,In_2248,N_376);
xnor U1024 (N_1024,In_22,In_2804);
nor U1025 (N_1025,N_591,In_2827);
xor U1026 (N_1026,In_2184,In_876);
xor U1027 (N_1027,In_1818,In_2323);
nand U1028 (N_1028,N_129,In_2094);
nand U1029 (N_1029,In_1927,In_2698);
nand U1030 (N_1030,In_1824,In_1013);
and U1031 (N_1031,N_507,In_2725);
xor U1032 (N_1032,In_682,In_1852);
and U1033 (N_1033,In_2807,In_2553);
nor U1034 (N_1034,In_1484,In_854);
xnor U1035 (N_1035,In_1251,In_1938);
and U1036 (N_1036,In_2679,N_273);
nand U1037 (N_1037,In_2590,In_2086);
nor U1038 (N_1038,N_187,N_531);
or U1039 (N_1039,In_2730,In_2895);
nand U1040 (N_1040,In_1635,In_584);
xnor U1041 (N_1041,In_604,In_2754);
nand U1042 (N_1042,In_662,In_184);
xor U1043 (N_1043,In_880,In_2358);
or U1044 (N_1044,N_491,In_305);
nor U1045 (N_1045,N_15,In_2468);
and U1046 (N_1046,In_802,In_1158);
xnor U1047 (N_1047,In_630,In_667);
nand U1048 (N_1048,In_203,N_411);
nor U1049 (N_1049,In_460,In_974);
or U1050 (N_1050,In_2533,In_2935);
nor U1051 (N_1051,N_469,In_2621);
xor U1052 (N_1052,In_1736,N_298);
and U1053 (N_1053,In_1760,N_88);
nor U1054 (N_1054,In_1709,In_1362);
and U1055 (N_1055,In_2061,In_1989);
nand U1056 (N_1056,In_2797,N_100);
and U1057 (N_1057,In_2158,In_512);
nand U1058 (N_1058,In_1112,In_2494);
xor U1059 (N_1059,N_266,In_1793);
nand U1060 (N_1060,N_235,In_497);
and U1061 (N_1061,In_892,In_8);
xnor U1062 (N_1062,In_1276,In_1607);
or U1063 (N_1063,In_1557,N_217);
or U1064 (N_1064,In_6,In_80);
and U1065 (N_1065,In_1295,In_783);
nand U1066 (N_1066,In_1696,In_2157);
xor U1067 (N_1067,In_995,N_354);
xnor U1068 (N_1068,In_620,N_75);
and U1069 (N_1069,N_210,In_1955);
xnor U1070 (N_1070,In_2677,In_1902);
nor U1071 (N_1071,In_168,In_2869);
or U1072 (N_1072,In_550,In_1541);
nor U1073 (N_1073,N_141,N_138);
or U1074 (N_1074,In_304,In_1939);
nor U1075 (N_1075,In_2579,In_953);
nor U1076 (N_1076,In_2210,N_414);
nor U1077 (N_1077,In_1723,N_194);
or U1078 (N_1078,In_2033,N_470);
xnor U1079 (N_1079,In_1321,In_1248);
nand U1080 (N_1080,In_242,In_651);
or U1081 (N_1081,In_1096,In_2536);
xor U1082 (N_1082,In_882,In_2544);
xor U1083 (N_1083,In_1616,In_1558);
nand U1084 (N_1084,In_453,In_915);
xnor U1085 (N_1085,In_1911,In_2660);
nand U1086 (N_1086,N_420,In_2684);
xnor U1087 (N_1087,N_461,N_150);
nor U1088 (N_1088,In_1145,N_161);
nor U1089 (N_1089,In_285,In_2397);
and U1090 (N_1090,In_1184,In_1380);
or U1091 (N_1091,In_1905,In_1001);
xnor U1092 (N_1092,In_2783,In_2977);
nor U1093 (N_1093,In_1937,In_1263);
and U1094 (N_1094,In_983,In_2125);
xnor U1095 (N_1095,In_1876,In_2477);
nand U1096 (N_1096,In_1478,In_94);
and U1097 (N_1097,In_860,N_477);
or U1098 (N_1098,In_2720,In_1763);
and U1099 (N_1099,N_7,In_2573);
nand U1100 (N_1100,In_1896,In_2422);
nor U1101 (N_1101,In_1325,In_64);
xor U1102 (N_1102,In_681,N_319);
nand U1103 (N_1103,N_548,N_415);
xor U1104 (N_1104,In_2524,N_464);
xor U1105 (N_1105,In_2460,In_2803);
nand U1106 (N_1106,In_1472,N_87);
nor U1107 (N_1107,N_257,In_2268);
xnor U1108 (N_1108,In_395,In_594);
xor U1109 (N_1109,In_1828,In_2883);
nand U1110 (N_1110,N_206,In_2923);
nand U1111 (N_1111,In_1537,N_115);
nand U1112 (N_1112,In_271,In_1721);
or U1113 (N_1113,N_132,N_40);
and U1114 (N_1114,N_441,In_641);
or U1115 (N_1115,N_495,In_730);
xor U1116 (N_1116,In_362,N_229);
nor U1117 (N_1117,In_1060,N_103);
nand U1118 (N_1118,N_185,In_1090);
xnor U1119 (N_1119,N_364,In_1359);
xor U1120 (N_1120,N_360,In_2188);
nand U1121 (N_1121,In_728,In_2591);
nand U1122 (N_1122,N_316,In_1354);
xor U1123 (N_1123,N_25,In_1301);
nand U1124 (N_1124,In_2342,N_377);
xor U1125 (N_1125,In_40,In_1360);
and U1126 (N_1126,In_2860,In_484);
or U1127 (N_1127,In_590,In_976);
nand U1128 (N_1128,In_1004,In_744);
nor U1129 (N_1129,In_894,In_2260);
or U1130 (N_1130,In_1506,In_1761);
xor U1131 (N_1131,N_565,In_2498);
and U1132 (N_1132,N_158,N_296);
nand U1133 (N_1133,In_2045,N_262);
nor U1134 (N_1134,N_435,In_292);
nor U1135 (N_1135,In_1913,In_1960);
nor U1136 (N_1136,In_2312,In_833);
xor U1137 (N_1137,In_42,In_1625);
nand U1138 (N_1138,N_342,In_2097);
nand U1139 (N_1139,In_320,In_582);
or U1140 (N_1140,In_426,In_796);
xnor U1141 (N_1141,N_179,In_906);
nor U1142 (N_1142,In_2892,N_547);
nor U1143 (N_1143,In_1959,N_570);
nor U1144 (N_1144,In_2736,N_500);
xor U1145 (N_1145,N_230,In_2111);
nand U1146 (N_1146,N_26,In_1430);
nand U1147 (N_1147,In_1124,In_1672);
and U1148 (N_1148,In_735,In_1168);
or U1149 (N_1149,In_2865,N_89);
nand U1150 (N_1150,In_1690,N_91);
and U1151 (N_1151,In_2946,N_313);
nand U1152 (N_1152,N_355,In_1461);
and U1153 (N_1153,In_84,N_532);
or U1154 (N_1154,In_956,In_996);
nor U1155 (N_1155,In_948,In_118);
xor U1156 (N_1156,N_227,In_355);
xor U1157 (N_1157,In_370,In_162);
or U1158 (N_1158,In_1401,In_1921);
xor U1159 (N_1159,In_758,N_527);
nor U1160 (N_1160,N_339,N_184);
and U1161 (N_1161,N_19,In_2393);
or U1162 (N_1162,N_39,In_2490);
and U1163 (N_1163,In_1685,In_2297);
or U1164 (N_1164,In_1566,In_2686);
xnor U1165 (N_1165,In_964,In_224);
xnor U1166 (N_1166,In_2816,In_1087);
nor U1167 (N_1167,In_2620,In_1863);
nor U1168 (N_1168,In_570,In_24);
nand U1169 (N_1169,In_2390,N_173);
and U1170 (N_1170,In_1606,In_1233);
or U1171 (N_1171,In_41,N_218);
nor U1172 (N_1172,In_1258,In_2672);
xnor U1173 (N_1173,N_462,In_119);
xor U1174 (N_1174,In_919,In_330);
nor U1175 (N_1175,In_2304,N_486);
and U1176 (N_1176,In_2043,N_523);
xor U1177 (N_1177,In_180,In_691);
nand U1178 (N_1178,In_1687,In_1945);
nor U1179 (N_1179,In_1382,In_275);
nor U1180 (N_1180,In_2516,In_1420);
nor U1181 (N_1181,In_1491,N_171);
or U1182 (N_1182,In_1247,In_1303);
nand U1183 (N_1183,N_238,In_1454);
and U1184 (N_1184,In_2491,In_221);
and U1185 (N_1185,In_731,In_1272);
nor U1186 (N_1186,In_1370,N_320);
xnor U1187 (N_1187,In_1651,N_417);
nor U1188 (N_1188,In_2688,In_2762);
nand U1189 (N_1189,N_595,In_276);
and U1190 (N_1190,In_1284,In_173);
or U1191 (N_1191,N_295,N_168);
and U1192 (N_1192,In_2156,In_1877);
xor U1193 (N_1193,In_2616,In_519);
and U1194 (N_1194,In_1146,In_133);
nor U1195 (N_1195,In_1447,In_344);
or U1196 (N_1196,In_2564,In_2171);
and U1197 (N_1197,In_1878,In_2501);
or U1198 (N_1198,In_2375,In_521);
or U1199 (N_1199,N_3,In_154);
xnor U1200 (N_1200,In_576,N_375);
or U1201 (N_1201,N_204,N_1184);
xor U1202 (N_1202,N_1098,In_788);
nor U1203 (N_1203,In_1780,In_1814);
nand U1204 (N_1204,N_616,N_615);
or U1205 (N_1205,In_539,In_2090);
and U1206 (N_1206,In_2300,In_733);
nor U1207 (N_1207,N_1154,N_1094);
nand U1208 (N_1208,N_819,N_707);
or U1209 (N_1209,In_1508,In_1662);
xnor U1210 (N_1210,In_137,N_374);
nor U1211 (N_1211,In_1832,In_2711);
nor U1212 (N_1212,N_975,In_644);
or U1213 (N_1213,N_828,N_1066);
or U1214 (N_1214,N_841,N_948);
nand U1215 (N_1215,N_991,In_1302);
nand U1216 (N_1216,N_992,N_1004);
xnor U1217 (N_1217,N_481,N_869);
and U1218 (N_1218,N_1048,N_528);
nand U1219 (N_1219,In_125,In_1409);
or U1220 (N_1220,In_2897,N_997);
nor U1221 (N_1221,In_1725,In_918);
nor U1222 (N_1222,N_545,N_857);
and U1223 (N_1223,N_946,N_36);
nor U1224 (N_1224,In_2613,N_1021);
and U1225 (N_1225,N_606,In_269);
nand U1226 (N_1226,N_1043,N_977);
xnor U1227 (N_1227,N_799,In_513);
xnor U1228 (N_1228,N_348,N_466);
and U1229 (N_1229,N_280,In_1622);
xor U1230 (N_1230,N_733,In_1727);
or U1231 (N_1231,In_1078,In_545);
nand U1232 (N_1232,In_2833,N_785);
or U1233 (N_1233,In_2680,In_1278);
xnor U1234 (N_1234,In_2683,In_1425);
nor U1235 (N_1235,N_276,N_628);
nor U1236 (N_1236,N_506,N_424);
xor U1237 (N_1237,N_865,N_1034);
nand U1238 (N_1238,In_599,In_844);
nand U1239 (N_1239,In_316,In_791);
xnor U1240 (N_1240,N_634,N_90);
or U1241 (N_1241,In_318,In_1890);
xnor U1242 (N_1242,In_683,N_202);
or U1243 (N_1243,N_118,In_837);
xnor U1244 (N_1244,N_772,N_766);
or U1245 (N_1245,In_121,N_837);
and U1246 (N_1246,In_1292,In_1503);
xor U1247 (N_1247,N_1166,N_632);
or U1248 (N_1248,N_357,In_646);
or U1249 (N_1249,In_1970,N_784);
or U1250 (N_1250,In_900,In_321);
nor U1251 (N_1251,N_1168,N_847);
nand U1252 (N_1252,N_662,In_1714);
nand U1253 (N_1253,In_697,In_950);
xnor U1254 (N_1254,In_2051,In_1629);
nand U1255 (N_1255,In_1334,In_1059);
or U1256 (N_1256,In_2882,N_700);
xnor U1257 (N_1257,In_2904,N_1101);
nand U1258 (N_1258,In_150,In_538);
nor U1259 (N_1259,In_324,N_559);
and U1260 (N_1260,N_473,N_777);
nor U1261 (N_1261,N_1093,N_829);
nor U1262 (N_1262,In_1812,In_1034);
or U1263 (N_1263,N_982,N_878);
xor U1264 (N_1264,In_1028,N_734);
nor U1265 (N_1265,N_543,In_2109);
nor U1266 (N_1266,In_779,In_1564);
nor U1267 (N_1267,In_2752,N_131);
and U1268 (N_1268,N_1148,N_618);
nor U1269 (N_1269,In_2916,In_491);
and U1270 (N_1270,N_1061,In_2369);
nand U1271 (N_1271,N_608,In_717);
or U1272 (N_1272,In_1628,N_338);
xor U1273 (N_1273,N_969,N_494);
or U1274 (N_1274,In_1906,In_656);
and U1275 (N_1275,In_2515,N_67);
xor U1276 (N_1276,In_1882,N_556);
nand U1277 (N_1277,In_26,N_538);
xnor U1278 (N_1278,In_2611,In_2928);
xor U1279 (N_1279,In_1505,In_2052);
or U1280 (N_1280,In_2175,In_300);
xnor U1281 (N_1281,N_673,N_688);
and U1282 (N_1282,In_1976,In_2519);
xor U1283 (N_1283,In_1385,N_771);
nand U1284 (N_1284,N_791,In_237);
nand U1285 (N_1285,In_1133,In_1187);
and U1286 (N_1286,N_1180,N_925);
nor U1287 (N_1287,In_904,In_1205);
or U1288 (N_1288,N_487,N_213);
xnor U1289 (N_1289,N_1144,N_795);
nor U1290 (N_1290,In_564,N_679);
nand U1291 (N_1291,In_1720,In_622);
xnor U1292 (N_1292,N_586,N_642);
and U1293 (N_1293,N_330,In_2019);
or U1294 (N_1294,N_613,In_1645);
or U1295 (N_1295,In_647,N_560);
nand U1296 (N_1296,N_620,In_1898);
or U1297 (N_1297,In_1468,In_2739);
and U1298 (N_1298,In_1137,N_1133);
or U1299 (N_1299,N_718,In_2899);
or U1300 (N_1300,In_2577,N_268);
nor U1301 (N_1301,N_451,N_986);
xnor U1302 (N_1302,N_14,In_745);
and U1303 (N_1303,N_1018,In_2550);
and U1304 (N_1304,N_1007,N_1189);
xnor U1305 (N_1305,N_933,In_1032);
xor U1306 (N_1306,In_113,N_601);
and U1307 (N_1307,In_2914,In_2054);
or U1308 (N_1308,N_990,In_463);
and U1309 (N_1309,In_781,N_69);
nand U1310 (N_1310,N_219,N_1125);
and U1311 (N_1311,N_697,In_785);
or U1312 (N_1312,In_2950,In_2985);
nand U1313 (N_1313,N_1197,In_2211);
xor U1314 (N_1314,In_461,N_580);
xnor U1315 (N_1315,N_33,N_465);
nand U1316 (N_1316,N_1049,In_2413);
xnor U1317 (N_1317,In_944,N_344);
nor U1318 (N_1318,N_896,N_796);
nor U1319 (N_1319,N_1027,In_771);
or U1320 (N_1320,N_1062,N_874);
nor U1321 (N_1321,N_351,N_830);
nand U1322 (N_1322,In_2226,N_237);
xnor U1323 (N_1323,N_460,N_1025);
nor U1324 (N_1324,In_2625,In_1413);
nor U1325 (N_1325,N_1117,N_1091);
xor U1326 (N_1326,In_1019,N_629);
xnor U1327 (N_1327,In_1677,In_2507);
and U1328 (N_1328,In_2908,N_1047);
nand U1329 (N_1329,N_1112,In_2810);
nor U1330 (N_1330,In_503,In_810);
and U1331 (N_1331,In_2131,N_960);
or U1332 (N_1332,In_1182,In_1173);
or U1333 (N_1333,N_645,In_569);
xnor U1334 (N_1334,In_766,N_996);
and U1335 (N_1335,N_1083,N_906);
nor U1336 (N_1336,N_576,In_2834);
xnor U1337 (N_1337,In_913,N_1116);
nand U1338 (N_1338,N_1063,In_715);
xor U1339 (N_1339,N_940,N_643);
or U1340 (N_1340,N_1033,In_1091);
nand U1341 (N_1341,N_1128,In_387);
or U1342 (N_1342,In_327,N_1028);
nand U1343 (N_1343,N_603,N_911);
or U1344 (N_1344,N_1196,In_529);
nand U1345 (N_1345,In_591,In_2199);
nand U1346 (N_1346,In_1652,In_2585);
xor U1347 (N_1347,N_806,N_1181);
nor U1348 (N_1348,In_973,In_2644);
nor U1349 (N_1349,In_2823,In_310);
nor U1350 (N_1350,In_2176,N_515);
nor U1351 (N_1351,In_2906,N_1163);
or U1352 (N_1352,N_749,N_277);
or U1353 (N_1353,In_530,N_169);
nor U1354 (N_1354,In_429,In_2265);
nor U1355 (N_1355,N_722,N_716);
nor U1356 (N_1356,In_2980,N_24);
nand U1357 (N_1357,N_463,N_926);
xor U1358 (N_1358,In_2328,In_2012);
nor U1359 (N_1359,In_581,N_478);
nand U1360 (N_1360,In_332,N_188);
nand U1361 (N_1361,N_1080,N_687);
or U1362 (N_1362,N_621,In_1340);
or U1363 (N_1363,In_2197,In_2003);
or U1364 (N_1364,N_903,N_957);
xnor U1365 (N_1365,In_2398,N_959);
xnor U1366 (N_1366,In_1316,In_2624);
and U1367 (N_1367,N_1055,In_1734);
and U1368 (N_1368,In_2565,In_2984);
xnor U1369 (N_1369,N_921,In_1005);
or U1370 (N_1370,In_2986,N_901);
nor U1371 (N_1371,In_807,In_2500);
nor U1372 (N_1372,In_797,In_2428);
nand U1373 (N_1373,In_1891,N_637);
nand U1374 (N_1374,In_1132,In_444);
nand U1375 (N_1375,N_225,In_385);
nand U1376 (N_1376,N_78,In_2776);
nor U1377 (N_1377,N_430,In_1070);
nor U1378 (N_1378,N_468,N_843);
xnor U1379 (N_1379,N_713,In_1515);
xor U1380 (N_1380,N_517,In_1648);
and U1381 (N_1381,In_1600,In_2842);
or U1382 (N_1382,In_12,In_1269);
and U1383 (N_1383,In_1864,N_488);
xnor U1384 (N_1384,In_1917,In_2742);
nor U1385 (N_1385,In_1701,N_699);
xnor U1386 (N_1386,In_922,N_952);
nand U1387 (N_1387,In_889,In_2193);
nand U1388 (N_1388,In_2182,N_431);
and U1389 (N_1389,N_447,In_1398);
xor U1390 (N_1390,N_783,In_1274);
or U1391 (N_1391,In_348,In_152);
and U1392 (N_1392,N_383,In_384);
nand U1393 (N_1393,N_526,N_861);
xnor U1394 (N_1394,N_9,N_321);
nor U1395 (N_1395,In_1933,N_706);
xnor U1396 (N_1396,In_1977,N_963);
nand U1397 (N_1397,In_596,In_2761);
xor U1398 (N_1398,In_2508,In_2166);
xor U1399 (N_1399,In_1638,In_1442);
and U1400 (N_1400,In_874,In_2506);
xnor U1401 (N_1401,N_445,In_1982);
or U1402 (N_1402,N_271,N_484);
nor U1403 (N_1403,N_1,N_988);
or U1404 (N_1404,In_1395,N_972);
or U1405 (N_1405,In_1225,In_2352);
and U1406 (N_1406,N_391,N_1135);
and U1407 (N_1407,N_197,In_1355);
and U1408 (N_1408,In_1056,In_402);
nor U1409 (N_1409,N_597,In_2793);
and U1410 (N_1410,N_553,In_2952);
or U1411 (N_1411,N_851,In_2785);
and U1412 (N_1412,N_899,N_683);
nor U1413 (N_1413,N_593,N_647);
or U1414 (N_1414,N_113,N_924);
and U1415 (N_1415,N_1178,N_867);
or U1416 (N_1416,N_702,N_654);
and U1417 (N_1417,N_1143,N_732);
or U1418 (N_1418,In_417,In_75);
nor U1419 (N_1419,In_2747,In_1103);
or U1420 (N_1420,N_909,N_498);
xor U1421 (N_1421,In_2504,In_1925);
or U1422 (N_1422,In_159,N_979);
and U1423 (N_1423,In_1465,N_1113);
nor U1424 (N_1424,N_757,N_530);
or U1425 (N_1425,N_1079,N_846);
and U1426 (N_1426,N_1059,N_1190);
and U1427 (N_1427,In_2778,N_1167);
or U1428 (N_1428,In_1914,In_2493);
xor U1429 (N_1429,In_616,In_1064);
or U1430 (N_1430,In_274,N_516);
nand U1431 (N_1431,In_401,N_882);
nor U1432 (N_1432,In_2112,N_804);
nor U1433 (N_1433,N_279,N_842);
and U1434 (N_1434,N_522,In_2781);
nor U1435 (N_1435,In_841,In_1743);
and U1436 (N_1436,N_34,In_1872);
nand U1437 (N_1437,In_2789,N_1198);
nand U1438 (N_1438,N_684,In_404);
nand U1439 (N_1439,In_1259,N_29);
xor U1440 (N_1440,In_2790,N_1058);
or U1441 (N_1441,In_2879,In_1109);
xor U1442 (N_1442,N_1022,In_2186);
xnor U1443 (N_1443,N_939,In_469);
xor U1444 (N_1444,In_949,In_30);
nor U1445 (N_1445,In_943,N_976);
and U1446 (N_1446,N_935,N_1032);
and U1447 (N_1447,N_1065,N_410);
and U1448 (N_1448,In_2223,N_755);
and U1449 (N_1449,In_2307,N_1089);
xor U1450 (N_1450,N_1035,In_110);
and U1451 (N_1451,In_2178,N_166);
nand U1452 (N_1452,In_608,In_1131);
and U1453 (N_1453,N_1124,In_1636);
or U1454 (N_1454,In_1423,N_1132);
xnor U1455 (N_1455,N_1029,In_2963);
xor U1456 (N_1456,N_696,N_336);
and U1457 (N_1457,N_1044,In_5);
xnor U1458 (N_1458,In_183,N_1171);
and U1459 (N_1459,In_354,N_326);
nor U1460 (N_1460,In_1488,N_433);
nor U1461 (N_1461,N_1077,In_2671);
and U1462 (N_1462,In_787,N_917);
nor U1463 (N_1463,In_1427,In_1332);
nor U1464 (N_1464,N_1123,N_886);
or U1465 (N_1465,In_433,N_665);
nand U1466 (N_1466,In_1675,In_103);
or U1467 (N_1467,In_1803,In_2836);
xnor U1468 (N_1468,N_879,In_2344);
nor U1469 (N_1469,N_121,N_822);
xor U1470 (N_1470,N_254,N_738);
xor U1471 (N_1471,N_1090,N_1075);
nor U1472 (N_1472,N_1120,In_2502);
or U1473 (N_1473,In_428,In_559);
and U1474 (N_1474,In_2699,N_1191);
and U1475 (N_1475,N_1160,N_125);
nand U1476 (N_1476,In_1689,N_503);
and U1477 (N_1477,In_1159,N_720);
nand U1478 (N_1478,N_607,N_222);
and U1479 (N_1479,N_1102,In_1483);
or U1480 (N_1480,In_1966,In_1885);
nand U1481 (N_1481,N_1060,In_16);
or U1482 (N_1482,In_2073,N_1070);
and U1483 (N_1483,N_754,N_686);
nand U1484 (N_1484,N_192,N_1140);
or U1485 (N_1485,In_1543,N_998);
and U1486 (N_1486,N_630,N_659);
nor U1487 (N_1487,N_329,In_1713);
nand U1488 (N_1488,In_593,N_936);
nand U1489 (N_1489,In_2703,In_2901);
nor U1490 (N_1490,N_648,In_1201);
xor U1491 (N_1491,In_71,N_1186);
and U1492 (N_1492,N_1096,N_915);
and U1493 (N_1493,In_2165,N_743);
nor U1494 (N_1494,N_402,N_452);
and U1495 (N_1495,N_912,N_989);
xnor U1496 (N_1496,N_511,In_991);
nor U1497 (N_1497,N_1082,In_1892);
or U1498 (N_1498,In_167,N_1012);
or U1499 (N_1499,In_345,In_1067);
nand U1500 (N_1500,N_564,In_377);
and U1501 (N_1501,N_244,N_1152);
and U1502 (N_1502,N_521,In_2316);
xor U1503 (N_1503,N_221,N_807);
or U1504 (N_1504,In_302,N_877);
and U1505 (N_1505,In_1181,N_938);
or U1506 (N_1506,N_315,N_769);
nand U1507 (N_1507,N_762,In_67);
and U1508 (N_1508,In_859,N_1172);
and U1509 (N_1509,In_1513,N_868);
or U1510 (N_1510,In_1416,N_1000);
nand U1511 (N_1511,N_729,In_371);
nand U1512 (N_1512,In_1999,In_2697);
or U1513 (N_1513,In_2299,In_2362);
and U1514 (N_1514,In_72,In_122);
nor U1515 (N_1515,In_2529,In_2741);
nand U1516 (N_1516,N_1176,N_143);
or U1517 (N_1517,N_1106,N_1005);
and U1518 (N_1518,N_209,N_1159);
xor U1519 (N_1519,N_1037,N_892);
nand U1520 (N_1520,N_554,In_813);
nand U1521 (N_1521,In_2719,N_1014);
and U1522 (N_1522,N_589,In_2594);
nand U1523 (N_1523,N_612,N_765);
xnor U1524 (N_1524,In_1974,N_561);
nor U1525 (N_1525,N_930,N_922);
or U1526 (N_1526,N_1174,In_1012);
nor U1527 (N_1527,In_2313,In_2459);
nand U1528 (N_1528,In_725,In_2692);
and U1529 (N_1529,In_510,N_459);
nor U1530 (N_1530,In_2844,N_394);
nand U1531 (N_1531,In_2330,In_258);
or U1532 (N_1532,In_1317,In_90);
nor U1533 (N_1533,In_2303,N_73);
and U1534 (N_1534,In_970,N_779);
or U1535 (N_1535,N_885,In_440);
or U1536 (N_1536,In_456,In_2517);
nand U1537 (N_1537,N_967,N_274);
or U1538 (N_1538,N_134,In_1845);
nor U1539 (N_1539,N_639,In_603);
xor U1540 (N_1540,N_790,In_940);
nand U1541 (N_1541,N_1187,N_1131);
xnor U1542 (N_1542,In_1655,In_2845);
and U1543 (N_1543,In_2549,N_1074);
nand U1544 (N_1544,N_361,N_859);
nor U1545 (N_1545,N_436,In_1731);
xnor U1546 (N_1546,N_476,N_814);
xnor U1547 (N_1547,N_228,In_2001);
nor U1548 (N_1548,In_883,N_1177);
and U1549 (N_1549,In_2526,In_2559);
nand U1550 (N_1550,In_82,In_172);
or U1551 (N_1551,In_380,N_705);
nand U1552 (N_1552,In_2521,In_2414);
nor U1553 (N_1553,In_2915,N_965);
nand U1554 (N_1554,In_2893,N_537);
or U1555 (N_1555,In_1893,In_621);
xnor U1556 (N_1556,In_1022,In_1532);
and U1557 (N_1557,In_2858,N_727);
and U1558 (N_1558,N_780,In_1189);
or U1559 (N_1559,N_47,N_721);
xor U1560 (N_1560,N_735,In_2920);
nor U1561 (N_1561,N_1016,N_529);
nand U1562 (N_1562,In_1250,In_869);
nor U1563 (N_1563,N_692,N_895);
or U1564 (N_1564,In_1120,N_1121);
nand U1565 (N_1565,In_2835,N_1017);
nand U1566 (N_1566,N_482,N_1137);
and U1567 (N_1567,N_193,In_1476);
xor U1568 (N_1568,In_2825,N_327);
and U1569 (N_1569,N_504,N_314);
xnor U1570 (N_1570,N_943,N_251);
nand U1571 (N_1571,In_1372,In_1660);
nor U1572 (N_1572,N_492,In_2421);
xnor U1573 (N_1573,N_1150,In_1627);
nand U1574 (N_1574,In_789,In_1176);
xor U1575 (N_1575,N_962,N_920);
nand U1576 (N_1576,N_584,In_2829);
xor U1577 (N_1577,In_978,In_393);
nand U1578 (N_1578,In_2987,N_698);
nand U1579 (N_1579,N_778,In_1550);
and U1580 (N_1580,N_704,N_782);
xnor U1581 (N_1581,In_2000,In_1781);
nand U1582 (N_1582,In_2715,In_2900);
nand U1583 (N_1583,In_1496,N_130);
xnor U1584 (N_1584,N_880,In_2689);
and U1585 (N_1585,In_2567,N_539);
xnor U1586 (N_1586,In_334,N_442);
xnor U1587 (N_1587,In_1764,N_968);
and U1588 (N_1588,In_313,N_1175);
and U1589 (N_1589,N_871,In_1549);
or U1590 (N_1590,In_2596,In_2732);
nand U1591 (N_1591,N_1085,In_1705);
nand U1592 (N_1592,In_2870,N_626);
or U1593 (N_1593,N_753,In_1281);
and U1594 (N_1594,N_1046,In_602);
nor U1595 (N_1595,N_1109,N_739);
and U1596 (N_1596,N_839,N_305);
and U1597 (N_1597,N_0,In_535);
or U1598 (N_1598,In_4,In_2622);
or U1599 (N_1599,In_358,In_689);
nor U1600 (N_1600,N_817,In_714);
nor U1601 (N_1601,In_2822,In_2065);
and U1602 (N_1602,N_1192,In_2880);
and U1603 (N_1603,N_311,N_81);
and U1604 (N_1604,N_1179,N_736);
or U1605 (N_1605,In_1195,In_148);
or U1606 (N_1606,N_1024,N_525);
nand U1607 (N_1607,In_1538,In_2828);
or U1608 (N_1608,N_866,N_950);
nand U1609 (N_1609,N_695,N_602);
nor U1610 (N_1610,N_764,N_283);
nand U1611 (N_1611,In_39,N_1087);
nand U1612 (N_1612,N_818,N_958);
xor U1613 (N_1613,In_1699,In_2523);
or U1614 (N_1614,In_2449,In_2627);
nand U1615 (N_1615,N_54,In_2034);
nor U1616 (N_1616,N_864,In_592);
xor U1617 (N_1617,N_905,N_900);
nor U1618 (N_1618,In_580,N_291);
nand U1619 (N_1619,N_638,In_1719);
nor U1620 (N_1620,In_273,In_204);
or U1621 (N_1621,N_1169,N_63);
xor U1622 (N_1622,N_1084,N_332);
or U1623 (N_1623,N_984,In_1439);
nand U1624 (N_1624,In_1485,N_650);
or U1625 (N_1625,N_434,N_77);
nand U1626 (N_1626,N_703,In_1686);
nand U1627 (N_1627,In_1122,In_476);
nor U1628 (N_1628,N_675,N_849);
nand U1629 (N_1629,N_30,N_835);
nand U1630 (N_1630,In_372,N_761);
nand U1631 (N_1631,In_2011,In_924);
and U1632 (N_1632,N_758,N_947);
nor U1633 (N_1633,N_397,In_2322);
xnor U1634 (N_1634,N_1155,N_1103);
or U1635 (N_1635,In_548,In_2337);
or U1636 (N_1636,In_587,N_163);
nor U1637 (N_1637,In_637,In_557);
nor U1638 (N_1638,N_694,In_415);
xor U1639 (N_1639,N_928,N_763);
nor U1640 (N_1640,In_2029,N_746);
nor U1641 (N_1641,In_9,N_824);
nor U1642 (N_1642,In_1421,In_1610);
and U1643 (N_1643,In_53,In_1665);
and U1644 (N_1644,N_862,In_2096);
nand U1645 (N_1645,N_388,N_1134);
xor U1646 (N_1646,In_790,In_218);
nand U1647 (N_1647,In_2263,In_908);
or U1648 (N_1648,In_2643,In_1324);
and U1649 (N_1649,In_2081,In_2907);
nor U1650 (N_1650,N_1013,N_951);
xor U1651 (N_1651,N_652,N_747);
or U1652 (N_1652,In_1846,N_44);
nor U1653 (N_1653,In_2527,In_2021);
xnor U1654 (N_1654,In_1239,N_624);
and U1655 (N_1655,In_1897,N_737);
nor U1656 (N_1656,In_1683,N_496);
and U1657 (N_1657,In_1745,In_2872);
or U1658 (N_1658,In_1698,N_1069);
nand U1659 (N_1659,In_1191,In_1300);
or U1660 (N_1660,N_1141,In_2233);
xor U1661 (N_1661,N_399,In_2853);
xnor U1662 (N_1662,N_440,N_1145);
or U1663 (N_1663,N_760,In_99);
nor U1664 (N_1664,N_955,In_2499);
or U1665 (N_1665,In_2772,In_439);
or U1666 (N_1666,N_821,In_1837);
xnor U1667 (N_1667,In_2586,In_437);
and U1668 (N_1668,In_762,N_929);
or U1669 (N_1669,N_793,N_292);
or U1670 (N_1670,N_421,N_927);
xor U1671 (N_1671,N_577,In_1407);
xor U1672 (N_1672,N_808,In_2592);
or U1673 (N_1673,In_487,N_1139);
or U1674 (N_1674,In_1585,N_1162);
xor U1675 (N_1675,In_2510,N_367);
nor U1676 (N_1676,N_1118,In_806);
and U1677 (N_1677,N_672,N_775);
and U1678 (N_1678,N_1040,In_1033);
and U1679 (N_1679,In_1117,N_981);
or U1680 (N_1680,In_2070,In_312);
nor U1681 (N_1681,N_625,N_263);
xor U1682 (N_1682,N_681,In_413);
xor U1683 (N_1683,N_428,N_518);
or U1684 (N_1684,N_207,In_962);
xor U1685 (N_1685,N_60,N_365);
or U1686 (N_1686,In_1676,N_350);
or U1687 (N_1687,N_1095,N_913);
and U1688 (N_1688,N_308,In_2443);
xnor U1689 (N_1689,In_1270,In_309);
and U1690 (N_1690,N_557,In_1384);
xor U1691 (N_1691,N_1071,N_250);
xor U1692 (N_1692,In_2283,N_711);
or U1693 (N_1693,In_611,N_536);
nand U1694 (N_1694,In_1411,N_1003);
and U1695 (N_1695,In_398,N_971);
nand U1696 (N_1696,N_827,In_2246);
or U1697 (N_1697,N_825,In_1172);
nor U1698 (N_1698,In_1587,N_1182);
nand U1699 (N_1699,N_1076,In_1026);
and U1700 (N_1700,In_219,N_823);
nor U1701 (N_1701,N_728,N_51);
and U1702 (N_1702,In_1043,In_2254);
xnor U1703 (N_1703,In_633,N_405);
nand U1704 (N_1704,N_888,In_1268);
nor U1705 (N_1705,In_2650,N_619);
and U1706 (N_1706,N_1183,In_2142);
xnor U1707 (N_1707,In_2733,In_2333);
and U1708 (N_1708,N_741,N_614);
or U1709 (N_1709,In_2069,N_1136);
and U1710 (N_1710,In_1104,N_715);
and U1711 (N_1711,In_1313,N_970);
nor U1712 (N_1712,In_2572,N_1149);
and U1713 (N_1713,In_993,In_2925);
and U1714 (N_1714,In_1153,In_1750);
and U1715 (N_1715,In_1171,N_883);
and U1716 (N_1716,N_691,In_2532);
and U1717 (N_1717,N_891,In_2942);
nand U1718 (N_1718,In_2191,In_890);
nand U1719 (N_1719,In_2261,In_246);
nor U1720 (N_1720,In_342,In_2379);
xnor U1721 (N_1721,N_386,In_2400);
nand U1722 (N_1722,N_62,In_1586);
or U1723 (N_1723,In_317,N_714);
xnor U1724 (N_1724,N_562,N_444);
or U1725 (N_1725,N_910,N_1073);
or U1726 (N_1726,N_569,In_157);
nor U1727 (N_1727,N_1002,In_2528);
or U1728 (N_1728,In_2439,N_1099);
nand U1729 (N_1729,In_1194,In_1363);
nand U1730 (N_1730,N_812,In_2201);
or U1731 (N_1731,N_742,N_139);
or U1732 (N_1732,In_2830,N_144);
nand U1733 (N_1733,In_1618,In_303);
or U1734 (N_1734,In_338,In_2881);
and U1735 (N_1735,In_245,N_20);
and U1736 (N_1736,N_31,In_1804);
or U1737 (N_1737,N_505,In_669);
or U1738 (N_1738,In_2291,In_382);
nand U1739 (N_1739,In_1368,In_1632);
or U1740 (N_1740,In_1016,In_2071);
and U1741 (N_1741,In_1265,N_396);
and U1742 (N_1742,In_1144,In_734);
nand U1743 (N_1743,In_2760,In_326);
nor U1744 (N_1744,In_1183,In_473);
and U1745 (N_1745,In_1234,In_1165);
xor U1746 (N_1746,N_651,N_767);
xor U1747 (N_1747,N_176,N_1015);
and U1748 (N_1748,N_798,N_644);
nor U1749 (N_1749,N_372,N_1010);
nand U1750 (N_1750,In_2077,N_281);
and U1751 (N_1751,N_949,In_989);
nand U1752 (N_1752,N_641,In_526);
xnor U1753 (N_1753,In_1931,N_1067);
or U1754 (N_1754,In_373,N_493);
or U1755 (N_1755,N_811,N_1068);
nand U1756 (N_1756,In_1932,In_760);
nand U1757 (N_1757,In_865,N_284);
or U1758 (N_1758,In_1567,In_170);
or U1759 (N_1759,N_1119,N_708);
or U1760 (N_1760,In_638,In_1957);
nand U1761 (N_1761,In_1192,N_306);
nand U1762 (N_1762,N_792,N_956);
nand U1763 (N_1763,N_750,N_994);
and U1764 (N_1764,In_98,In_687);
nor U1765 (N_1765,In_163,N_200);
nor U1766 (N_1766,N_600,N_640);
nor U1767 (N_1767,N_1104,In_2497);
nor U1768 (N_1768,In_885,In_241);
and U1769 (N_1769,In_2800,In_62);
nand U1770 (N_1770,In_1178,In_1024);
nor U1771 (N_1771,In_431,In_412);
or U1772 (N_1772,In_2944,In_690);
nor U1773 (N_1773,N_497,In_1044);
nor U1774 (N_1774,In_1573,In_2973);
nand U1775 (N_1775,In_1667,In_615);
nor U1776 (N_1776,In_2503,N_1056);
or U1777 (N_1777,In_2722,In_2943);
xnor U1778 (N_1778,N_571,N_581);
xor U1779 (N_1779,N_983,N_1185);
nor U1780 (N_1780,In_2075,In_2905);
nand U1781 (N_1781,In_1071,N_400);
xor U1782 (N_1782,In_937,In_2152);
and U1783 (N_1783,N_1001,N_631);
or U1784 (N_1784,N_203,In_1511);
nand U1785 (N_1785,In_254,N_1052);
nor U1786 (N_1786,In_1710,In_1470);
nand U1787 (N_1787,In_2039,In_2338);
nor U1788 (N_1788,N_893,N_38);
or U1789 (N_1789,In_664,N_802);
or U1790 (N_1790,N_788,N_786);
xnor U1791 (N_1791,In_2194,In_818);
and U1792 (N_1792,N_916,N_1042);
xnor U1793 (N_1793,In_175,In_1633);
xor U1794 (N_1794,N_717,N_1110);
nand U1795 (N_1795,In_2909,In_2023);
nor U1796 (N_1796,In_1246,In_862);
nand U1797 (N_1797,In_2177,N_489);
nand U1798 (N_1798,N_366,In_2941);
xor U1799 (N_1799,In_1445,In_361);
nand U1800 (N_1800,N_774,N_1345);
or U1801 (N_1801,In_325,N_1211);
or U1802 (N_1802,In_1730,N_61);
nand U1803 (N_1803,N_934,N_347);
or U1804 (N_1804,In_2408,N_1655);
nand U1805 (N_1805,N_1746,N_810);
xor U1806 (N_1806,In_2285,N_406);
and U1807 (N_1807,N_1357,In_2884);
or U1808 (N_1808,N_1796,In_1840);
nand U1809 (N_1809,N_1464,N_1497);
and U1810 (N_1810,In_2740,N_1740);
xor U1811 (N_1811,N_1449,In_425);
and U1812 (N_1812,N_1686,N_1698);
and U1813 (N_1813,In_1534,In_1924);
nor U1814 (N_1814,N_964,N_768);
and U1815 (N_1815,N_1794,N_897);
and U1816 (N_1816,N_1513,N_1335);
xor U1817 (N_1817,N_781,N_1658);
nor U1818 (N_1818,N_838,In_2910);
nor U1819 (N_1819,In_2074,N_1036);
and U1820 (N_1820,N_1313,N_1712);
nor U1821 (N_1821,N_1210,N_1276);
nand U1822 (N_1822,N_432,In_1554);
xor U1823 (N_1823,N_1485,N_1151);
xor U1824 (N_1824,N_341,N_1402);
and U1825 (N_1825,In_1252,N_856);
nor U1826 (N_1826,In_945,N_167);
xnor U1827 (N_1827,In_138,N_599);
nor U1828 (N_1828,N_1347,N_1153);
or U1829 (N_1829,N_1528,In_1951);
nand U1830 (N_1830,N_195,N_1667);
or U1831 (N_1831,N_1405,N_1605);
xnor U1832 (N_1832,In_2214,In_139);
nand U1833 (N_1833,N_1165,N_1598);
nor U1834 (N_1834,In_1352,N_1298);
or U1835 (N_1835,In_2955,N_1235);
nor U1836 (N_1836,In_2936,In_1930);
or U1837 (N_1837,N_1483,N_797);
or U1838 (N_1838,In_1978,In_514);
nand U1839 (N_1839,In_2078,N_1576);
or U1840 (N_1840,N_1506,N_1566);
nor U1841 (N_1841,N_1250,In_1670);
nor U1842 (N_1842,N_1487,N_499);
nand U1843 (N_1843,N_172,N_1224);
nand U1844 (N_1844,N_1450,N_605);
or U1845 (N_1845,N_148,N_1239);
nor U1846 (N_1846,N_10,N_776);
and U1847 (N_1847,N_1535,N_1736);
nand U1848 (N_1848,N_1249,N_1525);
nand U1849 (N_1849,In_1520,N_685);
nor U1850 (N_1850,N_1316,N_1423);
and U1851 (N_1851,N_246,N_1504);
nand U1852 (N_1852,N_1651,In_1236);
nand U1853 (N_1853,N_1762,N_1045);
nand U1854 (N_1854,In_1644,N_147);
nand U1855 (N_1855,N_1759,N_999);
or U1856 (N_1856,N_1256,N_731);
and U1857 (N_1857,N_937,N_1554);
or U1858 (N_1858,N_1469,N_1439);
or U1859 (N_1859,N_1649,N_1719);
and U1860 (N_1860,N_1390,N_1318);
nand U1861 (N_1861,N_1718,N_146);
nand U1862 (N_1862,N_875,N_1374);
xor U1863 (N_1863,In_774,N_636);
and U1864 (N_1864,N_1616,N_1523);
xor U1865 (N_1865,In_341,N_124);
xor U1866 (N_1866,N_1766,N_858);
nand U1867 (N_1867,In_1865,N_1730);
nor U1868 (N_1868,N_1367,N_1650);
and U1869 (N_1869,N_604,In_1577);
nand U1870 (N_1870,N_1635,N_1403);
xor U1871 (N_1871,In_1871,N_1427);
nor U1872 (N_1872,In_2605,N_443);
nand U1873 (N_1873,N_1733,In_1658);
nor U1874 (N_1874,N_1257,N_1491);
xnor U1875 (N_1875,In_1226,In_2384);
xor U1876 (N_1876,N_1670,N_1366);
and U1877 (N_1877,N_1767,N_1088);
xnor U1878 (N_1878,N_800,N_1568);
or U1879 (N_1879,N_1587,N_1446);
nor U1880 (N_1880,In_1085,N_1509);
xnor U1881 (N_1881,N_1280,N_1575);
and U1882 (N_1882,N_1314,N_189);
and U1883 (N_1883,N_1320,In_505);
or U1884 (N_1884,N_1678,N_1115);
xor U1885 (N_1885,N_224,N_980);
nand U1886 (N_1886,In_2873,N_1344);
xnor U1887 (N_1887,N_1285,In_1572);
nor U1888 (N_1888,N_853,In_1948);
nor U1889 (N_1889,N_1507,N_1748);
or U1890 (N_1890,N_745,In_1987);
and U1891 (N_1891,N_1674,N_1753);
and U1892 (N_1892,In_1329,N_1632);
nor U1893 (N_1893,In_2076,N_1758);
and U1894 (N_1894,In_968,In_1894);
nor U1895 (N_1895,N_1663,N_833);
nor U1896 (N_1896,In_2386,In_1036);
nor U1897 (N_1897,N_1422,N_1309);
nand U1898 (N_1898,N_751,N_805);
or U1899 (N_1899,In_2159,N_1613);
nand U1900 (N_1900,N_1623,In_1429);
and U1901 (N_1901,N_1567,N_908);
nor U1902 (N_1902,In_1770,N_1786);
and U1903 (N_1903,N_1519,N_109);
and U1904 (N_1904,In_1547,N_832);
xor U1905 (N_1905,In_2228,N_1466);
nand U1906 (N_1906,N_1785,N_1039);
xor U1907 (N_1907,N_966,N_76);
nand U1908 (N_1908,In_2170,N_944);
nand U1909 (N_1909,N_1330,N_1275);
nor U1910 (N_1910,N_1679,N_1307);
and U1911 (N_1911,N_1333,In_1174);
xor U1912 (N_1912,In_101,N_1735);
or U1913 (N_1913,N_1370,N_1768);
or U1914 (N_1914,N_787,In_1581);
nand U1915 (N_1915,In_1356,N_666);
nor U1916 (N_1916,N_1092,N_1326);
and U1917 (N_1917,In_2587,N_1626);
nor U1918 (N_1918,N_587,N_1726);
nand U1919 (N_1919,N_1463,In_435);
nor U1920 (N_1920,N_1300,N_1493);
or U1921 (N_1921,In_583,In_2885);
nor U1922 (N_1922,In_2469,In_2399);
or U1923 (N_1923,N_1409,N_1362);
and U1924 (N_1924,N_1361,In_2314);
or U1925 (N_1925,N_1421,N_730);
nand U1926 (N_1926,N_1299,In_711);
and U1927 (N_1927,N_1452,N_1011);
or U1928 (N_1928,In_191,N_657);
and U1929 (N_1929,N_1435,N_863);
and U1930 (N_1930,N_1516,N_1225);
nand U1931 (N_1931,In_1881,N_724);
nor U1932 (N_1932,In_2121,N_1205);
xor U1933 (N_1933,In_278,N_1627);
and U1934 (N_1934,N_1228,N_1688);
xnor U1935 (N_1935,N_649,N_1383);
or U1936 (N_1936,In_2115,N_1400);
or U1937 (N_1937,In_135,In_1943);
or U1938 (N_1938,N_1207,N_1350);
or U1939 (N_1939,N_1247,N_1661);
nand U1940 (N_1940,N_1732,N_1558);
nand U1941 (N_1941,In_143,N_1780);
nand U1942 (N_1942,N_1301,N_726);
xnor U1943 (N_1943,N_1170,In_2085);
nor U1944 (N_1944,N_719,N_1694);
or U1945 (N_1945,In_1507,N_1395);
nor U1946 (N_1946,N_1653,N_1274);
nor U1947 (N_1947,N_1772,N_1206);
nand U1948 (N_1948,N_1244,N_1440);
xor U1949 (N_1949,In_2145,In_836);
or U1950 (N_1950,N_744,N_1792);
or U1951 (N_1951,In_1105,N_1706);
nand U1952 (N_1952,In_252,In_61);
nand U1953 (N_1953,N_1521,N_1763);
and U1954 (N_1954,N_1492,N_1157);
xnor U1955 (N_1955,N_1524,N_661);
nor U1956 (N_1956,N_1020,In_934);
or U1957 (N_1957,N_1188,N_789);
xor U1958 (N_1958,N_183,N_413);
or U1959 (N_1959,N_1305,In_1073);
nand U1960 (N_1960,N_1358,In_932);
xnor U1961 (N_1961,In_764,N_1557);
or U1962 (N_1962,N_1332,N_1739);
nand U1963 (N_1963,In_1232,N_1417);
nand U1964 (N_1964,N_1253,N_1473);
xor U1965 (N_1965,In_2780,N_1551);
xor U1966 (N_1966,In_1595,N_660);
nor U1967 (N_1967,N_84,N_932);
or U1968 (N_1968,N_1503,N_1750);
nand U1969 (N_1969,N_1714,In_49);
xor U1970 (N_1970,N_1371,In_479);
nor U1971 (N_1971,N_942,N_1646);
or U1972 (N_1972,N_836,In_2724);
nand U1973 (N_1973,N_1418,N_1193);
and U1974 (N_1974,N_1622,N_1683);
xor U1975 (N_1975,N_941,N_1747);
nand U1976 (N_1976,N_1574,N_1217);
and U1977 (N_1977,N_1634,In_1715);
and U1978 (N_1978,N_1541,N_1227);
xnor U1979 (N_1979,N_1614,In_2623);
nand U1980 (N_1980,N_1243,N_1306);
and U1981 (N_1981,N_855,N_1212);
and U1982 (N_1982,N_1619,N_1533);
and U1983 (N_1983,N_1705,N_1490);
and U1984 (N_1984,N_813,In_2945);
and U1985 (N_1985,N_1480,In_1081);
nand U1986 (N_1986,N_1343,N_42);
or U1987 (N_1987,N_1610,N_378);
nor U1988 (N_1988,N_1208,N_1743);
and U1989 (N_1989,N_609,In_2614);
and U1990 (N_1990,N_1637,In_2470);
or U1991 (N_1991,N_45,N_1222);
or U1992 (N_1992,N_1562,N_55);
xor U1993 (N_1993,N_1286,In_1027);
nand U1994 (N_1994,N_1245,In_998);
and U1995 (N_1995,N_1475,N_1388);
nand U1996 (N_1996,N_1770,N_1050);
and U1997 (N_1997,N_1142,N_1233);
and U1998 (N_1998,N_1431,N_1372);
nor U1999 (N_1999,N_1008,In_2391);
nand U2000 (N_2000,In_1972,N_1559);
nand U2001 (N_2001,N_1547,N_1689);
or U2002 (N_2002,N_1720,N_1476);
xnor U2003 (N_2003,In_920,In_418);
nand U2004 (N_2004,N_1744,In_1441);
xnor U2005 (N_2005,N_1411,N_961);
xnor U2006 (N_2006,In_2036,N_1246);
xnor U2007 (N_2007,N_1267,N_1363);
or U2008 (N_2008,N_1460,N_1601);
xnor U2009 (N_2009,N_1223,N_914);
nand U2010 (N_2010,N_1264,N_49);
or U2011 (N_2011,N_1671,In_2461);
nand U2012 (N_2012,N_1586,N_1742);
and U2013 (N_2013,In_2135,N_801);
xor U2014 (N_2014,N_1229,N_1488);
nand U2015 (N_2015,N_1356,N_1006);
nor U2016 (N_2016,In_849,In_2298);
and U2017 (N_2017,N_1288,N_1755);
nor U2018 (N_2018,N_1693,In_1535);
xnor U2019 (N_2019,N_1401,N_840);
nand U2020 (N_2020,In_506,In_2609);
nor U2021 (N_2021,In_1020,N_889);
nor U2022 (N_2022,In_2854,In_2974);
xor U2023 (N_2023,N_1442,In_868);
nor U2024 (N_2024,N_1455,N_1540);
nor U2025 (N_2025,N_1030,N_57);
xor U2026 (N_2026,N_1277,N_677);
nand U2027 (N_2027,N_1546,In_2281);
xor U2028 (N_2028,In_2765,N_1038);
xor U2029 (N_2029,N_1216,In_2185);
nor U2030 (N_2030,N_1349,N_1387);
nor U2031 (N_2031,N_633,N_1572);
xnor U2032 (N_2032,N_1081,In_156);
nor U2033 (N_2033,N_1617,N_37);
nor U2034 (N_2034,N_598,N_175);
xnor U2035 (N_2035,N_1579,N_1782);
nand U2036 (N_2036,In_1082,N_1214);
nand U2037 (N_2037,N_359,N_588);
nor U2038 (N_2038,N_872,In_2327);
or U2039 (N_2039,N_653,In_839);
nor U2040 (N_2040,N_1472,N_1474);
nor U2041 (N_2041,N_1728,N_1684);
and U2042 (N_2042,N_1408,N_1652);
nor U2043 (N_2043,N_1434,N_748);
xnor U2044 (N_2044,In_2629,N_1373);
and U2045 (N_2045,N_1323,N_22);
or U2046 (N_2046,N_1284,In_2476);
and U2047 (N_2047,N_1379,N_56);
nor U2048 (N_2048,In_1114,In_1796);
xor U2049 (N_2049,N_845,N_1252);
nor U2050 (N_2050,In_1431,N_610);
xnor U2051 (N_2051,N_454,N_1364);
and U2052 (N_2052,N_1478,N_395);
nor U2053 (N_2053,In_202,N_1700);
xnor U2054 (N_2054,N_1199,N_1756);
or U2055 (N_2055,N_1051,N_1009);
nand U2056 (N_2056,N_1232,N_99);
and U2057 (N_2057,N_1534,N_1641);
and U2058 (N_2058,N_1470,N_1164);
or U2059 (N_2059,N_1263,N_1105);
xor U2060 (N_2060,N_226,N_701);
nor U2061 (N_2061,N_211,In_1850);
nor U2062 (N_2062,In_366,In_1057);
xor U2063 (N_2063,N_848,N_1202);
nand U2064 (N_2064,In_335,N_1231);
or U2065 (N_2065,In_1802,In_1650);
and U2066 (N_2066,N_669,N_1638);
xnor U2067 (N_2067,In_2356,In_416);
nand U2068 (N_2068,In_1379,N_759);
or U2069 (N_2069,N_1437,N_756);
nor U2070 (N_2070,N_1668,In_1612);
and U2071 (N_2071,N_1640,N_850);
nand U2072 (N_2072,N_854,N_1681);
and U2073 (N_2073,In_2681,N_1471);
and U2074 (N_2074,N_1108,N_1426);
or U2075 (N_2075,N_1315,In_2801);
nand U2076 (N_2076,N_1548,N_1642);
or U2077 (N_2077,N_594,N_894);
nand U2078 (N_2078,N_1173,In_805);
nand U2079 (N_2079,N_1778,N_1268);
or U2080 (N_2080,In_314,N_1194);
and U2081 (N_2081,N_1549,N_655);
nor U2082 (N_2082,In_489,N_1593);
or U2083 (N_2083,In_1217,In_540);
nor U2084 (N_2084,N_1502,In_1072);
or U2085 (N_2085,N_1644,N_809);
nand U2086 (N_2086,In_881,N_1447);
or U2087 (N_2087,N_1514,N_1327);
nor U2088 (N_2088,N_676,In_1048);
nor U2089 (N_2089,In_988,In_130);
nor U2090 (N_2090,N_1775,N_1287);
and U2091 (N_2091,N_1781,In_2415);
nor U2092 (N_2092,N_1624,N_1588);
and U2093 (N_2093,N_1695,N_1773);
nor U2094 (N_2094,In_1296,N_667);
nand U2095 (N_2095,N_1413,N_1377);
xor U2096 (N_2096,In_1888,N_1230);
nor U2097 (N_2097,N_1242,N_931);
nand U2098 (N_2098,In_451,N_1129);
nor U2099 (N_2099,N_1310,N_1236);
and U2100 (N_2100,In_2640,N_1621);
and U2101 (N_2101,N_1293,In_457);
nor U2102 (N_2102,N_322,In_2964);
and U2103 (N_2103,N_1353,N_1351);
xor U2104 (N_2104,In_1151,N_1752);
xor U2105 (N_2105,N_627,N_510);
and U2106 (N_2106,N_1690,N_1448);
nor U2107 (N_2107,N_1592,N_622);
or U2108 (N_2108,N_1324,N_1329);
nor U2109 (N_2109,N_269,In_2287);
xnor U2110 (N_2110,N_1708,N_346);
or U2111 (N_2111,In_2509,N_1078);
or U2112 (N_2112,N_1352,In_238);
nand U2113 (N_2113,N_1789,In_1314);
nand U2114 (N_2114,N_907,N_1799);
or U2115 (N_2115,N_1325,N_1454);
and U2116 (N_2116,In_1023,N_1585);
or U2117 (N_2117,In_1816,N_1779);
xor U2118 (N_2118,N_954,N_1368);
xnor U2119 (N_2119,N_1553,N_1334);
xor U2120 (N_2120,N_1425,N_509);
xnor U2121 (N_2121,N_1702,N_1282);
xnor U2122 (N_2122,N_1765,In_872);
xnor U2123 (N_2123,N_1532,N_1290);
and U2124 (N_2124,In_2932,In_319);
nor U2125 (N_2125,N_1057,N_233);
xnor U2126 (N_2126,In_634,In_1668);
nand U2127 (N_2127,In_2593,N_1479);
nand U2128 (N_2128,N_1258,N_1737);
xnor U2129 (N_2129,N_1114,N_1468);
or U2130 (N_2130,N_1654,In_1732);
xnor U2131 (N_2131,N_1218,In_1569);
and U2132 (N_2132,In_124,In_1077);
nor U2133 (N_2133,N_1701,N_387);
and U2134 (N_2134,N_1270,N_1026);
xor U2135 (N_2135,N_1526,N_1611);
xor U2136 (N_2136,N_1604,In_2617);
nor U2137 (N_2137,N_120,In_1353);
and U2138 (N_2138,In_2053,In_1418);
and U2139 (N_2139,N_1221,In_2714);
nor U2140 (N_2140,N_1724,In_2225);
or U2141 (N_2141,N_97,In_2657);
nand U2142 (N_2142,N_1272,N_1517);
or U2143 (N_2143,N_1754,N_1629);
nand U2144 (N_2144,N_1777,N_353);
nand U2145 (N_2145,N_890,N_671);
and U2146 (N_2146,In_1843,N_712);
nand U2147 (N_2147,N_1738,N_1636);
nand U2148 (N_2148,N_709,N_1620);
nor U2149 (N_2149,N_458,N_1336);
nor U2150 (N_2150,N_438,N_1589);
nand U2151 (N_2151,N_1392,In_95);
and U2152 (N_2152,N_1443,N_1615);
xor U2153 (N_2153,In_1971,N_1369);
nand U2154 (N_2154,N_1385,N_1481);
nor U2155 (N_2155,N_1685,N_216);
and U2156 (N_2156,N_1462,N_1791);
nand U2157 (N_2157,In_2365,N_1582);
xor U2158 (N_2158,N_710,N_1451);
or U2159 (N_2159,N_1319,N_212);
nor U2160 (N_2160,N_1639,N_1031);
nor U2161 (N_2161,N_568,In_579);
xor U2162 (N_2162,N_381,N_1433);
nand U2163 (N_2163,N_1511,N_145);
or U2164 (N_2164,In_2442,N_1444);
or U2165 (N_2165,In_1614,N_1130);
or U2166 (N_2166,N_1355,N_1203);
nor U2167 (N_2167,In_1521,N_1699);
nor U2168 (N_2168,In_2949,In_1079);
and U2169 (N_2169,N_1382,In_1788);
or U2170 (N_2170,In_2588,N_1259);
nor U2171 (N_2171,N_1465,N_1359);
and U2172 (N_2172,N_1322,N_1769);
xnor U2173 (N_2173,N_1672,N_1711);
or U2174 (N_2174,In_2569,N_1542);
or U2175 (N_2175,N_844,N_1657);
or U2176 (N_2176,N_1494,N_1261);
nand U2177 (N_2177,N_1354,N_1584);
or U2178 (N_2178,N_1571,N_664);
nand U2179 (N_2179,N_116,N_1722);
nand U2180 (N_2180,N_1543,In_28);
nand U2181 (N_2181,N_1453,In_171);
xor U2182 (N_2182,N_1544,N_1484);
nand U2183 (N_2183,N_1677,In_2808);
or U2184 (N_2184,N_773,N_1391);
xor U2185 (N_2185,N_152,N_1297);
or U2186 (N_2186,In_235,In_1294);
or U2187 (N_2187,In_1791,In_2676);
nand U2188 (N_2188,N_1458,N_1687);
nor U2189 (N_2189,N_1565,N_1577);
xor U2190 (N_2190,In_1568,N_1793);
or U2191 (N_2191,In_2189,In_25);
nand U2192 (N_2192,N_1461,N_1560);
or U2193 (N_2193,In_301,N_1321);
xnor U2194 (N_2194,N_1398,N_1341);
and U2195 (N_2195,In_528,N_1664);
or U2196 (N_2196,N_1745,N_83);
xnor U2197 (N_2197,N_1774,N_1215);
xnor U2198 (N_2198,N_1303,N_1432);
or U2199 (N_2199,N_923,In_2546);
and U2200 (N_2200,N_82,In_2405);
nand U2201 (N_2201,N_887,N_815);
and U2202 (N_2202,N_1380,N_1220);
and U2203 (N_2203,N_898,N_1420);
and U2204 (N_2204,N_1328,N_177);
nor U2205 (N_2205,N_1406,N_1643);
nor U2206 (N_2206,In_179,N_1456);
and U2207 (N_2207,N_1757,N_1240);
nor U2208 (N_2208,N_1414,N_1669);
xnor U2209 (N_2209,N_723,N_1254);
or U2210 (N_2210,N_1311,In_508);
and U2211 (N_2211,N_1338,N_1213);
or U2212 (N_2212,N_663,N_674);
nand U2213 (N_2213,In_2820,N_1292);
or U2214 (N_2214,N_1707,N_1662);
xor U2215 (N_2215,N_1570,N_1251);
or U2216 (N_2216,N_1709,In_281);
nor U2217 (N_2217,N_1122,N_1404);
xnor U2218 (N_2218,N_369,N_333);
nand U2219 (N_2219,N_1340,In_360);
nand U2220 (N_2220,N_1147,N_1331);
nor U2221 (N_2221,N_1086,N_1378);
nor U2222 (N_2222,N_945,N_1410);
nor U2223 (N_2223,N_752,In_879);
nand U2224 (N_2224,In_1123,N_876);
xnor U2225 (N_2225,In_2876,N_1271);
nand U2226 (N_2226,N_1630,N_1527);
nand U2227 (N_2227,In_2841,N_1496);
and U2228 (N_2228,N_1580,N_690);
xnor U2229 (N_2229,N_1710,N_1339);
or U2230 (N_2230,N_1749,In_2696);
and U2231 (N_2231,In_1021,N_162);
nor U2232 (N_2232,In_2195,N_27);
nor U2233 (N_2233,In_1591,N_1628);
or U2234 (N_2234,N_1656,N_1407);
nand U2235 (N_2235,N_1416,N_1761);
xnor U2236 (N_2236,N_953,In_1949);
or U2237 (N_2237,N_1647,In_1514);
and U2238 (N_2238,N_1278,In_2187);
xnor U2239 (N_2239,In_1990,N_1696);
nand U2240 (N_2240,N_1508,N_1510);
and U2241 (N_2241,N_1219,N_1054);
nand U2242 (N_2242,N_1501,N_1430);
or U2243 (N_2243,In_2209,N_1600);
nor U2244 (N_2244,N_1578,N_1489);
nor U2245 (N_2245,N_1608,N_974);
nor U2246 (N_2246,N_670,N_1552);
nor U2247 (N_2247,In_794,N_1760);
nand U2248 (N_2248,N_1625,N_1603);
xnor U2249 (N_2249,N_1375,N_1764);
nand U2250 (N_2250,N_12,N_1308);
and U2251 (N_2251,N_1659,N_617);
nor U2252 (N_2252,In_1459,N_1697);
nor U2253 (N_2253,N_1304,N_1041);
nand U2254 (N_2254,N_404,N_1317);
or U2255 (N_2255,N_831,N_1539);
nor U2256 (N_2256,In_350,N_1204);
and U2257 (N_2257,N_1665,N_437);
nor U2258 (N_2258,In_2416,N_1704);
and U2259 (N_2259,In_606,N_1459);
and U2260 (N_2260,N_1515,N_1660);
and U2261 (N_2261,In_2653,In_311);
and U2262 (N_2262,In_2141,N_1741);
nand U2263 (N_2263,N_1072,N_1397);
nand U2264 (N_2264,N_401,In_2992);
xnor U2265 (N_2265,N_1751,N_1522);
or U2266 (N_2266,N_1158,N_309);
nor U2267 (N_2267,In_2831,In_835);
xor U2268 (N_2268,N_1337,N_285);
or U2269 (N_2269,N_1618,N_1691);
nor U2270 (N_2270,N_1680,N_1607);
nand U2271 (N_2271,N_987,N_1127);
xor U2272 (N_2272,N_1381,In_46);
nor U2273 (N_2273,N_1556,In_2292);
and U2274 (N_2274,N_1365,N_156);
or U2275 (N_2275,N_1512,N_1790);
nor U2276 (N_2276,In_2274,In_243);
nor U2277 (N_2277,N_689,In_907);
xnor U2278 (N_2278,N_1260,In_1338);
nor U2279 (N_2279,N_1281,N_1146);
xnor U2280 (N_2280,In_911,N_668);
nand U2281 (N_2281,N_1594,N_1520);
and U2282 (N_2282,In_782,In_2969);
xor U2283 (N_2283,N_1599,In_2994);
nor U2284 (N_2284,In_2598,N_1788);
or U2285 (N_2285,N_1429,N_1536);
nor U2286 (N_2286,N_1609,N_1597);
and U2287 (N_2287,In_228,N_85);
nor U2288 (N_2288,N_1097,N_1731);
or U2289 (N_2289,N_693,N_1234);
nor U2290 (N_2290,N_1100,N_1262);
nand U2291 (N_2291,In_903,N_1053);
nor U2292 (N_2292,N_1342,In_1744);
or U2293 (N_2293,N_1428,N_678);
nand U2294 (N_2294,N_1273,N_1734);
nor U2295 (N_2295,N_356,N_658);
or U2296 (N_2296,N_1666,In_2229);
or U2297 (N_2297,N_635,N_1727);
nand U2298 (N_2298,N_1111,N_1457);
nand U2299 (N_2299,N_1389,N_1348);
and U2300 (N_2300,N_1396,N_1797);
nor U2301 (N_2301,N_1209,N_884);
nand U2302 (N_2302,N_1393,N_1673);
nor U2303 (N_2303,N_1237,N_1445);
and U2304 (N_2304,In_1847,In_1735);
and U2305 (N_2305,N_1200,N_1482);
or U2306 (N_2306,N_1424,In_546);
or U2307 (N_2307,In_1985,N_973);
nand U2308 (N_2308,N_258,N_1550);
nor U2309 (N_2309,N_860,In_536);
or U2310 (N_2310,N_919,N_1415);
and U2311 (N_2311,In_784,In_2432);
nand U2312 (N_2312,N_1569,N_1386);
xnor U2313 (N_2313,N_1645,N_1784);
nor U2314 (N_2314,N_1126,N_820);
xnor U2315 (N_2315,In_1039,N_95);
or U2316 (N_2316,N_340,N_1467);
and U2317 (N_2317,In_2496,In_531);
nand U2318 (N_2318,N_1648,N_816);
xor U2319 (N_2319,In_89,N_656);
nand U2320 (N_2320,N_1716,N_725);
or U2321 (N_2321,In_609,N_1561);
nand U2322 (N_2322,N_870,N_1499);
or U2323 (N_2323,N_1531,N_1717);
xnor U2324 (N_2324,N_1596,N_904);
nor U2325 (N_2325,N_72,N_1675);
xnor U2326 (N_2326,N_1591,N_317);
or U2327 (N_2327,N_1787,N_1692);
or U2328 (N_2328,N_1595,N_1486);
nand U2329 (N_2329,N_1682,In_2996);
nor U2330 (N_2330,N_1529,N_403);
or U2331 (N_2331,N_1530,N_1226);
or U2332 (N_2332,N_467,N_392);
and U2333 (N_2333,N_1161,N_1241);
nand U2334 (N_2334,N_1312,N_770);
nor U2335 (N_2335,In_2639,In_2581);
xor U2336 (N_2336,N_1573,N_646);
and U2337 (N_2337,N_1294,N_834);
nand U2338 (N_2338,N_1498,N_918);
nand U2339 (N_2339,N_1612,In_2938);
nor U2340 (N_2340,N_1518,N_1436);
or U2341 (N_2341,In_2438,In_1463);
nand U2342 (N_2342,N_1798,N_1266);
or U2343 (N_2343,N_94,N_1419);
xor U2344 (N_2344,In_1746,In_346);
or U2345 (N_2345,N_1725,N_803);
and U2346 (N_2346,N_1713,N_1676);
nor U2347 (N_2347,N_1394,N_534);
or U2348 (N_2348,In_27,N_682);
or U2349 (N_2349,In_1245,N_1581);
nor U2350 (N_2350,In_2079,N_1606);
nand U2351 (N_2351,In_720,N_1729);
xor U2352 (N_2352,N_1248,N_151);
xnor U2353 (N_2353,N_993,In_287);
or U2354 (N_2354,N_1412,In_1774);
nor U2355 (N_2355,N_1283,In_1035);
and U2356 (N_2356,N_514,N_1269);
nor U2357 (N_2357,N_826,N_1201);
and U2358 (N_2358,N_1399,N_1477);
xnor U2359 (N_2359,N_1302,In_2513);
and U2360 (N_2360,N_288,N_1545);
or U2361 (N_2361,In_659,In_2891);
or U2362 (N_2362,In_2700,N_873);
and U2363 (N_2363,N_1289,N_1771);
and U2364 (N_2364,N_1795,N_985);
nand U2365 (N_2365,In_2902,N_1723);
or U2366 (N_2366,In_873,In_2471);
and U2367 (N_2367,In_1769,N_1783);
xor U2368 (N_2368,N_1295,In_2566);
xnor U2369 (N_2369,N_1776,N_1631);
xor U2370 (N_2370,N_1441,N_1107);
xnor U2371 (N_2371,N_1537,N_1500);
nand U2372 (N_2372,N_1346,N_1715);
xor U2373 (N_2373,N_1064,N_740);
nand U2374 (N_2374,N_1583,N_540);
xnor U2375 (N_2375,In_2113,In_829);
and U2376 (N_2376,In_1280,N_1156);
and U2377 (N_2377,N_1023,N_1563);
nor U2378 (N_2378,N_881,N_794);
xnor U2379 (N_2379,N_1384,N_623);
and U2380 (N_2380,N_1633,In_1438);
or U2381 (N_2381,N_1376,N_1238);
xor U2382 (N_2382,N_1505,In_893);
and U2383 (N_2383,N_1195,N_1138);
nand U2384 (N_2384,In_266,N_1265);
nor U2385 (N_2385,N_1555,N_1564);
or U2386 (N_2386,N_1438,N_1590);
and U2387 (N_2387,In_2968,N_611);
and U2388 (N_2388,N_1703,N_427);
nor U2389 (N_2389,In_1318,N_1255);
and U2390 (N_2390,N_1291,N_1602);
and U2391 (N_2391,N_1538,N_1360);
xor U2392 (N_2392,N_1019,In_2373);
xor U2393 (N_2393,N_902,N_978);
nand U2394 (N_2394,N_1495,N_995);
nand U2395 (N_2395,N_255,In_1038);
or U2396 (N_2396,In_853,N_1721);
nand U2397 (N_2397,N_1279,N_852);
xnor U2398 (N_2398,N_1296,In_2282);
nand U2399 (N_2399,N_680,In_704);
xor U2400 (N_2400,N_1960,N_2059);
and U2401 (N_2401,N_1869,N_2222);
nor U2402 (N_2402,N_2194,N_2012);
and U2403 (N_2403,N_2296,N_1953);
or U2404 (N_2404,N_2021,N_2195);
nand U2405 (N_2405,N_2058,N_2193);
xnor U2406 (N_2406,N_2113,N_2117);
and U2407 (N_2407,N_1959,N_1966);
xor U2408 (N_2408,N_1996,N_2197);
nor U2409 (N_2409,N_2251,N_1933);
nand U2410 (N_2410,N_1870,N_2125);
and U2411 (N_2411,N_2147,N_1859);
or U2412 (N_2412,N_2019,N_2110);
or U2413 (N_2413,N_1817,N_2280);
nor U2414 (N_2414,N_1812,N_2250);
nand U2415 (N_2415,N_2100,N_2300);
xor U2416 (N_2416,N_1882,N_2144);
and U2417 (N_2417,N_1905,N_2173);
nor U2418 (N_2418,N_2078,N_1855);
nor U2419 (N_2419,N_1989,N_2281);
nor U2420 (N_2420,N_1874,N_2308);
or U2421 (N_2421,N_1974,N_2364);
nand U2422 (N_2422,N_2156,N_2084);
and U2423 (N_2423,N_2092,N_2027);
and U2424 (N_2424,N_1920,N_2130);
or U2425 (N_2425,N_1861,N_2180);
nor U2426 (N_2426,N_2097,N_1913);
xnor U2427 (N_2427,N_2020,N_2052);
or U2428 (N_2428,N_1884,N_1810);
xor U2429 (N_2429,N_2140,N_1973);
xor U2430 (N_2430,N_1946,N_2157);
xor U2431 (N_2431,N_2391,N_2079);
nor U2432 (N_2432,N_2284,N_2234);
and U2433 (N_2433,N_1995,N_2361);
or U2434 (N_2434,N_2323,N_1878);
and U2435 (N_2435,N_1942,N_2080);
or U2436 (N_2436,N_2353,N_2388);
nor U2437 (N_2437,N_2282,N_1820);
nor U2438 (N_2438,N_1956,N_2287);
or U2439 (N_2439,N_2396,N_2082);
nand U2440 (N_2440,N_2236,N_2273);
nor U2441 (N_2441,N_2106,N_2261);
xnor U2442 (N_2442,N_2056,N_2008);
xor U2443 (N_2443,N_1868,N_1807);
or U2444 (N_2444,N_2153,N_1916);
nand U2445 (N_2445,N_2270,N_2238);
nand U2446 (N_2446,N_2395,N_1952);
and U2447 (N_2447,N_2062,N_1890);
nor U2448 (N_2448,N_2101,N_2057);
and U2449 (N_2449,N_2038,N_2049);
or U2450 (N_2450,N_1816,N_1990);
xnor U2451 (N_2451,N_2136,N_2346);
nand U2452 (N_2452,N_1903,N_2112);
or U2453 (N_2453,N_1912,N_2329);
or U2454 (N_2454,N_2002,N_2149);
xor U2455 (N_2455,N_2132,N_2143);
nor U2456 (N_2456,N_2174,N_2202);
and U2457 (N_2457,N_2286,N_2335);
nand U2458 (N_2458,N_1899,N_2216);
xor U2459 (N_2459,N_2349,N_1840);
and U2460 (N_2460,N_2217,N_2248);
xnor U2461 (N_2461,N_2184,N_2225);
nor U2462 (N_2462,N_2294,N_2321);
xnor U2463 (N_2463,N_2145,N_2375);
or U2464 (N_2464,N_2191,N_2179);
nor U2465 (N_2465,N_2382,N_1934);
or U2466 (N_2466,N_2182,N_2271);
xnor U2467 (N_2467,N_2289,N_2133);
or U2468 (N_2468,N_1944,N_2172);
xnor U2469 (N_2469,N_2000,N_1997);
or U2470 (N_2470,N_2047,N_2029);
and U2471 (N_2471,N_1876,N_2275);
and U2472 (N_2472,N_2011,N_1802);
nand U2473 (N_2473,N_2360,N_2031);
and U2474 (N_2474,N_2071,N_2241);
and U2475 (N_2475,N_1862,N_2231);
and U2476 (N_2476,N_1842,N_2098);
nor U2477 (N_2477,N_2381,N_1814);
xnor U2478 (N_2478,N_2355,N_1830);
nor U2479 (N_2479,N_1845,N_1841);
or U2480 (N_2480,N_1945,N_1888);
xnor U2481 (N_2481,N_1809,N_2091);
xnor U2482 (N_2482,N_1894,N_2336);
nand U2483 (N_2483,N_2229,N_1887);
and U2484 (N_2484,N_2134,N_2189);
nand U2485 (N_2485,N_1914,N_1927);
nor U2486 (N_2486,N_2066,N_2010);
or U2487 (N_2487,N_2154,N_2207);
and U2488 (N_2488,N_2164,N_2218);
or U2489 (N_2489,N_1972,N_1836);
or U2490 (N_2490,N_2030,N_2311);
nand U2491 (N_2491,N_1801,N_2252);
and U2492 (N_2492,N_2256,N_2373);
nor U2493 (N_2493,N_2387,N_2032);
or U2494 (N_2494,N_2260,N_2116);
nand U2495 (N_2495,N_1994,N_1804);
or U2496 (N_2496,N_1929,N_2070);
nand U2497 (N_2497,N_2259,N_1950);
nand U2498 (N_2498,N_2269,N_1900);
and U2499 (N_2499,N_1980,N_1993);
xnor U2500 (N_2500,N_2095,N_2240);
and U2501 (N_2501,N_1850,N_2114);
or U2502 (N_2502,N_1825,N_1856);
nor U2503 (N_2503,N_2288,N_2239);
and U2504 (N_2504,N_2334,N_1981);
xor U2505 (N_2505,N_2371,N_2013);
nand U2506 (N_2506,N_2188,N_2087);
and U2507 (N_2507,N_1827,N_1925);
xnor U2508 (N_2508,N_1977,N_2036);
nand U2509 (N_2509,N_2190,N_2043);
nor U2510 (N_2510,N_2158,N_2046);
nand U2511 (N_2511,N_2226,N_2119);
or U2512 (N_2512,N_2312,N_2099);
nor U2513 (N_2513,N_2139,N_2293);
xnor U2514 (N_2514,N_2061,N_2257);
nor U2515 (N_2515,N_2331,N_2210);
and U2516 (N_2516,N_2372,N_2244);
nor U2517 (N_2517,N_1931,N_2050);
nor U2518 (N_2518,N_1898,N_1935);
nand U2519 (N_2519,N_2276,N_2384);
or U2520 (N_2520,N_2150,N_1938);
nor U2521 (N_2521,N_2024,N_1979);
xnor U2522 (N_2522,N_2040,N_1808);
and U2523 (N_2523,N_2304,N_2185);
nand U2524 (N_2524,N_2333,N_1860);
xor U2525 (N_2525,N_2128,N_1853);
or U2526 (N_2526,N_2124,N_2378);
nand U2527 (N_2527,N_2295,N_2068);
xnor U2528 (N_2528,N_2390,N_2298);
and U2529 (N_2529,N_2303,N_1919);
xor U2530 (N_2530,N_2351,N_2060);
or U2531 (N_2531,N_1928,N_2332);
nand U2532 (N_2532,N_2186,N_2096);
xor U2533 (N_2533,N_1881,N_2392);
or U2534 (N_2534,N_1984,N_2368);
and U2535 (N_2535,N_2352,N_2007);
or U2536 (N_2536,N_2268,N_2039);
and U2537 (N_2537,N_2135,N_1987);
xor U2538 (N_2538,N_2350,N_1922);
or U2539 (N_2539,N_2033,N_2347);
or U2540 (N_2540,N_1969,N_2126);
nand U2541 (N_2541,N_2115,N_1924);
and U2542 (N_2542,N_1883,N_2196);
nor U2543 (N_2543,N_2363,N_2192);
xnor U2544 (N_2544,N_2200,N_2077);
or U2545 (N_2545,N_1964,N_1967);
or U2546 (N_2546,N_2067,N_1937);
and U2547 (N_2547,N_2305,N_1958);
nor U2548 (N_2548,N_2072,N_2069);
and U2549 (N_2549,N_1858,N_2309);
xor U2550 (N_2550,N_2328,N_2083);
nand U2551 (N_2551,N_2121,N_1803);
nand U2552 (N_2552,N_2063,N_2205);
and U2553 (N_2553,N_2314,N_2074);
or U2554 (N_2554,N_1819,N_2064);
nor U2555 (N_2555,N_1889,N_2006);
nand U2556 (N_2556,N_1811,N_1940);
nand U2557 (N_2557,N_2348,N_2004);
or U2558 (N_2558,N_1828,N_2341);
or U2559 (N_2559,N_2003,N_2243);
or U2560 (N_2560,N_2223,N_2340);
nor U2561 (N_2561,N_1831,N_2111);
or U2562 (N_2562,N_2208,N_1902);
or U2563 (N_2563,N_2397,N_1951);
or U2564 (N_2564,N_2255,N_2247);
or U2565 (N_2565,N_2263,N_2262);
and U2566 (N_2566,N_2264,N_1955);
xnor U2567 (N_2567,N_2142,N_2224);
or U2568 (N_2568,N_1849,N_2160);
or U2569 (N_2569,N_2338,N_2344);
or U2570 (N_2570,N_2141,N_2317);
and U2571 (N_2571,N_1926,N_2380);
xnor U2572 (N_2572,N_2310,N_1908);
or U2573 (N_2573,N_2118,N_1833);
nand U2574 (N_2574,N_2151,N_2389);
xor U2575 (N_2575,N_2237,N_2242);
nand U2576 (N_2576,N_2206,N_1854);
and U2577 (N_2577,N_1843,N_2102);
and U2578 (N_2578,N_1896,N_1906);
xnor U2579 (N_2579,N_1901,N_2266);
nor U2580 (N_2580,N_2176,N_2219);
nor U2581 (N_2581,N_1975,N_2122);
nor U2582 (N_2582,N_2028,N_1839);
nor U2583 (N_2583,N_2175,N_2204);
nor U2584 (N_2584,N_2162,N_2220);
xor U2585 (N_2585,N_1948,N_1939);
and U2586 (N_2586,N_2386,N_2367);
nor U2587 (N_2587,N_2094,N_2358);
and U2588 (N_2588,N_1872,N_1991);
or U2589 (N_2589,N_2227,N_2327);
or U2590 (N_2590,N_2169,N_1863);
nor U2591 (N_2591,N_2283,N_1879);
nor U2592 (N_2592,N_2107,N_2325);
and U2593 (N_2593,N_2265,N_2369);
xor U2594 (N_2594,N_1886,N_2258);
or U2595 (N_2595,N_2354,N_1986);
xnor U2596 (N_2596,N_2177,N_2076);
nand U2597 (N_2597,N_2167,N_2155);
nand U2598 (N_2598,N_2320,N_2277);
and U2599 (N_2599,N_2088,N_1821);
xnor U2600 (N_2600,N_1805,N_1982);
nor U2601 (N_2601,N_1992,N_2326);
nor U2602 (N_2602,N_2221,N_2009);
xnor U2603 (N_2603,N_1909,N_1943);
or U2604 (N_2604,N_2018,N_2103);
nand U2605 (N_2605,N_1880,N_2137);
xnor U2606 (N_2606,N_2232,N_2399);
and U2607 (N_2607,N_2307,N_2365);
or U2608 (N_2608,N_1985,N_2345);
nor U2609 (N_2609,N_2376,N_2214);
xor U2610 (N_2610,N_2356,N_2168);
and U2611 (N_2611,N_1970,N_1852);
or U2612 (N_2612,N_2171,N_2291);
nand U2613 (N_2613,N_2198,N_2152);
and U2614 (N_2614,N_2212,N_2343);
nand U2615 (N_2615,N_2104,N_2090);
nand U2616 (N_2616,N_2051,N_1893);
nand U2617 (N_2617,N_2374,N_2274);
nor U2618 (N_2618,N_2123,N_1947);
xor U2619 (N_2619,N_1978,N_2035);
nor U2620 (N_2620,N_2015,N_2319);
nor U2621 (N_2621,N_2394,N_1941);
or U2622 (N_2622,N_2215,N_1961);
xor U2623 (N_2623,N_2054,N_2301);
and U2624 (N_2624,N_2235,N_2163);
nor U2625 (N_2625,N_2086,N_2034);
or U2626 (N_2626,N_2302,N_2249);
nand U2627 (N_2627,N_1949,N_1954);
nand U2628 (N_2628,N_2203,N_2201);
and U2629 (N_2629,N_2048,N_1846);
nand U2630 (N_2630,N_2045,N_2016);
and U2631 (N_2631,N_1822,N_1848);
nor U2632 (N_2632,N_1871,N_2127);
nor U2633 (N_2633,N_2362,N_2005);
nor U2634 (N_2634,N_1865,N_1968);
and U2635 (N_2635,N_1907,N_1818);
or U2636 (N_2636,N_1867,N_2272);
or U2637 (N_2637,N_2120,N_2254);
nor U2638 (N_2638,N_2379,N_2209);
and U2639 (N_2639,N_1832,N_2278);
nand U2640 (N_2640,N_1963,N_2181);
nor U2641 (N_2641,N_1838,N_2089);
and U2642 (N_2642,N_2285,N_2297);
or U2643 (N_2643,N_2159,N_2318);
or U2644 (N_2644,N_2041,N_1976);
xor U2645 (N_2645,N_2148,N_1835);
or U2646 (N_2646,N_2245,N_1813);
or U2647 (N_2647,N_2267,N_2037);
xor U2648 (N_2648,N_1800,N_1965);
or U2649 (N_2649,N_2383,N_2053);
or U2650 (N_2650,N_2183,N_2025);
nand U2651 (N_2651,N_1891,N_1844);
xor U2652 (N_2652,N_2366,N_2138);
or U2653 (N_2653,N_1999,N_1851);
nor U2654 (N_2654,N_1904,N_2306);
or U2655 (N_2655,N_2055,N_2023);
xor U2656 (N_2656,N_1877,N_2017);
xor U2657 (N_2657,N_2165,N_2001);
or U2658 (N_2658,N_2131,N_1915);
or U2659 (N_2659,N_2290,N_2044);
nor U2660 (N_2660,N_2075,N_2315);
nand U2661 (N_2661,N_1936,N_2246);
nand U2662 (N_2662,N_2211,N_1917);
or U2663 (N_2663,N_1875,N_1988);
or U2664 (N_2664,N_2393,N_2370);
nor U2665 (N_2665,N_1918,N_1873);
xnor U2666 (N_2666,N_2178,N_2166);
nand U2667 (N_2667,N_2316,N_1895);
nand U2668 (N_2668,N_2199,N_1932);
nand U2669 (N_2669,N_1834,N_1971);
nor U2670 (N_2670,N_1857,N_2337);
nor U2671 (N_2671,N_2279,N_1864);
nand U2672 (N_2672,N_1923,N_2299);
xnor U2673 (N_2673,N_2292,N_2170);
xnor U2674 (N_2674,N_2065,N_2109);
nand U2675 (N_2675,N_2022,N_1911);
and U2676 (N_2676,N_1837,N_1866);
and U2677 (N_2677,N_2377,N_2085);
or U2678 (N_2678,N_2233,N_1962);
xor U2679 (N_2679,N_2339,N_2105);
nor U2680 (N_2680,N_2357,N_2228);
or U2681 (N_2681,N_1815,N_2398);
xor U2682 (N_2682,N_1806,N_2253);
nand U2683 (N_2683,N_2330,N_2093);
or U2684 (N_2684,N_1885,N_1892);
nor U2685 (N_2685,N_1921,N_1930);
nor U2686 (N_2686,N_1897,N_2073);
or U2687 (N_2687,N_2342,N_2146);
or U2688 (N_2688,N_2359,N_2313);
and U2689 (N_2689,N_1998,N_2230);
or U2690 (N_2690,N_1824,N_2385);
or U2691 (N_2691,N_2081,N_2108);
xor U2692 (N_2692,N_2213,N_1829);
nor U2693 (N_2693,N_2129,N_2187);
xor U2694 (N_2694,N_1823,N_2026);
nor U2695 (N_2695,N_1957,N_2042);
and U2696 (N_2696,N_1847,N_2324);
or U2697 (N_2697,N_1910,N_1826);
xnor U2698 (N_2698,N_2322,N_2014);
xnor U2699 (N_2699,N_2161,N_1983);
nor U2700 (N_2700,N_1848,N_2209);
and U2701 (N_2701,N_2310,N_1997);
and U2702 (N_2702,N_2166,N_1971);
and U2703 (N_2703,N_2169,N_2186);
nand U2704 (N_2704,N_2300,N_2216);
or U2705 (N_2705,N_2243,N_2277);
xnor U2706 (N_2706,N_2288,N_1943);
or U2707 (N_2707,N_2298,N_1916);
or U2708 (N_2708,N_1913,N_2052);
xor U2709 (N_2709,N_1806,N_2026);
xor U2710 (N_2710,N_2161,N_2265);
nor U2711 (N_2711,N_2392,N_1976);
and U2712 (N_2712,N_1981,N_1872);
xor U2713 (N_2713,N_1998,N_1888);
and U2714 (N_2714,N_2071,N_1937);
and U2715 (N_2715,N_1821,N_1985);
nand U2716 (N_2716,N_2289,N_2346);
nand U2717 (N_2717,N_2030,N_1835);
xor U2718 (N_2718,N_2396,N_1807);
or U2719 (N_2719,N_1984,N_1910);
nor U2720 (N_2720,N_1853,N_2218);
and U2721 (N_2721,N_2268,N_2145);
or U2722 (N_2722,N_1885,N_2026);
and U2723 (N_2723,N_2349,N_2362);
or U2724 (N_2724,N_2194,N_1983);
or U2725 (N_2725,N_2116,N_1835);
and U2726 (N_2726,N_2380,N_2124);
xor U2727 (N_2727,N_2373,N_2079);
or U2728 (N_2728,N_2148,N_2261);
or U2729 (N_2729,N_2298,N_1848);
nand U2730 (N_2730,N_1899,N_1970);
nor U2731 (N_2731,N_2321,N_2006);
nor U2732 (N_2732,N_2200,N_2286);
xnor U2733 (N_2733,N_1851,N_2316);
or U2734 (N_2734,N_1979,N_2279);
xor U2735 (N_2735,N_2001,N_2130);
xor U2736 (N_2736,N_1838,N_2041);
and U2737 (N_2737,N_1986,N_2225);
nand U2738 (N_2738,N_2252,N_2198);
or U2739 (N_2739,N_1886,N_2177);
and U2740 (N_2740,N_2031,N_2272);
and U2741 (N_2741,N_1946,N_2376);
nand U2742 (N_2742,N_2323,N_2109);
or U2743 (N_2743,N_2239,N_1978);
nand U2744 (N_2744,N_1947,N_2325);
xnor U2745 (N_2745,N_2322,N_1879);
and U2746 (N_2746,N_2114,N_1958);
or U2747 (N_2747,N_1830,N_2310);
and U2748 (N_2748,N_2096,N_1880);
and U2749 (N_2749,N_2115,N_1996);
xnor U2750 (N_2750,N_2386,N_2258);
xor U2751 (N_2751,N_2338,N_2184);
nor U2752 (N_2752,N_2376,N_1865);
xor U2753 (N_2753,N_1819,N_2032);
nand U2754 (N_2754,N_2009,N_2334);
nor U2755 (N_2755,N_2009,N_2387);
nor U2756 (N_2756,N_1961,N_1837);
nor U2757 (N_2757,N_2010,N_2069);
nand U2758 (N_2758,N_2302,N_2299);
or U2759 (N_2759,N_2102,N_1910);
nor U2760 (N_2760,N_2194,N_2168);
xnor U2761 (N_2761,N_2090,N_2051);
nand U2762 (N_2762,N_2229,N_2136);
nor U2763 (N_2763,N_2046,N_2000);
or U2764 (N_2764,N_2204,N_2163);
and U2765 (N_2765,N_1920,N_1923);
or U2766 (N_2766,N_1800,N_2122);
and U2767 (N_2767,N_1847,N_2317);
nand U2768 (N_2768,N_1899,N_2246);
nor U2769 (N_2769,N_2024,N_2175);
nor U2770 (N_2770,N_2381,N_2063);
nor U2771 (N_2771,N_2174,N_1985);
or U2772 (N_2772,N_2308,N_1885);
nor U2773 (N_2773,N_2164,N_1915);
nand U2774 (N_2774,N_2261,N_1957);
xor U2775 (N_2775,N_2144,N_1996);
xor U2776 (N_2776,N_1906,N_2216);
and U2777 (N_2777,N_1903,N_2341);
nand U2778 (N_2778,N_1840,N_1961);
and U2779 (N_2779,N_2089,N_2232);
and U2780 (N_2780,N_2267,N_2295);
xor U2781 (N_2781,N_1869,N_1935);
and U2782 (N_2782,N_2027,N_1989);
nor U2783 (N_2783,N_2363,N_2058);
nor U2784 (N_2784,N_2249,N_2145);
nor U2785 (N_2785,N_2188,N_2041);
xnor U2786 (N_2786,N_2019,N_1971);
xnor U2787 (N_2787,N_2212,N_2333);
nand U2788 (N_2788,N_2203,N_2138);
and U2789 (N_2789,N_2287,N_1965);
and U2790 (N_2790,N_1982,N_2247);
xnor U2791 (N_2791,N_2146,N_2000);
and U2792 (N_2792,N_2181,N_1807);
nand U2793 (N_2793,N_2032,N_2021);
and U2794 (N_2794,N_1927,N_2120);
or U2795 (N_2795,N_2220,N_1817);
nor U2796 (N_2796,N_2099,N_1943);
and U2797 (N_2797,N_2370,N_2211);
xor U2798 (N_2798,N_2198,N_1856);
and U2799 (N_2799,N_2166,N_1807);
xnor U2800 (N_2800,N_1912,N_2065);
and U2801 (N_2801,N_1886,N_1883);
xnor U2802 (N_2802,N_2151,N_1800);
nor U2803 (N_2803,N_2329,N_2319);
and U2804 (N_2804,N_2273,N_1972);
nor U2805 (N_2805,N_2307,N_2052);
xnor U2806 (N_2806,N_2046,N_2348);
or U2807 (N_2807,N_2177,N_1996);
nor U2808 (N_2808,N_2194,N_2379);
xnor U2809 (N_2809,N_2390,N_1907);
nand U2810 (N_2810,N_1806,N_1975);
xnor U2811 (N_2811,N_2346,N_2032);
nor U2812 (N_2812,N_1839,N_2199);
xnor U2813 (N_2813,N_2088,N_2394);
nand U2814 (N_2814,N_1877,N_1923);
and U2815 (N_2815,N_1984,N_2280);
nand U2816 (N_2816,N_2063,N_2056);
nor U2817 (N_2817,N_2374,N_2013);
nor U2818 (N_2818,N_2192,N_2050);
or U2819 (N_2819,N_2040,N_1851);
nand U2820 (N_2820,N_2388,N_2082);
nor U2821 (N_2821,N_2399,N_1919);
nand U2822 (N_2822,N_2141,N_2069);
nor U2823 (N_2823,N_1945,N_2315);
or U2824 (N_2824,N_2312,N_2229);
nand U2825 (N_2825,N_2070,N_2033);
xor U2826 (N_2826,N_1800,N_1876);
nor U2827 (N_2827,N_2324,N_2168);
nand U2828 (N_2828,N_1933,N_1939);
xnor U2829 (N_2829,N_1834,N_2217);
nor U2830 (N_2830,N_2134,N_2398);
and U2831 (N_2831,N_1812,N_2084);
or U2832 (N_2832,N_1975,N_2000);
xor U2833 (N_2833,N_1867,N_2383);
nor U2834 (N_2834,N_1917,N_2333);
and U2835 (N_2835,N_2185,N_2067);
xnor U2836 (N_2836,N_2318,N_2024);
or U2837 (N_2837,N_2350,N_1867);
nor U2838 (N_2838,N_2159,N_2258);
nand U2839 (N_2839,N_2141,N_2133);
nor U2840 (N_2840,N_2096,N_2250);
or U2841 (N_2841,N_2165,N_1898);
xor U2842 (N_2842,N_2037,N_2173);
and U2843 (N_2843,N_2022,N_2162);
and U2844 (N_2844,N_2338,N_2106);
and U2845 (N_2845,N_1900,N_2207);
xor U2846 (N_2846,N_2144,N_2022);
or U2847 (N_2847,N_2252,N_1806);
and U2848 (N_2848,N_1895,N_2313);
and U2849 (N_2849,N_2251,N_1837);
xor U2850 (N_2850,N_2079,N_2294);
or U2851 (N_2851,N_2068,N_2297);
or U2852 (N_2852,N_2002,N_2015);
or U2853 (N_2853,N_2372,N_1890);
nor U2854 (N_2854,N_1912,N_1973);
nor U2855 (N_2855,N_1910,N_2241);
nor U2856 (N_2856,N_2363,N_2316);
nand U2857 (N_2857,N_2328,N_1827);
nor U2858 (N_2858,N_2085,N_2380);
or U2859 (N_2859,N_2219,N_2201);
and U2860 (N_2860,N_2210,N_2287);
nand U2861 (N_2861,N_2085,N_2304);
nor U2862 (N_2862,N_1976,N_1874);
xnor U2863 (N_2863,N_2219,N_2041);
xor U2864 (N_2864,N_2271,N_2330);
xnor U2865 (N_2865,N_1870,N_1809);
or U2866 (N_2866,N_1803,N_2081);
nor U2867 (N_2867,N_2010,N_2156);
and U2868 (N_2868,N_2076,N_2344);
and U2869 (N_2869,N_2134,N_2222);
and U2870 (N_2870,N_2115,N_1958);
xnor U2871 (N_2871,N_2148,N_1814);
and U2872 (N_2872,N_2053,N_1836);
nand U2873 (N_2873,N_2172,N_2238);
or U2874 (N_2874,N_1851,N_2337);
and U2875 (N_2875,N_1893,N_1828);
nor U2876 (N_2876,N_2364,N_2036);
or U2877 (N_2877,N_2163,N_1928);
or U2878 (N_2878,N_2119,N_1826);
or U2879 (N_2879,N_1843,N_2028);
nand U2880 (N_2880,N_1850,N_1837);
xnor U2881 (N_2881,N_2334,N_2046);
or U2882 (N_2882,N_1980,N_1904);
or U2883 (N_2883,N_1855,N_2305);
nor U2884 (N_2884,N_1951,N_1995);
nand U2885 (N_2885,N_1884,N_2084);
or U2886 (N_2886,N_2078,N_2054);
or U2887 (N_2887,N_2158,N_2110);
nand U2888 (N_2888,N_2016,N_2015);
and U2889 (N_2889,N_2145,N_2000);
nor U2890 (N_2890,N_1865,N_1809);
nand U2891 (N_2891,N_2339,N_2397);
or U2892 (N_2892,N_2007,N_2353);
xor U2893 (N_2893,N_1820,N_1928);
nand U2894 (N_2894,N_1841,N_2272);
nand U2895 (N_2895,N_2395,N_1828);
nand U2896 (N_2896,N_1905,N_2176);
nand U2897 (N_2897,N_2318,N_1884);
nand U2898 (N_2898,N_2117,N_2179);
and U2899 (N_2899,N_2230,N_1955);
and U2900 (N_2900,N_2081,N_2042);
nand U2901 (N_2901,N_1812,N_1817);
nor U2902 (N_2902,N_1998,N_2089);
nand U2903 (N_2903,N_2361,N_2137);
or U2904 (N_2904,N_2198,N_1911);
nor U2905 (N_2905,N_2344,N_2296);
nor U2906 (N_2906,N_1869,N_1987);
and U2907 (N_2907,N_2201,N_2322);
nor U2908 (N_2908,N_1885,N_2249);
or U2909 (N_2909,N_2266,N_2219);
nand U2910 (N_2910,N_2245,N_2120);
nand U2911 (N_2911,N_2173,N_1895);
xor U2912 (N_2912,N_1934,N_2217);
xor U2913 (N_2913,N_2306,N_2132);
and U2914 (N_2914,N_2150,N_2032);
nand U2915 (N_2915,N_2037,N_2199);
xnor U2916 (N_2916,N_1919,N_2344);
xor U2917 (N_2917,N_2055,N_1809);
nand U2918 (N_2918,N_1991,N_2209);
nor U2919 (N_2919,N_2189,N_1895);
nand U2920 (N_2920,N_2052,N_2339);
nand U2921 (N_2921,N_2230,N_2004);
nor U2922 (N_2922,N_1803,N_2023);
or U2923 (N_2923,N_2177,N_2304);
and U2924 (N_2924,N_1860,N_1837);
nor U2925 (N_2925,N_1824,N_1908);
nor U2926 (N_2926,N_1821,N_2195);
nor U2927 (N_2927,N_2062,N_2365);
xnor U2928 (N_2928,N_2137,N_2133);
xnor U2929 (N_2929,N_2285,N_2040);
xor U2930 (N_2930,N_2311,N_1851);
or U2931 (N_2931,N_2271,N_2096);
or U2932 (N_2932,N_2145,N_2043);
nor U2933 (N_2933,N_1823,N_2399);
and U2934 (N_2934,N_2283,N_2337);
xor U2935 (N_2935,N_1800,N_2125);
nand U2936 (N_2936,N_2330,N_2216);
xnor U2937 (N_2937,N_2151,N_1829);
nand U2938 (N_2938,N_2025,N_2021);
and U2939 (N_2939,N_2306,N_1853);
nand U2940 (N_2940,N_1931,N_2143);
or U2941 (N_2941,N_2024,N_2147);
nor U2942 (N_2942,N_1806,N_2266);
nand U2943 (N_2943,N_1948,N_2114);
nor U2944 (N_2944,N_1872,N_2211);
and U2945 (N_2945,N_2058,N_2191);
or U2946 (N_2946,N_2337,N_2392);
or U2947 (N_2947,N_2246,N_1980);
xnor U2948 (N_2948,N_2309,N_1907);
nor U2949 (N_2949,N_2340,N_2209);
nand U2950 (N_2950,N_2092,N_1802);
and U2951 (N_2951,N_1869,N_2299);
and U2952 (N_2952,N_2306,N_1991);
or U2953 (N_2953,N_2234,N_2362);
or U2954 (N_2954,N_2031,N_1933);
xor U2955 (N_2955,N_1807,N_1979);
xnor U2956 (N_2956,N_1829,N_1827);
or U2957 (N_2957,N_2196,N_2199);
or U2958 (N_2958,N_2242,N_2284);
xnor U2959 (N_2959,N_1942,N_2133);
xnor U2960 (N_2960,N_2073,N_2224);
or U2961 (N_2961,N_2246,N_2328);
nand U2962 (N_2962,N_2286,N_2226);
xor U2963 (N_2963,N_2001,N_2159);
or U2964 (N_2964,N_2331,N_1980);
or U2965 (N_2965,N_2115,N_2216);
and U2966 (N_2966,N_2246,N_2270);
xor U2967 (N_2967,N_2019,N_2227);
nand U2968 (N_2968,N_2148,N_1944);
nor U2969 (N_2969,N_2102,N_1804);
or U2970 (N_2970,N_1935,N_1985);
and U2971 (N_2971,N_2164,N_2180);
or U2972 (N_2972,N_2015,N_1948);
nand U2973 (N_2973,N_2250,N_2028);
xor U2974 (N_2974,N_1800,N_2059);
xnor U2975 (N_2975,N_1909,N_2205);
and U2976 (N_2976,N_1935,N_2114);
nor U2977 (N_2977,N_2261,N_2213);
xor U2978 (N_2978,N_1992,N_2189);
nand U2979 (N_2979,N_1899,N_2161);
nand U2980 (N_2980,N_2241,N_2224);
nor U2981 (N_2981,N_2207,N_2011);
xnor U2982 (N_2982,N_1832,N_1856);
nand U2983 (N_2983,N_1807,N_2272);
nand U2984 (N_2984,N_2099,N_1863);
xor U2985 (N_2985,N_1974,N_2363);
nor U2986 (N_2986,N_2170,N_2163);
or U2987 (N_2987,N_2042,N_2123);
and U2988 (N_2988,N_1801,N_1961);
nor U2989 (N_2989,N_2174,N_2066);
or U2990 (N_2990,N_2211,N_2149);
nor U2991 (N_2991,N_2043,N_2033);
nand U2992 (N_2992,N_2084,N_1878);
or U2993 (N_2993,N_2011,N_1929);
nor U2994 (N_2994,N_1931,N_1930);
and U2995 (N_2995,N_2259,N_2378);
nand U2996 (N_2996,N_1942,N_2288);
nand U2997 (N_2997,N_2346,N_2096);
and U2998 (N_2998,N_1854,N_1822);
or U2999 (N_2999,N_1931,N_2094);
nand U3000 (N_3000,N_2951,N_2883);
xnor U3001 (N_3001,N_2434,N_2522);
nand U3002 (N_3002,N_2449,N_2657);
nand U3003 (N_3003,N_2581,N_2727);
nor U3004 (N_3004,N_2945,N_2811);
xor U3005 (N_3005,N_2898,N_2903);
nor U3006 (N_3006,N_2450,N_2674);
xnor U3007 (N_3007,N_2567,N_2623);
nor U3008 (N_3008,N_2912,N_2768);
xnor U3009 (N_3009,N_2471,N_2443);
xor U3010 (N_3010,N_2534,N_2608);
and U3011 (N_3011,N_2855,N_2685);
or U3012 (N_3012,N_2654,N_2720);
or U3013 (N_3013,N_2592,N_2820);
and U3014 (N_3014,N_2762,N_2920);
or U3015 (N_3015,N_2829,N_2607);
xor U3016 (N_3016,N_2761,N_2990);
xnor U3017 (N_3017,N_2813,N_2456);
nor U3018 (N_3018,N_2459,N_2454);
xor U3019 (N_3019,N_2462,N_2864);
or U3020 (N_3020,N_2564,N_2747);
xor U3021 (N_3021,N_2474,N_2796);
and U3022 (N_3022,N_2957,N_2644);
or U3023 (N_3023,N_2691,N_2642);
and U3024 (N_3024,N_2987,N_2435);
and U3025 (N_3025,N_2686,N_2639);
nor U3026 (N_3026,N_2599,N_2514);
and U3027 (N_3027,N_2809,N_2986);
nor U3028 (N_3028,N_2413,N_2615);
nor U3029 (N_3029,N_2563,N_2844);
nor U3030 (N_3030,N_2962,N_2453);
xor U3031 (N_3031,N_2724,N_2437);
nand U3032 (N_3032,N_2753,N_2881);
xor U3033 (N_3033,N_2910,N_2847);
or U3034 (N_3034,N_2426,N_2465);
xor U3035 (N_3035,N_2635,N_2513);
xor U3036 (N_3036,N_2925,N_2452);
xnor U3037 (N_3037,N_2839,N_2963);
nor U3038 (N_3038,N_2973,N_2786);
nor U3039 (N_3039,N_2626,N_2735);
or U3040 (N_3040,N_2767,N_2923);
and U3041 (N_3041,N_2680,N_2841);
or U3042 (N_3042,N_2542,N_2823);
nand U3043 (N_3043,N_2784,N_2979);
nand U3044 (N_3044,N_2613,N_2645);
nand U3045 (N_3045,N_2827,N_2492);
nor U3046 (N_3046,N_2417,N_2464);
and U3047 (N_3047,N_2602,N_2916);
nand U3048 (N_3048,N_2715,N_2414);
nand U3049 (N_3049,N_2968,N_2650);
or U3050 (N_3050,N_2947,N_2476);
or U3051 (N_3051,N_2693,N_2953);
or U3052 (N_3052,N_2928,N_2905);
nand U3053 (N_3053,N_2653,N_2935);
and U3054 (N_3054,N_2755,N_2890);
nor U3055 (N_3055,N_2914,N_2909);
and U3056 (N_3056,N_2868,N_2942);
and U3057 (N_3057,N_2853,N_2984);
and U3058 (N_3058,N_2468,N_2852);
nand U3059 (N_3059,N_2477,N_2529);
or U3060 (N_3060,N_2961,N_2489);
nand U3061 (N_3061,N_2588,N_2577);
and U3062 (N_3062,N_2954,N_2763);
and U3063 (N_3063,N_2965,N_2511);
nor U3064 (N_3064,N_2992,N_2931);
nor U3065 (N_3065,N_2774,N_2901);
nor U3066 (N_3066,N_2836,N_2833);
and U3067 (N_3067,N_2593,N_2779);
xnor U3068 (N_3068,N_2463,N_2550);
and U3069 (N_3069,N_2988,N_2889);
or U3070 (N_3070,N_2746,N_2738);
nor U3071 (N_3071,N_2663,N_2533);
and U3072 (N_3072,N_2643,N_2950);
or U3073 (N_3073,N_2669,N_2525);
and U3074 (N_3074,N_2991,N_2557);
nor U3075 (N_3075,N_2817,N_2497);
nor U3076 (N_3076,N_2749,N_2573);
xor U3077 (N_3077,N_2980,N_2740);
nor U3078 (N_3078,N_2505,N_2444);
xor U3079 (N_3079,N_2771,N_2553);
or U3080 (N_3080,N_2407,N_2457);
or U3081 (N_3081,N_2429,N_2978);
and U3082 (N_3082,N_2467,N_2496);
xor U3083 (N_3083,N_2851,N_2981);
and U3084 (N_3084,N_2830,N_2696);
or U3085 (N_3085,N_2876,N_2554);
or U3086 (N_3086,N_2598,N_2636);
and U3087 (N_3087,N_2741,N_2846);
nor U3088 (N_3088,N_2549,N_2911);
nand U3089 (N_3089,N_2859,N_2586);
nand U3090 (N_3090,N_2939,N_2568);
nand U3091 (N_3091,N_2617,N_2430);
nand U3092 (N_3092,N_2587,N_2624);
nor U3093 (N_3093,N_2926,N_2930);
and U3094 (N_3094,N_2879,N_2486);
xor U3095 (N_3095,N_2997,N_2656);
nor U3096 (N_3096,N_2538,N_2871);
nor U3097 (N_3097,N_2610,N_2956);
nand U3098 (N_3098,N_2484,N_2678);
nor U3099 (N_3099,N_2424,N_2507);
or U3100 (N_3100,N_2932,N_2714);
nor U3101 (N_3101,N_2500,N_2673);
or U3102 (N_3102,N_2527,N_2433);
xnor U3103 (N_3103,N_2810,N_2485);
and U3104 (N_3104,N_2619,N_2744);
xor U3105 (N_3105,N_2439,N_2488);
and U3106 (N_3106,N_2819,N_2479);
xor U3107 (N_3107,N_2604,N_2532);
nand U3108 (N_3108,N_2498,N_2662);
nand U3109 (N_3109,N_2493,N_2949);
or U3110 (N_3110,N_2828,N_2758);
nor U3111 (N_3111,N_2616,N_2440);
nand U3112 (N_3112,N_2929,N_2770);
nor U3113 (N_3113,N_2428,N_2442);
or U3114 (N_3114,N_2585,N_2700);
nor U3115 (N_3115,N_2825,N_2712);
nor U3116 (N_3116,N_2952,N_2732);
nor U3117 (N_3117,N_2789,N_2897);
xor U3118 (N_3118,N_2609,N_2475);
xor U3119 (N_3119,N_2873,N_2652);
nand U3120 (N_3120,N_2702,N_2606);
xnor U3121 (N_3121,N_2405,N_2692);
and U3122 (N_3122,N_2551,N_2821);
or U3123 (N_3123,N_2870,N_2861);
or U3124 (N_3124,N_2423,N_2967);
nand U3125 (N_3125,N_2793,N_2941);
xnor U3126 (N_3126,N_2893,N_2756);
nand U3127 (N_3127,N_2989,N_2526);
or U3128 (N_3128,N_2600,N_2971);
nor U3129 (N_3129,N_2638,N_2863);
nand U3130 (N_3130,N_2541,N_2869);
or U3131 (N_3131,N_2412,N_2518);
or U3132 (N_3132,N_2483,N_2765);
xnor U3133 (N_3133,N_2797,N_2614);
and U3134 (N_3134,N_2546,N_2591);
nand U3135 (N_3135,N_2832,N_2713);
or U3136 (N_3136,N_2848,N_2955);
or U3137 (N_3137,N_2690,N_2427);
nand U3138 (N_3138,N_2575,N_2629);
nor U3139 (N_3139,N_2561,N_2802);
and U3140 (N_3140,N_2535,N_2537);
nand U3141 (N_3141,N_2733,N_2502);
nor U3142 (N_3142,N_2687,N_2743);
nand U3143 (N_3143,N_2640,N_2540);
nand U3144 (N_3144,N_2469,N_2865);
and U3145 (N_3145,N_2734,N_2804);
xor U3146 (N_3146,N_2566,N_2775);
xnor U3147 (N_3147,N_2676,N_2637);
nor U3148 (N_3148,N_2785,N_2501);
nand U3149 (N_3149,N_2432,N_2545);
nand U3150 (N_3150,N_2976,N_2706);
or U3151 (N_3151,N_2583,N_2408);
and U3152 (N_3152,N_2547,N_2709);
and U3153 (N_3153,N_2704,N_2866);
nand U3154 (N_3154,N_2737,N_2900);
nand U3155 (N_3155,N_2603,N_2622);
nand U3156 (N_3156,N_2748,N_2915);
nand U3157 (N_3157,N_2560,N_2421);
nor U3158 (N_3158,N_2933,N_2699);
nand U3159 (N_3159,N_2887,N_2504);
and U3160 (N_3160,N_2728,N_2831);
or U3161 (N_3161,N_2751,N_2875);
nand U3162 (N_3162,N_2778,N_2888);
xnor U3163 (N_3163,N_2896,N_2975);
nand U3164 (N_3164,N_2460,N_2589);
nor U3165 (N_3165,N_2966,N_2499);
xnor U3166 (N_3166,N_2794,N_2618);
or U3167 (N_3167,N_2999,N_2630);
or U3168 (N_3168,N_2491,N_2441);
or U3169 (N_3169,N_2461,N_2760);
nand U3170 (N_3170,N_2482,N_2596);
nand U3171 (N_3171,N_2904,N_2776);
xnor U3172 (N_3172,N_2729,N_2739);
and U3173 (N_3173,N_2725,N_2531);
nand U3174 (N_3174,N_2985,N_2574);
xor U3175 (N_3175,N_2446,N_2695);
nor U3176 (N_3176,N_2509,N_2816);
xnor U3177 (N_3177,N_2882,N_2899);
nand U3178 (N_3178,N_2548,N_2647);
and U3179 (N_3179,N_2944,N_2788);
nor U3180 (N_3180,N_2917,N_2982);
xnor U3181 (N_3181,N_2675,N_2523);
or U3182 (N_3182,N_2908,N_2854);
xor U3183 (N_3183,N_2969,N_2641);
and U3184 (N_3184,N_2922,N_2711);
xnor U3185 (N_3185,N_2555,N_2708);
and U3186 (N_3186,N_2777,N_2448);
nand U3187 (N_3187,N_2977,N_2891);
xor U3188 (N_3188,N_2536,N_2480);
xor U3189 (N_3189,N_2672,N_2666);
nor U3190 (N_3190,N_2668,N_2661);
nand U3191 (N_3191,N_2694,N_2487);
and U3192 (N_3192,N_2582,N_2838);
and U3193 (N_3193,N_2438,N_2418);
nand U3194 (N_3194,N_2632,N_2562);
nor U3195 (N_3195,N_2840,N_2716);
nor U3196 (N_3196,N_2472,N_2835);
nand U3197 (N_3197,N_2478,N_2572);
or U3198 (N_3198,N_2697,N_2579);
nor U3199 (N_3199,N_2422,N_2934);
xor U3200 (N_3200,N_2558,N_2913);
nand U3201 (N_3201,N_2812,N_2894);
nor U3202 (N_3202,N_2565,N_2402);
nand U3203 (N_3203,N_2425,N_2808);
or U3204 (N_3204,N_2906,N_2959);
nand U3205 (N_3205,N_2570,N_2850);
or U3206 (N_3206,N_2946,N_2791);
and U3207 (N_3207,N_2721,N_2938);
nor U3208 (N_3208,N_2494,N_2877);
and U3209 (N_3209,N_2936,N_2818);
nor U3210 (N_3210,N_2921,N_2837);
and U3211 (N_3211,N_2458,N_2845);
nand U3212 (N_3212,N_2544,N_2506);
nand U3213 (N_3213,N_2803,N_2958);
nand U3214 (N_3214,N_2764,N_2658);
nor U3215 (N_3215,N_2406,N_2431);
and U3216 (N_3216,N_2798,N_2718);
nor U3217 (N_3217,N_2508,N_2569);
nand U3218 (N_3218,N_2872,N_2769);
nor U3219 (N_3219,N_2528,N_2948);
or U3220 (N_3220,N_2634,N_2578);
nand U3221 (N_3221,N_2404,N_2717);
or U3222 (N_3222,N_2445,N_2689);
and U3223 (N_3223,N_2736,N_2726);
nand U3224 (N_3224,N_2670,N_2473);
xor U3225 (N_3225,N_2655,N_2605);
or U3226 (N_3226,N_2495,N_2862);
nand U3227 (N_3227,N_2772,N_2671);
nand U3228 (N_3228,N_2842,N_2648);
xnor U3229 (N_3229,N_2843,N_2520);
and U3230 (N_3230,N_2665,N_2517);
nand U3231 (N_3231,N_2415,N_2594);
nand U3232 (N_3232,N_2400,N_2684);
nor U3233 (N_3233,N_2805,N_2539);
nor U3234 (N_3234,N_2892,N_2710);
or U3235 (N_3235,N_2651,N_2664);
nor U3236 (N_3236,N_2927,N_2974);
nand U3237 (N_3237,N_2874,N_2503);
nor U3238 (N_3238,N_2681,N_2612);
or U3239 (N_3239,N_2682,N_2886);
or U3240 (N_3240,N_2705,N_2807);
and U3241 (N_3241,N_2860,N_2795);
nand U3242 (N_3242,N_2742,N_2679);
xor U3243 (N_3243,N_2409,N_2722);
nand U3244 (N_3244,N_2515,N_2822);
and U3245 (N_3245,N_2576,N_2983);
nand U3246 (N_3246,N_2683,N_2701);
xor U3247 (N_3247,N_2416,N_2521);
xnor U3248 (N_3248,N_2996,N_2937);
nor U3249 (N_3249,N_2436,N_2698);
and U3250 (N_3250,N_2516,N_2918);
or U3251 (N_3251,N_2590,N_2780);
and U3252 (N_3252,N_2620,N_2878);
xor U3253 (N_3253,N_2824,N_2419);
nor U3254 (N_3254,N_2754,N_2806);
nor U3255 (N_3255,N_2907,N_2943);
nand U3256 (N_3256,N_2597,N_2451);
xor U3257 (N_3257,N_2857,N_2885);
nand U3258 (N_3258,N_2601,N_2660);
nor U3259 (N_3259,N_2752,N_2703);
nand U3260 (N_3260,N_2783,N_2649);
or U3261 (N_3261,N_2970,N_2834);
xor U3262 (N_3262,N_2571,N_2552);
and U3263 (N_3263,N_2584,N_2800);
xnor U3264 (N_3264,N_2447,N_2902);
nor U3265 (N_3265,N_2646,N_2995);
nand U3266 (N_3266,N_2543,N_2455);
xor U3267 (N_3267,N_2611,N_2633);
or U3268 (N_3268,N_2972,N_2964);
and U3269 (N_3269,N_2677,N_2858);
or U3270 (N_3270,N_2401,N_2814);
nor U3271 (N_3271,N_2627,N_2998);
nor U3272 (N_3272,N_2512,N_2659);
or U3273 (N_3273,N_2826,N_2667);
xnor U3274 (N_3274,N_2688,N_2707);
xnor U3275 (N_3275,N_2559,N_2792);
nor U3276 (N_3276,N_2750,N_2867);
nor U3277 (N_3277,N_2524,N_2766);
xor U3278 (N_3278,N_2787,N_2730);
xnor U3279 (N_3279,N_2919,N_2884);
or U3280 (N_3280,N_2745,N_2940);
nand U3281 (N_3281,N_2781,N_2519);
or U3282 (N_3282,N_2410,N_2723);
and U3283 (N_3283,N_2490,N_2470);
nand U3284 (N_3284,N_2924,N_2481);
or U3285 (N_3285,N_2759,N_2420);
nand U3286 (N_3286,N_2773,N_2993);
xnor U3287 (N_3287,N_2719,N_2790);
and U3288 (N_3288,N_2556,N_2595);
and U3289 (N_3289,N_2895,N_2621);
xor U3290 (N_3290,N_2782,N_2403);
and U3291 (N_3291,N_2960,N_2631);
nand U3292 (N_3292,N_2510,N_2799);
xor U3293 (N_3293,N_2757,N_2994);
and U3294 (N_3294,N_2815,N_2530);
nand U3295 (N_3295,N_2466,N_2625);
xor U3296 (N_3296,N_2801,N_2856);
nor U3297 (N_3297,N_2411,N_2849);
xor U3298 (N_3298,N_2731,N_2628);
nor U3299 (N_3299,N_2880,N_2580);
and U3300 (N_3300,N_2522,N_2919);
or U3301 (N_3301,N_2842,N_2510);
or U3302 (N_3302,N_2651,N_2723);
xnor U3303 (N_3303,N_2987,N_2818);
or U3304 (N_3304,N_2691,N_2460);
and U3305 (N_3305,N_2910,N_2892);
xnor U3306 (N_3306,N_2822,N_2836);
nor U3307 (N_3307,N_2778,N_2883);
nor U3308 (N_3308,N_2511,N_2990);
xor U3309 (N_3309,N_2737,N_2823);
nor U3310 (N_3310,N_2435,N_2467);
nor U3311 (N_3311,N_2924,N_2726);
or U3312 (N_3312,N_2862,N_2750);
xor U3313 (N_3313,N_2617,N_2436);
xor U3314 (N_3314,N_2502,N_2661);
xor U3315 (N_3315,N_2931,N_2733);
or U3316 (N_3316,N_2668,N_2489);
nand U3317 (N_3317,N_2529,N_2676);
nand U3318 (N_3318,N_2752,N_2597);
or U3319 (N_3319,N_2503,N_2625);
or U3320 (N_3320,N_2989,N_2724);
and U3321 (N_3321,N_2561,N_2826);
nor U3322 (N_3322,N_2450,N_2492);
nand U3323 (N_3323,N_2992,N_2704);
xnor U3324 (N_3324,N_2727,N_2508);
or U3325 (N_3325,N_2586,N_2793);
and U3326 (N_3326,N_2895,N_2637);
xor U3327 (N_3327,N_2928,N_2687);
xnor U3328 (N_3328,N_2643,N_2699);
or U3329 (N_3329,N_2537,N_2570);
and U3330 (N_3330,N_2573,N_2465);
xor U3331 (N_3331,N_2624,N_2880);
or U3332 (N_3332,N_2423,N_2534);
and U3333 (N_3333,N_2922,N_2408);
nand U3334 (N_3334,N_2725,N_2604);
and U3335 (N_3335,N_2885,N_2728);
or U3336 (N_3336,N_2748,N_2403);
and U3337 (N_3337,N_2999,N_2719);
and U3338 (N_3338,N_2564,N_2693);
and U3339 (N_3339,N_2803,N_2529);
nor U3340 (N_3340,N_2761,N_2533);
nand U3341 (N_3341,N_2772,N_2490);
and U3342 (N_3342,N_2594,N_2584);
and U3343 (N_3343,N_2583,N_2422);
nor U3344 (N_3344,N_2429,N_2869);
xnor U3345 (N_3345,N_2793,N_2756);
nor U3346 (N_3346,N_2931,N_2689);
or U3347 (N_3347,N_2760,N_2534);
nor U3348 (N_3348,N_2546,N_2897);
nand U3349 (N_3349,N_2980,N_2979);
nor U3350 (N_3350,N_2546,N_2845);
or U3351 (N_3351,N_2985,N_2986);
xnor U3352 (N_3352,N_2453,N_2933);
or U3353 (N_3353,N_2719,N_2513);
nand U3354 (N_3354,N_2414,N_2766);
and U3355 (N_3355,N_2620,N_2725);
xnor U3356 (N_3356,N_2563,N_2574);
or U3357 (N_3357,N_2984,N_2687);
xor U3358 (N_3358,N_2508,N_2421);
and U3359 (N_3359,N_2442,N_2970);
nand U3360 (N_3360,N_2920,N_2442);
and U3361 (N_3361,N_2954,N_2583);
and U3362 (N_3362,N_2433,N_2797);
or U3363 (N_3363,N_2662,N_2617);
or U3364 (N_3364,N_2821,N_2876);
nor U3365 (N_3365,N_2576,N_2488);
nand U3366 (N_3366,N_2733,N_2471);
nand U3367 (N_3367,N_2565,N_2905);
nor U3368 (N_3368,N_2560,N_2794);
or U3369 (N_3369,N_2934,N_2997);
and U3370 (N_3370,N_2470,N_2925);
or U3371 (N_3371,N_2679,N_2591);
and U3372 (N_3372,N_2838,N_2572);
xnor U3373 (N_3373,N_2838,N_2923);
and U3374 (N_3374,N_2885,N_2803);
or U3375 (N_3375,N_2949,N_2523);
and U3376 (N_3376,N_2966,N_2842);
or U3377 (N_3377,N_2818,N_2459);
xnor U3378 (N_3378,N_2830,N_2559);
xor U3379 (N_3379,N_2571,N_2753);
nor U3380 (N_3380,N_2462,N_2674);
xor U3381 (N_3381,N_2787,N_2697);
nor U3382 (N_3382,N_2954,N_2631);
or U3383 (N_3383,N_2973,N_2763);
nand U3384 (N_3384,N_2642,N_2958);
nand U3385 (N_3385,N_2667,N_2460);
xor U3386 (N_3386,N_2615,N_2547);
xor U3387 (N_3387,N_2921,N_2749);
or U3388 (N_3388,N_2679,N_2921);
or U3389 (N_3389,N_2643,N_2958);
or U3390 (N_3390,N_2827,N_2604);
and U3391 (N_3391,N_2484,N_2606);
nor U3392 (N_3392,N_2832,N_2963);
or U3393 (N_3393,N_2611,N_2465);
and U3394 (N_3394,N_2932,N_2538);
or U3395 (N_3395,N_2931,N_2451);
or U3396 (N_3396,N_2564,N_2821);
xor U3397 (N_3397,N_2824,N_2742);
nor U3398 (N_3398,N_2841,N_2502);
nor U3399 (N_3399,N_2995,N_2796);
or U3400 (N_3400,N_2570,N_2560);
xnor U3401 (N_3401,N_2729,N_2523);
or U3402 (N_3402,N_2818,N_2646);
and U3403 (N_3403,N_2421,N_2923);
or U3404 (N_3404,N_2732,N_2864);
and U3405 (N_3405,N_2619,N_2655);
nand U3406 (N_3406,N_2724,N_2658);
and U3407 (N_3407,N_2489,N_2478);
nand U3408 (N_3408,N_2748,N_2665);
nor U3409 (N_3409,N_2810,N_2827);
nand U3410 (N_3410,N_2968,N_2832);
nor U3411 (N_3411,N_2892,N_2677);
nor U3412 (N_3412,N_2852,N_2770);
nor U3413 (N_3413,N_2439,N_2572);
or U3414 (N_3414,N_2678,N_2797);
nand U3415 (N_3415,N_2939,N_2517);
nand U3416 (N_3416,N_2653,N_2682);
xor U3417 (N_3417,N_2875,N_2843);
xnor U3418 (N_3418,N_2973,N_2700);
xnor U3419 (N_3419,N_2656,N_2545);
xor U3420 (N_3420,N_2547,N_2881);
nand U3421 (N_3421,N_2834,N_2637);
and U3422 (N_3422,N_2720,N_2476);
and U3423 (N_3423,N_2478,N_2672);
and U3424 (N_3424,N_2535,N_2488);
and U3425 (N_3425,N_2684,N_2867);
xor U3426 (N_3426,N_2745,N_2562);
or U3427 (N_3427,N_2620,N_2974);
nand U3428 (N_3428,N_2775,N_2771);
or U3429 (N_3429,N_2692,N_2796);
and U3430 (N_3430,N_2493,N_2917);
and U3431 (N_3431,N_2587,N_2601);
and U3432 (N_3432,N_2476,N_2936);
xnor U3433 (N_3433,N_2428,N_2922);
or U3434 (N_3434,N_2520,N_2833);
xor U3435 (N_3435,N_2771,N_2788);
or U3436 (N_3436,N_2839,N_2846);
and U3437 (N_3437,N_2694,N_2769);
xor U3438 (N_3438,N_2884,N_2731);
xor U3439 (N_3439,N_2513,N_2907);
xnor U3440 (N_3440,N_2427,N_2485);
xor U3441 (N_3441,N_2467,N_2629);
and U3442 (N_3442,N_2815,N_2459);
or U3443 (N_3443,N_2602,N_2644);
nor U3444 (N_3444,N_2723,N_2763);
xnor U3445 (N_3445,N_2726,N_2913);
nand U3446 (N_3446,N_2586,N_2595);
nor U3447 (N_3447,N_2928,N_2573);
and U3448 (N_3448,N_2709,N_2450);
nor U3449 (N_3449,N_2782,N_2897);
nand U3450 (N_3450,N_2767,N_2886);
or U3451 (N_3451,N_2706,N_2535);
xor U3452 (N_3452,N_2410,N_2810);
nor U3453 (N_3453,N_2675,N_2921);
nand U3454 (N_3454,N_2848,N_2779);
nand U3455 (N_3455,N_2617,N_2554);
nand U3456 (N_3456,N_2780,N_2771);
and U3457 (N_3457,N_2780,N_2603);
or U3458 (N_3458,N_2708,N_2410);
nor U3459 (N_3459,N_2527,N_2791);
or U3460 (N_3460,N_2659,N_2696);
xnor U3461 (N_3461,N_2619,N_2905);
nand U3462 (N_3462,N_2764,N_2781);
nand U3463 (N_3463,N_2499,N_2445);
nand U3464 (N_3464,N_2449,N_2727);
nand U3465 (N_3465,N_2799,N_2571);
or U3466 (N_3466,N_2589,N_2695);
xor U3467 (N_3467,N_2999,N_2455);
nor U3468 (N_3468,N_2583,N_2778);
nand U3469 (N_3469,N_2643,N_2602);
or U3470 (N_3470,N_2759,N_2635);
or U3471 (N_3471,N_2573,N_2407);
xnor U3472 (N_3472,N_2918,N_2795);
nand U3473 (N_3473,N_2686,N_2935);
or U3474 (N_3474,N_2588,N_2987);
and U3475 (N_3475,N_2977,N_2795);
and U3476 (N_3476,N_2795,N_2420);
nand U3477 (N_3477,N_2567,N_2552);
nor U3478 (N_3478,N_2846,N_2584);
nand U3479 (N_3479,N_2627,N_2583);
nand U3480 (N_3480,N_2853,N_2551);
or U3481 (N_3481,N_2847,N_2684);
nor U3482 (N_3482,N_2702,N_2842);
or U3483 (N_3483,N_2941,N_2847);
or U3484 (N_3484,N_2479,N_2816);
nand U3485 (N_3485,N_2974,N_2657);
or U3486 (N_3486,N_2916,N_2627);
nand U3487 (N_3487,N_2573,N_2524);
xor U3488 (N_3488,N_2926,N_2771);
or U3489 (N_3489,N_2474,N_2891);
nor U3490 (N_3490,N_2581,N_2710);
or U3491 (N_3491,N_2549,N_2762);
and U3492 (N_3492,N_2660,N_2912);
nor U3493 (N_3493,N_2776,N_2468);
nor U3494 (N_3494,N_2640,N_2850);
and U3495 (N_3495,N_2845,N_2928);
xnor U3496 (N_3496,N_2996,N_2429);
and U3497 (N_3497,N_2772,N_2794);
nor U3498 (N_3498,N_2580,N_2473);
xor U3499 (N_3499,N_2696,N_2523);
nand U3500 (N_3500,N_2677,N_2540);
nor U3501 (N_3501,N_2517,N_2884);
xor U3502 (N_3502,N_2852,N_2564);
or U3503 (N_3503,N_2431,N_2777);
or U3504 (N_3504,N_2877,N_2754);
xor U3505 (N_3505,N_2408,N_2836);
xnor U3506 (N_3506,N_2921,N_2515);
nand U3507 (N_3507,N_2661,N_2982);
or U3508 (N_3508,N_2930,N_2556);
and U3509 (N_3509,N_2668,N_2791);
or U3510 (N_3510,N_2913,N_2711);
or U3511 (N_3511,N_2526,N_2971);
nand U3512 (N_3512,N_2545,N_2414);
nor U3513 (N_3513,N_2410,N_2492);
or U3514 (N_3514,N_2743,N_2558);
nor U3515 (N_3515,N_2784,N_2704);
xor U3516 (N_3516,N_2783,N_2631);
and U3517 (N_3517,N_2427,N_2590);
nand U3518 (N_3518,N_2922,N_2456);
and U3519 (N_3519,N_2559,N_2400);
xor U3520 (N_3520,N_2485,N_2791);
or U3521 (N_3521,N_2462,N_2616);
or U3522 (N_3522,N_2629,N_2920);
nor U3523 (N_3523,N_2714,N_2419);
nor U3524 (N_3524,N_2883,N_2416);
or U3525 (N_3525,N_2761,N_2958);
xnor U3526 (N_3526,N_2737,N_2789);
nor U3527 (N_3527,N_2822,N_2575);
or U3528 (N_3528,N_2464,N_2528);
nand U3529 (N_3529,N_2763,N_2545);
or U3530 (N_3530,N_2440,N_2516);
xnor U3531 (N_3531,N_2970,N_2603);
nor U3532 (N_3532,N_2789,N_2955);
and U3533 (N_3533,N_2759,N_2693);
and U3534 (N_3534,N_2739,N_2590);
or U3535 (N_3535,N_2678,N_2558);
or U3536 (N_3536,N_2540,N_2744);
xnor U3537 (N_3537,N_2893,N_2763);
and U3538 (N_3538,N_2425,N_2702);
nor U3539 (N_3539,N_2704,N_2856);
nor U3540 (N_3540,N_2446,N_2610);
nor U3541 (N_3541,N_2452,N_2421);
xor U3542 (N_3542,N_2789,N_2976);
nor U3543 (N_3543,N_2768,N_2561);
nand U3544 (N_3544,N_2650,N_2819);
nand U3545 (N_3545,N_2882,N_2809);
and U3546 (N_3546,N_2508,N_2499);
nor U3547 (N_3547,N_2784,N_2701);
xnor U3548 (N_3548,N_2956,N_2837);
nand U3549 (N_3549,N_2463,N_2754);
and U3550 (N_3550,N_2779,N_2643);
or U3551 (N_3551,N_2529,N_2494);
and U3552 (N_3552,N_2687,N_2900);
or U3553 (N_3553,N_2571,N_2944);
or U3554 (N_3554,N_2566,N_2666);
and U3555 (N_3555,N_2568,N_2836);
xnor U3556 (N_3556,N_2996,N_2442);
nand U3557 (N_3557,N_2732,N_2637);
nor U3558 (N_3558,N_2860,N_2476);
xnor U3559 (N_3559,N_2824,N_2930);
or U3560 (N_3560,N_2784,N_2461);
and U3561 (N_3561,N_2763,N_2745);
nand U3562 (N_3562,N_2488,N_2875);
or U3563 (N_3563,N_2693,N_2981);
nor U3564 (N_3564,N_2826,N_2745);
nand U3565 (N_3565,N_2457,N_2667);
nor U3566 (N_3566,N_2588,N_2759);
nor U3567 (N_3567,N_2673,N_2654);
nand U3568 (N_3568,N_2886,N_2881);
or U3569 (N_3569,N_2461,N_2418);
nor U3570 (N_3570,N_2427,N_2705);
nor U3571 (N_3571,N_2972,N_2673);
nor U3572 (N_3572,N_2591,N_2940);
and U3573 (N_3573,N_2722,N_2890);
xor U3574 (N_3574,N_2744,N_2556);
nor U3575 (N_3575,N_2915,N_2631);
nor U3576 (N_3576,N_2434,N_2904);
and U3577 (N_3577,N_2626,N_2541);
and U3578 (N_3578,N_2591,N_2481);
or U3579 (N_3579,N_2546,N_2427);
nand U3580 (N_3580,N_2562,N_2482);
or U3581 (N_3581,N_2991,N_2993);
nand U3582 (N_3582,N_2431,N_2427);
xnor U3583 (N_3583,N_2666,N_2688);
xnor U3584 (N_3584,N_2747,N_2600);
xor U3585 (N_3585,N_2407,N_2492);
or U3586 (N_3586,N_2951,N_2483);
and U3587 (N_3587,N_2439,N_2693);
and U3588 (N_3588,N_2648,N_2421);
xnor U3589 (N_3589,N_2979,N_2616);
and U3590 (N_3590,N_2500,N_2501);
nor U3591 (N_3591,N_2610,N_2830);
nor U3592 (N_3592,N_2802,N_2612);
nor U3593 (N_3593,N_2742,N_2958);
and U3594 (N_3594,N_2854,N_2939);
and U3595 (N_3595,N_2459,N_2507);
and U3596 (N_3596,N_2509,N_2427);
nand U3597 (N_3597,N_2501,N_2862);
nor U3598 (N_3598,N_2869,N_2849);
xor U3599 (N_3599,N_2646,N_2402);
and U3600 (N_3600,N_3373,N_3359);
nand U3601 (N_3601,N_3333,N_3048);
nand U3602 (N_3602,N_3232,N_3343);
nor U3603 (N_3603,N_3484,N_3397);
nand U3604 (N_3604,N_3086,N_3561);
xnor U3605 (N_3605,N_3241,N_3138);
xnor U3606 (N_3606,N_3012,N_3065);
and U3607 (N_3607,N_3572,N_3124);
nor U3608 (N_3608,N_3193,N_3275);
or U3609 (N_3609,N_3271,N_3510);
nand U3610 (N_3610,N_3418,N_3369);
nor U3611 (N_3611,N_3311,N_3464);
xnor U3612 (N_3612,N_3051,N_3229);
and U3613 (N_3613,N_3169,N_3254);
and U3614 (N_3614,N_3548,N_3570);
or U3615 (N_3615,N_3074,N_3030);
or U3616 (N_3616,N_3218,N_3262);
nand U3617 (N_3617,N_3263,N_3084);
or U3618 (N_3618,N_3095,N_3010);
xor U3619 (N_3619,N_3137,N_3072);
or U3620 (N_3620,N_3047,N_3270);
xnor U3621 (N_3621,N_3145,N_3059);
and U3622 (N_3622,N_3289,N_3123);
and U3623 (N_3623,N_3313,N_3211);
nor U3624 (N_3624,N_3290,N_3368);
nand U3625 (N_3625,N_3321,N_3535);
nor U3626 (N_3626,N_3214,N_3280);
nand U3627 (N_3627,N_3425,N_3136);
xnor U3628 (N_3628,N_3203,N_3285);
nor U3629 (N_3629,N_3399,N_3528);
or U3630 (N_3630,N_3175,N_3332);
nand U3631 (N_3631,N_3331,N_3268);
or U3632 (N_3632,N_3238,N_3101);
and U3633 (N_3633,N_3581,N_3341);
nand U3634 (N_3634,N_3436,N_3043);
nor U3635 (N_3635,N_3108,N_3213);
nand U3636 (N_3636,N_3549,N_3508);
xor U3637 (N_3637,N_3061,N_3093);
or U3638 (N_3638,N_3182,N_3122);
xor U3639 (N_3639,N_3252,N_3062);
nor U3640 (N_3640,N_3517,N_3091);
nor U3641 (N_3641,N_3015,N_3000);
nor U3642 (N_3642,N_3292,N_3477);
nand U3643 (N_3643,N_3109,N_3454);
and U3644 (N_3644,N_3345,N_3230);
nor U3645 (N_3645,N_3599,N_3562);
nand U3646 (N_3646,N_3547,N_3387);
xor U3647 (N_3647,N_3294,N_3512);
and U3648 (N_3648,N_3054,N_3307);
and U3649 (N_3649,N_3465,N_3557);
or U3650 (N_3650,N_3092,N_3105);
nor U3651 (N_3651,N_3117,N_3079);
nor U3652 (N_3652,N_3023,N_3318);
nor U3653 (N_3653,N_3001,N_3173);
or U3654 (N_3654,N_3494,N_3448);
or U3655 (N_3655,N_3468,N_3146);
and U3656 (N_3656,N_3440,N_3410);
xnor U3657 (N_3657,N_3550,N_3038);
nand U3658 (N_3658,N_3090,N_3305);
nor U3659 (N_3659,N_3041,N_3019);
or U3660 (N_3660,N_3140,N_3130);
nor U3661 (N_3661,N_3469,N_3080);
or U3662 (N_3662,N_3050,N_3488);
or U3663 (N_3663,N_3071,N_3427);
and U3664 (N_3664,N_3190,N_3304);
and U3665 (N_3665,N_3184,N_3049);
and U3666 (N_3666,N_3310,N_3330);
xnor U3667 (N_3667,N_3029,N_3404);
nor U3668 (N_3668,N_3513,N_3595);
and U3669 (N_3669,N_3301,N_3526);
xor U3670 (N_3670,N_3162,N_3206);
nand U3671 (N_3671,N_3185,N_3367);
or U3672 (N_3672,N_3361,N_3558);
nand U3673 (N_3673,N_3186,N_3007);
and U3674 (N_3674,N_3199,N_3174);
nor U3675 (N_3675,N_3246,N_3383);
nor U3676 (N_3676,N_3208,N_3461);
xnor U3677 (N_3677,N_3165,N_3258);
xor U3678 (N_3678,N_3155,N_3264);
and U3679 (N_3679,N_3594,N_3514);
or U3680 (N_3680,N_3302,N_3350);
nand U3681 (N_3681,N_3088,N_3422);
or U3682 (N_3682,N_3402,N_3243);
or U3683 (N_3683,N_3286,N_3445);
nand U3684 (N_3684,N_3125,N_3168);
nor U3685 (N_3685,N_3194,N_3196);
and U3686 (N_3686,N_3154,N_3308);
or U3687 (N_3687,N_3249,N_3014);
nand U3688 (N_3688,N_3348,N_3257);
and U3689 (N_3689,N_3351,N_3336);
nand U3690 (N_3690,N_3156,N_3297);
nand U3691 (N_3691,N_3273,N_3374);
nand U3692 (N_3692,N_3044,N_3344);
nand U3693 (N_3693,N_3278,N_3040);
or U3694 (N_3694,N_3008,N_3189);
nand U3695 (N_3695,N_3377,N_3157);
or U3696 (N_3696,N_3215,N_3272);
and U3697 (N_3697,N_3391,N_3167);
and U3698 (N_3698,N_3452,N_3543);
and U3699 (N_3699,N_3159,N_3544);
and U3700 (N_3700,N_3319,N_3151);
nand U3701 (N_3701,N_3586,N_3118);
xnor U3702 (N_3702,N_3565,N_3476);
nand U3703 (N_3703,N_3063,N_3166);
and U3704 (N_3704,N_3293,N_3085);
nand U3705 (N_3705,N_3417,N_3147);
nand U3706 (N_3706,N_3020,N_3375);
nor U3707 (N_3707,N_3180,N_3487);
nand U3708 (N_3708,N_3200,N_3385);
or U3709 (N_3709,N_3267,N_3106);
xor U3710 (N_3710,N_3300,N_3390);
nand U3711 (N_3711,N_3055,N_3354);
xor U3712 (N_3712,N_3531,N_3017);
or U3713 (N_3713,N_3111,N_3435);
or U3714 (N_3714,N_3409,N_3421);
xor U3715 (N_3715,N_3067,N_3335);
and U3716 (N_3716,N_3069,N_3120);
and U3717 (N_3717,N_3276,N_3068);
nor U3718 (N_3718,N_3400,N_3475);
or U3719 (N_3719,N_3027,N_3456);
xor U3720 (N_3720,N_3337,N_3161);
nor U3721 (N_3721,N_3392,N_3471);
nand U3722 (N_3722,N_3573,N_3314);
nand U3723 (N_3723,N_3433,N_3187);
nor U3724 (N_3724,N_3066,N_3009);
nand U3725 (N_3725,N_3450,N_3260);
nand U3726 (N_3726,N_3323,N_3378);
nand U3727 (N_3727,N_3303,N_3459);
nand U3728 (N_3728,N_3083,N_3149);
nand U3729 (N_3729,N_3470,N_3505);
nand U3730 (N_3730,N_3416,N_3371);
nor U3731 (N_3731,N_3281,N_3287);
nand U3732 (N_3732,N_3533,N_3515);
nand U3733 (N_3733,N_3220,N_3204);
nand U3734 (N_3734,N_3466,N_3447);
or U3735 (N_3735,N_3100,N_3366);
nand U3736 (N_3736,N_3455,N_3589);
and U3737 (N_3737,N_3004,N_3560);
nand U3738 (N_3738,N_3121,N_3474);
nor U3739 (N_3739,N_3247,N_3472);
xor U3740 (N_3740,N_3536,N_3462);
xnor U3741 (N_3741,N_3568,N_3128);
xnor U3742 (N_3742,N_3236,N_3396);
nand U3743 (N_3743,N_3362,N_3179);
and U3744 (N_3744,N_3315,N_3582);
and U3745 (N_3745,N_3401,N_3590);
or U3746 (N_3746,N_3207,N_3329);
nand U3747 (N_3747,N_3542,N_3546);
nand U3748 (N_3748,N_3235,N_3511);
nand U3749 (N_3749,N_3439,N_3002);
and U3750 (N_3750,N_3288,N_3250);
xor U3751 (N_3751,N_3210,N_3518);
xor U3752 (N_3752,N_3198,N_3143);
xor U3753 (N_3753,N_3496,N_3567);
and U3754 (N_3754,N_3274,N_3177);
nand U3755 (N_3755,N_3411,N_3089);
or U3756 (N_3756,N_3504,N_3265);
nand U3757 (N_3757,N_3324,N_3078);
or U3758 (N_3758,N_3357,N_3559);
or U3759 (N_3759,N_3490,N_3255);
nor U3760 (N_3760,N_3036,N_3132);
or U3761 (N_3761,N_3491,N_3114);
nor U3762 (N_3762,N_3192,N_3449);
or U3763 (N_3763,N_3394,N_3429);
or U3764 (N_3764,N_3405,N_3597);
and U3765 (N_3765,N_3003,N_3188);
or U3766 (N_3766,N_3160,N_3389);
or U3767 (N_3767,N_3356,N_3564);
nand U3768 (N_3768,N_3408,N_3413);
or U3769 (N_3769,N_3224,N_3591);
nand U3770 (N_3770,N_3058,N_3178);
xor U3771 (N_3771,N_3152,N_3501);
or U3772 (N_3772,N_3219,N_3493);
xnor U3773 (N_3773,N_3566,N_3588);
nor U3774 (N_3774,N_3284,N_3443);
xor U3775 (N_3775,N_3372,N_3463);
or U3776 (N_3776,N_3099,N_3516);
nor U3777 (N_3777,N_3395,N_3191);
nor U3778 (N_3778,N_3441,N_3056);
nor U3779 (N_3779,N_3453,N_3251);
nor U3780 (N_3780,N_3415,N_3347);
xnor U3781 (N_3781,N_3153,N_3028);
and U3782 (N_3782,N_3110,N_3098);
nor U3783 (N_3783,N_3212,N_3346);
nand U3784 (N_3784,N_3103,N_3025);
nand U3785 (N_3785,N_3529,N_3553);
nand U3786 (N_3786,N_3164,N_3525);
nand U3787 (N_3787,N_3340,N_3352);
xnor U3788 (N_3788,N_3242,N_3052);
and U3789 (N_3789,N_3438,N_3296);
or U3790 (N_3790,N_3502,N_3419);
nand U3791 (N_3791,N_3201,N_3306);
or U3792 (N_3792,N_3585,N_3370);
xor U3793 (N_3793,N_3139,N_3216);
nand U3794 (N_3794,N_3176,N_3571);
nor U3795 (N_3795,N_3593,N_3225);
nor U3796 (N_3796,N_3342,N_3171);
nor U3797 (N_3797,N_3320,N_3327);
nand U3798 (N_3798,N_3328,N_3498);
xor U3799 (N_3799,N_3231,N_3045);
nand U3800 (N_3800,N_3414,N_3298);
and U3801 (N_3801,N_3442,N_3024);
nor U3802 (N_3802,N_3388,N_3217);
and U3803 (N_3803,N_3202,N_3485);
and U3804 (N_3804,N_3349,N_3506);
nand U3805 (N_3805,N_3282,N_3011);
or U3806 (N_3806,N_3382,N_3077);
and U3807 (N_3807,N_3432,N_3393);
or U3808 (N_3808,N_3579,N_3039);
and U3809 (N_3809,N_3584,N_3545);
nor U3810 (N_3810,N_3412,N_3150);
nor U3811 (N_3811,N_3424,N_3060);
or U3812 (N_3812,N_3384,N_3587);
and U3813 (N_3813,N_3540,N_3205);
nor U3814 (N_3814,N_3037,N_3569);
or U3815 (N_3815,N_3523,N_3234);
nand U3816 (N_3816,N_3142,N_3181);
xnor U3817 (N_3817,N_3119,N_3530);
xnor U3818 (N_3818,N_3042,N_3163);
nand U3819 (N_3819,N_3478,N_3596);
and U3820 (N_3820,N_3133,N_3102);
xnor U3821 (N_3821,N_3221,N_3222);
and U3822 (N_3822,N_3021,N_3053);
nand U3823 (N_3823,N_3299,N_3034);
or U3824 (N_3824,N_3428,N_3134);
xnor U3825 (N_3825,N_3261,N_3295);
and U3826 (N_3826,N_3407,N_3483);
nand U3827 (N_3827,N_3376,N_3227);
nand U3828 (N_3828,N_3426,N_3519);
or U3829 (N_3829,N_3073,N_3170);
and U3830 (N_3830,N_3446,N_3495);
nand U3831 (N_3831,N_3075,N_3482);
nand U3832 (N_3832,N_3598,N_3148);
or U3833 (N_3833,N_3226,N_3026);
nor U3834 (N_3834,N_3195,N_3437);
and U3835 (N_3835,N_3183,N_3116);
nor U3836 (N_3836,N_3228,N_3420);
nand U3837 (N_3837,N_3578,N_3430);
and U3838 (N_3838,N_3334,N_3423);
and U3839 (N_3839,N_3094,N_3312);
and U3840 (N_3840,N_3309,N_3097);
xor U3841 (N_3841,N_3458,N_3035);
nor U3842 (N_3842,N_3339,N_3279);
and U3843 (N_3843,N_3580,N_3005);
or U3844 (N_3844,N_3431,N_3380);
or U3845 (N_3845,N_3554,N_3500);
nand U3846 (N_3846,N_3057,N_3358);
xnor U3847 (N_3847,N_3209,N_3244);
and U3848 (N_3848,N_3381,N_3325);
nand U3849 (N_3849,N_3135,N_3046);
or U3850 (N_3850,N_3457,N_3522);
xor U3851 (N_3851,N_3406,N_3239);
or U3852 (N_3852,N_3509,N_3486);
nor U3853 (N_3853,N_3006,N_3365);
and U3854 (N_3854,N_3338,N_3363);
nand U3855 (N_3855,N_3016,N_3480);
nand U3856 (N_3856,N_3444,N_3115);
nor U3857 (N_3857,N_3556,N_3256);
and U3858 (N_3858,N_3489,N_3364);
nand U3859 (N_3859,N_3022,N_3551);
or U3860 (N_3860,N_3592,N_3266);
nand U3861 (N_3861,N_3576,N_3492);
nor U3862 (N_3862,N_3322,N_3031);
or U3863 (N_3863,N_3233,N_3112);
xnor U3864 (N_3864,N_3481,N_3479);
xnor U3865 (N_3865,N_3538,N_3583);
or U3866 (N_3866,N_3141,N_3316);
xor U3867 (N_3867,N_3473,N_3240);
xnor U3868 (N_3868,N_3096,N_3563);
xnor U3869 (N_3869,N_3555,N_3317);
or U3870 (N_3870,N_3575,N_3434);
nor U3871 (N_3871,N_3237,N_3104);
nor U3872 (N_3872,N_3503,N_3532);
nand U3873 (N_3873,N_3277,N_3283);
or U3874 (N_3874,N_3087,N_3129);
nor U3875 (N_3875,N_3539,N_3520);
xor U3876 (N_3876,N_3013,N_3499);
or U3877 (N_3877,N_3534,N_3460);
nand U3878 (N_3878,N_3070,N_3259);
or U3879 (N_3879,N_3527,N_3064);
or U3880 (N_3880,N_3248,N_3126);
nor U3881 (N_3881,N_3032,N_3018);
nand U3882 (N_3882,N_3326,N_3082);
and U3883 (N_3883,N_3524,N_3552);
xor U3884 (N_3884,N_3467,N_3253);
xnor U3885 (N_3885,N_3269,N_3076);
nand U3886 (N_3886,N_3245,N_3541);
xor U3887 (N_3887,N_3081,N_3360);
or U3888 (N_3888,N_3113,N_3197);
and U3889 (N_3889,N_3107,N_3158);
xnor U3890 (N_3890,N_3379,N_3537);
and U3891 (N_3891,N_3574,N_3398);
xor U3892 (N_3892,N_3386,N_3403);
nor U3893 (N_3893,N_3127,N_3223);
nand U3894 (N_3894,N_3131,N_3144);
nor U3895 (N_3895,N_3521,N_3355);
and U3896 (N_3896,N_3451,N_3172);
xnor U3897 (N_3897,N_3353,N_3577);
nor U3898 (N_3898,N_3507,N_3291);
xnor U3899 (N_3899,N_3497,N_3033);
nand U3900 (N_3900,N_3313,N_3340);
nand U3901 (N_3901,N_3583,N_3271);
xnor U3902 (N_3902,N_3152,N_3469);
and U3903 (N_3903,N_3210,N_3147);
nand U3904 (N_3904,N_3328,N_3555);
nor U3905 (N_3905,N_3351,N_3489);
xnor U3906 (N_3906,N_3152,N_3252);
and U3907 (N_3907,N_3184,N_3160);
or U3908 (N_3908,N_3514,N_3565);
and U3909 (N_3909,N_3301,N_3066);
xor U3910 (N_3910,N_3327,N_3065);
nand U3911 (N_3911,N_3195,N_3288);
nor U3912 (N_3912,N_3202,N_3372);
nand U3913 (N_3913,N_3118,N_3198);
nand U3914 (N_3914,N_3296,N_3241);
nor U3915 (N_3915,N_3334,N_3360);
nand U3916 (N_3916,N_3000,N_3259);
and U3917 (N_3917,N_3598,N_3256);
nand U3918 (N_3918,N_3344,N_3530);
xor U3919 (N_3919,N_3394,N_3258);
xnor U3920 (N_3920,N_3125,N_3203);
xnor U3921 (N_3921,N_3100,N_3233);
nor U3922 (N_3922,N_3582,N_3062);
and U3923 (N_3923,N_3264,N_3330);
or U3924 (N_3924,N_3248,N_3148);
and U3925 (N_3925,N_3440,N_3260);
nor U3926 (N_3926,N_3592,N_3154);
xor U3927 (N_3927,N_3459,N_3291);
nand U3928 (N_3928,N_3326,N_3243);
and U3929 (N_3929,N_3375,N_3104);
nand U3930 (N_3930,N_3217,N_3408);
nor U3931 (N_3931,N_3081,N_3111);
or U3932 (N_3932,N_3256,N_3533);
and U3933 (N_3933,N_3059,N_3523);
and U3934 (N_3934,N_3350,N_3494);
xnor U3935 (N_3935,N_3371,N_3519);
nand U3936 (N_3936,N_3076,N_3144);
xor U3937 (N_3937,N_3295,N_3369);
nor U3938 (N_3938,N_3542,N_3294);
nor U3939 (N_3939,N_3312,N_3329);
nand U3940 (N_3940,N_3522,N_3442);
nor U3941 (N_3941,N_3272,N_3545);
xor U3942 (N_3942,N_3567,N_3111);
nor U3943 (N_3943,N_3183,N_3054);
nand U3944 (N_3944,N_3562,N_3414);
or U3945 (N_3945,N_3154,N_3549);
nand U3946 (N_3946,N_3037,N_3010);
nor U3947 (N_3947,N_3388,N_3500);
and U3948 (N_3948,N_3151,N_3019);
and U3949 (N_3949,N_3407,N_3135);
nor U3950 (N_3950,N_3456,N_3062);
nor U3951 (N_3951,N_3548,N_3358);
or U3952 (N_3952,N_3560,N_3470);
nor U3953 (N_3953,N_3416,N_3304);
nor U3954 (N_3954,N_3271,N_3085);
nor U3955 (N_3955,N_3115,N_3308);
xnor U3956 (N_3956,N_3004,N_3210);
or U3957 (N_3957,N_3323,N_3177);
nor U3958 (N_3958,N_3502,N_3077);
or U3959 (N_3959,N_3265,N_3593);
and U3960 (N_3960,N_3336,N_3361);
and U3961 (N_3961,N_3484,N_3326);
nor U3962 (N_3962,N_3140,N_3169);
nor U3963 (N_3963,N_3312,N_3432);
nand U3964 (N_3964,N_3215,N_3015);
or U3965 (N_3965,N_3183,N_3141);
nor U3966 (N_3966,N_3151,N_3005);
xor U3967 (N_3967,N_3048,N_3177);
or U3968 (N_3968,N_3416,N_3032);
and U3969 (N_3969,N_3087,N_3231);
and U3970 (N_3970,N_3028,N_3390);
or U3971 (N_3971,N_3016,N_3501);
nor U3972 (N_3972,N_3561,N_3463);
nand U3973 (N_3973,N_3191,N_3079);
nor U3974 (N_3974,N_3242,N_3209);
and U3975 (N_3975,N_3491,N_3494);
nand U3976 (N_3976,N_3592,N_3301);
nand U3977 (N_3977,N_3433,N_3011);
or U3978 (N_3978,N_3074,N_3139);
nor U3979 (N_3979,N_3413,N_3597);
and U3980 (N_3980,N_3239,N_3364);
xor U3981 (N_3981,N_3403,N_3512);
nor U3982 (N_3982,N_3532,N_3165);
nand U3983 (N_3983,N_3251,N_3314);
nand U3984 (N_3984,N_3026,N_3254);
nor U3985 (N_3985,N_3457,N_3567);
xnor U3986 (N_3986,N_3444,N_3143);
nor U3987 (N_3987,N_3043,N_3087);
and U3988 (N_3988,N_3524,N_3344);
or U3989 (N_3989,N_3100,N_3449);
nor U3990 (N_3990,N_3278,N_3594);
nand U3991 (N_3991,N_3579,N_3519);
or U3992 (N_3992,N_3211,N_3332);
or U3993 (N_3993,N_3492,N_3510);
nor U3994 (N_3994,N_3107,N_3021);
nor U3995 (N_3995,N_3185,N_3164);
xor U3996 (N_3996,N_3099,N_3076);
nand U3997 (N_3997,N_3035,N_3418);
nand U3998 (N_3998,N_3373,N_3173);
xnor U3999 (N_3999,N_3299,N_3335);
and U4000 (N_4000,N_3447,N_3449);
and U4001 (N_4001,N_3016,N_3094);
or U4002 (N_4002,N_3048,N_3578);
and U4003 (N_4003,N_3178,N_3458);
xnor U4004 (N_4004,N_3009,N_3093);
or U4005 (N_4005,N_3530,N_3421);
nor U4006 (N_4006,N_3210,N_3159);
xor U4007 (N_4007,N_3244,N_3013);
and U4008 (N_4008,N_3433,N_3387);
xnor U4009 (N_4009,N_3305,N_3360);
or U4010 (N_4010,N_3333,N_3376);
nand U4011 (N_4011,N_3075,N_3557);
and U4012 (N_4012,N_3111,N_3454);
or U4013 (N_4013,N_3253,N_3440);
xor U4014 (N_4014,N_3050,N_3137);
and U4015 (N_4015,N_3592,N_3090);
or U4016 (N_4016,N_3028,N_3057);
nor U4017 (N_4017,N_3164,N_3388);
and U4018 (N_4018,N_3560,N_3520);
or U4019 (N_4019,N_3261,N_3544);
xnor U4020 (N_4020,N_3508,N_3082);
and U4021 (N_4021,N_3370,N_3410);
nor U4022 (N_4022,N_3131,N_3343);
xor U4023 (N_4023,N_3574,N_3094);
xnor U4024 (N_4024,N_3551,N_3259);
or U4025 (N_4025,N_3511,N_3135);
nand U4026 (N_4026,N_3048,N_3148);
xnor U4027 (N_4027,N_3081,N_3401);
nor U4028 (N_4028,N_3491,N_3498);
and U4029 (N_4029,N_3290,N_3521);
xor U4030 (N_4030,N_3270,N_3557);
xnor U4031 (N_4031,N_3210,N_3056);
nand U4032 (N_4032,N_3083,N_3118);
nand U4033 (N_4033,N_3356,N_3157);
nor U4034 (N_4034,N_3373,N_3567);
or U4035 (N_4035,N_3389,N_3562);
nor U4036 (N_4036,N_3139,N_3564);
xor U4037 (N_4037,N_3444,N_3133);
nand U4038 (N_4038,N_3347,N_3150);
xnor U4039 (N_4039,N_3157,N_3542);
xnor U4040 (N_4040,N_3289,N_3599);
nor U4041 (N_4041,N_3579,N_3046);
nor U4042 (N_4042,N_3465,N_3214);
or U4043 (N_4043,N_3134,N_3269);
and U4044 (N_4044,N_3581,N_3495);
or U4045 (N_4045,N_3384,N_3320);
or U4046 (N_4046,N_3029,N_3012);
xor U4047 (N_4047,N_3158,N_3049);
xor U4048 (N_4048,N_3533,N_3161);
or U4049 (N_4049,N_3071,N_3102);
nand U4050 (N_4050,N_3347,N_3139);
xor U4051 (N_4051,N_3548,N_3271);
nand U4052 (N_4052,N_3196,N_3453);
nor U4053 (N_4053,N_3057,N_3180);
nor U4054 (N_4054,N_3508,N_3403);
xnor U4055 (N_4055,N_3425,N_3161);
or U4056 (N_4056,N_3040,N_3073);
xnor U4057 (N_4057,N_3118,N_3391);
or U4058 (N_4058,N_3568,N_3557);
nand U4059 (N_4059,N_3064,N_3359);
or U4060 (N_4060,N_3360,N_3185);
nor U4061 (N_4061,N_3220,N_3568);
xnor U4062 (N_4062,N_3214,N_3297);
or U4063 (N_4063,N_3349,N_3368);
nor U4064 (N_4064,N_3064,N_3343);
and U4065 (N_4065,N_3408,N_3390);
nand U4066 (N_4066,N_3317,N_3453);
or U4067 (N_4067,N_3143,N_3460);
or U4068 (N_4068,N_3157,N_3004);
nand U4069 (N_4069,N_3261,N_3220);
nor U4070 (N_4070,N_3231,N_3401);
xor U4071 (N_4071,N_3297,N_3581);
xor U4072 (N_4072,N_3098,N_3327);
or U4073 (N_4073,N_3051,N_3184);
xnor U4074 (N_4074,N_3131,N_3566);
nand U4075 (N_4075,N_3426,N_3155);
and U4076 (N_4076,N_3540,N_3091);
or U4077 (N_4077,N_3595,N_3140);
or U4078 (N_4078,N_3305,N_3451);
or U4079 (N_4079,N_3433,N_3194);
nand U4080 (N_4080,N_3015,N_3450);
nor U4081 (N_4081,N_3423,N_3173);
nand U4082 (N_4082,N_3089,N_3261);
or U4083 (N_4083,N_3053,N_3134);
or U4084 (N_4084,N_3442,N_3182);
or U4085 (N_4085,N_3593,N_3080);
nand U4086 (N_4086,N_3105,N_3396);
xnor U4087 (N_4087,N_3381,N_3187);
or U4088 (N_4088,N_3519,N_3235);
nand U4089 (N_4089,N_3326,N_3054);
and U4090 (N_4090,N_3219,N_3511);
or U4091 (N_4091,N_3311,N_3217);
and U4092 (N_4092,N_3278,N_3300);
nor U4093 (N_4093,N_3365,N_3361);
or U4094 (N_4094,N_3178,N_3008);
and U4095 (N_4095,N_3378,N_3367);
xor U4096 (N_4096,N_3559,N_3515);
or U4097 (N_4097,N_3402,N_3466);
and U4098 (N_4098,N_3210,N_3040);
nor U4099 (N_4099,N_3061,N_3489);
nand U4100 (N_4100,N_3263,N_3208);
nand U4101 (N_4101,N_3161,N_3165);
and U4102 (N_4102,N_3135,N_3047);
nand U4103 (N_4103,N_3485,N_3559);
nor U4104 (N_4104,N_3499,N_3218);
nand U4105 (N_4105,N_3271,N_3264);
xor U4106 (N_4106,N_3005,N_3307);
nor U4107 (N_4107,N_3022,N_3587);
or U4108 (N_4108,N_3220,N_3176);
and U4109 (N_4109,N_3467,N_3176);
or U4110 (N_4110,N_3160,N_3068);
or U4111 (N_4111,N_3087,N_3142);
xnor U4112 (N_4112,N_3015,N_3489);
or U4113 (N_4113,N_3078,N_3283);
or U4114 (N_4114,N_3315,N_3287);
and U4115 (N_4115,N_3092,N_3178);
or U4116 (N_4116,N_3009,N_3380);
and U4117 (N_4117,N_3044,N_3107);
nand U4118 (N_4118,N_3483,N_3075);
nor U4119 (N_4119,N_3129,N_3116);
and U4120 (N_4120,N_3302,N_3363);
nand U4121 (N_4121,N_3382,N_3414);
or U4122 (N_4122,N_3250,N_3592);
nand U4123 (N_4123,N_3105,N_3303);
nand U4124 (N_4124,N_3145,N_3210);
nor U4125 (N_4125,N_3264,N_3192);
or U4126 (N_4126,N_3302,N_3420);
nor U4127 (N_4127,N_3567,N_3428);
nor U4128 (N_4128,N_3310,N_3160);
xnor U4129 (N_4129,N_3153,N_3029);
or U4130 (N_4130,N_3374,N_3515);
and U4131 (N_4131,N_3213,N_3167);
or U4132 (N_4132,N_3168,N_3204);
nand U4133 (N_4133,N_3079,N_3158);
nor U4134 (N_4134,N_3420,N_3187);
nand U4135 (N_4135,N_3521,N_3128);
xor U4136 (N_4136,N_3135,N_3448);
nand U4137 (N_4137,N_3465,N_3122);
or U4138 (N_4138,N_3150,N_3245);
xnor U4139 (N_4139,N_3076,N_3559);
xor U4140 (N_4140,N_3581,N_3232);
nor U4141 (N_4141,N_3086,N_3149);
and U4142 (N_4142,N_3122,N_3082);
and U4143 (N_4143,N_3336,N_3267);
xnor U4144 (N_4144,N_3358,N_3496);
nor U4145 (N_4145,N_3288,N_3554);
and U4146 (N_4146,N_3581,N_3267);
xor U4147 (N_4147,N_3019,N_3258);
nand U4148 (N_4148,N_3511,N_3579);
nand U4149 (N_4149,N_3469,N_3275);
nor U4150 (N_4150,N_3449,N_3406);
xor U4151 (N_4151,N_3225,N_3456);
xor U4152 (N_4152,N_3340,N_3431);
and U4153 (N_4153,N_3568,N_3160);
nand U4154 (N_4154,N_3596,N_3459);
xnor U4155 (N_4155,N_3159,N_3062);
nand U4156 (N_4156,N_3471,N_3317);
xor U4157 (N_4157,N_3470,N_3492);
xnor U4158 (N_4158,N_3162,N_3269);
and U4159 (N_4159,N_3290,N_3031);
xor U4160 (N_4160,N_3223,N_3349);
nor U4161 (N_4161,N_3339,N_3080);
nor U4162 (N_4162,N_3233,N_3299);
xor U4163 (N_4163,N_3405,N_3104);
nor U4164 (N_4164,N_3349,N_3213);
nor U4165 (N_4165,N_3564,N_3478);
or U4166 (N_4166,N_3029,N_3460);
or U4167 (N_4167,N_3367,N_3243);
nor U4168 (N_4168,N_3498,N_3392);
or U4169 (N_4169,N_3314,N_3028);
xor U4170 (N_4170,N_3578,N_3432);
or U4171 (N_4171,N_3146,N_3007);
and U4172 (N_4172,N_3170,N_3266);
xor U4173 (N_4173,N_3208,N_3310);
xor U4174 (N_4174,N_3028,N_3459);
nand U4175 (N_4175,N_3336,N_3200);
nand U4176 (N_4176,N_3397,N_3039);
nor U4177 (N_4177,N_3198,N_3510);
and U4178 (N_4178,N_3098,N_3278);
or U4179 (N_4179,N_3357,N_3069);
nand U4180 (N_4180,N_3082,N_3084);
nand U4181 (N_4181,N_3131,N_3110);
and U4182 (N_4182,N_3429,N_3305);
nand U4183 (N_4183,N_3242,N_3504);
or U4184 (N_4184,N_3191,N_3559);
xor U4185 (N_4185,N_3412,N_3434);
and U4186 (N_4186,N_3081,N_3297);
nor U4187 (N_4187,N_3120,N_3099);
or U4188 (N_4188,N_3476,N_3371);
xnor U4189 (N_4189,N_3217,N_3354);
nand U4190 (N_4190,N_3587,N_3394);
xor U4191 (N_4191,N_3056,N_3307);
xnor U4192 (N_4192,N_3070,N_3444);
nand U4193 (N_4193,N_3497,N_3575);
xor U4194 (N_4194,N_3334,N_3161);
or U4195 (N_4195,N_3089,N_3519);
nor U4196 (N_4196,N_3005,N_3271);
and U4197 (N_4197,N_3079,N_3078);
or U4198 (N_4198,N_3239,N_3346);
and U4199 (N_4199,N_3011,N_3009);
xnor U4200 (N_4200,N_4192,N_3770);
or U4201 (N_4201,N_3798,N_3912);
nand U4202 (N_4202,N_4097,N_4063);
nor U4203 (N_4203,N_4127,N_4069);
xor U4204 (N_4204,N_3651,N_4002);
and U4205 (N_4205,N_3750,N_3742);
or U4206 (N_4206,N_4081,N_3849);
xor U4207 (N_4207,N_3623,N_4102);
xor U4208 (N_4208,N_3963,N_3974);
or U4209 (N_4209,N_4100,N_3661);
and U4210 (N_4210,N_4130,N_3642);
xor U4211 (N_4211,N_3757,N_3611);
or U4212 (N_4212,N_3650,N_4095);
xor U4213 (N_4213,N_4070,N_3762);
and U4214 (N_4214,N_4174,N_3712);
nand U4215 (N_4215,N_4111,N_3881);
and U4216 (N_4216,N_3747,N_3619);
and U4217 (N_4217,N_3633,N_3786);
and U4218 (N_4218,N_4010,N_4165);
nor U4219 (N_4219,N_3810,N_3797);
or U4220 (N_4220,N_3721,N_4006);
or U4221 (N_4221,N_3740,N_3732);
and U4222 (N_4222,N_3718,N_3877);
nand U4223 (N_4223,N_3784,N_4123);
nor U4224 (N_4224,N_3741,N_3918);
and U4225 (N_4225,N_3787,N_3905);
nor U4226 (N_4226,N_3645,N_3959);
or U4227 (N_4227,N_3907,N_4046);
or U4228 (N_4228,N_4128,N_3771);
nand U4229 (N_4229,N_4159,N_3823);
or U4230 (N_4230,N_4151,N_3856);
or U4231 (N_4231,N_4021,N_4037);
and U4232 (N_4232,N_3977,N_3956);
nor U4233 (N_4233,N_3711,N_3602);
nor U4234 (N_4234,N_4169,N_4098);
or U4235 (N_4235,N_4049,N_3998);
or U4236 (N_4236,N_3708,N_4008);
and U4237 (N_4237,N_4089,N_3818);
xor U4238 (N_4238,N_4149,N_3719);
xnor U4239 (N_4239,N_3900,N_3863);
nand U4240 (N_4240,N_3846,N_3824);
xnor U4241 (N_4241,N_4059,N_4142);
xnor U4242 (N_4242,N_3945,N_3821);
nand U4243 (N_4243,N_4076,N_4164);
nor U4244 (N_4244,N_4023,N_3731);
or U4245 (N_4245,N_3892,N_3940);
or U4246 (N_4246,N_3816,N_3826);
or U4247 (N_4247,N_3903,N_3815);
xnor U4248 (N_4248,N_3802,N_3928);
nor U4249 (N_4249,N_3803,N_3865);
and U4250 (N_4250,N_3957,N_4012);
nor U4251 (N_4251,N_3922,N_3795);
or U4252 (N_4252,N_4009,N_3831);
or U4253 (N_4253,N_4042,N_3639);
nor U4254 (N_4254,N_4162,N_4168);
nor U4255 (N_4255,N_3871,N_3689);
nor U4256 (N_4256,N_3668,N_3748);
nor U4257 (N_4257,N_4029,N_4099);
and U4258 (N_4258,N_3769,N_3904);
nand U4259 (N_4259,N_3614,N_3669);
nand U4260 (N_4260,N_3999,N_3657);
or U4261 (N_4261,N_4020,N_3788);
or U4262 (N_4262,N_3717,N_3931);
and U4263 (N_4263,N_3613,N_4040);
and U4264 (N_4264,N_3997,N_3898);
nand U4265 (N_4265,N_4190,N_3923);
xor U4266 (N_4266,N_4024,N_3857);
nor U4267 (N_4267,N_3671,N_3832);
and U4268 (N_4268,N_4178,N_4141);
and U4269 (N_4269,N_3807,N_3801);
or U4270 (N_4270,N_3701,N_3683);
nand U4271 (N_4271,N_3709,N_3843);
xnor U4272 (N_4272,N_3682,N_4167);
and U4273 (N_4273,N_3860,N_4093);
nor U4274 (N_4274,N_3775,N_3728);
xnor U4275 (N_4275,N_3972,N_3906);
nand U4276 (N_4276,N_4031,N_4054);
nand U4277 (N_4277,N_4073,N_3858);
or U4278 (N_4278,N_3799,N_3993);
nand U4279 (N_4279,N_3791,N_3636);
nor U4280 (N_4280,N_3938,N_4157);
nand U4281 (N_4281,N_4147,N_4041);
nor U4282 (N_4282,N_3745,N_3899);
nor U4283 (N_4283,N_3790,N_3943);
nor U4284 (N_4284,N_3941,N_3896);
xor U4285 (N_4285,N_4148,N_3984);
or U4286 (N_4286,N_3975,N_4087);
xnor U4287 (N_4287,N_3612,N_3820);
nand U4288 (N_4288,N_3631,N_3991);
nand U4289 (N_4289,N_4060,N_3654);
xor U4290 (N_4290,N_3618,N_3814);
nand U4291 (N_4291,N_4000,N_3765);
and U4292 (N_4292,N_3674,N_3944);
nor U4293 (N_4293,N_4194,N_3796);
nor U4294 (N_4294,N_3994,N_4119);
nor U4295 (N_4295,N_3764,N_4110);
nand U4296 (N_4296,N_3932,N_3793);
or U4297 (N_4297,N_4121,N_3847);
and U4298 (N_4298,N_4027,N_3686);
nand U4299 (N_4299,N_3607,N_3872);
xor U4300 (N_4300,N_4072,N_3656);
or U4301 (N_4301,N_3838,N_3722);
xnor U4302 (N_4302,N_4005,N_3679);
nor U4303 (N_4303,N_3664,N_3973);
or U4304 (N_4304,N_3780,N_3610);
or U4305 (N_4305,N_3926,N_4105);
or U4306 (N_4306,N_3879,N_4101);
and U4307 (N_4307,N_3919,N_4039);
nand U4308 (N_4308,N_4077,N_4177);
or U4309 (N_4309,N_3707,N_3996);
and U4310 (N_4310,N_3658,N_4187);
or U4311 (N_4311,N_3672,N_3734);
or U4312 (N_4312,N_4064,N_4195);
or U4313 (N_4313,N_3710,N_4183);
xor U4314 (N_4314,N_4026,N_4172);
nor U4315 (N_4315,N_3884,N_3894);
or U4316 (N_4316,N_3813,N_3874);
xor U4317 (N_4317,N_4090,N_3681);
nor U4318 (N_4318,N_4103,N_3729);
or U4319 (N_4319,N_4083,N_3714);
xor U4320 (N_4320,N_3976,N_3883);
or U4321 (N_4321,N_4156,N_3962);
nor U4322 (N_4322,N_3634,N_3933);
xnor U4323 (N_4323,N_4084,N_3696);
nand U4324 (N_4324,N_3949,N_4061);
and U4325 (N_4325,N_3692,N_3632);
and U4326 (N_4326,N_3864,N_3951);
nand U4327 (N_4327,N_3715,N_3897);
xnor U4328 (N_4328,N_3659,N_3617);
or U4329 (N_4329,N_3827,N_3893);
xnor U4330 (N_4330,N_4135,N_3836);
nand U4331 (N_4331,N_3990,N_4025);
xnor U4332 (N_4332,N_3646,N_3759);
xor U4333 (N_4333,N_4197,N_3806);
nor U4334 (N_4334,N_3822,N_4139);
xnor U4335 (N_4335,N_3667,N_3861);
nor U4336 (N_4336,N_4136,N_4001);
xnor U4337 (N_4337,N_3809,N_3862);
and U4338 (N_4338,N_3624,N_3675);
nor U4339 (N_4339,N_3605,N_4011);
and U4340 (N_4340,N_3615,N_3804);
xor U4341 (N_4341,N_3635,N_3687);
and U4342 (N_4342,N_3867,N_4088);
nand U4343 (N_4343,N_4131,N_4045);
or U4344 (N_4344,N_4092,N_4066);
xnor U4345 (N_4345,N_3890,N_3819);
or U4346 (N_4346,N_3678,N_3660);
or U4347 (N_4347,N_3965,N_3727);
and U4348 (N_4348,N_3979,N_4004);
or U4349 (N_4349,N_3968,N_3915);
nor U4350 (N_4350,N_4052,N_3980);
or U4351 (N_4351,N_3684,N_3758);
and U4352 (N_4352,N_3697,N_3653);
and U4353 (N_4353,N_4138,N_3604);
or U4354 (N_4354,N_3924,N_3781);
and U4355 (N_4355,N_3737,N_4118);
nand U4356 (N_4356,N_3774,N_4079);
nor U4357 (N_4357,N_4150,N_3950);
or U4358 (N_4358,N_3842,N_3772);
and U4359 (N_4359,N_3992,N_3647);
and U4360 (N_4360,N_3695,N_3670);
or U4361 (N_4361,N_4146,N_3783);
nand U4362 (N_4362,N_4182,N_3828);
nor U4363 (N_4363,N_3730,N_4199);
nand U4364 (N_4364,N_4188,N_3855);
or U4365 (N_4365,N_3920,N_4155);
nor U4366 (N_4366,N_4067,N_4114);
nand U4367 (N_4367,N_3886,N_4158);
nand U4368 (N_4368,N_3985,N_4122);
nand U4369 (N_4369,N_3725,N_4152);
and U4370 (N_4370,N_3735,N_4137);
or U4371 (N_4371,N_3913,N_4003);
and U4372 (N_4372,N_4030,N_3776);
and U4373 (N_4373,N_4016,N_3811);
and U4374 (N_4374,N_4189,N_3960);
and U4375 (N_4375,N_3794,N_3887);
xnor U4376 (N_4376,N_3700,N_3603);
or U4377 (N_4377,N_4019,N_3652);
xor U4378 (N_4378,N_3724,N_4104);
nand U4379 (N_4379,N_3850,N_4056);
nand U4380 (N_4380,N_3812,N_4120);
and U4381 (N_4381,N_3702,N_3703);
nand U4382 (N_4382,N_3763,N_3627);
nand U4383 (N_4383,N_3889,N_3981);
nor U4384 (N_4384,N_4198,N_3964);
xnor U4385 (N_4385,N_4062,N_3989);
or U4386 (N_4386,N_4048,N_3649);
or U4387 (N_4387,N_3914,N_3917);
nand U4388 (N_4388,N_3738,N_4065);
xor U4389 (N_4389,N_3937,N_4171);
nand U4390 (N_4390,N_3640,N_4175);
nor U4391 (N_4391,N_4106,N_3644);
nand U4392 (N_4392,N_3978,N_3666);
and U4393 (N_4393,N_3676,N_3609);
nor U4394 (N_4394,N_4126,N_4028);
and U4395 (N_4395,N_3726,N_3921);
nand U4396 (N_4396,N_3885,N_3746);
nor U4397 (N_4397,N_4166,N_3854);
or U4398 (N_4398,N_3739,N_3983);
or U4399 (N_4399,N_4068,N_3637);
and U4400 (N_4400,N_3625,N_3608);
or U4401 (N_4401,N_3995,N_3853);
and U4402 (N_4402,N_3648,N_4038);
and U4403 (N_4403,N_4108,N_3680);
nor U4404 (N_4404,N_4047,N_3955);
nand U4405 (N_4405,N_4057,N_3888);
and U4406 (N_4406,N_4112,N_3840);
xnor U4407 (N_4407,N_4109,N_3800);
and U4408 (N_4408,N_3839,N_3939);
nor U4409 (N_4409,N_3848,N_3751);
and U4410 (N_4410,N_3835,N_3982);
or U4411 (N_4411,N_4132,N_3690);
and U4412 (N_4412,N_3643,N_4154);
and U4413 (N_4413,N_3691,N_4191);
and U4414 (N_4414,N_3936,N_4078);
or U4415 (N_4415,N_3971,N_4161);
and U4416 (N_4416,N_3902,N_3778);
and U4417 (N_4417,N_3952,N_3916);
or U4418 (N_4418,N_3930,N_3673);
or U4419 (N_4419,N_3880,N_3789);
or U4420 (N_4420,N_3833,N_3895);
nor U4421 (N_4421,N_3622,N_3935);
and U4422 (N_4422,N_3626,N_3875);
or U4423 (N_4423,N_4032,N_3829);
nand U4424 (N_4424,N_4170,N_3629);
nor U4425 (N_4425,N_4186,N_3754);
nand U4426 (N_4426,N_3954,N_4050);
nand U4427 (N_4427,N_4051,N_3948);
xor U4428 (N_4428,N_3841,N_3852);
nand U4429 (N_4429,N_3706,N_3878);
xnor U4430 (N_4430,N_3616,N_4145);
or U4431 (N_4431,N_3630,N_4033);
nand U4432 (N_4432,N_4080,N_3699);
or U4433 (N_4433,N_3688,N_4144);
xnor U4434 (N_4434,N_4185,N_3792);
nor U4435 (N_4435,N_4053,N_4176);
or U4436 (N_4436,N_3986,N_3723);
or U4437 (N_4437,N_4115,N_3870);
or U4438 (N_4438,N_3663,N_3934);
nand U4439 (N_4439,N_4140,N_3621);
xnor U4440 (N_4440,N_3693,N_3744);
nor U4441 (N_4441,N_4036,N_3805);
nand U4442 (N_4442,N_3743,N_4129);
nor U4443 (N_4443,N_3641,N_3677);
or U4444 (N_4444,N_3779,N_3851);
xor U4445 (N_4445,N_4116,N_3736);
xor U4446 (N_4446,N_3910,N_4117);
nand U4447 (N_4447,N_3837,N_3698);
and U4448 (N_4448,N_4134,N_3876);
or U4449 (N_4449,N_3755,N_3908);
or U4450 (N_4450,N_3966,N_4071);
or U4451 (N_4451,N_3777,N_3901);
and U4452 (N_4452,N_4153,N_3942);
and U4453 (N_4453,N_3752,N_4018);
xor U4454 (N_4454,N_3859,N_3825);
nor U4455 (N_4455,N_4055,N_3768);
nor U4456 (N_4456,N_3665,N_3704);
xor U4457 (N_4457,N_4082,N_3873);
xnor U4458 (N_4458,N_3705,N_4035);
nand U4459 (N_4459,N_4007,N_3946);
or U4460 (N_4460,N_4133,N_3909);
nor U4461 (N_4461,N_4086,N_3845);
nor U4462 (N_4462,N_3601,N_4034);
or U4463 (N_4463,N_4058,N_3749);
nand U4464 (N_4464,N_4075,N_3600);
or U4465 (N_4465,N_3628,N_4181);
or U4466 (N_4466,N_4094,N_4091);
nor U4467 (N_4467,N_3756,N_4143);
xnor U4468 (N_4468,N_3760,N_3685);
or U4469 (N_4469,N_4193,N_3988);
nor U4470 (N_4470,N_3961,N_3716);
xnor U4471 (N_4471,N_3970,N_3868);
and U4472 (N_4472,N_4173,N_3844);
and U4473 (N_4473,N_3638,N_4013);
xor U4474 (N_4474,N_3620,N_3817);
nor U4475 (N_4475,N_4085,N_3655);
xor U4476 (N_4476,N_3891,N_3830);
or U4477 (N_4477,N_4044,N_4125);
or U4478 (N_4478,N_3958,N_4196);
nand U4479 (N_4479,N_4124,N_4179);
xor U4480 (N_4480,N_3987,N_3866);
and U4481 (N_4481,N_4096,N_3766);
nand U4482 (N_4482,N_3927,N_3929);
nand U4483 (N_4483,N_3782,N_4184);
or U4484 (N_4484,N_4107,N_3969);
xnor U4485 (N_4485,N_4113,N_4074);
or U4486 (N_4486,N_3785,N_3967);
or U4487 (N_4487,N_3911,N_3753);
and U4488 (N_4488,N_3947,N_3720);
or U4489 (N_4489,N_3662,N_4043);
xor U4490 (N_4490,N_3694,N_3773);
and U4491 (N_4491,N_3767,N_4014);
and U4492 (N_4492,N_4022,N_4015);
and U4493 (N_4493,N_3869,N_3606);
or U4494 (N_4494,N_4160,N_4017);
and U4495 (N_4495,N_3713,N_3761);
or U4496 (N_4496,N_3925,N_4163);
and U4497 (N_4497,N_3834,N_3882);
xnor U4498 (N_4498,N_3953,N_3733);
xnor U4499 (N_4499,N_3808,N_4180);
nor U4500 (N_4500,N_3969,N_3696);
xnor U4501 (N_4501,N_3607,N_3809);
or U4502 (N_4502,N_4030,N_3723);
nand U4503 (N_4503,N_3666,N_3649);
or U4504 (N_4504,N_3919,N_3861);
xor U4505 (N_4505,N_3756,N_3721);
or U4506 (N_4506,N_3778,N_4021);
nand U4507 (N_4507,N_3902,N_3692);
xnor U4508 (N_4508,N_3865,N_3992);
nand U4509 (N_4509,N_3971,N_3822);
nand U4510 (N_4510,N_3869,N_3617);
or U4511 (N_4511,N_4130,N_3974);
nor U4512 (N_4512,N_4191,N_3775);
and U4513 (N_4513,N_4113,N_3811);
and U4514 (N_4514,N_3944,N_3763);
nor U4515 (N_4515,N_3933,N_3953);
nand U4516 (N_4516,N_4158,N_4007);
or U4517 (N_4517,N_3605,N_3774);
or U4518 (N_4518,N_3822,N_3631);
and U4519 (N_4519,N_3901,N_3603);
or U4520 (N_4520,N_3616,N_3839);
or U4521 (N_4521,N_3781,N_3706);
and U4522 (N_4522,N_3631,N_3982);
nand U4523 (N_4523,N_3812,N_3821);
and U4524 (N_4524,N_4126,N_4083);
and U4525 (N_4525,N_3850,N_4096);
xnor U4526 (N_4526,N_3641,N_3979);
or U4527 (N_4527,N_3913,N_3601);
nand U4528 (N_4528,N_3884,N_3661);
xor U4529 (N_4529,N_4093,N_3904);
xnor U4530 (N_4530,N_3794,N_4034);
nand U4531 (N_4531,N_3757,N_4185);
or U4532 (N_4532,N_3781,N_3768);
nand U4533 (N_4533,N_3742,N_4037);
and U4534 (N_4534,N_3966,N_4157);
or U4535 (N_4535,N_3649,N_3868);
or U4536 (N_4536,N_3990,N_3718);
or U4537 (N_4537,N_3756,N_3663);
or U4538 (N_4538,N_4177,N_4199);
nand U4539 (N_4539,N_4030,N_4058);
nand U4540 (N_4540,N_3838,N_4130);
or U4541 (N_4541,N_3859,N_3804);
xor U4542 (N_4542,N_3691,N_4067);
nor U4543 (N_4543,N_4105,N_3839);
or U4544 (N_4544,N_3847,N_3658);
and U4545 (N_4545,N_3692,N_3608);
or U4546 (N_4546,N_4058,N_3797);
nor U4547 (N_4547,N_3710,N_3902);
nor U4548 (N_4548,N_3966,N_4171);
nor U4549 (N_4549,N_3689,N_4090);
nand U4550 (N_4550,N_4127,N_4077);
and U4551 (N_4551,N_3925,N_3936);
or U4552 (N_4552,N_4149,N_4185);
nand U4553 (N_4553,N_3806,N_4050);
and U4554 (N_4554,N_4196,N_4173);
xor U4555 (N_4555,N_3638,N_3643);
and U4556 (N_4556,N_3787,N_3892);
nor U4557 (N_4557,N_3827,N_4099);
nand U4558 (N_4558,N_3920,N_3884);
nor U4559 (N_4559,N_4079,N_4129);
or U4560 (N_4560,N_4154,N_4041);
nor U4561 (N_4561,N_3810,N_4013);
and U4562 (N_4562,N_3782,N_3605);
xnor U4563 (N_4563,N_4074,N_3642);
nand U4564 (N_4564,N_3827,N_3984);
and U4565 (N_4565,N_3966,N_3941);
nor U4566 (N_4566,N_3716,N_3655);
xnor U4567 (N_4567,N_3901,N_3708);
or U4568 (N_4568,N_4137,N_4196);
or U4569 (N_4569,N_3925,N_3749);
nand U4570 (N_4570,N_3759,N_4042);
nand U4571 (N_4571,N_3638,N_3905);
or U4572 (N_4572,N_3684,N_4118);
or U4573 (N_4573,N_3640,N_4042);
nand U4574 (N_4574,N_3866,N_3898);
xnor U4575 (N_4575,N_3891,N_4029);
xor U4576 (N_4576,N_3965,N_3784);
xor U4577 (N_4577,N_3884,N_4086);
and U4578 (N_4578,N_3647,N_3646);
xor U4579 (N_4579,N_3715,N_3710);
nor U4580 (N_4580,N_4131,N_3822);
nand U4581 (N_4581,N_3734,N_4114);
xnor U4582 (N_4582,N_3654,N_4091);
nor U4583 (N_4583,N_3911,N_4117);
or U4584 (N_4584,N_4069,N_3655);
xor U4585 (N_4585,N_4176,N_4143);
and U4586 (N_4586,N_3743,N_4080);
nor U4587 (N_4587,N_3866,N_3735);
or U4588 (N_4588,N_3780,N_3776);
xnor U4589 (N_4589,N_3631,N_4067);
and U4590 (N_4590,N_3788,N_3979);
nand U4591 (N_4591,N_3976,N_4057);
nand U4592 (N_4592,N_4060,N_3854);
and U4593 (N_4593,N_3816,N_3954);
and U4594 (N_4594,N_4083,N_4009);
xnor U4595 (N_4595,N_3934,N_3606);
and U4596 (N_4596,N_4048,N_3617);
nand U4597 (N_4597,N_4083,N_3844);
and U4598 (N_4598,N_3940,N_4130);
nand U4599 (N_4599,N_3923,N_3773);
nand U4600 (N_4600,N_3797,N_3686);
or U4601 (N_4601,N_4152,N_3978);
and U4602 (N_4602,N_4118,N_3946);
or U4603 (N_4603,N_4166,N_3732);
nor U4604 (N_4604,N_3818,N_3690);
xor U4605 (N_4605,N_3990,N_3647);
nor U4606 (N_4606,N_4194,N_3702);
and U4607 (N_4607,N_3804,N_3851);
nor U4608 (N_4608,N_4186,N_4069);
nor U4609 (N_4609,N_3746,N_4155);
nor U4610 (N_4610,N_3890,N_3610);
or U4611 (N_4611,N_4084,N_4075);
nand U4612 (N_4612,N_4111,N_4049);
nand U4613 (N_4613,N_4081,N_3629);
xnor U4614 (N_4614,N_3739,N_3810);
nand U4615 (N_4615,N_4100,N_4171);
nor U4616 (N_4616,N_3693,N_4172);
xnor U4617 (N_4617,N_3752,N_3715);
and U4618 (N_4618,N_3776,N_3787);
xnor U4619 (N_4619,N_4002,N_3928);
and U4620 (N_4620,N_4198,N_3761);
and U4621 (N_4621,N_3648,N_4035);
nor U4622 (N_4622,N_4121,N_4157);
and U4623 (N_4623,N_3708,N_3911);
or U4624 (N_4624,N_3882,N_4197);
or U4625 (N_4625,N_3678,N_3694);
nor U4626 (N_4626,N_3651,N_3908);
or U4627 (N_4627,N_3672,N_4094);
nor U4628 (N_4628,N_3615,N_4089);
and U4629 (N_4629,N_3833,N_3753);
and U4630 (N_4630,N_4086,N_3867);
nor U4631 (N_4631,N_4086,N_3643);
nor U4632 (N_4632,N_4116,N_3933);
xnor U4633 (N_4633,N_3861,N_3713);
or U4634 (N_4634,N_4013,N_3794);
nand U4635 (N_4635,N_3732,N_4003);
and U4636 (N_4636,N_3856,N_3915);
and U4637 (N_4637,N_4092,N_4183);
or U4638 (N_4638,N_3732,N_3639);
and U4639 (N_4639,N_3713,N_3921);
nor U4640 (N_4640,N_4004,N_3746);
nand U4641 (N_4641,N_4158,N_3728);
or U4642 (N_4642,N_3776,N_3676);
or U4643 (N_4643,N_3753,N_4108);
and U4644 (N_4644,N_4025,N_4115);
and U4645 (N_4645,N_4124,N_3978);
or U4646 (N_4646,N_3880,N_4066);
and U4647 (N_4647,N_3955,N_3841);
nand U4648 (N_4648,N_4072,N_4138);
xnor U4649 (N_4649,N_4110,N_4153);
nand U4650 (N_4650,N_3736,N_3710);
xor U4651 (N_4651,N_4155,N_3864);
and U4652 (N_4652,N_3825,N_3687);
xor U4653 (N_4653,N_3889,N_4194);
nor U4654 (N_4654,N_3668,N_3666);
or U4655 (N_4655,N_3676,N_4134);
nor U4656 (N_4656,N_3731,N_4152);
or U4657 (N_4657,N_3900,N_3781);
or U4658 (N_4658,N_3626,N_3635);
and U4659 (N_4659,N_3844,N_3843);
nand U4660 (N_4660,N_3985,N_3716);
nand U4661 (N_4661,N_3806,N_3894);
and U4662 (N_4662,N_4094,N_3843);
or U4663 (N_4663,N_3824,N_3735);
nor U4664 (N_4664,N_3997,N_4185);
and U4665 (N_4665,N_3651,N_3823);
nand U4666 (N_4666,N_3970,N_3932);
nand U4667 (N_4667,N_3857,N_4033);
nand U4668 (N_4668,N_4191,N_4181);
and U4669 (N_4669,N_3822,N_4040);
nor U4670 (N_4670,N_3879,N_4157);
or U4671 (N_4671,N_4107,N_3876);
and U4672 (N_4672,N_3882,N_4093);
xor U4673 (N_4673,N_3653,N_4032);
or U4674 (N_4674,N_3692,N_3909);
and U4675 (N_4675,N_4069,N_3779);
xnor U4676 (N_4676,N_3980,N_3601);
and U4677 (N_4677,N_3701,N_3611);
and U4678 (N_4678,N_4071,N_3942);
and U4679 (N_4679,N_4143,N_3808);
nor U4680 (N_4680,N_4070,N_3909);
or U4681 (N_4681,N_3945,N_3908);
nor U4682 (N_4682,N_4145,N_3926);
nand U4683 (N_4683,N_4133,N_4008);
and U4684 (N_4684,N_3980,N_3855);
and U4685 (N_4685,N_4139,N_4084);
and U4686 (N_4686,N_3631,N_3829);
xnor U4687 (N_4687,N_4193,N_3844);
and U4688 (N_4688,N_3876,N_3893);
nand U4689 (N_4689,N_3961,N_4030);
and U4690 (N_4690,N_3736,N_3922);
and U4691 (N_4691,N_3662,N_3823);
or U4692 (N_4692,N_4167,N_4195);
nor U4693 (N_4693,N_4120,N_4109);
nor U4694 (N_4694,N_3993,N_4160);
and U4695 (N_4695,N_4164,N_3603);
or U4696 (N_4696,N_3969,N_4145);
nand U4697 (N_4697,N_4120,N_3956);
xnor U4698 (N_4698,N_3764,N_4059);
nand U4699 (N_4699,N_4106,N_4105);
and U4700 (N_4700,N_3820,N_3856);
or U4701 (N_4701,N_3643,N_4192);
and U4702 (N_4702,N_4014,N_4075);
and U4703 (N_4703,N_3701,N_4062);
or U4704 (N_4704,N_3685,N_3967);
or U4705 (N_4705,N_4160,N_3755);
and U4706 (N_4706,N_3872,N_4083);
nor U4707 (N_4707,N_3802,N_4006);
nor U4708 (N_4708,N_4176,N_3646);
or U4709 (N_4709,N_3979,N_3947);
nand U4710 (N_4710,N_4193,N_3643);
xor U4711 (N_4711,N_3930,N_3946);
nor U4712 (N_4712,N_3614,N_4150);
nor U4713 (N_4713,N_3703,N_3995);
or U4714 (N_4714,N_3810,N_4007);
nor U4715 (N_4715,N_3736,N_3928);
nand U4716 (N_4716,N_4122,N_4060);
nand U4717 (N_4717,N_3794,N_3918);
nand U4718 (N_4718,N_4068,N_3896);
xnor U4719 (N_4719,N_3670,N_4117);
nand U4720 (N_4720,N_4030,N_3710);
xnor U4721 (N_4721,N_3601,N_3685);
nand U4722 (N_4722,N_3703,N_3828);
nor U4723 (N_4723,N_3776,N_4144);
or U4724 (N_4724,N_4182,N_3740);
nand U4725 (N_4725,N_3678,N_4015);
and U4726 (N_4726,N_3640,N_4054);
xor U4727 (N_4727,N_3817,N_3637);
xnor U4728 (N_4728,N_4124,N_3746);
xnor U4729 (N_4729,N_3650,N_4170);
nand U4730 (N_4730,N_3660,N_4146);
xnor U4731 (N_4731,N_3887,N_3608);
and U4732 (N_4732,N_4148,N_3833);
xnor U4733 (N_4733,N_3990,N_3711);
nor U4734 (N_4734,N_4144,N_4037);
or U4735 (N_4735,N_3879,N_3622);
and U4736 (N_4736,N_3834,N_3935);
nor U4737 (N_4737,N_3641,N_3815);
xnor U4738 (N_4738,N_3864,N_3874);
nor U4739 (N_4739,N_3738,N_3877);
or U4740 (N_4740,N_3866,N_4104);
or U4741 (N_4741,N_3755,N_3891);
or U4742 (N_4742,N_4197,N_3600);
nor U4743 (N_4743,N_3631,N_3712);
nor U4744 (N_4744,N_3683,N_3834);
or U4745 (N_4745,N_4131,N_3966);
nor U4746 (N_4746,N_4033,N_3666);
nand U4747 (N_4747,N_4105,N_4167);
xnor U4748 (N_4748,N_4034,N_3822);
and U4749 (N_4749,N_3646,N_3693);
nor U4750 (N_4750,N_3774,N_3753);
xnor U4751 (N_4751,N_3858,N_4003);
xor U4752 (N_4752,N_3806,N_3829);
and U4753 (N_4753,N_3959,N_3699);
xor U4754 (N_4754,N_3632,N_3691);
nor U4755 (N_4755,N_4169,N_3706);
nand U4756 (N_4756,N_3722,N_3792);
or U4757 (N_4757,N_3785,N_4060);
nand U4758 (N_4758,N_3801,N_3697);
xor U4759 (N_4759,N_4164,N_3966);
nor U4760 (N_4760,N_3757,N_4111);
nor U4761 (N_4761,N_4183,N_4020);
xor U4762 (N_4762,N_3983,N_4106);
nand U4763 (N_4763,N_4102,N_3728);
or U4764 (N_4764,N_3857,N_3720);
or U4765 (N_4765,N_4145,N_3728);
or U4766 (N_4766,N_4066,N_3835);
nand U4767 (N_4767,N_4065,N_3940);
nor U4768 (N_4768,N_3604,N_4169);
xor U4769 (N_4769,N_3658,N_3775);
nor U4770 (N_4770,N_3770,N_4083);
nand U4771 (N_4771,N_3737,N_3781);
and U4772 (N_4772,N_3626,N_3912);
and U4773 (N_4773,N_3971,N_3751);
nor U4774 (N_4774,N_3799,N_3726);
or U4775 (N_4775,N_3700,N_4124);
and U4776 (N_4776,N_4080,N_3679);
and U4777 (N_4777,N_3632,N_3636);
xor U4778 (N_4778,N_3801,N_3854);
and U4779 (N_4779,N_3743,N_3957);
nand U4780 (N_4780,N_4092,N_4132);
and U4781 (N_4781,N_3946,N_4088);
xor U4782 (N_4782,N_4194,N_4071);
xnor U4783 (N_4783,N_3645,N_4049);
nor U4784 (N_4784,N_4069,N_3650);
nor U4785 (N_4785,N_3647,N_3982);
or U4786 (N_4786,N_4106,N_4107);
or U4787 (N_4787,N_4063,N_4086);
and U4788 (N_4788,N_4102,N_3686);
nand U4789 (N_4789,N_3660,N_4193);
nand U4790 (N_4790,N_4093,N_4091);
xnor U4791 (N_4791,N_4070,N_4050);
or U4792 (N_4792,N_4176,N_3728);
xnor U4793 (N_4793,N_4169,N_3986);
xnor U4794 (N_4794,N_3826,N_4068);
nor U4795 (N_4795,N_3707,N_3758);
or U4796 (N_4796,N_3763,N_3606);
xor U4797 (N_4797,N_4002,N_3757);
nor U4798 (N_4798,N_3769,N_4116);
nor U4799 (N_4799,N_4073,N_3965);
and U4800 (N_4800,N_4788,N_4585);
or U4801 (N_4801,N_4286,N_4666);
and U4802 (N_4802,N_4789,N_4553);
or U4803 (N_4803,N_4589,N_4477);
and U4804 (N_4804,N_4658,N_4257);
xnor U4805 (N_4805,N_4695,N_4757);
or U4806 (N_4806,N_4224,N_4519);
nor U4807 (N_4807,N_4292,N_4772);
nand U4808 (N_4808,N_4603,N_4685);
nand U4809 (N_4809,N_4366,N_4750);
and U4810 (N_4810,N_4451,N_4416);
xnor U4811 (N_4811,N_4299,N_4435);
nand U4812 (N_4812,N_4475,N_4221);
or U4813 (N_4813,N_4582,N_4333);
or U4814 (N_4814,N_4775,N_4216);
and U4815 (N_4815,N_4497,N_4574);
nand U4816 (N_4816,N_4243,N_4262);
nor U4817 (N_4817,N_4365,N_4456);
nand U4818 (N_4818,N_4326,N_4638);
or U4819 (N_4819,N_4552,N_4606);
or U4820 (N_4820,N_4222,N_4373);
nor U4821 (N_4821,N_4533,N_4662);
nand U4822 (N_4822,N_4282,N_4646);
nor U4823 (N_4823,N_4278,N_4315);
xor U4824 (N_4824,N_4454,N_4537);
or U4825 (N_4825,N_4626,N_4424);
xnor U4826 (N_4826,N_4488,N_4781);
or U4827 (N_4827,N_4432,N_4518);
nand U4828 (N_4828,N_4705,N_4710);
or U4829 (N_4829,N_4521,N_4590);
nor U4830 (N_4830,N_4235,N_4226);
xor U4831 (N_4831,N_4461,N_4274);
or U4832 (N_4832,N_4479,N_4682);
and U4833 (N_4833,N_4740,N_4650);
xor U4834 (N_4834,N_4391,N_4717);
or U4835 (N_4835,N_4276,N_4527);
xor U4836 (N_4836,N_4669,N_4546);
and U4837 (N_4837,N_4382,N_4607);
and U4838 (N_4838,N_4377,N_4609);
and U4839 (N_4839,N_4792,N_4237);
or U4840 (N_4840,N_4207,N_4594);
nand U4841 (N_4841,N_4616,N_4399);
nor U4842 (N_4842,N_4450,N_4718);
xor U4843 (N_4843,N_4752,N_4200);
xnor U4844 (N_4844,N_4770,N_4637);
nor U4845 (N_4845,N_4393,N_4783);
xnor U4846 (N_4846,N_4564,N_4690);
nand U4847 (N_4847,N_4334,N_4671);
or U4848 (N_4848,N_4211,N_4431);
or U4849 (N_4849,N_4766,N_4360);
nor U4850 (N_4850,N_4608,N_4634);
nor U4851 (N_4851,N_4556,N_4245);
xor U4852 (N_4852,N_4641,N_4762);
nor U4853 (N_4853,N_4507,N_4723);
nor U4854 (N_4854,N_4768,N_4532);
or U4855 (N_4855,N_4268,N_4485);
and U4856 (N_4856,N_4653,N_4390);
and U4857 (N_4857,N_4678,N_4396);
nor U4858 (N_4858,N_4329,N_4541);
nand U4859 (N_4859,N_4376,N_4426);
xnor U4860 (N_4860,N_4528,N_4271);
and U4861 (N_4861,N_4332,N_4595);
xor U4862 (N_4862,N_4331,N_4526);
or U4863 (N_4863,N_4795,N_4489);
and U4864 (N_4864,N_4625,N_4511);
nor U4865 (N_4865,N_4765,N_4478);
nor U4866 (N_4866,N_4417,N_4720);
and U4867 (N_4867,N_4255,N_4675);
xnor U4868 (N_4868,N_4277,N_4597);
and U4869 (N_4869,N_4463,N_4645);
and U4870 (N_4870,N_4706,N_4505);
or U4871 (N_4871,N_4520,N_4325);
xor U4872 (N_4872,N_4305,N_4580);
nand U4873 (N_4873,N_4627,N_4324);
nand U4874 (N_4874,N_4313,N_4438);
nor U4875 (N_4875,N_4730,N_4676);
and U4876 (N_4876,N_4384,N_4364);
xnor U4877 (N_4877,N_4615,N_4764);
or U4878 (N_4878,N_4667,N_4492);
or U4879 (N_4879,N_4576,N_4794);
and U4880 (N_4880,N_4735,N_4458);
or U4881 (N_4881,N_4452,N_4363);
nor U4882 (N_4882,N_4756,N_4240);
and U4883 (N_4883,N_4287,N_4400);
xnor U4884 (N_4884,N_4696,N_4686);
and U4885 (N_4885,N_4445,N_4515);
xnor U4886 (N_4886,N_4535,N_4529);
xor U4887 (N_4887,N_4408,N_4231);
nor U4888 (N_4888,N_4621,N_4579);
and U4889 (N_4889,N_4578,N_4655);
and U4890 (N_4890,N_4563,N_4714);
or U4891 (N_4891,N_4449,N_4623);
nor U4892 (N_4892,N_4525,N_4264);
nand U4893 (N_4893,N_4244,N_4584);
nor U4894 (N_4894,N_4354,N_4620);
nor U4895 (N_4895,N_4760,N_4322);
or U4896 (N_4896,N_4692,N_4350);
xnor U4897 (N_4897,N_4447,N_4374);
nor U4898 (N_4898,N_4241,N_4504);
nand U4899 (N_4899,N_4266,N_4203);
nand U4900 (N_4900,N_4425,N_4739);
nor U4901 (N_4901,N_4462,N_4403);
or U4902 (N_4902,N_4743,N_4443);
or U4903 (N_4903,N_4596,N_4261);
or U4904 (N_4904,N_4547,N_4630);
and U4905 (N_4905,N_4604,N_4440);
and U4906 (N_4906,N_4567,N_4272);
or U4907 (N_4907,N_4367,N_4279);
and U4908 (N_4908,N_4651,N_4633);
nand U4909 (N_4909,N_4742,N_4407);
nand U4910 (N_4910,N_4737,N_4549);
nor U4911 (N_4911,N_4383,N_4728);
nand U4912 (N_4912,N_4668,N_4771);
nor U4913 (N_4913,N_4665,N_4618);
nand U4914 (N_4914,N_4388,N_4265);
xnor U4915 (N_4915,N_4712,N_4540);
nor U4916 (N_4916,N_4412,N_4751);
or U4917 (N_4917,N_4748,N_4711);
xnor U4918 (N_4918,N_4500,N_4729);
nor U4919 (N_4919,N_4288,N_4738);
or U4920 (N_4920,N_4782,N_4531);
nor U4921 (N_4921,N_4514,N_4444);
nand U4922 (N_4922,N_4734,N_4337);
nand U4923 (N_4923,N_4746,N_4275);
xor U4924 (N_4924,N_4709,N_4797);
and U4925 (N_4925,N_4430,N_4679);
nor U4926 (N_4926,N_4465,N_4508);
and U4927 (N_4927,N_4311,N_4640);
or U4928 (N_4928,N_4306,N_4428);
xnor U4929 (N_4929,N_4759,N_4591);
and U4930 (N_4930,N_4427,N_4600);
nand U4931 (N_4931,N_4569,N_4283);
nor U4932 (N_4932,N_4524,N_4660);
xnor U4933 (N_4933,N_4523,N_4688);
nand U4934 (N_4934,N_4559,N_4309);
or U4935 (N_4935,N_4338,N_4494);
nor U4936 (N_4936,N_4753,N_4544);
nor U4937 (N_4937,N_4217,N_4318);
nor U4938 (N_4938,N_4548,N_4251);
or U4939 (N_4939,N_4555,N_4530);
nor U4940 (N_4940,N_4586,N_4205);
or U4941 (N_4941,N_4716,N_4588);
and U4942 (N_4942,N_4345,N_4468);
nor U4943 (N_4943,N_4545,N_4767);
or U4944 (N_4944,N_4232,N_4259);
nor U4945 (N_4945,N_4395,N_4340);
nand U4946 (N_4946,N_4405,N_4575);
nor U4947 (N_4947,N_4436,N_4242);
nand U4948 (N_4948,N_4225,N_4538);
and U4949 (N_4949,N_4247,N_4694);
and U4950 (N_4950,N_4347,N_4674);
or U4951 (N_4951,N_4258,N_4605);
and U4952 (N_4952,N_4239,N_4301);
xnor U4953 (N_4953,N_4280,N_4601);
nand U4954 (N_4954,N_4236,N_4294);
or U4955 (N_4955,N_4330,N_4565);
nor U4956 (N_4956,N_4698,N_4715);
nand U4957 (N_4957,N_4414,N_4420);
and U4958 (N_4958,N_4534,N_4721);
xnor U4959 (N_4959,N_4446,N_4342);
or U4960 (N_4960,N_4471,N_4273);
xor U4961 (N_4961,N_4270,N_4693);
nor U4962 (N_4962,N_4482,N_4300);
or U4963 (N_4963,N_4230,N_4370);
and U4964 (N_4964,N_4780,N_4719);
nand U4965 (N_4965,N_4592,N_4246);
xor U4966 (N_4966,N_4375,N_4453);
and U4967 (N_4967,N_4672,N_4394);
and U4968 (N_4968,N_4214,N_4212);
or U4969 (N_4969,N_4201,N_4442);
xnor U4970 (N_4970,N_4402,N_4689);
nor U4971 (N_4971,N_4464,N_4368);
and U4972 (N_4972,N_4419,N_4577);
or U4973 (N_4973,N_4745,N_4799);
nand U4974 (N_4974,N_4204,N_4281);
nor U4975 (N_4975,N_4699,N_4228);
nand U4976 (N_4976,N_4724,N_4303);
nor U4977 (N_4977,N_4392,N_4381);
nor U4978 (N_4978,N_4339,N_4635);
and U4979 (N_4979,N_4252,N_4314);
xor U4980 (N_4980,N_4701,N_4639);
nand U4981 (N_4981,N_4501,N_4610);
or U4982 (N_4982,N_4202,N_4657);
or U4983 (N_4983,N_4320,N_4543);
nor U4984 (N_4984,N_4713,N_4248);
nand U4985 (N_4985,N_4786,N_4308);
or U4986 (N_4986,N_4773,N_4316);
or U4987 (N_4987,N_4429,N_4409);
and U4988 (N_4988,N_4573,N_4778);
xor U4989 (N_4989,N_4754,N_4351);
nand U4990 (N_4990,N_4581,N_4327);
xnor U4991 (N_4991,N_4379,N_4260);
nor U4992 (N_4992,N_4359,N_4406);
xnor U4993 (N_4993,N_4539,N_4380);
or U4994 (N_4994,N_4229,N_4362);
xor U4995 (N_4995,N_4472,N_4680);
and U4996 (N_4996,N_4557,N_4774);
nor U4997 (N_4997,N_4321,N_4483);
nand U4998 (N_4998,N_4628,N_4697);
nor U4999 (N_4999,N_4551,N_4704);
and U5000 (N_5000,N_4598,N_4502);
nor U5001 (N_5001,N_4208,N_4323);
nor U5002 (N_5002,N_4448,N_4643);
and U5003 (N_5003,N_4725,N_4480);
and U5004 (N_5004,N_4499,N_4344);
nand U5005 (N_5005,N_4647,N_4371);
xnor U5006 (N_5006,N_4476,N_4572);
nand U5007 (N_5007,N_4550,N_4469);
nor U5008 (N_5008,N_4421,N_4583);
or U5009 (N_5009,N_4568,N_4310);
nor U5010 (N_5010,N_4624,N_4290);
xnor U5011 (N_5011,N_4566,N_4386);
and U5012 (N_5012,N_4787,N_4536);
nor U5013 (N_5013,N_4289,N_4732);
or U5014 (N_5014,N_4560,N_4681);
nand U5015 (N_5015,N_4510,N_4328);
and U5016 (N_5016,N_4473,N_4747);
or U5017 (N_5017,N_4215,N_4673);
or U5018 (N_5018,N_4517,N_4219);
xnor U5019 (N_5019,N_4798,N_4353);
xnor U5020 (N_5020,N_4554,N_4389);
nand U5021 (N_5021,N_4487,N_4256);
and U5022 (N_5022,N_4632,N_4295);
xnor U5023 (N_5023,N_4210,N_4415);
and U5024 (N_5024,N_4369,N_4490);
nand U5025 (N_5025,N_4385,N_4223);
nand U5026 (N_5026,N_4250,N_4474);
nor U5027 (N_5027,N_4659,N_4355);
or U5028 (N_5028,N_4790,N_4763);
and U5029 (N_5029,N_4785,N_4677);
xnor U5030 (N_5030,N_4726,N_4631);
nor U5031 (N_5031,N_4460,N_4284);
nand U5032 (N_5032,N_4459,N_4796);
nor U5033 (N_5033,N_4227,N_4358);
nand U5034 (N_5034,N_4558,N_4777);
nor U5035 (N_5035,N_4410,N_4769);
xnor U5036 (N_5036,N_4467,N_4602);
and U5037 (N_5037,N_4617,N_4652);
or U5038 (N_5038,N_4707,N_4404);
or U5039 (N_5039,N_4495,N_4296);
xor U5040 (N_5040,N_4542,N_4570);
xor U5041 (N_5041,N_4470,N_4493);
nor U5042 (N_5042,N_4263,N_4304);
nor U5043 (N_5043,N_4437,N_4522);
xnor U5044 (N_5044,N_4319,N_4512);
or U5045 (N_5045,N_4661,N_4612);
nor U5046 (N_5046,N_4312,N_4664);
nand U5047 (N_5047,N_4317,N_4361);
nand U5048 (N_5048,N_4491,N_4708);
or U5049 (N_5049,N_4341,N_4749);
nand U5050 (N_5050,N_4398,N_4636);
nand U5051 (N_5051,N_4513,N_4561);
or U5052 (N_5052,N_4761,N_4336);
or U5053 (N_5053,N_4422,N_4684);
nand U5054 (N_5054,N_4691,N_4562);
xnor U5055 (N_5055,N_4307,N_4656);
xnor U5056 (N_5056,N_4571,N_4779);
or U5057 (N_5057,N_4434,N_4758);
xor U5058 (N_5058,N_4587,N_4614);
nor U5059 (N_5059,N_4776,N_4209);
nand U5060 (N_5060,N_4455,N_4267);
or U5061 (N_5061,N_4220,N_4349);
or U5062 (N_5062,N_4649,N_4648);
nor U5063 (N_5063,N_4298,N_4206);
and U5064 (N_5064,N_4343,N_4441);
nor U5065 (N_5065,N_4722,N_4644);
xnor U5066 (N_5066,N_4498,N_4249);
and U5067 (N_5067,N_4413,N_4611);
nor U5068 (N_5068,N_4357,N_4629);
or U5069 (N_5069,N_4397,N_4702);
and U5070 (N_5070,N_4736,N_4683);
or U5071 (N_5071,N_4291,N_4670);
and U5072 (N_5072,N_4744,N_4486);
xor U5073 (N_5073,N_4213,N_4793);
xnor U5074 (N_5074,N_4727,N_4297);
nand U5075 (N_5075,N_4253,N_4418);
nand U5076 (N_5076,N_4755,N_4218);
nand U5077 (N_5077,N_4509,N_4285);
and U5078 (N_5078,N_4234,N_4703);
xor U5079 (N_5079,N_4516,N_4654);
nand U5080 (N_5080,N_4741,N_4269);
xnor U5081 (N_5081,N_4411,N_4619);
or U5082 (N_5082,N_4784,N_4457);
or U5083 (N_5083,N_4433,N_4496);
and U5084 (N_5084,N_4733,N_4466);
nand U5085 (N_5085,N_4503,N_4622);
xor U5086 (N_5086,N_4593,N_4663);
and U5087 (N_5087,N_4700,N_4346);
xor U5088 (N_5088,N_4791,N_4348);
nand U5089 (N_5089,N_4387,N_4335);
and U5090 (N_5090,N_4731,N_4613);
and U5091 (N_5091,N_4238,N_4233);
or U5092 (N_5092,N_4352,N_4642);
nor U5093 (N_5093,N_4293,N_4506);
or U5094 (N_5094,N_4378,N_4439);
nor U5095 (N_5095,N_4302,N_4423);
xor U5096 (N_5096,N_4484,N_4372);
nand U5097 (N_5097,N_4481,N_4599);
nor U5098 (N_5098,N_4687,N_4401);
xor U5099 (N_5099,N_4254,N_4356);
or U5100 (N_5100,N_4675,N_4711);
and U5101 (N_5101,N_4248,N_4583);
nand U5102 (N_5102,N_4778,N_4261);
and U5103 (N_5103,N_4514,N_4786);
and U5104 (N_5104,N_4725,N_4626);
xnor U5105 (N_5105,N_4683,N_4636);
and U5106 (N_5106,N_4259,N_4681);
or U5107 (N_5107,N_4574,N_4413);
xnor U5108 (N_5108,N_4269,N_4271);
xnor U5109 (N_5109,N_4768,N_4368);
or U5110 (N_5110,N_4553,N_4659);
xnor U5111 (N_5111,N_4366,N_4406);
xor U5112 (N_5112,N_4306,N_4770);
and U5113 (N_5113,N_4222,N_4524);
or U5114 (N_5114,N_4348,N_4210);
or U5115 (N_5115,N_4332,N_4413);
xor U5116 (N_5116,N_4264,N_4688);
nand U5117 (N_5117,N_4442,N_4510);
or U5118 (N_5118,N_4743,N_4644);
xor U5119 (N_5119,N_4404,N_4554);
nand U5120 (N_5120,N_4657,N_4235);
or U5121 (N_5121,N_4242,N_4228);
xnor U5122 (N_5122,N_4396,N_4378);
xor U5123 (N_5123,N_4260,N_4263);
nor U5124 (N_5124,N_4392,N_4720);
nor U5125 (N_5125,N_4755,N_4317);
xor U5126 (N_5126,N_4594,N_4600);
and U5127 (N_5127,N_4484,N_4321);
or U5128 (N_5128,N_4290,N_4406);
and U5129 (N_5129,N_4455,N_4634);
xor U5130 (N_5130,N_4770,N_4760);
nor U5131 (N_5131,N_4795,N_4526);
nand U5132 (N_5132,N_4615,N_4595);
nor U5133 (N_5133,N_4543,N_4709);
nand U5134 (N_5134,N_4319,N_4292);
nand U5135 (N_5135,N_4590,N_4349);
and U5136 (N_5136,N_4778,N_4497);
nor U5137 (N_5137,N_4369,N_4381);
and U5138 (N_5138,N_4671,N_4720);
nor U5139 (N_5139,N_4709,N_4518);
nor U5140 (N_5140,N_4344,N_4571);
and U5141 (N_5141,N_4381,N_4653);
nor U5142 (N_5142,N_4760,N_4764);
xor U5143 (N_5143,N_4724,N_4339);
nor U5144 (N_5144,N_4401,N_4554);
xor U5145 (N_5145,N_4614,N_4406);
or U5146 (N_5146,N_4568,N_4216);
nand U5147 (N_5147,N_4206,N_4597);
nand U5148 (N_5148,N_4250,N_4370);
or U5149 (N_5149,N_4510,N_4645);
xor U5150 (N_5150,N_4264,N_4436);
or U5151 (N_5151,N_4299,N_4784);
xnor U5152 (N_5152,N_4270,N_4787);
nor U5153 (N_5153,N_4703,N_4559);
and U5154 (N_5154,N_4348,N_4473);
and U5155 (N_5155,N_4552,N_4532);
nand U5156 (N_5156,N_4654,N_4727);
and U5157 (N_5157,N_4728,N_4602);
nor U5158 (N_5158,N_4565,N_4521);
nor U5159 (N_5159,N_4230,N_4777);
nor U5160 (N_5160,N_4315,N_4429);
nand U5161 (N_5161,N_4436,N_4600);
or U5162 (N_5162,N_4659,N_4757);
nor U5163 (N_5163,N_4549,N_4660);
nor U5164 (N_5164,N_4432,N_4355);
or U5165 (N_5165,N_4361,N_4698);
and U5166 (N_5166,N_4269,N_4757);
and U5167 (N_5167,N_4237,N_4514);
or U5168 (N_5168,N_4557,N_4561);
nand U5169 (N_5169,N_4531,N_4723);
xor U5170 (N_5170,N_4750,N_4251);
and U5171 (N_5171,N_4582,N_4783);
nor U5172 (N_5172,N_4743,N_4737);
nor U5173 (N_5173,N_4479,N_4604);
and U5174 (N_5174,N_4369,N_4628);
xor U5175 (N_5175,N_4703,N_4640);
and U5176 (N_5176,N_4321,N_4344);
nor U5177 (N_5177,N_4751,N_4737);
and U5178 (N_5178,N_4254,N_4751);
or U5179 (N_5179,N_4750,N_4797);
nor U5180 (N_5180,N_4418,N_4351);
nor U5181 (N_5181,N_4796,N_4203);
xnor U5182 (N_5182,N_4751,N_4685);
or U5183 (N_5183,N_4319,N_4759);
xor U5184 (N_5184,N_4290,N_4368);
nand U5185 (N_5185,N_4437,N_4783);
or U5186 (N_5186,N_4351,N_4642);
xor U5187 (N_5187,N_4406,N_4385);
xor U5188 (N_5188,N_4489,N_4228);
nand U5189 (N_5189,N_4581,N_4267);
nand U5190 (N_5190,N_4465,N_4482);
or U5191 (N_5191,N_4552,N_4488);
xnor U5192 (N_5192,N_4516,N_4378);
nand U5193 (N_5193,N_4221,N_4311);
nor U5194 (N_5194,N_4588,N_4718);
nor U5195 (N_5195,N_4297,N_4254);
and U5196 (N_5196,N_4454,N_4253);
nor U5197 (N_5197,N_4672,N_4547);
and U5198 (N_5198,N_4548,N_4560);
xnor U5199 (N_5199,N_4472,N_4287);
and U5200 (N_5200,N_4293,N_4743);
nand U5201 (N_5201,N_4436,N_4276);
or U5202 (N_5202,N_4529,N_4650);
nand U5203 (N_5203,N_4249,N_4693);
and U5204 (N_5204,N_4217,N_4793);
and U5205 (N_5205,N_4771,N_4315);
nor U5206 (N_5206,N_4540,N_4651);
nand U5207 (N_5207,N_4651,N_4513);
xor U5208 (N_5208,N_4384,N_4410);
or U5209 (N_5209,N_4619,N_4355);
nand U5210 (N_5210,N_4234,N_4786);
nand U5211 (N_5211,N_4244,N_4240);
nor U5212 (N_5212,N_4485,N_4557);
xnor U5213 (N_5213,N_4756,N_4772);
and U5214 (N_5214,N_4563,N_4346);
xnor U5215 (N_5215,N_4547,N_4608);
nand U5216 (N_5216,N_4691,N_4565);
and U5217 (N_5217,N_4736,N_4526);
and U5218 (N_5218,N_4733,N_4228);
xor U5219 (N_5219,N_4247,N_4261);
and U5220 (N_5220,N_4542,N_4425);
or U5221 (N_5221,N_4416,N_4780);
nand U5222 (N_5222,N_4679,N_4283);
or U5223 (N_5223,N_4498,N_4607);
nor U5224 (N_5224,N_4754,N_4255);
and U5225 (N_5225,N_4742,N_4502);
nand U5226 (N_5226,N_4335,N_4357);
xor U5227 (N_5227,N_4714,N_4551);
nand U5228 (N_5228,N_4519,N_4637);
xor U5229 (N_5229,N_4665,N_4433);
nand U5230 (N_5230,N_4327,N_4404);
and U5231 (N_5231,N_4715,N_4708);
or U5232 (N_5232,N_4613,N_4761);
xnor U5233 (N_5233,N_4342,N_4418);
nor U5234 (N_5234,N_4313,N_4748);
and U5235 (N_5235,N_4623,N_4387);
xnor U5236 (N_5236,N_4573,N_4334);
nand U5237 (N_5237,N_4540,N_4657);
xnor U5238 (N_5238,N_4381,N_4624);
or U5239 (N_5239,N_4263,N_4515);
nor U5240 (N_5240,N_4414,N_4653);
nor U5241 (N_5241,N_4456,N_4308);
and U5242 (N_5242,N_4402,N_4716);
or U5243 (N_5243,N_4720,N_4243);
nor U5244 (N_5244,N_4773,N_4306);
nor U5245 (N_5245,N_4558,N_4678);
or U5246 (N_5246,N_4741,N_4219);
nor U5247 (N_5247,N_4256,N_4200);
nor U5248 (N_5248,N_4621,N_4741);
xnor U5249 (N_5249,N_4620,N_4390);
and U5250 (N_5250,N_4467,N_4236);
nor U5251 (N_5251,N_4270,N_4724);
xor U5252 (N_5252,N_4200,N_4540);
or U5253 (N_5253,N_4523,N_4454);
or U5254 (N_5254,N_4347,N_4503);
and U5255 (N_5255,N_4264,N_4502);
and U5256 (N_5256,N_4786,N_4407);
and U5257 (N_5257,N_4556,N_4303);
nand U5258 (N_5258,N_4483,N_4242);
nor U5259 (N_5259,N_4247,N_4778);
xor U5260 (N_5260,N_4724,N_4694);
or U5261 (N_5261,N_4309,N_4403);
nor U5262 (N_5262,N_4506,N_4266);
nand U5263 (N_5263,N_4696,N_4645);
and U5264 (N_5264,N_4725,N_4520);
and U5265 (N_5265,N_4648,N_4270);
xor U5266 (N_5266,N_4516,N_4562);
and U5267 (N_5267,N_4364,N_4688);
or U5268 (N_5268,N_4241,N_4792);
nand U5269 (N_5269,N_4755,N_4529);
xnor U5270 (N_5270,N_4266,N_4503);
xnor U5271 (N_5271,N_4385,N_4436);
and U5272 (N_5272,N_4767,N_4615);
nand U5273 (N_5273,N_4381,N_4604);
nand U5274 (N_5274,N_4203,N_4668);
nor U5275 (N_5275,N_4478,N_4701);
nor U5276 (N_5276,N_4726,N_4731);
and U5277 (N_5277,N_4643,N_4275);
nor U5278 (N_5278,N_4665,N_4277);
xor U5279 (N_5279,N_4223,N_4439);
and U5280 (N_5280,N_4755,N_4209);
and U5281 (N_5281,N_4272,N_4464);
xor U5282 (N_5282,N_4692,N_4488);
nor U5283 (N_5283,N_4523,N_4399);
nand U5284 (N_5284,N_4419,N_4344);
and U5285 (N_5285,N_4686,N_4544);
nand U5286 (N_5286,N_4223,N_4699);
nand U5287 (N_5287,N_4319,N_4615);
xnor U5288 (N_5288,N_4260,N_4459);
nand U5289 (N_5289,N_4435,N_4462);
or U5290 (N_5290,N_4281,N_4714);
xnor U5291 (N_5291,N_4657,N_4528);
nand U5292 (N_5292,N_4495,N_4277);
nand U5293 (N_5293,N_4407,N_4599);
or U5294 (N_5294,N_4722,N_4640);
nor U5295 (N_5295,N_4382,N_4733);
nor U5296 (N_5296,N_4209,N_4560);
and U5297 (N_5297,N_4655,N_4516);
or U5298 (N_5298,N_4543,N_4316);
or U5299 (N_5299,N_4517,N_4281);
nor U5300 (N_5300,N_4479,N_4387);
or U5301 (N_5301,N_4427,N_4281);
nand U5302 (N_5302,N_4598,N_4379);
and U5303 (N_5303,N_4230,N_4715);
nand U5304 (N_5304,N_4635,N_4472);
nand U5305 (N_5305,N_4321,N_4228);
nand U5306 (N_5306,N_4508,N_4713);
or U5307 (N_5307,N_4744,N_4283);
nand U5308 (N_5308,N_4258,N_4652);
nor U5309 (N_5309,N_4482,N_4736);
xor U5310 (N_5310,N_4757,N_4455);
xnor U5311 (N_5311,N_4731,N_4569);
and U5312 (N_5312,N_4268,N_4763);
xnor U5313 (N_5313,N_4618,N_4713);
nor U5314 (N_5314,N_4206,N_4403);
xor U5315 (N_5315,N_4565,N_4575);
nor U5316 (N_5316,N_4591,N_4230);
or U5317 (N_5317,N_4309,N_4413);
or U5318 (N_5318,N_4566,N_4763);
nand U5319 (N_5319,N_4297,N_4466);
or U5320 (N_5320,N_4674,N_4422);
and U5321 (N_5321,N_4257,N_4245);
xnor U5322 (N_5322,N_4606,N_4270);
nor U5323 (N_5323,N_4781,N_4570);
nor U5324 (N_5324,N_4324,N_4251);
xor U5325 (N_5325,N_4219,N_4259);
nand U5326 (N_5326,N_4473,N_4761);
and U5327 (N_5327,N_4749,N_4334);
xnor U5328 (N_5328,N_4470,N_4613);
and U5329 (N_5329,N_4609,N_4607);
xnor U5330 (N_5330,N_4707,N_4393);
nor U5331 (N_5331,N_4607,N_4669);
or U5332 (N_5332,N_4764,N_4781);
and U5333 (N_5333,N_4363,N_4525);
and U5334 (N_5334,N_4425,N_4704);
xnor U5335 (N_5335,N_4444,N_4421);
nand U5336 (N_5336,N_4733,N_4386);
or U5337 (N_5337,N_4399,N_4234);
nor U5338 (N_5338,N_4399,N_4741);
nand U5339 (N_5339,N_4383,N_4785);
nor U5340 (N_5340,N_4254,N_4684);
nand U5341 (N_5341,N_4670,N_4225);
nand U5342 (N_5342,N_4543,N_4746);
or U5343 (N_5343,N_4268,N_4367);
xnor U5344 (N_5344,N_4307,N_4557);
and U5345 (N_5345,N_4434,N_4797);
and U5346 (N_5346,N_4762,N_4626);
and U5347 (N_5347,N_4279,N_4533);
nor U5348 (N_5348,N_4733,N_4425);
nor U5349 (N_5349,N_4684,N_4687);
nand U5350 (N_5350,N_4204,N_4253);
nor U5351 (N_5351,N_4405,N_4666);
or U5352 (N_5352,N_4419,N_4773);
or U5353 (N_5353,N_4395,N_4221);
or U5354 (N_5354,N_4628,N_4623);
xor U5355 (N_5355,N_4527,N_4744);
and U5356 (N_5356,N_4558,N_4254);
nor U5357 (N_5357,N_4261,N_4509);
and U5358 (N_5358,N_4473,N_4343);
and U5359 (N_5359,N_4530,N_4768);
and U5360 (N_5360,N_4768,N_4440);
xnor U5361 (N_5361,N_4476,N_4780);
nand U5362 (N_5362,N_4375,N_4565);
nor U5363 (N_5363,N_4392,N_4203);
and U5364 (N_5364,N_4285,N_4647);
xor U5365 (N_5365,N_4354,N_4512);
nor U5366 (N_5366,N_4566,N_4431);
nand U5367 (N_5367,N_4550,N_4298);
and U5368 (N_5368,N_4744,N_4336);
nor U5369 (N_5369,N_4286,N_4780);
xor U5370 (N_5370,N_4390,N_4717);
and U5371 (N_5371,N_4266,N_4278);
or U5372 (N_5372,N_4537,N_4504);
nor U5373 (N_5373,N_4519,N_4565);
xnor U5374 (N_5374,N_4308,N_4646);
nor U5375 (N_5375,N_4585,N_4300);
xor U5376 (N_5376,N_4619,N_4507);
nand U5377 (N_5377,N_4606,N_4554);
xor U5378 (N_5378,N_4302,N_4461);
xnor U5379 (N_5379,N_4582,N_4661);
nand U5380 (N_5380,N_4495,N_4381);
nand U5381 (N_5381,N_4521,N_4375);
and U5382 (N_5382,N_4335,N_4715);
and U5383 (N_5383,N_4518,N_4261);
or U5384 (N_5384,N_4540,N_4296);
or U5385 (N_5385,N_4544,N_4287);
and U5386 (N_5386,N_4464,N_4616);
or U5387 (N_5387,N_4291,N_4736);
nand U5388 (N_5388,N_4553,N_4460);
nand U5389 (N_5389,N_4406,N_4515);
xnor U5390 (N_5390,N_4678,N_4389);
and U5391 (N_5391,N_4510,N_4582);
and U5392 (N_5392,N_4445,N_4492);
or U5393 (N_5393,N_4621,N_4605);
or U5394 (N_5394,N_4333,N_4551);
xnor U5395 (N_5395,N_4779,N_4243);
or U5396 (N_5396,N_4470,N_4390);
xor U5397 (N_5397,N_4260,N_4542);
xnor U5398 (N_5398,N_4648,N_4736);
and U5399 (N_5399,N_4373,N_4523);
nor U5400 (N_5400,N_5049,N_4908);
nor U5401 (N_5401,N_5067,N_5153);
nor U5402 (N_5402,N_5372,N_5103);
nand U5403 (N_5403,N_4846,N_4822);
nor U5404 (N_5404,N_5283,N_5134);
or U5405 (N_5405,N_4857,N_5314);
xnor U5406 (N_5406,N_5257,N_5070);
nor U5407 (N_5407,N_5368,N_5076);
and U5408 (N_5408,N_4845,N_4906);
nor U5409 (N_5409,N_4803,N_5141);
xnor U5410 (N_5410,N_5385,N_5349);
nor U5411 (N_5411,N_5165,N_5003);
or U5412 (N_5412,N_5244,N_5102);
and U5413 (N_5413,N_5362,N_5233);
or U5414 (N_5414,N_5156,N_5116);
or U5415 (N_5415,N_5159,N_5021);
nand U5416 (N_5416,N_5277,N_5062);
nor U5417 (N_5417,N_5389,N_5051);
and U5418 (N_5418,N_4867,N_4933);
or U5419 (N_5419,N_5011,N_5230);
or U5420 (N_5420,N_5353,N_5327);
or U5421 (N_5421,N_5128,N_5221);
and U5422 (N_5422,N_4999,N_5295);
xnor U5423 (N_5423,N_5239,N_5009);
xor U5424 (N_5424,N_4823,N_5114);
nand U5425 (N_5425,N_5130,N_4863);
nand U5426 (N_5426,N_5319,N_5175);
xor U5427 (N_5427,N_4990,N_5286);
and U5428 (N_5428,N_4888,N_5182);
nand U5429 (N_5429,N_4947,N_4972);
or U5430 (N_5430,N_5088,N_4878);
nor U5431 (N_5431,N_4875,N_5273);
nand U5432 (N_5432,N_5058,N_4966);
nor U5433 (N_5433,N_5198,N_5187);
and U5434 (N_5434,N_5201,N_5267);
and U5435 (N_5435,N_5325,N_4930);
nor U5436 (N_5436,N_5043,N_5111);
nand U5437 (N_5437,N_5075,N_5005);
xnor U5438 (N_5438,N_5214,N_4953);
or U5439 (N_5439,N_4926,N_4948);
and U5440 (N_5440,N_4929,N_4979);
nand U5441 (N_5441,N_5074,N_4848);
nor U5442 (N_5442,N_4873,N_5316);
xor U5443 (N_5443,N_5265,N_4812);
nand U5444 (N_5444,N_4833,N_5154);
xnor U5445 (N_5445,N_5350,N_5369);
nand U5446 (N_5446,N_5227,N_4935);
xor U5447 (N_5447,N_5176,N_5363);
xnor U5448 (N_5448,N_4963,N_4861);
nor U5449 (N_5449,N_5259,N_4956);
xor U5450 (N_5450,N_5019,N_5066);
or U5451 (N_5451,N_5162,N_4837);
nor U5452 (N_5452,N_5004,N_5234);
xor U5453 (N_5453,N_5183,N_5301);
nand U5454 (N_5454,N_4959,N_4946);
nand U5455 (N_5455,N_5121,N_5331);
and U5456 (N_5456,N_5205,N_5192);
or U5457 (N_5457,N_5335,N_5324);
and U5458 (N_5458,N_5377,N_4944);
xnor U5459 (N_5459,N_5135,N_5376);
xnor U5460 (N_5460,N_4968,N_5367);
xor U5461 (N_5461,N_5247,N_5077);
or U5462 (N_5462,N_4923,N_4869);
nor U5463 (N_5463,N_4905,N_5091);
or U5464 (N_5464,N_4992,N_4996);
nor U5465 (N_5465,N_5072,N_4917);
nand U5466 (N_5466,N_5087,N_5242);
nand U5467 (N_5467,N_5379,N_5359);
nand U5468 (N_5468,N_4899,N_5297);
nand U5469 (N_5469,N_5226,N_5137);
and U5470 (N_5470,N_5123,N_5306);
xor U5471 (N_5471,N_4913,N_5012);
nor U5472 (N_5472,N_5032,N_4919);
nand U5473 (N_5473,N_5080,N_5022);
xnor U5474 (N_5474,N_5191,N_5215);
nor U5475 (N_5475,N_4891,N_5023);
nand U5476 (N_5476,N_5048,N_5108);
or U5477 (N_5477,N_5388,N_5199);
and U5478 (N_5478,N_4824,N_5168);
nand U5479 (N_5479,N_5133,N_5181);
xnor U5480 (N_5480,N_5232,N_5180);
nor U5481 (N_5481,N_5309,N_4800);
nor U5482 (N_5482,N_4862,N_5185);
nor U5483 (N_5483,N_5036,N_4811);
nor U5484 (N_5484,N_4872,N_4850);
nand U5485 (N_5485,N_4886,N_5039);
nor U5486 (N_5486,N_5293,N_4967);
or U5487 (N_5487,N_5202,N_5041);
xnor U5488 (N_5488,N_5042,N_5188);
nand U5489 (N_5489,N_4969,N_5261);
xnor U5490 (N_5490,N_5236,N_4849);
and U5491 (N_5491,N_5308,N_5276);
nor U5492 (N_5492,N_4957,N_5024);
nor U5493 (N_5493,N_4808,N_4909);
nand U5494 (N_5494,N_4907,N_4955);
or U5495 (N_5495,N_5000,N_4882);
and U5496 (N_5496,N_5063,N_5345);
and U5497 (N_5497,N_5107,N_4835);
nor U5498 (N_5498,N_5392,N_5352);
nand U5499 (N_5499,N_4897,N_5381);
nand U5500 (N_5500,N_5157,N_5222);
xnor U5501 (N_5501,N_5290,N_5375);
or U5502 (N_5502,N_4874,N_4920);
nor U5503 (N_5503,N_5330,N_5251);
nand U5504 (N_5504,N_5149,N_5069);
nor U5505 (N_5505,N_4815,N_5161);
or U5506 (N_5506,N_5373,N_5015);
nor U5507 (N_5507,N_5120,N_5364);
xnor U5508 (N_5508,N_4937,N_5253);
nor U5509 (N_5509,N_5173,N_4806);
or U5510 (N_5510,N_5053,N_5194);
xor U5511 (N_5511,N_4939,N_5101);
nor U5512 (N_5512,N_4854,N_5317);
or U5513 (N_5513,N_5361,N_4988);
nand U5514 (N_5514,N_5384,N_5167);
nand U5515 (N_5515,N_5278,N_5390);
xnor U5516 (N_5516,N_4981,N_5177);
nor U5517 (N_5517,N_4901,N_5347);
or U5518 (N_5518,N_5189,N_4973);
nand U5519 (N_5519,N_4847,N_5184);
and U5520 (N_5520,N_5034,N_5397);
nand U5521 (N_5521,N_5081,N_4989);
and U5522 (N_5522,N_5050,N_5395);
nand U5523 (N_5523,N_5115,N_5264);
and U5524 (N_5524,N_5303,N_5139);
nand U5525 (N_5525,N_5315,N_5071);
nand U5526 (N_5526,N_5240,N_5068);
nor U5527 (N_5527,N_5179,N_4830);
or U5528 (N_5528,N_5010,N_5002);
nor U5529 (N_5529,N_5144,N_4997);
and U5530 (N_5530,N_4995,N_5046);
or U5531 (N_5531,N_5279,N_5100);
nand U5532 (N_5532,N_5171,N_5085);
nor U5533 (N_5533,N_5346,N_4820);
and U5534 (N_5534,N_4827,N_5031);
nor U5535 (N_5535,N_5001,N_5035);
and U5536 (N_5536,N_5030,N_5125);
nor U5537 (N_5537,N_5095,N_5151);
and U5538 (N_5538,N_5274,N_5086);
xor U5539 (N_5539,N_5126,N_5055);
nand U5540 (N_5540,N_5145,N_4838);
nor U5541 (N_5541,N_5332,N_4994);
or U5542 (N_5542,N_5097,N_5148);
and U5543 (N_5543,N_5132,N_5344);
xor U5544 (N_5544,N_5294,N_5398);
xnor U5545 (N_5545,N_4802,N_5322);
xor U5546 (N_5546,N_5280,N_5163);
nor U5547 (N_5547,N_5170,N_4950);
nor U5548 (N_5548,N_5174,N_4965);
or U5549 (N_5549,N_5318,N_5219);
and U5550 (N_5550,N_5106,N_5288);
and U5551 (N_5551,N_5027,N_4851);
xnor U5552 (N_5552,N_4918,N_4977);
nand U5553 (N_5553,N_4986,N_5225);
nor U5554 (N_5554,N_4952,N_5186);
xor U5555 (N_5555,N_5136,N_5037);
nand U5556 (N_5556,N_4921,N_5224);
xor U5557 (N_5557,N_4978,N_5203);
and U5558 (N_5558,N_5339,N_5358);
xnor U5559 (N_5559,N_5117,N_5040);
or U5560 (N_5560,N_5266,N_4817);
nor U5561 (N_5561,N_4880,N_5272);
xor U5562 (N_5562,N_5371,N_4943);
or U5563 (N_5563,N_4971,N_5237);
or U5564 (N_5564,N_5052,N_5256);
nand U5565 (N_5565,N_5217,N_4982);
or U5566 (N_5566,N_5380,N_4893);
xor U5567 (N_5567,N_4951,N_4819);
nand U5568 (N_5568,N_5296,N_5311);
xor U5569 (N_5569,N_5155,N_4914);
xnor U5570 (N_5570,N_4980,N_5124);
or U5571 (N_5571,N_5083,N_4964);
xor U5572 (N_5572,N_5248,N_5218);
nand U5573 (N_5573,N_5018,N_5228);
nand U5574 (N_5574,N_5158,N_5033);
or U5575 (N_5575,N_5337,N_5146);
or U5576 (N_5576,N_5017,N_4871);
nor U5577 (N_5577,N_4836,N_5223);
and U5578 (N_5578,N_4832,N_5268);
nand U5579 (N_5579,N_5338,N_5143);
nor U5580 (N_5580,N_4804,N_5064);
nor U5581 (N_5581,N_4879,N_5044);
xnor U5582 (N_5582,N_4993,N_5235);
nor U5583 (N_5583,N_4805,N_5246);
and U5584 (N_5584,N_5321,N_4958);
and U5585 (N_5585,N_5310,N_4866);
nand U5586 (N_5586,N_5200,N_5038);
and U5587 (N_5587,N_4931,N_5211);
xor U5588 (N_5588,N_4976,N_4974);
xor U5589 (N_5589,N_4825,N_4916);
nand U5590 (N_5590,N_5008,N_4900);
nand U5591 (N_5591,N_5355,N_5399);
nand U5592 (N_5592,N_4928,N_5104);
nor U5593 (N_5593,N_5013,N_4881);
nand U5594 (N_5594,N_5197,N_5127);
and U5595 (N_5595,N_4936,N_5082);
and U5596 (N_5596,N_4885,N_4960);
or U5597 (N_5597,N_5269,N_5393);
nand U5598 (N_5598,N_5357,N_5020);
xnor U5599 (N_5599,N_5014,N_5370);
or U5600 (N_5600,N_5275,N_5300);
xnor U5601 (N_5601,N_4984,N_4975);
nor U5602 (N_5602,N_5061,N_5229);
nand U5603 (N_5603,N_5210,N_4841);
xor U5604 (N_5604,N_5340,N_4889);
nor U5605 (N_5605,N_5118,N_4940);
nand U5606 (N_5606,N_5207,N_5099);
and U5607 (N_5607,N_5282,N_5178);
xor U5608 (N_5608,N_5360,N_5094);
nand U5609 (N_5609,N_5193,N_4895);
xnor U5610 (N_5610,N_5336,N_5260);
or U5611 (N_5611,N_4927,N_4987);
or U5612 (N_5612,N_5354,N_4954);
or U5613 (N_5613,N_5394,N_4904);
xnor U5614 (N_5614,N_4932,N_5152);
xnor U5615 (N_5615,N_4902,N_4887);
or U5616 (N_5616,N_4945,N_5245);
xor U5617 (N_5617,N_5320,N_4810);
or U5618 (N_5618,N_5304,N_4962);
or U5619 (N_5619,N_5334,N_5351);
xnor U5620 (N_5620,N_5383,N_5029);
and U5621 (N_5621,N_5238,N_4844);
nor U5622 (N_5622,N_5323,N_4884);
xor U5623 (N_5623,N_5307,N_4831);
and U5624 (N_5624,N_5284,N_5092);
nand U5625 (N_5625,N_4898,N_5119);
or U5626 (N_5626,N_4839,N_4870);
and U5627 (N_5627,N_5328,N_4859);
or U5628 (N_5628,N_4843,N_4868);
nor U5629 (N_5629,N_4852,N_5382);
and U5630 (N_5630,N_4856,N_5090);
nor U5631 (N_5631,N_5252,N_4860);
xor U5632 (N_5632,N_5299,N_4991);
nand U5633 (N_5633,N_4998,N_5098);
nor U5634 (N_5634,N_5054,N_4894);
xnor U5635 (N_5635,N_5057,N_5342);
nand U5636 (N_5636,N_5333,N_4876);
xor U5637 (N_5637,N_5166,N_4801);
nand U5638 (N_5638,N_5056,N_5096);
and U5639 (N_5639,N_5045,N_5195);
or U5640 (N_5640,N_4818,N_5305);
xnor U5641 (N_5641,N_4826,N_5190);
nand U5642 (N_5642,N_5255,N_4883);
and U5643 (N_5643,N_4865,N_5026);
and U5644 (N_5644,N_5287,N_5289);
nand U5645 (N_5645,N_4814,N_5391);
or U5646 (N_5646,N_5006,N_4816);
or U5647 (N_5647,N_4985,N_5084);
nor U5648 (N_5648,N_4890,N_5263);
nand U5649 (N_5649,N_4840,N_4807);
nand U5650 (N_5650,N_5249,N_5025);
xnor U5651 (N_5651,N_5112,N_5164);
xnor U5652 (N_5652,N_5213,N_5140);
and U5653 (N_5653,N_5078,N_5220);
and U5654 (N_5654,N_5093,N_5298);
or U5655 (N_5655,N_5073,N_4809);
nand U5656 (N_5656,N_4828,N_5209);
xor U5657 (N_5657,N_4896,N_5204);
or U5658 (N_5658,N_5374,N_5348);
nor U5659 (N_5659,N_4912,N_4961);
nor U5660 (N_5660,N_5241,N_4983);
xnor U5661 (N_5661,N_5131,N_5016);
or U5662 (N_5662,N_5387,N_5216);
nand U5663 (N_5663,N_5312,N_5326);
nor U5664 (N_5664,N_4853,N_5341);
xor U5665 (N_5665,N_5196,N_4858);
or U5666 (N_5666,N_5065,N_5060);
or U5667 (N_5667,N_5386,N_4821);
xor U5668 (N_5668,N_4924,N_4911);
xnor U5669 (N_5669,N_5208,N_5250);
and U5670 (N_5670,N_5231,N_4922);
and U5671 (N_5671,N_5142,N_4934);
nand U5672 (N_5672,N_5285,N_5254);
and U5673 (N_5673,N_5109,N_5329);
and U5674 (N_5674,N_4938,N_5302);
nand U5675 (N_5675,N_5113,N_5079);
nor U5676 (N_5676,N_5281,N_4925);
or U5677 (N_5677,N_4813,N_4834);
xor U5678 (N_5678,N_5059,N_5138);
nor U5679 (N_5679,N_5047,N_5089);
nor U5680 (N_5680,N_5212,N_4915);
and U5681 (N_5681,N_5105,N_4970);
xor U5682 (N_5682,N_4942,N_5366);
xor U5683 (N_5683,N_5262,N_5110);
nand U5684 (N_5684,N_5147,N_4877);
nand U5685 (N_5685,N_4910,N_4941);
xnor U5686 (N_5686,N_5169,N_5396);
nor U5687 (N_5687,N_5150,N_5291);
nand U5688 (N_5688,N_5007,N_5258);
and U5689 (N_5689,N_4855,N_5313);
xor U5690 (N_5690,N_5271,N_5172);
or U5691 (N_5691,N_5129,N_5356);
or U5692 (N_5692,N_5122,N_5365);
nand U5693 (N_5693,N_5160,N_4903);
nor U5694 (N_5694,N_5378,N_5206);
and U5695 (N_5695,N_4864,N_5292);
or U5696 (N_5696,N_4842,N_4829);
nand U5697 (N_5697,N_5028,N_5343);
nand U5698 (N_5698,N_5270,N_4949);
or U5699 (N_5699,N_5243,N_4892);
nand U5700 (N_5700,N_5261,N_5029);
or U5701 (N_5701,N_4967,N_5321);
nor U5702 (N_5702,N_5147,N_4898);
nand U5703 (N_5703,N_4844,N_4852);
and U5704 (N_5704,N_4891,N_4944);
nand U5705 (N_5705,N_5164,N_4895);
nor U5706 (N_5706,N_5334,N_4906);
xnor U5707 (N_5707,N_4906,N_5335);
or U5708 (N_5708,N_5201,N_5165);
and U5709 (N_5709,N_5261,N_4918);
or U5710 (N_5710,N_5279,N_5226);
nor U5711 (N_5711,N_5260,N_5338);
nand U5712 (N_5712,N_4979,N_5368);
nor U5713 (N_5713,N_5203,N_4979);
nand U5714 (N_5714,N_4996,N_4950);
nand U5715 (N_5715,N_5294,N_4991);
and U5716 (N_5716,N_4951,N_5294);
or U5717 (N_5717,N_5348,N_5063);
and U5718 (N_5718,N_5284,N_4911);
or U5719 (N_5719,N_5022,N_5365);
nand U5720 (N_5720,N_5376,N_4964);
nor U5721 (N_5721,N_5202,N_4895);
nor U5722 (N_5722,N_5231,N_4812);
or U5723 (N_5723,N_5319,N_4866);
xor U5724 (N_5724,N_4986,N_4953);
nor U5725 (N_5725,N_4841,N_5322);
xor U5726 (N_5726,N_5127,N_5152);
nor U5727 (N_5727,N_5031,N_5177);
and U5728 (N_5728,N_5088,N_4959);
xnor U5729 (N_5729,N_5267,N_5104);
nor U5730 (N_5730,N_5278,N_5180);
nor U5731 (N_5731,N_5234,N_5209);
or U5732 (N_5732,N_4867,N_4942);
xor U5733 (N_5733,N_5391,N_5064);
xor U5734 (N_5734,N_4921,N_4830);
nor U5735 (N_5735,N_4868,N_5275);
and U5736 (N_5736,N_5243,N_4992);
or U5737 (N_5737,N_5398,N_5289);
xnor U5738 (N_5738,N_5160,N_4978);
nand U5739 (N_5739,N_5241,N_5399);
xnor U5740 (N_5740,N_4933,N_4910);
xor U5741 (N_5741,N_5047,N_5132);
nand U5742 (N_5742,N_5249,N_5189);
or U5743 (N_5743,N_4947,N_5154);
or U5744 (N_5744,N_4996,N_5182);
or U5745 (N_5745,N_5135,N_5109);
nor U5746 (N_5746,N_5326,N_5283);
xor U5747 (N_5747,N_4887,N_5093);
nor U5748 (N_5748,N_4934,N_5082);
nand U5749 (N_5749,N_5284,N_4995);
xor U5750 (N_5750,N_5373,N_5090);
nand U5751 (N_5751,N_4838,N_4951);
nor U5752 (N_5752,N_5066,N_5004);
nand U5753 (N_5753,N_5096,N_4871);
nor U5754 (N_5754,N_4899,N_4991);
nor U5755 (N_5755,N_5283,N_4979);
nand U5756 (N_5756,N_5124,N_4999);
xnor U5757 (N_5757,N_5101,N_5226);
xnor U5758 (N_5758,N_5199,N_5058);
nand U5759 (N_5759,N_4805,N_4949);
xor U5760 (N_5760,N_5115,N_5390);
nand U5761 (N_5761,N_4889,N_5188);
or U5762 (N_5762,N_5138,N_5121);
nor U5763 (N_5763,N_4812,N_4904);
nor U5764 (N_5764,N_5156,N_4888);
or U5765 (N_5765,N_5388,N_5238);
or U5766 (N_5766,N_5125,N_5050);
and U5767 (N_5767,N_5367,N_5086);
and U5768 (N_5768,N_5014,N_5389);
or U5769 (N_5769,N_5071,N_4911);
nand U5770 (N_5770,N_5230,N_5369);
xnor U5771 (N_5771,N_5086,N_4814);
xor U5772 (N_5772,N_4909,N_5009);
or U5773 (N_5773,N_5394,N_5165);
or U5774 (N_5774,N_4914,N_4804);
or U5775 (N_5775,N_5330,N_5297);
and U5776 (N_5776,N_5063,N_5062);
nand U5777 (N_5777,N_5190,N_5339);
nor U5778 (N_5778,N_5174,N_5192);
xor U5779 (N_5779,N_5381,N_5237);
and U5780 (N_5780,N_5147,N_5226);
xnor U5781 (N_5781,N_5198,N_5013);
nand U5782 (N_5782,N_5110,N_4814);
nand U5783 (N_5783,N_4908,N_4983);
or U5784 (N_5784,N_4914,N_5063);
and U5785 (N_5785,N_5381,N_5023);
and U5786 (N_5786,N_5076,N_5045);
or U5787 (N_5787,N_5328,N_4880);
or U5788 (N_5788,N_5114,N_4897);
or U5789 (N_5789,N_5366,N_4880);
nand U5790 (N_5790,N_5391,N_4837);
nor U5791 (N_5791,N_5236,N_4858);
xor U5792 (N_5792,N_4801,N_5251);
nor U5793 (N_5793,N_4832,N_4950);
xnor U5794 (N_5794,N_5019,N_5093);
and U5795 (N_5795,N_4898,N_5299);
xor U5796 (N_5796,N_5283,N_5133);
and U5797 (N_5797,N_5275,N_4969);
or U5798 (N_5798,N_4831,N_5243);
nand U5799 (N_5799,N_4830,N_4850);
nand U5800 (N_5800,N_5244,N_5121);
or U5801 (N_5801,N_4941,N_5397);
nor U5802 (N_5802,N_5045,N_4850);
nor U5803 (N_5803,N_5216,N_5335);
and U5804 (N_5804,N_5372,N_5286);
nand U5805 (N_5805,N_5267,N_5164);
or U5806 (N_5806,N_4829,N_5262);
nor U5807 (N_5807,N_4916,N_5236);
nand U5808 (N_5808,N_5117,N_5156);
or U5809 (N_5809,N_4950,N_5109);
nor U5810 (N_5810,N_5360,N_5271);
or U5811 (N_5811,N_5190,N_4843);
nand U5812 (N_5812,N_4811,N_4835);
xnor U5813 (N_5813,N_5120,N_5031);
xnor U5814 (N_5814,N_5028,N_5340);
or U5815 (N_5815,N_4882,N_5185);
xor U5816 (N_5816,N_5333,N_5145);
or U5817 (N_5817,N_4862,N_5071);
or U5818 (N_5818,N_4923,N_4914);
nor U5819 (N_5819,N_5210,N_4949);
nor U5820 (N_5820,N_5139,N_5369);
and U5821 (N_5821,N_5173,N_4803);
nor U5822 (N_5822,N_5398,N_5077);
and U5823 (N_5823,N_5051,N_4928);
or U5824 (N_5824,N_4927,N_5004);
or U5825 (N_5825,N_5193,N_4855);
and U5826 (N_5826,N_5091,N_4845);
and U5827 (N_5827,N_5260,N_5197);
and U5828 (N_5828,N_5375,N_5354);
and U5829 (N_5829,N_5276,N_4984);
xor U5830 (N_5830,N_5256,N_5389);
nand U5831 (N_5831,N_4905,N_4984);
nor U5832 (N_5832,N_5164,N_5101);
nand U5833 (N_5833,N_4999,N_5357);
nor U5834 (N_5834,N_4940,N_4879);
or U5835 (N_5835,N_5082,N_4896);
xor U5836 (N_5836,N_4809,N_5297);
xor U5837 (N_5837,N_5380,N_5218);
or U5838 (N_5838,N_5333,N_5146);
nand U5839 (N_5839,N_5040,N_5312);
and U5840 (N_5840,N_4828,N_5291);
nand U5841 (N_5841,N_4891,N_5044);
or U5842 (N_5842,N_5042,N_5007);
nor U5843 (N_5843,N_4971,N_5235);
xor U5844 (N_5844,N_5084,N_4806);
xnor U5845 (N_5845,N_4913,N_4950);
or U5846 (N_5846,N_4853,N_4834);
nor U5847 (N_5847,N_5029,N_4929);
or U5848 (N_5848,N_5214,N_5374);
xnor U5849 (N_5849,N_5319,N_5343);
or U5850 (N_5850,N_5019,N_5063);
and U5851 (N_5851,N_4917,N_5314);
xor U5852 (N_5852,N_5293,N_5329);
and U5853 (N_5853,N_5271,N_5019);
or U5854 (N_5854,N_5218,N_4880);
nor U5855 (N_5855,N_5366,N_5351);
and U5856 (N_5856,N_5075,N_5218);
or U5857 (N_5857,N_4941,N_5275);
xnor U5858 (N_5858,N_5101,N_5177);
and U5859 (N_5859,N_5098,N_5255);
xor U5860 (N_5860,N_4928,N_4907);
nand U5861 (N_5861,N_4850,N_4888);
xor U5862 (N_5862,N_5031,N_5299);
xor U5863 (N_5863,N_5200,N_4936);
nor U5864 (N_5864,N_5346,N_5249);
nand U5865 (N_5865,N_4954,N_4858);
nand U5866 (N_5866,N_4809,N_5184);
nand U5867 (N_5867,N_5044,N_4999);
xnor U5868 (N_5868,N_5065,N_5122);
or U5869 (N_5869,N_5018,N_4918);
nor U5870 (N_5870,N_4931,N_5167);
or U5871 (N_5871,N_5199,N_4854);
nor U5872 (N_5872,N_5027,N_5331);
nor U5873 (N_5873,N_4934,N_5055);
and U5874 (N_5874,N_5178,N_4816);
or U5875 (N_5875,N_5153,N_4975);
and U5876 (N_5876,N_4858,N_5153);
nor U5877 (N_5877,N_5307,N_5103);
nor U5878 (N_5878,N_5296,N_5276);
xor U5879 (N_5879,N_5270,N_5208);
or U5880 (N_5880,N_5313,N_5262);
nor U5881 (N_5881,N_5163,N_4828);
or U5882 (N_5882,N_4947,N_5021);
and U5883 (N_5883,N_4927,N_5095);
nand U5884 (N_5884,N_5020,N_5291);
nor U5885 (N_5885,N_5171,N_5158);
and U5886 (N_5886,N_5250,N_5259);
or U5887 (N_5887,N_4978,N_4846);
and U5888 (N_5888,N_4974,N_5040);
xnor U5889 (N_5889,N_5046,N_5379);
xnor U5890 (N_5890,N_5275,N_4926);
and U5891 (N_5891,N_5078,N_5135);
nor U5892 (N_5892,N_4911,N_5340);
or U5893 (N_5893,N_5311,N_5077);
xor U5894 (N_5894,N_5155,N_5312);
and U5895 (N_5895,N_5073,N_5186);
nor U5896 (N_5896,N_5116,N_4817);
or U5897 (N_5897,N_5034,N_4927);
or U5898 (N_5898,N_5206,N_5360);
nor U5899 (N_5899,N_5242,N_5330);
xor U5900 (N_5900,N_5123,N_5289);
nor U5901 (N_5901,N_4886,N_4966);
nor U5902 (N_5902,N_4942,N_4865);
nor U5903 (N_5903,N_5172,N_5304);
and U5904 (N_5904,N_5079,N_5027);
or U5905 (N_5905,N_5008,N_4869);
or U5906 (N_5906,N_4874,N_5174);
and U5907 (N_5907,N_4964,N_5364);
xor U5908 (N_5908,N_5178,N_5313);
nor U5909 (N_5909,N_5396,N_5008);
xnor U5910 (N_5910,N_4801,N_5162);
nor U5911 (N_5911,N_5048,N_5279);
nand U5912 (N_5912,N_5106,N_5281);
and U5913 (N_5913,N_5362,N_5238);
nor U5914 (N_5914,N_4953,N_4974);
and U5915 (N_5915,N_5310,N_5140);
xnor U5916 (N_5916,N_5110,N_4809);
xor U5917 (N_5917,N_5350,N_5353);
and U5918 (N_5918,N_5152,N_5234);
and U5919 (N_5919,N_4942,N_5219);
or U5920 (N_5920,N_5352,N_5150);
xnor U5921 (N_5921,N_5153,N_5133);
or U5922 (N_5922,N_5066,N_5087);
nand U5923 (N_5923,N_5099,N_5090);
or U5924 (N_5924,N_4857,N_5301);
or U5925 (N_5925,N_4979,N_5379);
nand U5926 (N_5926,N_4857,N_5356);
xor U5927 (N_5927,N_5194,N_5132);
nand U5928 (N_5928,N_5218,N_5221);
nand U5929 (N_5929,N_5172,N_5396);
or U5930 (N_5930,N_5021,N_4804);
and U5931 (N_5931,N_5210,N_5045);
or U5932 (N_5932,N_5298,N_4909);
or U5933 (N_5933,N_5134,N_5018);
xor U5934 (N_5934,N_4985,N_5064);
xnor U5935 (N_5935,N_4929,N_5164);
nand U5936 (N_5936,N_5127,N_5001);
and U5937 (N_5937,N_4840,N_5211);
or U5938 (N_5938,N_5156,N_4878);
or U5939 (N_5939,N_5164,N_4995);
and U5940 (N_5940,N_5169,N_5328);
xor U5941 (N_5941,N_5341,N_4889);
xor U5942 (N_5942,N_5278,N_4823);
or U5943 (N_5943,N_5314,N_5015);
xor U5944 (N_5944,N_5127,N_4839);
or U5945 (N_5945,N_5377,N_4979);
and U5946 (N_5946,N_5270,N_5113);
and U5947 (N_5947,N_4991,N_5227);
nand U5948 (N_5948,N_4813,N_5279);
or U5949 (N_5949,N_5260,N_5399);
nand U5950 (N_5950,N_5262,N_5069);
or U5951 (N_5951,N_5271,N_4900);
and U5952 (N_5952,N_5267,N_4906);
or U5953 (N_5953,N_5364,N_5323);
nand U5954 (N_5954,N_5332,N_4990);
xnor U5955 (N_5955,N_5298,N_5191);
nor U5956 (N_5956,N_5024,N_5384);
nand U5957 (N_5957,N_5022,N_5261);
nand U5958 (N_5958,N_5378,N_4852);
xnor U5959 (N_5959,N_4803,N_5155);
or U5960 (N_5960,N_5296,N_5083);
nand U5961 (N_5961,N_4851,N_5094);
nand U5962 (N_5962,N_4877,N_5059);
nor U5963 (N_5963,N_5329,N_5059);
and U5964 (N_5964,N_4822,N_4940);
or U5965 (N_5965,N_5357,N_5242);
or U5966 (N_5966,N_4879,N_5184);
nand U5967 (N_5967,N_5071,N_4976);
nor U5968 (N_5968,N_5366,N_5361);
nand U5969 (N_5969,N_4914,N_5276);
or U5970 (N_5970,N_4949,N_5063);
and U5971 (N_5971,N_5286,N_5330);
and U5972 (N_5972,N_5094,N_5165);
xor U5973 (N_5973,N_4831,N_4865);
nor U5974 (N_5974,N_5141,N_4837);
nand U5975 (N_5975,N_5060,N_5376);
nor U5976 (N_5976,N_4910,N_4852);
or U5977 (N_5977,N_5057,N_5276);
xor U5978 (N_5978,N_4829,N_5056);
or U5979 (N_5979,N_5344,N_5255);
or U5980 (N_5980,N_5387,N_4827);
or U5981 (N_5981,N_5096,N_5107);
nor U5982 (N_5982,N_5193,N_4843);
and U5983 (N_5983,N_4851,N_4965);
and U5984 (N_5984,N_4988,N_5183);
nor U5985 (N_5985,N_5226,N_4883);
and U5986 (N_5986,N_5232,N_4983);
or U5987 (N_5987,N_5345,N_5238);
nand U5988 (N_5988,N_5082,N_5119);
xor U5989 (N_5989,N_4979,N_4899);
and U5990 (N_5990,N_4993,N_5171);
nand U5991 (N_5991,N_5164,N_5292);
xnor U5992 (N_5992,N_5293,N_5163);
xor U5993 (N_5993,N_4849,N_4858);
xnor U5994 (N_5994,N_5173,N_5193);
nor U5995 (N_5995,N_4943,N_5126);
or U5996 (N_5996,N_4894,N_5228);
nor U5997 (N_5997,N_5149,N_5286);
nand U5998 (N_5998,N_4834,N_5308);
or U5999 (N_5999,N_4847,N_5051);
and U6000 (N_6000,N_5766,N_5814);
nor U6001 (N_6001,N_5566,N_5847);
xor U6002 (N_6002,N_5841,N_5874);
and U6003 (N_6003,N_5518,N_5717);
or U6004 (N_6004,N_5999,N_5650);
or U6005 (N_6005,N_5982,N_5969);
and U6006 (N_6006,N_5909,N_5776);
nand U6007 (N_6007,N_5634,N_5586);
or U6008 (N_6008,N_5989,N_5472);
nand U6009 (N_6009,N_5785,N_5689);
nand U6010 (N_6010,N_5535,N_5445);
or U6011 (N_6011,N_5711,N_5452);
nand U6012 (N_6012,N_5401,N_5805);
nand U6013 (N_6013,N_5879,N_5824);
nor U6014 (N_6014,N_5831,N_5896);
nor U6015 (N_6015,N_5778,N_5431);
nand U6016 (N_6016,N_5668,N_5756);
and U6017 (N_6017,N_5434,N_5638);
or U6018 (N_6018,N_5731,N_5440);
nand U6019 (N_6019,N_5605,N_5968);
and U6020 (N_6020,N_5426,N_5536);
or U6021 (N_6021,N_5584,N_5476);
or U6022 (N_6022,N_5642,N_5512);
nor U6023 (N_6023,N_5478,N_5862);
or U6024 (N_6024,N_5744,N_5905);
nand U6025 (N_6025,N_5457,N_5592);
or U6026 (N_6026,N_5780,N_5726);
nor U6027 (N_6027,N_5791,N_5754);
nor U6028 (N_6028,N_5527,N_5549);
xnor U6029 (N_6029,N_5855,N_5406);
nand U6030 (N_6030,N_5661,N_5800);
xor U6031 (N_6031,N_5825,N_5438);
nor U6032 (N_6032,N_5623,N_5444);
nand U6033 (N_6033,N_5593,N_5927);
and U6034 (N_6034,N_5648,N_5891);
and U6035 (N_6035,N_5953,N_5915);
nor U6036 (N_6036,N_5437,N_5657);
nor U6037 (N_6037,N_5410,N_5414);
nor U6038 (N_6038,N_5792,N_5494);
nand U6039 (N_6039,N_5815,N_5483);
nand U6040 (N_6040,N_5424,N_5553);
nand U6041 (N_6041,N_5746,N_5542);
nor U6042 (N_6042,N_5411,N_5501);
and U6043 (N_6043,N_5732,N_5649);
xnor U6044 (N_6044,N_5706,N_5893);
and U6045 (N_6045,N_5933,N_5946);
xor U6046 (N_6046,N_5409,N_5582);
and U6047 (N_6047,N_5930,N_5742);
nand U6048 (N_6048,N_5528,N_5521);
or U6049 (N_6049,N_5774,N_5965);
nor U6050 (N_6050,N_5807,N_5420);
nor U6051 (N_6051,N_5641,N_5954);
nand U6052 (N_6052,N_5902,N_5700);
xnor U6053 (N_6053,N_5773,N_5901);
or U6054 (N_6054,N_5950,N_5975);
xnor U6055 (N_6055,N_5448,N_5898);
xor U6056 (N_6056,N_5727,N_5851);
xnor U6057 (N_6057,N_5809,N_5979);
or U6058 (N_6058,N_5844,N_5629);
and U6059 (N_6059,N_5447,N_5614);
nor U6060 (N_6060,N_5442,N_5561);
nor U6061 (N_6061,N_5906,N_5658);
or U6062 (N_6062,N_5863,N_5552);
and U6063 (N_6063,N_5627,N_5961);
xnor U6064 (N_6064,N_5980,N_5644);
and U6065 (N_6065,N_5798,N_5990);
nand U6066 (N_6066,N_5567,N_5506);
xnor U6067 (N_6067,N_5601,N_5917);
nand U6068 (N_6068,N_5485,N_5720);
and U6069 (N_6069,N_5836,N_5405);
nor U6070 (N_6070,N_5616,N_5753);
xor U6071 (N_6071,N_5760,N_5663);
xnor U6072 (N_6072,N_5579,N_5850);
xor U6073 (N_6073,N_5704,N_5974);
nor U6074 (N_6074,N_5959,N_5861);
and U6075 (N_6075,N_5441,N_5775);
and U6076 (N_6076,N_5908,N_5610);
and U6077 (N_6077,N_5869,N_5443);
nor U6078 (N_6078,N_5956,N_5872);
nor U6079 (N_6079,N_5607,N_5867);
nand U6080 (N_6080,N_5932,N_5958);
nor U6081 (N_6081,N_5783,N_5734);
and U6082 (N_6082,N_5507,N_5517);
xor U6083 (N_6083,N_5964,N_5556);
nand U6084 (N_6084,N_5547,N_5575);
and U6085 (N_6085,N_5903,N_5523);
nor U6086 (N_6086,N_5781,N_5992);
nor U6087 (N_6087,N_5705,N_5671);
xor U6088 (N_6088,N_5515,N_5949);
and U6089 (N_6089,N_5733,N_5460);
and U6090 (N_6090,N_5635,N_5963);
nor U6091 (N_6091,N_5771,N_5462);
nand U6092 (N_6092,N_5839,N_5699);
or U6093 (N_6093,N_5913,N_5900);
nand U6094 (N_6094,N_5660,N_5925);
nand U6095 (N_6095,N_5984,N_5797);
nand U6096 (N_6096,N_5813,N_5695);
nand U6097 (N_6097,N_5533,N_5456);
nor U6098 (N_6098,N_5811,N_5854);
xor U6099 (N_6099,N_5449,N_5966);
nand U6100 (N_6100,N_5577,N_5539);
nand U6101 (N_6101,N_5928,N_5716);
nand U6102 (N_6102,N_5784,N_5779);
nand U6103 (N_6103,N_5425,N_5981);
and U6104 (N_6104,N_5960,N_5670);
nor U6105 (N_6105,N_5866,N_5500);
nor U6106 (N_6106,N_5681,N_5769);
nor U6107 (N_6107,N_5772,N_5739);
xnor U6108 (N_6108,N_5916,N_5599);
and U6109 (N_6109,N_5770,N_5838);
nand U6110 (N_6110,N_5883,N_5823);
nor U6111 (N_6111,N_5531,N_5842);
xor U6112 (N_6112,N_5802,N_5914);
nor U6113 (N_6113,N_5931,N_5691);
and U6114 (N_6114,N_5534,N_5985);
and U6115 (N_6115,N_5688,N_5947);
or U6116 (N_6116,N_5454,N_5759);
and U6117 (N_6117,N_5679,N_5666);
and U6118 (N_6118,N_5569,N_5459);
xor U6119 (N_6119,N_5453,N_5451);
and U6120 (N_6120,N_5557,N_5647);
nor U6121 (N_6121,N_5503,N_5938);
xor U6122 (N_6122,N_5793,N_5479);
nand U6123 (N_6123,N_5765,N_5583);
xnor U6124 (N_6124,N_5899,N_5948);
nor U6125 (N_6125,N_5718,N_5829);
nand U6126 (N_6126,N_5408,N_5646);
nand U6127 (N_6127,N_5543,N_5832);
nor U6128 (N_6128,N_5676,N_5608);
or U6129 (N_6129,N_5762,N_5612);
xor U6130 (N_6130,N_5892,N_5466);
nand U6131 (N_6131,N_5526,N_5574);
nand U6132 (N_6132,N_5555,N_5736);
nand U6133 (N_6133,N_5585,N_5617);
and U6134 (N_6134,N_5645,N_5846);
xor U6135 (N_6135,N_5429,N_5498);
nand U6136 (N_6136,N_5761,N_5816);
and U6137 (N_6137,N_5589,N_5600);
xnor U6138 (N_6138,N_5803,N_5432);
nand U6139 (N_6139,N_5697,N_5568);
or U6140 (N_6140,N_5419,N_5923);
nor U6141 (N_6141,N_5570,N_5516);
xnor U6142 (N_6142,N_5701,N_5853);
nor U6143 (N_6143,N_5745,N_5843);
xnor U6144 (N_6144,N_5482,N_5777);
and U6145 (N_6145,N_5672,N_5693);
nor U6146 (N_6146,N_5943,N_5477);
nand U6147 (N_6147,N_5677,N_5465);
xor U6148 (N_6148,N_5694,N_5464);
nor U6149 (N_6149,N_5828,N_5730);
xnor U6150 (N_6150,N_5496,N_5941);
xnor U6151 (N_6151,N_5991,N_5682);
xnor U6152 (N_6152,N_5976,N_5702);
nor U6153 (N_6153,N_5653,N_5422);
nor U6154 (N_6154,N_5764,N_5722);
nand U6155 (N_6155,N_5835,N_5873);
nand U6156 (N_6156,N_5972,N_5402);
xnor U6157 (N_6157,N_5665,N_5710);
xor U6158 (N_6158,N_5415,N_5509);
xor U6159 (N_6159,N_5446,N_5499);
and U6160 (N_6160,N_5551,N_5911);
nand U6161 (N_6161,N_5619,N_5970);
nor U6162 (N_6162,N_5513,N_5848);
nand U6163 (N_6163,N_5840,N_5725);
and U6164 (N_6164,N_5871,N_5708);
or U6165 (N_6165,N_5882,N_5737);
nor U6166 (N_6166,N_5707,N_5758);
nor U6167 (N_6167,N_5435,N_5428);
or U6168 (N_6168,N_5897,N_5430);
nor U6169 (N_6169,N_5606,N_5573);
nor U6170 (N_6170,N_5510,N_5490);
nor U6171 (N_6171,N_5995,N_5486);
xor U6172 (N_6172,N_5719,N_5436);
or U6173 (N_6173,N_5877,N_5545);
nand U6174 (N_6174,N_5944,N_5819);
or U6175 (N_6175,N_5626,N_5757);
nand U6176 (N_6176,N_5942,N_5469);
xor U6177 (N_6177,N_5998,N_5787);
xor U6178 (N_6178,N_5788,N_5571);
nor U6179 (N_6179,N_5667,N_5935);
and U6180 (N_6180,N_5587,N_5581);
nand U6181 (N_6181,N_5920,N_5878);
nor U6182 (N_6182,N_5541,N_5603);
nand U6183 (N_6183,N_5576,N_5921);
or U6184 (N_6184,N_5590,N_5427);
xor U6185 (N_6185,N_5618,N_5703);
or U6186 (N_6186,N_5678,N_5748);
or U6187 (N_6187,N_5817,N_5529);
nor U6188 (N_6188,N_5656,N_5421);
nor U6189 (N_6189,N_5735,N_5698);
nor U6190 (N_6190,N_5611,N_5636);
nand U6191 (N_6191,N_5580,N_5741);
or U6192 (N_6192,N_5715,N_5845);
nor U6193 (N_6193,N_5962,N_5728);
and U6194 (N_6194,N_5564,N_5594);
and U6195 (N_6195,N_5400,N_5690);
or U6196 (N_6196,N_5685,N_5747);
nor U6197 (N_6197,N_5994,N_5620);
xor U6198 (N_6198,N_5471,N_5664);
or U6199 (N_6199,N_5983,N_5631);
or U6200 (N_6200,N_5924,N_5504);
nand U6201 (N_6201,N_5786,N_5812);
or U6202 (N_6202,N_5834,N_5856);
or U6203 (N_6203,N_5952,N_5864);
and U6204 (N_6204,N_5895,N_5473);
or U6205 (N_6205,N_5480,N_5563);
nand U6206 (N_6206,N_5910,N_5562);
nor U6207 (N_6207,N_5484,N_5591);
nand U6208 (N_6208,N_5495,N_5808);
or U6209 (N_6209,N_5655,N_5596);
nand U6210 (N_6210,N_5602,N_5749);
and U6211 (N_6211,N_5538,N_5565);
nor U6212 (N_6212,N_5996,N_5530);
or U6213 (N_6213,N_5767,N_5532);
nor U6214 (N_6214,N_5977,N_5934);
nor U6215 (N_6215,N_5524,N_5907);
xnor U6216 (N_6216,N_5796,N_5578);
and U6217 (N_6217,N_5894,N_5651);
or U6218 (N_6218,N_5450,N_5885);
nor U6219 (N_6219,N_5837,N_5550);
nand U6220 (N_6220,N_5971,N_5673);
nor U6221 (N_6221,N_5609,N_5491);
nand U6222 (N_6222,N_5709,N_5884);
nand U6223 (N_6223,N_5858,N_5987);
xnor U6224 (N_6224,N_5826,N_5470);
and U6225 (N_6225,N_5801,N_5548);
xnor U6226 (N_6226,N_5595,N_5794);
xor U6227 (N_6227,N_5417,N_5922);
xnor U6228 (N_6228,N_5721,N_5822);
nand U6229 (N_6229,N_5714,N_5763);
nor U6230 (N_6230,N_5522,N_5505);
xnor U6231 (N_6231,N_5804,N_5439);
xnor U6232 (N_6232,N_5588,N_5455);
xnor U6233 (N_6233,N_5624,N_5738);
xnor U6234 (N_6234,N_5481,N_5919);
nand U6235 (N_6235,N_5652,N_5654);
and U6236 (N_6236,N_5986,N_5830);
or U6237 (N_6237,N_5696,N_5790);
nand U6238 (N_6238,N_5743,N_5560);
nand U6239 (N_6239,N_5493,N_5724);
and U6240 (N_6240,N_5615,N_5936);
nor U6241 (N_6241,N_5821,N_5752);
nor U6242 (N_6242,N_5433,N_5810);
nand U6243 (N_6243,N_5418,N_5537);
and U6244 (N_6244,N_5613,N_5868);
and U6245 (N_6245,N_5519,N_5997);
nand U6246 (N_6246,N_5630,N_5857);
and U6247 (N_6247,N_5880,N_5945);
and U6248 (N_6248,N_5461,N_5632);
nor U6249 (N_6249,N_5918,N_5740);
and U6250 (N_6250,N_5416,N_5488);
nand U6251 (N_6251,N_5755,N_5978);
nand U6252 (N_6252,N_5912,N_5554);
nor U6253 (N_6253,N_5889,N_5860);
xor U6254 (N_6254,N_5951,N_5621);
and U6255 (N_6255,N_5546,N_5937);
or U6256 (N_6256,N_5514,N_5904);
or U6257 (N_6257,N_5559,N_5604);
nor U6258 (N_6258,N_5795,N_5818);
nor U6259 (N_6259,N_5926,N_5467);
xnor U6260 (N_6260,N_5458,N_5540);
and U6261 (N_6261,N_5750,N_5887);
xnor U6262 (N_6262,N_5633,N_5598);
nand U6263 (N_6263,N_5659,N_5859);
xnor U6264 (N_6264,N_5497,N_5475);
and U6265 (N_6265,N_5712,N_5487);
and U6266 (N_6266,N_5511,N_5849);
xor U6267 (N_6267,N_5684,N_5508);
nand U6268 (N_6268,N_5993,N_5489);
and U6269 (N_6269,N_5939,N_5888);
nand U6270 (N_6270,N_5520,N_5572);
nand U6271 (N_6271,N_5852,N_5870);
or U6272 (N_6272,N_5973,N_5680);
or U6273 (N_6273,N_5886,N_5723);
and U6274 (N_6274,N_5404,N_5492);
nand U6275 (N_6275,N_5833,N_5628);
xor U6276 (N_6276,N_5955,N_5751);
nand U6277 (N_6277,N_5687,N_5423);
nand U6278 (N_6278,N_5729,N_5675);
and U6279 (N_6279,N_5865,N_5669);
and U6280 (N_6280,N_5544,N_5686);
nor U6281 (N_6281,N_5413,N_5597);
nor U6282 (N_6282,N_5782,N_5637);
nand U6283 (N_6283,N_5890,N_5403);
or U6284 (N_6284,N_5640,N_5806);
or U6285 (N_6285,N_5525,N_5625);
and U6286 (N_6286,N_5967,N_5468);
and U6287 (N_6287,N_5988,N_5876);
xor U6288 (N_6288,N_5957,N_5881);
or U6289 (N_6289,N_5407,N_5643);
and U6290 (N_6290,N_5502,N_5463);
xnor U6291 (N_6291,N_5929,N_5799);
or U6292 (N_6292,N_5875,N_5692);
nor U6293 (N_6293,N_5713,N_5768);
and U6294 (N_6294,N_5474,N_5412);
xor U6295 (N_6295,N_5639,N_5789);
xor U6296 (N_6296,N_5683,N_5940);
and U6297 (N_6297,N_5558,N_5820);
or U6298 (N_6298,N_5622,N_5674);
or U6299 (N_6299,N_5827,N_5662);
xor U6300 (N_6300,N_5481,N_5982);
nor U6301 (N_6301,N_5748,N_5780);
xor U6302 (N_6302,N_5967,N_5991);
xnor U6303 (N_6303,N_5958,N_5814);
and U6304 (N_6304,N_5869,N_5592);
and U6305 (N_6305,N_5908,N_5697);
nor U6306 (N_6306,N_5678,N_5947);
nand U6307 (N_6307,N_5551,N_5535);
nor U6308 (N_6308,N_5431,N_5718);
and U6309 (N_6309,N_5779,N_5776);
and U6310 (N_6310,N_5833,N_5776);
nand U6311 (N_6311,N_5880,N_5599);
and U6312 (N_6312,N_5873,N_5474);
xnor U6313 (N_6313,N_5426,N_5519);
nor U6314 (N_6314,N_5922,N_5892);
xnor U6315 (N_6315,N_5547,N_5622);
and U6316 (N_6316,N_5638,N_5714);
or U6317 (N_6317,N_5915,N_5522);
or U6318 (N_6318,N_5467,N_5403);
nand U6319 (N_6319,N_5804,N_5878);
or U6320 (N_6320,N_5898,N_5681);
and U6321 (N_6321,N_5539,N_5571);
nor U6322 (N_6322,N_5718,N_5956);
nand U6323 (N_6323,N_5819,N_5851);
nand U6324 (N_6324,N_5446,N_5798);
nor U6325 (N_6325,N_5779,N_5912);
and U6326 (N_6326,N_5875,N_5959);
nor U6327 (N_6327,N_5893,N_5792);
nand U6328 (N_6328,N_5857,N_5686);
or U6329 (N_6329,N_5735,N_5465);
nand U6330 (N_6330,N_5554,N_5790);
or U6331 (N_6331,N_5477,N_5424);
and U6332 (N_6332,N_5538,N_5638);
xor U6333 (N_6333,N_5416,N_5879);
nand U6334 (N_6334,N_5891,N_5415);
nand U6335 (N_6335,N_5463,N_5687);
or U6336 (N_6336,N_5443,N_5560);
xnor U6337 (N_6337,N_5470,N_5606);
or U6338 (N_6338,N_5616,N_5547);
nand U6339 (N_6339,N_5410,N_5598);
or U6340 (N_6340,N_5953,N_5903);
nand U6341 (N_6341,N_5631,N_5766);
or U6342 (N_6342,N_5626,N_5443);
xnor U6343 (N_6343,N_5714,N_5912);
nand U6344 (N_6344,N_5598,N_5779);
and U6345 (N_6345,N_5879,N_5652);
nand U6346 (N_6346,N_5424,N_5583);
and U6347 (N_6347,N_5527,N_5565);
or U6348 (N_6348,N_5547,N_5868);
or U6349 (N_6349,N_5802,N_5416);
and U6350 (N_6350,N_5445,N_5933);
xor U6351 (N_6351,N_5762,N_5432);
and U6352 (N_6352,N_5630,N_5795);
or U6353 (N_6353,N_5594,N_5770);
and U6354 (N_6354,N_5804,N_5747);
and U6355 (N_6355,N_5834,N_5741);
or U6356 (N_6356,N_5855,N_5599);
and U6357 (N_6357,N_5873,N_5497);
and U6358 (N_6358,N_5547,N_5527);
or U6359 (N_6359,N_5587,N_5929);
or U6360 (N_6360,N_5720,N_5530);
nor U6361 (N_6361,N_5648,N_5518);
and U6362 (N_6362,N_5961,N_5810);
or U6363 (N_6363,N_5782,N_5527);
xor U6364 (N_6364,N_5851,N_5572);
nand U6365 (N_6365,N_5798,N_5764);
xor U6366 (N_6366,N_5463,N_5944);
and U6367 (N_6367,N_5442,N_5877);
nor U6368 (N_6368,N_5572,N_5853);
nor U6369 (N_6369,N_5882,N_5641);
nand U6370 (N_6370,N_5763,N_5406);
xnor U6371 (N_6371,N_5501,N_5836);
nand U6372 (N_6372,N_5602,N_5668);
xnor U6373 (N_6373,N_5714,N_5471);
nor U6374 (N_6374,N_5433,N_5918);
and U6375 (N_6375,N_5518,N_5530);
nand U6376 (N_6376,N_5784,N_5407);
and U6377 (N_6377,N_5480,N_5897);
nor U6378 (N_6378,N_5793,N_5876);
nand U6379 (N_6379,N_5823,N_5731);
xor U6380 (N_6380,N_5657,N_5686);
nor U6381 (N_6381,N_5827,N_5520);
or U6382 (N_6382,N_5974,N_5455);
xor U6383 (N_6383,N_5858,N_5438);
or U6384 (N_6384,N_5843,N_5798);
nand U6385 (N_6385,N_5743,N_5716);
and U6386 (N_6386,N_5717,N_5687);
and U6387 (N_6387,N_5443,N_5773);
nor U6388 (N_6388,N_5927,N_5740);
nand U6389 (N_6389,N_5836,N_5854);
nand U6390 (N_6390,N_5759,N_5580);
or U6391 (N_6391,N_5608,N_5640);
nand U6392 (N_6392,N_5912,N_5627);
and U6393 (N_6393,N_5954,N_5547);
nor U6394 (N_6394,N_5428,N_5969);
xnor U6395 (N_6395,N_5774,N_5898);
or U6396 (N_6396,N_5428,N_5497);
and U6397 (N_6397,N_5857,N_5956);
nor U6398 (N_6398,N_5626,N_5589);
nor U6399 (N_6399,N_5946,N_5818);
or U6400 (N_6400,N_5455,N_5564);
nor U6401 (N_6401,N_5699,N_5400);
nand U6402 (N_6402,N_5776,N_5591);
and U6403 (N_6403,N_5762,N_5732);
or U6404 (N_6404,N_5517,N_5972);
xnor U6405 (N_6405,N_5708,N_5451);
and U6406 (N_6406,N_5464,N_5704);
xnor U6407 (N_6407,N_5642,N_5798);
and U6408 (N_6408,N_5491,N_5580);
xor U6409 (N_6409,N_5895,N_5497);
and U6410 (N_6410,N_5496,N_5573);
nor U6411 (N_6411,N_5674,N_5588);
nor U6412 (N_6412,N_5994,N_5818);
and U6413 (N_6413,N_5619,N_5977);
and U6414 (N_6414,N_5472,N_5506);
nand U6415 (N_6415,N_5510,N_5592);
nand U6416 (N_6416,N_5835,N_5938);
or U6417 (N_6417,N_5855,N_5814);
xor U6418 (N_6418,N_5815,N_5807);
nor U6419 (N_6419,N_5882,N_5668);
nand U6420 (N_6420,N_5998,N_5601);
nand U6421 (N_6421,N_5577,N_5472);
xnor U6422 (N_6422,N_5906,N_5801);
or U6423 (N_6423,N_5500,N_5910);
xor U6424 (N_6424,N_5706,N_5676);
nand U6425 (N_6425,N_5443,N_5609);
xnor U6426 (N_6426,N_5802,N_5959);
nand U6427 (N_6427,N_5645,N_5818);
nor U6428 (N_6428,N_5797,N_5724);
xor U6429 (N_6429,N_5411,N_5848);
nand U6430 (N_6430,N_5590,N_5941);
nor U6431 (N_6431,N_5417,N_5664);
xnor U6432 (N_6432,N_5841,N_5664);
xnor U6433 (N_6433,N_5941,N_5886);
and U6434 (N_6434,N_5998,N_5615);
nor U6435 (N_6435,N_5690,N_5647);
xnor U6436 (N_6436,N_5517,N_5629);
nor U6437 (N_6437,N_5542,N_5778);
or U6438 (N_6438,N_5605,N_5552);
nor U6439 (N_6439,N_5515,N_5458);
nor U6440 (N_6440,N_5517,N_5665);
xor U6441 (N_6441,N_5456,N_5479);
nor U6442 (N_6442,N_5757,N_5515);
and U6443 (N_6443,N_5583,N_5754);
xor U6444 (N_6444,N_5429,N_5493);
xnor U6445 (N_6445,N_5456,N_5656);
or U6446 (N_6446,N_5521,N_5876);
or U6447 (N_6447,N_5925,N_5558);
and U6448 (N_6448,N_5897,N_5994);
and U6449 (N_6449,N_5902,N_5619);
and U6450 (N_6450,N_5845,N_5535);
nor U6451 (N_6451,N_5794,N_5409);
and U6452 (N_6452,N_5671,N_5508);
nand U6453 (N_6453,N_5630,N_5647);
nand U6454 (N_6454,N_5836,N_5929);
and U6455 (N_6455,N_5462,N_5512);
nor U6456 (N_6456,N_5958,N_5911);
xor U6457 (N_6457,N_5905,N_5801);
nand U6458 (N_6458,N_5482,N_5567);
nor U6459 (N_6459,N_5841,N_5423);
and U6460 (N_6460,N_5733,N_5651);
nand U6461 (N_6461,N_5566,N_5432);
xnor U6462 (N_6462,N_5483,N_5664);
xor U6463 (N_6463,N_5840,N_5900);
and U6464 (N_6464,N_5792,N_5567);
or U6465 (N_6465,N_5595,N_5464);
xor U6466 (N_6466,N_5439,N_5673);
nor U6467 (N_6467,N_5611,N_5826);
nor U6468 (N_6468,N_5409,N_5402);
or U6469 (N_6469,N_5947,N_5535);
and U6470 (N_6470,N_5773,N_5940);
xor U6471 (N_6471,N_5731,N_5698);
nand U6472 (N_6472,N_5850,N_5836);
or U6473 (N_6473,N_5775,N_5989);
nor U6474 (N_6474,N_5574,N_5664);
and U6475 (N_6475,N_5588,N_5505);
xor U6476 (N_6476,N_5810,N_5544);
and U6477 (N_6477,N_5590,N_5655);
and U6478 (N_6478,N_5917,N_5880);
xor U6479 (N_6479,N_5900,N_5556);
nand U6480 (N_6480,N_5580,N_5902);
and U6481 (N_6481,N_5844,N_5530);
nor U6482 (N_6482,N_5416,N_5790);
nand U6483 (N_6483,N_5766,N_5565);
xor U6484 (N_6484,N_5419,N_5911);
and U6485 (N_6485,N_5535,N_5403);
or U6486 (N_6486,N_5479,N_5972);
or U6487 (N_6487,N_5803,N_5526);
nand U6488 (N_6488,N_5575,N_5791);
or U6489 (N_6489,N_5825,N_5831);
and U6490 (N_6490,N_5427,N_5654);
nand U6491 (N_6491,N_5979,N_5447);
nor U6492 (N_6492,N_5739,N_5811);
nor U6493 (N_6493,N_5935,N_5468);
nand U6494 (N_6494,N_5873,N_5629);
or U6495 (N_6495,N_5662,N_5900);
xnor U6496 (N_6496,N_5583,N_5759);
and U6497 (N_6497,N_5729,N_5657);
xor U6498 (N_6498,N_5407,N_5752);
or U6499 (N_6499,N_5844,N_5408);
nor U6500 (N_6500,N_5974,N_5654);
nand U6501 (N_6501,N_5931,N_5925);
xnor U6502 (N_6502,N_5707,N_5955);
nor U6503 (N_6503,N_5760,N_5890);
and U6504 (N_6504,N_5711,N_5639);
nor U6505 (N_6505,N_5680,N_5610);
nand U6506 (N_6506,N_5433,N_5655);
or U6507 (N_6507,N_5931,N_5720);
xnor U6508 (N_6508,N_5867,N_5526);
and U6509 (N_6509,N_5811,N_5567);
or U6510 (N_6510,N_5774,N_5454);
and U6511 (N_6511,N_5645,N_5768);
nor U6512 (N_6512,N_5994,N_5522);
xnor U6513 (N_6513,N_5464,N_5669);
and U6514 (N_6514,N_5976,N_5889);
xnor U6515 (N_6515,N_5457,N_5931);
nand U6516 (N_6516,N_5506,N_5584);
or U6517 (N_6517,N_5779,N_5619);
nor U6518 (N_6518,N_5736,N_5652);
xor U6519 (N_6519,N_5621,N_5833);
and U6520 (N_6520,N_5626,N_5799);
nand U6521 (N_6521,N_5851,N_5508);
and U6522 (N_6522,N_5705,N_5483);
xor U6523 (N_6523,N_5957,N_5578);
and U6524 (N_6524,N_5509,N_5691);
nand U6525 (N_6525,N_5551,N_5741);
nand U6526 (N_6526,N_5903,N_5521);
or U6527 (N_6527,N_5503,N_5561);
xor U6528 (N_6528,N_5891,N_5955);
and U6529 (N_6529,N_5729,N_5682);
nand U6530 (N_6530,N_5415,N_5546);
xnor U6531 (N_6531,N_5637,N_5555);
xnor U6532 (N_6532,N_5427,N_5530);
nor U6533 (N_6533,N_5491,N_5538);
xor U6534 (N_6534,N_5996,N_5687);
nand U6535 (N_6535,N_5600,N_5584);
nand U6536 (N_6536,N_5750,N_5999);
xor U6537 (N_6537,N_5776,N_5482);
and U6538 (N_6538,N_5738,N_5797);
or U6539 (N_6539,N_5725,N_5467);
and U6540 (N_6540,N_5755,N_5525);
and U6541 (N_6541,N_5863,N_5668);
xnor U6542 (N_6542,N_5978,N_5941);
or U6543 (N_6543,N_5899,N_5998);
xnor U6544 (N_6544,N_5400,N_5852);
nor U6545 (N_6545,N_5810,N_5785);
or U6546 (N_6546,N_5624,N_5765);
or U6547 (N_6547,N_5462,N_5977);
and U6548 (N_6548,N_5781,N_5496);
nor U6549 (N_6549,N_5484,N_5683);
and U6550 (N_6550,N_5980,N_5882);
nand U6551 (N_6551,N_5691,N_5920);
and U6552 (N_6552,N_5962,N_5851);
and U6553 (N_6553,N_5538,N_5478);
nand U6554 (N_6554,N_5404,N_5810);
nor U6555 (N_6555,N_5653,N_5869);
or U6556 (N_6556,N_5932,N_5804);
and U6557 (N_6557,N_5876,N_5801);
nor U6558 (N_6558,N_5596,N_5690);
and U6559 (N_6559,N_5983,N_5678);
nor U6560 (N_6560,N_5733,N_5996);
and U6561 (N_6561,N_5947,N_5483);
and U6562 (N_6562,N_5558,N_5692);
nand U6563 (N_6563,N_5761,N_5607);
nor U6564 (N_6564,N_5474,N_5794);
xnor U6565 (N_6565,N_5955,N_5567);
and U6566 (N_6566,N_5595,N_5591);
nor U6567 (N_6567,N_5563,N_5829);
xor U6568 (N_6568,N_5549,N_5466);
and U6569 (N_6569,N_5727,N_5991);
and U6570 (N_6570,N_5495,N_5650);
xnor U6571 (N_6571,N_5924,N_5904);
nand U6572 (N_6572,N_5627,N_5796);
nor U6573 (N_6573,N_5726,N_5723);
xor U6574 (N_6574,N_5636,N_5916);
or U6575 (N_6575,N_5848,N_5556);
and U6576 (N_6576,N_5829,N_5610);
or U6577 (N_6577,N_5436,N_5543);
and U6578 (N_6578,N_5846,N_5792);
nor U6579 (N_6579,N_5680,N_5822);
or U6580 (N_6580,N_5795,N_5455);
and U6581 (N_6581,N_5615,N_5851);
or U6582 (N_6582,N_5881,N_5417);
nor U6583 (N_6583,N_5781,N_5443);
xnor U6584 (N_6584,N_5759,N_5958);
and U6585 (N_6585,N_5759,N_5704);
xnor U6586 (N_6586,N_5637,N_5648);
nor U6587 (N_6587,N_5782,N_5950);
xor U6588 (N_6588,N_5927,N_5782);
or U6589 (N_6589,N_5609,N_5894);
and U6590 (N_6590,N_5406,N_5610);
xor U6591 (N_6591,N_5844,N_5586);
xor U6592 (N_6592,N_5445,N_5936);
nand U6593 (N_6593,N_5945,N_5807);
or U6594 (N_6594,N_5729,N_5627);
xnor U6595 (N_6595,N_5955,N_5614);
xnor U6596 (N_6596,N_5678,N_5545);
and U6597 (N_6597,N_5797,N_5403);
or U6598 (N_6598,N_5402,N_5709);
nand U6599 (N_6599,N_5488,N_5858);
or U6600 (N_6600,N_6221,N_6505);
nor U6601 (N_6601,N_6029,N_6477);
xor U6602 (N_6602,N_6511,N_6503);
xor U6603 (N_6603,N_6025,N_6297);
xnor U6604 (N_6604,N_6369,N_6561);
nand U6605 (N_6605,N_6204,N_6462);
and U6606 (N_6606,N_6243,N_6069);
nand U6607 (N_6607,N_6480,N_6510);
nand U6608 (N_6608,N_6016,N_6395);
or U6609 (N_6609,N_6015,N_6392);
and U6610 (N_6610,N_6402,N_6096);
and U6611 (N_6611,N_6496,N_6393);
xor U6612 (N_6612,N_6102,N_6523);
nor U6613 (N_6613,N_6301,N_6125);
xor U6614 (N_6614,N_6324,N_6407);
nor U6615 (N_6615,N_6061,N_6411);
xor U6616 (N_6616,N_6321,N_6295);
nand U6617 (N_6617,N_6450,N_6579);
nand U6618 (N_6618,N_6388,N_6544);
or U6619 (N_6619,N_6173,N_6192);
or U6620 (N_6620,N_6240,N_6304);
or U6621 (N_6621,N_6362,N_6430);
nor U6622 (N_6622,N_6489,N_6217);
nand U6623 (N_6623,N_6536,N_6030);
or U6624 (N_6624,N_6282,N_6339);
or U6625 (N_6625,N_6097,N_6002);
nand U6626 (N_6626,N_6250,N_6119);
nor U6627 (N_6627,N_6058,N_6584);
xor U6628 (N_6628,N_6279,N_6149);
and U6629 (N_6629,N_6524,N_6409);
and U6630 (N_6630,N_6436,N_6062);
nor U6631 (N_6631,N_6384,N_6386);
nor U6632 (N_6632,N_6468,N_6396);
and U6633 (N_6633,N_6162,N_6031);
xnor U6634 (N_6634,N_6049,N_6131);
or U6635 (N_6635,N_6228,N_6539);
or U6636 (N_6636,N_6146,N_6249);
and U6637 (N_6637,N_6086,N_6059);
and U6638 (N_6638,N_6020,N_6398);
nand U6639 (N_6639,N_6267,N_6599);
nor U6640 (N_6640,N_6458,N_6389);
xnor U6641 (N_6641,N_6134,N_6274);
nor U6642 (N_6642,N_6521,N_6072);
or U6643 (N_6643,N_6296,N_6068);
and U6644 (N_6644,N_6590,N_6547);
or U6645 (N_6645,N_6591,N_6229);
nor U6646 (N_6646,N_6050,N_6514);
or U6647 (N_6647,N_6311,N_6567);
xor U6648 (N_6648,N_6543,N_6472);
nand U6649 (N_6649,N_6042,N_6105);
nor U6650 (N_6650,N_6180,N_6326);
or U6651 (N_6651,N_6248,N_6285);
and U6652 (N_6652,N_6275,N_6508);
xor U6653 (N_6653,N_6222,N_6185);
nor U6654 (N_6654,N_6017,N_6094);
nand U6655 (N_6655,N_6383,N_6583);
nand U6656 (N_6656,N_6338,N_6004);
nor U6657 (N_6657,N_6492,N_6365);
xnor U6658 (N_6658,N_6137,N_6236);
xnor U6659 (N_6659,N_6112,N_6494);
nand U6660 (N_6660,N_6394,N_6196);
nor U6661 (N_6661,N_6466,N_6423);
nor U6662 (N_6662,N_6055,N_6447);
and U6663 (N_6663,N_6574,N_6063);
nor U6664 (N_6664,N_6560,N_6382);
nor U6665 (N_6665,N_6313,N_6417);
and U6666 (N_6666,N_6551,N_6310);
nand U6667 (N_6667,N_6372,N_6242);
or U6668 (N_6668,N_6107,N_6155);
or U6669 (N_6669,N_6272,N_6467);
or U6670 (N_6670,N_6405,N_6485);
nor U6671 (N_6671,N_6512,N_6057);
and U6672 (N_6672,N_6438,N_6408);
xnor U6673 (N_6673,N_6360,N_6404);
or U6674 (N_6674,N_6251,N_6182);
xnor U6675 (N_6675,N_6459,N_6165);
or U6676 (N_6676,N_6344,N_6197);
nor U6677 (N_6677,N_6569,N_6451);
and U6678 (N_6678,N_6400,N_6479);
nand U6679 (N_6679,N_6376,N_6186);
nor U6680 (N_6680,N_6470,N_6270);
xnor U6681 (N_6681,N_6586,N_6227);
nand U6682 (N_6682,N_6148,N_6070);
nor U6683 (N_6683,N_6435,N_6246);
xnor U6684 (N_6684,N_6527,N_6201);
nand U6685 (N_6685,N_6481,N_6047);
xor U6686 (N_6686,N_6212,N_6244);
nor U6687 (N_6687,N_6158,N_6128);
nand U6688 (N_6688,N_6261,N_6441);
xnor U6689 (N_6689,N_6150,N_6566);
xnor U6690 (N_6690,N_6126,N_6044);
xnor U6691 (N_6691,N_6167,N_6427);
nand U6692 (N_6692,N_6585,N_6516);
and U6693 (N_6693,N_6298,N_6009);
nor U6694 (N_6694,N_6314,N_6170);
or U6695 (N_6695,N_6499,N_6143);
xor U6696 (N_6696,N_6060,N_6537);
or U6697 (N_6697,N_6135,N_6533);
or U6698 (N_6698,N_6006,N_6136);
or U6699 (N_6699,N_6113,N_6426);
and U6700 (N_6700,N_6247,N_6198);
nor U6701 (N_6701,N_6399,N_6034);
xor U6702 (N_6702,N_6043,N_6218);
nor U6703 (N_6703,N_6147,N_6273);
and U6704 (N_6704,N_6159,N_6419);
nor U6705 (N_6705,N_6152,N_6488);
or U6706 (N_6706,N_6259,N_6406);
xor U6707 (N_6707,N_6140,N_6570);
or U6708 (N_6708,N_6163,N_6000);
or U6709 (N_6709,N_6429,N_6093);
xor U6710 (N_6710,N_6234,N_6100);
nor U6711 (N_6711,N_6346,N_6291);
or U6712 (N_6712,N_6495,N_6177);
nor U6713 (N_6713,N_6422,N_6587);
and U6714 (N_6714,N_6012,N_6509);
xor U6715 (N_6715,N_6067,N_6497);
xor U6716 (N_6716,N_6431,N_6139);
and U6717 (N_6717,N_6108,N_6293);
nor U6718 (N_6718,N_6255,N_6315);
nand U6719 (N_6719,N_6506,N_6142);
xnor U6720 (N_6720,N_6048,N_6144);
or U6721 (N_6721,N_6230,N_6118);
and U6722 (N_6722,N_6164,N_6073);
and U6723 (N_6723,N_6453,N_6367);
and U6724 (N_6724,N_6014,N_6556);
and U6725 (N_6725,N_6379,N_6548);
xnor U6726 (N_6726,N_6403,N_6518);
nand U6727 (N_6727,N_6424,N_6082);
xor U6728 (N_6728,N_6446,N_6265);
nor U6729 (N_6729,N_6575,N_6233);
nand U6730 (N_6730,N_6032,N_6323);
or U6731 (N_6731,N_6036,N_6329);
xnor U6732 (N_6732,N_6300,N_6239);
xor U6733 (N_6733,N_6565,N_6127);
nand U6734 (N_6734,N_6562,N_6117);
nor U6735 (N_6735,N_6361,N_6445);
xor U6736 (N_6736,N_6018,N_6373);
and U6737 (N_6737,N_6380,N_6111);
nand U6738 (N_6738,N_6178,N_6151);
or U6739 (N_6739,N_6349,N_6114);
and U6740 (N_6740,N_6377,N_6487);
nor U6741 (N_6741,N_6331,N_6303);
xor U6742 (N_6742,N_6317,N_6374);
xnor U6743 (N_6743,N_6200,N_6237);
xnor U6744 (N_6744,N_6166,N_6532);
nand U6745 (N_6745,N_6215,N_6104);
or U6746 (N_6746,N_6318,N_6541);
or U6747 (N_6747,N_6175,N_6368);
nand U6748 (N_6748,N_6254,N_6580);
nand U6749 (N_6749,N_6076,N_6263);
or U6750 (N_6750,N_6581,N_6482);
or U6751 (N_6751,N_6530,N_6428);
and U6752 (N_6752,N_6592,N_6594);
and U6753 (N_6753,N_6121,N_6235);
nor U6754 (N_6754,N_6037,N_6397);
and U6755 (N_6755,N_6335,N_6209);
nand U6756 (N_6756,N_6437,N_6474);
and U6757 (N_6757,N_6354,N_6553);
and U6758 (N_6758,N_6064,N_6224);
nor U6759 (N_6759,N_6262,N_6308);
and U6760 (N_6760,N_6110,N_6053);
xnor U6761 (N_6761,N_6101,N_6046);
nor U6762 (N_6762,N_6486,N_6231);
or U6763 (N_6763,N_6122,N_6171);
and U6764 (N_6764,N_6091,N_6271);
and U6765 (N_6765,N_6109,N_6007);
and U6766 (N_6766,N_6381,N_6309);
or U6767 (N_6767,N_6001,N_6095);
or U6768 (N_6768,N_6203,N_6054);
or U6769 (N_6769,N_6473,N_6056);
nand U6770 (N_6770,N_6005,N_6457);
nand U6771 (N_6771,N_6515,N_6455);
or U6772 (N_6772,N_6202,N_6195);
and U6773 (N_6773,N_6507,N_6520);
and U6774 (N_6774,N_6019,N_6522);
and U6775 (N_6775,N_6129,N_6535);
or U6776 (N_6776,N_6232,N_6568);
nand U6777 (N_6777,N_6563,N_6375);
or U6778 (N_6778,N_6041,N_6026);
or U6779 (N_6779,N_6206,N_6199);
or U6780 (N_6780,N_6442,N_6552);
nand U6781 (N_6781,N_6087,N_6258);
and U6782 (N_6782,N_6154,N_6410);
xor U6783 (N_6783,N_6421,N_6003);
nor U6784 (N_6784,N_6452,N_6328);
nor U6785 (N_6785,N_6189,N_6208);
or U6786 (N_6786,N_6174,N_6475);
xnor U6787 (N_6787,N_6546,N_6184);
or U6788 (N_6788,N_6210,N_6440);
or U6789 (N_6789,N_6130,N_6513);
nor U6790 (N_6790,N_6425,N_6207);
nor U6791 (N_6791,N_6359,N_6120);
nor U6792 (N_6792,N_6370,N_6035);
nor U6793 (N_6793,N_6010,N_6434);
xor U6794 (N_6794,N_6106,N_6416);
and U6795 (N_6795,N_6266,N_6588);
and U6796 (N_6796,N_6168,N_6460);
and U6797 (N_6797,N_6078,N_6132);
nand U6798 (N_6798,N_6577,N_6350);
nand U6799 (N_6799,N_6269,N_6099);
xor U6800 (N_6800,N_6220,N_6502);
nand U6801 (N_6801,N_6252,N_6219);
nor U6802 (N_6802,N_6433,N_6194);
and U6803 (N_6803,N_6519,N_6052);
and U6804 (N_6804,N_6549,N_6176);
or U6805 (N_6805,N_6325,N_6124);
nor U6806 (N_6806,N_6385,N_6593);
xor U6807 (N_6807,N_6312,N_6337);
xnor U6808 (N_6808,N_6491,N_6504);
nand U6809 (N_6809,N_6021,N_6500);
or U6810 (N_6810,N_6033,N_6075);
xor U6811 (N_6811,N_6531,N_6306);
xor U6812 (N_6812,N_6088,N_6299);
or U6813 (N_6813,N_6038,N_6596);
or U6814 (N_6814,N_6305,N_6065);
nor U6815 (N_6815,N_6336,N_6083);
or U6816 (N_6816,N_6045,N_6432);
and U6817 (N_6817,N_6223,N_6534);
nor U6818 (N_6818,N_6316,N_6322);
or U6819 (N_6819,N_6456,N_6342);
nand U6820 (N_6820,N_6559,N_6187);
and U6821 (N_6821,N_6448,N_6387);
or U6822 (N_6822,N_6412,N_6077);
xor U6823 (N_6823,N_6557,N_6191);
xnor U6824 (N_6824,N_6153,N_6378);
nor U6825 (N_6825,N_6169,N_6027);
nor U6826 (N_6826,N_6355,N_6141);
xnor U6827 (N_6827,N_6550,N_6283);
or U6828 (N_6828,N_6517,N_6225);
nor U6829 (N_6829,N_6528,N_6356);
nand U6830 (N_6830,N_6414,N_6011);
xnor U6831 (N_6831,N_6286,N_6598);
or U6832 (N_6832,N_6444,N_6501);
xor U6833 (N_6833,N_6090,N_6066);
or U6834 (N_6834,N_6276,N_6555);
nand U6835 (N_6835,N_6260,N_6319);
xnor U6836 (N_6836,N_6022,N_6092);
and U6837 (N_6837,N_6353,N_6526);
xnor U6838 (N_6838,N_6347,N_6554);
xor U6839 (N_6839,N_6116,N_6449);
nor U6840 (N_6840,N_6573,N_6363);
or U6841 (N_6841,N_6211,N_6478);
nand U6842 (N_6842,N_6542,N_6080);
or U6843 (N_6843,N_6277,N_6443);
xor U6844 (N_6844,N_6582,N_6074);
xor U6845 (N_6845,N_6348,N_6454);
xor U6846 (N_6846,N_6264,N_6278);
nor U6847 (N_6847,N_6545,N_6418);
and U6848 (N_6848,N_6213,N_6039);
or U6849 (N_6849,N_6190,N_6498);
and U6850 (N_6850,N_6558,N_6351);
nor U6851 (N_6851,N_6028,N_6538);
or U6852 (N_6852,N_6288,N_6597);
or U6853 (N_6853,N_6420,N_6307);
nor U6854 (N_6854,N_6290,N_6332);
and U6855 (N_6855,N_6085,N_6103);
and U6856 (N_6856,N_6160,N_6490);
or U6857 (N_6857,N_6156,N_6357);
nand U6858 (N_6858,N_6253,N_6115);
nor U6859 (N_6859,N_6008,N_6330);
and U6860 (N_6860,N_6302,N_6257);
or U6861 (N_6861,N_6364,N_6023);
nand U6862 (N_6862,N_6484,N_6133);
xor U6863 (N_6863,N_6327,N_6476);
nand U6864 (N_6864,N_6157,N_6071);
nand U6865 (N_6865,N_6013,N_6589);
or U6866 (N_6866,N_6292,N_6390);
nand U6867 (N_6867,N_6401,N_6098);
xor U6868 (N_6868,N_6179,N_6145);
nand U6869 (N_6869,N_6268,N_6352);
xnor U6870 (N_6870,N_6320,N_6289);
nor U6871 (N_6871,N_6483,N_6529);
nand U6872 (N_6872,N_6461,N_6464);
and U6873 (N_6873,N_6540,N_6341);
or U6874 (N_6874,N_6294,N_6334);
nand U6875 (N_6875,N_6366,N_6183);
nand U6876 (N_6876,N_6465,N_6238);
and U6877 (N_6877,N_6525,N_6205);
or U6878 (N_6878,N_6138,N_6415);
xor U6879 (N_6879,N_6172,N_6226);
and U6880 (N_6880,N_6343,N_6371);
xnor U6881 (N_6881,N_6333,N_6358);
xor U6882 (N_6882,N_6345,N_6051);
nand U6883 (N_6883,N_6193,N_6079);
or U6884 (N_6884,N_6571,N_6572);
and U6885 (N_6885,N_6391,N_6123);
and U6886 (N_6886,N_6284,N_6564);
nand U6887 (N_6887,N_6181,N_6576);
xor U6888 (N_6888,N_6280,N_6469);
xnor U6889 (N_6889,N_6024,N_6595);
nand U6890 (N_6890,N_6493,N_6471);
nand U6891 (N_6891,N_6578,N_6463);
nor U6892 (N_6892,N_6214,N_6245);
or U6893 (N_6893,N_6281,N_6084);
nor U6894 (N_6894,N_6340,N_6089);
and U6895 (N_6895,N_6241,N_6439);
or U6896 (N_6896,N_6161,N_6081);
and U6897 (N_6897,N_6256,N_6413);
xor U6898 (N_6898,N_6188,N_6040);
and U6899 (N_6899,N_6216,N_6287);
and U6900 (N_6900,N_6167,N_6361);
or U6901 (N_6901,N_6094,N_6315);
nand U6902 (N_6902,N_6285,N_6367);
xor U6903 (N_6903,N_6582,N_6052);
nand U6904 (N_6904,N_6001,N_6091);
and U6905 (N_6905,N_6306,N_6118);
nor U6906 (N_6906,N_6373,N_6141);
and U6907 (N_6907,N_6297,N_6490);
nor U6908 (N_6908,N_6466,N_6393);
nor U6909 (N_6909,N_6519,N_6006);
nor U6910 (N_6910,N_6300,N_6409);
nand U6911 (N_6911,N_6504,N_6541);
nand U6912 (N_6912,N_6581,N_6207);
nand U6913 (N_6913,N_6003,N_6511);
and U6914 (N_6914,N_6544,N_6237);
nor U6915 (N_6915,N_6469,N_6520);
xnor U6916 (N_6916,N_6308,N_6018);
xnor U6917 (N_6917,N_6333,N_6097);
and U6918 (N_6918,N_6374,N_6587);
nand U6919 (N_6919,N_6073,N_6288);
nand U6920 (N_6920,N_6203,N_6171);
nand U6921 (N_6921,N_6501,N_6200);
nor U6922 (N_6922,N_6238,N_6538);
or U6923 (N_6923,N_6014,N_6290);
or U6924 (N_6924,N_6389,N_6198);
nor U6925 (N_6925,N_6042,N_6033);
or U6926 (N_6926,N_6540,N_6391);
xnor U6927 (N_6927,N_6277,N_6444);
xnor U6928 (N_6928,N_6264,N_6488);
nand U6929 (N_6929,N_6002,N_6181);
and U6930 (N_6930,N_6156,N_6446);
nor U6931 (N_6931,N_6582,N_6517);
xnor U6932 (N_6932,N_6593,N_6511);
nand U6933 (N_6933,N_6375,N_6030);
and U6934 (N_6934,N_6571,N_6008);
or U6935 (N_6935,N_6243,N_6473);
nor U6936 (N_6936,N_6340,N_6490);
xor U6937 (N_6937,N_6312,N_6354);
or U6938 (N_6938,N_6325,N_6405);
nor U6939 (N_6939,N_6100,N_6105);
nor U6940 (N_6940,N_6343,N_6564);
nor U6941 (N_6941,N_6332,N_6524);
nand U6942 (N_6942,N_6323,N_6108);
xnor U6943 (N_6943,N_6284,N_6563);
nor U6944 (N_6944,N_6552,N_6309);
nor U6945 (N_6945,N_6410,N_6151);
nor U6946 (N_6946,N_6264,N_6474);
or U6947 (N_6947,N_6487,N_6425);
nand U6948 (N_6948,N_6403,N_6405);
nand U6949 (N_6949,N_6039,N_6464);
and U6950 (N_6950,N_6164,N_6309);
or U6951 (N_6951,N_6273,N_6158);
nand U6952 (N_6952,N_6163,N_6435);
or U6953 (N_6953,N_6512,N_6147);
and U6954 (N_6954,N_6218,N_6091);
or U6955 (N_6955,N_6436,N_6112);
xor U6956 (N_6956,N_6052,N_6589);
xor U6957 (N_6957,N_6434,N_6238);
nor U6958 (N_6958,N_6079,N_6051);
or U6959 (N_6959,N_6329,N_6233);
xnor U6960 (N_6960,N_6260,N_6272);
nor U6961 (N_6961,N_6506,N_6287);
xor U6962 (N_6962,N_6570,N_6300);
and U6963 (N_6963,N_6259,N_6525);
and U6964 (N_6964,N_6092,N_6374);
nand U6965 (N_6965,N_6575,N_6235);
and U6966 (N_6966,N_6200,N_6059);
xor U6967 (N_6967,N_6106,N_6571);
nor U6968 (N_6968,N_6069,N_6219);
or U6969 (N_6969,N_6518,N_6058);
and U6970 (N_6970,N_6568,N_6319);
nor U6971 (N_6971,N_6298,N_6024);
nor U6972 (N_6972,N_6453,N_6104);
nor U6973 (N_6973,N_6314,N_6301);
or U6974 (N_6974,N_6495,N_6283);
and U6975 (N_6975,N_6490,N_6386);
xor U6976 (N_6976,N_6122,N_6032);
or U6977 (N_6977,N_6528,N_6108);
or U6978 (N_6978,N_6541,N_6316);
or U6979 (N_6979,N_6310,N_6485);
nand U6980 (N_6980,N_6018,N_6412);
nand U6981 (N_6981,N_6243,N_6127);
nand U6982 (N_6982,N_6525,N_6359);
nor U6983 (N_6983,N_6449,N_6550);
nor U6984 (N_6984,N_6009,N_6247);
nand U6985 (N_6985,N_6498,N_6355);
nor U6986 (N_6986,N_6493,N_6473);
nor U6987 (N_6987,N_6214,N_6498);
nand U6988 (N_6988,N_6168,N_6314);
and U6989 (N_6989,N_6501,N_6198);
and U6990 (N_6990,N_6288,N_6400);
nand U6991 (N_6991,N_6270,N_6500);
xnor U6992 (N_6992,N_6373,N_6076);
or U6993 (N_6993,N_6551,N_6480);
nor U6994 (N_6994,N_6509,N_6008);
nor U6995 (N_6995,N_6373,N_6191);
or U6996 (N_6996,N_6113,N_6114);
or U6997 (N_6997,N_6483,N_6018);
and U6998 (N_6998,N_6364,N_6270);
and U6999 (N_6999,N_6526,N_6094);
or U7000 (N_7000,N_6414,N_6203);
xor U7001 (N_7001,N_6529,N_6123);
nor U7002 (N_7002,N_6501,N_6554);
xor U7003 (N_7003,N_6195,N_6487);
xnor U7004 (N_7004,N_6250,N_6352);
nor U7005 (N_7005,N_6202,N_6212);
and U7006 (N_7006,N_6149,N_6143);
or U7007 (N_7007,N_6474,N_6526);
xnor U7008 (N_7008,N_6478,N_6144);
nand U7009 (N_7009,N_6500,N_6192);
and U7010 (N_7010,N_6358,N_6464);
nor U7011 (N_7011,N_6228,N_6363);
nand U7012 (N_7012,N_6181,N_6036);
xnor U7013 (N_7013,N_6529,N_6044);
xnor U7014 (N_7014,N_6266,N_6120);
or U7015 (N_7015,N_6286,N_6297);
nand U7016 (N_7016,N_6042,N_6328);
xor U7017 (N_7017,N_6310,N_6254);
and U7018 (N_7018,N_6546,N_6306);
or U7019 (N_7019,N_6231,N_6493);
or U7020 (N_7020,N_6077,N_6386);
nand U7021 (N_7021,N_6174,N_6252);
and U7022 (N_7022,N_6511,N_6254);
xnor U7023 (N_7023,N_6336,N_6106);
and U7024 (N_7024,N_6154,N_6221);
and U7025 (N_7025,N_6299,N_6188);
nor U7026 (N_7026,N_6310,N_6394);
nand U7027 (N_7027,N_6244,N_6076);
xor U7028 (N_7028,N_6054,N_6526);
nor U7029 (N_7029,N_6395,N_6174);
and U7030 (N_7030,N_6332,N_6354);
nor U7031 (N_7031,N_6016,N_6401);
nand U7032 (N_7032,N_6125,N_6530);
and U7033 (N_7033,N_6297,N_6402);
or U7034 (N_7034,N_6494,N_6218);
or U7035 (N_7035,N_6392,N_6099);
and U7036 (N_7036,N_6468,N_6293);
nor U7037 (N_7037,N_6510,N_6088);
and U7038 (N_7038,N_6142,N_6194);
xnor U7039 (N_7039,N_6111,N_6292);
or U7040 (N_7040,N_6285,N_6340);
nor U7041 (N_7041,N_6323,N_6539);
or U7042 (N_7042,N_6208,N_6363);
and U7043 (N_7043,N_6239,N_6499);
xor U7044 (N_7044,N_6350,N_6541);
xor U7045 (N_7045,N_6191,N_6469);
or U7046 (N_7046,N_6380,N_6192);
nand U7047 (N_7047,N_6491,N_6353);
and U7048 (N_7048,N_6234,N_6270);
or U7049 (N_7049,N_6275,N_6188);
or U7050 (N_7050,N_6464,N_6192);
or U7051 (N_7051,N_6201,N_6212);
and U7052 (N_7052,N_6361,N_6075);
nor U7053 (N_7053,N_6379,N_6276);
nand U7054 (N_7054,N_6511,N_6349);
and U7055 (N_7055,N_6537,N_6055);
or U7056 (N_7056,N_6257,N_6283);
nor U7057 (N_7057,N_6291,N_6556);
nand U7058 (N_7058,N_6052,N_6551);
xor U7059 (N_7059,N_6204,N_6429);
or U7060 (N_7060,N_6205,N_6559);
nand U7061 (N_7061,N_6571,N_6324);
xor U7062 (N_7062,N_6317,N_6025);
nor U7063 (N_7063,N_6416,N_6041);
xnor U7064 (N_7064,N_6382,N_6595);
nor U7065 (N_7065,N_6389,N_6105);
or U7066 (N_7066,N_6432,N_6236);
xor U7067 (N_7067,N_6029,N_6580);
and U7068 (N_7068,N_6212,N_6283);
nor U7069 (N_7069,N_6382,N_6181);
xor U7070 (N_7070,N_6007,N_6335);
or U7071 (N_7071,N_6181,N_6111);
or U7072 (N_7072,N_6233,N_6191);
and U7073 (N_7073,N_6124,N_6281);
and U7074 (N_7074,N_6077,N_6267);
nor U7075 (N_7075,N_6025,N_6434);
xor U7076 (N_7076,N_6263,N_6335);
xnor U7077 (N_7077,N_6063,N_6319);
nor U7078 (N_7078,N_6075,N_6045);
xnor U7079 (N_7079,N_6391,N_6109);
nor U7080 (N_7080,N_6279,N_6269);
or U7081 (N_7081,N_6586,N_6201);
and U7082 (N_7082,N_6352,N_6019);
or U7083 (N_7083,N_6233,N_6512);
nand U7084 (N_7084,N_6410,N_6094);
nand U7085 (N_7085,N_6350,N_6351);
nor U7086 (N_7086,N_6221,N_6193);
and U7087 (N_7087,N_6047,N_6049);
nand U7088 (N_7088,N_6099,N_6138);
or U7089 (N_7089,N_6257,N_6565);
and U7090 (N_7090,N_6206,N_6123);
or U7091 (N_7091,N_6394,N_6534);
or U7092 (N_7092,N_6345,N_6075);
and U7093 (N_7093,N_6556,N_6463);
nand U7094 (N_7094,N_6445,N_6498);
xor U7095 (N_7095,N_6124,N_6145);
xor U7096 (N_7096,N_6487,N_6493);
or U7097 (N_7097,N_6008,N_6543);
or U7098 (N_7098,N_6316,N_6002);
xnor U7099 (N_7099,N_6567,N_6302);
xnor U7100 (N_7100,N_6033,N_6202);
xnor U7101 (N_7101,N_6128,N_6058);
and U7102 (N_7102,N_6168,N_6436);
xor U7103 (N_7103,N_6000,N_6347);
nand U7104 (N_7104,N_6366,N_6533);
and U7105 (N_7105,N_6012,N_6082);
and U7106 (N_7106,N_6358,N_6170);
or U7107 (N_7107,N_6552,N_6133);
or U7108 (N_7108,N_6145,N_6039);
or U7109 (N_7109,N_6278,N_6170);
or U7110 (N_7110,N_6274,N_6213);
nand U7111 (N_7111,N_6502,N_6544);
nor U7112 (N_7112,N_6045,N_6167);
nor U7113 (N_7113,N_6514,N_6158);
nor U7114 (N_7114,N_6096,N_6169);
nand U7115 (N_7115,N_6015,N_6055);
xor U7116 (N_7116,N_6256,N_6516);
nor U7117 (N_7117,N_6086,N_6137);
and U7118 (N_7118,N_6207,N_6536);
or U7119 (N_7119,N_6214,N_6393);
and U7120 (N_7120,N_6552,N_6054);
or U7121 (N_7121,N_6073,N_6327);
and U7122 (N_7122,N_6067,N_6218);
or U7123 (N_7123,N_6166,N_6563);
nand U7124 (N_7124,N_6044,N_6381);
xor U7125 (N_7125,N_6094,N_6312);
nand U7126 (N_7126,N_6001,N_6525);
and U7127 (N_7127,N_6416,N_6500);
xnor U7128 (N_7128,N_6574,N_6065);
nand U7129 (N_7129,N_6465,N_6282);
xor U7130 (N_7130,N_6383,N_6341);
and U7131 (N_7131,N_6312,N_6538);
and U7132 (N_7132,N_6034,N_6507);
xnor U7133 (N_7133,N_6386,N_6502);
and U7134 (N_7134,N_6287,N_6435);
nand U7135 (N_7135,N_6594,N_6595);
xor U7136 (N_7136,N_6567,N_6155);
nand U7137 (N_7137,N_6097,N_6380);
nand U7138 (N_7138,N_6467,N_6302);
xnor U7139 (N_7139,N_6523,N_6484);
xor U7140 (N_7140,N_6312,N_6326);
nor U7141 (N_7141,N_6580,N_6154);
nor U7142 (N_7142,N_6276,N_6298);
and U7143 (N_7143,N_6504,N_6096);
nor U7144 (N_7144,N_6544,N_6285);
xor U7145 (N_7145,N_6504,N_6374);
xnor U7146 (N_7146,N_6563,N_6204);
or U7147 (N_7147,N_6079,N_6547);
nand U7148 (N_7148,N_6550,N_6244);
xnor U7149 (N_7149,N_6315,N_6039);
nor U7150 (N_7150,N_6506,N_6376);
xnor U7151 (N_7151,N_6240,N_6106);
nand U7152 (N_7152,N_6170,N_6547);
and U7153 (N_7153,N_6112,N_6334);
and U7154 (N_7154,N_6175,N_6243);
xnor U7155 (N_7155,N_6264,N_6171);
or U7156 (N_7156,N_6269,N_6477);
xnor U7157 (N_7157,N_6022,N_6018);
nor U7158 (N_7158,N_6558,N_6378);
nor U7159 (N_7159,N_6526,N_6050);
xor U7160 (N_7160,N_6298,N_6479);
and U7161 (N_7161,N_6101,N_6420);
or U7162 (N_7162,N_6058,N_6540);
nor U7163 (N_7163,N_6088,N_6175);
nor U7164 (N_7164,N_6024,N_6342);
nand U7165 (N_7165,N_6043,N_6198);
or U7166 (N_7166,N_6194,N_6446);
and U7167 (N_7167,N_6519,N_6319);
nand U7168 (N_7168,N_6092,N_6380);
xnor U7169 (N_7169,N_6289,N_6207);
xor U7170 (N_7170,N_6562,N_6460);
or U7171 (N_7171,N_6117,N_6402);
and U7172 (N_7172,N_6045,N_6576);
or U7173 (N_7173,N_6277,N_6596);
or U7174 (N_7174,N_6172,N_6136);
nand U7175 (N_7175,N_6302,N_6007);
nand U7176 (N_7176,N_6490,N_6442);
nor U7177 (N_7177,N_6325,N_6042);
xnor U7178 (N_7178,N_6236,N_6191);
xnor U7179 (N_7179,N_6197,N_6489);
or U7180 (N_7180,N_6523,N_6152);
or U7181 (N_7181,N_6322,N_6456);
xnor U7182 (N_7182,N_6150,N_6019);
or U7183 (N_7183,N_6494,N_6457);
and U7184 (N_7184,N_6274,N_6035);
xnor U7185 (N_7185,N_6226,N_6291);
xnor U7186 (N_7186,N_6248,N_6133);
nand U7187 (N_7187,N_6233,N_6340);
nand U7188 (N_7188,N_6158,N_6481);
nor U7189 (N_7189,N_6473,N_6029);
and U7190 (N_7190,N_6182,N_6322);
and U7191 (N_7191,N_6357,N_6323);
or U7192 (N_7192,N_6124,N_6415);
and U7193 (N_7193,N_6076,N_6128);
and U7194 (N_7194,N_6103,N_6440);
nor U7195 (N_7195,N_6479,N_6160);
nand U7196 (N_7196,N_6598,N_6060);
or U7197 (N_7197,N_6341,N_6385);
nor U7198 (N_7198,N_6020,N_6206);
nor U7199 (N_7199,N_6069,N_6217);
xor U7200 (N_7200,N_6682,N_6637);
or U7201 (N_7201,N_7047,N_6776);
nand U7202 (N_7202,N_6835,N_7170);
xnor U7203 (N_7203,N_7117,N_7137);
xor U7204 (N_7204,N_6938,N_6923);
xnor U7205 (N_7205,N_6813,N_6827);
nor U7206 (N_7206,N_6777,N_6804);
xor U7207 (N_7207,N_6905,N_6935);
or U7208 (N_7208,N_6785,N_6801);
nand U7209 (N_7209,N_6947,N_6719);
xor U7210 (N_7210,N_7154,N_6657);
or U7211 (N_7211,N_6939,N_7178);
nor U7212 (N_7212,N_6646,N_6656);
or U7213 (N_7213,N_6618,N_6894);
or U7214 (N_7214,N_6742,N_7066);
nand U7215 (N_7215,N_6796,N_7120);
nand U7216 (N_7216,N_7151,N_6806);
nor U7217 (N_7217,N_6906,N_7173);
and U7218 (N_7218,N_6799,N_7184);
nand U7219 (N_7219,N_6899,N_6976);
or U7220 (N_7220,N_7199,N_6733);
nand U7221 (N_7221,N_6839,N_7038);
or U7222 (N_7222,N_7013,N_6864);
nand U7223 (N_7223,N_6921,N_6766);
nor U7224 (N_7224,N_6875,N_6717);
nor U7225 (N_7225,N_7093,N_6751);
nor U7226 (N_7226,N_6967,N_7022);
and U7227 (N_7227,N_6833,N_7048);
or U7228 (N_7228,N_6709,N_7046);
nor U7229 (N_7229,N_6701,N_6670);
or U7230 (N_7230,N_6746,N_6846);
and U7231 (N_7231,N_6659,N_6972);
or U7232 (N_7232,N_7024,N_7085);
and U7233 (N_7233,N_6830,N_6679);
nor U7234 (N_7234,N_7181,N_7018);
and U7235 (N_7235,N_7135,N_6941);
or U7236 (N_7236,N_7124,N_7052);
nor U7237 (N_7237,N_6778,N_6890);
and U7238 (N_7238,N_6980,N_6691);
or U7239 (N_7239,N_7180,N_6913);
and U7240 (N_7240,N_6997,N_6767);
or U7241 (N_7241,N_6606,N_6655);
and U7242 (N_7242,N_6848,N_7089);
or U7243 (N_7243,N_6869,N_7077);
nand U7244 (N_7244,N_6652,N_6993);
nor U7245 (N_7245,N_6800,N_6769);
and U7246 (N_7246,N_6886,N_7111);
xor U7247 (N_7247,N_6747,N_6603);
nor U7248 (N_7248,N_6915,N_6966);
nor U7249 (N_7249,N_7069,N_7198);
or U7250 (N_7250,N_6863,N_6852);
and U7251 (N_7251,N_7083,N_6953);
and U7252 (N_7252,N_6710,N_6889);
xnor U7253 (N_7253,N_6936,N_6721);
nand U7254 (N_7254,N_6819,N_6964);
nor U7255 (N_7255,N_7056,N_6841);
or U7256 (N_7256,N_7065,N_6859);
xor U7257 (N_7257,N_6832,N_6920);
xor U7258 (N_7258,N_7142,N_7001);
and U7259 (N_7259,N_6943,N_6712);
and U7260 (N_7260,N_7068,N_6698);
nand U7261 (N_7261,N_7175,N_6663);
nand U7262 (N_7262,N_6822,N_7019);
or U7263 (N_7263,N_7165,N_7185);
or U7264 (N_7264,N_6749,N_6836);
or U7265 (N_7265,N_7031,N_6803);
or U7266 (N_7266,N_7164,N_6825);
nand U7267 (N_7267,N_7098,N_6756);
xnor U7268 (N_7268,N_6826,N_7149);
nor U7269 (N_7269,N_6810,N_7009);
nand U7270 (N_7270,N_6881,N_6888);
xor U7271 (N_7271,N_6957,N_7010);
xnor U7272 (N_7272,N_7182,N_7110);
nand U7273 (N_7273,N_7051,N_7121);
or U7274 (N_7274,N_6786,N_7079);
nand U7275 (N_7275,N_6707,N_7166);
nor U7276 (N_7276,N_6926,N_6680);
and U7277 (N_7277,N_7186,N_6843);
xor U7278 (N_7278,N_7043,N_6954);
and U7279 (N_7279,N_6834,N_6688);
xnor U7280 (N_7280,N_7092,N_7067);
or U7281 (N_7281,N_7035,N_7057);
nor U7282 (N_7282,N_6909,N_7195);
and U7283 (N_7283,N_7062,N_6704);
nand U7284 (N_7284,N_6978,N_6610);
nand U7285 (N_7285,N_7141,N_6861);
or U7286 (N_7286,N_7127,N_7090);
nand U7287 (N_7287,N_6986,N_6621);
nor U7288 (N_7288,N_6683,N_6639);
nor U7289 (N_7289,N_6768,N_6837);
xor U7290 (N_7290,N_6728,N_6979);
xnor U7291 (N_7291,N_6672,N_6952);
nor U7292 (N_7292,N_6632,N_6794);
or U7293 (N_7293,N_6916,N_7136);
or U7294 (N_7294,N_7017,N_7116);
and U7295 (N_7295,N_6775,N_7033);
and U7296 (N_7296,N_6734,N_6615);
nand U7297 (N_7297,N_6658,N_6735);
xnor U7298 (N_7298,N_6754,N_7040);
xnor U7299 (N_7299,N_6674,N_7072);
or U7300 (N_7300,N_6622,N_7059);
or U7301 (N_7301,N_6607,N_7091);
nand U7302 (N_7302,N_6910,N_7063);
or U7303 (N_7303,N_6630,N_6629);
nand U7304 (N_7304,N_7000,N_7125);
nand U7305 (N_7305,N_6823,N_7122);
or U7306 (N_7306,N_6922,N_6865);
or U7307 (N_7307,N_6678,N_6608);
xnor U7308 (N_7308,N_7194,N_6809);
nor U7309 (N_7309,N_6872,N_7143);
xor U7310 (N_7310,N_6866,N_6628);
nor U7311 (N_7311,N_7167,N_7037);
nor U7312 (N_7312,N_6983,N_6958);
nand U7313 (N_7313,N_7179,N_7155);
xnor U7314 (N_7314,N_6811,N_6763);
or U7315 (N_7315,N_6697,N_6611);
xnor U7316 (N_7316,N_6927,N_6653);
nor U7317 (N_7317,N_6686,N_6732);
and U7318 (N_7318,N_6878,N_6929);
and U7319 (N_7319,N_6723,N_6940);
xor U7320 (N_7320,N_6605,N_6681);
nor U7321 (N_7321,N_7023,N_6668);
nand U7322 (N_7322,N_7100,N_6842);
and U7323 (N_7323,N_7026,N_7021);
and U7324 (N_7324,N_6812,N_7002);
xnor U7325 (N_7325,N_7115,N_7074);
and U7326 (N_7326,N_6675,N_7188);
and U7327 (N_7327,N_7160,N_6641);
xnor U7328 (N_7328,N_6781,N_6948);
xor U7329 (N_7329,N_6928,N_7109);
and U7330 (N_7330,N_7096,N_6987);
or U7331 (N_7331,N_6654,N_6755);
and U7332 (N_7332,N_6808,N_6759);
or U7333 (N_7333,N_6782,N_6762);
xnor U7334 (N_7334,N_6956,N_6614);
or U7335 (N_7335,N_7144,N_6911);
and U7336 (N_7336,N_6820,N_6669);
and U7337 (N_7337,N_6969,N_6933);
nand U7338 (N_7338,N_6696,N_7041);
or U7339 (N_7339,N_6714,N_6706);
or U7340 (N_7340,N_6792,N_7094);
and U7341 (N_7341,N_7025,N_6718);
or U7342 (N_7342,N_7139,N_7132);
nand U7343 (N_7343,N_7054,N_7020);
xor U7344 (N_7344,N_7118,N_6744);
xnor U7345 (N_7345,N_7045,N_6694);
xor U7346 (N_7346,N_6645,N_7133);
or U7347 (N_7347,N_6844,N_7106);
nand U7348 (N_7348,N_6761,N_7008);
and U7349 (N_7349,N_7140,N_6858);
xor U7350 (N_7350,N_7087,N_6883);
nor U7351 (N_7351,N_6748,N_6772);
or U7352 (N_7352,N_6789,N_6617);
or U7353 (N_7353,N_6838,N_6931);
xnor U7354 (N_7354,N_6725,N_6884);
xnor U7355 (N_7355,N_6612,N_6847);
and U7356 (N_7356,N_6798,N_7168);
xnor U7357 (N_7357,N_6787,N_6918);
xnor U7358 (N_7358,N_6937,N_7055);
xor U7359 (N_7359,N_6671,N_6887);
nand U7360 (N_7360,N_7145,N_6985);
and U7361 (N_7361,N_7028,N_6855);
xnor U7362 (N_7362,N_6739,N_6814);
and U7363 (N_7363,N_6649,N_6934);
and U7364 (N_7364,N_7053,N_6840);
nor U7365 (N_7365,N_7095,N_7119);
nand U7366 (N_7366,N_6616,N_6716);
or U7367 (N_7367,N_7191,N_6713);
xor U7368 (N_7368,N_7150,N_7006);
or U7369 (N_7369,N_7159,N_6973);
nand U7370 (N_7370,N_7003,N_7104);
nor U7371 (N_7371,N_6790,N_6635);
and U7372 (N_7372,N_6895,N_7086);
nand U7373 (N_7373,N_6879,N_6955);
or U7374 (N_7374,N_6908,N_7029);
nor U7375 (N_7375,N_7108,N_6689);
xnor U7376 (N_7376,N_6764,N_7039);
and U7377 (N_7377,N_6974,N_6930);
xor U7378 (N_7378,N_6856,N_6690);
xor U7379 (N_7379,N_7157,N_7058);
and U7380 (N_7380,N_6774,N_6873);
xor U7381 (N_7381,N_6722,N_6788);
nand U7382 (N_7382,N_6932,N_6984);
xor U7383 (N_7383,N_6631,N_6765);
xor U7384 (N_7384,N_6660,N_6780);
xor U7385 (N_7385,N_6850,N_6726);
and U7386 (N_7386,N_6912,N_6745);
or U7387 (N_7387,N_6949,N_6853);
xnor U7388 (N_7388,N_7158,N_7032);
nor U7389 (N_7389,N_6815,N_6602);
nand U7390 (N_7390,N_6893,N_7129);
nor U7391 (N_7391,N_6882,N_7177);
nand U7392 (N_7392,N_6676,N_6634);
nor U7393 (N_7393,N_7183,N_6651);
nand U7394 (N_7394,N_6901,N_7082);
or U7395 (N_7395,N_7004,N_6730);
and U7396 (N_7396,N_6999,N_6871);
nor U7397 (N_7397,N_7070,N_7156);
xnor U7398 (N_7398,N_6693,N_7016);
nor U7399 (N_7399,N_6942,N_6917);
xnor U7400 (N_7400,N_6990,N_6903);
or U7401 (N_7401,N_6977,N_7105);
or U7402 (N_7402,N_6925,N_6770);
nand U7403 (N_7403,N_6849,N_7102);
and U7404 (N_7404,N_7161,N_6867);
or U7405 (N_7405,N_6896,N_6989);
and U7406 (N_7406,N_6946,N_7034);
xor U7407 (N_7407,N_7114,N_7081);
and U7408 (N_7408,N_7097,N_6703);
nand U7409 (N_7409,N_7162,N_6845);
xnor U7410 (N_7410,N_6907,N_7187);
xnor U7411 (N_7411,N_6737,N_6902);
or U7412 (N_7412,N_6664,N_7148);
nor U7413 (N_7413,N_6626,N_6647);
or U7414 (N_7414,N_7075,N_6860);
and U7415 (N_7415,N_7012,N_7197);
nor U7416 (N_7416,N_6944,N_6897);
nor U7417 (N_7417,N_6818,N_6988);
or U7418 (N_7418,N_6880,N_6898);
nor U7419 (N_7419,N_6711,N_6831);
or U7420 (N_7420,N_6661,N_6876);
nor U7421 (N_7421,N_7071,N_6857);
nand U7422 (N_7422,N_6638,N_6817);
nand U7423 (N_7423,N_7131,N_6784);
nand U7424 (N_7424,N_7060,N_6961);
nand U7425 (N_7425,N_6960,N_6900);
nor U7426 (N_7426,N_6662,N_6760);
nor U7427 (N_7427,N_7103,N_6995);
xor U7428 (N_7428,N_6914,N_6919);
nor U7429 (N_7429,N_6684,N_6625);
nand U7430 (N_7430,N_6642,N_7011);
nand U7431 (N_7431,N_6797,N_7015);
xor U7432 (N_7432,N_6891,N_7036);
and U7433 (N_7433,N_6708,N_7169);
and U7434 (N_7434,N_7196,N_6724);
and U7435 (N_7435,N_7171,N_6965);
xnor U7436 (N_7436,N_6624,N_6795);
nor U7437 (N_7437,N_7172,N_6643);
nand U7438 (N_7438,N_7189,N_6620);
and U7439 (N_7439,N_6738,N_7005);
nor U7440 (N_7440,N_6633,N_6874);
and U7441 (N_7441,N_6673,N_6752);
nor U7442 (N_7442,N_6975,N_7163);
and U7443 (N_7443,N_7176,N_6828);
xor U7444 (N_7444,N_6687,N_6962);
and U7445 (N_7445,N_6623,N_6854);
or U7446 (N_7446,N_6779,N_7050);
or U7447 (N_7447,N_6996,N_7126);
or U7448 (N_7448,N_7112,N_6729);
or U7449 (N_7449,N_7049,N_7027);
or U7450 (N_7450,N_6991,N_6600);
nor U7451 (N_7451,N_6702,N_7123);
or U7452 (N_7452,N_6771,N_7044);
xnor U7453 (N_7453,N_6757,N_6720);
and U7454 (N_7454,N_7192,N_7030);
and U7455 (N_7455,N_6793,N_6982);
nor U7456 (N_7456,N_7088,N_7153);
and U7457 (N_7457,N_6971,N_6677);
nand U7458 (N_7458,N_6736,N_6644);
nor U7459 (N_7459,N_6758,N_7078);
nand U7460 (N_7460,N_6715,N_6892);
and U7461 (N_7461,N_6609,N_6731);
and U7462 (N_7462,N_7007,N_6877);
nor U7463 (N_7463,N_6970,N_6998);
and U7464 (N_7464,N_6753,N_6613);
or U7465 (N_7465,N_7174,N_6650);
and U7466 (N_7466,N_6945,N_7073);
and U7467 (N_7467,N_7113,N_7101);
nor U7468 (N_7468,N_6692,N_6695);
xor U7469 (N_7469,N_7146,N_6816);
xnor U7470 (N_7470,N_7128,N_6805);
xnor U7471 (N_7471,N_6741,N_7138);
xor U7472 (N_7472,N_6904,N_6627);
nor U7473 (N_7473,N_6705,N_7014);
nand U7474 (N_7474,N_6868,N_7064);
nand U7475 (N_7475,N_7147,N_6640);
and U7476 (N_7476,N_6601,N_7107);
xnor U7477 (N_7477,N_6791,N_6807);
xnor U7478 (N_7478,N_6665,N_7193);
or U7479 (N_7479,N_6862,N_6667);
nor U7480 (N_7480,N_6783,N_6648);
nor U7481 (N_7481,N_7190,N_6743);
nand U7482 (N_7482,N_6750,N_7152);
xnor U7483 (N_7483,N_6924,N_6802);
and U7484 (N_7484,N_6950,N_6700);
or U7485 (N_7485,N_7134,N_6968);
xnor U7486 (N_7486,N_6870,N_7042);
nand U7487 (N_7487,N_6740,N_7130);
xor U7488 (N_7488,N_6851,N_6829);
nand U7489 (N_7489,N_6699,N_6773);
xor U7490 (N_7490,N_7061,N_6821);
nand U7491 (N_7491,N_6959,N_6992);
or U7492 (N_7492,N_7099,N_6604);
nand U7493 (N_7493,N_6636,N_6981);
and U7494 (N_7494,N_7080,N_7076);
nand U7495 (N_7495,N_6727,N_6619);
nor U7496 (N_7496,N_6994,N_7084);
xor U7497 (N_7497,N_6685,N_6963);
nand U7498 (N_7498,N_6885,N_6824);
or U7499 (N_7499,N_6666,N_6951);
nor U7500 (N_7500,N_6814,N_6841);
nor U7501 (N_7501,N_6785,N_6889);
or U7502 (N_7502,N_6762,N_7117);
xor U7503 (N_7503,N_7094,N_6743);
nand U7504 (N_7504,N_7148,N_6677);
and U7505 (N_7505,N_7058,N_7015);
nand U7506 (N_7506,N_7050,N_6842);
xor U7507 (N_7507,N_7037,N_7029);
xor U7508 (N_7508,N_6829,N_6959);
or U7509 (N_7509,N_7068,N_7050);
xor U7510 (N_7510,N_6795,N_6905);
xnor U7511 (N_7511,N_6837,N_6608);
xor U7512 (N_7512,N_6925,N_7100);
nor U7513 (N_7513,N_6731,N_7105);
nand U7514 (N_7514,N_6993,N_6769);
and U7515 (N_7515,N_6892,N_7029);
or U7516 (N_7516,N_7038,N_6871);
and U7517 (N_7517,N_6979,N_6872);
xor U7518 (N_7518,N_6733,N_6769);
nand U7519 (N_7519,N_6729,N_6775);
nand U7520 (N_7520,N_7010,N_6855);
and U7521 (N_7521,N_6692,N_6915);
xnor U7522 (N_7522,N_6797,N_6900);
or U7523 (N_7523,N_6824,N_6721);
nor U7524 (N_7524,N_6807,N_6909);
or U7525 (N_7525,N_7063,N_6965);
nand U7526 (N_7526,N_6855,N_6900);
nand U7527 (N_7527,N_7021,N_6681);
nor U7528 (N_7528,N_6961,N_6935);
or U7529 (N_7529,N_7151,N_7163);
and U7530 (N_7530,N_6954,N_7036);
nand U7531 (N_7531,N_7135,N_6718);
xnor U7532 (N_7532,N_6780,N_6988);
xnor U7533 (N_7533,N_6937,N_6699);
nand U7534 (N_7534,N_6971,N_6833);
nor U7535 (N_7535,N_7191,N_7045);
nand U7536 (N_7536,N_6881,N_6621);
nand U7537 (N_7537,N_7144,N_6817);
and U7538 (N_7538,N_6883,N_7052);
xnor U7539 (N_7539,N_6647,N_6867);
nand U7540 (N_7540,N_6657,N_6749);
and U7541 (N_7541,N_6989,N_6902);
and U7542 (N_7542,N_6788,N_7130);
nand U7543 (N_7543,N_6645,N_6988);
and U7544 (N_7544,N_6951,N_7005);
or U7545 (N_7545,N_6737,N_6820);
nor U7546 (N_7546,N_6964,N_7134);
xor U7547 (N_7547,N_6734,N_7159);
xnor U7548 (N_7548,N_7168,N_6687);
xor U7549 (N_7549,N_7111,N_7150);
nor U7550 (N_7550,N_6947,N_6989);
xor U7551 (N_7551,N_7047,N_7154);
or U7552 (N_7552,N_7140,N_6998);
or U7553 (N_7553,N_6727,N_7002);
and U7554 (N_7554,N_7100,N_6644);
xor U7555 (N_7555,N_6832,N_6910);
and U7556 (N_7556,N_6669,N_7162);
nand U7557 (N_7557,N_7038,N_6624);
and U7558 (N_7558,N_6868,N_6684);
and U7559 (N_7559,N_6743,N_6861);
and U7560 (N_7560,N_6636,N_7129);
nand U7561 (N_7561,N_6640,N_6694);
or U7562 (N_7562,N_7006,N_6896);
nand U7563 (N_7563,N_6812,N_6608);
xor U7564 (N_7564,N_6981,N_6606);
nor U7565 (N_7565,N_7148,N_6948);
nand U7566 (N_7566,N_7103,N_6784);
xor U7567 (N_7567,N_6884,N_6802);
nor U7568 (N_7568,N_6751,N_6675);
or U7569 (N_7569,N_6739,N_7011);
nor U7570 (N_7570,N_6952,N_7019);
or U7571 (N_7571,N_7160,N_7126);
or U7572 (N_7572,N_7132,N_7172);
and U7573 (N_7573,N_6683,N_6945);
nor U7574 (N_7574,N_6648,N_6644);
or U7575 (N_7575,N_7128,N_6663);
or U7576 (N_7576,N_6988,N_6689);
nand U7577 (N_7577,N_6699,N_7083);
nor U7578 (N_7578,N_7145,N_7075);
nor U7579 (N_7579,N_6610,N_7057);
or U7580 (N_7580,N_7025,N_7134);
xor U7581 (N_7581,N_7161,N_7031);
nand U7582 (N_7582,N_6922,N_7163);
nor U7583 (N_7583,N_6806,N_6867);
nand U7584 (N_7584,N_6994,N_6697);
nor U7585 (N_7585,N_6731,N_6870);
and U7586 (N_7586,N_6651,N_6961);
nor U7587 (N_7587,N_6660,N_6959);
nor U7588 (N_7588,N_7019,N_7065);
nand U7589 (N_7589,N_6625,N_7134);
or U7590 (N_7590,N_6687,N_7029);
nand U7591 (N_7591,N_6942,N_6651);
xnor U7592 (N_7592,N_7154,N_7086);
nand U7593 (N_7593,N_7090,N_7140);
or U7594 (N_7594,N_7169,N_6781);
and U7595 (N_7595,N_6843,N_6930);
nand U7596 (N_7596,N_6937,N_6671);
or U7597 (N_7597,N_6718,N_6818);
nand U7598 (N_7598,N_7131,N_6906);
or U7599 (N_7599,N_7013,N_6977);
and U7600 (N_7600,N_6826,N_6825);
and U7601 (N_7601,N_6682,N_6640);
or U7602 (N_7602,N_6737,N_7079);
xnor U7603 (N_7603,N_6900,N_6787);
nand U7604 (N_7604,N_6823,N_7017);
or U7605 (N_7605,N_6652,N_6840);
or U7606 (N_7606,N_7124,N_6790);
nor U7607 (N_7607,N_7016,N_7012);
nor U7608 (N_7608,N_6753,N_6602);
xnor U7609 (N_7609,N_6749,N_6805);
nor U7610 (N_7610,N_6682,N_6723);
xnor U7611 (N_7611,N_7178,N_7047);
xnor U7612 (N_7612,N_6694,N_6821);
nand U7613 (N_7613,N_6707,N_7180);
nand U7614 (N_7614,N_7073,N_7100);
nand U7615 (N_7615,N_6690,N_7059);
or U7616 (N_7616,N_6890,N_7141);
nand U7617 (N_7617,N_6900,N_6905);
or U7618 (N_7618,N_6681,N_6893);
nor U7619 (N_7619,N_7036,N_6746);
nor U7620 (N_7620,N_7068,N_7112);
nor U7621 (N_7621,N_6932,N_7194);
and U7622 (N_7622,N_6600,N_7136);
and U7623 (N_7623,N_7046,N_7127);
and U7624 (N_7624,N_6605,N_6842);
and U7625 (N_7625,N_7037,N_7005);
nand U7626 (N_7626,N_6810,N_6840);
and U7627 (N_7627,N_6759,N_7160);
or U7628 (N_7628,N_6885,N_6965);
nor U7629 (N_7629,N_6603,N_6848);
nand U7630 (N_7630,N_6882,N_6952);
nor U7631 (N_7631,N_6678,N_6778);
nor U7632 (N_7632,N_7070,N_6918);
and U7633 (N_7633,N_6766,N_6747);
or U7634 (N_7634,N_6996,N_6601);
nor U7635 (N_7635,N_7010,N_7058);
or U7636 (N_7636,N_6618,N_6693);
xor U7637 (N_7637,N_7110,N_6637);
nand U7638 (N_7638,N_6976,N_6920);
xnor U7639 (N_7639,N_7044,N_6699);
xor U7640 (N_7640,N_6624,N_6929);
xnor U7641 (N_7641,N_6686,N_7099);
and U7642 (N_7642,N_7119,N_7072);
nand U7643 (N_7643,N_6720,N_6691);
and U7644 (N_7644,N_7077,N_7172);
xor U7645 (N_7645,N_6648,N_6870);
and U7646 (N_7646,N_6980,N_6666);
and U7647 (N_7647,N_7020,N_6779);
nor U7648 (N_7648,N_6918,N_6850);
nor U7649 (N_7649,N_6828,N_6793);
and U7650 (N_7650,N_6868,N_6998);
or U7651 (N_7651,N_6817,N_7046);
xnor U7652 (N_7652,N_6889,N_7049);
or U7653 (N_7653,N_6625,N_6916);
nand U7654 (N_7654,N_6973,N_6971);
or U7655 (N_7655,N_6789,N_6719);
and U7656 (N_7656,N_7115,N_6718);
nor U7657 (N_7657,N_6938,N_6790);
xor U7658 (N_7658,N_7053,N_7013);
or U7659 (N_7659,N_6837,N_6799);
or U7660 (N_7660,N_6934,N_6918);
or U7661 (N_7661,N_7141,N_6934);
nand U7662 (N_7662,N_6984,N_6819);
and U7663 (N_7663,N_6699,N_7063);
nand U7664 (N_7664,N_7073,N_6605);
and U7665 (N_7665,N_6826,N_7122);
xor U7666 (N_7666,N_6803,N_7131);
nor U7667 (N_7667,N_6911,N_6696);
and U7668 (N_7668,N_6962,N_7087);
nor U7669 (N_7669,N_7079,N_6732);
or U7670 (N_7670,N_6801,N_6855);
nand U7671 (N_7671,N_7174,N_6842);
or U7672 (N_7672,N_6870,N_6954);
nor U7673 (N_7673,N_6871,N_6856);
and U7674 (N_7674,N_6750,N_6650);
xnor U7675 (N_7675,N_6954,N_7066);
or U7676 (N_7676,N_6649,N_7044);
xor U7677 (N_7677,N_7058,N_6927);
or U7678 (N_7678,N_6635,N_6975);
or U7679 (N_7679,N_6976,N_6758);
nand U7680 (N_7680,N_6903,N_6874);
or U7681 (N_7681,N_7131,N_6639);
or U7682 (N_7682,N_7002,N_6883);
or U7683 (N_7683,N_6661,N_7074);
nor U7684 (N_7684,N_7096,N_7107);
xor U7685 (N_7685,N_7170,N_6782);
or U7686 (N_7686,N_7130,N_7146);
xnor U7687 (N_7687,N_6790,N_7167);
or U7688 (N_7688,N_6986,N_6609);
and U7689 (N_7689,N_6881,N_6969);
xnor U7690 (N_7690,N_6910,N_6646);
nand U7691 (N_7691,N_6643,N_6915);
xnor U7692 (N_7692,N_6727,N_6833);
or U7693 (N_7693,N_6623,N_7166);
nand U7694 (N_7694,N_7055,N_6619);
and U7695 (N_7695,N_7048,N_6896);
nand U7696 (N_7696,N_7084,N_6685);
and U7697 (N_7697,N_6708,N_6872);
nor U7698 (N_7698,N_7023,N_6971);
and U7699 (N_7699,N_6748,N_6605);
xnor U7700 (N_7700,N_6996,N_6717);
xnor U7701 (N_7701,N_7190,N_7001);
nand U7702 (N_7702,N_6752,N_6784);
nand U7703 (N_7703,N_6770,N_7133);
xor U7704 (N_7704,N_7142,N_6816);
xor U7705 (N_7705,N_6763,N_7174);
xnor U7706 (N_7706,N_7039,N_6694);
nand U7707 (N_7707,N_7118,N_7106);
nor U7708 (N_7708,N_7176,N_6888);
or U7709 (N_7709,N_6860,N_6829);
or U7710 (N_7710,N_6729,N_6984);
or U7711 (N_7711,N_7067,N_6869);
nand U7712 (N_7712,N_6750,N_6815);
or U7713 (N_7713,N_7162,N_7022);
xor U7714 (N_7714,N_6717,N_6936);
or U7715 (N_7715,N_7029,N_7052);
nor U7716 (N_7716,N_7047,N_6692);
or U7717 (N_7717,N_6989,N_6817);
nand U7718 (N_7718,N_7146,N_7078);
nand U7719 (N_7719,N_6647,N_7141);
and U7720 (N_7720,N_6632,N_6908);
xnor U7721 (N_7721,N_7104,N_6649);
nor U7722 (N_7722,N_6676,N_6824);
xnor U7723 (N_7723,N_6838,N_7003);
nor U7724 (N_7724,N_7145,N_6945);
nor U7725 (N_7725,N_7137,N_7020);
or U7726 (N_7726,N_6640,N_6925);
xor U7727 (N_7727,N_6849,N_6683);
and U7728 (N_7728,N_6762,N_6823);
nor U7729 (N_7729,N_6775,N_6914);
nor U7730 (N_7730,N_6666,N_7128);
or U7731 (N_7731,N_7115,N_6902);
nor U7732 (N_7732,N_7164,N_6979);
nor U7733 (N_7733,N_7059,N_6638);
or U7734 (N_7734,N_6931,N_6769);
and U7735 (N_7735,N_6848,N_6785);
and U7736 (N_7736,N_7083,N_6935);
xor U7737 (N_7737,N_6936,N_6720);
nand U7738 (N_7738,N_6979,N_7168);
nand U7739 (N_7739,N_7130,N_6936);
nand U7740 (N_7740,N_6932,N_7069);
or U7741 (N_7741,N_6739,N_6659);
xor U7742 (N_7742,N_6845,N_6932);
and U7743 (N_7743,N_7161,N_6632);
and U7744 (N_7744,N_7107,N_7060);
xnor U7745 (N_7745,N_7058,N_6970);
or U7746 (N_7746,N_7101,N_7197);
nor U7747 (N_7747,N_7032,N_7079);
nand U7748 (N_7748,N_6925,N_7029);
nand U7749 (N_7749,N_7089,N_7007);
or U7750 (N_7750,N_6744,N_7061);
and U7751 (N_7751,N_6814,N_6899);
and U7752 (N_7752,N_6873,N_7135);
nor U7753 (N_7753,N_6646,N_6692);
nand U7754 (N_7754,N_7023,N_6979);
and U7755 (N_7755,N_6782,N_7072);
nor U7756 (N_7756,N_6741,N_6778);
and U7757 (N_7757,N_6694,N_6866);
nor U7758 (N_7758,N_6664,N_6980);
and U7759 (N_7759,N_7142,N_6711);
xnor U7760 (N_7760,N_6686,N_7134);
nor U7761 (N_7761,N_6695,N_7010);
or U7762 (N_7762,N_6951,N_7111);
or U7763 (N_7763,N_6787,N_6605);
or U7764 (N_7764,N_7024,N_6603);
nor U7765 (N_7765,N_6775,N_6955);
nor U7766 (N_7766,N_6885,N_7017);
or U7767 (N_7767,N_7112,N_6942);
nor U7768 (N_7768,N_6681,N_7153);
nand U7769 (N_7769,N_6708,N_7082);
xnor U7770 (N_7770,N_7084,N_6668);
and U7771 (N_7771,N_7013,N_6607);
and U7772 (N_7772,N_6840,N_6780);
xnor U7773 (N_7773,N_6911,N_6759);
nor U7774 (N_7774,N_7013,N_6618);
or U7775 (N_7775,N_6619,N_7085);
nor U7776 (N_7776,N_7050,N_7089);
nand U7777 (N_7777,N_6679,N_6898);
or U7778 (N_7778,N_6722,N_6735);
or U7779 (N_7779,N_6616,N_6677);
and U7780 (N_7780,N_7164,N_7193);
xnor U7781 (N_7781,N_7135,N_7039);
nand U7782 (N_7782,N_6829,N_6703);
xor U7783 (N_7783,N_6883,N_6999);
nor U7784 (N_7784,N_7188,N_6799);
xnor U7785 (N_7785,N_6886,N_6784);
and U7786 (N_7786,N_6818,N_6874);
nor U7787 (N_7787,N_6930,N_6710);
nand U7788 (N_7788,N_6801,N_6724);
and U7789 (N_7789,N_6831,N_6759);
nor U7790 (N_7790,N_6959,N_6938);
nand U7791 (N_7791,N_6863,N_7089);
xor U7792 (N_7792,N_6618,N_6759);
nor U7793 (N_7793,N_7090,N_7151);
nand U7794 (N_7794,N_7012,N_6827);
xnor U7795 (N_7795,N_6940,N_6738);
nor U7796 (N_7796,N_6915,N_6812);
or U7797 (N_7797,N_6736,N_6623);
or U7798 (N_7798,N_6811,N_6815);
xnor U7799 (N_7799,N_6607,N_6662);
and U7800 (N_7800,N_7253,N_7772);
or U7801 (N_7801,N_7743,N_7278);
xnor U7802 (N_7802,N_7474,N_7704);
xnor U7803 (N_7803,N_7541,N_7555);
xnor U7804 (N_7804,N_7204,N_7207);
nand U7805 (N_7805,N_7619,N_7244);
nor U7806 (N_7806,N_7258,N_7450);
nor U7807 (N_7807,N_7586,N_7697);
or U7808 (N_7808,N_7436,N_7770);
or U7809 (N_7809,N_7352,N_7344);
nor U7810 (N_7810,N_7599,N_7625);
xnor U7811 (N_7811,N_7415,N_7326);
or U7812 (N_7812,N_7791,N_7659);
nor U7813 (N_7813,N_7446,N_7227);
nor U7814 (N_7814,N_7384,N_7543);
xor U7815 (N_7815,N_7329,N_7390);
nor U7816 (N_7816,N_7486,N_7705);
nor U7817 (N_7817,N_7714,N_7279);
and U7818 (N_7818,N_7289,N_7441);
and U7819 (N_7819,N_7476,N_7201);
or U7820 (N_7820,N_7414,N_7660);
xor U7821 (N_7821,N_7257,N_7623);
nor U7822 (N_7822,N_7669,N_7615);
and U7823 (N_7823,N_7638,N_7358);
or U7824 (N_7824,N_7229,N_7317);
xnor U7825 (N_7825,N_7367,N_7608);
and U7826 (N_7826,N_7387,N_7473);
and U7827 (N_7827,N_7311,N_7696);
nor U7828 (N_7828,N_7266,N_7688);
xor U7829 (N_7829,N_7342,N_7325);
and U7830 (N_7830,N_7375,N_7790);
nand U7831 (N_7831,N_7232,N_7652);
nor U7832 (N_7832,N_7636,N_7693);
nand U7833 (N_7833,N_7215,N_7685);
nor U7834 (N_7834,N_7760,N_7742);
and U7835 (N_7835,N_7573,N_7559);
nor U7836 (N_7836,N_7549,N_7618);
or U7837 (N_7837,N_7509,N_7613);
and U7838 (N_7838,N_7202,N_7241);
xnor U7839 (N_7839,N_7297,N_7340);
nand U7840 (N_7840,N_7260,N_7591);
and U7841 (N_7841,N_7456,N_7631);
and U7842 (N_7842,N_7723,N_7682);
nand U7843 (N_7843,N_7745,N_7418);
xor U7844 (N_7844,N_7264,N_7280);
nand U7845 (N_7845,N_7491,N_7489);
or U7846 (N_7846,N_7678,N_7356);
nor U7847 (N_7847,N_7656,N_7767);
xnor U7848 (N_7848,N_7233,N_7612);
xor U7849 (N_7849,N_7265,N_7649);
nand U7850 (N_7850,N_7262,N_7601);
or U7851 (N_7851,N_7210,N_7710);
nor U7852 (N_7852,N_7249,N_7251);
xor U7853 (N_7853,N_7464,N_7263);
nor U7854 (N_7854,N_7679,N_7381);
or U7855 (N_7855,N_7488,N_7468);
nor U7856 (N_7856,N_7518,N_7754);
and U7857 (N_7857,N_7411,N_7554);
xnor U7858 (N_7858,N_7577,N_7642);
or U7859 (N_7859,N_7434,N_7552);
xnor U7860 (N_7860,N_7235,N_7788);
or U7861 (N_7861,N_7479,N_7421);
or U7862 (N_7862,N_7350,N_7542);
xnor U7863 (N_7863,N_7359,N_7664);
nor U7864 (N_7864,N_7432,N_7724);
or U7865 (N_7865,N_7459,N_7548);
xnor U7866 (N_7866,N_7451,N_7399);
nor U7867 (N_7867,N_7789,N_7256);
nor U7868 (N_7868,N_7563,N_7515);
or U7869 (N_7869,N_7483,N_7400);
or U7870 (N_7870,N_7639,N_7501);
and U7871 (N_7871,N_7794,N_7331);
nor U7872 (N_7872,N_7602,N_7598);
xnor U7873 (N_7873,N_7547,N_7480);
nor U7874 (N_7874,N_7521,N_7394);
nor U7875 (N_7875,N_7334,N_7578);
or U7876 (N_7876,N_7620,N_7460);
nor U7877 (N_7877,N_7597,N_7644);
or U7878 (N_7878,N_7449,N_7301);
xor U7879 (N_7879,N_7641,N_7646);
or U7880 (N_7880,N_7707,N_7208);
nand U7881 (N_7881,N_7741,N_7269);
or U7882 (N_7882,N_7640,N_7778);
nand U7883 (N_7883,N_7309,N_7594);
and U7884 (N_7884,N_7799,N_7261);
nor U7885 (N_7885,N_7600,N_7429);
xnor U7886 (N_7886,N_7243,N_7252);
nand U7887 (N_7887,N_7274,N_7703);
nor U7888 (N_7888,N_7628,N_7445);
xor U7889 (N_7889,N_7545,N_7632);
and U7890 (N_7890,N_7226,N_7477);
nor U7891 (N_7891,N_7609,N_7593);
nor U7892 (N_7892,N_7712,N_7397);
xor U7893 (N_7893,N_7672,N_7512);
or U7894 (N_7894,N_7516,N_7708);
nor U7895 (N_7895,N_7439,N_7291);
nor U7896 (N_7896,N_7321,N_7223);
nor U7897 (N_7897,N_7647,N_7587);
nor U7898 (N_7898,N_7629,N_7428);
xor U7899 (N_7899,N_7268,N_7240);
nor U7900 (N_7900,N_7282,N_7690);
and U7901 (N_7901,N_7401,N_7295);
nor U7902 (N_7902,N_7348,N_7746);
and U7903 (N_7903,N_7292,N_7630);
xnor U7904 (N_7904,N_7315,N_7218);
nand U7905 (N_7905,N_7405,N_7306);
and U7906 (N_7906,N_7701,N_7654);
nand U7907 (N_7907,N_7270,N_7308);
nor U7908 (N_7908,N_7718,N_7404);
and U7909 (N_7909,N_7395,N_7335);
and U7910 (N_7910,N_7683,N_7485);
or U7911 (N_7911,N_7546,N_7569);
and U7912 (N_7912,N_7444,N_7376);
xor U7913 (N_7913,N_7389,N_7287);
or U7914 (N_7914,N_7369,N_7290);
nand U7915 (N_7915,N_7231,N_7592);
nand U7916 (N_7916,N_7667,N_7499);
xor U7917 (N_7917,N_7374,N_7737);
xnor U7918 (N_7918,N_7528,N_7595);
nor U7919 (N_7919,N_7753,N_7782);
xor U7920 (N_7920,N_7527,N_7795);
nand U7921 (N_7921,N_7645,N_7273);
and U7922 (N_7922,N_7379,N_7526);
nand U7923 (N_7923,N_7313,N_7302);
xnor U7924 (N_7924,N_7764,N_7493);
nor U7925 (N_7925,N_7506,N_7368);
nand U7926 (N_7926,N_7427,N_7779);
nand U7927 (N_7927,N_7582,N_7346);
nor U7928 (N_7928,N_7706,N_7420);
nor U7929 (N_7929,N_7467,N_7328);
nor U7930 (N_7930,N_7386,N_7382);
nor U7931 (N_7931,N_7700,N_7607);
or U7932 (N_7932,N_7373,N_7665);
and U7933 (N_7933,N_7637,N_7220);
xnor U7934 (N_7934,N_7378,N_7517);
xor U7935 (N_7935,N_7733,N_7663);
or U7936 (N_7936,N_7355,N_7787);
and U7937 (N_7937,N_7579,N_7729);
xnor U7938 (N_7938,N_7503,N_7716);
nand U7939 (N_7939,N_7206,N_7380);
nand U7940 (N_7940,N_7588,N_7440);
and U7941 (N_7941,N_7529,N_7622);
and U7942 (N_7942,N_7205,N_7730);
and U7943 (N_7943,N_7699,N_7761);
or U7944 (N_7944,N_7254,N_7353);
nand U7945 (N_7945,N_7551,N_7424);
and U7946 (N_7946,N_7722,N_7341);
xor U7947 (N_7947,N_7463,N_7447);
and U7948 (N_7948,N_7225,N_7633);
nor U7949 (N_7949,N_7316,N_7255);
nor U7950 (N_7950,N_7650,N_7371);
nand U7951 (N_7951,N_7417,N_7357);
or U7952 (N_7952,N_7203,N_7583);
and U7953 (N_7953,N_7366,N_7388);
or U7954 (N_7954,N_7423,N_7322);
or U7955 (N_7955,N_7361,N_7777);
or U7956 (N_7956,N_7475,N_7272);
xor U7957 (N_7957,N_7458,N_7466);
nand U7958 (N_7958,N_7532,N_7674);
nand U7959 (N_7959,N_7435,N_7748);
nand U7960 (N_7960,N_7259,N_7310);
xnor U7961 (N_7961,N_7749,N_7336);
and U7962 (N_7962,N_7500,N_7771);
nand U7963 (N_7963,N_7416,N_7568);
or U7964 (N_7964,N_7318,N_7481);
xnor U7965 (N_7965,N_7438,N_7616);
nand U7966 (N_7966,N_7585,N_7286);
and U7967 (N_7967,N_7472,N_7237);
and U7968 (N_7968,N_7453,N_7402);
xor U7969 (N_7969,N_7570,N_7731);
or U7970 (N_7970,N_7603,N_7792);
nand U7971 (N_7971,N_7673,N_7238);
nor U7972 (N_7972,N_7433,N_7363);
nor U7973 (N_7973,N_7413,N_7419);
nand U7974 (N_7974,N_7470,N_7497);
xor U7975 (N_7975,N_7455,N_7740);
nor U7976 (N_7976,N_7695,N_7755);
and U7977 (N_7977,N_7478,N_7285);
and U7978 (N_7978,N_7303,N_7756);
nand U7979 (N_7979,N_7412,N_7560);
nand U7980 (N_7980,N_7236,N_7702);
and U7981 (N_7981,N_7604,N_7393);
nand U7982 (N_7982,N_7377,N_7511);
xnor U7983 (N_7983,N_7635,N_7490);
nand U7984 (N_7984,N_7655,N_7200);
nor U7985 (N_7985,N_7530,N_7589);
and U7986 (N_7986,N_7362,N_7610);
nand U7987 (N_7987,N_7314,N_7648);
xnor U7988 (N_7988,N_7298,N_7747);
and U7989 (N_7989,N_7797,N_7658);
or U7990 (N_7990,N_7796,N_7343);
and U7991 (N_7991,N_7522,N_7495);
nand U7992 (N_7992,N_7752,N_7798);
nor U7993 (N_7993,N_7296,N_7567);
or U7994 (N_7994,N_7680,N_7276);
and U7995 (N_7995,N_7294,N_7461);
nor U7996 (N_7996,N_7535,N_7606);
and U7997 (N_7997,N_7250,N_7538);
and U7998 (N_7998,N_7735,N_7721);
nand U7999 (N_7999,N_7793,N_7662);
and U8000 (N_8000,N_7739,N_7245);
xor U8001 (N_8001,N_7768,N_7692);
nor U8002 (N_8002,N_7720,N_7626);
or U8003 (N_8003,N_7557,N_7507);
nor U8004 (N_8004,N_7784,N_7726);
and U8005 (N_8005,N_7514,N_7617);
and U8006 (N_8006,N_7719,N_7759);
and U8007 (N_8007,N_7339,N_7403);
nor U8008 (N_8008,N_7383,N_7327);
nor U8009 (N_8009,N_7406,N_7581);
nand U8010 (N_8010,N_7533,N_7725);
xor U8011 (N_8011,N_7769,N_7671);
or U8012 (N_8012,N_7482,N_7448);
and U8013 (N_8013,N_7324,N_7410);
xnor U8014 (N_8014,N_7687,N_7347);
or U8015 (N_8015,N_7305,N_7275);
or U8016 (N_8016,N_7525,N_7694);
or U8017 (N_8017,N_7624,N_7775);
and U8018 (N_8018,N_7561,N_7469);
nor U8019 (N_8019,N_7580,N_7409);
nor U8020 (N_8020,N_7364,N_7247);
and U8021 (N_8021,N_7681,N_7214);
xnor U8022 (N_8022,N_7452,N_7596);
xor U8023 (N_8023,N_7575,N_7283);
nand U8024 (N_8024,N_7426,N_7657);
nor U8025 (N_8025,N_7430,N_7698);
and U8026 (N_8026,N_7744,N_7323);
xor U8027 (N_8027,N_7653,N_7216);
nand U8028 (N_8028,N_7277,N_7536);
nand U8029 (N_8029,N_7462,N_7300);
xor U8030 (N_8030,N_7571,N_7246);
nor U8031 (N_8031,N_7727,N_7565);
or U8032 (N_8032,N_7267,N_7299);
nand U8033 (N_8033,N_7677,N_7763);
nor U8034 (N_8034,N_7407,N_7312);
and U8035 (N_8035,N_7354,N_7540);
nor U8036 (N_8036,N_7239,N_7553);
or U8037 (N_8037,N_7751,N_7242);
or U8038 (N_8038,N_7709,N_7392);
or U8039 (N_8039,N_7562,N_7513);
or U8040 (N_8040,N_7457,N_7614);
or U8041 (N_8041,N_7684,N_7284);
nand U8042 (N_8042,N_7213,N_7398);
and U8043 (N_8043,N_7391,N_7487);
and U8044 (N_8044,N_7785,N_7307);
or U8045 (N_8045,N_7519,N_7711);
and U8046 (N_8046,N_7564,N_7550);
xor U8047 (N_8047,N_7750,N_7337);
nand U8048 (N_8048,N_7734,N_7271);
nand U8049 (N_8049,N_7627,N_7502);
xnor U8050 (N_8050,N_7661,N_7523);
and U8051 (N_8051,N_7209,N_7691);
nor U8052 (N_8052,N_7281,N_7780);
nor U8053 (N_8053,N_7576,N_7773);
nor U8054 (N_8054,N_7230,N_7496);
and U8055 (N_8055,N_7492,N_7221);
nand U8056 (N_8056,N_7320,N_7385);
nand U8057 (N_8057,N_7471,N_7670);
and U8058 (N_8058,N_7776,N_7634);
and U8059 (N_8059,N_7224,N_7572);
and U8060 (N_8060,N_7370,N_7584);
nand U8061 (N_8061,N_7228,N_7781);
or U8062 (N_8062,N_7234,N_7666);
or U8063 (N_8063,N_7715,N_7786);
nor U8064 (N_8064,N_7574,N_7349);
nor U8065 (N_8065,N_7766,N_7774);
or U8066 (N_8066,N_7211,N_7333);
nand U8067 (N_8067,N_7222,N_7504);
nand U8068 (N_8068,N_7425,N_7611);
and U8069 (N_8069,N_7676,N_7360);
nor U8070 (N_8070,N_7465,N_7408);
or U8071 (N_8071,N_7686,N_7544);
xor U8072 (N_8072,N_7248,N_7498);
xnor U8073 (N_8073,N_7304,N_7713);
nor U8074 (N_8074,N_7765,N_7484);
nor U8075 (N_8075,N_7288,N_7728);
nor U8076 (N_8076,N_7330,N_7442);
xor U8077 (N_8077,N_7605,N_7621);
and U8078 (N_8078,N_7422,N_7351);
or U8079 (N_8079,N_7431,N_7556);
xnor U8080 (N_8080,N_7531,N_7675);
nor U8081 (N_8081,N_7437,N_7293);
xnor U8082 (N_8082,N_7668,N_7365);
and U8083 (N_8083,N_7520,N_7396);
and U8084 (N_8084,N_7510,N_7534);
xnor U8085 (N_8085,N_7783,N_7643);
or U8086 (N_8086,N_7494,N_7508);
nand U8087 (N_8087,N_7558,N_7590);
nor U8088 (N_8088,N_7717,N_7372);
nand U8089 (N_8089,N_7338,N_7332);
nand U8090 (N_8090,N_7732,N_7219);
nor U8091 (N_8091,N_7319,N_7217);
and U8092 (N_8092,N_7762,N_7689);
or U8093 (N_8093,N_7524,N_7736);
nand U8094 (N_8094,N_7757,N_7505);
or U8095 (N_8095,N_7443,N_7539);
nor U8096 (N_8096,N_7738,N_7345);
nor U8097 (N_8097,N_7212,N_7758);
nor U8098 (N_8098,N_7651,N_7454);
or U8099 (N_8099,N_7566,N_7537);
nor U8100 (N_8100,N_7423,N_7799);
and U8101 (N_8101,N_7710,N_7504);
or U8102 (N_8102,N_7295,N_7484);
and U8103 (N_8103,N_7433,N_7704);
and U8104 (N_8104,N_7759,N_7723);
or U8105 (N_8105,N_7428,N_7602);
or U8106 (N_8106,N_7396,N_7420);
xor U8107 (N_8107,N_7286,N_7797);
nand U8108 (N_8108,N_7592,N_7282);
and U8109 (N_8109,N_7538,N_7720);
xor U8110 (N_8110,N_7778,N_7334);
and U8111 (N_8111,N_7412,N_7744);
nand U8112 (N_8112,N_7587,N_7767);
or U8113 (N_8113,N_7493,N_7262);
nand U8114 (N_8114,N_7415,N_7330);
nor U8115 (N_8115,N_7648,N_7409);
xor U8116 (N_8116,N_7450,N_7498);
nand U8117 (N_8117,N_7252,N_7429);
or U8118 (N_8118,N_7480,N_7479);
and U8119 (N_8119,N_7390,N_7737);
nand U8120 (N_8120,N_7307,N_7583);
xnor U8121 (N_8121,N_7324,N_7386);
xnor U8122 (N_8122,N_7534,N_7420);
nand U8123 (N_8123,N_7772,N_7464);
and U8124 (N_8124,N_7517,N_7715);
and U8125 (N_8125,N_7745,N_7571);
nand U8126 (N_8126,N_7704,N_7388);
xnor U8127 (N_8127,N_7635,N_7688);
nand U8128 (N_8128,N_7753,N_7275);
nand U8129 (N_8129,N_7328,N_7440);
or U8130 (N_8130,N_7603,N_7368);
nor U8131 (N_8131,N_7655,N_7452);
or U8132 (N_8132,N_7488,N_7446);
nand U8133 (N_8133,N_7679,N_7462);
and U8134 (N_8134,N_7257,N_7353);
nand U8135 (N_8135,N_7259,N_7496);
nor U8136 (N_8136,N_7226,N_7202);
or U8137 (N_8137,N_7242,N_7323);
nand U8138 (N_8138,N_7206,N_7734);
xor U8139 (N_8139,N_7441,N_7507);
nand U8140 (N_8140,N_7552,N_7791);
or U8141 (N_8141,N_7761,N_7379);
nor U8142 (N_8142,N_7601,N_7415);
and U8143 (N_8143,N_7552,N_7673);
nand U8144 (N_8144,N_7576,N_7327);
xor U8145 (N_8145,N_7256,N_7578);
nor U8146 (N_8146,N_7474,N_7224);
xor U8147 (N_8147,N_7599,N_7593);
nor U8148 (N_8148,N_7259,N_7605);
or U8149 (N_8149,N_7743,N_7638);
nor U8150 (N_8150,N_7690,N_7547);
xnor U8151 (N_8151,N_7577,N_7736);
or U8152 (N_8152,N_7369,N_7367);
xnor U8153 (N_8153,N_7580,N_7628);
xnor U8154 (N_8154,N_7362,N_7518);
nor U8155 (N_8155,N_7248,N_7342);
nor U8156 (N_8156,N_7513,N_7258);
xor U8157 (N_8157,N_7535,N_7588);
or U8158 (N_8158,N_7521,N_7772);
and U8159 (N_8159,N_7393,N_7581);
or U8160 (N_8160,N_7633,N_7362);
nor U8161 (N_8161,N_7397,N_7674);
nor U8162 (N_8162,N_7757,N_7496);
xor U8163 (N_8163,N_7404,N_7254);
and U8164 (N_8164,N_7249,N_7446);
or U8165 (N_8165,N_7627,N_7595);
and U8166 (N_8166,N_7267,N_7419);
and U8167 (N_8167,N_7791,N_7715);
or U8168 (N_8168,N_7400,N_7613);
nor U8169 (N_8169,N_7658,N_7657);
nand U8170 (N_8170,N_7717,N_7553);
nor U8171 (N_8171,N_7345,N_7734);
xnor U8172 (N_8172,N_7721,N_7797);
nand U8173 (N_8173,N_7775,N_7614);
xor U8174 (N_8174,N_7556,N_7791);
nor U8175 (N_8175,N_7367,N_7704);
and U8176 (N_8176,N_7459,N_7370);
and U8177 (N_8177,N_7519,N_7441);
nor U8178 (N_8178,N_7572,N_7764);
xnor U8179 (N_8179,N_7609,N_7783);
nand U8180 (N_8180,N_7378,N_7776);
nor U8181 (N_8181,N_7296,N_7585);
and U8182 (N_8182,N_7280,N_7605);
xor U8183 (N_8183,N_7620,N_7462);
and U8184 (N_8184,N_7677,N_7799);
or U8185 (N_8185,N_7700,N_7296);
xor U8186 (N_8186,N_7620,N_7738);
and U8187 (N_8187,N_7374,N_7556);
and U8188 (N_8188,N_7476,N_7355);
nor U8189 (N_8189,N_7702,N_7284);
or U8190 (N_8190,N_7227,N_7619);
nand U8191 (N_8191,N_7720,N_7762);
xor U8192 (N_8192,N_7483,N_7401);
and U8193 (N_8193,N_7511,N_7210);
xnor U8194 (N_8194,N_7282,N_7307);
nor U8195 (N_8195,N_7268,N_7454);
xnor U8196 (N_8196,N_7355,N_7384);
nor U8197 (N_8197,N_7446,N_7267);
xor U8198 (N_8198,N_7562,N_7291);
nand U8199 (N_8199,N_7643,N_7237);
xnor U8200 (N_8200,N_7641,N_7342);
nor U8201 (N_8201,N_7434,N_7371);
nand U8202 (N_8202,N_7440,N_7219);
nand U8203 (N_8203,N_7289,N_7688);
or U8204 (N_8204,N_7388,N_7316);
nor U8205 (N_8205,N_7428,N_7460);
or U8206 (N_8206,N_7644,N_7245);
and U8207 (N_8207,N_7261,N_7601);
nand U8208 (N_8208,N_7364,N_7422);
nand U8209 (N_8209,N_7436,N_7520);
or U8210 (N_8210,N_7631,N_7245);
or U8211 (N_8211,N_7743,N_7757);
nand U8212 (N_8212,N_7357,N_7365);
xnor U8213 (N_8213,N_7795,N_7474);
nand U8214 (N_8214,N_7491,N_7242);
nor U8215 (N_8215,N_7382,N_7539);
nor U8216 (N_8216,N_7337,N_7520);
or U8217 (N_8217,N_7620,N_7652);
xor U8218 (N_8218,N_7576,N_7603);
or U8219 (N_8219,N_7398,N_7320);
or U8220 (N_8220,N_7769,N_7335);
nand U8221 (N_8221,N_7676,N_7569);
nand U8222 (N_8222,N_7686,N_7308);
and U8223 (N_8223,N_7406,N_7370);
xnor U8224 (N_8224,N_7741,N_7773);
nor U8225 (N_8225,N_7655,N_7214);
nor U8226 (N_8226,N_7437,N_7713);
and U8227 (N_8227,N_7588,N_7759);
nor U8228 (N_8228,N_7696,N_7598);
and U8229 (N_8229,N_7310,N_7358);
and U8230 (N_8230,N_7437,N_7249);
and U8231 (N_8231,N_7731,N_7763);
xnor U8232 (N_8232,N_7650,N_7583);
and U8233 (N_8233,N_7553,N_7315);
or U8234 (N_8234,N_7615,N_7511);
nor U8235 (N_8235,N_7589,N_7268);
xor U8236 (N_8236,N_7790,N_7546);
nand U8237 (N_8237,N_7636,N_7724);
nand U8238 (N_8238,N_7243,N_7212);
nand U8239 (N_8239,N_7576,N_7542);
nor U8240 (N_8240,N_7217,N_7637);
and U8241 (N_8241,N_7695,N_7448);
nand U8242 (N_8242,N_7581,N_7304);
and U8243 (N_8243,N_7258,N_7437);
or U8244 (N_8244,N_7250,N_7398);
and U8245 (N_8245,N_7614,N_7317);
nand U8246 (N_8246,N_7554,N_7567);
or U8247 (N_8247,N_7672,N_7657);
xnor U8248 (N_8248,N_7281,N_7397);
nand U8249 (N_8249,N_7215,N_7428);
or U8250 (N_8250,N_7549,N_7535);
nand U8251 (N_8251,N_7391,N_7397);
nand U8252 (N_8252,N_7757,N_7303);
nand U8253 (N_8253,N_7671,N_7795);
nor U8254 (N_8254,N_7659,N_7363);
nand U8255 (N_8255,N_7630,N_7537);
nand U8256 (N_8256,N_7455,N_7725);
and U8257 (N_8257,N_7356,N_7641);
nand U8258 (N_8258,N_7283,N_7416);
xnor U8259 (N_8259,N_7296,N_7574);
nor U8260 (N_8260,N_7325,N_7396);
and U8261 (N_8261,N_7679,N_7585);
and U8262 (N_8262,N_7315,N_7296);
nor U8263 (N_8263,N_7426,N_7544);
and U8264 (N_8264,N_7709,N_7743);
or U8265 (N_8265,N_7288,N_7606);
nand U8266 (N_8266,N_7751,N_7777);
nand U8267 (N_8267,N_7580,N_7326);
or U8268 (N_8268,N_7624,N_7352);
xnor U8269 (N_8269,N_7420,N_7250);
and U8270 (N_8270,N_7303,N_7518);
or U8271 (N_8271,N_7567,N_7338);
nand U8272 (N_8272,N_7613,N_7314);
nor U8273 (N_8273,N_7701,N_7477);
nand U8274 (N_8274,N_7752,N_7223);
nand U8275 (N_8275,N_7313,N_7675);
nor U8276 (N_8276,N_7633,N_7414);
or U8277 (N_8277,N_7544,N_7521);
nand U8278 (N_8278,N_7526,N_7468);
or U8279 (N_8279,N_7650,N_7266);
or U8280 (N_8280,N_7519,N_7751);
xor U8281 (N_8281,N_7261,N_7233);
nor U8282 (N_8282,N_7738,N_7395);
xnor U8283 (N_8283,N_7482,N_7254);
xnor U8284 (N_8284,N_7570,N_7775);
nor U8285 (N_8285,N_7553,N_7236);
xnor U8286 (N_8286,N_7430,N_7545);
nand U8287 (N_8287,N_7603,N_7532);
nor U8288 (N_8288,N_7220,N_7600);
or U8289 (N_8289,N_7574,N_7482);
or U8290 (N_8290,N_7292,N_7228);
and U8291 (N_8291,N_7371,N_7454);
nor U8292 (N_8292,N_7357,N_7709);
and U8293 (N_8293,N_7366,N_7485);
nand U8294 (N_8294,N_7570,N_7341);
xnor U8295 (N_8295,N_7376,N_7402);
xor U8296 (N_8296,N_7570,N_7716);
nand U8297 (N_8297,N_7456,N_7479);
or U8298 (N_8298,N_7613,N_7476);
nor U8299 (N_8299,N_7735,N_7383);
and U8300 (N_8300,N_7630,N_7711);
nor U8301 (N_8301,N_7417,N_7484);
nor U8302 (N_8302,N_7395,N_7456);
xnor U8303 (N_8303,N_7408,N_7538);
and U8304 (N_8304,N_7438,N_7554);
and U8305 (N_8305,N_7288,N_7761);
or U8306 (N_8306,N_7383,N_7713);
xnor U8307 (N_8307,N_7406,N_7225);
nor U8308 (N_8308,N_7569,N_7404);
nor U8309 (N_8309,N_7293,N_7727);
nor U8310 (N_8310,N_7723,N_7261);
xor U8311 (N_8311,N_7346,N_7211);
nor U8312 (N_8312,N_7295,N_7696);
nor U8313 (N_8313,N_7501,N_7385);
and U8314 (N_8314,N_7468,N_7603);
xnor U8315 (N_8315,N_7612,N_7446);
and U8316 (N_8316,N_7373,N_7355);
or U8317 (N_8317,N_7439,N_7614);
or U8318 (N_8318,N_7389,N_7519);
xor U8319 (N_8319,N_7612,N_7746);
or U8320 (N_8320,N_7405,N_7594);
and U8321 (N_8321,N_7258,N_7669);
or U8322 (N_8322,N_7798,N_7403);
nand U8323 (N_8323,N_7454,N_7647);
and U8324 (N_8324,N_7325,N_7426);
nand U8325 (N_8325,N_7448,N_7411);
nor U8326 (N_8326,N_7230,N_7568);
nand U8327 (N_8327,N_7558,N_7402);
nand U8328 (N_8328,N_7758,N_7203);
xnor U8329 (N_8329,N_7756,N_7738);
xor U8330 (N_8330,N_7347,N_7653);
and U8331 (N_8331,N_7792,N_7536);
and U8332 (N_8332,N_7634,N_7397);
or U8333 (N_8333,N_7776,N_7794);
and U8334 (N_8334,N_7648,N_7713);
nor U8335 (N_8335,N_7719,N_7276);
xnor U8336 (N_8336,N_7300,N_7628);
or U8337 (N_8337,N_7388,N_7607);
xnor U8338 (N_8338,N_7768,N_7714);
xnor U8339 (N_8339,N_7342,N_7513);
nor U8340 (N_8340,N_7526,N_7461);
nor U8341 (N_8341,N_7608,N_7443);
or U8342 (N_8342,N_7447,N_7457);
or U8343 (N_8343,N_7321,N_7663);
and U8344 (N_8344,N_7410,N_7757);
nand U8345 (N_8345,N_7661,N_7501);
and U8346 (N_8346,N_7778,N_7575);
nor U8347 (N_8347,N_7410,N_7345);
and U8348 (N_8348,N_7645,N_7513);
xnor U8349 (N_8349,N_7312,N_7399);
nand U8350 (N_8350,N_7210,N_7543);
nor U8351 (N_8351,N_7397,N_7275);
nor U8352 (N_8352,N_7734,N_7326);
nand U8353 (N_8353,N_7586,N_7725);
nor U8354 (N_8354,N_7683,N_7599);
nor U8355 (N_8355,N_7762,N_7312);
or U8356 (N_8356,N_7433,N_7654);
nand U8357 (N_8357,N_7795,N_7581);
nor U8358 (N_8358,N_7693,N_7386);
nand U8359 (N_8359,N_7758,N_7750);
or U8360 (N_8360,N_7388,N_7510);
nand U8361 (N_8361,N_7204,N_7513);
or U8362 (N_8362,N_7536,N_7206);
and U8363 (N_8363,N_7584,N_7329);
nand U8364 (N_8364,N_7490,N_7424);
nor U8365 (N_8365,N_7671,N_7644);
xnor U8366 (N_8366,N_7440,N_7500);
xnor U8367 (N_8367,N_7623,N_7408);
or U8368 (N_8368,N_7440,N_7239);
or U8369 (N_8369,N_7390,N_7704);
nand U8370 (N_8370,N_7667,N_7405);
or U8371 (N_8371,N_7450,N_7549);
nand U8372 (N_8372,N_7381,N_7324);
and U8373 (N_8373,N_7700,N_7688);
nor U8374 (N_8374,N_7708,N_7312);
or U8375 (N_8375,N_7490,N_7367);
xor U8376 (N_8376,N_7744,N_7421);
xnor U8377 (N_8377,N_7281,N_7415);
nor U8378 (N_8378,N_7506,N_7372);
xnor U8379 (N_8379,N_7486,N_7450);
xnor U8380 (N_8380,N_7508,N_7317);
or U8381 (N_8381,N_7556,N_7644);
and U8382 (N_8382,N_7467,N_7667);
nand U8383 (N_8383,N_7520,N_7498);
xor U8384 (N_8384,N_7453,N_7345);
and U8385 (N_8385,N_7769,N_7483);
xnor U8386 (N_8386,N_7478,N_7315);
xnor U8387 (N_8387,N_7295,N_7359);
and U8388 (N_8388,N_7281,N_7525);
and U8389 (N_8389,N_7738,N_7654);
xnor U8390 (N_8390,N_7724,N_7240);
nor U8391 (N_8391,N_7745,N_7343);
nor U8392 (N_8392,N_7613,N_7406);
nand U8393 (N_8393,N_7522,N_7500);
xor U8394 (N_8394,N_7727,N_7788);
nand U8395 (N_8395,N_7377,N_7659);
nor U8396 (N_8396,N_7636,N_7331);
nor U8397 (N_8397,N_7748,N_7545);
or U8398 (N_8398,N_7494,N_7700);
nand U8399 (N_8399,N_7651,N_7482);
or U8400 (N_8400,N_8157,N_8070);
and U8401 (N_8401,N_8236,N_8101);
nand U8402 (N_8402,N_7813,N_8183);
xor U8403 (N_8403,N_7838,N_7989);
xor U8404 (N_8404,N_7879,N_7950);
xnor U8405 (N_8405,N_8340,N_8328);
xnor U8406 (N_8406,N_8282,N_7849);
and U8407 (N_8407,N_8300,N_8208);
or U8408 (N_8408,N_7916,N_8376);
xor U8409 (N_8409,N_8377,N_8167);
or U8410 (N_8410,N_8156,N_8017);
nor U8411 (N_8411,N_8230,N_7816);
or U8412 (N_8412,N_8108,N_7968);
nor U8413 (N_8413,N_7945,N_8105);
xnor U8414 (N_8414,N_7818,N_8139);
or U8415 (N_8415,N_7851,N_8096);
nand U8416 (N_8416,N_7856,N_8109);
nor U8417 (N_8417,N_8014,N_7943);
and U8418 (N_8418,N_7853,N_8241);
nand U8419 (N_8419,N_8333,N_8146);
nand U8420 (N_8420,N_7895,N_8052);
nand U8421 (N_8421,N_8055,N_8189);
xor U8422 (N_8422,N_7861,N_8242);
xor U8423 (N_8423,N_8291,N_7926);
nand U8424 (N_8424,N_7827,N_8152);
nor U8425 (N_8425,N_8395,N_8392);
nand U8426 (N_8426,N_8283,N_8325);
and U8427 (N_8427,N_8310,N_7868);
nor U8428 (N_8428,N_8323,N_8299);
and U8429 (N_8429,N_7899,N_8194);
nand U8430 (N_8430,N_8364,N_8324);
or U8431 (N_8431,N_8080,N_7886);
or U8432 (N_8432,N_8149,N_8011);
nand U8433 (N_8433,N_8046,N_7935);
and U8434 (N_8434,N_8073,N_8025);
or U8435 (N_8435,N_7932,N_8274);
or U8436 (N_8436,N_8125,N_7803);
nor U8437 (N_8437,N_8275,N_8272);
xnor U8438 (N_8438,N_8092,N_8042);
nand U8439 (N_8439,N_8319,N_8345);
and U8440 (N_8440,N_7985,N_8220);
xor U8441 (N_8441,N_8175,N_8172);
nor U8442 (N_8442,N_8393,N_7878);
or U8443 (N_8443,N_8278,N_8251);
nor U8444 (N_8444,N_8249,N_7801);
and U8445 (N_8445,N_8036,N_8214);
nor U8446 (N_8446,N_8027,N_8264);
xor U8447 (N_8447,N_7815,N_8204);
nor U8448 (N_8448,N_8169,N_8031);
nor U8449 (N_8449,N_8255,N_7930);
and U8450 (N_8450,N_8240,N_8084);
or U8451 (N_8451,N_8260,N_8018);
xor U8452 (N_8452,N_8131,N_8126);
xnor U8453 (N_8453,N_8159,N_8331);
nor U8454 (N_8454,N_8262,N_8099);
nand U8455 (N_8455,N_8396,N_8034);
nor U8456 (N_8456,N_7951,N_8062);
nand U8457 (N_8457,N_8045,N_7959);
xnor U8458 (N_8458,N_8199,N_8243);
xnor U8459 (N_8459,N_7890,N_8353);
nor U8460 (N_8460,N_8170,N_8254);
and U8461 (N_8461,N_7919,N_8357);
nand U8462 (N_8462,N_7971,N_8124);
xnor U8463 (N_8463,N_8305,N_7986);
xor U8464 (N_8464,N_7877,N_8234);
nor U8465 (N_8465,N_8112,N_7978);
xor U8466 (N_8466,N_8228,N_8206);
nor U8467 (N_8467,N_8344,N_8129);
nor U8468 (N_8468,N_8119,N_7914);
nor U8469 (N_8469,N_8285,N_8238);
xnor U8470 (N_8470,N_7947,N_8284);
nand U8471 (N_8471,N_8259,N_7921);
xor U8472 (N_8472,N_7896,N_7873);
nand U8473 (N_8473,N_8095,N_8226);
nand U8474 (N_8474,N_7824,N_8153);
xnor U8475 (N_8475,N_8193,N_8040);
and U8476 (N_8476,N_7979,N_7889);
nand U8477 (N_8477,N_7936,N_7942);
nor U8478 (N_8478,N_8181,N_7952);
or U8479 (N_8479,N_7810,N_7987);
or U8480 (N_8480,N_7966,N_8387);
and U8481 (N_8481,N_8104,N_7940);
and U8482 (N_8482,N_8212,N_8160);
nand U8483 (N_8483,N_8177,N_8269);
or U8484 (N_8484,N_8003,N_8338);
nor U8485 (N_8485,N_8192,N_8245);
and U8486 (N_8486,N_8120,N_8314);
nor U8487 (N_8487,N_8111,N_8320);
and U8488 (N_8488,N_7850,N_8021);
or U8489 (N_8489,N_8277,N_8075);
nor U8490 (N_8490,N_7912,N_8221);
nand U8491 (N_8491,N_8217,N_8135);
nor U8492 (N_8492,N_7997,N_8394);
xnor U8493 (N_8493,N_8163,N_8090);
nor U8494 (N_8494,N_8281,N_8134);
and U8495 (N_8495,N_8056,N_8168);
or U8496 (N_8496,N_7956,N_7931);
nand U8497 (N_8497,N_7867,N_8094);
nand U8498 (N_8498,N_7990,N_8267);
xor U8499 (N_8499,N_8133,N_7831);
nor U8500 (N_8500,N_8289,N_7880);
nor U8501 (N_8501,N_8022,N_8038);
nand U8502 (N_8502,N_8351,N_8037);
or U8503 (N_8503,N_7922,N_8235);
and U8504 (N_8504,N_8150,N_7905);
nor U8505 (N_8505,N_8128,N_7819);
nand U8506 (N_8506,N_7829,N_8142);
nand U8507 (N_8507,N_8178,N_8077);
and U8508 (N_8508,N_8297,N_8063);
nor U8509 (N_8509,N_8225,N_8127);
xnor U8510 (N_8510,N_7820,N_8363);
and U8511 (N_8511,N_8081,N_8020);
nand U8512 (N_8512,N_7929,N_7894);
nor U8513 (N_8513,N_8334,N_7939);
xor U8514 (N_8514,N_8078,N_7802);
nand U8515 (N_8515,N_8312,N_7884);
or U8516 (N_8516,N_7998,N_7907);
or U8517 (N_8517,N_8203,N_8008);
xnor U8518 (N_8518,N_8100,N_8360);
nand U8519 (N_8519,N_8082,N_7937);
nand U8520 (N_8520,N_7949,N_7812);
and U8521 (N_8521,N_8389,N_8019);
xnor U8522 (N_8522,N_7844,N_7839);
and U8523 (N_8523,N_8359,N_8304);
and U8524 (N_8524,N_7904,N_7814);
or U8525 (N_8525,N_7821,N_8143);
nand U8526 (N_8526,N_8064,N_7837);
and U8527 (N_8527,N_7876,N_7917);
nor U8528 (N_8528,N_7981,N_7903);
xor U8529 (N_8529,N_8270,N_8076);
and U8530 (N_8530,N_8085,N_8138);
or U8531 (N_8531,N_8044,N_8332);
or U8532 (N_8532,N_8051,N_7908);
nor U8533 (N_8533,N_7822,N_8263);
and U8534 (N_8534,N_8012,N_8370);
or U8535 (N_8535,N_8116,N_8329);
or U8536 (N_8536,N_8246,N_7836);
nor U8537 (N_8537,N_8313,N_8381);
xnor U8538 (N_8538,N_8294,N_7944);
nor U8539 (N_8539,N_8253,N_7869);
nor U8540 (N_8540,N_8180,N_7928);
nand U8541 (N_8541,N_8010,N_7954);
nor U8542 (N_8542,N_8301,N_8290);
nand U8543 (N_8543,N_8252,N_7855);
nand U8544 (N_8544,N_7900,N_8215);
xor U8545 (N_8545,N_7911,N_7883);
and U8546 (N_8546,N_8186,N_8107);
or U8547 (N_8547,N_8050,N_7892);
and U8548 (N_8548,N_8271,N_7885);
nand U8549 (N_8549,N_7965,N_8043);
and U8550 (N_8550,N_7924,N_8355);
xor U8551 (N_8551,N_8211,N_7962);
nand U8552 (N_8552,N_8088,N_7974);
xnor U8553 (N_8553,N_8117,N_8074);
nand U8554 (N_8554,N_8141,N_8071);
xor U8555 (N_8555,N_7994,N_7863);
xor U8556 (N_8556,N_8322,N_8026);
xnor U8557 (N_8557,N_8348,N_7955);
xor U8558 (N_8558,N_8144,N_8093);
and U8559 (N_8559,N_8342,N_8229);
nor U8560 (N_8560,N_8083,N_8059);
nand U8561 (N_8561,N_8326,N_7825);
and U8562 (N_8562,N_8231,N_7866);
nor U8563 (N_8563,N_8151,N_7857);
nand U8564 (N_8564,N_7860,N_8106);
or U8565 (N_8565,N_8369,N_8384);
nor U8566 (N_8566,N_7972,N_8047);
xnor U8567 (N_8567,N_7901,N_7913);
nand U8568 (N_8568,N_8379,N_7973);
or U8569 (N_8569,N_7870,N_8388);
nand U8570 (N_8570,N_8336,N_7842);
nand U8571 (N_8571,N_8158,N_8016);
or U8572 (N_8572,N_8197,N_7834);
or U8573 (N_8573,N_7817,N_8202);
nor U8574 (N_8574,N_8306,N_7871);
and U8575 (N_8575,N_8265,N_8239);
or U8576 (N_8576,N_7977,N_8182);
or U8577 (N_8577,N_8013,N_8200);
nand U8578 (N_8578,N_8001,N_8224);
xnor U8579 (N_8579,N_8161,N_8383);
xnor U8580 (N_8580,N_8009,N_7991);
or U8581 (N_8581,N_7845,N_8209);
xnor U8582 (N_8582,N_7961,N_8399);
nor U8583 (N_8583,N_7862,N_8247);
xnor U8584 (N_8584,N_7830,N_8347);
or U8585 (N_8585,N_8257,N_8205);
nand U8586 (N_8586,N_8223,N_7957);
or U8587 (N_8587,N_8198,N_8196);
nor U8588 (N_8588,N_8136,N_8123);
or U8589 (N_8589,N_8171,N_8176);
nand U8590 (N_8590,N_8187,N_8165);
nand U8591 (N_8591,N_8261,N_7888);
nand U8592 (N_8592,N_8232,N_7970);
xor U8593 (N_8593,N_8137,N_8250);
xor U8594 (N_8594,N_8179,N_7804);
or U8595 (N_8595,N_8362,N_8258);
nor U8596 (N_8596,N_8339,N_8057);
xnor U8597 (N_8597,N_7881,N_8091);
or U8598 (N_8598,N_8385,N_8352);
nor U8599 (N_8599,N_8216,N_8201);
nor U8600 (N_8600,N_7805,N_8110);
nor U8601 (N_8601,N_8308,N_8030);
xor U8602 (N_8602,N_8140,N_8188);
nand U8603 (N_8603,N_8041,N_8373);
and U8604 (N_8604,N_8061,N_7807);
nor U8605 (N_8605,N_7958,N_7902);
or U8606 (N_8606,N_8341,N_8007);
and U8607 (N_8607,N_8227,N_8173);
or U8608 (N_8608,N_7846,N_7933);
xnor U8609 (N_8609,N_8023,N_7847);
xor U8610 (N_8610,N_7946,N_8367);
nand U8611 (N_8611,N_8330,N_8321);
and U8612 (N_8612,N_7854,N_8327);
nand U8613 (N_8613,N_8317,N_8154);
and U8614 (N_8614,N_8122,N_8065);
nor U8615 (N_8615,N_8054,N_7843);
nor U8616 (N_8616,N_7828,N_7841);
nor U8617 (N_8617,N_8397,N_8248);
nor U8618 (N_8618,N_7923,N_8391);
xnor U8619 (N_8619,N_8296,N_8273);
and U8620 (N_8620,N_8287,N_8033);
or U8621 (N_8621,N_8293,N_7809);
xnor U8622 (N_8622,N_8166,N_8118);
or U8623 (N_8623,N_7858,N_8280);
or U8624 (N_8624,N_8184,N_8311);
nor U8625 (N_8625,N_7925,N_8002);
or U8626 (N_8626,N_8315,N_8102);
nor U8627 (N_8627,N_8130,N_7910);
and U8628 (N_8628,N_8114,N_7875);
nor U8629 (N_8629,N_8222,N_7865);
nand U8630 (N_8630,N_7975,N_8266);
nand U8631 (N_8631,N_8380,N_8368);
nor U8632 (N_8632,N_8268,N_8256);
nor U8633 (N_8633,N_8162,N_8365);
nand U8634 (N_8634,N_8115,N_8032);
nand U8635 (N_8635,N_8219,N_7941);
and U8636 (N_8636,N_8356,N_8349);
xnor U8637 (N_8637,N_7826,N_8148);
nor U8638 (N_8638,N_8210,N_7918);
nor U8639 (N_8639,N_8398,N_8279);
and U8640 (N_8640,N_8029,N_8087);
or U8641 (N_8641,N_8035,N_8098);
nor U8642 (N_8642,N_8079,N_7874);
xnor U8643 (N_8643,N_7835,N_8069);
and U8644 (N_8644,N_7920,N_7953);
xnor U8645 (N_8645,N_8086,N_8039);
nor U8646 (N_8646,N_7963,N_7964);
or U8647 (N_8647,N_8288,N_7927);
or U8648 (N_8648,N_7967,N_7808);
and U8649 (N_8649,N_8006,N_8207);
xor U8650 (N_8650,N_8354,N_8318);
and U8651 (N_8651,N_8185,N_8147);
or U8652 (N_8652,N_8372,N_8005);
nor U8653 (N_8653,N_8233,N_8058);
nor U8654 (N_8654,N_8164,N_7882);
nand U8655 (N_8655,N_8366,N_7995);
nand U8656 (N_8656,N_8303,N_8048);
nor U8657 (N_8657,N_7915,N_8295);
nor U8658 (N_8658,N_8072,N_8004);
nand U8659 (N_8659,N_8195,N_8068);
nor U8660 (N_8660,N_7893,N_7872);
nor U8661 (N_8661,N_8067,N_7898);
nand U8662 (N_8662,N_7984,N_8386);
nand U8663 (N_8663,N_7852,N_8309);
xor U8664 (N_8664,N_7811,N_8132);
or U8665 (N_8665,N_7983,N_7976);
or U8666 (N_8666,N_8015,N_8097);
xor U8667 (N_8667,N_8024,N_7934);
nand U8668 (N_8668,N_8382,N_8343);
nand U8669 (N_8669,N_8145,N_8374);
or U8670 (N_8670,N_8286,N_7992);
xor U8671 (N_8671,N_8066,N_7864);
and U8672 (N_8672,N_7891,N_8060);
and U8673 (N_8673,N_7960,N_8053);
nand U8674 (N_8674,N_7948,N_8191);
and U8675 (N_8675,N_7823,N_7988);
nor U8676 (N_8676,N_8335,N_8361);
and U8677 (N_8677,N_7999,N_7833);
nand U8678 (N_8678,N_7832,N_8378);
or U8679 (N_8679,N_8028,N_7800);
and U8680 (N_8680,N_7840,N_8390);
and U8681 (N_8681,N_8371,N_7909);
nand U8682 (N_8682,N_7859,N_8307);
and U8683 (N_8683,N_8358,N_7806);
or U8684 (N_8684,N_8346,N_7969);
and U8685 (N_8685,N_8350,N_8292);
or U8686 (N_8686,N_8244,N_7980);
nor U8687 (N_8687,N_7993,N_8089);
nand U8688 (N_8688,N_7996,N_8337);
xnor U8689 (N_8689,N_8302,N_8121);
xnor U8690 (N_8690,N_8375,N_8000);
or U8691 (N_8691,N_8113,N_8218);
nor U8692 (N_8692,N_7897,N_8276);
nand U8693 (N_8693,N_7887,N_7982);
nor U8694 (N_8694,N_8155,N_7848);
and U8695 (N_8695,N_8316,N_7906);
xnor U8696 (N_8696,N_8049,N_8174);
nand U8697 (N_8697,N_7938,N_8298);
and U8698 (N_8698,N_8190,N_8103);
and U8699 (N_8699,N_8213,N_8237);
nor U8700 (N_8700,N_8262,N_8125);
nand U8701 (N_8701,N_7993,N_8359);
or U8702 (N_8702,N_7962,N_8368);
xnor U8703 (N_8703,N_8229,N_8125);
and U8704 (N_8704,N_7924,N_8365);
nor U8705 (N_8705,N_8036,N_8090);
nor U8706 (N_8706,N_8179,N_8274);
nand U8707 (N_8707,N_8197,N_8180);
nand U8708 (N_8708,N_8191,N_8347);
nor U8709 (N_8709,N_8128,N_8172);
nor U8710 (N_8710,N_8133,N_8145);
xor U8711 (N_8711,N_8123,N_8243);
nand U8712 (N_8712,N_8330,N_8369);
and U8713 (N_8713,N_7838,N_7834);
nand U8714 (N_8714,N_8140,N_8032);
xor U8715 (N_8715,N_7896,N_8350);
nor U8716 (N_8716,N_7988,N_8324);
nand U8717 (N_8717,N_8385,N_8287);
or U8718 (N_8718,N_8291,N_7927);
or U8719 (N_8719,N_7912,N_7828);
or U8720 (N_8720,N_7898,N_8002);
xor U8721 (N_8721,N_7890,N_8202);
or U8722 (N_8722,N_8003,N_8261);
nand U8723 (N_8723,N_8301,N_8042);
and U8724 (N_8724,N_8195,N_7939);
nor U8725 (N_8725,N_8290,N_8175);
or U8726 (N_8726,N_8120,N_7861);
or U8727 (N_8727,N_7971,N_8170);
and U8728 (N_8728,N_8158,N_7803);
nor U8729 (N_8729,N_7892,N_8193);
or U8730 (N_8730,N_7985,N_8242);
nand U8731 (N_8731,N_8346,N_7869);
or U8732 (N_8732,N_7962,N_7865);
nor U8733 (N_8733,N_7937,N_7949);
and U8734 (N_8734,N_8380,N_8149);
xor U8735 (N_8735,N_7812,N_8083);
or U8736 (N_8736,N_8277,N_8127);
or U8737 (N_8737,N_8044,N_8282);
xor U8738 (N_8738,N_8167,N_8032);
xor U8739 (N_8739,N_8162,N_7876);
nor U8740 (N_8740,N_8032,N_8262);
xnor U8741 (N_8741,N_8292,N_8116);
nand U8742 (N_8742,N_8148,N_7813);
or U8743 (N_8743,N_8165,N_7919);
nor U8744 (N_8744,N_8100,N_7858);
and U8745 (N_8745,N_8336,N_7951);
or U8746 (N_8746,N_8093,N_7888);
xnor U8747 (N_8747,N_7998,N_8121);
nor U8748 (N_8748,N_8244,N_7964);
and U8749 (N_8749,N_7983,N_7867);
xor U8750 (N_8750,N_8295,N_8173);
or U8751 (N_8751,N_8087,N_8241);
and U8752 (N_8752,N_8064,N_7905);
xor U8753 (N_8753,N_7922,N_8029);
nor U8754 (N_8754,N_8288,N_8136);
xor U8755 (N_8755,N_8208,N_7901);
nor U8756 (N_8756,N_8217,N_7854);
xnor U8757 (N_8757,N_7871,N_7946);
xnor U8758 (N_8758,N_8381,N_8097);
and U8759 (N_8759,N_8351,N_8028);
and U8760 (N_8760,N_8195,N_8057);
xnor U8761 (N_8761,N_8128,N_8289);
or U8762 (N_8762,N_7881,N_8294);
nand U8763 (N_8763,N_8034,N_7933);
and U8764 (N_8764,N_8198,N_7830);
and U8765 (N_8765,N_8280,N_7954);
xnor U8766 (N_8766,N_7941,N_8316);
nor U8767 (N_8767,N_8211,N_7835);
and U8768 (N_8768,N_7996,N_8316);
or U8769 (N_8769,N_8353,N_8154);
nand U8770 (N_8770,N_7893,N_8200);
xor U8771 (N_8771,N_8174,N_7852);
nor U8772 (N_8772,N_8079,N_7936);
nand U8773 (N_8773,N_8050,N_7954);
nor U8774 (N_8774,N_8380,N_8359);
nor U8775 (N_8775,N_8121,N_7880);
xor U8776 (N_8776,N_8275,N_8327);
nor U8777 (N_8777,N_8386,N_7921);
or U8778 (N_8778,N_7937,N_7914);
xor U8779 (N_8779,N_8299,N_8147);
or U8780 (N_8780,N_7829,N_8107);
or U8781 (N_8781,N_8159,N_7887);
or U8782 (N_8782,N_8211,N_8340);
or U8783 (N_8783,N_8010,N_8002);
and U8784 (N_8784,N_8003,N_8216);
and U8785 (N_8785,N_8011,N_7989);
and U8786 (N_8786,N_8368,N_7913);
xnor U8787 (N_8787,N_7982,N_8227);
and U8788 (N_8788,N_8302,N_7898);
and U8789 (N_8789,N_8085,N_7869);
and U8790 (N_8790,N_8122,N_8079);
or U8791 (N_8791,N_7805,N_7847);
nand U8792 (N_8792,N_8308,N_7829);
or U8793 (N_8793,N_8144,N_8084);
or U8794 (N_8794,N_7925,N_8248);
or U8795 (N_8795,N_8282,N_8090);
and U8796 (N_8796,N_8364,N_7949);
and U8797 (N_8797,N_8064,N_8227);
nor U8798 (N_8798,N_8071,N_7973);
nor U8799 (N_8799,N_8120,N_8288);
and U8800 (N_8800,N_8314,N_8035);
xnor U8801 (N_8801,N_8124,N_8300);
nand U8802 (N_8802,N_8331,N_8211);
nor U8803 (N_8803,N_8175,N_8197);
xnor U8804 (N_8804,N_8242,N_8117);
nor U8805 (N_8805,N_7950,N_8038);
nor U8806 (N_8806,N_8080,N_8047);
or U8807 (N_8807,N_8307,N_7863);
or U8808 (N_8808,N_8105,N_8046);
xor U8809 (N_8809,N_8377,N_8325);
xor U8810 (N_8810,N_7859,N_8178);
xnor U8811 (N_8811,N_7956,N_8261);
or U8812 (N_8812,N_8171,N_8257);
nand U8813 (N_8813,N_8092,N_8318);
xor U8814 (N_8814,N_8370,N_8353);
xnor U8815 (N_8815,N_8365,N_8011);
nand U8816 (N_8816,N_8025,N_7915);
or U8817 (N_8817,N_7860,N_8092);
and U8818 (N_8818,N_8343,N_8296);
or U8819 (N_8819,N_7953,N_8209);
or U8820 (N_8820,N_8330,N_8161);
xnor U8821 (N_8821,N_8371,N_8353);
nor U8822 (N_8822,N_7997,N_8039);
xor U8823 (N_8823,N_8272,N_8280);
nor U8824 (N_8824,N_7942,N_8285);
or U8825 (N_8825,N_8264,N_8186);
nand U8826 (N_8826,N_8123,N_7943);
or U8827 (N_8827,N_7963,N_8209);
and U8828 (N_8828,N_8312,N_7865);
nor U8829 (N_8829,N_7859,N_8329);
or U8830 (N_8830,N_8042,N_7929);
nor U8831 (N_8831,N_8179,N_8018);
xor U8832 (N_8832,N_8325,N_7892);
nor U8833 (N_8833,N_7935,N_7909);
nor U8834 (N_8834,N_7838,N_7973);
or U8835 (N_8835,N_8045,N_8164);
nor U8836 (N_8836,N_7859,N_8089);
nand U8837 (N_8837,N_8359,N_8098);
nand U8838 (N_8838,N_7840,N_8118);
nand U8839 (N_8839,N_8173,N_8339);
or U8840 (N_8840,N_8072,N_7936);
xor U8841 (N_8841,N_7901,N_8131);
xor U8842 (N_8842,N_8101,N_8008);
xor U8843 (N_8843,N_8081,N_8174);
xor U8844 (N_8844,N_8190,N_8157);
nand U8845 (N_8845,N_7977,N_8300);
and U8846 (N_8846,N_7820,N_7888);
nand U8847 (N_8847,N_7807,N_7931);
or U8848 (N_8848,N_8328,N_8325);
xnor U8849 (N_8849,N_8208,N_7989);
nand U8850 (N_8850,N_7900,N_8006);
nor U8851 (N_8851,N_8054,N_8394);
or U8852 (N_8852,N_8175,N_7835);
nand U8853 (N_8853,N_8056,N_8088);
nor U8854 (N_8854,N_8113,N_8030);
nor U8855 (N_8855,N_7918,N_7823);
or U8856 (N_8856,N_7853,N_8389);
or U8857 (N_8857,N_7877,N_7823);
xor U8858 (N_8858,N_7930,N_8013);
nand U8859 (N_8859,N_8190,N_8112);
and U8860 (N_8860,N_8394,N_7880);
nand U8861 (N_8861,N_7883,N_8011);
nor U8862 (N_8862,N_7813,N_8308);
nor U8863 (N_8863,N_8289,N_7977);
or U8864 (N_8864,N_8292,N_8099);
or U8865 (N_8865,N_7811,N_8202);
nand U8866 (N_8866,N_7820,N_8373);
and U8867 (N_8867,N_8193,N_8276);
nand U8868 (N_8868,N_7939,N_7930);
or U8869 (N_8869,N_8335,N_8284);
and U8870 (N_8870,N_7844,N_8056);
or U8871 (N_8871,N_7991,N_8359);
nor U8872 (N_8872,N_8028,N_8029);
xnor U8873 (N_8873,N_7810,N_7890);
and U8874 (N_8874,N_7856,N_8352);
or U8875 (N_8875,N_8147,N_8199);
xnor U8876 (N_8876,N_7899,N_7980);
xor U8877 (N_8877,N_8322,N_8064);
and U8878 (N_8878,N_8340,N_8251);
nand U8879 (N_8879,N_8138,N_8102);
and U8880 (N_8880,N_8292,N_7861);
nand U8881 (N_8881,N_8182,N_8022);
xnor U8882 (N_8882,N_7968,N_8314);
nand U8883 (N_8883,N_8343,N_8380);
and U8884 (N_8884,N_7808,N_8194);
or U8885 (N_8885,N_7888,N_7808);
and U8886 (N_8886,N_8376,N_7871);
nand U8887 (N_8887,N_7969,N_8330);
nand U8888 (N_8888,N_7871,N_7992);
nor U8889 (N_8889,N_8394,N_7839);
or U8890 (N_8890,N_8394,N_8216);
nand U8891 (N_8891,N_7855,N_8064);
xor U8892 (N_8892,N_8039,N_8206);
nand U8893 (N_8893,N_8317,N_8327);
or U8894 (N_8894,N_8179,N_8375);
or U8895 (N_8895,N_7898,N_7960);
or U8896 (N_8896,N_7883,N_8277);
and U8897 (N_8897,N_7945,N_7867);
or U8898 (N_8898,N_8206,N_7871);
nand U8899 (N_8899,N_8276,N_8194);
and U8900 (N_8900,N_8287,N_8360);
xnor U8901 (N_8901,N_7857,N_8002);
nor U8902 (N_8902,N_7906,N_7803);
nor U8903 (N_8903,N_7842,N_7878);
nor U8904 (N_8904,N_7986,N_8332);
nand U8905 (N_8905,N_8372,N_7881);
nor U8906 (N_8906,N_7886,N_8182);
xor U8907 (N_8907,N_8215,N_8158);
or U8908 (N_8908,N_8088,N_8142);
xor U8909 (N_8909,N_8348,N_8178);
nor U8910 (N_8910,N_8054,N_8300);
and U8911 (N_8911,N_7998,N_8069);
xor U8912 (N_8912,N_8097,N_8338);
or U8913 (N_8913,N_8337,N_7884);
nor U8914 (N_8914,N_7835,N_8396);
nand U8915 (N_8915,N_8048,N_7990);
and U8916 (N_8916,N_8072,N_8101);
xor U8917 (N_8917,N_8266,N_8079);
or U8918 (N_8918,N_8241,N_7912);
or U8919 (N_8919,N_7960,N_7857);
and U8920 (N_8920,N_8369,N_8087);
or U8921 (N_8921,N_8327,N_8120);
nor U8922 (N_8922,N_8089,N_7847);
xnor U8923 (N_8923,N_7895,N_8270);
nor U8924 (N_8924,N_8044,N_8325);
nand U8925 (N_8925,N_8230,N_7931);
and U8926 (N_8926,N_8099,N_8055);
or U8927 (N_8927,N_7850,N_8308);
nor U8928 (N_8928,N_8030,N_7829);
and U8929 (N_8929,N_8398,N_7830);
nor U8930 (N_8930,N_8158,N_8147);
or U8931 (N_8931,N_7830,N_7880);
nor U8932 (N_8932,N_8230,N_8332);
or U8933 (N_8933,N_8320,N_8327);
nand U8934 (N_8934,N_7932,N_8355);
and U8935 (N_8935,N_8354,N_8187);
xor U8936 (N_8936,N_8137,N_8246);
nor U8937 (N_8937,N_8211,N_7982);
nand U8938 (N_8938,N_8394,N_8254);
and U8939 (N_8939,N_7827,N_7896);
nor U8940 (N_8940,N_7832,N_8248);
nand U8941 (N_8941,N_8399,N_7917);
and U8942 (N_8942,N_7929,N_8291);
nand U8943 (N_8943,N_7991,N_7826);
nand U8944 (N_8944,N_7953,N_7840);
or U8945 (N_8945,N_7903,N_7921);
nand U8946 (N_8946,N_8344,N_7953);
or U8947 (N_8947,N_8365,N_8299);
and U8948 (N_8948,N_8342,N_7997);
nand U8949 (N_8949,N_8040,N_7826);
and U8950 (N_8950,N_8331,N_8376);
nor U8951 (N_8951,N_7806,N_8335);
or U8952 (N_8952,N_8361,N_8329);
xor U8953 (N_8953,N_7802,N_7846);
and U8954 (N_8954,N_7807,N_8295);
xnor U8955 (N_8955,N_7970,N_8200);
nand U8956 (N_8956,N_7957,N_8022);
and U8957 (N_8957,N_7959,N_8081);
and U8958 (N_8958,N_8196,N_8013);
nand U8959 (N_8959,N_8358,N_7902);
nand U8960 (N_8960,N_7965,N_7959);
xor U8961 (N_8961,N_7949,N_7954);
xor U8962 (N_8962,N_7825,N_8315);
nand U8963 (N_8963,N_8350,N_8172);
nand U8964 (N_8964,N_8209,N_8301);
nand U8965 (N_8965,N_8237,N_8371);
nand U8966 (N_8966,N_8289,N_8041);
nand U8967 (N_8967,N_8164,N_8036);
or U8968 (N_8968,N_7810,N_8169);
xor U8969 (N_8969,N_8336,N_8183);
or U8970 (N_8970,N_8003,N_8013);
and U8971 (N_8971,N_8321,N_8090);
and U8972 (N_8972,N_7888,N_7914);
nor U8973 (N_8973,N_7810,N_8323);
nor U8974 (N_8974,N_8326,N_7873);
and U8975 (N_8975,N_8169,N_7921);
xor U8976 (N_8976,N_8142,N_7923);
and U8977 (N_8977,N_7954,N_8276);
xnor U8978 (N_8978,N_8179,N_8047);
xnor U8979 (N_8979,N_8027,N_8325);
xor U8980 (N_8980,N_8284,N_7872);
and U8981 (N_8981,N_8166,N_8140);
nand U8982 (N_8982,N_8073,N_8159);
xnor U8983 (N_8983,N_7811,N_8092);
nor U8984 (N_8984,N_8312,N_7936);
xor U8985 (N_8985,N_8077,N_8273);
nand U8986 (N_8986,N_8248,N_8338);
or U8987 (N_8987,N_7958,N_7957);
nor U8988 (N_8988,N_8273,N_8067);
xor U8989 (N_8989,N_8105,N_7956);
and U8990 (N_8990,N_8077,N_8316);
nor U8991 (N_8991,N_8242,N_8060);
or U8992 (N_8992,N_7810,N_8391);
and U8993 (N_8993,N_8163,N_8358);
nor U8994 (N_8994,N_7922,N_8052);
nor U8995 (N_8995,N_8030,N_8028);
nand U8996 (N_8996,N_7854,N_7844);
or U8997 (N_8997,N_8194,N_7994);
and U8998 (N_8998,N_8203,N_8319);
or U8999 (N_8999,N_8325,N_8294);
or U9000 (N_9000,N_8887,N_8824);
or U9001 (N_9001,N_8822,N_8919);
xor U9002 (N_9002,N_8871,N_8811);
nand U9003 (N_9003,N_8609,N_8860);
xnor U9004 (N_9004,N_8830,N_8627);
or U9005 (N_9005,N_8633,N_8743);
xor U9006 (N_9006,N_8455,N_8404);
nand U9007 (N_9007,N_8996,N_8877);
and U9008 (N_9008,N_8915,N_8695);
xor U9009 (N_9009,N_8835,N_8604);
nand U9010 (N_9010,N_8848,N_8571);
nor U9011 (N_9011,N_8726,N_8599);
xor U9012 (N_9012,N_8753,N_8967);
nor U9013 (N_9013,N_8954,N_8817);
and U9014 (N_9014,N_8629,N_8761);
or U9015 (N_9015,N_8456,N_8563);
or U9016 (N_9016,N_8809,N_8662);
xor U9017 (N_9017,N_8494,N_8555);
nand U9018 (N_9018,N_8833,N_8600);
and U9019 (N_9019,N_8984,N_8828);
nor U9020 (N_9020,N_8713,N_8696);
and U9021 (N_9021,N_8978,N_8553);
nand U9022 (N_9022,N_8861,N_8651);
and U9023 (N_9023,N_8565,N_8714);
or U9024 (N_9024,N_8927,N_8794);
or U9025 (N_9025,N_8656,N_8453);
nand U9026 (N_9026,N_8950,N_8879);
nand U9027 (N_9027,N_8905,N_8483);
nor U9028 (N_9028,N_8853,N_8434);
or U9029 (N_9029,N_8839,N_8519);
nor U9030 (N_9030,N_8963,N_8735);
nand U9031 (N_9031,N_8500,N_8411);
xor U9032 (N_9032,N_8512,N_8574);
or U9033 (N_9033,N_8851,N_8469);
nor U9034 (N_9034,N_8829,N_8891);
or U9035 (N_9035,N_8660,N_8790);
and U9036 (N_9036,N_8744,N_8748);
and U9037 (N_9037,N_8682,N_8678);
nor U9038 (N_9038,N_8890,N_8466);
nor U9039 (N_9039,N_8872,N_8614);
nor U9040 (N_9040,N_8775,N_8424);
nor U9041 (N_9041,N_8441,N_8987);
and U9042 (N_9042,N_8994,N_8777);
nand U9043 (N_9043,N_8725,N_8903);
nand U9044 (N_9044,N_8670,N_8489);
nand U9045 (N_9045,N_8669,N_8935);
nand U9046 (N_9046,N_8737,N_8405);
xor U9047 (N_9047,N_8586,N_8698);
or U9048 (N_9048,N_8492,N_8918);
or U9049 (N_9049,N_8475,N_8542);
nand U9050 (N_9050,N_8827,N_8896);
and U9051 (N_9051,N_8423,N_8868);
or U9052 (N_9052,N_8813,N_8899);
and U9053 (N_9053,N_8533,N_8977);
and U9054 (N_9054,N_8831,N_8438);
xnor U9055 (N_9055,N_8610,N_8823);
nand U9056 (N_9056,N_8976,N_8981);
and U9057 (N_9057,N_8941,N_8757);
and U9058 (N_9058,N_8582,N_8747);
nor U9059 (N_9059,N_8807,N_8968);
nor U9060 (N_9060,N_8874,N_8920);
nand U9061 (N_9061,N_8888,N_8457);
and U9062 (N_9062,N_8523,N_8755);
or U9063 (N_9063,N_8878,N_8815);
nand U9064 (N_9064,N_8717,N_8841);
nor U9065 (N_9065,N_8547,N_8646);
nand U9066 (N_9066,N_8679,N_8573);
nand U9067 (N_9067,N_8693,N_8739);
or U9068 (N_9068,N_8955,N_8847);
and U9069 (N_9069,N_8762,N_8842);
nor U9070 (N_9070,N_8710,N_8495);
nand U9071 (N_9071,N_8689,N_8487);
xnor U9072 (N_9072,N_8583,N_8703);
nor U9073 (N_9073,N_8718,N_8538);
nor U9074 (N_9074,N_8485,N_8606);
nor U9075 (N_9075,N_8562,N_8499);
xnor U9076 (N_9076,N_8673,N_8889);
nand U9077 (N_9077,N_8684,N_8998);
nand U9078 (N_9078,N_8722,N_8468);
and U9079 (N_9079,N_8638,N_8699);
nand U9080 (N_9080,N_8576,N_8417);
xor U9081 (N_9081,N_8951,N_8778);
xnor U9082 (N_9082,N_8785,N_8467);
nor U9083 (N_9083,N_8581,N_8862);
nor U9084 (N_9084,N_8480,N_8578);
nand U9085 (N_9085,N_8621,N_8593);
and U9086 (N_9086,N_8838,N_8639);
nand U9087 (N_9087,N_8972,N_8625);
nor U9088 (N_9088,N_8849,N_8789);
nor U9089 (N_9089,N_8979,N_8892);
xor U9090 (N_9090,N_8788,N_8766);
nand U9091 (N_9091,N_8588,N_8858);
or U9092 (N_9092,N_8772,N_8429);
or U9093 (N_9093,N_8445,N_8866);
nand U9094 (N_9094,N_8465,N_8448);
or U9095 (N_9095,N_8731,N_8685);
nor U9096 (N_9096,N_8402,N_8647);
nor U9097 (N_9097,N_8940,N_8926);
and U9098 (N_9098,N_8784,N_8650);
xnor U9099 (N_9099,N_8936,N_8530);
or U9100 (N_9100,N_8432,N_8746);
or U9101 (N_9101,N_8708,N_8661);
and U9102 (N_9102,N_8900,N_8444);
nand U9103 (N_9103,N_8765,N_8724);
nand U9104 (N_9104,N_8461,N_8464);
nand U9105 (N_9105,N_8974,N_8933);
nor U9106 (N_9106,N_8907,N_8534);
nand U9107 (N_9107,N_8886,N_8760);
nand U9108 (N_9108,N_8750,N_8721);
nand U9109 (N_9109,N_8914,N_8846);
nand U9110 (N_9110,N_8529,N_8601);
xor U9111 (N_9111,N_8518,N_8836);
xor U9112 (N_9112,N_8692,N_8628);
or U9113 (N_9113,N_8814,N_8473);
or U9114 (N_9114,N_8431,N_8999);
or U9115 (N_9115,N_8754,N_8472);
nand U9116 (N_9116,N_8452,N_8497);
xor U9117 (N_9117,N_8439,N_8507);
or U9118 (N_9118,N_8677,N_8501);
nand U9119 (N_9119,N_8742,N_8420);
or U9120 (N_9120,N_8644,N_8554);
or U9121 (N_9121,N_8882,N_8592);
and U9122 (N_9122,N_8732,N_8636);
and U9123 (N_9123,N_8667,N_8594);
nor U9124 (N_9124,N_8482,N_8970);
or U9125 (N_9125,N_8973,N_8910);
and U9126 (N_9126,N_8883,N_8447);
or U9127 (N_9127,N_8934,N_8613);
nor U9128 (N_9128,N_8840,N_8597);
nor U9129 (N_9129,N_8821,N_8983);
nor U9130 (N_9130,N_8570,N_8442);
nand U9131 (N_9131,N_8427,N_8412);
and U9132 (N_9132,N_8819,N_8770);
xnor U9133 (N_9133,N_8937,N_8885);
and U9134 (N_9134,N_8691,N_8577);
and U9135 (N_9135,N_8605,N_8906);
or U9136 (N_9136,N_8738,N_8705);
xnor U9137 (N_9137,N_8930,N_8478);
nor U9138 (N_9138,N_8720,N_8749);
xnor U9139 (N_9139,N_8686,N_8558);
nand U9140 (N_9140,N_8802,N_8654);
nand U9141 (N_9141,N_8645,N_8490);
or U9142 (N_9142,N_8990,N_8537);
or U9143 (N_9143,N_8969,N_8481);
xor U9144 (N_9144,N_8635,N_8881);
xnor U9145 (N_9145,N_8652,N_8917);
nor U9146 (N_9146,N_8855,N_8741);
nor U9147 (N_9147,N_8707,N_8414);
nor U9148 (N_9148,N_8857,N_8532);
nor U9149 (N_9149,N_8630,N_8929);
nand U9150 (N_9150,N_8767,N_8723);
and U9151 (N_9151,N_8818,N_8702);
nor U9152 (N_9152,N_8992,N_8806);
nand U9153 (N_9153,N_8779,N_8585);
and U9154 (N_9154,N_8908,N_8763);
and U9155 (N_9155,N_8869,N_8734);
and U9156 (N_9156,N_8843,N_8663);
and U9157 (N_9157,N_8911,N_8607);
xnor U9158 (N_9158,N_8460,N_8719);
or U9159 (N_9159,N_8709,N_8854);
nor U9160 (N_9160,N_8774,N_8956);
nand U9161 (N_9161,N_8852,N_8596);
xnor U9162 (N_9162,N_8561,N_8488);
nor U9163 (N_9163,N_8510,N_8572);
or U9164 (N_9164,N_8948,N_8557);
and U9165 (N_9165,N_8975,N_8611);
and U9166 (N_9166,N_8535,N_8664);
nor U9167 (N_9167,N_8642,N_8711);
and U9168 (N_9168,N_8904,N_8640);
and U9169 (N_9169,N_8844,N_8520);
nand U9170 (N_9170,N_8704,N_8801);
nand U9171 (N_9171,N_8493,N_8524);
nor U9172 (N_9172,N_8419,N_8945);
nor U9173 (N_9173,N_8608,N_8780);
xor U9174 (N_9174,N_8961,N_8567);
nand U9175 (N_9175,N_8437,N_8623);
nand U9176 (N_9176,N_8550,N_8958);
or U9177 (N_9177,N_8856,N_8820);
or U9178 (N_9178,N_8971,N_8873);
or U9179 (N_9179,N_8944,N_8740);
or U9180 (N_9180,N_8952,N_8957);
nor U9181 (N_9181,N_8546,N_8845);
and U9182 (N_9182,N_8422,N_8932);
nor U9183 (N_9183,N_8808,N_8913);
or U9184 (N_9184,N_8566,N_8752);
nand U9185 (N_9185,N_8459,N_8579);
nand U9186 (N_9186,N_8834,N_8458);
and U9187 (N_9187,N_8643,N_8690);
xor U9188 (N_9188,N_8997,N_8986);
nor U9189 (N_9189,N_8867,N_8786);
nand U9190 (N_9190,N_8922,N_8618);
xor U9191 (N_9191,N_8800,N_8421);
nand U9192 (N_9192,N_8825,N_8504);
nand U9193 (N_9193,N_8942,N_8924);
or U9194 (N_9194,N_8476,N_8470);
and U9195 (N_9195,N_8568,N_8751);
nor U9196 (N_9196,N_8960,N_8527);
nor U9197 (N_9197,N_8508,N_8666);
nor U9198 (N_9198,N_8884,N_8551);
nor U9199 (N_9199,N_8587,N_8773);
nand U9200 (N_9200,N_8706,N_8416);
xor U9201 (N_9201,N_8536,N_8985);
nand U9202 (N_9202,N_8528,N_8634);
nor U9203 (N_9203,N_8659,N_8521);
nand U9204 (N_9204,N_8559,N_8804);
nor U9205 (N_9205,N_8671,N_8943);
nand U9206 (N_9206,N_8649,N_8850);
nor U9207 (N_9207,N_8436,N_8474);
or U9208 (N_9208,N_8989,N_8771);
xor U9209 (N_9209,N_8805,N_8712);
xor U9210 (N_9210,N_8543,N_8701);
xnor U9211 (N_9211,N_8540,N_8632);
xor U9212 (N_9212,N_8443,N_8728);
nand U9213 (N_9213,N_8575,N_8966);
xnor U9214 (N_9214,N_8876,N_8622);
nand U9215 (N_9215,N_8672,N_8515);
or U9216 (N_9216,N_8631,N_8864);
or U9217 (N_9217,N_8946,N_8991);
and U9218 (N_9218,N_8406,N_8988);
and U9219 (N_9219,N_8511,N_8893);
nor U9220 (N_9220,N_8418,N_8683);
xnor U9221 (N_9221,N_8513,N_8727);
or U9222 (N_9222,N_8736,N_8923);
nand U9223 (N_9223,N_8595,N_8502);
nand U9224 (N_9224,N_8616,N_8484);
xor U9225 (N_9225,N_8653,N_8451);
xnor U9226 (N_9226,N_8916,N_8939);
or U9227 (N_9227,N_8798,N_8556);
nor U9228 (N_9228,N_8791,N_8584);
nand U9229 (N_9229,N_8598,N_8928);
nand U9230 (N_9230,N_8938,N_8810);
or U9231 (N_9231,N_8496,N_8962);
nor U9232 (N_9232,N_8863,N_8549);
nand U9233 (N_9233,N_8674,N_8545);
xor U9234 (N_9234,N_8425,N_8799);
and U9235 (N_9235,N_8641,N_8668);
nand U9236 (N_9236,N_8446,N_8995);
or U9237 (N_9237,N_8463,N_8400);
nor U9238 (N_9238,N_8875,N_8506);
and U9239 (N_9239,N_8912,N_8716);
and U9240 (N_9240,N_8517,N_8953);
nor U9241 (N_9241,N_8894,N_8655);
or U9242 (N_9242,N_8745,N_8965);
and U9243 (N_9243,N_8898,N_8797);
nand U9244 (N_9244,N_8479,N_8759);
nor U9245 (N_9245,N_8787,N_8803);
or U9246 (N_9246,N_8964,N_8832);
nor U9247 (N_9247,N_8730,N_8694);
nand U9248 (N_9248,N_8491,N_8590);
or U9249 (N_9249,N_8902,N_8688);
and U9250 (N_9250,N_8617,N_8925);
nor U9251 (N_9251,N_8548,N_8410);
and U9252 (N_9252,N_8681,N_8993);
nand U9253 (N_9253,N_8407,N_8783);
nor U9254 (N_9254,N_8769,N_8580);
nor U9255 (N_9255,N_8676,N_8837);
and U9256 (N_9256,N_8826,N_8782);
nor U9257 (N_9257,N_8462,N_8413);
xnor U9258 (N_9258,N_8525,N_8615);
and U9259 (N_9259,N_8509,N_8796);
nand U9260 (N_9260,N_8870,N_8931);
or U9261 (N_9261,N_8865,N_8776);
nand U9262 (N_9262,N_8959,N_8697);
nand U9263 (N_9263,N_8526,N_8816);
nor U9264 (N_9264,N_8700,N_8792);
and U9265 (N_9265,N_8665,N_8560);
and U9266 (N_9266,N_8505,N_8901);
xor U9267 (N_9267,N_8612,N_8603);
xor U9268 (N_9268,N_8569,N_8450);
and U9269 (N_9269,N_8729,N_8675);
xor U9270 (N_9270,N_8658,N_8909);
nor U9271 (N_9271,N_8471,N_8503);
xnor U9272 (N_9272,N_8949,N_8620);
nor U9273 (N_9273,N_8433,N_8680);
nand U9274 (N_9274,N_8758,N_8648);
or U9275 (N_9275,N_8531,N_8921);
or U9276 (N_9276,N_8687,N_8793);
nor U9277 (N_9277,N_8426,N_8880);
nor U9278 (N_9278,N_8539,N_8795);
nand U9279 (N_9279,N_8401,N_8764);
or U9280 (N_9280,N_8449,N_8514);
and U9281 (N_9281,N_8781,N_8715);
nor U9282 (N_9282,N_8768,N_8947);
xnor U9283 (N_9283,N_8516,N_8982);
and U9284 (N_9284,N_8409,N_8756);
nor U9285 (N_9285,N_8415,N_8980);
or U9286 (N_9286,N_8602,N_8552);
and U9287 (N_9287,N_8544,N_8541);
or U9288 (N_9288,N_8486,N_8626);
nand U9289 (N_9289,N_8522,N_8498);
nand U9290 (N_9290,N_8454,N_8589);
xor U9291 (N_9291,N_8733,N_8897);
or U9292 (N_9292,N_8435,N_8440);
nor U9293 (N_9293,N_8430,N_8591);
nand U9294 (N_9294,N_8637,N_8657);
nor U9295 (N_9295,N_8564,N_8619);
nor U9296 (N_9296,N_8408,N_8859);
xor U9297 (N_9297,N_8624,N_8477);
or U9298 (N_9298,N_8403,N_8895);
nand U9299 (N_9299,N_8428,N_8812);
and U9300 (N_9300,N_8821,N_8844);
or U9301 (N_9301,N_8942,N_8670);
and U9302 (N_9302,N_8757,N_8722);
nand U9303 (N_9303,N_8539,N_8932);
xnor U9304 (N_9304,N_8651,N_8795);
nor U9305 (N_9305,N_8494,N_8449);
nand U9306 (N_9306,N_8968,N_8735);
xnor U9307 (N_9307,N_8732,N_8879);
xor U9308 (N_9308,N_8449,N_8597);
and U9309 (N_9309,N_8731,N_8493);
nor U9310 (N_9310,N_8527,N_8833);
xor U9311 (N_9311,N_8968,N_8729);
or U9312 (N_9312,N_8459,N_8735);
and U9313 (N_9313,N_8810,N_8852);
nand U9314 (N_9314,N_8789,N_8416);
nand U9315 (N_9315,N_8427,N_8752);
xor U9316 (N_9316,N_8566,N_8471);
nand U9317 (N_9317,N_8449,N_8999);
xor U9318 (N_9318,N_8641,N_8630);
or U9319 (N_9319,N_8522,N_8566);
or U9320 (N_9320,N_8610,N_8622);
xor U9321 (N_9321,N_8537,N_8630);
xor U9322 (N_9322,N_8792,N_8912);
nand U9323 (N_9323,N_8873,N_8455);
and U9324 (N_9324,N_8865,N_8563);
xnor U9325 (N_9325,N_8519,N_8760);
and U9326 (N_9326,N_8663,N_8617);
or U9327 (N_9327,N_8426,N_8815);
xnor U9328 (N_9328,N_8703,N_8424);
nor U9329 (N_9329,N_8607,N_8855);
nor U9330 (N_9330,N_8483,N_8639);
nand U9331 (N_9331,N_8933,N_8868);
and U9332 (N_9332,N_8675,N_8432);
xnor U9333 (N_9333,N_8645,N_8911);
and U9334 (N_9334,N_8573,N_8947);
nor U9335 (N_9335,N_8605,N_8955);
or U9336 (N_9336,N_8895,N_8987);
or U9337 (N_9337,N_8758,N_8452);
nor U9338 (N_9338,N_8400,N_8525);
and U9339 (N_9339,N_8989,N_8533);
and U9340 (N_9340,N_8899,N_8972);
nor U9341 (N_9341,N_8855,N_8903);
and U9342 (N_9342,N_8577,N_8933);
nand U9343 (N_9343,N_8472,N_8685);
and U9344 (N_9344,N_8844,N_8513);
xnor U9345 (N_9345,N_8669,N_8558);
and U9346 (N_9346,N_8619,N_8707);
and U9347 (N_9347,N_8563,N_8547);
nor U9348 (N_9348,N_8765,N_8469);
nor U9349 (N_9349,N_8478,N_8815);
xnor U9350 (N_9350,N_8786,N_8609);
nor U9351 (N_9351,N_8927,N_8810);
nand U9352 (N_9352,N_8415,N_8889);
or U9353 (N_9353,N_8817,N_8862);
or U9354 (N_9354,N_8690,N_8448);
nand U9355 (N_9355,N_8708,N_8621);
nand U9356 (N_9356,N_8943,N_8967);
or U9357 (N_9357,N_8915,N_8952);
nand U9358 (N_9358,N_8612,N_8785);
or U9359 (N_9359,N_8930,N_8450);
or U9360 (N_9360,N_8422,N_8938);
nand U9361 (N_9361,N_8752,N_8429);
and U9362 (N_9362,N_8610,N_8718);
xnor U9363 (N_9363,N_8909,N_8619);
and U9364 (N_9364,N_8423,N_8503);
nand U9365 (N_9365,N_8728,N_8893);
and U9366 (N_9366,N_8753,N_8808);
and U9367 (N_9367,N_8993,N_8633);
nor U9368 (N_9368,N_8447,N_8966);
nor U9369 (N_9369,N_8464,N_8774);
and U9370 (N_9370,N_8655,N_8839);
xnor U9371 (N_9371,N_8925,N_8464);
nand U9372 (N_9372,N_8821,N_8817);
nor U9373 (N_9373,N_8540,N_8526);
xnor U9374 (N_9374,N_8831,N_8440);
xnor U9375 (N_9375,N_8711,N_8899);
xor U9376 (N_9376,N_8957,N_8627);
nor U9377 (N_9377,N_8950,N_8491);
nor U9378 (N_9378,N_8798,N_8843);
nand U9379 (N_9379,N_8678,N_8629);
xnor U9380 (N_9380,N_8789,N_8659);
nor U9381 (N_9381,N_8464,N_8937);
or U9382 (N_9382,N_8773,N_8670);
and U9383 (N_9383,N_8585,N_8991);
nand U9384 (N_9384,N_8404,N_8615);
and U9385 (N_9385,N_8473,N_8848);
and U9386 (N_9386,N_8714,N_8682);
xor U9387 (N_9387,N_8694,N_8474);
nand U9388 (N_9388,N_8426,N_8525);
and U9389 (N_9389,N_8876,N_8475);
nand U9390 (N_9390,N_8955,N_8519);
xor U9391 (N_9391,N_8686,N_8642);
nor U9392 (N_9392,N_8995,N_8965);
xor U9393 (N_9393,N_8624,N_8740);
nand U9394 (N_9394,N_8783,N_8707);
xor U9395 (N_9395,N_8485,N_8869);
xor U9396 (N_9396,N_8520,N_8555);
xor U9397 (N_9397,N_8529,N_8656);
nor U9398 (N_9398,N_8462,N_8810);
or U9399 (N_9399,N_8700,N_8781);
xnor U9400 (N_9400,N_8925,N_8493);
or U9401 (N_9401,N_8830,N_8785);
and U9402 (N_9402,N_8719,N_8851);
xnor U9403 (N_9403,N_8541,N_8493);
or U9404 (N_9404,N_8818,N_8925);
or U9405 (N_9405,N_8600,N_8764);
or U9406 (N_9406,N_8794,N_8896);
xor U9407 (N_9407,N_8831,N_8819);
and U9408 (N_9408,N_8711,N_8493);
nand U9409 (N_9409,N_8792,N_8518);
and U9410 (N_9410,N_8617,N_8692);
or U9411 (N_9411,N_8846,N_8621);
and U9412 (N_9412,N_8728,N_8645);
xnor U9413 (N_9413,N_8738,N_8443);
nor U9414 (N_9414,N_8766,N_8512);
or U9415 (N_9415,N_8696,N_8458);
nand U9416 (N_9416,N_8604,N_8595);
nor U9417 (N_9417,N_8854,N_8942);
nor U9418 (N_9418,N_8690,N_8478);
or U9419 (N_9419,N_8884,N_8715);
and U9420 (N_9420,N_8979,N_8573);
nor U9421 (N_9421,N_8755,N_8851);
xnor U9422 (N_9422,N_8438,N_8738);
nor U9423 (N_9423,N_8521,N_8431);
and U9424 (N_9424,N_8762,N_8953);
xor U9425 (N_9425,N_8678,N_8686);
or U9426 (N_9426,N_8974,N_8873);
nor U9427 (N_9427,N_8495,N_8867);
xor U9428 (N_9428,N_8720,N_8854);
xor U9429 (N_9429,N_8812,N_8929);
nor U9430 (N_9430,N_8969,N_8644);
or U9431 (N_9431,N_8495,N_8441);
nand U9432 (N_9432,N_8443,N_8827);
xor U9433 (N_9433,N_8626,N_8714);
xor U9434 (N_9434,N_8800,N_8444);
xnor U9435 (N_9435,N_8759,N_8426);
or U9436 (N_9436,N_8659,N_8463);
xor U9437 (N_9437,N_8400,N_8567);
nor U9438 (N_9438,N_8733,N_8993);
and U9439 (N_9439,N_8811,N_8781);
nor U9440 (N_9440,N_8969,N_8734);
xnor U9441 (N_9441,N_8431,N_8544);
or U9442 (N_9442,N_8426,N_8508);
nand U9443 (N_9443,N_8623,N_8551);
nor U9444 (N_9444,N_8902,N_8674);
nor U9445 (N_9445,N_8728,N_8491);
and U9446 (N_9446,N_8422,N_8598);
and U9447 (N_9447,N_8423,N_8549);
xor U9448 (N_9448,N_8443,N_8852);
nor U9449 (N_9449,N_8797,N_8820);
or U9450 (N_9450,N_8452,N_8750);
xnor U9451 (N_9451,N_8784,N_8592);
nor U9452 (N_9452,N_8917,N_8939);
xnor U9453 (N_9453,N_8789,N_8679);
nor U9454 (N_9454,N_8435,N_8675);
and U9455 (N_9455,N_8467,N_8476);
nand U9456 (N_9456,N_8954,N_8509);
or U9457 (N_9457,N_8430,N_8818);
nand U9458 (N_9458,N_8993,N_8936);
xnor U9459 (N_9459,N_8782,N_8909);
xnor U9460 (N_9460,N_8852,N_8605);
nand U9461 (N_9461,N_8943,N_8805);
and U9462 (N_9462,N_8447,N_8662);
and U9463 (N_9463,N_8850,N_8786);
nand U9464 (N_9464,N_8633,N_8554);
nand U9465 (N_9465,N_8599,N_8782);
nor U9466 (N_9466,N_8558,N_8925);
nor U9467 (N_9467,N_8418,N_8989);
nand U9468 (N_9468,N_8421,N_8812);
nand U9469 (N_9469,N_8735,N_8576);
nor U9470 (N_9470,N_8574,N_8491);
nand U9471 (N_9471,N_8713,N_8882);
nand U9472 (N_9472,N_8486,N_8474);
and U9473 (N_9473,N_8863,N_8683);
or U9474 (N_9474,N_8455,N_8607);
or U9475 (N_9475,N_8619,N_8452);
or U9476 (N_9476,N_8644,N_8415);
and U9477 (N_9477,N_8683,N_8408);
xnor U9478 (N_9478,N_8569,N_8947);
and U9479 (N_9479,N_8442,N_8438);
nand U9480 (N_9480,N_8556,N_8871);
nor U9481 (N_9481,N_8650,N_8423);
nor U9482 (N_9482,N_8995,N_8884);
nand U9483 (N_9483,N_8452,N_8547);
nand U9484 (N_9484,N_8677,N_8667);
nand U9485 (N_9485,N_8751,N_8448);
xnor U9486 (N_9486,N_8431,N_8976);
or U9487 (N_9487,N_8874,N_8968);
nand U9488 (N_9488,N_8616,N_8844);
nor U9489 (N_9489,N_8547,N_8606);
nand U9490 (N_9490,N_8454,N_8779);
and U9491 (N_9491,N_8732,N_8473);
xnor U9492 (N_9492,N_8540,N_8550);
or U9493 (N_9493,N_8875,N_8837);
or U9494 (N_9494,N_8916,N_8932);
and U9495 (N_9495,N_8961,N_8590);
xnor U9496 (N_9496,N_8620,N_8479);
and U9497 (N_9497,N_8872,N_8402);
xnor U9498 (N_9498,N_8831,N_8815);
and U9499 (N_9499,N_8559,N_8513);
xor U9500 (N_9500,N_8497,N_8443);
nand U9501 (N_9501,N_8732,N_8563);
or U9502 (N_9502,N_8541,N_8723);
nor U9503 (N_9503,N_8946,N_8739);
and U9504 (N_9504,N_8465,N_8510);
nand U9505 (N_9505,N_8806,N_8743);
nand U9506 (N_9506,N_8499,N_8411);
xnor U9507 (N_9507,N_8910,N_8897);
and U9508 (N_9508,N_8864,N_8622);
and U9509 (N_9509,N_8859,N_8930);
xor U9510 (N_9510,N_8419,N_8632);
xor U9511 (N_9511,N_8529,N_8550);
nor U9512 (N_9512,N_8547,N_8675);
and U9513 (N_9513,N_8790,N_8558);
and U9514 (N_9514,N_8705,N_8906);
and U9515 (N_9515,N_8959,N_8877);
nor U9516 (N_9516,N_8961,N_8549);
or U9517 (N_9517,N_8676,N_8696);
or U9518 (N_9518,N_8495,N_8764);
nand U9519 (N_9519,N_8555,N_8724);
xnor U9520 (N_9520,N_8480,N_8892);
nor U9521 (N_9521,N_8588,N_8406);
nor U9522 (N_9522,N_8873,N_8760);
xor U9523 (N_9523,N_8891,N_8649);
nor U9524 (N_9524,N_8670,N_8738);
xor U9525 (N_9525,N_8850,N_8778);
or U9526 (N_9526,N_8842,N_8641);
and U9527 (N_9527,N_8495,N_8718);
xor U9528 (N_9528,N_8404,N_8849);
or U9529 (N_9529,N_8820,N_8879);
or U9530 (N_9530,N_8493,N_8452);
xor U9531 (N_9531,N_8614,N_8576);
or U9532 (N_9532,N_8729,N_8471);
and U9533 (N_9533,N_8403,N_8772);
nor U9534 (N_9534,N_8668,N_8541);
nor U9535 (N_9535,N_8699,N_8822);
nor U9536 (N_9536,N_8934,N_8764);
xnor U9537 (N_9537,N_8806,N_8796);
and U9538 (N_9538,N_8488,N_8467);
nand U9539 (N_9539,N_8799,N_8995);
xor U9540 (N_9540,N_8553,N_8598);
or U9541 (N_9541,N_8704,N_8690);
nand U9542 (N_9542,N_8506,N_8411);
or U9543 (N_9543,N_8637,N_8828);
nand U9544 (N_9544,N_8702,N_8416);
and U9545 (N_9545,N_8968,N_8811);
and U9546 (N_9546,N_8723,N_8918);
or U9547 (N_9547,N_8450,N_8905);
and U9548 (N_9548,N_8924,N_8530);
or U9549 (N_9549,N_8430,N_8637);
nand U9550 (N_9550,N_8966,N_8944);
xnor U9551 (N_9551,N_8577,N_8775);
nand U9552 (N_9552,N_8405,N_8720);
or U9553 (N_9553,N_8846,N_8663);
and U9554 (N_9554,N_8632,N_8953);
xnor U9555 (N_9555,N_8964,N_8713);
and U9556 (N_9556,N_8457,N_8725);
and U9557 (N_9557,N_8567,N_8632);
or U9558 (N_9558,N_8847,N_8912);
xor U9559 (N_9559,N_8728,N_8588);
or U9560 (N_9560,N_8609,N_8529);
nor U9561 (N_9561,N_8931,N_8896);
xnor U9562 (N_9562,N_8615,N_8884);
xor U9563 (N_9563,N_8563,N_8546);
and U9564 (N_9564,N_8405,N_8908);
xnor U9565 (N_9565,N_8884,N_8915);
xnor U9566 (N_9566,N_8927,N_8655);
xor U9567 (N_9567,N_8750,N_8562);
nand U9568 (N_9568,N_8584,N_8826);
nor U9569 (N_9569,N_8496,N_8754);
nor U9570 (N_9570,N_8469,N_8749);
nor U9571 (N_9571,N_8418,N_8750);
xnor U9572 (N_9572,N_8573,N_8531);
nor U9573 (N_9573,N_8570,N_8436);
or U9574 (N_9574,N_8689,N_8936);
and U9575 (N_9575,N_8924,N_8975);
and U9576 (N_9576,N_8791,N_8690);
xor U9577 (N_9577,N_8806,N_8563);
xor U9578 (N_9578,N_8449,N_8828);
and U9579 (N_9579,N_8516,N_8795);
or U9580 (N_9580,N_8536,N_8927);
nor U9581 (N_9581,N_8795,N_8425);
xor U9582 (N_9582,N_8703,N_8796);
xnor U9583 (N_9583,N_8610,N_8716);
or U9584 (N_9584,N_8648,N_8623);
or U9585 (N_9585,N_8919,N_8415);
xor U9586 (N_9586,N_8732,N_8409);
nor U9587 (N_9587,N_8935,N_8757);
xnor U9588 (N_9588,N_8728,N_8966);
and U9589 (N_9589,N_8872,N_8865);
nand U9590 (N_9590,N_8609,N_8421);
nand U9591 (N_9591,N_8479,N_8418);
or U9592 (N_9592,N_8966,N_8861);
nor U9593 (N_9593,N_8742,N_8955);
or U9594 (N_9594,N_8955,N_8642);
nor U9595 (N_9595,N_8428,N_8926);
nand U9596 (N_9596,N_8751,N_8893);
or U9597 (N_9597,N_8741,N_8519);
nor U9598 (N_9598,N_8873,N_8948);
xnor U9599 (N_9599,N_8462,N_8649);
xor U9600 (N_9600,N_9348,N_9030);
and U9601 (N_9601,N_9451,N_9188);
or U9602 (N_9602,N_9059,N_9102);
and U9603 (N_9603,N_9118,N_9191);
nand U9604 (N_9604,N_9501,N_9584);
nor U9605 (N_9605,N_9496,N_9493);
and U9606 (N_9606,N_9548,N_9042);
and U9607 (N_9607,N_9587,N_9016);
xor U9608 (N_9608,N_9307,N_9519);
nand U9609 (N_9609,N_9260,N_9511);
xor U9610 (N_9610,N_9043,N_9359);
xnor U9611 (N_9611,N_9277,N_9061);
xor U9612 (N_9612,N_9007,N_9342);
nand U9613 (N_9613,N_9055,N_9251);
nor U9614 (N_9614,N_9082,N_9326);
nor U9615 (N_9615,N_9269,N_9179);
nor U9616 (N_9616,N_9427,N_9202);
nor U9617 (N_9617,N_9544,N_9418);
and U9618 (N_9618,N_9457,N_9370);
and U9619 (N_9619,N_9015,N_9445);
xnor U9620 (N_9620,N_9454,N_9396);
and U9621 (N_9621,N_9143,N_9324);
nand U9622 (N_9622,N_9442,N_9489);
nand U9623 (N_9623,N_9539,N_9432);
or U9624 (N_9624,N_9368,N_9469);
xor U9625 (N_9625,N_9154,N_9001);
or U9626 (N_9626,N_9570,N_9170);
or U9627 (N_9627,N_9431,N_9062);
nand U9628 (N_9628,N_9379,N_9239);
or U9629 (N_9629,N_9228,N_9258);
nor U9630 (N_9630,N_9175,N_9421);
xnor U9631 (N_9631,N_9448,N_9416);
or U9632 (N_9632,N_9337,N_9483);
nand U9633 (N_9633,N_9000,N_9381);
nor U9634 (N_9634,N_9299,N_9078);
xor U9635 (N_9635,N_9279,N_9098);
nor U9636 (N_9636,N_9031,N_9210);
and U9637 (N_9637,N_9458,N_9585);
nor U9638 (N_9638,N_9088,N_9012);
nor U9639 (N_9639,N_9259,N_9306);
nand U9640 (N_9640,N_9387,N_9116);
and U9641 (N_9641,N_9119,N_9275);
nand U9642 (N_9642,N_9014,N_9415);
xnor U9643 (N_9643,N_9231,N_9545);
nand U9644 (N_9644,N_9339,N_9124);
nor U9645 (N_9645,N_9140,N_9192);
nor U9646 (N_9646,N_9595,N_9047);
xor U9647 (N_9647,N_9443,N_9298);
xor U9648 (N_9648,N_9166,N_9343);
nor U9649 (N_9649,N_9171,N_9336);
xnor U9650 (N_9650,N_9321,N_9005);
nand U9651 (N_9651,N_9477,N_9598);
and U9652 (N_9652,N_9543,N_9145);
nor U9653 (N_9653,N_9214,N_9033);
and U9654 (N_9654,N_9487,N_9159);
xnor U9655 (N_9655,N_9104,N_9195);
nor U9656 (N_9656,N_9495,N_9280);
or U9657 (N_9657,N_9472,N_9450);
nor U9658 (N_9658,N_9232,N_9045);
or U9659 (N_9659,N_9272,N_9108);
nand U9660 (N_9660,N_9129,N_9211);
and U9661 (N_9661,N_9024,N_9224);
xnor U9662 (N_9662,N_9329,N_9041);
or U9663 (N_9663,N_9026,N_9138);
or U9664 (N_9664,N_9546,N_9254);
and U9665 (N_9665,N_9130,N_9486);
xnor U9666 (N_9666,N_9360,N_9578);
nand U9667 (N_9667,N_9237,N_9407);
and U9668 (N_9668,N_9067,N_9048);
xnor U9669 (N_9669,N_9468,N_9592);
or U9670 (N_9670,N_9131,N_9074);
and U9671 (N_9671,N_9392,N_9494);
nor U9672 (N_9672,N_9182,N_9185);
or U9673 (N_9673,N_9221,N_9293);
nor U9674 (N_9674,N_9471,N_9250);
or U9675 (N_9675,N_9412,N_9169);
and U9676 (N_9676,N_9080,N_9184);
and U9677 (N_9677,N_9025,N_9564);
nor U9678 (N_9678,N_9513,N_9435);
nand U9679 (N_9679,N_9066,N_9197);
and U9680 (N_9680,N_9127,N_9245);
nor U9681 (N_9681,N_9597,N_9424);
nand U9682 (N_9682,N_9373,N_9036);
or U9683 (N_9683,N_9401,N_9400);
or U9684 (N_9684,N_9155,N_9346);
nand U9685 (N_9685,N_9205,N_9198);
nor U9686 (N_9686,N_9302,N_9094);
or U9687 (N_9687,N_9527,N_9109);
and U9688 (N_9688,N_9242,N_9203);
xor U9689 (N_9689,N_9573,N_9463);
nor U9690 (N_9690,N_9535,N_9453);
nor U9691 (N_9691,N_9426,N_9163);
nand U9692 (N_9692,N_9518,N_9478);
nand U9693 (N_9693,N_9183,N_9485);
nor U9694 (N_9694,N_9404,N_9219);
or U9695 (N_9695,N_9332,N_9399);
and U9696 (N_9696,N_9069,N_9551);
and U9697 (N_9697,N_9114,N_9167);
nand U9698 (N_9698,N_9514,N_9086);
or U9699 (N_9699,N_9218,N_9054);
and U9700 (N_9700,N_9582,N_9206);
nand U9701 (N_9701,N_9561,N_9452);
nand U9702 (N_9702,N_9390,N_9523);
xnor U9703 (N_9703,N_9319,N_9460);
nand U9704 (N_9704,N_9076,N_9576);
or U9705 (N_9705,N_9349,N_9240);
xnor U9706 (N_9706,N_9344,N_9097);
and U9707 (N_9707,N_9049,N_9236);
xor U9708 (N_9708,N_9509,N_9320);
nand U9709 (N_9709,N_9436,N_9158);
xor U9710 (N_9710,N_9372,N_9276);
or U9711 (N_9711,N_9227,N_9017);
and U9712 (N_9712,N_9134,N_9382);
nor U9713 (N_9713,N_9071,N_9503);
nor U9714 (N_9714,N_9340,N_9393);
xnor U9715 (N_9715,N_9287,N_9540);
and U9716 (N_9716,N_9314,N_9538);
xor U9717 (N_9717,N_9365,N_9222);
and U9718 (N_9718,N_9318,N_9084);
or U9719 (N_9719,N_9103,N_9447);
xor U9720 (N_9720,N_9056,N_9357);
nor U9721 (N_9721,N_9482,N_9196);
nand U9722 (N_9722,N_9207,N_9402);
or U9723 (N_9723,N_9374,N_9225);
xor U9724 (N_9724,N_9208,N_9316);
nor U9725 (N_9725,N_9006,N_9310);
nor U9726 (N_9726,N_9201,N_9480);
and U9727 (N_9727,N_9586,N_9520);
or U9728 (N_9728,N_9052,N_9364);
xor U9729 (N_9729,N_9438,N_9474);
xnor U9730 (N_9730,N_9051,N_9212);
xor U9731 (N_9731,N_9593,N_9353);
xor U9732 (N_9732,N_9274,N_9273);
nor U9733 (N_9733,N_9467,N_9408);
nand U9734 (N_9734,N_9488,N_9093);
and U9735 (N_9735,N_9281,N_9405);
xor U9736 (N_9736,N_9554,N_9568);
nand U9737 (N_9737,N_9216,N_9040);
nand U9738 (N_9738,N_9362,N_9238);
nor U9739 (N_9739,N_9456,N_9200);
or U9740 (N_9740,N_9013,N_9296);
and U9741 (N_9741,N_9252,N_9283);
and U9742 (N_9742,N_9376,N_9128);
nor U9743 (N_9743,N_9367,N_9434);
xnor U9744 (N_9744,N_9220,N_9092);
or U9745 (N_9745,N_9149,N_9068);
nor U9746 (N_9746,N_9429,N_9046);
and U9747 (N_9747,N_9057,N_9534);
and U9748 (N_9748,N_9596,N_9053);
and U9749 (N_9749,N_9085,N_9304);
and U9750 (N_9750,N_9562,N_9479);
nand U9751 (N_9751,N_9151,N_9526);
xor U9752 (N_9752,N_9204,N_9464);
or U9753 (N_9753,N_9571,N_9136);
xnor U9754 (N_9754,N_9120,N_9035);
and U9755 (N_9755,N_9446,N_9162);
or U9756 (N_9756,N_9403,N_9270);
xnor U9757 (N_9757,N_9261,N_9023);
and U9758 (N_9758,N_9515,N_9249);
nand U9759 (N_9759,N_9366,N_9462);
nor U9760 (N_9760,N_9498,N_9060);
or U9761 (N_9761,N_9579,N_9234);
and U9762 (N_9762,N_9223,N_9099);
nor U9763 (N_9763,N_9027,N_9572);
xor U9764 (N_9764,N_9009,N_9248);
xnor U9765 (N_9765,N_9301,N_9284);
or U9766 (N_9766,N_9157,N_9411);
or U9767 (N_9767,N_9389,N_9461);
and U9768 (N_9768,N_9377,N_9504);
or U9769 (N_9769,N_9295,N_9107);
nand U9770 (N_9770,N_9029,N_9090);
nor U9771 (N_9771,N_9081,N_9294);
or U9772 (N_9772,N_9020,N_9430);
and U9773 (N_9773,N_9406,N_9288);
and U9774 (N_9774,N_9338,N_9268);
or U9775 (N_9775,N_9285,N_9358);
and U9776 (N_9776,N_9063,N_9309);
and U9777 (N_9777,N_9531,N_9363);
and U9778 (N_9778,N_9075,N_9492);
nor U9779 (N_9779,N_9428,N_9002);
nand U9780 (N_9780,N_9133,N_9557);
or U9781 (N_9781,N_9065,N_9152);
or U9782 (N_9782,N_9267,N_9559);
or U9783 (N_9783,N_9325,N_9034);
or U9784 (N_9784,N_9290,N_9345);
nand U9785 (N_9785,N_9150,N_9126);
nand U9786 (N_9786,N_9541,N_9575);
nor U9787 (N_9787,N_9064,N_9213);
nor U9788 (N_9788,N_9186,N_9165);
xor U9789 (N_9789,N_9555,N_9289);
xor U9790 (N_9790,N_9044,N_9141);
nand U9791 (N_9791,N_9230,N_9437);
nor U9792 (N_9792,N_9282,N_9502);
xor U9793 (N_9793,N_9278,N_9187);
and U9794 (N_9794,N_9079,N_9466);
nand U9795 (N_9795,N_9243,N_9414);
nand U9796 (N_9796,N_9148,N_9160);
or U9797 (N_9797,N_9137,N_9308);
or U9798 (N_9798,N_9199,N_9022);
or U9799 (N_9799,N_9004,N_9524);
or U9800 (N_9800,N_9083,N_9265);
and U9801 (N_9801,N_9423,N_9589);
nand U9802 (N_9802,N_9476,N_9386);
nand U9803 (N_9803,N_9096,N_9574);
xnor U9804 (N_9804,N_9491,N_9413);
or U9805 (N_9805,N_9566,N_9588);
nand U9806 (N_9806,N_9369,N_9533);
or U9807 (N_9807,N_9591,N_9522);
nor U9808 (N_9808,N_9139,N_9590);
xor U9809 (N_9809,N_9072,N_9341);
and U9810 (N_9810,N_9173,N_9172);
xor U9811 (N_9811,N_9422,N_9168);
xor U9812 (N_9812,N_9244,N_9560);
nand U9813 (N_9813,N_9410,N_9322);
or U9814 (N_9814,N_9567,N_9398);
or U9815 (N_9815,N_9516,N_9180);
nor U9816 (N_9816,N_9475,N_9193);
or U9817 (N_9817,N_9153,N_9100);
nand U9818 (N_9818,N_9132,N_9111);
nand U9819 (N_9819,N_9356,N_9003);
and U9820 (N_9820,N_9508,N_9256);
and U9821 (N_9821,N_9217,N_9444);
xor U9822 (N_9822,N_9537,N_9105);
xnor U9823 (N_9823,N_9176,N_9313);
nor U9824 (N_9824,N_9021,N_9305);
nor U9825 (N_9825,N_9383,N_9552);
or U9826 (N_9826,N_9178,N_9510);
nand U9827 (N_9827,N_9378,N_9490);
xnor U9828 (N_9828,N_9121,N_9384);
or U9829 (N_9829,N_9528,N_9297);
and U9830 (N_9830,N_9433,N_9556);
nand U9831 (N_9831,N_9599,N_9292);
xor U9832 (N_9832,N_9312,N_9594);
or U9833 (N_9833,N_9323,N_9095);
and U9834 (N_9834,N_9300,N_9465);
nor U9835 (N_9835,N_9380,N_9529);
or U9836 (N_9836,N_9473,N_9011);
or U9837 (N_9837,N_9177,N_9558);
nor U9838 (N_9838,N_9583,N_9209);
nor U9839 (N_9839,N_9091,N_9512);
or U9840 (N_9840,N_9229,N_9164);
nor U9841 (N_9841,N_9101,N_9135);
nor U9842 (N_9842,N_9507,N_9439);
or U9843 (N_9843,N_9500,N_9263);
and U9844 (N_9844,N_9241,N_9147);
xor U9845 (N_9845,N_9351,N_9089);
and U9846 (N_9846,N_9361,N_9246);
nand U9847 (N_9847,N_9459,N_9073);
and U9848 (N_9848,N_9580,N_9335);
nand U9849 (N_9849,N_9577,N_9255);
nor U9850 (N_9850,N_9506,N_9194);
nor U9851 (N_9851,N_9455,N_9536);
and U9852 (N_9852,N_9233,N_9032);
xor U9853 (N_9853,N_9257,N_9350);
and U9854 (N_9854,N_9530,N_9226);
nand U9855 (N_9855,N_9122,N_9481);
xor U9856 (N_9856,N_9247,N_9355);
or U9857 (N_9857,N_9028,N_9550);
xnor U9858 (N_9858,N_9517,N_9395);
nor U9859 (N_9859,N_9497,N_9058);
nor U9860 (N_9860,N_9328,N_9334);
nor U9861 (N_9861,N_9581,N_9266);
nor U9862 (N_9862,N_9235,N_9070);
xor U9863 (N_9863,N_9125,N_9253);
or U9864 (N_9864,N_9008,N_9569);
xnor U9865 (N_9865,N_9038,N_9375);
and U9866 (N_9866,N_9330,N_9315);
nor U9867 (N_9867,N_9394,N_9037);
nand U9868 (N_9868,N_9333,N_9050);
nand U9869 (N_9869,N_9391,N_9142);
or U9870 (N_9870,N_9449,N_9117);
nor U9871 (N_9871,N_9317,N_9417);
or U9872 (N_9872,N_9542,N_9420);
nand U9873 (N_9873,N_9019,N_9553);
and U9874 (N_9874,N_9397,N_9010);
nor U9875 (N_9875,N_9156,N_9264);
nand U9876 (N_9876,N_9499,N_9347);
or U9877 (N_9877,N_9371,N_9505);
nor U9878 (N_9878,N_9388,N_9087);
nor U9879 (N_9879,N_9291,N_9215);
nand U9880 (N_9880,N_9262,N_9271);
nor U9881 (N_9881,N_9440,N_9525);
nand U9882 (N_9882,N_9484,N_9521);
or U9883 (N_9883,N_9425,N_9409);
nor U9884 (N_9884,N_9115,N_9077);
or U9885 (N_9885,N_9113,N_9331);
and U9886 (N_9886,N_9112,N_9123);
xor U9887 (N_9887,N_9385,N_9106);
nor U9888 (N_9888,N_9146,N_9470);
nand U9889 (N_9889,N_9018,N_9286);
nand U9890 (N_9890,N_9327,N_9110);
and U9891 (N_9891,N_9532,N_9441);
and U9892 (N_9892,N_9190,N_9419);
nand U9893 (N_9893,N_9354,N_9303);
nand U9894 (N_9894,N_9181,N_9352);
and U9895 (N_9895,N_9144,N_9311);
xor U9896 (N_9896,N_9039,N_9565);
nor U9897 (N_9897,N_9563,N_9161);
nor U9898 (N_9898,N_9189,N_9174);
nor U9899 (N_9899,N_9547,N_9549);
nand U9900 (N_9900,N_9016,N_9041);
xnor U9901 (N_9901,N_9267,N_9587);
nor U9902 (N_9902,N_9094,N_9061);
xnor U9903 (N_9903,N_9417,N_9247);
or U9904 (N_9904,N_9097,N_9509);
nand U9905 (N_9905,N_9339,N_9499);
and U9906 (N_9906,N_9004,N_9256);
nor U9907 (N_9907,N_9428,N_9194);
or U9908 (N_9908,N_9449,N_9452);
nand U9909 (N_9909,N_9030,N_9375);
or U9910 (N_9910,N_9494,N_9384);
nand U9911 (N_9911,N_9054,N_9284);
nor U9912 (N_9912,N_9166,N_9148);
xor U9913 (N_9913,N_9069,N_9516);
xnor U9914 (N_9914,N_9556,N_9021);
xor U9915 (N_9915,N_9366,N_9536);
xor U9916 (N_9916,N_9557,N_9222);
and U9917 (N_9917,N_9577,N_9375);
nand U9918 (N_9918,N_9174,N_9285);
and U9919 (N_9919,N_9569,N_9229);
xnor U9920 (N_9920,N_9573,N_9498);
nand U9921 (N_9921,N_9572,N_9075);
xor U9922 (N_9922,N_9364,N_9521);
xor U9923 (N_9923,N_9050,N_9014);
or U9924 (N_9924,N_9575,N_9491);
or U9925 (N_9925,N_9287,N_9272);
nand U9926 (N_9926,N_9261,N_9504);
nor U9927 (N_9927,N_9544,N_9249);
xor U9928 (N_9928,N_9216,N_9539);
xor U9929 (N_9929,N_9296,N_9468);
or U9930 (N_9930,N_9171,N_9294);
or U9931 (N_9931,N_9417,N_9369);
nand U9932 (N_9932,N_9221,N_9125);
or U9933 (N_9933,N_9570,N_9194);
xnor U9934 (N_9934,N_9064,N_9137);
nand U9935 (N_9935,N_9008,N_9273);
nor U9936 (N_9936,N_9201,N_9394);
or U9937 (N_9937,N_9359,N_9271);
and U9938 (N_9938,N_9214,N_9122);
nor U9939 (N_9939,N_9516,N_9360);
and U9940 (N_9940,N_9483,N_9215);
nor U9941 (N_9941,N_9175,N_9343);
nand U9942 (N_9942,N_9420,N_9127);
xor U9943 (N_9943,N_9406,N_9377);
and U9944 (N_9944,N_9135,N_9380);
nand U9945 (N_9945,N_9452,N_9227);
and U9946 (N_9946,N_9401,N_9041);
xnor U9947 (N_9947,N_9318,N_9256);
xnor U9948 (N_9948,N_9289,N_9436);
nand U9949 (N_9949,N_9007,N_9596);
or U9950 (N_9950,N_9079,N_9248);
xnor U9951 (N_9951,N_9025,N_9193);
and U9952 (N_9952,N_9146,N_9003);
nand U9953 (N_9953,N_9083,N_9327);
or U9954 (N_9954,N_9081,N_9554);
xnor U9955 (N_9955,N_9125,N_9559);
or U9956 (N_9956,N_9226,N_9389);
and U9957 (N_9957,N_9508,N_9087);
or U9958 (N_9958,N_9242,N_9214);
nor U9959 (N_9959,N_9595,N_9504);
xnor U9960 (N_9960,N_9118,N_9551);
xnor U9961 (N_9961,N_9578,N_9102);
xor U9962 (N_9962,N_9227,N_9543);
or U9963 (N_9963,N_9213,N_9339);
xnor U9964 (N_9964,N_9554,N_9249);
and U9965 (N_9965,N_9067,N_9263);
and U9966 (N_9966,N_9568,N_9534);
or U9967 (N_9967,N_9059,N_9377);
and U9968 (N_9968,N_9020,N_9374);
nand U9969 (N_9969,N_9043,N_9065);
nand U9970 (N_9970,N_9460,N_9569);
and U9971 (N_9971,N_9039,N_9023);
or U9972 (N_9972,N_9580,N_9541);
xor U9973 (N_9973,N_9031,N_9315);
xor U9974 (N_9974,N_9344,N_9247);
nor U9975 (N_9975,N_9299,N_9016);
nor U9976 (N_9976,N_9098,N_9538);
nor U9977 (N_9977,N_9399,N_9031);
or U9978 (N_9978,N_9379,N_9034);
or U9979 (N_9979,N_9128,N_9595);
nand U9980 (N_9980,N_9599,N_9238);
or U9981 (N_9981,N_9192,N_9223);
xnor U9982 (N_9982,N_9588,N_9328);
xnor U9983 (N_9983,N_9348,N_9136);
and U9984 (N_9984,N_9038,N_9172);
nand U9985 (N_9985,N_9392,N_9168);
and U9986 (N_9986,N_9173,N_9238);
xnor U9987 (N_9987,N_9099,N_9118);
xor U9988 (N_9988,N_9532,N_9095);
or U9989 (N_9989,N_9194,N_9372);
xnor U9990 (N_9990,N_9566,N_9468);
nor U9991 (N_9991,N_9428,N_9453);
nand U9992 (N_9992,N_9131,N_9241);
and U9993 (N_9993,N_9535,N_9126);
and U9994 (N_9994,N_9566,N_9280);
or U9995 (N_9995,N_9042,N_9241);
nor U9996 (N_9996,N_9031,N_9156);
nor U9997 (N_9997,N_9218,N_9431);
nor U9998 (N_9998,N_9557,N_9049);
and U9999 (N_9999,N_9077,N_9287);
and U10000 (N_10000,N_9240,N_9157);
or U10001 (N_10001,N_9551,N_9196);
nor U10002 (N_10002,N_9357,N_9476);
xnor U10003 (N_10003,N_9093,N_9529);
xnor U10004 (N_10004,N_9141,N_9578);
and U10005 (N_10005,N_9152,N_9522);
and U10006 (N_10006,N_9355,N_9324);
nor U10007 (N_10007,N_9289,N_9089);
and U10008 (N_10008,N_9257,N_9599);
nor U10009 (N_10009,N_9432,N_9013);
or U10010 (N_10010,N_9598,N_9168);
nand U10011 (N_10011,N_9024,N_9223);
nor U10012 (N_10012,N_9002,N_9287);
or U10013 (N_10013,N_9062,N_9087);
nand U10014 (N_10014,N_9402,N_9131);
nor U10015 (N_10015,N_9324,N_9523);
xnor U10016 (N_10016,N_9393,N_9285);
xnor U10017 (N_10017,N_9275,N_9511);
nor U10018 (N_10018,N_9459,N_9078);
nor U10019 (N_10019,N_9003,N_9159);
xnor U10020 (N_10020,N_9214,N_9505);
xnor U10021 (N_10021,N_9291,N_9222);
nand U10022 (N_10022,N_9395,N_9305);
or U10023 (N_10023,N_9279,N_9411);
or U10024 (N_10024,N_9457,N_9189);
xor U10025 (N_10025,N_9327,N_9092);
nor U10026 (N_10026,N_9167,N_9482);
and U10027 (N_10027,N_9418,N_9370);
or U10028 (N_10028,N_9133,N_9300);
nor U10029 (N_10029,N_9131,N_9465);
nor U10030 (N_10030,N_9583,N_9037);
xnor U10031 (N_10031,N_9117,N_9148);
xor U10032 (N_10032,N_9276,N_9169);
xor U10033 (N_10033,N_9151,N_9475);
or U10034 (N_10034,N_9043,N_9278);
xnor U10035 (N_10035,N_9084,N_9259);
nand U10036 (N_10036,N_9058,N_9582);
nand U10037 (N_10037,N_9561,N_9319);
xnor U10038 (N_10038,N_9313,N_9220);
nand U10039 (N_10039,N_9329,N_9081);
or U10040 (N_10040,N_9048,N_9246);
or U10041 (N_10041,N_9495,N_9175);
xnor U10042 (N_10042,N_9579,N_9403);
nand U10043 (N_10043,N_9144,N_9077);
nor U10044 (N_10044,N_9006,N_9296);
nand U10045 (N_10045,N_9072,N_9058);
nor U10046 (N_10046,N_9137,N_9299);
nor U10047 (N_10047,N_9320,N_9474);
or U10048 (N_10048,N_9579,N_9502);
nor U10049 (N_10049,N_9006,N_9271);
or U10050 (N_10050,N_9028,N_9483);
and U10051 (N_10051,N_9224,N_9582);
and U10052 (N_10052,N_9213,N_9016);
nor U10053 (N_10053,N_9490,N_9304);
xnor U10054 (N_10054,N_9025,N_9520);
nand U10055 (N_10055,N_9315,N_9273);
xor U10056 (N_10056,N_9040,N_9315);
xor U10057 (N_10057,N_9398,N_9068);
or U10058 (N_10058,N_9364,N_9556);
xnor U10059 (N_10059,N_9446,N_9072);
nor U10060 (N_10060,N_9493,N_9275);
and U10061 (N_10061,N_9573,N_9090);
and U10062 (N_10062,N_9107,N_9347);
or U10063 (N_10063,N_9000,N_9170);
nor U10064 (N_10064,N_9474,N_9350);
and U10065 (N_10065,N_9166,N_9467);
nand U10066 (N_10066,N_9133,N_9554);
or U10067 (N_10067,N_9344,N_9145);
and U10068 (N_10068,N_9525,N_9520);
or U10069 (N_10069,N_9151,N_9444);
or U10070 (N_10070,N_9137,N_9162);
xnor U10071 (N_10071,N_9479,N_9450);
nor U10072 (N_10072,N_9057,N_9438);
xor U10073 (N_10073,N_9484,N_9336);
or U10074 (N_10074,N_9179,N_9131);
xnor U10075 (N_10075,N_9385,N_9311);
or U10076 (N_10076,N_9337,N_9258);
xnor U10077 (N_10077,N_9195,N_9253);
nor U10078 (N_10078,N_9436,N_9019);
or U10079 (N_10079,N_9599,N_9154);
and U10080 (N_10080,N_9378,N_9251);
or U10081 (N_10081,N_9261,N_9242);
and U10082 (N_10082,N_9302,N_9027);
nand U10083 (N_10083,N_9564,N_9079);
xor U10084 (N_10084,N_9529,N_9514);
nand U10085 (N_10085,N_9187,N_9153);
nor U10086 (N_10086,N_9036,N_9561);
nand U10087 (N_10087,N_9566,N_9447);
and U10088 (N_10088,N_9468,N_9047);
nand U10089 (N_10089,N_9407,N_9564);
nor U10090 (N_10090,N_9264,N_9429);
or U10091 (N_10091,N_9466,N_9118);
xor U10092 (N_10092,N_9473,N_9162);
xor U10093 (N_10093,N_9526,N_9268);
and U10094 (N_10094,N_9363,N_9380);
nor U10095 (N_10095,N_9091,N_9462);
xor U10096 (N_10096,N_9207,N_9233);
and U10097 (N_10097,N_9133,N_9084);
nor U10098 (N_10098,N_9324,N_9375);
nor U10099 (N_10099,N_9590,N_9545);
xnor U10100 (N_10100,N_9336,N_9575);
nor U10101 (N_10101,N_9327,N_9446);
nor U10102 (N_10102,N_9230,N_9312);
nand U10103 (N_10103,N_9064,N_9528);
and U10104 (N_10104,N_9566,N_9188);
and U10105 (N_10105,N_9363,N_9587);
nor U10106 (N_10106,N_9306,N_9155);
or U10107 (N_10107,N_9062,N_9506);
xnor U10108 (N_10108,N_9559,N_9544);
and U10109 (N_10109,N_9204,N_9240);
nand U10110 (N_10110,N_9088,N_9103);
nand U10111 (N_10111,N_9089,N_9193);
or U10112 (N_10112,N_9575,N_9408);
nor U10113 (N_10113,N_9555,N_9254);
nor U10114 (N_10114,N_9146,N_9070);
and U10115 (N_10115,N_9353,N_9166);
nor U10116 (N_10116,N_9425,N_9315);
xor U10117 (N_10117,N_9196,N_9219);
nor U10118 (N_10118,N_9174,N_9597);
and U10119 (N_10119,N_9487,N_9238);
and U10120 (N_10120,N_9391,N_9569);
or U10121 (N_10121,N_9294,N_9431);
and U10122 (N_10122,N_9465,N_9026);
nand U10123 (N_10123,N_9326,N_9599);
xor U10124 (N_10124,N_9415,N_9544);
or U10125 (N_10125,N_9152,N_9010);
and U10126 (N_10126,N_9543,N_9544);
nor U10127 (N_10127,N_9121,N_9015);
nor U10128 (N_10128,N_9172,N_9547);
nor U10129 (N_10129,N_9165,N_9366);
nand U10130 (N_10130,N_9531,N_9302);
nor U10131 (N_10131,N_9194,N_9525);
and U10132 (N_10132,N_9545,N_9002);
nor U10133 (N_10133,N_9324,N_9549);
nor U10134 (N_10134,N_9064,N_9542);
nor U10135 (N_10135,N_9532,N_9419);
xor U10136 (N_10136,N_9009,N_9352);
nand U10137 (N_10137,N_9290,N_9434);
nor U10138 (N_10138,N_9460,N_9154);
xor U10139 (N_10139,N_9556,N_9360);
xnor U10140 (N_10140,N_9282,N_9020);
nand U10141 (N_10141,N_9127,N_9201);
nor U10142 (N_10142,N_9109,N_9169);
nor U10143 (N_10143,N_9415,N_9164);
nor U10144 (N_10144,N_9357,N_9149);
xor U10145 (N_10145,N_9248,N_9143);
nor U10146 (N_10146,N_9031,N_9115);
xnor U10147 (N_10147,N_9418,N_9416);
xor U10148 (N_10148,N_9575,N_9327);
and U10149 (N_10149,N_9544,N_9595);
xnor U10150 (N_10150,N_9028,N_9388);
nand U10151 (N_10151,N_9538,N_9134);
and U10152 (N_10152,N_9096,N_9415);
xnor U10153 (N_10153,N_9054,N_9123);
xor U10154 (N_10154,N_9193,N_9039);
xnor U10155 (N_10155,N_9259,N_9300);
nand U10156 (N_10156,N_9324,N_9259);
or U10157 (N_10157,N_9505,N_9402);
and U10158 (N_10158,N_9482,N_9037);
xnor U10159 (N_10159,N_9063,N_9411);
or U10160 (N_10160,N_9490,N_9025);
xor U10161 (N_10161,N_9050,N_9182);
nor U10162 (N_10162,N_9035,N_9249);
nand U10163 (N_10163,N_9365,N_9347);
nor U10164 (N_10164,N_9510,N_9162);
xor U10165 (N_10165,N_9342,N_9264);
or U10166 (N_10166,N_9353,N_9315);
or U10167 (N_10167,N_9361,N_9059);
nor U10168 (N_10168,N_9376,N_9263);
xnor U10169 (N_10169,N_9548,N_9053);
and U10170 (N_10170,N_9448,N_9571);
xnor U10171 (N_10171,N_9063,N_9532);
nand U10172 (N_10172,N_9007,N_9349);
or U10173 (N_10173,N_9159,N_9170);
nor U10174 (N_10174,N_9026,N_9275);
nor U10175 (N_10175,N_9133,N_9513);
and U10176 (N_10176,N_9480,N_9395);
xnor U10177 (N_10177,N_9100,N_9279);
or U10178 (N_10178,N_9006,N_9400);
and U10179 (N_10179,N_9310,N_9418);
and U10180 (N_10180,N_9508,N_9533);
and U10181 (N_10181,N_9329,N_9394);
or U10182 (N_10182,N_9565,N_9257);
nor U10183 (N_10183,N_9360,N_9305);
or U10184 (N_10184,N_9358,N_9491);
and U10185 (N_10185,N_9211,N_9324);
or U10186 (N_10186,N_9042,N_9549);
or U10187 (N_10187,N_9148,N_9449);
xor U10188 (N_10188,N_9216,N_9428);
or U10189 (N_10189,N_9388,N_9061);
nor U10190 (N_10190,N_9218,N_9098);
nand U10191 (N_10191,N_9115,N_9245);
and U10192 (N_10192,N_9342,N_9069);
nor U10193 (N_10193,N_9475,N_9562);
nand U10194 (N_10194,N_9402,N_9298);
or U10195 (N_10195,N_9095,N_9021);
xor U10196 (N_10196,N_9301,N_9318);
nand U10197 (N_10197,N_9230,N_9362);
xor U10198 (N_10198,N_9066,N_9095);
and U10199 (N_10199,N_9507,N_9401);
nand U10200 (N_10200,N_9852,N_9783);
or U10201 (N_10201,N_9623,N_10185);
and U10202 (N_10202,N_10004,N_9695);
or U10203 (N_10203,N_10163,N_9671);
and U10204 (N_10204,N_9771,N_9950);
nand U10205 (N_10205,N_10048,N_9890);
or U10206 (N_10206,N_9955,N_10002);
xor U10207 (N_10207,N_9896,N_9888);
or U10208 (N_10208,N_10084,N_9702);
nor U10209 (N_10209,N_9629,N_9863);
and U10210 (N_10210,N_9989,N_9869);
and U10211 (N_10211,N_10190,N_10134);
nand U10212 (N_10212,N_10189,N_9934);
or U10213 (N_10213,N_10058,N_9690);
or U10214 (N_10214,N_9954,N_10107);
nand U10215 (N_10215,N_9871,N_9670);
nand U10216 (N_10216,N_10138,N_9612);
and U10217 (N_10217,N_9699,N_9902);
or U10218 (N_10218,N_10060,N_9642);
and U10219 (N_10219,N_9901,N_9772);
and U10220 (N_10220,N_10149,N_9785);
nor U10221 (N_10221,N_10197,N_10109);
nor U10222 (N_10222,N_10122,N_10156);
and U10223 (N_10223,N_9745,N_9880);
and U10224 (N_10224,N_10074,N_9668);
and U10225 (N_10225,N_9627,N_9641);
and U10226 (N_10226,N_10100,N_9821);
and U10227 (N_10227,N_9606,N_9932);
or U10228 (N_10228,N_9698,N_9601);
xor U10229 (N_10229,N_9618,N_9680);
xor U10230 (N_10230,N_9966,N_10042);
and U10231 (N_10231,N_10115,N_9971);
and U10232 (N_10232,N_9986,N_9972);
nor U10233 (N_10233,N_10151,N_10033);
nand U10234 (N_10234,N_9632,N_9631);
xnor U10235 (N_10235,N_10059,N_9761);
nand U10236 (N_10236,N_9640,N_10013);
nor U10237 (N_10237,N_9970,N_10136);
or U10238 (N_10238,N_9665,N_9732);
nor U10239 (N_10239,N_9874,N_9851);
or U10240 (N_10240,N_9870,N_10153);
or U10241 (N_10241,N_9674,N_10086);
and U10242 (N_10242,N_9963,N_9770);
and U10243 (N_10243,N_10167,N_10025);
nor U10244 (N_10244,N_10199,N_9700);
or U10245 (N_10245,N_9886,N_10066);
nor U10246 (N_10246,N_9750,N_10145);
and U10247 (N_10247,N_9915,N_9815);
nor U10248 (N_10248,N_9639,N_9913);
nand U10249 (N_10249,N_10028,N_9843);
nand U10250 (N_10250,N_10106,N_10077);
and U10251 (N_10251,N_9687,N_9756);
and U10252 (N_10252,N_9957,N_10160);
or U10253 (N_10253,N_9914,N_10010);
nor U10254 (N_10254,N_9751,N_9709);
xor U10255 (N_10255,N_10159,N_9602);
xnor U10256 (N_10256,N_9694,N_10112);
nand U10257 (N_10257,N_10079,N_10067);
nor U10258 (N_10258,N_9697,N_9712);
or U10259 (N_10259,N_9620,N_9861);
nor U10260 (N_10260,N_10006,N_9766);
xor U10261 (N_10261,N_10078,N_9867);
xor U10262 (N_10262,N_9776,N_10011);
xnor U10263 (N_10263,N_10144,N_9689);
nor U10264 (N_10264,N_10031,N_10170);
xnor U10265 (N_10265,N_9939,N_10147);
nand U10266 (N_10266,N_9844,N_9795);
or U10267 (N_10267,N_10198,N_9806);
or U10268 (N_10268,N_10009,N_10047);
nand U10269 (N_10269,N_9959,N_9820);
xor U10270 (N_10270,N_9845,N_9824);
xor U10271 (N_10271,N_9865,N_9958);
xnor U10272 (N_10272,N_9762,N_10101);
or U10273 (N_10273,N_9866,N_9946);
xor U10274 (N_10274,N_10049,N_9881);
nand U10275 (N_10275,N_9782,N_9802);
or U10276 (N_10276,N_9969,N_9916);
nor U10277 (N_10277,N_9705,N_9838);
nand U10278 (N_10278,N_9898,N_9884);
and U10279 (N_10279,N_9839,N_9784);
nor U10280 (N_10280,N_10034,N_10166);
nand U10281 (N_10281,N_9685,N_9974);
and U10282 (N_10282,N_9683,N_9610);
and U10283 (N_10283,N_10113,N_10018);
or U10284 (N_10284,N_9737,N_9703);
and U10285 (N_10285,N_10164,N_9625);
nand U10286 (N_10286,N_9895,N_9662);
xor U10287 (N_10287,N_9922,N_9691);
and U10288 (N_10288,N_10098,N_9962);
or U10289 (N_10289,N_10186,N_9764);
or U10290 (N_10290,N_9834,N_10015);
nor U10291 (N_10291,N_9830,N_9677);
or U10292 (N_10292,N_10005,N_10108);
nor U10293 (N_10293,N_9979,N_9775);
nand U10294 (N_10294,N_9807,N_9981);
nand U10295 (N_10295,N_10085,N_9805);
nor U10296 (N_10296,N_10127,N_10021);
and U10297 (N_10297,N_9835,N_9996);
nor U10298 (N_10298,N_10056,N_10125);
and U10299 (N_10299,N_10075,N_9692);
nand U10300 (N_10300,N_10117,N_10082);
nor U10301 (N_10301,N_9853,N_9717);
nor U10302 (N_10302,N_9803,N_10162);
nor U10303 (N_10303,N_9905,N_9603);
nor U10304 (N_10304,N_9749,N_9722);
nor U10305 (N_10305,N_10143,N_10176);
or U10306 (N_10306,N_9657,N_10040);
and U10307 (N_10307,N_9804,N_10137);
xor U10308 (N_10308,N_10099,N_9711);
or U10309 (N_10309,N_9636,N_10169);
nor U10310 (N_10310,N_10173,N_10053);
xnor U10311 (N_10311,N_9800,N_10041);
nand U10312 (N_10312,N_9660,N_9965);
xnor U10313 (N_10313,N_9716,N_9763);
or U10314 (N_10314,N_9667,N_10155);
xnor U10315 (N_10315,N_9681,N_9799);
or U10316 (N_10316,N_10114,N_9726);
and U10317 (N_10317,N_9925,N_9653);
or U10318 (N_10318,N_9897,N_10032);
nand U10319 (N_10319,N_9810,N_9862);
xnor U10320 (N_10320,N_10063,N_9889);
or U10321 (N_10321,N_10126,N_9779);
nor U10322 (N_10322,N_9829,N_10045);
xnor U10323 (N_10323,N_9836,N_9875);
nor U10324 (N_10324,N_10062,N_10168);
nand U10325 (N_10325,N_10121,N_9973);
nand U10326 (N_10326,N_9812,N_9633);
and U10327 (N_10327,N_9611,N_9725);
nor U10328 (N_10328,N_10046,N_10051);
xor U10329 (N_10329,N_9893,N_9651);
xor U10330 (N_10330,N_9634,N_10142);
or U10331 (N_10331,N_10174,N_9891);
or U10332 (N_10332,N_9952,N_9917);
nor U10333 (N_10333,N_9847,N_10179);
xor U10334 (N_10334,N_9757,N_10110);
and U10335 (N_10335,N_10008,N_10129);
and U10336 (N_10336,N_9994,N_9672);
nor U10337 (N_10337,N_9947,N_9936);
nand U10338 (N_10338,N_9985,N_9991);
xnor U10339 (N_10339,N_10080,N_9794);
nand U10340 (N_10340,N_9811,N_9797);
xnor U10341 (N_10341,N_9613,N_9876);
nor U10342 (N_10342,N_9744,N_9935);
nand U10343 (N_10343,N_10183,N_9760);
and U10344 (N_10344,N_9828,N_10123);
nand U10345 (N_10345,N_9968,N_10014);
or U10346 (N_10346,N_9903,N_10068);
or U10347 (N_10347,N_10035,N_9630);
and U10348 (N_10348,N_10003,N_10001);
nand U10349 (N_10349,N_10027,N_9928);
nand U10350 (N_10350,N_9645,N_9964);
or U10351 (N_10351,N_10081,N_9748);
or U10352 (N_10352,N_10096,N_9747);
and U10353 (N_10353,N_9792,N_9988);
nor U10354 (N_10354,N_10091,N_10193);
or U10355 (N_10355,N_9825,N_9999);
or U10356 (N_10356,N_10050,N_10037);
or U10357 (N_10357,N_9953,N_9643);
xnor U10358 (N_10358,N_10039,N_9727);
xor U10359 (N_10359,N_9808,N_10157);
nand U10360 (N_10360,N_9605,N_9659);
xor U10361 (N_10361,N_9849,N_9773);
xor U10362 (N_10362,N_9855,N_9848);
xnor U10363 (N_10363,N_9707,N_10135);
or U10364 (N_10364,N_9600,N_10029);
xnor U10365 (N_10365,N_10150,N_9984);
nor U10366 (N_10366,N_9734,N_9937);
xor U10367 (N_10367,N_9621,N_9837);
nor U10368 (N_10368,N_9663,N_9796);
or U10369 (N_10369,N_9607,N_9728);
xnor U10370 (N_10370,N_10104,N_10097);
and U10371 (N_10371,N_10152,N_9669);
xor U10372 (N_10372,N_10119,N_9904);
nand U10373 (N_10373,N_10089,N_9791);
xnor U10374 (N_10374,N_9759,N_9774);
nand U10375 (N_10375,N_9912,N_10161);
nand U10376 (N_10376,N_9842,N_9608);
xnor U10377 (N_10377,N_9765,N_9833);
xnor U10378 (N_10378,N_9942,N_9822);
and U10379 (N_10379,N_9872,N_9877);
or U10380 (N_10380,N_9735,N_9755);
xnor U10381 (N_10381,N_10175,N_9993);
nand U10382 (N_10382,N_9649,N_9648);
or U10383 (N_10383,N_9752,N_9857);
and U10384 (N_10384,N_9731,N_9995);
and U10385 (N_10385,N_9723,N_9879);
nand U10386 (N_10386,N_9992,N_10191);
and U10387 (N_10387,N_9684,N_9908);
xor U10388 (N_10388,N_9786,N_9816);
xor U10389 (N_10389,N_9656,N_10148);
nor U10390 (N_10390,N_9793,N_9961);
nor U10391 (N_10391,N_10146,N_9650);
or U10392 (N_10392,N_10103,N_10043);
and U10393 (N_10393,N_9967,N_10069);
xor U10394 (N_10394,N_9624,N_9931);
xor U10395 (N_10395,N_10092,N_9933);
nor U10396 (N_10396,N_10130,N_9854);
nand U10397 (N_10397,N_10057,N_9696);
and U10398 (N_10398,N_10088,N_9713);
nor U10399 (N_10399,N_9921,N_9714);
or U10400 (N_10400,N_9635,N_9754);
or U10401 (N_10401,N_9990,N_9982);
and U10402 (N_10402,N_9769,N_9742);
nand U10403 (N_10403,N_9885,N_9927);
nor U10404 (N_10404,N_9658,N_9892);
nor U10405 (N_10405,N_9823,N_9738);
nor U10406 (N_10406,N_9941,N_9675);
xnor U10407 (N_10407,N_9883,N_10195);
and U10408 (N_10408,N_9923,N_9858);
and U10409 (N_10409,N_9978,N_10055);
or U10410 (N_10410,N_9778,N_10128);
and U10411 (N_10411,N_9646,N_9619);
xnor U10412 (N_10412,N_9622,N_10030);
and U10413 (N_10413,N_10023,N_9617);
xor U10414 (N_10414,N_9819,N_9980);
nor U10415 (N_10415,N_10180,N_10133);
and U10416 (N_10416,N_9887,N_10154);
and U10417 (N_10417,N_10022,N_9790);
and U10418 (N_10418,N_9987,N_9604);
or U10419 (N_10419,N_10070,N_10182);
nand U10420 (N_10420,N_10116,N_10187);
xor U10421 (N_10421,N_9719,N_9686);
xor U10422 (N_10422,N_10131,N_10024);
and U10423 (N_10423,N_9873,N_10083);
and U10424 (N_10424,N_9720,N_9626);
xor U10425 (N_10425,N_10184,N_9746);
and U10426 (N_10426,N_9721,N_10020);
or U10427 (N_10427,N_9878,N_9637);
xnor U10428 (N_10428,N_9907,N_9780);
or U10429 (N_10429,N_9951,N_9846);
nor U10430 (N_10430,N_9900,N_9906);
or U10431 (N_10431,N_9983,N_9882);
or U10432 (N_10432,N_9673,N_9976);
nor U10433 (N_10433,N_9868,N_9826);
xor U10434 (N_10434,N_9704,N_9801);
xor U10435 (N_10435,N_9864,N_10192);
nor U10436 (N_10436,N_9929,N_9827);
or U10437 (N_10437,N_9944,N_10181);
nand U10438 (N_10438,N_9918,N_10140);
xor U10439 (N_10439,N_10118,N_10036);
nand U10440 (N_10440,N_10087,N_10064);
xor U10441 (N_10441,N_9817,N_9789);
xor U10442 (N_10442,N_9688,N_9661);
nor U10443 (N_10443,N_9814,N_10090);
nor U10444 (N_10444,N_10073,N_10102);
xor U10445 (N_10445,N_9924,N_9652);
or U10446 (N_10446,N_10038,N_9730);
nor U10447 (N_10447,N_10165,N_9777);
or U10448 (N_10448,N_9664,N_10105);
xor U10449 (N_10449,N_9781,N_10120);
or U10450 (N_10450,N_9609,N_9841);
or U10451 (N_10451,N_9813,N_9956);
nor U10452 (N_10452,N_9960,N_10124);
xnor U10453 (N_10453,N_10044,N_9948);
xnor U10454 (N_10454,N_9655,N_9943);
nor U10455 (N_10455,N_9798,N_9647);
xnor U10456 (N_10456,N_9679,N_9911);
nor U10457 (N_10457,N_9753,N_10196);
or U10458 (N_10458,N_9615,N_9682);
nand U10459 (N_10459,N_10095,N_9831);
and U10460 (N_10460,N_9919,N_10007);
nand U10461 (N_10461,N_10065,N_10000);
nor U10462 (N_10462,N_10139,N_10158);
or U10463 (N_10463,N_10071,N_9997);
xnor U10464 (N_10464,N_9616,N_9638);
and U10465 (N_10465,N_10141,N_9809);
and U10466 (N_10466,N_10132,N_9678);
xnor U10467 (N_10467,N_10172,N_9977);
nand U10468 (N_10468,N_10177,N_9710);
and U10469 (N_10469,N_9767,N_9741);
xnor U10470 (N_10470,N_10093,N_10111);
nor U10471 (N_10471,N_9945,N_9758);
xor U10472 (N_10472,N_9708,N_10094);
nor U10473 (N_10473,N_9998,N_9743);
and U10474 (N_10474,N_10061,N_9718);
and U10475 (N_10475,N_10188,N_10178);
or U10476 (N_10476,N_9740,N_9949);
xnor U10477 (N_10477,N_9729,N_9676);
nor U10478 (N_10478,N_9701,N_9654);
xor U10479 (N_10479,N_9788,N_9899);
nand U10480 (N_10480,N_9938,N_9840);
or U10481 (N_10481,N_9787,N_9894);
nand U10482 (N_10482,N_9910,N_9614);
and U10483 (N_10483,N_10016,N_9666);
and U10484 (N_10484,N_9768,N_10012);
and U10485 (N_10485,N_10054,N_9628);
nor U10486 (N_10486,N_9733,N_9920);
nand U10487 (N_10487,N_10026,N_9736);
or U10488 (N_10488,N_9706,N_9860);
or U10489 (N_10489,N_9909,N_9832);
nor U10490 (N_10490,N_9739,N_9724);
nand U10491 (N_10491,N_9644,N_10019);
nor U10492 (N_10492,N_9930,N_10194);
and U10493 (N_10493,N_10072,N_10017);
nor U10494 (N_10494,N_10052,N_9850);
xor U10495 (N_10495,N_9926,N_9818);
nand U10496 (N_10496,N_9715,N_9859);
or U10497 (N_10497,N_9693,N_9856);
nand U10498 (N_10498,N_9940,N_9975);
nand U10499 (N_10499,N_10076,N_10171);
or U10500 (N_10500,N_9766,N_10179);
nor U10501 (N_10501,N_10090,N_10138);
or U10502 (N_10502,N_9921,N_10096);
and U10503 (N_10503,N_9940,N_9961);
and U10504 (N_10504,N_10020,N_9774);
or U10505 (N_10505,N_9627,N_9863);
xnor U10506 (N_10506,N_10050,N_9914);
and U10507 (N_10507,N_9850,N_9648);
nand U10508 (N_10508,N_9604,N_10120);
and U10509 (N_10509,N_10004,N_10072);
or U10510 (N_10510,N_9621,N_9746);
nor U10511 (N_10511,N_9878,N_9938);
xor U10512 (N_10512,N_10155,N_10021);
xor U10513 (N_10513,N_9678,N_10170);
or U10514 (N_10514,N_9661,N_9604);
xor U10515 (N_10515,N_9975,N_9623);
or U10516 (N_10516,N_9742,N_10068);
nor U10517 (N_10517,N_9907,N_9985);
or U10518 (N_10518,N_9985,N_10138);
and U10519 (N_10519,N_9696,N_9958);
nor U10520 (N_10520,N_9755,N_9732);
and U10521 (N_10521,N_9662,N_10096);
nor U10522 (N_10522,N_10138,N_9936);
xnor U10523 (N_10523,N_9683,N_9827);
xnor U10524 (N_10524,N_10161,N_10104);
nand U10525 (N_10525,N_9731,N_9740);
xor U10526 (N_10526,N_9756,N_10042);
or U10527 (N_10527,N_9994,N_9945);
or U10528 (N_10528,N_10178,N_10190);
nand U10529 (N_10529,N_9997,N_9750);
nand U10530 (N_10530,N_9714,N_10067);
nor U10531 (N_10531,N_10126,N_10144);
nand U10532 (N_10532,N_9900,N_9688);
and U10533 (N_10533,N_9710,N_9604);
or U10534 (N_10534,N_9898,N_10153);
and U10535 (N_10535,N_9802,N_9856);
nand U10536 (N_10536,N_9866,N_9747);
nand U10537 (N_10537,N_9887,N_9988);
or U10538 (N_10538,N_10184,N_10056);
xor U10539 (N_10539,N_10024,N_9678);
xnor U10540 (N_10540,N_9961,N_9729);
xor U10541 (N_10541,N_9684,N_9770);
xor U10542 (N_10542,N_9911,N_9823);
nand U10543 (N_10543,N_9957,N_10015);
or U10544 (N_10544,N_10154,N_9712);
nand U10545 (N_10545,N_9659,N_9926);
and U10546 (N_10546,N_9884,N_9663);
or U10547 (N_10547,N_10183,N_10167);
nand U10548 (N_10548,N_9615,N_9987);
nand U10549 (N_10549,N_10131,N_10173);
and U10550 (N_10550,N_9738,N_9602);
and U10551 (N_10551,N_9615,N_9966);
or U10552 (N_10552,N_10068,N_9690);
xor U10553 (N_10553,N_9818,N_9948);
and U10554 (N_10554,N_10097,N_9779);
xor U10555 (N_10555,N_9705,N_9783);
nand U10556 (N_10556,N_9707,N_10058);
nor U10557 (N_10557,N_9737,N_10187);
xnor U10558 (N_10558,N_9931,N_9747);
nor U10559 (N_10559,N_9881,N_9656);
nand U10560 (N_10560,N_10172,N_10115);
and U10561 (N_10561,N_10063,N_9662);
nand U10562 (N_10562,N_10114,N_10090);
nor U10563 (N_10563,N_9750,N_9882);
and U10564 (N_10564,N_9741,N_10174);
nand U10565 (N_10565,N_9614,N_9911);
or U10566 (N_10566,N_9919,N_10127);
and U10567 (N_10567,N_9895,N_9722);
and U10568 (N_10568,N_9783,N_10065);
nor U10569 (N_10569,N_9733,N_9653);
and U10570 (N_10570,N_9873,N_9672);
nand U10571 (N_10571,N_9770,N_9935);
or U10572 (N_10572,N_10067,N_10131);
nand U10573 (N_10573,N_9859,N_9888);
nor U10574 (N_10574,N_9977,N_9747);
nand U10575 (N_10575,N_9998,N_9794);
nand U10576 (N_10576,N_9848,N_9791);
xor U10577 (N_10577,N_9782,N_10108);
xnor U10578 (N_10578,N_10027,N_9948);
and U10579 (N_10579,N_9678,N_9832);
nand U10580 (N_10580,N_10087,N_9648);
nand U10581 (N_10581,N_9815,N_9775);
nand U10582 (N_10582,N_9713,N_9700);
xor U10583 (N_10583,N_10170,N_9916);
xor U10584 (N_10584,N_10044,N_9903);
and U10585 (N_10585,N_9952,N_9941);
nand U10586 (N_10586,N_9784,N_10011);
or U10587 (N_10587,N_9868,N_9629);
and U10588 (N_10588,N_9964,N_10102);
nand U10589 (N_10589,N_9632,N_9682);
nand U10590 (N_10590,N_9696,N_10073);
or U10591 (N_10591,N_9828,N_10039);
and U10592 (N_10592,N_9659,N_9890);
nor U10593 (N_10593,N_9771,N_9806);
and U10594 (N_10594,N_9792,N_9935);
nor U10595 (N_10595,N_9942,N_9605);
nand U10596 (N_10596,N_9820,N_9621);
and U10597 (N_10597,N_9618,N_10117);
and U10598 (N_10598,N_9838,N_9859);
nand U10599 (N_10599,N_9810,N_10059);
nor U10600 (N_10600,N_10062,N_9788);
xnor U10601 (N_10601,N_9625,N_9853);
and U10602 (N_10602,N_9780,N_9929);
xnor U10603 (N_10603,N_9807,N_10167);
or U10604 (N_10604,N_10070,N_9982);
and U10605 (N_10605,N_9838,N_9908);
xnor U10606 (N_10606,N_10118,N_10046);
xor U10607 (N_10607,N_9711,N_9934);
or U10608 (N_10608,N_10093,N_9883);
nand U10609 (N_10609,N_10135,N_10141);
nand U10610 (N_10610,N_10069,N_10176);
or U10611 (N_10611,N_10111,N_9815);
and U10612 (N_10612,N_9671,N_9757);
nand U10613 (N_10613,N_9905,N_9703);
nor U10614 (N_10614,N_9696,N_10192);
xor U10615 (N_10615,N_10012,N_9805);
or U10616 (N_10616,N_9885,N_9960);
nor U10617 (N_10617,N_10084,N_9850);
and U10618 (N_10618,N_9712,N_9845);
or U10619 (N_10619,N_10093,N_9865);
nand U10620 (N_10620,N_10033,N_9710);
and U10621 (N_10621,N_9765,N_9971);
xnor U10622 (N_10622,N_9828,N_10047);
and U10623 (N_10623,N_9745,N_10111);
nor U10624 (N_10624,N_9916,N_10137);
nand U10625 (N_10625,N_9698,N_9791);
or U10626 (N_10626,N_9974,N_9858);
and U10627 (N_10627,N_10175,N_9815);
nor U10628 (N_10628,N_9926,N_10110);
nor U10629 (N_10629,N_10187,N_9991);
nor U10630 (N_10630,N_9706,N_10019);
and U10631 (N_10631,N_9734,N_10139);
and U10632 (N_10632,N_9659,N_10137);
xnor U10633 (N_10633,N_9954,N_10092);
nor U10634 (N_10634,N_9614,N_9698);
or U10635 (N_10635,N_10106,N_9600);
nand U10636 (N_10636,N_9784,N_9630);
xor U10637 (N_10637,N_10038,N_9804);
and U10638 (N_10638,N_9749,N_10090);
nand U10639 (N_10639,N_9841,N_10112);
nand U10640 (N_10640,N_9831,N_9736);
xnor U10641 (N_10641,N_9703,N_9859);
xor U10642 (N_10642,N_10126,N_9618);
xor U10643 (N_10643,N_10060,N_9795);
and U10644 (N_10644,N_10041,N_10147);
and U10645 (N_10645,N_9742,N_10101);
or U10646 (N_10646,N_9818,N_10073);
and U10647 (N_10647,N_9992,N_10074);
and U10648 (N_10648,N_9899,N_10143);
and U10649 (N_10649,N_10052,N_10026);
xor U10650 (N_10650,N_9647,N_10008);
xnor U10651 (N_10651,N_10012,N_9670);
or U10652 (N_10652,N_9675,N_9850);
xnor U10653 (N_10653,N_9804,N_9822);
and U10654 (N_10654,N_9761,N_9814);
or U10655 (N_10655,N_10115,N_9751);
xnor U10656 (N_10656,N_10190,N_9924);
nand U10657 (N_10657,N_9697,N_9991);
and U10658 (N_10658,N_9987,N_9789);
or U10659 (N_10659,N_10085,N_9614);
nand U10660 (N_10660,N_9937,N_10137);
nand U10661 (N_10661,N_9744,N_10034);
and U10662 (N_10662,N_9930,N_9721);
nand U10663 (N_10663,N_10026,N_9820);
or U10664 (N_10664,N_10106,N_9735);
nand U10665 (N_10665,N_10043,N_9830);
nor U10666 (N_10666,N_9772,N_10121);
nand U10667 (N_10667,N_9772,N_9935);
xnor U10668 (N_10668,N_9971,N_9726);
nand U10669 (N_10669,N_10149,N_9652);
nand U10670 (N_10670,N_9900,N_10039);
nand U10671 (N_10671,N_9704,N_10020);
nor U10672 (N_10672,N_9739,N_9740);
nand U10673 (N_10673,N_9837,N_10083);
and U10674 (N_10674,N_9885,N_9956);
nand U10675 (N_10675,N_10110,N_9664);
nand U10676 (N_10676,N_10083,N_10124);
nand U10677 (N_10677,N_9612,N_9665);
or U10678 (N_10678,N_10135,N_9847);
and U10679 (N_10679,N_9997,N_9757);
or U10680 (N_10680,N_10144,N_9891);
and U10681 (N_10681,N_10164,N_10166);
xnor U10682 (N_10682,N_10086,N_9947);
nand U10683 (N_10683,N_9986,N_9827);
nand U10684 (N_10684,N_10149,N_9951);
xnor U10685 (N_10685,N_10085,N_9823);
and U10686 (N_10686,N_9734,N_10177);
and U10687 (N_10687,N_9811,N_10046);
or U10688 (N_10688,N_9625,N_9824);
or U10689 (N_10689,N_9970,N_9633);
xnor U10690 (N_10690,N_9780,N_9804);
or U10691 (N_10691,N_9814,N_9635);
nor U10692 (N_10692,N_9823,N_9910);
and U10693 (N_10693,N_9702,N_10013);
nor U10694 (N_10694,N_9607,N_9709);
xor U10695 (N_10695,N_9722,N_10121);
nand U10696 (N_10696,N_10160,N_9608);
or U10697 (N_10697,N_10115,N_10031);
and U10698 (N_10698,N_9969,N_9881);
nand U10699 (N_10699,N_9784,N_9827);
and U10700 (N_10700,N_9947,N_9901);
nand U10701 (N_10701,N_9933,N_9628);
nor U10702 (N_10702,N_9746,N_10147);
xor U10703 (N_10703,N_9866,N_9625);
or U10704 (N_10704,N_9713,N_9727);
and U10705 (N_10705,N_9900,N_10065);
xnor U10706 (N_10706,N_9978,N_9716);
or U10707 (N_10707,N_9864,N_9811);
nor U10708 (N_10708,N_10029,N_9879);
or U10709 (N_10709,N_9857,N_9928);
or U10710 (N_10710,N_9675,N_10149);
nor U10711 (N_10711,N_10017,N_10028);
and U10712 (N_10712,N_9764,N_9731);
nor U10713 (N_10713,N_10025,N_9831);
and U10714 (N_10714,N_10078,N_10146);
and U10715 (N_10715,N_9733,N_9896);
nor U10716 (N_10716,N_9971,N_9869);
or U10717 (N_10717,N_9872,N_9644);
nor U10718 (N_10718,N_9993,N_9648);
nand U10719 (N_10719,N_9802,N_10011);
or U10720 (N_10720,N_9872,N_9604);
nor U10721 (N_10721,N_10000,N_10167);
xnor U10722 (N_10722,N_9948,N_9940);
or U10723 (N_10723,N_10128,N_10193);
nand U10724 (N_10724,N_9802,N_9859);
and U10725 (N_10725,N_10125,N_10098);
and U10726 (N_10726,N_9818,N_10090);
nand U10727 (N_10727,N_9632,N_10115);
nand U10728 (N_10728,N_10149,N_10089);
or U10729 (N_10729,N_9951,N_9791);
nand U10730 (N_10730,N_9627,N_10073);
xnor U10731 (N_10731,N_9860,N_10100);
and U10732 (N_10732,N_9627,N_10076);
nand U10733 (N_10733,N_9772,N_9950);
xor U10734 (N_10734,N_10078,N_10111);
nor U10735 (N_10735,N_10153,N_10038);
xor U10736 (N_10736,N_9917,N_10130);
nand U10737 (N_10737,N_9716,N_9929);
nand U10738 (N_10738,N_9841,N_9791);
nor U10739 (N_10739,N_10169,N_9930);
xnor U10740 (N_10740,N_9769,N_10057);
nand U10741 (N_10741,N_10079,N_10093);
nand U10742 (N_10742,N_9769,N_9743);
nor U10743 (N_10743,N_9874,N_9777);
or U10744 (N_10744,N_10030,N_9923);
nor U10745 (N_10745,N_9871,N_9686);
xor U10746 (N_10746,N_9980,N_10136);
or U10747 (N_10747,N_9875,N_10135);
xor U10748 (N_10748,N_9692,N_10054);
and U10749 (N_10749,N_9981,N_9609);
and U10750 (N_10750,N_9852,N_9753);
or U10751 (N_10751,N_9831,N_9615);
xor U10752 (N_10752,N_9782,N_10129);
or U10753 (N_10753,N_10163,N_9772);
nand U10754 (N_10754,N_9690,N_9781);
or U10755 (N_10755,N_10023,N_10158);
nor U10756 (N_10756,N_10009,N_9656);
and U10757 (N_10757,N_9884,N_10009);
or U10758 (N_10758,N_10097,N_10026);
nor U10759 (N_10759,N_9737,N_10144);
xor U10760 (N_10760,N_9793,N_9887);
nand U10761 (N_10761,N_9750,N_9611);
and U10762 (N_10762,N_9627,N_10017);
nand U10763 (N_10763,N_9925,N_9961);
nand U10764 (N_10764,N_9908,N_10189);
xor U10765 (N_10765,N_9824,N_10169);
xor U10766 (N_10766,N_10163,N_9618);
xnor U10767 (N_10767,N_9992,N_10179);
and U10768 (N_10768,N_10157,N_10167);
xor U10769 (N_10769,N_10036,N_10156);
nor U10770 (N_10770,N_9992,N_9798);
xnor U10771 (N_10771,N_9604,N_9748);
nand U10772 (N_10772,N_9789,N_9634);
and U10773 (N_10773,N_9740,N_10026);
nand U10774 (N_10774,N_9949,N_10062);
nor U10775 (N_10775,N_10170,N_9682);
xnor U10776 (N_10776,N_9832,N_9808);
nor U10777 (N_10777,N_10067,N_10197);
nor U10778 (N_10778,N_9825,N_10121);
nor U10779 (N_10779,N_10175,N_9984);
xor U10780 (N_10780,N_9923,N_9849);
nand U10781 (N_10781,N_9604,N_10041);
nor U10782 (N_10782,N_9824,N_9799);
or U10783 (N_10783,N_10183,N_9720);
xor U10784 (N_10784,N_9761,N_10183);
or U10785 (N_10785,N_10105,N_10026);
and U10786 (N_10786,N_9637,N_9923);
xor U10787 (N_10787,N_9774,N_9985);
nand U10788 (N_10788,N_9971,N_10072);
or U10789 (N_10789,N_9911,N_10047);
and U10790 (N_10790,N_9644,N_10181);
xor U10791 (N_10791,N_10128,N_9901);
or U10792 (N_10792,N_10124,N_9902);
nand U10793 (N_10793,N_9938,N_10141);
nand U10794 (N_10794,N_9908,N_10185);
or U10795 (N_10795,N_9642,N_9668);
nand U10796 (N_10796,N_9877,N_10149);
and U10797 (N_10797,N_9845,N_9630);
nand U10798 (N_10798,N_10063,N_9874);
nor U10799 (N_10799,N_9946,N_10007);
xor U10800 (N_10800,N_10677,N_10374);
or U10801 (N_10801,N_10503,N_10464);
and U10802 (N_10802,N_10550,N_10349);
nand U10803 (N_10803,N_10473,N_10461);
and U10804 (N_10804,N_10277,N_10208);
or U10805 (N_10805,N_10331,N_10292);
nor U10806 (N_10806,N_10584,N_10565);
nor U10807 (N_10807,N_10325,N_10211);
nor U10808 (N_10808,N_10476,N_10674);
nand U10809 (N_10809,N_10704,N_10434);
nand U10810 (N_10810,N_10749,N_10221);
nand U10811 (N_10811,N_10556,N_10533);
nor U10812 (N_10812,N_10306,N_10387);
nor U10813 (N_10813,N_10781,N_10265);
and U10814 (N_10814,N_10239,N_10611);
xnor U10815 (N_10815,N_10564,N_10339);
nand U10816 (N_10816,N_10701,N_10432);
and U10817 (N_10817,N_10559,N_10517);
xnor U10818 (N_10818,N_10435,N_10290);
and U10819 (N_10819,N_10684,N_10402);
xnor U10820 (N_10820,N_10705,N_10694);
and U10821 (N_10821,N_10596,N_10735);
and U10822 (N_10822,N_10445,N_10593);
xnor U10823 (N_10823,N_10516,N_10602);
or U10824 (N_10824,N_10351,N_10238);
nand U10825 (N_10825,N_10377,N_10577);
nand U10826 (N_10826,N_10285,N_10532);
xor U10827 (N_10827,N_10304,N_10367);
xor U10828 (N_10828,N_10608,N_10469);
nand U10829 (N_10829,N_10569,N_10723);
and U10830 (N_10830,N_10686,N_10336);
and U10831 (N_10831,N_10798,N_10530);
nor U10832 (N_10832,N_10715,N_10787);
xnor U10833 (N_10833,N_10284,N_10629);
nand U10834 (N_10834,N_10606,N_10492);
and U10835 (N_10835,N_10248,N_10386);
or U10836 (N_10836,N_10460,N_10352);
xnor U10837 (N_10837,N_10465,N_10499);
and U10838 (N_10838,N_10744,N_10310);
or U10839 (N_10839,N_10784,N_10390);
or U10840 (N_10840,N_10298,N_10441);
nor U10841 (N_10841,N_10363,N_10706);
nor U10842 (N_10842,N_10515,N_10630);
or U10843 (N_10843,N_10718,N_10250);
nor U10844 (N_10844,N_10538,N_10741);
xnor U10845 (N_10845,N_10586,N_10685);
xnor U10846 (N_10846,N_10788,N_10202);
xor U10847 (N_10847,N_10578,N_10682);
nand U10848 (N_10848,N_10262,N_10266);
and U10849 (N_10849,N_10734,N_10431);
xor U10850 (N_10850,N_10338,N_10257);
xor U10851 (N_10851,N_10279,N_10603);
nor U10852 (N_10852,N_10254,N_10716);
and U10853 (N_10853,N_10496,N_10767);
xnor U10854 (N_10854,N_10411,N_10612);
or U10855 (N_10855,N_10752,N_10378);
and U10856 (N_10856,N_10635,N_10521);
or U10857 (N_10857,N_10703,N_10348);
or U10858 (N_10858,N_10796,N_10407);
nand U10859 (N_10859,N_10406,N_10536);
nor U10860 (N_10860,N_10247,N_10707);
or U10861 (N_10861,N_10779,N_10452);
nor U10862 (N_10862,N_10592,N_10637);
or U10863 (N_10863,N_10664,N_10625);
or U10864 (N_10864,N_10678,N_10252);
nor U10865 (N_10865,N_10563,N_10772);
xnor U10866 (N_10866,N_10655,N_10327);
xnor U10867 (N_10867,N_10324,N_10750);
and U10868 (N_10868,N_10646,N_10360);
xnor U10869 (N_10869,N_10769,N_10792);
nor U10870 (N_10870,N_10361,N_10332);
and U10871 (N_10871,N_10708,N_10766);
nor U10872 (N_10872,N_10307,N_10448);
and U10873 (N_10873,N_10553,N_10401);
nand U10874 (N_10874,N_10757,N_10312);
nand U10875 (N_10875,N_10218,N_10638);
nor U10876 (N_10876,N_10580,N_10626);
xnor U10877 (N_10877,N_10233,N_10690);
and U10878 (N_10878,N_10234,N_10366);
xnor U10879 (N_10879,N_10249,N_10283);
nor U10880 (N_10880,N_10620,N_10313);
and U10881 (N_10881,N_10719,N_10730);
or U10882 (N_10882,N_10791,N_10692);
nor U10883 (N_10883,N_10342,N_10617);
nand U10884 (N_10884,N_10486,N_10300);
nor U10885 (N_10885,N_10227,N_10455);
and U10886 (N_10886,N_10551,N_10599);
nand U10887 (N_10887,N_10272,N_10573);
or U10888 (N_10888,N_10729,N_10774);
or U10889 (N_10889,N_10627,N_10241);
nand U10890 (N_10890,N_10797,N_10299);
nor U10891 (N_10891,N_10665,N_10511);
nor U10892 (N_10892,N_10699,N_10246);
xor U10893 (N_10893,N_10598,N_10588);
xnor U10894 (N_10894,N_10333,N_10673);
or U10895 (N_10895,N_10418,N_10437);
nor U10896 (N_10896,N_10489,N_10373);
xor U10897 (N_10897,N_10264,N_10323);
nand U10898 (N_10898,N_10380,N_10205);
xnor U10899 (N_10899,N_10451,N_10540);
xor U10900 (N_10900,N_10488,N_10354);
nor U10901 (N_10901,N_10413,N_10255);
nand U10902 (N_10902,N_10760,N_10656);
or U10903 (N_10903,N_10364,N_10459);
nor U10904 (N_10904,N_10442,N_10326);
or U10905 (N_10905,N_10773,N_10243);
nor U10906 (N_10906,N_10423,N_10547);
nand U10907 (N_10907,N_10281,N_10231);
or U10908 (N_10908,N_10616,N_10793);
xor U10909 (N_10909,N_10543,N_10375);
and U10910 (N_10910,N_10725,N_10581);
or U10911 (N_10911,N_10383,N_10671);
xor U10912 (N_10912,N_10585,N_10320);
nand U10913 (N_10913,N_10397,N_10275);
xor U10914 (N_10914,N_10764,N_10237);
xnor U10915 (N_10915,N_10739,N_10783);
nor U10916 (N_10916,N_10650,N_10615);
or U10917 (N_10917,N_10661,N_10724);
xor U10918 (N_10918,N_10462,N_10263);
nand U10919 (N_10919,N_10557,N_10681);
nor U10920 (N_10920,N_10754,N_10355);
xnor U10921 (N_10921,N_10583,N_10537);
nand U10922 (N_10922,N_10356,N_10698);
and U10923 (N_10923,N_10427,N_10329);
xnor U10924 (N_10924,N_10645,N_10649);
nor U10925 (N_10925,N_10498,N_10371);
nand U10926 (N_10926,N_10634,N_10415);
nor U10927 (N_10927,N_10605,N_10315);
xnor U10928 (N_10928,N_10412,N_10497);
or U10929 (N_10929,N_10341,N_10506);
nand U10930 (N_10930,N_10711,N_10381);
nand U10931 (N_10931,N_10222,N_10505);
or U10932 (N_10932,N_10353,N_10544);
nor U10933 (N_10933,N_10282,N_10491);
nand U10934 (N_10934,N_10509,N_10370);
or U10935 (N_10935,N_10523,N_10269);
and U10936 (N_10936,N_10662,N_10225);
nand U10937 (N_10937,N_10676,N_10301);
nor U10938 (N_10938,N_10242,N_10235);
or U10939 (N_10939,N_10785,N_10429);
nor U10940 (N_10940,N_10405,N_10641);
nor U10941 (N_10941,N_10500,N_10594);
or U10942 (N_10942,N_10474,N_10765);
nor U10943 (N_10943,N_10410,N_10552);
nand U10944 (N_10944,N_10293,N_10542);
nor U10945 (N_10945,N_10520,N_10228);
and U10946 (N_10946,N_10261,N_10314);
nor U10947 (N_10947,N_10396,N_10574);
nor U10948 (N_10948,N_10663,N_10270);
nand U10949 (N_10949,N_10288,N_10504);
nor U10950 (N_10950,N_10549,N_10591);
xor U10951 (N_10951,N_10382,N_10527);
or U10952 (N_10952,N_10771,N_10691);
xor U10953 (N_10953,N_10713,N_10748);
and U10954 (N_10954,N_10369,N_10541);
or U10955 (N_10955,N_10394,N_10717);
and U10956 (N_10956,N_10278,N_10659);
nand U10957 (N_10957,N_10642,N_10346);
and U10958 (N_10958,N_10693,N_10660);
nor U10959 (N_10959,N_10514,N_10319);
xor U10960 (N_10960,N_10466,N_10669);
nand U10961 (N_10961,N_10291,N_10482);
nand U10962 (N_10962,N_10675,N_10762);
and U10963 (N_10963,N_10420,N_10738);
and U10964 (N_10964,N_10294,N_10614);
or U10965 (N_10965,N_10654,N_10359);
and U10966 (N_10966,N_10484,N_10778);
nand U10967 (N_10967,N_10575,N_10385);
nor U10968 (N_10968,N_10695,N_10732);
or U10969 (N_10969,N_10216,N_10350);
and U10970 (N_10970,N_10643,N_10518);
nand U10971 (N_10971,N_10740,N_10444);
or U10972 (N_10972,N_10733,N_10624);
and U10973 (N_10973,N_10322,N_10622);
xor U10974 (N_10974,N_10493,N_10404);
nor U10975 (N_10975,N_10430,N_10582);
nand U10976 (N_10976,N_10204,N_10728);
nand U10977 (N_10977,N_10276,N_10609);
and U10978 (N_10978,N_10274,N_10389);
and U10979 (N_10979,N_10309,N_10790);
and U10980 (N_10980,N_10416,N_10560);
or U10981 (N_10981,N_10742,N_10480);
or U10982 (N_10982,N_10758,N_10494);
xor U10983 (N_10983,N_10590,N_10226);
nor U10984 (N_10984,N_10207,N_10528);
nand U10985 (N_10985,N_10457,N_10631);
nand U10986 (N_10986,N_10456,N_10513);
nor U10987 (N_10987,N_10311,N_10251);
or U10988 (N_10988,N_10539,N_10534);
nand U10989 (N_10989,N_10731,N_10743);
nand U10990 (N_10990,N_10794,N_10700);
nand U10991 (N_10991,N_10424,N_10328);
or U10992 (N_10992,N_10502,N_10720);
nand U10993 (N_10993,N_10510,N_10756);
and U10994 (N_10994,N_10621,N_10570);
nand U10995 (N_10995,N_10408,N_10712);
or U10996 (N_10996,N_10316,N_10613);
xnor U10997 (N_10997,N_10321,N_10240);
nor U10998 (N_10998,N_10368,N_10362);
xor U10999 (N_10999,N_10303,N_10524);
nand U11000 (N_11000,N_10213,N_10253);
and U11001 (N_11001,N_10260,N_10400);
nand U11002 (N_11002,N_10343,N_10618);
nand U11003 (N_11003,N_10280,N_10286);
or U11004 (N_11004,N_10666,N_10210);
nand U11005 (N_11005,N_10639,N_10597);
xor U11006 (N_11006,N_10463,N_10628);
nand U11007 (N_11007,N_10753,N_10212);
xnor U11008 (N_11008,N_10232,N_10289);
or U11009 (N_11009,N_10443,N_10376);
nand U11010 (N_11010,N_10670,N_10347);
nor U11011 (N_11011,N_10722,N_10688);
nand U11012 (N_11012,N_10714,N_10372);
and U11013 (N_11013,N_10651,N_10633);
or U11014 (N_11014,N_10214,N_10230);
xnor U11015 (N_11015,N_10640,N_10782);
and U11016 (N_11016,N_10483,N_10571);
and U11017 (N_11017,N_10317,N_10558);
nor U11018 (N_11018,N_10726,N_10657);
and U11019 (N_11019,N_10220,N_10258);
nor U11020 (N_11020,N_10679,N_10710);
xor U11021 (N_11021,N_10422,N_10330);
or U11022 (N_11022,N_10302,N_10653);
or U11023 (N_11023,N_10721,N_10409);
nand U11024 (N_11024,N_10395,N_10697);
nand U11025 (N_11025,N_10403,N_10644);
or U11026 (N_11026,N_10799,N_10689);
nor U11027 (N_11027,N_10295,N_10548);
and U11028 (N_11028,N_10229,N_10224);
xor U11029 (N_11029,N_10471,N_10450);
xor U11030 (N_11030,N_10296,N_10759);
or U11031 (N_11031,N_10393,N_10776);
and U11032 (N_11032,N_10454,N_10398);
nand U11033 (N_11033,N_10522,N_10485);
nor U11034 (N_11034,N_10702,N_10334);
nor U11035 (N_11035,N_10428,N_10271);
nor U11036 (N_11036,N_10391,N_10223);
nor U11037 (N_11037,N_10206,N_10217);
nand U11038 (N_11038,N_10267,N_10259);
or U11039 (N_11039,N_10417,N_10297);
or U11040 (N_11040,N_10425,N_10399);
nor U11041 (N_11041,N_10388,N_10467);
nor U11042 (N_11042,N_10576,N_10786);
and U11043 (N_11043,N_10268,N_10636);
xnor U11044 (N_11044,N_10554,N_10392);
nor U11045 (N_11045,N_10607,N_10379);
or U11046 (N_11046,N_10438,N_10236);
nor U11047 (N_11047,N_10453,N_10209);
nor U11048 (N_11048,N_10495,N_10421);
or U11049 (N_11049,N_10273,N_10668);
or U11050 (N_11050,N_10648,N_10357);
nand U11051 (N_11051,N_10755,N_10414);
nand U11052 (N_11052,N_10696,N_10305);
or U11053 (N_11053,N_10795,N_10439);
nor U11054 (N_11054,N_10545,N_10610);
nor U11055 (N_11055,N_10487,N_10761);
nand U11056 (N_11056,N_10589,N_10751);
or U11057 (N_11057,N_10318,N_10344);
nand U11058 (N_11058,N_10587,N_10470);
nand U11059 (N_11059,N_10619,N_10763);
and U11060 (N_11060,N_10426,N_10479);
xor U11061 (N_11061,N_10365,N_10680);
nor U11062 (N_11062,N_10436,N_10475);
nand U11063 (N_11063,N_10245,N_10531);
or U11064 (N_11064,N_10632,N_10308);
xnor U11065 (N_11065,N_10478,N_10358);
and U11066 (N_11066,N_10440,N_10604);
nor U11067 (N_11067,N_10468,N_10561);
or U11068 (N_11068,N_10709,N_10472);
and U11069 (N_11069,N_10525,N_10746);
nand U11070 (N_11070,N_10770,N_10340);
and U11071 (N_11071,N_10449,N_10203);
or U11072 (N_11072,N_10447,N_10745);
nor U11073 (N_11073,N_10683,N_10477);
xor U11074 (N_11074,N_10579,N_10652);
nor U11075 (N_11075,N_10287,N_10244);
xnor U11076 (N_11076,N_10384,N_10419);
nor U11077 (N_11077,N_10658,N_10727);
xor U11078 (N_11078,N_10775,N_10667);
nor U11079 (N_11079,N_10512,N_10595);
nand U11080 (N_11080,N_10623,N_10768);
and U11081 (N_11081,N_10546,N_10535);
nand U11082 (N_11082,N_10736,N_10777);
xnor U11083 (N_11083,N_10555,N_10507);
and U11084 (N_11084,N_10215,N_10337);
nor U11085 (N_11085,N_10200,N_10737);
xor U11086 (N_11086,N_10562,N_10335);
or U11087 (N_11087,N_10256,N_10481);
xor U11088 (N_11088,N_10201,N_10672);
nand U11089 (N_11089,N_10529,N_10572);
xor U11090 (N_11090,N_10501,N_10687);
and U11091 (N_11091,N_10446,N_10647);
xnor U11092 (N_11092,N_10219,N_10526);
and U11093 (N_11093,N_10508,N_10789);
xor U11094 (N_11094,N_10567,N_10747);
nor U11095 (N_11095,N_10433,N_10566);
xor U11096 (N_11096,N_10490,N_10568);
nand U11097 (N_11097,N_10601,N_10519);
xor U11098 (N_11098,N_10458,N_10600);
xor U11099 (N_11099,N_10345,N_10780);
and U11100 (N_11100,N_10729,N_10674);
nand U11101 (N_11101,N_10333,N_10620);
xnor U11102 (N_11102,N_10411,N_10610);
or U11103 (N_11103,N_10344,N_10323);
nand U11104 (N_11104,N_10373,N_10628);
or U11105 (N_11105,N_10778,N_10413);
and U11106 (N_11106,N_10244,N_10681);
xnor U11107 (N_11107,N_10278,N_10723);
or U11108 (N_11108,N_10648,N_10780);
or U11109 (N_11109,N_10301,N_10450);
nand U11110 (N_11110,N_10770,N_10471);
nor U11111 (N_11111,N_10571,N_10549);
nor U11112 (N_11112,N_10564,N_10433);
nand U11113 (N_11113,N_10716,N_10294);
nor U11114 (N_11114,N_10506,N_10373);
and U11115 (N_11115,N_10260,N_10291);
and U11116 (N_11116,N_10665,N_10316);
nand U11117 (N_11117,N_10216,N_10662);
and U11118 (N_11118,N_10706,N_10442);
nor U11119 (N_11119,N_10394,N_10446);
nor U11120 (N_11120,N_10344,N_10698);
nand U11121 (N_11121,N_10532,N_10421);
nor U11122 (N_11122,N_10692,N_10652);
or U11123 (N_11123,N_10533,N_10515);
xnor U11124 (N_11124,N_10440,N_10459);
and U11125 (N_11125,N_10626,N_10326);
nor U11126 (N_11126,N_10632,N_10716);
nor U11127 (N_11127,N_10510,N_10757);
xnor U11128 (N_11128,N_10778,N_10365);
or U11129 (N_11129,N_10748,N_10676);
or U11130 (N_11130,N_10428,N_10628);
or U11131 (N_11131,N_10505,N_10502);
and U11132 (N_11132,N_10556,N_10545);
nand U11133 (N_11133,N_10796,N_10266);
xor U11134 (N_11134,N_10749,N_10249);
nand U11135 (N_11135,N_10736,N_10455);
or U11136 (N_11136,N_10363,N_10521);
and U11137 (N_11137,N_10588,N_10624);
nand U11138 (N_11138,N_10554,N_10715);
nor U11139 (N_11139,N_10267,N_10657);
xnor U11140 (N_11140,N_10762,N_10221);
nor U11141 (N_11141,N_10550,N_10501);
nor U11142 (N_11142,N_10510,N_10780);
and U11143 (N_11143,N_10241,N_10323);
or U11144 (N_11144,N_10313,N_10251);
or U11145 (N_11145,N_10538,N_10674);
or U11146 (N_11146,N_10365,N_10468);
xor U11147 (N_11147,N_10308,N_10252);
nor U11148 (N_11148,N_10301,N_10325);
nand U11149 (N_11149,N_10689,N_10254);
and U11150 (N_11150,N_10306,N_10460);
xnor U11151 (N_11151,N_10268,N_10202);
or U11152 (N_11152,N_10261,N_10750);
nor U11153 (N_11153,N_10662,N_10249);
nor U11154 (N_11154,N_10363,N_10344);
and U11155 (N_11155,N_10323,N_10233);
nand U11156 (N_11156,N_10330,N_10487);
or U11157 (N_11157,N_10747,N_10308);
nand U11158 (N_11158,N_10586,N_10200);
nor U11159 (N_11159,N_10641,N_10595);
nand U11160 (N_11160,N_10545,N_10595);
and U11161 (N_11161,N_10531,N_10298);
or U11162 (N_11162,N_10590,N_10558);
xnor U11163 (N_11163,N_10238,N_10410);
xor U11164 (N_11164,N_10369,N_10263);
xnor U11165 (N_11165,N_10221,N_10368);
and U11166 (N_11166,N_10222,N_10438);
and U11167 (N_11167,N_10467,N_10600);
nor U11168 (N_11168,N_10737,N_10525);
xnor U11169 (N_11169,N_10202,N_10780);
and U11170 (N_11170,N_10507,N_10584);
or U11171 (N_11171,N_10271,N_10287);
and U11172 (N_11172,N_10567,N_10474);
and U11173 (N_11173,N_10430,N_10521);
xor U11174 (N_11174,N_10591,N_10536);
and U11175 (N_11175,N_10284,N_10289);
or U11176 (N_11176,N_10330,N_10728);
nand U11177 (N_11177,N_10749,N_10519);
or U11178 (N_11178,N_10331,N_10743);
and U11179 (N_11179,N_10521,N_10416);
and U11180 (N_11180,N_10560,N_10739);
or U11181 (N_11181,N_10698,N_10420);
xnor U11182 (N_11182,N_10664,N_10348);
nand U11183 (N_11183,N_10702,N_10635);
and U11184 (N_11184,N_10671,N_10725);
nor U11185 (N_11185,N_10488,N_10244);
xor U11186 (N_11186,N_10308,N_10690);
or U11187 (N_11187,N_10320,N_10733);
nand U11188 (N_11188,N_10687,N_10554);
or U11189 (N_11189,N_10501,N_10209);
xor U11190 (N_11190,N_10437,N_10535);
or U11191 (N_11191,N_10556,N_10668);
and U11192 (N_11192,N_10334,N_10514);
xnor U11193 (N_11193,N_10751,N_10417);
nor U11194 (N_11194,N_10577,N_10235);
or U11195 (N_11195,N_10612,N_10340);
nor U11196 (N_11196,N_10282,N_10576);
and U11197 (N_11197,N_10382,N_10234);
or U11198 (N_11198,N_10361,N_10683);
xnor U11199 (N_11199,N_10416,N_10780);
xor U11200 (N_11200,N_10314,N_10357);
nor U11201 (N_11201,N_10280,N_10766);
and U11202 (N_11202,N_10786,N_10794);
and U11203 (N_11203,N_10486,N_10720);
nor U11204 (N_11204,N_10534,N_10414);
nor U11205 (N_11205,N_10486,N_10562);
xnor U11206 (N_11206,N_10472,N_10389);
nand U11207 (N_11207,N_10408,N_10662);
nand U11208 (N_11208,N_10590,N_10560);
nand U11209 (N_11209,N_10458,N_10753);
nor U11210 (N_11210,N_10415,N_10787);
xnor U11211 (N_11211,N_10716,N_10779);
and U11212 (N_11212,N_10730,N_10452);
nand U11213 (N_11213,N_10501,N_10625);
xnor U11214 (N_11214,N_10559,N_10633);
xor U11215 (N_11215,N_10308,N_10241);
and U11216 (N_11216,N_10557,N_10692);
or U11217 (N_11217,N_10574,N_10648);
or U11218 (N_11218,N_10609,N_10659);
and U11219 (N_11219,N_10639,N_10582);
xnor U11220 (N_11220,N_10332,N_10735);
nand U11221 (N_11221,N_10775,N_10483);
and U11222 (N_11222,N_10497,N_10685);
nand U11223 (N_11223,N_10492,N_10425);
or U11224 (N_11224,N_10713,N_10451);
nor U11225 (N_11225,N_10763,N_10414);
and U11226 (N_11226,N_10353,N_10463);
and U11227 (N_11227,N_10507,N_10405);
xor U11228 (N_11228,N_10501,N_10778);
xnor U11229 (N_11229,N_10477,N_10340);
xnor U11230 (N_11230,N_10605,N_10552);
or U11231 (N_11231,N_10604,N_10776);
nand U11232 (N_11232,N_10308,N_10616);
nor U11233 (N_11233,N_10627,N_10407);
or U11234 (N_11234,N_10536,N_10242);
xor U11235 (N_11235,N_10314,N_10380);
and U11236 (N_11236,N_10674,N_10394);
nor U11237 (N_11237,N_10279,N_10707);
nor U11238 (N_11238,N_10362,N_10219);
xnor U11239 (N_11239,N_10689,N_10652);
and U11240 (N_11240,N_10619,N_10688);
nor U11241 (N_11241,N_10334,N_10634);
or U11242 (N_11242,N_10654,N_10379);
and U11243 (N_11243,N_10471,N_10251);
and U11244 (N_11244,N_10782,N_10384);
or U11245 (N_11245,N_10427,N_10624);
nand U11246 (N_11246,N_10243,N_10573);
xor U11247 (N_11247,N_10231,N_10212);
or U11248 (N_11248,N_10583,N_10471);
xnor U11249 (N_11249,N_10622,N_10296);
and U11250 (N_11250,N_10477,N_10403);
xnor U11251 (N_11251,N_10265,N_10264);
nor U11252 (N_11252,N_10332,N_10227);
xor U11253 (N_11253,N_10485,N_10555);
xor U11254 (N_11254,N_10711,N_10748);
and U11255 (N_11255,N_10683,N_10390);
nor U11256 (N_11256,N_10499,N_10562);
nand U11257 (N_11257,N_10400,N_10306);
xor U11258 (N_11258,N_10261,N_10422);
nand U11259 (N_11259,N_10677,N_10637);
or U11260 (N_11260,N_10717,N_10757);
xor U11261 (N_11261,N_10691,N_10348);
nand U11262 (N_11262,N_10619,N_10715);
or U11263 (N_11263,N_10506,N_10463);
nor U11264 (N_11264,N_10315,N_10328);
or U11265 (N_11265,N_10219,N_10529);
xor U11266 (N_11266,N_10697,N_10319);
nand U11267 (N_11267,N_10332,N_10646);
and U11268 (N_11268,N_10521,N_10346);
and U11269 (N_11269,N_10416,N_10284);
or U11270 (N_11270,N_10536,N_10402);
nor U11271 (N_11271,N_10502,N_10461);
nand U11272 (N_11272,N_10206,N_10276);
or U11273 (N_11273,N_10471,N_10656);
or U11274 (N_11274,N_10343,N_10700);
nand U11275 (N_11275,N_10486,N_10624);
xnor U11276 (N_11276,N_10370,N_10617);
or U11277 (N_11277,N_10349,N_10221);
or U11278 (N_11278,N_10321,N_10272);
or U11279 (N_11279,N_10629,N_10304);
and U11280 (N_11280,N_10293,N_10665);
nand U11281 (N_11281,N_10511,N_10313);
nor U11282 (N_11282,N_10300,N_10713);
nor U11283 (N_11283,N_10325,N_10457);
or U11284 (N_11284,N_10488,N_10307);
nand U11285 (N_11285,N_10630,N_10363);
or U11286 (N_11286,N_10603,N_10766);
and U11287 (N_11287,N_10454,N_10324);
and U11288 (N_11288,N_10740,N_10508);
and U11289 (N_11289,N_10627,N_10540);
or U11290 (N_11290,N_10328,N_10630);
nand U11291 (N_11291,N_10656,N_10230);
xor U11292 (N_11292,N_10280,N_10357);
xnor U11293 (N_11293,N_10715,N_10460);
nor U11294 (N_11294,N_10226,N_10433);
nor U11295 (N_11295,N_10640,N_10238);
nand U11296 (N_11296,N_10200,N_10304);
and U11297 (N_11297,N_10233,N_10314);
xor U11298 (N_11298,N_10272,N_10735);
or U11299 (N_11299,N_10755,N_10693);
nand U11300 (N_11300,N_10209,N_10333);
xor U11301 (N_11301,N_10371,N_10511);
nand U11302 (N_11302,N_10469,N_10577);
and U11303 (N_11303,N_10353,N_10449);
nor U11304 (N_11304,N_10712,N_10409);
or U11305 (N_11305,N_10439,N_10719);
and U11306 (N_11306,N_10551,N_10328);
and U11307 (N_11307,N_10287,N_10481);
nor U11308 (N_11308,N_10267,N_10508);
nand U11309 (N_11309,N_10378,N_10345);
or U11310 (N_11310,N_10254,N_10415);
nor U11311 (N_11311,N_10773,N_10799);
or U11312 (N_11312,N_10386,N_10365);
or U11313 (N_11313,N_10267,N_10252);
nor U11314 (N_11314,N_10784,N_10601);
nor U11315 (N_11315,N_10431,N_10374);
xnor U11316 (N_11316,N_10744,N_10670);
and U11317 (N_11317,N_10461,N_10449);
xnor U11318 (N_11318,N_10756,N_10294);
xnor U11319 (N_11319,N_10745,N_10249);
and U11320 (N_11320,N_10234,N_10794);
or U11321 (N_11321,N_10423,N_10472);
or U11322 (N_11322,N_10216,N_10786);
or U11323 (N_11323,N_10784,N_10254);
nor U11324 (N_11324,N_10759,N_10417);
nand U11325 (N_11325,N_10389,N_10570);
nand U11326 (N_11326,N_10209,N_10757);
nand U11327 (N_11327,N_10652,N_10749);
and U11328 (N_11328,N_10783,N_10662);
xnor U11329 (N_11329,N_10766,N_10325);
nor U11330 (N_11330,N_10414,N_10591);
nand U11331 (N_11331,N_10492,N_10712);
nor U11332 (N_11332,N_10315,N_10531);
xnor U11333 (N_11333,N_10205,N_10390);
xor U11334 (N_11334,N_10262,N_10645);
or U11335 (N_11335,N_10304,N_10320);
nor U11336 (N_11336,N_10494,N_10320);
xnor U11337 (N_11337,N_10552,N_10227);
or U11338 (N_11338,N_10376,N_10477);
nand U11339 (N_11339,N_10668,N_10435);
or U11340 (N_11340,N_10602,N_10291);
or U11341 (N_11341,N_10657,N_10360);
and U11342 (N_11342,N_10442,N_10477);
nand U11343 (N_11343,N_10279,N_10590);
nor U11344 (N_11344,N_10226,N_10390);
nor U11345 (N_11345,N_10518,N_10416);
xor U11346 (N_11346,N_10727,N_10492);
and U11347 (N_11347,N_10609,N_10411);
nor U11348 (N_11348,N_10461,N_10318);
or U11349 (N_11349,N_10576,N_10436);
nor U11350 (N_11350,N_10741,N_10379);
or U11351 (N_11351,N_10519,N_10538);
and U11352 (N_11352,N_10214,N_10653);
xnor U11353 (N_11353,N_10795,N_10345);
and U11354 (N_11354,N_10657,N_10521);
or U11355 (N_11355,N_10476,N_10258);
xor U11356 (N_11356,N_10678,N_10539);
and U11357 (N_11357,N_10759,N_10657);
or U11358 (N_11358,N_10553,N_10656);
or U11359 (N_11359,N_10539,N_10215);
nor U11360 (N_11360,N_10411,N_10558);
or U11361 (N_11361,N_10372,N_10697);
or U11362 (N_11362,N_10530,N_10674);
and U11363 (N_11363,N_10295,N_10428);
nand U11364 (N_11364,N_10414,N_10745);
nor U11365 (N_11365,N_10502,N_10795);
nand U11366 (N_11366,N_10250,N_10451);
and U11367 (N_11367,N_10736,N_10672);
nand U11368 (N_11368,N_10539,N_10419);
and U11369 (N_11369,N_10659,N_10795);
nor U11370 (N_11370,N_10453,N_10505);
and U11371 (N_11371,N_10496,N_10799);
nor U11372 (N_11372,N_10287,N_10201);
and U11373 (N_11373,N_10374,N_10583);
nor U11374 (N_11374,N_10626,N_10649);
nand U11375 (N_11375,N_10237,N_10392);
and U11376 (N_11376,N_10711,N_10693);
nor U11377 (N_11377,N_10690,N_10612);
nand U11378 (N_11378,N_10548,N_10325);
and U11379 (N_11379,N_10499,N_10775);
or U11380 (N_11380,N_10226,N_10533);
and U11381 (N_11381,N_10725,N_10338);
nand U11382 (N_11382,N_10727,N_10220);
or U11383 (N_11383,N_10706,N_10261);
nand U11384 (N_11384,N_10747,N_10643);
nor U11385 (N_11385,N_10511,N_10523);
and U11386 (N_11386,N_10521,N_10419);
and U11387 (N_11387,N_10636,N_10311);
xnor U11388 (N_11388,N_10676,N_10377);
nand U11389 (N_11389,N_10757,N_10247);
and U11390 (N_11390,N_10236,N_10619);
nor U11391 (N_11391,N_10798,N_10598);
and U11392 (N_11392,N_10355,N_10679);
xnor U11393 (N_11393,N_10471,N_10794);
nor U11394 (N_11394,N_10785,N_10397);
nand U11395 (N_11395,N_10649,N_10606);
nor U11396 (N_11396,N_10465,N_10672);
xnor U11397 (N_11397,N_10660,N_10215);
xor U11398 (N_11398,N_10361,N_10496);
nor U11399 (N_11399,N_10759,N_10293);
nand U11400 (N_11400,N_10854,N_11274);
nor U11401 (N_11401,N_10844,N_11023);
nand U11402 (N_11402,N_10903,N_11368);
and U11403 (N_11403,N_11364,N_11084);
nand U11404 (N_11404,N_11395,N_11133);
nor U11405 (N_11405,N_11048,N_10954);
and U11406 (N_11406,N_10908,N_10824);
or U11407 (N_11407,N_11359,N_10809);
nand U11408 (N_11408,N_11076,N_10963);
nand U11409 (N_11409,N_11032,N_11194);
nor U11410 (N_11410,N_10898,N_10803);
or U11411 (N_11411,N_11270,N_10975);
or U11412 (N_11412,N_11268,N_11132);
nor U11413 (N_11413,N_11309,N_11393);
nand U11414 (N_11414,N_11341,N_11147);
nand U11415 (N_11415,N_11233,N_11107);
nor U11416 (N_11416,N_11079,N_11123);
and U11417 (N_11417,N_10909,N_11092);
xnor U11418 (N_11418,N_11174,N_11288);
xor U11419 (N_11419,N_11322,N_10902);
xnor U11420 (N_11420,N_11355,N_10845);
or U11421 (N_11421,N_10862,N_11386);
nand U11422 (N_11422,N_11223,N_10956);
xnor U11423 (N_11423,N_11303,N_11319);
xor U11424 (N_11424,N_11176,N_10828);
nand U11425 (N_11425,N_10891,N_11028);
or U11426 (N_11426,N_11086,N_11228);
nor U11427 (N_11427,N_11334,N_11247);
and U11428 (N_11428,N_11162,N_11356);
or U11429 (N_11429,N_11090,N_10804);
xnor U11430 (N_11430,N_11367,N_11034);
nand U11431 (N_11431,N_11281,N_11026);
nor U11432 (N_11432,N_11054,N_11128);
and U11433 (N_11433,N_11057,N_10887);
and U11434 (N_11434,N_11178,N_10806);
and U11435 (N_11435,N_10964,N_10812);
nor U11436 (N_11436,N_10955,N_10833);
nor U11437 (N_11437,N_11089,N_11015);
nor U11438 (N_11438,N_10872,N_11203);
xor U11439 (N_11439,N_11343,N_10999);
nor U11440 (N_11440,N_11141,N_10938);
and U11441 (N_11441,N_11192,N_11312);
or U11442 (N_11442,N_11031,N_11308);
nor U11443 (N_11443,N_11397,N_10935);
or U11444 (N_11444,N_11295,N_11314);
xor U11445 (N_11445,N_11232,N_10949);
nor U11446 (N_11446,N_10888,N_10879);
or U11447 (N_11447,N_10811,N_10852);
and U11448 (N_11448,N_11020,N_10974);
nor U11449 (N_11449,N_11243,N_11213);
xor U11450 (N_11450,N_11014,N_11065);
and U11451 (N_11451,N_11017,N_11399);
or U11452 (N_11452,N_11333,N_11197);
nor U11453 (N_11453,N_10966,N_11159);
xor U11454 (N_11454,N_11067,N_11053);
nor U11455 (N_11455,N_11383,N_10830);
nor U11456 (N_11456,N_11069,N_10931);
xor U11457 (N_11457,N_11236,N_11221);
xnor U11458 (N_11458,N_11182,N_11164);
and U11459 (N_11459,N_11366,N_11245);
or U11460 (N_11460,N_11006,N_11184);
or U11461 (N_11461,N_11160,N_11198);
and U11462 (N_11462,N_11169,N_10855);
and U11463 (N_11463,N_10962,N_10926);
or U11464 (N_11464,N_11384,N_11305);
and U11465 (N_11465,N_11254,N_10875);
nand U11466 (N_11466,N_10947,N_11306);
xnor U11467 (N_11467,N_11394,N_10894);
or U11468 (N_11468,N_11344,N_10937);
xnor U11469 (N_11469,N_11296,N_10985);
or U11470 (N_11470,N_11099,N_11326);
and U11471 (N_11471,N_11029,N_11064);
and U11472 (N_11472,N_11142,N_11177);
or U11473 (N_11473,N_11327,N_11339);
and U11474 (N_11474,N_11199,N_10936);
xnor U11475 (N_11475,N_11137,N_11004);
nand U11476 (N_11476,N_11003,N_11350);
xnor U11477 (N_11477,N_10823,N_10896);
nand U11478 (N_11478,N_10969,N_11362);
nor U11479 (N_11479,N_10991,N_10876);
xnor U11480 (N_11480,N_11082,N_10993);
xor U11481 (N_11481,N_11220,N_11127);
nor U11482 (N_11482,N_11136,N_10960);
or U11483 (N_11483,N_11300,N_10929);
nand U11484 (N_11484,N_10822,N_11181);
xnor U11485 (N_11485,N_11385,N_10987);
and U11486 (N_11486,N_11098,N_11338);
nand U11487 (N_11487,N_10815,N_10881);
nand U11488 (N_11488,N_11321,N_10972);
and U11489 (N_11489,N_11250,N_11037);
or U11490 (N_11490,N_11377,N_11258);
xor U11491 (N_11491,N_10976,N_11150);
xnor U11492 (N_11492,N_11371,N_10910);
xnor U11493 (N_11493,N_11242,N_11323);
and U11494 (N_11494,N_11106,N_11072);
nand U11495 (N_11495,N_11271,N_11167);
xnor U11496 (N_11496,N_11075,N_11055);
xnor U11497 (N_11497,N_10818,N_11110);
nand U11498 (N_11498,N_10856,N_11349);
nor U11499 (N_11499,N_11033,N_10873);
nor U11500 (N_11500,N_11298,N_10846);
nor U11501 (N_11501,N_10980,N_11313);
or U11502 (N_11502,N_11325,N_11279);
and U11503 (N_11503,N_11390,N_11013);
and U11504 (N_11504,N_11264,N_11130);
nor U11505 (N_11505,N_11149,N_11116);
xnor U11506 (N_11506,N_11140,N_11117);
and U11507 (N_11507,N_11345,N_11216);
or U11508 (N_11508,N_10821,N_10890);
and U11509 (N_11509,N_10829,N_10988);
nor U11510 (N_11510,N_10904,N_10843);
or U11511 (N_11511,N_11027,N_11318);
nor U11512 (N_11512,N_11387,N_10942);
nor U11513 (N_11513,N_10978,N_11108);
xnor U11514 (N_11514,N_10912,N_11139);
or U11515 (N_11515,N_10866,N_10897);
xor U11516 (N_11516,N_10899,N_11148);
and U11517 (N_11517,N_11294,N_11052);
nand U11518 (N_11518,N_10944,N_10906);
nand U11519 (N_11519,N_11277,N_11261);
and U11520 (N_11520,N_11155,N_11074);
nor U11521 (N_11521,N_11389,N_11269);
or U11522 (N_11522,N_11043,N_11201);
or U11523 (N_11523,N_10895,N_11248);
nor U11524 (N_11524,N_11091,N_11179);
and U11525 (N_11525,N_11024,N_11267);
nor U11526 (N_11526,N_11287,N_10940);
or U11527 (N_11527,N_11154,N_10917);
nand U11528 (N_11528,N_11129,N_11146);
nor U11529 (N_11529,N_10847,N_11195);
xor U11530 (N_11530,N_11378,N_11022);
and U11531 (N_11531,N_10934,N_10877);
or U11532 (N_11532,N_11114,N_10826);
xnor U11533 (N_11533,N_11101,N_11212);
nor U11534 (N_11534,N_11060,N_11219);
nand U11535 (N_11535,N_10870,N_11105);
nand U11536 (N_11536,N_11125,N_11068);
xnor U11537 (N_11537,N_11234,N_11392);
xor U11538 (N_11538,N_11097,N_11342);
and U11539 (N_11539,N_10907,N_11376);
nor U11540 (N_11540,N_10957,N_10827);
or U11541 (N_11541,N_11070,N_10983);
xor U11542 (N_11542,N_10863,N_11189);
xnor U11543 (N_11543,N_10914,N_11008);
nand U11544 (N_11544,N_11200,N_11347);
xor U11545 (N_11545,N_11044,N_10807);
nand U11546 (N_11546,N_11235,N_11265);
or U11547 (N_11547,N_11340,N_11175);
or U11548 (N_11548,N_11187,N_11357);
nand U11549 (N_11549,N_10842,N_11291);
nor U11550 (N_11550,N_11163,N_11286);
nor U11551 (N_11551,N_11227,N_10998);
nor U11552 (N_11552,N_11172,N_11225);
or U11553 (N_11553,N_10885,N_11310);
or U11554 (N_11554,N_10820,N_11276);
xnor U11555 (N_11555,N_10990,N_11257);
and U11556 (N_11556,N_10973,N_10825);
nor U11557 (N_11557,N_11215,N_11019);
nand U11558 (N_11558,N_10950,N_11369);
and U11559 (N_11559,N_11186,N_10816);
nand U11560 (N_11560,N_11238,N_11188);
xnor U11561 (N_11561,N_11217,N_11002);
nand U11562 (N_11562,N_11165,N_11100);
nor U11563 (N_11563,N_11205,N_11185);
nor U11564 (N_11564,N_11051,N_10831);
xor U11565 (N_11565,N_10933,N_11204);
or U11566 (N_11566,N_11373,N_10860);
and U11567 (N_11567,N_11280,N_11348);
nor U11568 (N_11568,N_10921,N_11253);
and U11569 (N_11569,N_11284,N_11104);
nor U11570 (N_11570,N_11226,N_11039);
xnor U11571 (N_11571,N_10892,N_11040);
nand U11572 (N_11572,N_11030,N_10851);
xnor U11573 (N_11573,N_10995,N_11272);
nand U11574 (N_11574,N_11061,N_11007);
nor U11575 (N_11575,N_11011,N_11244);
or U11576 (N_11576,N_11056,N_11191);
nor U11577 (N_11577,N_10883,N_10943);
and U11578 (N_11578,N_11012,N_11038);
nor U11579 (N_11579,N_11046,N_11208);
nand U11580 (N_11580,N_10819,N_10836);
and U11581 (N_11581,N_10874,N_11211);
nor U11582 (N_11582,N_11374,N_11352);
nor U11583 (N_11583,N_10832,N_11047);
nor U11584 (N_11584,N_11207,N_11237);
and U11585 (N_11585,N_11094,N_10878);
xnor U11586 (N_11586,N_10981,N_10850);
xnor U11587 (N_11587,N_10901,N_11266);
xor U11588 (N_11588,N_10932,N_10853);
nor U11589 (N_11589,N_11260,N_10849);
or U11590 (N_11590,N_11001,N_11126);
nor U11591 (N_11591,N_11025,N_11379);
or U11592 (N_11592,N_11124,N_11157);
xnor U11593 (N_11593,N_11170,N_10841);
xnor U11594 (N_11594,N_11190,N_11088);
and U11595 (N_11595,N_11336,N_11398);
and U11596 (N_11596,N_11131,N_11346);
nor U11597 (N_11597,N_11171,N_11290);
nand U11598 (N_11598,N_10808,N_11121);
nor U11599 (N_11599,N_10967,N_11381);
and U11600 (N_11600,N_11222,N_11256);
and U11601 (N_11601,N_11283,N_10979);
nand U11602 (N_11602,N_10858,N_10882);
or U11603 (N_11603,N_11358,N_11144);
and U11604 (N_11604,N_11380,N_11016);
or U11605 (N_11605,N_10864,N_11302);
nand U11606 (N_11606,N_10994,N_10986);
nand U11607 (N_11607,N_11293,N_11331);
nand U11608 (N_11608,N_11118,N_11173);
and U11609 (N_11609,N_11263,N_11289);
or U11610 (N_11610,N_10837,N_10840);
nor U11611 (N_11611,N_10884,N_11050);
xor U11612 (N_11612,N_11009,N_11388);
nand U11613 (N_11613,N_11229,N_11005);
and U11614 (N_11614,N_11071,N_11351);
nor U11615 (N_11615,N_10839,N_11360);
nand U11616 (N_11616,N_11196,N_11093);
or U11617 (N_11617,N_10930,N_10923);
or U11618 (N_11618,N_11145,N_10977);
nand U11619 (N_11619,N_10971,N_10848);
or U11620 (N_11620,N_11249,N_11241);
nor U11621 (N_11621,N_10997,N_11275);
nand U11622 (N_11622,N_11143,N_11297);
nand U11623 (N_11623,N_11063,N_11224);
xnor U11624 (N_11624,N_11375,N_11119);
or U11625 (N_11625,N_11328,N_10900);
nand U11626 (N_11626,N_11396,N_10817);
xor U11627 (N_11627,N_10889,N_11354);
and U11628 (N_11628,N_11335,N_11151);
nor U11629 (N_11629,N_10810,N_10838);
or U11630 (N_11630,N_10922,N_10968);
nor U11631 (N_11631,N_11301,N_11320);
nand U11632 (N_11632,N_11304,N_10868);
and U11633 (N_11633,N_10802,N_11035);
nand U11634 (N_11634,N_11218,N_10859);
and U11635 (N_11635,N_10919,N_11231);
nor U11636 (N_11636,N_11083,N_11214);
or U11637 (N_11637,N_11021,N_11087);
nand U11638 (N_11638,N_11096,N_10913);
nor U11639 (N_11639,N_11282,N_11042);
or U11640 (N_11640,N_11041,N_11202);
and U11641 (N_11641,N_11183,N_11246);
or U11642 (N_11642,N_10805,N_10813);
nor U11643 (N_11643,N_11134,N_10893);
and U11644 (N_11644,N_10982,N_11018);
or U11645 (N_11645,N_11077,N_11209);
nand U11646 (N_11646,N_11112,N_10918);
nor U11647 (N_11647,N_11259,N_11109);
or U11648 (N_11648,N_11315,N_10916);
xor U11649 (N_11649,N_11156,N_11206);
nor U11650 (N_11650,N_11252,N_11158);
and U11651 (N_11651,N_10992,N_10801);
and U11652 (N_11652,N_10965,N_11103);
xor U11653 (N_11653,N_11251,N_10880);
nand U11654 (N_11654,N_11166,N_11311);
or U11655 (N_11655,N_11080,N_11078);
or U11656 (N_11656,N_10945,N_10996);
and U11657 (N_11657,N_11193,N_10952);
or U11658 (N_11658,N_10915,N_10911);
and U11659 (N_11659,N_10920,N_11330);
xnor U11660 (N_11660,N_11210,N_10905);
xor U11661 (N_11661,N_11168,N_10946);
nor U11662 (N_11662,N_11081,N_11161);
nand U11663 (N_11663,N_11135,N_11239);
nor U11664 (N_11664,N_11332,N_10800);
xor U11665 (N_11665,N_10886,N_11307);
xor U11666 (N_11666,N_11122,N_11152);
nor U11667 (N_11667,N_11316,N_11058);
nor U11668 (N_11668,N_10959,N_11230);
nor U11669 (N_11669,N_11353,N_10924);
or U11670 (N_11670,N_11066,N_10867);
or U11671 (N_11671,N_11382,N_11045);
and U11672 (N_11672,N_11317,N_10925);
or U11673 (N_11673,N_11391,N_11062);
nor U11674 (N_11674,N_10857,N_11180);
nand U11675 (N_11675,N_11278,N_11273);
nor U11676 (N_11676,N_11115,N_10989);
nand U11677 (N_11677,N_11153,N_11095);
and U11678 (N_11678,N_11085,N_11111);
nor U11679 (N_11679,N_10869,N_10865);
and U11680 (N_11680,N_10927,N_10984);
xnor U11681 (N_11681,N_10939,N_10970);
xor U11682 (N_11682,N_11329,N_11000);
and U11683 (N_11683,N_10941,N_11120);
and U11684 (N_11684,N_11262,N_11113);
xnor U11685 (N_11685,N_10928,N_11292);
xor U11686 (N_11686,N_11036,N_10861);
nand U11687 (N_11687,N_11059,N_11102);
nand U11688 (N_11688,N_11010,N_11365);
xor U11689 (N_11689,N_11240,N_11138);
and U11690 (N_11690,N_10834,N_11049);
and U11691 (N_11691,N_10814,N_10835);
xor U11692 (N_11692,N_10958,N_11073);
or U11693 (N_11693,N_11372,N_11363);
nor U11694 (N_11694,N_11285,N_10871);
xnor U11695 (N_11695,N_11324,N_10953);
nor U11696 (N_11696,N_11361,N_11370);
and U11697 (N_11697,N_11337,N_10951);
and U11698 (N_11698,N_10961,N_11299);
xor U11699 (N_11699,N_11255,N_10948);
xnor U11700 (N_11700,N_11394,N_11098);
xnor U11701 (N_11701,N_10912,N_10879);
nand U11702 (N_11702,N_11367,N_11154);
xnor U11703 (N_11703,N_11024,N_11378);
and U11704 (N_11704,N_10864,N_10947);
or U11705 (N_11705,N_11281,N_11359);
and U11706 (N_11706,N_11347,N_11286);
xor U11707 (N_11707,N_11349,N_11219);
nand U11708 (N_11708,N_10987,N_11014);
nor U11709 (N_11709,N_11114,N_11040);
nand U11710 (N_11710,N_11029,N_10970);
nand U11711 (N_11711,N_10820,N_10891);
or U11712 (N_11712,N_11152,N_10815);
xor U11713 (N_11713,N_11113,N_11172);
xnor U11714 (N_11714,N_11355,N_11258);
nor U11715 (N_11715,N_11365,N_11132);
nor U11716 (N_11716,N_11144,N_11029);
nor U11717 (N_11717,N_11057,N_10903);
or U11718 (N_11718,N_11294,N_10968);
nand U11719 (N_11719,N_10875,N_11252);
xor U11720 (N_11720,N_10966,N_10821);
nor U11721 (N_11721,N_10921,N_10805);
nor U11722 (N_11722,N_11210,N_11286);
nor U11723 (N_11723,N_11188,N_11113);
nor U11724 (N_11724,N_11074,N_11371);
or U11725 (N_11725,N_10806,N_11085);
nand U11726 (N_11726,N_11016,N_11292);
nand U11727 (N_11727,N_10994,N_10846);
or U11728 (N_11728,N_11295,N_11115);
or U11729 (N_11729,N_11393,N_11347);
and U11730 (N_11730,N_10869,N_10913);
xnor U11731 (N_11731,N_10828,N_11121);
and U11732 (N_11732,N_10939,N_11050);
and U11733 (N_11733,N_10832,N_10816);
nand U11734 (N_11734,N_11358,N_10855);
and U11735 (N_11735,N_11049,N_10977);
nor U11736 (N_11736,N_11114,N_11265);
nor U11737 (N_11737,N_11080,N_11291);
or U11738 (N_11738,N_11242,N_11184);
nor U11739 (N_11739,N_11259,N_11110);
nor U11740 (N_11740,N_11152,N_11232);
xnor U11741 (N_11741,N_10813,N_11309);
and U11742 (N_11742,N_11363,N_11008);
xor U11743 (N_11743,N_11338,N_11208);
nand U11744 (N_11744,N_10812,N_11108);
or U11745 (N_11745,N_11065,N_11015);
and U11746 (N_11746,N_11220,N_11225);
and U11747 (N_11747,N_11373,N_11126);
or U11748 (N_11748,N_11266,N_11052);
and U11749 (N_11749,N_10927,N_10994);
xnor U11750 (N_11750,N_10832,N_10841);
and U11751 (N_11751,N_10922,N_11215);
and U11752 (N_11752,N_11284,N_11142);
nor U11753 (N_11753,N_11012,N_10962);
nor U11754 (N_11754,N_10942,N_11333);
xor U11755 (N_11755,N_10832,N_11099);
xor U11756 (N_11756,N_11373,N_10951);
xnor U11757 (N_11757,N_10933,N_11314);
or U11758 (N_11758,N_11386,N_10881);
or U11759 (N_11759,N_11254,N_11350);
and U11760 (N_11760,N_11285,N_10802);
and U11761 (N_11761,N_11319,N_11210);
nand U11762 (N_11762,N_10862,N_11144);
nor U11763 (N_11763,N_11138,N_11062);
and U11764 (N_11764,N_11290,N_11080);
and U11765 (N_11765,N_11062,N_10842);
nand U11766 (N_11766,N_11338,N_11234);
or U11767 (N_11767,N_11169,N_11213);
and U11768 (N_11768,N_11227,N_10825);
nand U11769 (N_11769,N_11371,N_11152);
or U11770 (N_11770,N_10985,N_10999);
nand U11771 (N_11771,N_11099,N_10806);
and U11772 (N_11772,N_11194,N_10968);
or U11773 (N_11773,N_10802,N_10981);
xnor U11774 (N_11774,N_11121,N_11175);
nor U11775 (N_11775,N_10934,N_11058);
or U11776 (N_11776,N_11113,N_11120);
nor U11777 (N_11777,N_11013,N_11384);
nand U11778 (N_11778,N_10847,N_11332);
xnor U11779 (N_11779,N_11306,N_11026);
nor U11780 (N_11780,N_11252,N_11082);
nor U11781 (N_11781,N_11198,N_11190);
xor U11782 (N_11782,N_10823,N_11154);
and U11783 (N_11783,N_11205,N_10910);
xor U11784 (N_11784,N_10816,N_11211);
nor U11785 (N_11785,N_11331,N_10807);
nor U11786 (N_11786,N_10836,N_10886);
nand U11787 (N_11787,N_11216,N_10900);
and U11788 (N_11788,N_11366,N_11205);
xor U11789 (N_11789,N_11376,N_11256);
or U11790 (N_11790,N_11058,N_11348);
and U11791 (N_11791,N_10901,N_11176);
and U11792 (N_11792,N_11268,N_11237);
or U11793 (N_11793,N_11242,N_11337);
and U11794 (N_11794,N_11131,N_11069);
or U11795 (N_11795,N_11137,N_11254);
nor U11796 (N_11796,N_10817,N_11018);
nor U11797 (N_11797,N_11257,N_10989);
or U11798 (N_11798,N_10892,N_11301);
nor U11799 (N_11799,N_10954,N_10863);
xnor U11800 (N_11800,N_11228,N_11014);
nand U11801 (N_11801,N_11103,N_10832);
or U11802 (N_11802,N_10892,N_11111);
and U11803 (N_11803,N_11089,N_11389);
xnor U11804 (N_11804,N_11370,N_10987);
and U11805 (N_11805,N_11265,N_10844);
xnor U11806 (N_11806,N_11309,N_10900);
or U11807 (N_11807,N_11240,N_11104);
nand U11808 (N_11808,N_11333,N_11292);
nor U11809 (N_11809,N_11266,N_11248);
or U11810 (N_11810,N_10914,N_11177);
xnor U11811 (N_11811,N_11306,N_11285);
xnor U11812 (N_11812,N_11369,N_11250);
nor U11813 (N_11813,N_11234,N_11197);
nand U11814 (N_11814,N_11042,N_11378);
and U11815 (N_11815,N_11323,N_11142);
and U11816 (N_11816,N_10972,N_11056);
or U11817 (N_11817,N_10855,N_10912);
xnor U11818 (N_11818,N_11343,N_11338);
xor U11819 (N_11819,N_10807,N_10815);
nor U11820 (N_11820,N_11270,N_10881);
or U11821 (N_11821,N_10913,N_10886);
or U11822 (N_11822,N_11334,N_11085);
nand U11823 (N_11823,N_11067,N_10924);
xnor U11824 (N_11824,N_11235,N_11081);
nand U11825 (N_11825,N_10985,N_10974);
and U11826 (N_11826,N_10902,N_11264);
and U11827 (N_11827,N_11367,N_10822);
nand U11828 (N_11828,N_11214,N_11280);
xor U11829 (N_11829,N_10870,N_11148);
and U11830 (N_11830,N_11098,N_11392);
and U11831 (N_11831,N_11322,N_10861);
xnor U11832 (N_11832,N_11082,N_10981);
xnor U11833 (N_11833,N_11114,N_11250);
nand U11834 (N_11834,N_11259,N_11389);
nor U11835 (N_11835,N_11366,N_11253);
xnor U11836 (N_11836,N_10936,N_11267);
nand U11837 (N_11837,N_11168,N_10830);
xor U11838 (N_11838,N_11202,N_11214);
or U11839 (N_11839,N_11274,N_11085);
nor U11840 (N_11840,N_10802,N_10872);
and U11841 (N_11841,N_11374,N_10823);
xor U11842 (N_11842,N_10871,N_11050);
or U11843 (N_11843,N_10877,N_11328);
and U11844 (N_11844,N_11165,N_10832);
or U11845 (N_11845,N_10928,N_11028);
nand U11846 (N_11846,N_11258,N_11097);
or U11847 (N_11847,N_11237,N_11296);
nor U11848 (N_11848,N_11309,N_11031);
nor U11849 (N_11849,N_11169,N_11296);
xor U11850 (N_11850,N_11308,N_10858);
nand U11851 (N_11851,N_10840,N_10959);
or U11852 (N_11852,N_11033,N_11303);
xor U11853 (N_11853,N_11094,N_10997);
xor U11854 (N_11854,N_10958,N_11106);
xnor U11855 (N_11855,N_10828,N_10947);
xnor U11856 (N_11856,N_11264,N_11298);
and U11857 (N_11857,N_11230,N_11284);
xnor U11858 (N_11858,N_11249,N_11321);
or U11859 (N_11859,N_10890,N_10854);
xnor U11860 (N_11860,N_11242,N_11133);
xnor U11861 (N_11861,N_11342,N_10994);
nor U11862 (N_11862,N_10826,N_11373);
or U11863 (N_11863,N_11199,N_10810);
nor U11864 (N_11864,N_11080,N_10943);
or U11865 (N_11865,N_11165,N_11323);
and U11866 (N_11866,N_11153,N_11044);
nor U11867 (N_11867,N_11001,N_11056);
nor U11868 (N_11868,N_11051,N_10889);
or U11869 (N_11869,N_10834,N_11180);
xor U11870 (N_11870,N_10849,N_10824);
nand U11871 (N_11871,N_11358,N_11212);
nor U11872 (N_11872,N_11384,N_11243);
nand U11873 (N_11873,N_10845,N_11153);
nor U11874 (N_11874,N_11236,N_11184);
nand U11875 (N_11875,N_10865,N_10864);
or U11876 (N_11876,N_11134,N_11326);
and U11877 (N_11877,N_11059,N_11113);
and U11878 (N_11878,N_10872,N_11231);
or U11879 (N_11879,N_11000,N_11237);
nand U11880 (N_11880,N_11000,N_11312);
nand U11881 (N_11881,N_10848,N_11233);
xnor U11882 (N_11882,N_11088,N_10852);
nand U11883 (N_11883,N_11161,N_10986);
and U11884 (N_11884,N_11349,N_11376);
and U11885 (N_11885,N_10858,N_11108);
nand U11886 (N_11886,N_11277,N_11057);
nor U11887 (N_11887,N_11096,N_11139);
nor U11888 (N_11888,N_10950,N_11081);
or U11889 (N_11889,N_10917,N_10866);
or U11890 (N_11890,N_11292,N_11300);
or U11891 (N_11891,N_11204,N_10845);
nor U11892 (N_11892,N_11198,N_10866);
xnor U11893 (N_11893,N_11308,N_10955);
nor U11894 (N_11894,N_11251,N_11358);
xnor U11895 (N_11895,N_10982,N_11129);
xnor U11896 (N_11896,N_11310,N_11287);
and U11897 (N_11897,N_11194,N_11051);
nor U11898 (N_11898,N_11221,N_11012);
and U11899 (N_11899,N_10818,N_10911);
and U11900 (N_11900,N_11007,N_11320);
xor U11901 (N_11901,N_11140,N_10890);
or U11902 (N_11902,N_10961,N_11390);
nand U11903 (N_11903,N_11007,N_11107);
nand U11904 (N_11904,N_11203,N_10906);
xor U11905 (N_11905,N_10946,N_11159);
nand U11906 (N_11906,N_11347,N_11333);
xnor U11907 (N_11907,N_11209,N_10884);
nor U11908 (N_11908,N_10954,N_11108);
nor U11909 (N_11909,N_10833,N_11392);
nor U11910 (N_11910,N_11236,N_11000);
or U11911 (N_11911,N_11374,N_10984);
and U11912 (N_11912,N_11078,N_11189);
nor U11913 (N_11913,N_11302,N_11097);
nand U11914 (N_11914,N_11092,N_10863);
and U11915 (N_11915,N_11185,N_10900);
and U11916 (N_11916,N_10851,N_11314);
nand U11917 (N_11917,N_11123,N_10899);
or U11918 (N_11918,N_11268,N_10839);
nor U11919 (N_11919,N_10973,N_10827);
nor U11920 (N_11920,N_10916,N_10810);
xnor U11921 (N_11921,N_11079,N_10818);
nor U11922 (N_11922,N_11301,N_11038);
and U11923 (N_11923,N_11094,N_11144);
and U11924 (N_11924,N_10953,N_11234);
nand U11925 (N_11925,N_10976,N_11182);
nand U11926 (N_11926,N_11290,N_10886);
xor U11927 (N_11927,N_10974,N_10905);
nor U11928 (N_11928,N_11066,N_10820);
or U11929 (N_11929,N_11053,N_11377);
and U11930 (N_11930,N_10995,N_11135);
and U11931 (N_11931,N_10890,N_11025);
or U11932 (N_11932,N_11016,N_11331);
nor U11933 (N_11933,N_11189,N_11274);
or U11934 (N_11934,N_11125,N_11161);
nor U11935 (N_11935,N_11353,N_10841);
or U11936 (N_11936,N_10885,N_11348);
or U11937 (N_11937,N_11269,N_11177);
nand U11938 (N_11938,N_11253,N_11177);
nor U11939 (N_11939,N_11062,N_11109);
xor U11940 (N_11940,N_11255,N_10935);
nand U11941 (N_11941,N_11303,N_11225);
and U11942 (N_11942,N_10816,N_11055);
xor U11943 (N_11943,N_11318,N_10991);
and U11944 (N_11944,N_11224,N_11118);
or U11945 (N_11945,N_10894,N_10994);
nor U11946 (N_11946,N_11307,N_11037);
nand U11947 (N_11947,N_11391,N_11000);
nand U11948 (N_11948,N_10827,N_11218);
or U11949 (N_11949,N_11230,N_10906);
nor U11950 (N_11950,N_11138,N_11398);
xnor U11951 (N_11951,N_11319,N_11391);
nand U11952 (N_11952,N_11184,N_11397);
nand U11953 (N_11953,N_11174,N_11125);
xor U11954 (N_11954,N_11316,N_11124);
or U11955 (N_11955,N_10968,N_10955);
nor U11956 (N_11956,N_10831,N_11359);
nand U11957 (N_11957,N_11114,N_10993);
or U11958 (N_11958,N_11207,N_11120);
xnor U11959 (N_11959,N_11066,N_11361);
or U11960 (N_11960,N_11219,N_10880);
or U11961 (N_11961,N_11047,N_11367);
and U11962 (N_11962,N_11172,N_11361);
xor U11963 (N_11963,N_10803,N_10875);
nand U11964 (N_11964,N_11067,N_10901);
nand U11965 (N_11965,N_10904,N_10920);
and U11966 (N_11966,N_10891,N_11140);
xnor U11967 (N_11967,N_11243,N_10848);
or U11968 (N_11968,N_11369,N_10976);
and U11969 (N_11969,N_11059,N_10980);
xor U11970 (N_11970,N_11359,N_11181);
or U11971 (N_11971,N_11037,N_11239);
or U11972 (N_11972,N_11132,N_11362);
xor U11973 (N_11973,N_11092,N_11240);
nor U11974 (N_11974,N_10994,N_10955);
nor U11975 (N_11975,N_11293,N_11385);
and U11976 (N_11976,N_10876,N_11375);
nor U11977 (N_11977,N_11380,N_10957);
nand U11978 (N_11978,N_10814,N_11005);
and U11979 (N_11979,N_11014,N_10894);
nand U11980 (N_11980,N_11378,N_11212);
or U11981 (N_11981,N_10982,N_11205);
or U11982 (N_11982,N_11292,N_10837);
or U11983 (N_11983,N_10968,N_10954);
and U11984 (N_11984,N_10909,N_11127);
nor U11985 (N_11985,N_11317,N_11181);
nor U11986 (N_11986,N_10897,N_11260);
nor U11987 (N_11987,N_10869,N_11347);
nand U11988 (N_11988,N_11028,N_11274);
nand U11989 (N_11989,N_10910,N_10883);
xnor U11990 (N_11990,N_10814,N_11139);
and U11991 (N_11991,N_10839,N_10999);
or U11992 (N_11992,N_11267,N_11153);
nand U11993 (N_11993,N_11042,N_10903);
nand U11994 (N_11994,N_11075,N_10875);
nand U11995 (N_11995,N_10963,N_11174);
nand U11996 (N_11996,N_10812,N_10925);
nand U11997 (N_11997,N_11239,N_11301);
nor U11998 (N_11998,N_10986,N_11399);
and U11999 (N_11999,N_11079,N_10899);
xor U12000 (N_12000,N_11575,N_11946);
or U12001 (N_12001,N_11495,N_11621);
and U12002 (N_12002,N_11602,N_11985);
and U12003 (N_12003,N_11958,N_11537);
nor U12004 (N_12004,N_11791,N_11923);
or U12005 (N_12005,N_11699,N_11926);
nor U12006 (N_12006,N_11645,N_11956);
nand U12007 (N_12007,N_11641,N_11427);
and U12008 (N_12008,N_11994,N_11919);
or U12009 (N_12009,N_11802,N_11516);
nor U12010 (N_12010,N_11662,N_11734);
and U12011 (N_12011,N_11903,N_11932);
nor U12012 (N_12012,N_11543,N_11770);
nor U12013 (N_12013,N_11873,N_11678);
or U12014 (N_12014,N_11927,N_11717);
nor U12015 (N_12015,N_11786,N_11401);
or U12016 (N_12016,N_11476,N_11400);
xor U12017 (N_12017,N_11521,N_11478);
xnor U12018 (N_12018,N_11584,N_11744);
and U12019 (N_12019,N_11862,N_11914);
xnor U12020 (N_12020,N_11829,N_11644);
nor U12021 (N_12021,N_11954,N_11413);
or U12022 (N_12022,N_11680,N_11733);
or U12023 (N_12023,N_11855,N_11485);
and U12024 (N_12024,N_11850,N_11664);
or U12025 (N_12025,N_11816,N_11824);
and U12026 (N_12026,N_11606,N_11812);
xor U12027 (N_12027,N_11568,N_11623);
nand U12028 (N_12028,N_11686,N_11777);
or U12029 (N_12029,N_11940,N_11555);
xnor U12030 (N_12030,N_11915,N_11975);
nand U12031 (N_12031,N_11481,N_11809);
and U12032 (N_12032,N_11587,N_11776);
nand U12033 (N_12033,N_11920,N_11806);
nor U12034 (N_12034,N_11719,N_11986);
nor U12035 (N_12035,N_11789,N_11752);
or U12036 (N_12036,N_11827,N_11962);
and U12037 (N_12037,N_11529,N_11968);
and U12038 (N_12038,N_11679,N_11412);
nand U12039 (N_12039,N_11609,N_11909);
nor U12040 (N_12040,N_11727,N_11911);
nand U12041 (N_12041,N_11947,N_11710);
nor U12042 (N_12042,N_11561,N_11805);
nor U12043 (N_12043,N_11819,N_11488);
nand U12044 (N_12044,N_11432,N_11665);
xor U12045 (N_12045,N_11430,N_11886);
or U12046 (N_12046,N_11825,N_11702);
xor U12047 (N_12047,N_11512,N_11657);
nand U12048 (N_12048,N_11963,N_11953);
nand U12049 (N_12049,N_11640,N_11965);
or U12050 (N_12050,N_11961,N_11999);
nand U12051 (N_12051,N_11670,N_11697);
xnor U12052 (N_12052,N_11878,N_11472);
nor U12053 (N_12053,N_11658,N_11605);
nor U12054 (N_12054,N_11450,N_11864);
xnor U12055 (N_12055,N_11499,N_11936);
nor U12056 (N_12056,N_11627,N_11434);
and U12057 (N_12057,N_11804,N_11790);
and U12058 (N_12058,N_11580,N_11964);
xor U12059 (N_12059,N_11728,N_11939);
xnor U12060 (N_12060,N_11960,N_11766);
nand U12061 (N_12061,N_11690,N_11726);
nor U12062 (N_12062,N_11851,N_11970);
nor U12063 (N_12063,N_11496,N_11706);
nor U12064 (N_12064,N_11466,N_11979);
nor U12065 (N_12065,N_11801,N_11889);
nand U12066 (N_12066,N_11813,N_11504);
nor U12067 (N_12067,N_11431,N_11693);
or U12068 (N_12068,N_11474,N_11541);
nand U12069 (N_12069,N_11781,N_11406);
nand U12070 (N_12070,N_11411,N_11462);
nor U12071 (N_12071,N_11765,N_11608);
xnor U12072 (N_12072,N_11437,N_11562);
and U12073 (N_12073,N_11443,N_11426);
and U12074 (N_12074,N_11826,N_11684);
nand U12075 (N_12075,N_11856,N_11634);
nand U12076 (N_12076,N_11967,N_11546);
xor U12077 (N_12077,N_11736,N_11457);
or U12078 (N_12078,N_11872,N_11489);
nand U12079 (N_12079,N_11676,N_11542);
xor U12080 (N_12080,N_11796,N_11471);
nand U12081 (N_12081,N_11688,N_11773);
and U12082 (N_12082,N_11607,N_11797);
nor U12083 (N_12083,N_11746,N_11749);
and U12084 (N_12084,N_11757,N_11581);
xor U12085 (N_12085,N_11907,N_11464);
nand U12086 (N_12086,N_11660,N_11635);
xnor U12087 (N_12087,N_11540,N_11763);
xnor U12088 (N_12088,N_11571,N_11828);
and U12089 (N_12089,N_11778,N_11506);
nor U12090 (N_12090,N_11800,N_11852);
or U12091 (N_12091,N_11737,N_11724);
and U12092 (N_12092,N_11556,N_11754);
nor U12093 (N_12093,N_11547,N_11897);
nand U12094 (N_12094,N_11654,N_11458);
and U12095 (N_12095,N_11906,N_11971);
nand U12096 (N_12096,N_11990,N_11814);
nor U12097 (N_12097,N_11928,N_11811);
and U12098 (N_12098,N_11685,N_11890);
or U12099 (N_12099,N_11675,N_11439);
or U12100 (N_12100,N_11545,N_11616);
or U12101 (N_12101,N_11854,N_11667);
nand U12102 (N_12102,N_11977,N_11637);
or U12103 (N_12103,N_11483,N_11425);
nor U12104 (N_12104,N_11579,N_11424);
xor U12105 (N_12105,N_11845,N_11505);
and U12106 (N_12106,N_11815,N_11701);
nand U12107 (N_12107,N_11625,N_11905);
nor U12108 (N_12108,N_11576,N_11553);
xnor U12109 (N_12109,N_11972,N_11740);
xor U12110 (N_12110,N_11721,N_11577);
and U12111 (N_12111,N_11560,N_11593);
xor U12112 (N_12112,N_11973,N_11433);
nand U12113 (N_12113,N_11867,N_11421);
xor U12114 (N_12114,N_11966,N_11894);
nor U12115 (N_12115,N_11762,N_11570);
or U12116 (N_12116,N_11924,N_11944);
or U12117 (N_12117,N_11910,N_11803);
nor U12118 (N_12118,N_11788,N_11494);
and U12119 (N_12119,N_11729,N_11624);
or U12120 (N_12120,N_11987,N_11751);
or U12121 (N_12121,N_11617,N_11984);
and U12122 (N_12122,N_11687,N_11822);
xnor U12123 (N_12123,N_11524,N_11632);
and U12124 (N_12124,N_11900,N_11892);
or U12125 (N_12125,N_11525,N_11860);
xnor U12126 (N_12126,N_11991,N_11917);
nand U12127 (N_12127,N_11951,N_11950);
and U12128 (N_12128,N_11438,N_11414);
nor U12129 (N_12129,N_11422,N_11743);
nand U12130 (N_12130,N_11417,N_11651);
nand U12131 (N_12131,N_11768,N_11514);
nor U12132 (N_12132,N_11866,N_11707);
and U12133 (N_12133,N_11882,N_11509);
and U12134 (N_12134,N_11848,N_11595);
and U12135 (N_12135,N_11588,N_11718);
nand U12136 (N_12136,N_11487,N_11930);
nor U12137 (N_12137,N_11614,N_11952);
xnor U12138 (N_12138,N_11544,N_11650);
xnor U12139 (N_12139,N_11780,N_11731);
or U12140 (N_12140,N_11933,N_11831);
nor U12141 (N_12141,N_11441,N_11569);
nor U12142 (N_12142,N_11877,N_11722);
nor U12143 (N_12143,N_11705,N_11647);
and U12144 (N_12144,N_11779,N_11563);
xnor U12145 (N_12145,N_11620,N_11596);
nand U12146 (N_12146,N_11633,N_11709);
nor U12147 (N_12147,N_11683,N_11934);
and U12148 (N_12148,N_11567,N_11549);
and U12149 (N_12149,N_11913,N_11823);
or U12150 (N_12150,N_11612,N_11446);
or U12151 (N_12151,N_11698,N_11613);
nor U12152 (N_12152,N_11774,N_11594);
nor U12153 (N_12153,N_11918,N_11448);
nand U12154 (N_12154,N_11460,N_11630);
nor U12155 (N_12155,N_11618,N_11677);
xor U12156 (N_12156,N_11477,N_11573);
nand U12157 (N_12157,N_11817,N_11528);
and U12158 (N_12158,N_11454,N_11611);
nor U12159 (N_12159,N_11871,N_11469);
or U12160 (N_12160,N_11849,N_11761);
xnor U12161 (N_12161,N_11452,N_11558);
xor U12162 (N_12162,N_11475,N_11771);
nor U12163 (N_12163,N_11883,N_11652);
and U12164 (N_12164,N_11793,N_11482);
or U12165 (N_12165,N_11782,N_11767);
or U12166 (N_12166,N_11470,N_11753);
or U12167 (N_12167,N_11552,N_11794);
nand U12168 (N_12168,N_11583,N_11735);
and U12169 (N_12169,N_11695,N_11480);
nor U12170 (N_12170,N_11957,N_11444);
or U12171 (N_12171,N_11989,N_11655);
xor U12172 (N_12172,N_11490,N_11639);
and U12173 (N_12173,N_11898,N_11503);
xor U12174 (N_12174,N_11978,N_11837);
xor U12175 (N_12175,N_11747,N_11626);
xor U12176 (N_12176,N_11868,N_11517);
nand U12177 (N_12177,N_11473,N_11410);
nand U12178 (N_12178,N_11535,N_11519);
or U12179 (N_12179,N_11844,N_11993);
nand U12180 (N_12180,N_11597,N_11574);
or U12181 (N_12181,N_11732,N_11730);
nor U12182 (N_12182,N_11513,N_11980);
nand U12183 (N_12183,N_11716,N_11810);
nor U12184 (N_12184,N_11785,N_11861);
xor U12185 (N_12185,N_11420,N_11592);
or U12186 (N_12186,N_11586,N_11451);
nor U12187 (N_12187,N_11689,N_11879);
nor U12188 (N_12188,N_11997,N_11486);
xnor U12189 (N_12189,N_11712,N_11755);
or U12190 (N_12190,N_11598,N_11520);
and U12191 (N_12191,N_11880,N_11557);
or U12192 (N_12192,N_11842,N_11619);
nand U12193 (N_12193,N_11772,N_11696);
nor U12194 (N_12194,N_11601,N_11692);
nand U12195 (N_12195,N_11461,N_11566);
nand U12196 (N_12196,N_11518,N_11834);
or U12197 (N_12197,N_11564,N_11578);
nand U12198 (N_12198,N_11671,N_11589);
or U12199 (N_12199,N_11741,N_11955);
and U12200 (N_12200,N_11901,N_11419);
nand U12201 (N_12201,N_11832,N_11600);
xor U12202 (N_12202,N_11840,N_11784);
or U12203 (N_12203,N_11534,N_11551);
nand U12204 (N_12204,N_11491,N_11714);
and U12205 (N_12205,N_11673,N_11533);
xor U12206 (N_12206,N_11453,N_11526);
and U12207 (N_12207,N_11591,N_11976);
nand U12208 (N_12208,N_11646,N_11929);
nor U12209 (N_12209,N_11604,N_11682);
nor U12210 (N_12210,N_11603,N_11539);
and U12211 (N_12211,N_11631,N_11428);
xnor U12212 (N_12212,N_11497,N_11447);
nand U12213 (N_12213,N_11830,N_11713);
and U12214 (N_12214,N_11500,N_11493);
nor U12215 (N_12215,N_11942,N_11715);
nand U12216 (N_12216,N_11442,N_11416);
nor U12217 (N_12217,N_11656,N_11925);
nand U12218 (N_12218,N_11636,N_11904);
or U12219 (N_12219,N_11895,N_11902);
nand U12220 (N_12220,N_11996,N_11838);
nor U12221 (N_12221,N_11893,N_11459);
nor U12222 (N_12222,N_11402,N_11445);
or U12223 (N_12223,N_11981,N_11661);
and U12224 (N_12224,N_11436,N_11649);
nor U12225 (N_12225,N_11982,N_11405);
xnor U12226 (N_12226,N_11629,N_11723);
xnor U12227 (N_12227,N_11703,N_11759);
xnor U12228 (N_12228,N_11764,N_11615);
or U12229 (N_12229,N_11666,N_11559);
and U12230 (N_12230,N_11870,N_11523);
xnor U12231 (N_12231,N_11691,N_11532);
or U12232 (N_12232,N_11935,N_11787);
nor U12233 (N_12233,N_11511,N_11648);
and U12234 (N_12234,N_11792,N_11429);
or U12235 (N_12235,N_11865,N_11467);
xor U12236 (N_12236,N_11863,N_11507);
nor U12237 (N_12237,N_11643,N_11403);
or U12238 (N_12238,N_11449,N_11843);
or U12239 (N_12239,N_11404,N_11498);
xnor U12240 (N_12240,N_11998,N_11463);
nor U12241 (N_12241,N_11610,N_11875);
xor U12242 (N_12242,N_11599,N_11912);
xnor U12243 (N_12243,N_11821,N_11992);
xnor U12244 (N_12244,N_11653,N_11440);
nor U12245 (N_12245,N_11694,N_11674);
nor U12246 (N_12246,N_11502,N_11492);
nor U12247 (N_12247,N_11858,N_11869);
nor U12248 (N_12248,N_11775,N_11758);
nand U12249 (N_12249,N_11554,N_11921);
xnor U12250 (N_12250,N_11409,N_11969);
nor U12251 (N_12251,N_11415,N_11945);
xnor U12252 (N_12252,N_11949,N_11515);
nand U12253 (N_12253,N_11876,N_11530);
xnor U12254 (N_12254,N_11884,N_11681);
xor U12255 (N_12255,N_11548,N_11659);
nor U12256 (N_12256,N_11839,N_11853);
nor U12257 (N_12257,N_11465,N_11550);
nor U12258 (N_12258,N_11888,N_11527);
xnor U12259 (N_12259,N_11841,N_11820);
and U12260 (N_12260,N_11468,N_11846);
xnor U12261 (N_12261,N_11938,N_11590);
or U12262 (N_12262,N_11669,N_11748);
or U12263 (N_12263,N_11738,N_11941);
nand U12264 (N_12264,N_11899,N_11808);
nand U12265 (N_12265,N_11407,N_11423);
or U12266 (N_12266,N_11983,N_11418);
xnor U12267 (N_12267,N_11484,N_11622);
and U12268 (N_12268,N_11916,N_11859);
nand U12269 (N_12269,N_11742,N_11585);
nand U12270 (N_12270,N_11501,N_11937);
or U12271 (N_12271,N_11725,N_11510);
or U12272 (N_12272,N_11835,N_11795);
and U12273 (N_12273,N_11672,N_11668);
and U12274 (N_12274,N_11931,N_11756);
nor U12275 (N_12275,N_11943,N_11857);
xnor U12276 (N_12276,N_11538,N_11565);
xor U12277 (N_12277,N_11455,N_11887);
nor U12278 (N_12278,N_11974,N_11799);
or U12279 (N_12279,N_11807,N_11847);
nand U12280 (N_12280,N_11522,N_11642);
nand U12281 (N_12281,N_11536,N_11435);
or U12282 (N_12282,N_11995,N_11663);
nand U12283 (N_12283,N_11769,N_11720);
xnor U12284 (N_12284,N_11891,N_11628);
or U12285 (N_12285,N_11833,N_11456);
and U12286 (N_12286,N_11874,N_11836);
or U12287 (N_12287,N_11760,N_11948);
nand U12288 (N_12288,N_11508,N_11959);
or U12289 (N_12289,N_11704,N_11988);
nand U12290 (N_12290,N_11711,N_11885);
nor U12291 (N_12291,N_11798,N_11739);
nor U12292 (N_12292,N_11922,N_11572);
and U12293 (N_12293,N_11896,N_11750);
xor U12294 (N_12294,N_11881,N_11783);
xnor U12295 (N_12295,N_11408,N_11818);
and U12296 (N_12296,N_11479,N_11582);
or U12297 (N_12297,N_11531,N_11908);
nand U12298 (N_12298,N_11708,N_11638);
xnor U12299 (N_12299,N_11745,N_11700);
nor U12300 (N_12300,N_11856,N_11803);
nor U12301 (N_12301,N_11727,N_11638);
xor U12302 (N_12302,N_11422,N_11951);
or U12303 (N_12303,N_11772,N_11408);
and U12304 (N_12304,N_11750,N_11969);
nand U12305 (N_12305,N_11448,N_11703);
nor U12306 (N_12306,N_11881,N_11761);
nand U12307 (N_12307,N_11519,N_11743);
and U12308 (N_12308,N_11722,N_11459);
or U12309 (N_12309,N_11481,N_11853);
nand U12310 (N_12310,N_11431,N_11893);
nor U12311 (N_12311,N_11658,N_11719);
xor U12312 (N_12312,N_11947,N_11482);
xnor U12313 (N_12313,N_11637,N_11565);
and U12314 (N_12314,N_11520,N_11907);
xor U12315 (N_12315,N_11623,N_11552);
xor U12316 (N_12316,N_11423,N_11841);
or U12317 (N_12317,N_11436,N_11742);
nand U12318 (N_12318,N_11992,N_11979);
and U12319 (N_12319,N_11483,N_11939);
xnor U12320 (N_12320,N_11564,N_11496);
xnor U12321 (N_12321,N_11931,N_11543);
and U12322 (N_12322,N_11934,N_11770);
nor U12323 (N_12323,N_11795,N_11862);
xnor U12324 (N_12324,N_11582,N_11671);
xnor U12325 (N_12325,N_11871,N_11888);
and U12326 (N_12326,N_11509,N_11480);
xor U12327 (N_12327,N_11660,N_11986);
or U12328 (N_12328,N_11780,N_11421);
and U12329 (N_12329,N_11441,N_11628);
xor U12330 (N_12330,N_11799,N_11836);
xnor U12331 (N_12331,N_11789,N_11563);
nor U12332 (N_12332,N_11609,N_11547);
nor U12333 (N_12333,N_11406,N_11557);
xnor U12334 (N_12334,N_11773,N_11438);
nand U12335 (N_12335,N_11923,N_11750);
nand U12336 (N_12336,N_11657,N_11860);
or U12337 (N_12337,N_11767,N_11896);
and U12338 (N_12338,N_11979,N_11796);
nor U12339 (N_12339,N_11466,N_11448);
nand U12340 (N_12340,N_11950,N_11645);
nand U12341 (N_12341,N_11445,N_11492);
or U12342 (N_12342,N_11647,N_11866);
nand U12343 (N_12343,N_11596,N_11980);
and U12344 (N_12344,N_11511,N_11919);
and U12345 (N_12345,N_11753,N_11909);
nor U12346 (N_12346,N_11864,N_11729);
xnor U12347 (N_12347,N_11899,N_11774);
and U12348 (N_12348,N_11846,N_11669);
or U12349 (N_12349,N_11818,N_11450);
nand U12350 (N_12350,N_11798,N_11855);
nand U12351 (N_12351,N_11814,N_11742);
and U12352 (N_12352,N_11993,N_11889);
nor U12353 (N_12353,N_11488,N_11541);
xor U12354 (N_12354,N_11962,N_11499);
and U12355 (N_12355,N_11557,N_11776);
xnor U12356 (N_12356,N_11776,N_11404);
or U12357 (N_12357,N_11571,N_11948);
and U12358 (N_12358,N_11850,N_11773);
and U12359 (N_12359,N_11779,N_11437);
nor U12360 (N_12360,N_11934,N_11782);
nand U12361 (N_12361,N_11449,N_11478);
and U12362 (N_12362,N_11403,N_11958);
xor U12363 (N_12363,N_11794,N_11737);
nand U12364 (N_12364,N_11999,N_11609);
or U12365 (N_12365,N_11727,N_11533);
xor U12366 (N_12366,N_11930,N_11600);
nand U12367 (N_12367,N_11453,N_11765);
and U12368 (N_12368,N_11814,N_11633);
nand U12369 (N_12369,N_11725,N_11656);
or U12370 (N_12370,N_11407,N_11870);
or U12371 (N_12371,N_11859,N_11853);
xnor U12372 (N_12372,N_11671,N_11622);
or U12373 (N_12373,N_11547,N_11578);
or U12374 (N_12374,N_11912,N_11519);
or U12375 (N_12375,N_11549,N_11887);
nand U12376 (N_12376,N_11489,N_11824);
nand U12377 (N_12377,N_11684,N_11467);
nand U12378 (N_12378,N_11954,N_11571);
xnor U12379 (N_12379,N_11759,N_11770);
xor U12380 (N_12380,N_11452,N_11846);
nand U12381 (N_12381,N_11798,N_11889);
or U12382 (N_12382,N_11624,N_11902);
xor U12383 (N_12383,N_11900,N_11717);
nor U12384 (N_12384,N_11540,N_11638);
nor U12385 (N_12385,N_11456,N_11860);
nor U12386 (N_12386,N_11556,N_11806);
nor U12387 (N_12387,N_11931,N_11755);
and U12388 (N_12388,N_11572,N_11701);
xnor U12389 (N_12389,N_11870,N_11899);
nor U12390 (N_12390,N_11440,N_11739);
nand U12391 (N_12391,N_11474,N_11549);
or U12392 (N_12392,N_11920,N_11758);
and U12393 (N_12393,N_11662,N_11403);
nor U12394 (N_12394,N_11844,N_11992);
xnor U12395 (N_12395,N_11412,N_11541);
or U12396 (N_12396,N_11960,N_11553);
or U12397 (N_12397,N_11913,N_11654);
nor U12398 (N_12398,N_11977,N_11499);
and U12399 (N_12399,N_11761,N_11801);
and U12400 (N_12400,N_11802,N_11745);
or U12401 (N_12401,N_11636,N_11451);
and U12402 (N_12402,N_11884,N_11823);
nand U12403 (N_12403,N_11934,N_11884);
or U12404 (N_12404,N_11645,N_11729);
nand U12405 (N_12405,N_11489,N_11429);
or U12406 (N_12406,N_11737,N_11488);
xnor U12407 (N_12407,N_11527,N_11639);
xor U12408 (N_12408,N_11770,N_11562);
nand U12409 (N_12409,N_11898,N_11893);
nand U12410 (N_12410,N_11602,N_11436);
nand U12411 (N_12411,N_11891,N_11422);
or U12412 (N_12412,N_11795,N_11770);
nand U12413 (N_12413,N_11788,N_11723);
or U12414 (N_12414,N_11990,N_11823);
nor U12415 (N_12415,N_11855,N_11848);
or U12416 (N_12416,N_11980,N_11833);
xnor U12417 (N_12417,N_11651,N_11471);
nand U12418 (N_12418,N_11514,N_11465);
xnor U12419 (N_12419,N_11733,N_11437);
xnor U12420 (N_12420,N_11516,N_11826);
and U12421 (N_12421,N_11716,N_11859);
or U12422 (N_12422,N_11403,N_11883);
xnor U12423 (N_12423,N_11714,N_11690);
xor U12424 (N_12424,N_11854,N_11446);
nand U12425 (N_12425,N_11874,N_11607);
or U12426 (N_12426,N_11811,N_11806);
nor U12427 (N_12427,N_11430,N_11699);
nand U12428 (N_12428,N_11912,N_11712);
and U12429 (N_12429,N_11455,N_11409);
xor U12430 (N_12430,N_11920,N_11976);
nor U12431 (N_12431,N_11702,N_11477);
and U12432 (N_12432,N_11486,N_11520);
nor U12433 (N_12433,N_11895,N_11593);
or U12434 (N_12434,N_11648,N_11615);
xor U12435 (N_12435,N_11538,N_11959);
or U12436 (N_12436,N_11546,N_11410);
or U12437 (N_12437,N_11847,N_11695);
nor U12438 (N_12438,N_11656,N_11788);
and U12439 (N_12439,N_11955,N_11861);
nor U12440 (N_12440,N_11899,N_11418);
or U12441 (N_12441,N_11646,N_11455);
and U12442 (N_12442,N_11949,N_11616);
and U12443 (N_12443,N_11897,N_11444);
or U12444 (N_12444,N_11771,N_11726);
and U12445 (N_12445,N_11693,N_11817);
nand U12446 (N_12446,N_11497,N_11516);
or U12447 (N_12447,N_11415,N_11758);
nand U12448 (N_12448,N_11841,N_11452);
nor U12449 (N_12449,N_11805,N_11547);
or U12450 (N_12450,N_11485,N_11628);
or U12451 (N_12451,N_11438,N_11769);
nor U12452 (N_12452,N_11928,N_11433);
nand U12453 (N_12453,N_11855,N_11945);
nand U12454 (N_12454,N_11822,N_11633);
or U12455 (N_12455,N_11878,N_11560);
xor U12456 (N_12456,N_11905,N_11744);
or U12457 (N_12457,N_11697,N_11924);
or U12458 (N_12458,N_11498,N_11781);
nor U12459 (N_12459,N_11521,N_11476);
or U12460 (N_12460,N_11557,N_11402);
and U12461 (N_12461,N_11535,N_11692);
xnor U12462 (N_12462,N_11782,N_11916);
and U12463 (N_12463,N_11605,N_11844);
nor U12464 (N_12464,N_11985,N_11854);
or U12465 (N_12465,N_11768,N_11667);
xnor U12466 (N_12466,N_11420,N_11729);
or U12467 (N_12467,N_11893,N_11497);
nor U12468 (N_12468,N_11602,N_11960);
xor U12469 (N_12469,N_11587,N_11872);
and U12470 (N_12470,N_11703,N_11652);
xnor U12471 (N_12471,N_11707,N_11458);
nor U12472 (N_12472,N_11992,N_11425);
and U12473 (N_12473,N_11515,N_11731);
xnor U12474 (N_12474,N_11460,N_11533);
nor U12475 (N_12475,N_11673,N_11983);
nor U12476 (N_12476,N_11855,N_11834);
xnor U12477 (N_12477,N_11683,N_11930);
xor U12478 (N_12478,N_11428,N_11915);
nor U12479 (N_12479,N_11919,N_11498);
and U12480 (N_12480,N_11610,N_11448);
nand U12481 (N_12481,N_11635,N_11596);
nor U12482 (N_12482,N_11404,N_11405);
xor U12483 (N_12483,N_11959,N_11475);
nor U12484 (N_12484,N_11668,N_11504);
nor U12485 (N_12485,N_11416,N_11800);
xnor U12486 (N_12486,N_11507,N_11992);
nand U12487 (N_12487,N_11904,N_11447);
xnor U12488 (N_12488,N_11511,N_11942);
nand U12489 (N_12489,N_11516,N_11618);
nor U12490 (N_12490,N_11945,N_11426);
and U12491 (N_12491,N_11645,N_11736);
nand U12492 (N_12492,N_11819,N_11598);
nand U12493 (N_12493,N_11594,N_11909);
and U12494 (N_12494,N_11525,N_11973);
nand U12495 (N_12495,N_11543,N_11921);
xnor U12496 (N_12496,N_11460,N_11948);
nand U12497 (N_12497,N_11993,N_11515);
and U12498 (N_12498,N_11414,N_11441);
and U12499 (N_12499,N_11602,N_11774);
nor U12500 (N_12500,N_11669,N_11851);
or U12501 (N_12501,N_11654,N_11843);
nor U12502 (N_12502,N_11406,N_11889);
nand U12503 (N_12503,N_11654,N_11958);
xnor U12504 (N_12504,N_11422,N_11588);
nand U12505 (N_12505,N_11472,N_11776);
xor U12506 (N_12506,N_11441,N_11946);
or U12507 (N_12507,N_11509,N_11823);
nor U12508 (N_12508,N_11671,N_11908);
and U12509 (N_12509,N_11652,N_11483);
nor U12510 (N_12510,N_11895,N_11485);
nand U12511 (N_12511,N_11959,N_11496);
or U12512 (N_12512,N_11410,N_11421);
xor U12513 (N_12513,N_11578,N_11827);
nand U12514 (N_12514,N_11842,N_11559);
or U12515 (N_12515,N_11517,N_11407);
nor U12516 (N_12516,N_11877,N_11639);
and U12517 (N_12517,N_11919,N_11982);
xnor U12518 (N_12518,N_11479,N_11706);
and U12519 (N_12519,N_11678,N_11463);
xor U12520 (N_12520,N_11756,N_11475);
nand U12521 (N_12521,N_11836,N_11412);
xor U12522 (N_12522,N_11503,N_11965);
xnor U12523 (N_12523,N_11641,N_11814);
xor U12524 (N_12524,N_11687,N_11660);
nor U12525 (N_12525,N_11496,N_11649);
or U12526 (N_12526,N_11424,N_11942);
xnor U12527 (N_12527,N_11632,N_11522);
and U12528 (N_12528,N_11480,N_11952);
or U12529 (N_12529,N_11448,N_11803);
nand U12530 (N_12530,N_11433,N_11403);
xor U12531 (N_12531,N_11679,N_11580);
or U12532 (N_12532,N_11740,N_11612);
or U12533 (N_12533,N_11643,N_11910);
and U12534 (N_12534,N_11677,N_11819);
nand U12535 (N_12535,N_11863,N_11912);
nand U12536 (N_12536,N_11882,N_11933);
or U12537 (N_12537,N_11503,N_11978);
and U12538 (N_12538,N_11594,N_11601);
xor U12539 (N_12539,N_11466,N_11802);
nor U12540 (N_12540,N_11924,N_11820);
xor U12541 (N_12541,N_11526,N_11501);
xnor U12542 (N_12542,N_11545,N_11633);
or U12543 (N_12543,N_11904,N_11693);
xor U12544 (N_12544,N_11547,N_11999);
nor U12545 (N_12545,N_11756,N_11712);
or U12546 (N_12546,N_11550,N_11685);
nand U12547 (N_12547,N_11780,N_11412);
or U12548 (N_12548,N_11524,N_11883);
or U12549 (N_12549,N_11983,N_11908);
or U12550 (N_12550,N_11535,N_11561);
nor U12551 (N_12551,N_11470,N_11781);
and U12552 (N_12552,N_11978,N_11401);
nand U12553 (N_12553,N_11627,N_11876);
xor U12554 (N_12554,N_11654,N_11906);
or U12555 (N_12555,N_11694,N_11405);
or U12556 (N_12556,N_11503,N_11870);
nand U12557 (N_12557,N_11821,N_11410);
or U12558 (N_12558,N_11716,N_11985);
nand U12559 (N_12559,N_11766,N_11942);
nor U12560 (N_12560,N_11606,N_11592);
xnor U12561 (N_12561,N_11943,N_11803);
nand U12562 (N_12562,N_11729,N_11846);
and U12563 (N_12563,N_11612,N_11886);
and U12564 (N_12564,N_11987,N_11720);
and U12565 (N_12565,N_11988,N_11883);
nand U12566 (N_12566,N_11705,N_11868);
or U12567 (N_12567,N_11495,N_11895);
or U12568 (N_12568,N_11505,N_11689);
and U12569 (N_12569,N_11574,N_11661);
or U12570 (N_12570,N_11803,N_11531);
or U12571 (N_12571,N_11554,N_11873);
and U12572 (N_12572,N_11572,N_11702);
xor U12573 (N_12573,N_11490,N_11638);
nor U12574 (N_12574,N_11501,N_11557);
xor U12575 (N_12575,N_11423,N_11803);
xor U12576 (N_12576,N_11582,N_11508);
and U12577 (N_12577,N_11895,N_11479);
nor U12578 (N_12578,N_11633,N_11454);
and U12579 (N_12579,N_11902,N_11859);
nand U12580 (N_12580,N_11437,N_11847);
and U12581 (N_12581,N_11768,N_11854);
nand U12582 (N_12582,N_11881,N_11878);
nor U12583 (N_12583,N_11987,N_11801);
xnor U12584 (N_12584,N_11709,N_11508);
and U12585 (N_12585,N_11530,N_11880);
xnor U12586 (N_12586,N_11436,N_11927);
xor U12587 (N_12587,N_11967,N_11755);
xnor U12588 (N_12588,N_11727,N_11777);
and U12589 (N_12589,N_11884,N_11519);
or U12590 (N_12590,N_11970,N_11467);
xnor U12591 (N_12591,N_11609,N_11965);
or U12592 (N_12592,N_11875,N_11761);
or U12593 (N_12593,N_11991,N_11785);
and U12594 (N_12594,N_11864,N_11876);
xnor U12595 (N_12595,N_11452,N_11434);
or U12596 (N_12596,N_11916,N_11601);
nor U12597 (N_12597,N_11847,N_11758);
and U12598 (N_12598,N_11977,N_11505);
xnor U12599 (N_12599,N_11656,N_11457);
and U12600 (N_12600,N_12307,N_12440);
nand U12601 (N_12601,N_12163,N_12482);
xor U12602 (N_12602,N_12193,N_12271);
and U12603 (N_12603,N_12591,N_12558);
and U12604 (N_12604,N_12218,N_12075);
or U12605 (N_12605,N_12103,N_12403);
or U12606 (N_12606,N_12070,N_12287);
nor U12607 (N_12607,N_12593,N_12003);
or U12608 (N_12608,N_12044,N_12050);
or U12609 (N_12609,N_12568,N_12544);
xor U12610 (N_12610,N_12504,N_12013);
xnor U12611 (N_12611,N_12101,N_12205);
or U12612 (N_12612,N_12320,N_12132);
or U12613 (N_12613,N_12083,N_12134);
nand U12614 (N_12614,N_12356,N_12241);
nand U12615 (N_12615,N_12378,N_12268);
nor U12616 (N_12616,N_12485,N_12470);
and U12617 (N_12617,N_12308,N_12446);
and U12618 (N_12618,N_12093,N_12095);
nor U12619 (N_12619,N_12138,N_12459);
nand U12620 (N_12620,N_12563,N_12326);
or U12621 (N_12621,N_12305,N_12337);
nand U12622 (N_12622,N_12123,N_12561);
or U12623 (N_12623,N_12180,N_12110);
and U12624 (N_12624,N_12399,N_12435);
or U12625 (N_12625,N_12115,N_12158);
and U12626 (N_12626,N_12196,N_12588);
or U12627 (N_12627,N_12160,N_12582);
nand U12628 (N_12628,N_12031,N_12513);
nand U12629 (N_12629,N_12560,N_12579);
nor U12630 (N_12630,N_12144,N_12040);
or U12631 (N_12631,N_12049,N_12497);
nor U12632 (N_12632,N_12455,N_12245);
or U12633 (N_12633,N_12443,N_12082);
or U12634 (N_12634,N_12165,N_12157);
xnor U12635 (N_12635,N_12206,N_12397);
xnor U12636 (N_12636,N_12018,N_12359);
or U12637 (N_12637,N_12599,N_12436);
xor U12638 (N_12638,N_12100,N_12432);
nor U12639 (N_12639,N_12516,N_12267);
xnor U12640 (N_12640,N_12159,N_12032);
nor U12641 (N_12641,N_12025,N_12415);
or U12642 (N_12642,N_12086,N_12143);
and U12643 (N_12643,N_12188,N_12204);
and U12644 (N_12644,N_12189,N_12475);
xnor U12645 (N_12645,N_12057,N_12011);
or U12646 (N_12646,N_12358,N_12441);
nand U12647 (N_12647,N_12096,N_12171);
xnor U12648 (N_12648,N_12445,N_12312);
and U12649 (N_12649,N_12304,N_12195);
and U12650 (N_12650,N_12572,N_12332);
or U12651 (N_12651,N_12395,N_12221);
nor U12652 (N_12652,N_12448,N_12198);
xor U12653 (N_12653,N_12302,N_12152);
or U12654 (N_12654,N_12251,N_12087);
nand U12655 (N_12655,N_12369,N_12175);
or U12656 (N_12656,N_12000,N_12349);
xnor U12657 (N_12657,N_12249,N_12092);
xor U12658 (N_12658,N_12517,N_12421);
nor U12659 (N_12659,N_12061,N_12231);
nor U12660 (N_12660,N_12466,N_12429);
and U12661 (N_12661,N_12077,N_12004);
nor U12662 (N_12662,N_12148,N_12174);
nand U12663 (N_12663,N_12137,N_12037);
xor U12664 (N_12664,N_12376,N_12553);
or U12665 (N_12665,N_12139,N_12185);
xnor U12666 (N_12666,N_12564,N_12007);
xnor U12667 (N_12667,N_12129,N_12442);
nand U12668 (N_12668,N_12453,N_12434);
nand U12669 (N_12669,N_12041,N_12407);
or U12670 (N_12670,N_12454,N_12401);
nand U12671 (N_12671,N_12278,N_12480);
or U12672 (N_12672,N_12197,N_12255);
or U12673 (N_12673,N_12045,N_12089);
and U12674 (N_12674,N_12292,N_12094);
nand U12675 (N_12675,N_12541,N_12114);
or U12676 (N_12676,N_12507,N_12474);
nor U12677 (N_12677,N_12362,N_12364);
nor U12678 (N_12678,N_12254,N_12225);
nor U12679 (N_12679,N_12047,N_12106);
and U12680 (N_12680,N_12021,N_12472);
and U12681 (N_12681,N_12363,N_12514);
nand U12682 (N_12682,N_12012,N_12334);
nor U12683 (N_12683,N_12573,N_12024);
or U12684 (N_12684,N_12357,N_12091);
nor U12685 (N_12685,N_12353,N_12140);
xor U12686 (N_12686,N_12431,N_12203);
nor U12687 (N_12687,N_12065,N_12154);
xnor U12688 (N_12688,N_12523,N_12232);
and U12689 (N_12689,N_12272,N_12336);
xor U12690 (N_12690,N_12317,N_12284);
or U12691 (N_12691,N_12539,N_12084);
xor U12692 (N_12692,N_12394,N_12348);
or U12693 (N_12693,N_12515,N_12355);
nor U12694 (N_12694,N_12398,N_12405);
xor U12695 (N_12695,N_12492,N_12276);
and U12696 (N_12696,N_12277,N_12079);
nand U12697 (N_12697,N_12371,N_12595);
nand U12698 (N_12698,N_12496,N_12131);
or U12699 (N_12699,N_12210,N_12023);
nand U12700 (N_12700,N_12549,N_12019);
xnor U12701 (N_12701,N_12330,N_12104);
or U12702 (N_12702,N_12462,N_12053);
nor U12703 (N_12703,N_12263,N_12344);
or U12704 (N_12704,N_12461,N_12223);
and U12705 (N_12705,N_12486,N_12427);
nand U12706 (N_12706,N_12479,N_12379);
nand U12707 (N_12707,N_12450,N_12266);
nand U12708 (N_12708,N_12173,N_12176);
and U12709 (N_12709,N_12275,N_12183);
nand U12710 (N_12710,N_12166,N_12509);
or U12711 (N_12711,N_12338,N_12476);
nor U12712 (N_12712,N_12341,N_12048);
nor U12713 (N_12713,N_12130,N_12518);
xor U12714 (N_12714,N_12512,N_12335);
or U12715 (N_12715,N_12543,N_12471);
nor U12716 (N_12716,N_12238,N_12331);
xor U12717 (N_12717,N_12122,N_12488);
or U12718 (N_12718,N_12107,N_12527);
xor U12719 (N_12719,N_12162,N_12531);
or U12720 (N_12720,N_12499,N_12460);
nor U12721 (N_12721,N_12433,N_12002);
xnor U12722 (N_12722,N_12098,N_12033);
nor U12723 (N_12723,N_12182,N_12178);
nand U12724 (N_12724,N_12009,N_12283);
nor U12725 (N_12725,N_12124,N_12146);
xor U12726 (N_12726,N_12483,N_12316);
nor U12727 (N_12727,N_12298,N_12248);
and U12728 (N_12728,N_12246,N_12410);
nand U12729 (N_12729,N_12493,N_12102);
xnor U12730 (N_12730,N_12244,N_12309);
nor U12731 (N_12731,N_12256,N_12406);
nand U12732 (N_12732,N_12449,N_12285);
nand U12733 (N_12733,N_12511,N_12265);
xnor U12734 (N_12734,N_12554,N_12575);
nand U12735 (N_12735,N_12375,N_12141);
nor U12736 (N_12736,N_12001,N_12209);
xor U12737 (N_12737,N_12417,N_12169);
nand U12738 (N_12738,N_12522,N_12273);
or U12739 (N_12739,N_12027,N_12250);
nor U12740 (N_12740,N_12333,N_12351);
xor U12741 (N_12741,N_12022,N_12161);
nand U12742 (N_12742,N_12097,N_12329);
or U12743 (N_12743,N_12465,N_12199);
nor U12744 (N_12744,N_12192,N_12393);
nor U12745 (N_12745,N_12542,N_12062);
xor U12746 (N_12746,N_12313,N_12528);
xor U12747 (N_12747,N_12211,N_12212);
nor U12748 (N_12748,N_12236,N_12119);
nor U12749 (N_12749,N_12574,N_12444);
nand U12750 (N_12750,N_12490,N_12227);
nand U12751 (N_12751,N_12036,N_12237);
nor U12752 (N_12752,N_12402,N_12219);
nand U12753 (N_12753,N_12447,N_12319);
and U12754 (N_12754,N_12008,N_12396);
and U12755 (N_12755,N_12194,N_12301);
or U12756 (N_12756,N_12386,N_12350);
nand U12757 (N_12757,N_12294,N_12257);
nor U12758 (N_12758,N_12150,N_12280);
nand U12759 (N_12759,N_12252,N_12030);
or U12760 (N_12760,N_12584,N_12594);
or U12761 (N_12761,N_12533,N_12177);
nor U12762 (N_12762,N_12216,N_12015);
nor U12763 (N_12763,N_12073,N_12367);
or U12764 (N_12764,N_12133,N_12478);
nor U12765 (N_12765,N_12121,N_12566);
nor U12766 (N_12766,N_12260,N_12042);
or U12767 (N_12767,N_12167,N_12457);
or U12768 (N_12768,N_12262,N_12366);
or U12769 (N_12769,N_12290,N_12587);
and U12770 (N_12770,N_12063,N_12577);
and U12771 (N_12771,N_12506,N_12439);
or U12772 (N_12772,N_12422,N_12377);
xor U12773 (N_12773,N_12562,N_12072);
nor U12774 (N_12774,N_12530,N_12170);
nor U12775 (N_12775,N_12213,N_12099);
nor U12776 (N_12776,N_12214,N_12220);
and U12777 (N_12777,N_12535,N_12202);
or U12778 (N_12778,N_12014,N_12127);
and U12779 (N_12779,N_12519,N_12361);
nand U12780 (N_12780,N_12525,N_12108);
nand U12781 (N_12781,N_12058,N_12054);
or U12782 (N_12782,N_12570,N_12286);
xnor U12783 (N_12783,N_12325,N_12327);
nor U12784 (N_12784,N_12310,N_12229);
nand U12785 (N_12785,N_12253,N_12491);
nor U12786 (N_12786,N_12067,N_12296);
nand U12787 (N_12787,N_12400,N_12322);
and U12788 (N_12788,N_12311,N_12026);
nand U12789 (N_12789,N_12452,N_12164);
nor U12790 (N_12790,N_12464,N_12117);
nor U12791 (N_12791,N_12264,N_12306);
or U12792 (N_12792,N_12016,N_12473);
or U12793 (N_12793,N_12430,N_12051);
or U12794 (N_12794,N_12389,N_12583);
xor U12795 (N_12795,N_12555,N_12318);
nand U12796 (N_12796,N_12234,N_12424);
or U12797 (N_12797,N_12501,N_12038);
nor U12798 (N_12798,N_12571,N_12228);
nand U12799 (N_12799,N_12419,N_12112);
xor U12800 (N_12800,N_12113,N_12168);
xnor U12801 (N_12801,N_12384,N_12552);
nand U12802 (N_12802,N_12116,N_12391);
nand U12803 (N_12803,N_12181,N_12080);
nand U12804 (N_12804,N_12324,N_12388);
or U12805 (N_12805,N_12060,N_12315);
xnor U12806 (N_12806,N_12226,N_12346);
nand U12807 (N_12807,N_12293,N_12385);
and U12808 (N_12808,N_12589,N_12006);
nand U12809 (N_12809,N_12569,N_12020);
and U12810 (N_12810,N_12526,N_12428);
xnor U12811 (N_12811,N_12314,N_12387);
nor U12812 (N_12812,N_12261,N_12529);
xor U12813 (N_12813,N_12437,N_12423);
nand U12814 (N_12814,N_12043,N_12039);
xnor U12815 (N_12815,N_12145,N_12064);
and U12816 (N_12816,N_12365,N_12111);
xor U12817 (N_12817,N_12414,N_12556);
nor U12818 (N_12818,N_12597,N_12151);
or U12819 (N_12819,N_12208,N_12240);
nor U12820 (N_12820,N_12187,N_12532);
and U12821 (N_12821,N_12425,N_12586);
nor U12822 (N_12822,N_12536,N_12200);
xnor U12823 (N_12823,N_12592,N_12463);
nand U12824 (N_12824,N_12239,N_12495);
and U12825 (N_12825,N_12370,N_12297);
nor U12826 (N_12826,N_12372,N_12340);
or U12827 (N_12827,N_12380,N_12147);
nor U12828 (N_12828,N_12282,N_12413);
nand U12829 (N_12829,N_12247,N_12534);
xor U12830 (N_12830,N_12299,N_12494);
and U12831 (N_12831,N_12068,N_12081);
nor U12832 (N_12832,N_12550,N_12300);
nand U12833 (N_12833,N_12416,N_12230);
and U12834 (N_12834,N_12217,N_12545);
xor U12835 (N_12835,N_12418,N_12005);
nor U12836 (N_12836,N_12069,N_12510);
nand U12837 (N_12837,N_12017,N_12323);
and U12838 (N_12838,N_12179,N_12295);
nand U12839 (N_12839,N_12382,N_12078);
nand U12840 (N_12840,N_12347,N_12565);
nand U12841 (N_12841,N_12035,N_12125);
nor U12842 (N_12842,N_12489,N_12469);
nand U12843 (N_12843,N_12288,N_12088);
or U12844 (N_12844,N_12557,N_12508);
nor U12845 (N_12845,N_12059,N_12368);
nor U12846 (N_12846,N_12477,N_12224);
and U12847 (N_12847,N_12270,N_12590);
nand U12848 (N_12848,N_12155,N_12551);
or U12849 (N_12849,N_12052,N_12390);
nand U12850 (N_12850,N_12426,N_12343);
nor U12851 (N_12851,N_12411,N_12281);
nand U12852 (N_12852,N_12585,N_12328);
nand U12853 (N_12853,N_12259,N_12408);
xor U12854 (N_12854,N_12274,N_12136);
nand U12855 (N_12855,N_12354,N_12578);
xnor U12856 (N_12856,N_12269,N_12502);
or U12857 (N_12857,N_12374,N_12481);
nor U12858 (N_12858,N_12546,N_12242);
nor U12859 (N_12859,N_12321,N_12190);
nor U12860 (N_12860,N_12524,N_12596);
xnor U12861 (N_12861,N_12505,N_12105);
nor U12862 (N_12862,N_12207,N_12201);
nor U12863 (N_12863,N_12279,N_12235);
and U12864 (N_12864,N_12135,N_12420);
nor U12865 (N_12865,N_12373,N_12120);
nand U12866 (N_12866,N_12156,N_12046);
nor U12867 (N_12867,N_12258,N_12191);
nor U12868 (N_12868,N_12487,N_12503);
and U12869 (N_12869,N_12383,N_12109);
or U12870 (N_12870,N_12360,N_12128);
or U12871 (N_12871,N_12153,N_12458);
or U12872 (N_12872,N_12055,N_12456);
nand U12873 (N_12873,N_12451,N_12567);
nor U12874 (N_12874,N_12090,N_12029);
nor U12875 (N_12875,N_12484,N_12339);
nand U12876 (N_12876,N_12074,N_12559);
or U12877 (N_12877,N_12520,N_12303);
and U12878 (N_12878,N_12500,N_12381);
xor U12879 (N_12879,N_12034,N_12548);
and U12880 (N_12880,N_12468,N_12233);
xor U12881 (N_12881,N_12404,N_12184);
or U12882 (N_12882,N_12345,N_12056);
and U12883 (N_12883,N_12222,N_12467);
xnor U12884 (N_12884,N_12540,N_12172);
xnor U12885 (N_12885,N_12438,N_12118);
and U12886 (N_12886,N_12598,N_12215);
nor U12887 (N_12887,N_12412,N_12149);
or U12888 (N_12888,N_12010,N_12547);
nor U12889 (N_12889,N_12537,N_12581);
nor U12890 (N_12890,N_12085,N_12498);
or U12891 (N_12891,N_12342,N_12538);
nor U12892 (N_12892,N_12071,N_12066);
xor U12893 (N_12893,N_12142,N_12392);
and U12894 (N_12894,N_12186,N_12076);
or U12895 (N_12895,N_12521,N_12580);
nor U12896 (N_12896,N_12291,N_12243);
nor U12897 (N_12897,N_12028,N_12576);
or U12898 (N_12898,N_12126,N_12289);
nand U12899 (N_12899,N_12409,N_12352);
nor U12900 (N_12900,N_12094,N_12047);
and U12901 (N_12901,N_12238,N_12214);
xor U12902 (N_12902,N_12348,N_12205);
or U12903 (N_12903,N_12302,N_12051);
nand U12904 (N_12904,N_12439,N_12236);
nor U12905 (N_12905,N_12335,N_12006);
xnor U12906 (N_12906,N_12298,N_12140);
and U12907 (N_12907,N_12097,N_12217);
or U12908 (N_12908,N_12149,N_12353);
xor U12909 (N_12909,N_12284,N_12258);
or U12910 (N_12910,N_12564,N_12449);
nand U12911 (N_12911,N_12280,N_12117);
xnor U12912 (N_12912,N_12342,N_12192);
and U12913 (N_12913,N_12246,N_12519);
xor U12914 (N_12914,N_12053,N_12520);
xor U12915 (N_12915,N_12155,N_12262);
nor U12916 (N_12916,N_12335,N_12085);
xor U12917 (N_12917,N_12150,N_12012);
or U12918 (N_12918,N_12470,N_12017);
nor U12919 (N_12919,N_12560,N_12135);
and U12920 (N_12920,N_12301,N_12453);
and U12921 (N_12921,N_12249,N_12234);
and U12922 (N_12922,N_12235,N_12293);
xor U12923 (N_12923,N_12262,N_12362);
nand U12924 (N_12924,N_12199,N_12378);
xnor U12925 (N_12925,N_12530,N_12153);
nand U12926 (N_12926,N_12587,N_12009);
or U12927 (N_12927,N_12103,N_12174);
xnor U12928 (N_12928,N_12262,N_12517);
xnor U12929 (N_12929,N_12445,N_12428);
nand U12930 (N_12930,N_12151,N_12137);
nand U12931 (N_12931,N_12075,N_12440);
nor U12932 (N_12932,N_12519,N_12206);
nor U12933 (N_12933,N_12459,N_12176);
and U12934 (N_12934,N_12578,N_12379);
xor U12935 (N_12935,N_12367,N_12482);
xnor U12936 (N_12936,N_12382,N_12240);
xnor U12937 (N_12937,N_12088,N_12580);
xnor U12938 (N_12938,N_12289,N_12498);
xor U12939 (N_12939,N_12343,N_12300);
xor U12940 (N_12940,N_12548,N_12166);
xnor U12941 (N_12941,N_12333,N_12181);
nor U12942 (N_12942,N_12352,N_12003);
or U12943 (N_12943,N_12480,N_12113);
or U12944 (N_12944,N_12450,N_12403);
nand U12945 (N_12945,N_12494,N_12314);
and U12946 (N_12946,N_12295,N_12246);
nor U12947 (N_12947,N_12311,N_12075);
nand U12948 (N_12948,N_12257,N_12287);
and U12949 (N_12949,N_12492,N_12147);
or U12950 (N_12950,N_12110,N_12351);
and U12951 (N_12951,N_12380,N_12073);
and U12952 (N_12952,N_12243,N_12137);
or U12953 (N_12953,N_12525,N_12294);
nor U12954 (N_12954,N_12416,N_12481);
xnor U12955 (N_12955,N_12098,N_12228);
nand U12956 (N_12956,N_12581,N_12431);
xor U12957 (N_12957,N_12480,N_12090);
xnor U12958 (N_12958,N_12380,N_12225);
xnor U12959 (N_12959,N_12349,N_12213);
nand U12960 (N_12960,N_12327,N_12416);
or U12961 (N_12961,N_12554,N_12293);
and U12962 (N_12962,N_12368,N_12510);
and U12963 (N_12963,N_12037,N_12043);
nand U12964 (N_12964,N_12379,N_12006);
and U12965 (N_12965,N_12219,N_12287);
xor U12966 (N_12966,N_12181,N_12580);
or U12967 (N_12967,N_12395,N_12468);
nand U12968 (N_12968,N_12081,N_12409);
nand U12969 (N_12969,N_12581,N_12426);
xnor U12970 (N_12970,N_12355,N_12566);
xor U12971 (N_12971,N_12121,N_12457);
and U12972 (N_12972,N_12105,N_12411);
or U12973 (N_12973,N_12573,N_12439);
nor U12974 (N_12974,N_12268,N_12036);
xor U12975 (N_12975,N_12367,N_12355);
or U12976 (N_12976,N_12583,N_12090);
nor U12977 (N_12977,N_12030,N_12472);
xnor U12978 (N_12978,N_12578,N_12573);
nand U12979 (N_12979,N_12268,N_12505);
xor U12980 (N_12980,N_12562,N_12351);
and U12981 (N_12981,N_12152,N_12270);
or U12982 (N_12982,N_12409,N_12091);
and U12983 (N_12983,N_12222,N_12155);
nand U12984 (N_12984,N_12128,N_12207);
nor U12985 (N_12985,N_12415,N_12020);
or U12986 (N_12986,N_12523,N_12312);
nand U12987 (N_12987,N_12507,N_12135);
or U12988 (N_12988,N_12115,N_12320);
and U12989 (N_12989,N_12451,N_12057);
nand U12990 (N_12990,N_12120,N_12242);
nor U12991 (N_12991,N_12131,N_12492);
or U12992 (N_12992,N_12507,N_12361);
and U12993 (N_12993,N_12325,N_12548);
nand U12994 (N_12994,N_12521,N_12233);
xor U12995 (N_12995,N_12263,N_12153);
xor U12996 (N_12996,N_12162,N_12054);
or U12997 (N_12997,N_12536,N_12583);
nor U12998 (N_12998,N_12261,N_12143);
and U12999 (N_12999,N_12294,N_12412);
nand U13000 (N_13000,N_12311,N_12297);
nand U13001 (N_13001,N_12438,N_12444);
and U13002 (N_13002,N_12463,N_12445);
xnor U13003 (N_13003,N_12082,N_12257);
nand U13004 (N_13004,N_12419,N_12287);
xnor U13005 (N_13005,N_12439,N_12486);
nor U13006 (N_13006,N_12228,N_12014);
xor U13007 (N_13007,N_12274,N_12239);
or U13008 (N_13008,N_12548,N_12336);
and U13009 (N_13009,N_12127,N_12404);
nand U13010 (N_13010,N_12506,N_12557);
and U13011 (N_13011,N_12043,N_12271);
xnor U13012 (N_13012,N_12053,N_12138);
or U13013 (N_13013,N_12553,N_12509);
or U13014 (N_13014,N_12181,N_12330);
nor U13015 (N_13015,N_12443,N_12264);
and U13016 (N_13016,N_12061,N_12411);
nor U13017 (N_13017,N_12407,N_12477);
xnor U13018 (N_13018,N_12313,N_12530);
and U13019 (N_13019,N_12031,N_12300);
or U13020 (N_13020,N_12481,N_12434);
or U13021 (N_13021,N_12437,N_12242);
or U13022 (N_13022,N_12031,N_12427);
nor U13023 (N_13023,N_12146,N_12048);
xnor U13024 (N_13024,N_12578,N_12417);
xnor U13025 (N_13025,N_12475,N_12568);
nand U13026 (N_13026,N_12371,N_12388);
nor U13027 (N_13027,N_12436,N_12043);
xnor U13028 (N_13028,N_12175,N_12456);
and U13029 (N_13029,N_12280,N_12446);
and U13030 (N_13030,N_12482,N_12236);
nor U13031 (N_13031,N_12116,N_12031);
and U13032 (N_13032,N_12520,N_12557);
nor U13033 (N_13033,N_12400,N_12326);
nor U13034 (N_13034,N_12591,N_12441);
and U13035 (N_13035,N_12522,N_12349);
nor U13036 (N_13036,N_12093,N_12182);
nor U13037 (N_13037,N_12102,N_12261);
nand U13038 (N_13038,N_12309,N_12324);
nand U13039 (N_13039,N_12331,N_12042);
or U13040 (N_13040,N_12074,N_12242);
xor U13041 (N_13041,N_12061,N_12424);
nand U13042 (N_13042,N_12314,N_12526);
or U13043 (N_13043,N_12491,N_12252);
or U13044 (N_13044,N_12426,N_12510);
nand U13045 (N_13045,N_12213,N_12255);
xnor U13046 (N_13046,N_12090,N_12085);
nor U13047 (N_13047,N_12057,N_12382);
or U13048 (N_13048,N_12433,N_12240);
nor U13049 (N_13049,N_12413,N_12418);
nand U13050 (N_13050,N_12377,N_12284);
xnor U13051 (N_13051,N_12412,N_12122);
and U13052 (N_13052,N_12579,N_12166);
and U13053 (N_13053,N_12030,N_12587);
nor U13054 (N_13054,N_12210,N_12018);
or U13055 (N_13055,N_12099,N_12344);
nand U13056 (N_13056,N_12266,N_12506);
nand U13057 (N_13057,N_12367,N_12005);
xnor U13058 (N_13058,N_12323,N_12039);
xor U13059 (N_13059,N_12561,N_12360);
xor U13060 (N_13060,N_12299,N_12409);
and U13061 (N_13061,N_12258,N_12522);
and U13062 (N_13062,N_12037,N_12259);
nand U13063 (N_13063,N_12110,N_12587);
or U13064 (N_13064,N_12043,N_12401);
nand U13065 (N_13065,N_12462,N_12247);
and U13066 (N_13066,N_12301,N_12210);
nand U13067 (N_13067,N_12579,N_12522);
nand U13068 (N_13068,N_12456,N_12376);
or U13069 (N_13069,N_12536,N_12112);
or U13070 (N_13070,N_12156,N_12341);
nor U13071 (N_13071,N_12396,N_12568);
or U13072 (N_13072,N_12353,N_12399);
or U13073 (N_13073,N_12505,N_12166);
or U13074 (N_13074,N_12240,N_12087);
nor U13075 (N_13075,N_12338,N_12192);
xor U13076 (N_13076,N_12326,N_12203);
or U13077 (N_13077,N_12264,N_12291);
xor U13078 (N_13078,N_12090,N_12124);
nor U13079 (N_13079,N_12121,N_12489);
xor U13080 (N_13080,N_12506,N_12201);
nand U13081 (N_13081,N_12249,N_12123);
nand U13082 (N_13082,N_12547,N_12546);
and U13083 (N_13083,N_12104,N_12556);
nand U13084 (N_13084,N_12572,N_12329);
or U13085 (N_13085,N_12592,N_12596);
nand U13086 (N_13086,N_12579,N_12094);
nor U13087 (N_13087,N_12227,N_12495);
nor U13088 (N_13088,N_12326,N_12321);
nor U13089 (N_13089,N_12556,N_12337);
or U13090 (N_13090,N_12378,N_12338);
or U13091 (N_13091,N_12181,N_12037);
and U13092 (N_13092,N_12174,N_12593);
xnor U13093 (N_13093,N_12268,N_12491);
xor U13094 (N_13094,N_12277,N_12564);
and U13095 (N_13095,N_12407,N_12428);
xor U13096 (N_13096,N_12482,N_12285);
and U13097 (N_13097,N_12169,N_12282);
or U13098 (N_13098,N_12107,N_12353);
or U13099 (N_13099,N_12240,N_12420);
and U13100 (N_13100,N_12131,N_12351);
nor U13101 (N_13101,N_12405,N_12048);
nor U13102 (N_13102,N_12279,N_12347);
xor U13103 (N_13103,N_12052,N_12518);
nor U13104 (N_13104,N_12342,N_12420);
and U13105 (N_13105,N_12437,N_12486);
and U13106 (N_13106,N_12087,N_12525);
or U13107 (N_13107,N_12379,N_12420);
nor U13108 (N_13108,N_12366,N_12282);
and U13109 (N_13109,N_12571,N_12381);
nor U13110 (N_13110,N_12250,N_12184);
nand U13111 (N_13111,N_12537,N_12114);
and U13112 (N_13112,N_12329,N_12578);
or U13113 (N_13113,N_12190,N_12358);
and U13114 (N_13114,N_12052,N_12395);
or U13115 (N_13115,N_12385,N_12161);
nor U13116 (N_13116,N_12581,N_12189);
and U13117 (N_13117,N_12059,N_12167);
nand U13118 (N_13118,N_12450,N_12199);
xor U13119 (N_13119,N_12047,N_12399);
nor U13120 (N_13120,N_12240,N_12031);
nor U13121 (N_13121,N_12154,N_12101);
nor U13122 (N_13122,N_12199,N_12316);
xor U13123 (N_13123,N_12329,N_12204);
and U13124 (N_13124,N_12164,N_12035);
xor U13125 (N_13125,N_12237,N_12284);
and U13126 (N_13126,N_12341,N_12575);
nand U13127 (N_13127,N_12394,N_12516);
or U13128 (N_13128,N_12509,N_12123);
nor U13129 (N_13129,N_12303,N_12126);
or U13130 (N_13130,N_12555,N_12255);
or U13131 (N_13131,N_12596,N_12525);
xor U13132 (N_13132,N_12284,N_12337);
and U13133 (N_13133,N_12069,N_12595);
nand U13134 (N_13134,N_12103,N_12441);
nor U13135 (N_13135,N_12175,N_12493);
nand U13136 (N_13136,N_12180,N_12552);
or U13137 (N_13137,N_12452,N_12068);
and U13138 (N_13138,N_12319,N_12431);
and U13139 (N_13139,N_12016,N_12413);
xnor U13140 (N_13140,N_12364,N_12297);
or U13141 (N_13141,N_12482,N_12378);
and U13142 (N_13142,N_12091,N_12394);
nand U13143 (N_13143,N_12548,N_12346);
nor U13144 (N_13144,N_12288,N_12461);
nand U13145 (N_13145,N_12022,N_12248);
nand U13146 (N_13146,N_12397,N_12598);
or U13147 (N_13147,N_12112,N_12119);
nor U13148 (N_13148,N_12196,N_12173);
nor U13149 (N_13149,N_12386,N_12004);
xnor U13150 (N_13150,N_12000,N_12486);
or U13151 (N_13151,N_12065,N_12159);
nand U13152 (N_13152,N_12550,N_12359);
nand U13153 (N_13153,N_12292,N_12488);
xnor U13154 (N_13154,N_12014,N_12008);
or U13155 (N_13155,N_12272,N_12429);
and U13156 (N_13156,N_12336,N_12056);
or U13157 (N_13157,N_12355,N_12009);
nand U13158 (N_13158,N_12192,N_12521);
and U13159 (N_13159,N_12226,N_12435);
and U13160 (N_13160,N_12263,N_12296);
and U13161 (N_13161,N_12002,N_12208);
xnor U13162 (N_13162,N_12476,N_12010);
and U13163 (N_13163,N_12567,N_12066);
xnor U13164 (N_13164,N_12021,N_12369);
xnor U13165 (N_13165,N_12063,N_12076);
and U13166 (N_13166,N_12135,N_12460);
xnor U13167 (N_13167,N_12025,N_12044);
and U13168 (N_13168,N_12185,N_12299);
nand U13169 (N_13169,N_12397,N_12372);
and U13170 (N_13170,N_12438,N_12256);
xor U13171 (N_13171,N_12257,N_12485);
nor U13172 (N_13172,N_12134,N_12405);
nor U13173 (N_13173,N_12085,N_12113);
or U13174 (N_13174,N_12360,N_12396);
xnor U13175 (N_13175,N_12592,N_12471);
nor U13176 (N_13176,N_12171,N_12291);
xnor U13177 (N_13177,N_12466,N_12478);
nor U13178 (N_13178,N_12245,N_12473);
and U13179 (N_13179,N_12157,N_12436);
nand U13180 (N_13180,N_12065,N_12057);
nand U13181 (N_13181,N_12521,N_12179);
and U13182 (N_13182,N_12161,N_12049);
nor U13183 (N_13183,N_12261,N_12097);
nand U13184 (N_13184,N_12380,N_12509);
xor U13185 (N_13185,N_12327,N_12580);
and U13186 (N_13186,N_12508,N_12427);
xnor U13187 (N_13187,N_12116,N_12328);
nor U13188 (N_13188,N_12395,N_12230);
or U13189 (N_13189,N_12120,N_12059);
or U13190 (N_13190,N_12598,N_12379);
xnor U13191 (N_13191,N_12254,N_12505);
nor U13192 (N_13192,N_12445,N_12443);
xnor U13193 (N_13193,N_12577,N_12251);
nand U13194 (N_13194,N_12066,N_12459);
nand U13195 (N_13195,N_12489,N_12009);
xnor U13196 (N_13196,N_12564,N_12092);
xor U13197 (N_13197,N_12257,N_12421);
and U13198 (N_13198,N_12129,N_12423);
xor U13199 (N_13199,N_12027,N_12354);
nand U13200 (N_13200,N_12912,N_12941);
nor U13201 (N_13201,N_12781,N_13163);
nor U13202 (N_13202,N_13188,N_12614);
and U13203 (N_13203,N_13077,N_12718);
nand U13204 (N_13204,N_12782,N_12814);
xor U13205 (N_13205,N_12848,N_12921);
nor U13206 (N_13206,N_12974,N_13183);
nand U13207 (N_13207,N_12824,N_13113);
xnor U13208 (N_13208,N_12706,N_12699);
nor U13209 (N_13209,N_13018,N_12661);
or U13210 (N_13210,N_12634,N_12864);
xnor U13211 (N_13211,N_12958,N_13051);
and U13212 (N_13212,N_12601,N_13123);
nor U13213 (N_13213,N_12820,N_12847);
nor U13214 (N_13214,N_13076,N_12604);
or U13215 (N_13215,N_13100,N_13120);
or U13216 (N_13216,N_13105,N_13061);
nor U13217 (N_13217,N_12806,N_13191);
xor U13218 (N_13218,N_12966,N_13186);
nand U13219 (N_13219,N_13132,N_13166);
xor U13220 (N_13220,N_12929,N_13092);
and U13221 (N_13221,N_12896,N_13124);
nor U13222 (N_13222,N_13145,N_12995);
or U13223 (N_13223,N_13146,N_12705);
xnor U13224 (N_13224,N_13083,N_12830);
xor U13225 (N_13225,N_12952,N_12967);
or U13226 (N_13226,N_12815,N_13174);
xor U13227 (N_13227,N_12660,N_13025);
xnor U13228 (N_13228,N_12887,N_12905);
or U13229 (N_13229,N_13130,N_12695);
nand U13230 (N_13230,N_13161,N_13023);
nor U13231 (N_13231,N_12858,N_12642);
or U13232 (N_13232,N_12882,N_13171);
and U13233 (N_13233,N_12656,N_13015);
or U13234 (N_13234,N_12652,N_13040);
and U13235 (N_13235,N_13032,N_13075);
nor U13236 (N_13236,N_12627,N_13164);
nand U13237 (N_13237,N_12962,N_12742);
xor U13238 (N_13238,N_12648,N_12777);
nor U13239 (N_13239,N_12790,N_12846);
or U13240 (N_13240,N_13139,N_13176);
xnor U13241 (N_13241,N_13177,N_12982);
or U13242 (N_13242,N_12667,N_12681);
or U13243 (N_13243,N_12850,N_12776);
or U13244 (N_13244,N_13080,N_13147);
or U13245 (N_13245,N_13064,N_13005);
and U13246 (N_13246,N_12693,N_13106);
nor U13247 (N_13247,N_13110,N_13059);
or U13248 (N_13248,N_12877,N_13078);
xor U13249 (N_13249,N_13199,N_13062);
or U13250 (N_13250,N_12791,N_12712);
or U13251 (N_13251,N_12602,N_13019);
and U13252 (N_13252,N_12906,N_13028);
nor U13253 (N_13253,N_12978,N_12639);
xor U13254 (N_13254,N_12630,N_13006);
nand U13255 (N_13255,N_13138,N_13141);
or U13256 (N_13256,N_13049,N_12694);
or U13257 (N_13257,N_12725,N_12653);
nand U13258 (N_13258,N_12907,N_12988);
nand U13259 (N_13259,N_12881,N_12828);
and U13260 (N_13260,N_13085,N_13156);
or U13261 (N_13261,N_13116,N_12747);
and U13262 (N_13262,N_12735,N_12943);
xor U13263 (N_13263,N_13185,N_12731);
nand U13264 (N_13264,N_13112,N_13095);
xnor U13265 (N_13265,N_12924,N_12893);
nand U13266 (N_13266,N_12947,N_12778);
nand U13267 (N_13267,N_13155,N_12779);
xor U13268 (N_13268,N_13187,N_12857);
nand U13269 (N_13269,N_12873,N_12679);
nand U13270 (N_13270,N_13071,N_13068);
nand U13271 (N_13271,N_13194,N_12964);
and U13272 (N_13272,N_12972,N_13158);
and U13273 (N_13273,N_12839,N_12672);
xor U13274 (N_13274,N_12853,N_13157);
or U13275 (N_13275,N_12981,N_12913);
nor U13276 (N_13276,N_12620,N_12700);
or U13277 (N_13277,N_13197,N_12714);
nand U13278 (N_13278,N_12757,N_12840);
xor U13279 (N_13279,N_12668,N_13087);
or U13280 (N_13280,N_12788,N_12826);
xor U13281 (N_13281,N_12861,N_12666);
nand U13282 (N_13282,N_12741,N_12698);
or U13283 (N_13283,N_12629,N_13024);
or U13284 (N_13284,N_12745,N_12686);
nor U13285 (N_13285,N_12810,N_13125);
and U13286 (N_13286,N_12692,N_12944);
and U13287 (N_13287,N_13043,N_12968);
or U13288 (N_13288,N_13081,N_12608);
xnor U13289 (N_13289,N_12677,N_13119);
nor U13290 (N_13290,N_13126,N_12662);
nor U13291 (N_13291,N_13091,N_12934);
and U13292 (N_13292,N_13039,N_12876);
and U13293 (N_13293,N_12751,N_13181);
or U13294 (N_13294,N_12697,N_12983);
and U13295 (N_13295,N_13063,N_12622);
and U13296 (N_13296,N_13094,N_13111);
nand U13297 (N_13297,N_13060,N_13152);
xnor U13298 (N_13298,N_12657,N_12902);
nand U13299 (N_13299,N_13027,N_12768);
and U13300 (N_13300,N_12991,N_12770);
xor U13301 (N_13301,N_12856,N_12923);
nand U13302 (N_13302,N_12859,N_12865);
xor U13303 (N_13303,N_12663,N_12603);
xnor U13304 (N_13304,N_12960,N_13122);
nand U13305 (N_13305,N_12640,N_13137);
nand U13306 (N_13306,N_13021,N_12899);
nand U13307 (N_13307,N_12746,N_12628);
nand U13308 (N_13308,N_12959,N_13096);
nor U13309 (N_13309,N_13117,N_12842);
or U13310 (N_13310,N_12726,N_13131);
xor U13311 (N_13311,N_13148,N_12973);
and U13312 (N_13312,N_12756,N_12739);
nand U13313 (N_13313,N_12932,N_13001);
xor U13314 (N_13314,N_12678,N_13048);
nor U13315 (N_13315,N_12612,N_13151);
or U13316 (N_13316,N_12794,N_12797);
xnor U13317 (N_13317,N_13196,N_13073);
nand U13318 (N_13318,N_12682,N_12691);
nand U13319 (N_13319,N_12975,N_12910);
or U13320 (N_13320,N_12619,N_13057);
nor U13321 (N_13321,N_13162,N_12792);
or U13322 (N_13322,N_12615,N_13102);
and U13323 (N_13323,N_12898,N_13114);
xor U13324 (N_13324,N_13144,N_13056);
xor U13325 (N_13325,N_12970,N_12780);
and U13326 (N_13326,N_12939,N_12606);
nor U13327 (N_13327,N_13090,N_12651);
nand U13328 (N_13328,N_12733,N_13031);
nand U13329 (N_13329,N_12696,N_12727);
xor U13330 (N_13330,N_12675,N_12811);
nand U13331 (N_13331,N_12673,N_12940);
nand U13332 (N_13332,N_13029,N_12827);
nand U13333 (N_13333,N_13093,N_13115);
xnor U13334 (N_13334,N_13010,N_13189);
nor U13335 (N_13335,N_12717,N_13045);
nand U13336 (N_13336,N_13067,N_12774);
or U13337 (N_13337,N_12875,N_13182);
and U13338 (N_13338,N_13030,N_13101);
nand U13339 (N_13339,N_13099,N_12720);
xor U13340 (N_13340,N_12644,N_12605);
nand U13341 (N_13341,N_13150,N_13153);
nand U13342 (N_13342,N_12843,N_12948);
or U13343 (N_13343,N_12909,N_12834);
xor U13344 (N_13344,N_12795,N_13170);
nor U13345 (N_13345,N_12759,N_13033);
xnor U13346 (N_13346,N_12665,N_12637);
and U13347 (N_13347,N_13014,N_12938);
or U13348 (N_13348,N_12617,N_12680);
nor U13349 (N_13349,N_12734,N_13172);
nand U13350 (N_13350,N_12635,N_12730);
xor U13351 (N_13351,N_12738,N_13046);
or U13352 (N_13352,N_12710,N_13074);
nor U13353 (N_13353,N_12674,N_13097);
and U13354 (N_13354,N_13178,N_12796);
nor U13355 (N_13355,N_12645,N_12946);
nor U13356 (N_13356,N_12748,N_12928);
nand U13357 (N_13357,N_13160,N_12987);
nor U13358 (N_13358,N_12767,N_13193);
or U13359 (N_13359,N_12872,N_13053);
nand U13360 (N_13360,N_12892,N_12953);
xnor U13361 (N_13361,N_12916,N_12744);
nor U13362 (N_13362,N_13044,N_13104);
xnor U13363 (N_13363,N_13195,N_12999);
or U13364 (N_13364,N_12787,N_12769);
nand U13365 (N_13365,N_12880,N_12819);
or U13366 (N_13366,N_13017,N_12927);
or U13367 (N_13367,N_12990,N_13107);
and U13368 (N_13368,N_12989,N_12931);
xor U13369 (N_13369,N_12849,N_12807);
xnor U13370 (N_13370,N_13084,N_13037);
nand U13371 (N_13371,N_12930,N_12996);
or U13372 (N_13372,N_12954,N_12891);
xor U13373 (N_13373,N_13020,N_12998);
nor U13374 (N_13374,N_12878,N_12701);
nor U13375 (N_13375,N_12707,N_13069);
and U13376 (N_13376,N_13052,N_12789);
or U13377 (N_13377,N_12646,N_13175);
and U13378 (N_13378,N_13003,N_12979);
nor U13379 (N_13379,N_12659,N_12841);
xnor U13380 (N_13380,N_12736,N_12754);
and U13381 (N_13381,N_12676,N_12831);
xor U13382 (N_13382,N_12869,N_13066);
or U13383 (N_13383,N_13086,N_12874);
xor U13384 (N_13384,N_12749,N_12838);
xnor U13385 (N_13385,N_12715,N_12955);
nand U13386 (N_13386,N_13184,N_12925);
xor U13387 (N_13387,N_12808,N_12713);
xor U13388 (N_13388,N_12616,N_12821);
or U13389 (N_13389,N_13149,N_12851);
nor U13390 (N_13390,N_12980,N_12845);
or U13391 (N_13391,N_13159,N_12740);
nor U13392 (N_13392,N_12649,N_12702);
or U13393 (N_13393,N_13173,N_12613);
xnor U13394 (N_13394,N_12610,N_12772);
and U13395 (N_13395,N_12817,N_12920);
nand U13396 (N_13396,N_13180,N_13108);
or U13397 (N_13397,N_13072,N_12993);
or U13398 (N_13398,N_12836,N_12632);
nand U13399 (N_13399,N_12723,N_12854);
nand U13400 (N_13400,N_12658,N_12753);
xor U13401 (N_13401,N_12607,N_12655);
nand U13402 (N_13402,N_13169,N_12965);
and U13403 (N_13403,N_13002,N_12600);
nor U13404 (N_13404,N_12901,N_13167);
xor U13405 (N_13405,N_12800,N_13136);
or U13406 (N_13406,N_12870,N_12886);
or U13407 (N_13407,N_12863,N_12883);
nor U13408 (N_13408,N_12625,N_13098);
nand U13409 (N_13409,N_12957,N_12922);
nand U13410 (N_13410,N_12915,N_12623);
nor U13411 (N_13411,N_12631,N_12908);
xor U13412 (N_13412,N_12728,N_12664);
or U13413 (N_13413,N_12911,N_12650);
or U13414 (N_13414,N_12670,N_12773);
nand U13415 (N_13415,N_13026,N_12812);
and U13416 (N_13416,N_12885,N_13013);
and U13417 (N_13417,N_13089,N_12683);
nor U13418 (N_13418,N_13103,N_12813);
nor U13419 (N_13419,N_13042,N_13088);
and U13420 (N_13420,N_12684,N_12784);
xnor U13421 (N_13421,N_12709,N_12862);
or U13422 (N_13422,N_12889,N_12937);
xor U13423 (N_13423,N_12933,N_13054);
nor U13424 (N_13424,N_13036,N_12798);
or U13425 (N_13425,N_13022,N_12618);
or U13426 (N_13426,N_13007,N_12956);
and U13427 (N_13427,N_12994,N_12685);
nand U13428 (N_13428,N_12866,N_13121);
or U13429 (N_13429,N_12837,N_13008);
nor U13430 (N_13430,N_13109,N_12722);
nor U13431 (N_13431,N_12708,N_12833);
xor U13432 (N_13432,N_12626,N_13134);
or U13433 (N_13433,N_12844,N_12961);
nor U13434 (N_13434,N_13034,N_12816);
xor U13435 (N_13435,N_12903,N_13009);
nand U13436 (N_13436,N_13168,N_13058);
or U13437 (N_13437,N_12624,N_12763);
nor U13438 (N_13438,N_12732,N_12969);
or U13439 (N_13439,N_12823,N_12690);
nor U13440 (N_13440,N_12647,N_12633);
and U13441 (N_13441,N_12805,N_12765);
xor U13442 (N_13442,N_12719,N_12868);
or U13443 (N_13443,N_12704,N_12802);
nor U13444 (N_13444,N_13011,N_12724);
and U13445 (N_13445,N_13179,N_12786);
nor U13446 (N_13446,N_12766,N_12771);
and U13447 (N_13447,N_12867,N_12783);
xnor U13448 (N_13448,N_13135,N_13129);
nand U13449 (N_13449,N_12638,N_13050);
xor U13450 (N_13450,N_13079,N_12755);
and U13451 (N_13451,N_12992,N_13154);
and U13452 (N_13452,N_12703,N_12643);
nand U13453 (N_13453,N_12871,N_12621);
or U13454 (N_13454,N_12895,N_13055);
and U13455 (N_13455,N_12945,N_12793);
nand U13456 (N_13456,N_12818,N_13198);
and U13457 (N_13457,N_12669,N_12799);
and U13458 (N_13458,N_13016,N_12986);
nand U13459 (N_13459,N_12809,N_13038);
nand U13460 (N_13460,N_12985,N_12904);
and U13461 (N_13461,N_12888,N_12884);
nand U13462 (N_13462,N_13128,N_12926);
nand U13463 (N_13463,N_12919,N_13041);
and U13464 (N_13464,N_12801,N_13004);
xor U13465 (N_13465,N_12829,N_12654);
or U13466 (N_13466,N_12976,N_13142);
or U13467 (N_13467,N_13127,N_12997);
nand U13468 (N_13468,N_12949,N_13118);
nand U13469 (N_13469,N_12977,N_12914);
nor U13470 (N_13470,N_12729,N_12711);
xnor U13471 (N_13471,N_12936,N_12890);
nand U13472 (N_13472,N_12971,N_12825);
and U13473 (N_13473,N_12917,N_12687);
nor U13474 (N_13474,N_12611,N_12636);
and U13475 (N_13475,N_12860,N_12879);
nor U13476 (N_13476,N_12671,N_12758);
nor U13477 (N_13477,N_12942,N_12855);
and U13478 (N_13478,N_12951,N_12609);
xor U13479 (N_13479,N_12852,N_13035);
nor U13480 (N_13480,N_13047,N_12764);
nor U13481 (N_13481,N_12963,N_12761);
nor U13482 (N_13482,N_12785,N_12918);
or U13483 (N_13483,N_12716,N_13165);
xnor U13484 (N_13484,N_12689,N_12935);
nand U13485 (N_13485,N_12752,N_12822);
nor U13486 (N_13486,N_12803,N_12721);
nor U13487 (N_13487,N_12900,N_12775);
and U13488 (N_13488,N_12743,N_13012);
nor U13489 (N_13489,N_12641,N_12760);
or U13490 (N_13490,N_13082,N_12897);
nor U13491 (N_13491,N_12950,N_12750);
and U13492 (N_13492,N_12835,N_13192);
and U13493 (N_13493,N_12804,N_13133);
or U13494 (N_13494,N_12737,N_12984);
nor U13495 (N_13495,N_13143,N_13065);
and U13496 (N_13496,N_12894,N_13190);
and U13497 (N_13497,N_13070,N_13000);
xnor U13498 (N_13498,N_12832,N_12688);
and U13499 (N_13499,N_13140,N_12762);
xor U13500 (N_13500,N_13125,N_13067);
nand U13501 (N_13501,N_12612,N_12928);
nand U13502 (N_13502,N_12745,N_13156);
nand U13503 (N_13503,N_12713,N_13089);
nand U13504 (N_13504,N_12928,N_12822);
or U13505 (N_13505,N_12858,N_12740);
xnor U13506 (N_13506,N_13134,N_12889);
xor U13507 (N_13507,N_12793,N_12760);
nor U13508 (N_13508,N_13142,N_12926);
xnor U13509 (N_13509,N_12695,N_13097);
xor U13510 (N_13510,N_12949,N_13185);
xor U13511 (N_13511,N_12963,N_12923);
nand U13512 (N_13512,N_12762,N_12799);
or U13513 (N_13513,N_12892,N_12916);
nand U13514 (N_13514,N_12905,N_12904);
nand U13515 (N_13515,N_12959,N_12879);
or U13516 (N_13516,N_13169,N_12799);
and U13517 (N_13517,N_12737,N_12787);
nor U13518 (N_13518,N_12901,N_12741);
nor U13519 (N_13519,N_12770,N_12733);
or U13520 (N_13520,N_12787,N_12614);
nor U13521 (N_13521,N_12963,N_13042);
and U13522 (N_13522,N_12715,N_13125);
nand U13523 (N_13523,N_13020,N_12970);
nor U13524 (N_13524,N_12603,N_12704);
xnor U13525 (N_13525,N_12693,N_13011);
nand U13526 (N_13526,N_12679,N_12965);
xor U13527 (N_13527,N_12920,N_12707);
and U13528 (N_13528,N_13034,N_12829);
nand U13529 (N_13529,N_13094,N_12738);
and U13530 (N_13530,N_13099,N_13154);
nand U13531 (N_13531,N_12985,N_13145);
and U13532 (N_13532,N_12859,N_12872);
or U13533 (N_13533,N_13111,N_12896);
or U13534 (N_13534,N_12874,N_12891);
nor U13535 (N_13535,N_13163,N_13191);
nand U13536 (N_13536,N_12982,N_12724);
nand U13537 (N_13537,N_13141,N_12909);
nand U13538 (N_13538,N_13115,N_12767);
nor U13539 (N_13539,N_13002,N_12813);
or U13540 (N_13540,N_13191,N_12915);
xor U13541 (N_13541,N_12975,N_12836);
and U13542 (N_13542,N_13169,N_12792);
xor U13543 (N_13543,N_13059,N_13178);
xnor U13544 (N_13544,N_12923,N_12982);
and U13545 (N_13545,N_12706,N_13182);
or U13546 (N_13546,N_12932,N_12935);
nand U13547 (N_13547,N_12648,N_12791);
or U13548 (N_13548,N_12974,N_12703);
nor U13549 (N_13549,N_12923,N_12616);
nand U13550 (N_13550,N_12733,N_13102);
nor U13551 (N_13551,N_12937,N_12844);
nand U13552 (N_13552,N_13189,N_13127);
and U13553 (N_13553,N_12905,N_12675);
nand U13554 (N_13554,N_12912,N_12881);
nor U13555 (N_13555,N_13022,N_12771);
xor U13556 (N_13556,N_13171,N_12963);
xnor U13557 (N_13557,N_13077,N_12662);
nor U13558 (N_13558,N_12635,N_12870);
nand U13559 (N_13559,N_12876,N_12822);
or U13560 (N_13560,N_12702,N_12664);
or U13561 (N_13561,N_12916,N_13113);
xnor U13562 (N_13562,N_13175,N_12679);
nor U13563 (N_13563,N_13190,N_13046);
or U13564 (N_13564,N_12910,N_12611);
nor U13565 (N_13565,N_12902,N_12719);
nor U13566 (N_13566,N_12915,N_12680);
nand U13567 (N_13567,N_12700,N_12736);
and U13568 (N_13568,N_12872,N_12989);
xor U13569 (N_13569,N_13102,N_12708);
or U13570 (N_13570,N_12875,N_12732);
nor U13571 (N_13571,N_12949,N_12693);
nand U13572 (N_13572,N_13136,N_12660);
nand U13573 (N_13573,N_13191,N_13138);
nor U13574 (N_13574,N_13146,N_12803);
and U13575 (N_13575,N_12600,N_13033);
nand U13576 (N_13576,N_12652,N_12925);
and U13577 (N_13577,N_12629,N_12892);
or U13578 (N_13578,N_12892,N_13006);
or U13579 (N_13579,N_13092,N_13000);
and U13580 (N_13580,N_12955,N_12894);
and U13581 (N_13581,N_13022,N_12674);
or U13582 (N_13582,N_12618,N_12935);
and U13583 (N_13583,N_12893,N_13174);
nand U13584 (N_13584,N_12964,N_13082);
and U13585 (N_13585,N_13120,N_12841);
or U13586 (N_13586,N_13148,N_12666);
nor U13587 (N_13587,N_13095,N_13020);
and U13588 (N_13588,N_13197,N_12898);
and U13589 (N_13589,N_12930,N_12671);
nand U13590 (N_13590,N_13156,N_12886);
xnor U13591 (N_13591,N_12601,N_12873);
nand U13592 (N_13592,N_12601,N_12715);
xor U13593 (N_13593,N_12994,N_12801);
xnor U13594 (N_13594,N_13187,N_12919);
or U13595 (N_13595,N_12646,N_12619);
or U13596 (N_13596,N_12691,N_12923);
and U13597 (N_13597,N_12788,N_13063);
or U13598 (N_13598,N_12974,N_13032);
nand U13599 (N_13599,N_13108,N_13193);
and U13600 (N_13600,N_12663,N_13061);
and U13601 (N_13601,N_12927,N_13116);
nand U13602 (N_13602,N_12703,N_13174);
xnor U13603 (N_13603,N_12936,N_13050);
xor U13604 (N_13604,N_12910,N_12713);
and U13605 (N_13605,N_13124,N_12909);
nand U13606 (N_13606,N_12685,N_12958);
nand U13607 (N_13607,N_12662,N_12942);
nand U13608 (N_13608,N_13008,N_13037);
nand U13609 (N_13609,N_12625,N_12702);
nor U13610 (N_13610,N_13101,N_13174);
nor U13611 (N_13611,N_12946,N_12821);
and U13612 (N_13612,N_13102,N_13120);
nor U13613 (N_13613,N_12980,N_12866);
or U13614 (N_13614,N_13132,N_12823);
nor U13615 (N_13615,N_13023,N_13086);
nor U13616 (N_13616,N_12746,N_12900);
nand U13617 (N_13617,N_12778,N_12917);
nand U13618 (N_13618,N_13018,N_12763);
and U13619 (N_13619,N_12776,N_12698);
and U13620 (N_13620,N_13151,N_13175);
xor U13621 (N_13621,N_13017,N_12860);
xor U13622 (N_13622,N_12793,N_13181);
and U13623 (N_13623,N_12808,N_12813);
xnor U13624 (N_13624,N_12933,N_12758);
nor U13625 (N_13625,N_12645,N_12744);
xnor U13626 (N_13626,N_12674,N_12617);
nor U13627 (N_13627,N_12667,N_13062);
and U13628 (N_13628,N_12669,N_13025);
xnor U13629 (N_13629,N_12720,N_13103);
xor U13630 (N_13630,N_13119,N_12716);
xor U13631 (N_13631,N_12851,N_13098);
xor U13632 (N_13632,N_12786,N_12600);
nand U13633 (N_13633,N_12827,N_13096);
or U13634 (N_13634,N_12678,N_12840);
nand U13635 (N_13635,N_13193,N_12751);
or U13636 (N_13636,N_12674,N_12983);
nand U13637 (N_13637,N_12897,N_12688);
xnor U13638 (N_13638,N_12995,N_13041);
xor U13639 (N_13639,N_13099,N_12603);
nor U13640 (N_13640,N_13130,N_13106);
nor U13641 (N_13641,N_13001,N_12665);
and U13642 (N_13642,N_12838,N_12645);
and U13643 (N_13643,N_13185,N_12944);
or U13644 (N_13644,N_12946,N_13064);
xor U13645 (N_13645,N_12632,N_12977);
nand U13646 (N_13646,N_13045,N_13166);
and U13647 (N_13647,N_13163,N_13027);
nand U13648 (N_13648,N_12906,N_12750);
and U13649 (N_13649,N_12693,N_12674);
xnor U13650 (N_13650,N_12661,N_12955);
xor U13651 (N_13651,N_12873,N_13010);
xor U13652 (N_13652,N_12688,N_12829);
xor U13653 (N_13653,N_12856,N_12781);
or U13654 (N_13654,N_12771,N_13060);
and U13655 (N_13655,N_12795,N_12765);
nor U13656 (N_13656,N_12958,N_12676);
nand U13657 (N_13657,N_12976,N_13187);
or U13658 (N_13658,N_12843,N_13125);
xor U13659 (N_13659,N_13149,N_12718);
and U13660 (N_13660,N_12694,N_13197);
xor U13661 (N_13661,N_13005,N_12647);
and U13662 (N_13662,N_12605,N_12722);
xnor U13663 (N_13663,N_12924,N_12618);
nand U13664 (N_13664,N_13047,N_13162);
and U13665 (N_13665,N_13125,N_12676);
xor U13666 (N_13666,N_12710,N_13019);
or U13667 (N_13667,N_12762,N_12989);
nand U13668 (N_13668,N_13020,N_13171);
and U13669 (N_13669,N_12851,N_12646);
nand U13670 (N_13670,N_12908,N_12873);
and U13671 (N_13671,N_12885,N_12801);
and U13672 (N_13672,N_13045,N_13169);
nor U13673 (N_13673,N_13074,N_12747);
and U13674 (N_13674,N_12927,N_12728);
or U13675 (N_13675,N_13051,N_12925);
nor U13676 (N_13676,N_13156,N_12919);
nor U13677 (N_13677,N_13091,N_13160);
or U13678 (N_13678,N_12775,N_12795);
xnor U13679 (N_13679,N_12676,N_12888);
and U13680 (N_13680,N_13051,N_12809);
nand U13681 (N_13681,N_12976,N_13084);
nor U13682 (N_13682,N_12632,N_12746);
and U13683 (N_13683,N_12968,N_12638);
nor U13684 (N_13684,N_12950,N_12986);
and U13685 (N_13685,N_12648,N_12674);
nor U13686 (N_13686,N_13003,N_13195);
nand U13687 (N_13687,N_13041,N_12794);
xnor U13688 (N_13688,N_12803,N_13109);
xor U13689 (N_13689,N_13026,N_12667);
or U13690 (N_13690,N_13151,N_13120);
xnor U13691 (N_13691,N_13066,N_13003);
nand U13692 (N_13692,N_12822,N_12832);
nand U13693 (N_13693,N_12739,N_13130);
nand U13694 (N_13694,N_13050,N_13046);
nor U13695 (N_13695,N_12825,N_12790);
and U13696 (N_13696,N_13189,N_13164);
nand U13697 (N_13697,N_12608,N_13095);
xnor U13698 (N_13698,N_12653,N_12866);
or U13699 (N_13699,N_13193,N_12921);
xnor U13700 (N_13700,N_12886,N_12771);
or U13701 (N_13701,N_13062,N_12937);
or U13702 (N_13702,N_12863,N_12741);
nor U13703 (N_13703,N_12813,N_12723);
and U13704 (N_13704,N_12974,N_12928);
and U13705 (N_13705,N_13152,N_12831);
nor U13706 (N_13706,N_12903,N_12920);
xnor U13707 (N_13707,N_12720,N_12677);
nand U13708 (N_13708,N_12852,N_12764);
or U13709 (N_13709,N_13071,N_13056);
nand U13710 (N_13710,N_12927,N_12925);
and U13711 (N_13711,N_12664,N_12628);
and U13712 (N_13712,N_12957,N_12702);
nor U13713 (N_13713,N_12866,N_13102);
and U13714 (N_13714,N_12948,N_12801);
xor U13715 (N_13715,N_12762,N_12601);
xnor U13716 (N_13716,N_12875,N_13003);
or U13717 (N_13717,N_12688,N_13067);
and U13718 (N_13718,N_12668,N_12712);
and U13719 (N_13719,N_12615,N_12712);
or U13720 (N_13720,N_13122,N_13069);
and U13721 (N_13721,N_12663,N_12639);
or U13722 (N_13722,N_12837,N_12970);
nor U13723 (N_13723,N_12766,N_12945);
nand U13724 (N_13724,N_12890,N_12656);
xor U13725 (N_13725,N_13054,N_12652);
nor U13726 (N_13726,N_12732,N_12817);
nand U13727 (N_13727,N_12768,N_12604);
xnor U13728 (N_13728,N_12894,N_13028);
nor U13729 (N_13729,N_12744,N_13179);
nand U13730 (N_13730,N_12737,N_12724);
or U13731 (N_13731,N_12731,N_13034);
or U13732 (N_13732,N_12870,N_12811);
nor U13733 (N_13733,N_13087,N_12843);
nand U13734 (N_13734,N_12848,N_12612);
and U13735 (N_13735,N_12637,N_12762);
nor U13736 (N_13736,N_12986,N_12717);
and U13737 (N_13737,N_12700,N_12874);
or U13738 (N_13738,N_13092,N_12903);
nand U13739 (N_13739,N_12666,N_12804);
nor U13740 (N_13740,N_12770,N_12686);
or U13741 (N_13741,N_12805,N_13032);
xor U13742 (N_13742,N_12955,N_13015);
nand U13743 (N_13743,N_12772,N_12940);
or U13744 (N_13744,N_13031,N_12712);
nand U13745 (N_13745,N_12713,N_12782);
or U13746 (N_13746,N_13061,N_12852);
and U13747 (N_13747,N_12706,N_13027);
xnor U13748 (N_13748,N_12704,N_12849);
and U13749 (N_13749,N_12682,N_12602);
xnor U13750 (N_13750,N_13094,N_12633);
nand U13751 (N_13751,N_13048,N_13027);
or U13752 (N_13752,N_12758,N_12891);
xnor U13753 (N_13753,N_12938,N_12911);
xnor U13754 (N_13754,N_12671,N_13027);
xnor U13755 (N_13755,N_12613,N_12665);
nand U13756 (N_13756,N_13115,N_12674);
xor U13757 (N_13757,N_12815,N_13085);
or U13758 (N_13758,N_12616,N_12899);
or U13759 (N_13759,N_13058,N_12698);
nand U13760 (N_13760,N_13065,N_12813);
nor U13761 (N_13761,N_12649,N_13066);
or U13762 (N_13762,N_13020,N_12973);
or U13763 (N_13763,N_12679,N_13099);
and U13764 (N_13764,N_12921,N_12763);
nor U13765 (N_13765,N_12792,N_13042);
xnor U13766 (N_13766,N_12980,N_13101);
xor U13767 (N_13767,N_12895,N_12990);
nor U13768 (N_13768,N_13185,N_12990);
nor U13769 (N_13769,N_12637,N_12952);
nand U13770 (N_13770,N_12859,N_12937);
and U13771 (N_13771,N_13035,N_12867);
nand U13772 (N_13772,N_12775,N_12783);
and U13773 (N_13773,N_13075,N_12793);
nand U13774 (N_13774,N_12774,N_12924);
nand U13775 (N_13775,N_12973,N_13153);
nand U13776 (N_13776,N_12955,N_12730);
and U13777 (N_13777,N_12945,N_13103);
nand U13778 (N_13778,N_12766,N_12999);
nor U13779 (N_13779,N_13063,N_13165);
or U13780 (N_13780,N_12727,N_12990);
nor U13781 (N_13781,N_12679,N_12896);
nand U13782 (N_13782,N_12823,N_12853);
and U13783 (N_13783,N_12854,N_12628);
nand U13784 (N_13784,N_13016,N_13020);
nor U13785 (N_13785,N_13021,N_12736);
and U13786 (N_13786,N_12626,N_12668);
nor U13787 (N_13787,N_12772,N_12626);
nor U13788 (N_13788,N_12793,N_13128);
xor U13789 (N_13789,N_13183,N_12753);
or U13790 (N_13790,N_12782,N_13008);
nand U13791 (N_13791,N_12695,N_13128);
and U13792 (N_13792,N_12740,N_12952);
or U13793 (N_13793,N_12819,N_12814);
nor U13794 (N_13794,N_12829,N_12888);
nor U13795 (N_13795,N_12643,N_12952);
nor U13796 (N_13796,N_12874,N_13018);
or U13797 (N_13797,N_12648,N_12827);
nor U13798 (N_13798,N_12600,N_12735);
nor U13799 (N_13799,N_12918,N_12812);
nand U13800 (N_13800,N_13265,N_13415);
xor U13801 (N_13801,N_13781,N_13399);
or U13802 (N_13802,N_13201,N_13290);
or U13803 (N_13803,N_13683,N_13378);
or U13804 (N_13804,N_13605,N_13280);
nand U13805 (N_13805,N_13461,N_13629);
or U13806 (N_13806,N_13436,N_13516);
xnor U13807 (N_13807,N_13510,N_13546);
nand U13808 (N_13808,N_13653,N_13323);
or U13809 (N_13809,N_13440,N_13754);
xor U13810 (N_13810,N_13585,N_13608);
and U13811 (N_13811,N_13661,N_13619);
nor U13812 (N_13812,N_13594,N_13662);
and U13813 (N_13813,N_13581,N_13272);
nand U13814 (N_13814,N_13237,N_13634);
and U13815 (N_13815,N_13344,N_13509);
and U13816 (N_13816,N_13479,N_13632);
and U13817 (N_13817,N_13268,N_13222);
and U13818 (N_13818,N_13622,N_13665);
and U13819 (N_13819,N_13286,N_13716);
xor U13820 (N_13820,N_13587,N_13664);
and U13821 (N_13821,N_13707,N_13687);
xor U13822 (N_13822,N_13756,N_13238);
xnor U13823 (N_13823,N_13469,N_13447);
and U13824 (N_13824,N_13251,N_13441);
and U13825 (N_13825,N_13458,N_13519);
xor U13826 (N_13826,N_13226,N_13274);
nand U13827 (N_13827,N_13410,N_13452);
nand U13828 (N_13828,N_13429,N_13604);
nand U13829 (N_13829,N_13395,N_13554);
or U13830 (N_13830,N_13545,N_13439);
nand U13831 (N_13831,N_13285,N_13695);
xnor U13832 (N_13832,N_13721,N_13644);
and U13833 (N_13833,N_13468,N_13224);
nor U13834 (N_13834,N_13732,N_13531);
nor U13835 (N_13835,N_13267,N_13232);
nand U13836 (N_13836,N_13673,N_13544);
and U13837 (N_13837,N_13621,N_13693);
and U13838 (N_13838,N_13351,N_13291);
xor U13839 (N_13839,N_13462,N_13618);
nor U13840 (N_13840,N_13787,N_13580);
or U13841 (N_13841,N_13365,N_13339);
and U13842 (N_13842,N_13329,N_13616);
and U13843 (N_13843,N_13748,N_13557);
nand U13844 (N_13844,N_13211,N_13537);
or U13845 (N_13845,N_13586,N_13614);
nand U13846 (N_13846,N_13451,N_13243);
nand U13847 (N_13847,N_13353,N_13369);
nand U13848 (N_13848,N_13709,N_13242);
or U13849 (N_13849,N_13637,N_13487);
and U13850 (N_13850,N_13514,N_13476);
nand U13851 (N_13851,N_13209,N_13527);
nor U13852 (N_13852,N_13720,N_13633);
nand U13853 (N_13853,N_13488,N_13692);
nand U13854 (N_13854,N_13655,N_13314);
or U13855 (N_13855,N_13743,N_13795);
and U13856 (N_13856,N_13266,N_13646);
and U13857 (N_13857,N_13538,N_13437);
or U13858 (N_13858,N_13791,N_13259);
and U13859 (N_13859,N_13292,N_13304);
or U13860 (N_13860,N_13698,N_13471);
nor U13861 (N_13861,N_13563,N_13595);
and U13862 (N_13862,N_13725,N_13249);
nor U13863 (N_13863,N_13303,N_13680);
and U13864 (N_13864,N_13635,N_13525);
or U13865 (N_13865,N_13566,N_13689);
or U13866 (N_13866,N_13230,N_13744);
and U13867 (N_13867,N_13783,N_13567);
xor U13868 (N_13868,N_13326,N_13796);
nor U13869 (N_13869,N_13533,N_13360);
xnor U13870 (N_13870,N_13349,N_13278);
nor U13871 (N_13871,N_13387,N_13416);
and U13872 (N_13872,N_13247,N_13651);
nor U13873 (N_13873,N_13374,N_13388);
and U13874 (N_13874,N_13660,N_13785);
nand U13875 (N_13875,N_13738,N_13472);
nor U13876 (N_13876,N_13240,N_13542);
xnor U13877 (N_13877,N_13375,N_13790);
and U13878 (N_13878,N_13475,N_13385);
xor U13879 (N_13879,N_13455,N_13253);
or U13880 (N_13880,N_13504,N_13681);
nand U13881 (N_13881,N_13438,N_13256);
xor U13882 (N_13882,N_13766,N_13562);
and U13883 (N_13883,N_13317,N_13464);
xnor U13884 (N_13884,N_13245,N_13667);
and U13885 (N_13885,N_13448,N_13298);
and U13886 (N_13886,N_13467,N_13702);
nand U13887 (N_13887,N_13383,N_13508);
xor U13888 (N_13888,N_13481,N_13578);
xor U13889 (N_13889,N_13221,N_13381);
and U13890 (N_13890,N_13423,N_13271);
or U13891 (N_13891,N_13417,N_13645);
or U13892 (N_13892,N_13491,N_13737);
and U13893 (N_13893,N_13677,N_13778);
or U13894 (N_13894,N_13214,N_13348);
and U13895 (N_13895,N_13712,N_13282);
nand U13896 (N_13896,N_13564,N_13493);
nor U13897 (N_13897,N_13302,N_13456);
or U13898 (N_13898,N_13362,N_13498);
nor U13899 (N_13899,N_13729,N_13406);
and U13900 (N_13900,N_13411,N_13218);
or U13901 (N_13901,N_13305,N_13257);
nor U13902 (N_13902,N_13733,N_13370);
nand U13903 (N_13903,N_13705,N_13799);
nand U13904 (N_13904,N_13200,N_13691);
nor U13905 (N_13905,N_13283,N_13270);
nand U13906 (N_13906,N_13293,N_13570);
or U13907 (N_13907,N_13718,N_13773);
nand U13908 (N_13908,N_13223,N_13255);
xnor U13909 (N_13909,N_13706,N_13246);
nor U13910 (N_13910,N_13552,N_13534);
nand U13911 (N_13911,N_13335,N_13625);
or U13912 (N_13912,N_13584,N_13768);
or U13913 (N_13913,N_13669,N_13688);
nand U13914 (N_13914,N_13524,N_13396);
nor U13915 (N_13915,N_13483,N_13239);
nand U13916 (N_13916,N_13289,N_13306);
xnor U13917 (N_13917,N_13575,N_13338);
xnor U13918 (N_13918,N_13658,N_13607);
nand U13919 (N_13919,N_13728,N_13319);
nand U13920 (N_13920,N_13643,N_13572);
or U13921 (N_13921,N_13789,N_13397);
xnor U13922 (N_13922,N_13609,N_13758);
nand U13923 (N_13923,N_13354,N_13394);
and U13924 (N_13924,N_13241,N_13296);
nor U13925 (N_13925,N_13358,N_13672);
nand U13926 (N_13926,N_13424,N_13393);
nand U13927 (N_13927,N_13315,N_13433);
nand U13928 (N_13928,N_13412,N_13343);
or U13929 (N_13929,N_13261,N_13526);
and U13930 (N_13930,N_13231,N_13495);
and U13931 (N_13931,N_13421,N_13589);
or U13932 (N_13932,N_13250,N_13719);
or U13933 (N_13933,N_13565,N_13699);
nor U13934 (N_13934,N_13392,N_13690);
or U13935 (N_13935,N_13505,N_13228);
or U13936 (N_13936,N_13640,N_13435);
xnor U13937 (N_13937,N_13742,N_13460);
and U13938 (N_13938,N_13626,N_13675);
and U13939 (N_13939,N_13263,N_13597);
or U13940 (N_13940,N_13484,N_13599);
nor U13941 (N_13941,N_13694,N_13715);
xnor U13942 (N_13942,N_13213,N_13372);
nor U13943 (N_13943,N_13316,N_13615);
xnor U13944 (N_13944,N_13420,N_13308);
or U13945 (N_13945,N_13312,N_13398);
and U13946 (N_13946,N_13610,N_13409);
nand U13947 (N_13947,N_13761,N_13666);
or U13948 (N_13948,N_13294,N_13523);
nand U13949 (N_13949,N_13300,N_13219);
xnor U13950 (N_13950,N_13755,N_13624);
or U13951 (N_13951,N_13485,N_13321);
xor U13952 (N_13952,N_13337,N_13442);
xnor U13953 (N_13953,N_13740,N_13384);
nand U13954 (N_13954,N_13422,N_13331);
nor U13955 (N_13955,N_13671,N_13408);
or U13956 (N_13956,N_13553,N_13639);
and U13957 (N_13957,N_13212,N_13361);
nand U13958 (N_13958,N_13547,N_13473);
xor U13959 (N_13959,N_13678,N_13356);
nor U13960 (N_13960,N_13390,N_13714);
or U13961 (N_13961,N_13638,N_13497);
nand U13962 (N_13962,N_13430,N_13735);
or U13963 (N_13963,N_13753,N_13465);
xor U13964 (N_13964,N_13466,N_13613);
and U13965 (N_13965,N_13401,N_13577);
or U13966 (N_13966,N_13457,N_13543);
nand U13967 (N_13967,N_13764,N_13478);
or U13968 (N_13968,N_13264,N_13551);
nand U13969 (N_13969,N_13324,N_13446);
nand U13970 (N_13970,N_13382,N_13431);
xor U13971 (N_13971,N_13407,N_13373);
xnor U13972 (N_13972,N_13490,N_13459);
xor U13973 (N_13973,N_13269,N_13334);
nand U13974 (N_13974,N_13606,N_13262);
and U13975 (N_13975,N_13454,N_13359);
or U13976 (N_13976,N_13751,N_13696);
xnor U13977 (N_13977,N_13797,N_13434);
xor U13978 (N_13978,N_13571,N_13593);
nand U13979 (N_13979,N_13203,N_13333);
xor U13980 (N_13980,N_13512,N_13647);
xnor U13981 (N_13981,N_13277,N_13731);
or U13982 (N_13982,N_13309,N_13528);
nor U13983 (N_13983,N_13413,N_13463);
nor U13984 (N_13984,N_13276,N_13786);
and U13985 (N_13985,N_13765,N_13336);
nand U13986 (N_13986,N_13404,N_13225);
and U13987 (N_13987,N_13367,N_13656);
and U13988 (N_13988,N_13573,N_13518);
or U13989 (N_13989,N_13503,N_13535);
nand U13990 (N_13990,N_13313,N_13601);
nor U13991 (N_13991,N_13379,N_13650);
nand U13992 (N_13992,N_13657,N_13684);
xnor U13993 (N_13993,N_13583,N_13494);
and U13994 (N_13994,N_13569,N_13363);
or U13995 (N_13995,N_13496,N_13701);
or U13996 (N_13996,N_13548,N_13414);
nand U13997 (N_13997,N_13474,N_13549);
xor U13998 (N_13998,N_13244,N_13749);
or U13999 (N_13999,N_13784,N_13704);
or U14000 (N_14000,N_13780,N_13341);
nor U14001 (N_14001,N_13260,N_13206);
or U14002 (N_14002,N_13450,N_13652);
nand U14003 (N_14003,N_13679,N_13654);
and U14004 (N_14004,N_13521,N_13760);
or U14005 (N_14005,N_13210,N_13301);
nand U14006 (N_14006,N_13529,N_13402);
or U14007 (N_14007,N_13770,N_13710);
xor U14008 (N_14008,N_13376,N_13555);
or U14009 (N_14009,N_13628,N_13642);
xor U14010 (N_14010,N_13330,N_13470);
nor U14011 (N_14011,N_13350,N_13730);
nand U14012 (N_14012,N_13582,N_13310);
nand U14013 (N_14013,N_13697,N_13328);
nand U14014 (N_14014,N_13425,N_13327);
xnor U14015 (N_14015,N_13480,N_13346);
nor U14016 (N_14016,N_13332,N_13631);
nor U14017 (N_14017,N_13234,N_13596);
nand U14018 (N_14018,N_13522,N_13746);
nand U14019 (N_14019,N_13603,N_13641);
and U14020 (N_14020,N_13774,N_13258);
and U14021 (N_14021,N_13530,N_13726);
or U14022 (N_14022,N_13769,N_13443);
nor U14023 (N_14023,N_13736,N_13284);
xor U14024 (N_14024,N_13297,N_13419);
or U14025 (N_14025,N_13205,N_13745);
nor U14026 (N_14026,N_13287,N_13352);
xnor U14027 (N_14027,N_13482,N_13727);
nor U14028 (N_14028,N_13275,N_13506);
or U14029 (N_14029,N_13762,N_13320);
xnor U14030 (N_14030,N_13368,N_13739);
or U14031 (N_14031,N_13747,N_13576);
xnor U14032 (N_14032,N_13636,N_13711);
xor U14033 (N_14033,N_13611,N_13602);
xnor U14034 (N_14034,N_13322,N_13630);
nand U14035 (N_14035,N_13685,N_13325);
xor U14036 (N_14036,N_13788,N_13345);
nor U14037 (N_14037,N_13511,N_13612);
or U14038 (N_14038,N_13617,N_13500);
xnor U14039 (N_14039,N_13713,N_13340);
nor U14040 (N_14040,N_13386,N_13590);
nand U14041 (N_14041,N_13568,N_13204);
xor U14042 (N_14042,N_13486,N_13389);
nand U14043 (N_14043,N_13579,N_13515);
nand U14044 (N_14044,N_13295,N_13380);
and U14045 (N_14045,N_13777,N_13600);
nor U14046 (N_14046,N_13507,N_13347);
xor U14047 (N_14047,N_13377,N_13536);
xnor U14048 (N_14048,N_13792,N_13371);
and U14049 (N_14049,N_13532,N_13752);
and U14050 (N_14050,N_13556,N_13794);
xor U14051 (N_14051,N_13489,N_13772);
nand U14052 (N_14052,N_13355,N_13559);
xor U14053 (N_14053,N_13307,N_13288);
nand U14054 (N_14054,N_13432,N_13703);
xnor U14055 (N_14055,N_13750,N_13428);
nor U14056 (N_14056,N_13229,N_13623);
xnor U14057 (N_14057,N_13798,N_13318);
or U14058 (N_14058,N_13252,N_13235);
xnor U14059 (N_14059,N_13722,N_13560);
or U14060 (N_14060,N_13620,N_13273);
nand U14061 (N_14061,N_13757,N_13686);
and U14062 (N_14062,N_13453,N_13311);
nor U14063 (N_14063,N_13591,N_13492);
nand U14064 (N_14064,N_13682,N_13364);
or U14065 (N_14065,N_13391,N_13649);
nor U14066 (N_14066,N_13299,N_13734);
nor U14067 (N_14067,N_13202,N_13763);
nor U14068 (N_14068,N_13499,N_13207);
nor U14069 (N_14069,N_13708,N_13771);
xor U14070 (N_14070,N_13598,N_13659);
and U14071 (N_14071,N_13405,N_13668);
and U14072 (N_14072,N_13775,N_13588);
xor U14073 (N_14073,N_13342,N_13220);
nor U14074 (N_14074,N_13502,N_13627);
xnor U14075 (N_14075,N_13208,N_13724);
or U14076 (N_14076,N_13444,N_13670);
and U14077 (N_14077,N_13254,N_13663);
and U14078 (N_14078,N_13782,N_13366);
nand U14079 (N_14079,N_13248,N_13592);
nor U14080 (N_14080,N_13648,N_13550);
xor U14081 (N_14081,N_13561,N_13574);
and U14082 (N_14082,N_13674,N_13477);
and U14083 (N_14083,N_13513,N_13400);
xnor U14084 (N_14084,N_13449,N_13779);
xor U14085 (N_14085,N_13520,N_13558);
or U14086 (N_14086,N_13767,N_13776);
or U14087 (N_14087,N_13281,N_13418);
or U14088 (N_14088,N_13793,N_13426);
or U14089 (N_14089,N_13445,N_13741);
nand U14090 (N_14090,N_13236,N_13403);
or U14091 (N_14091,N_13700,N_13723);
nor U14092 (N_14092,N_13759,N_13233);
and U14093 (N_14093,N_13427,N_13541);
and U14094 (N_14094,N_13517,N_13215);
nand U14095 (N_14095,N_13540,N_13676);
nor U14096 (N_14096,N_13279,N_13217);
nand U14097 (N_14097,N_13539,N_13357);
and U14098 (N_14098,N_13216,N_13501);
nor U14099 (N_14099,N_13717,N_13227);
nand U14100 (N_14100,N_13767,N_13256);
and U14101 (N_14101,N_13452,N_13762);
nand U14102 (N_14102,N_13410,N_13440);
nand U14103 (N_14103,N_13305,N_13721);
nand U14104 (N_14104,N_13495,N_13715);
and U14105 (N_14105,N_13398,N_13784);
nor U14106 (N_14106,N_13754,N_13334);
and U14107 (N_14107,N_13731,N_13756);
and U14108 (N_14108,N_13701,N_13380);
xor U14109 (N_14109,N_13337,N_13517);
and U14110 (N_14110,N_13799,N_13258);
nor U14111 (N_14111,N_13405,N_13714);
nand U14112 (N_14112,N_13602,N_13337);
and U14113 (N_14113,N_13768,N_13268);
or U14114 (N_14114,N_13607,N_13790);
or U14115 (N_14115,N_13737,N_13681);
or U14116 (N_14116,N_13413,N_13578);
nand U14117 (N_14117,N_13282,N_13750);
nor U14118 (N_14118,N_13284,N_13613);
nor U14119 (N_14119,N_13454,N_13367);
nand U14120 (N_14120,N_13524,N_13446);
nand U14121 (N_14121,N_13637,N_13708);
or U14122 (N_14122,N_13723,N_13346);
and U14123 (N_14123,N_13426,N_13630);
nor U14124 (N_14124,N_13650,N_13320);
and U14125 (N_14125,N_13468,N_13465);
xnor U14126 (N_14126,N_13566,N_13437);
or U14127 (N_14127,N_13630,N_13627);
nand U14128 (N_14128,N_13340,N_13776);
xnor U14129 (N_14129,N_13636,N_13486);
and U14130 (N_14130,N_13746,N_13262);
nand U14131 (N_14131,N_13692,N_13602);
nand U14132 (N_14132,N_13505,N_13707);
xnor U14133 (N_14133,N_13616,N_13314);
or U14134 (N_14134,N_13729,N_13237);
nor U14135 (N_14135,N_13773,N_13736);
xnor U14136 (N_14136,N_13389,N_13350);
and U14137 (N_14137,N_13593,N_13471);
nor U14138 (N_14138,N_13363,N_13731);
and U14139 (N_14139,N_13583,N_13496);
and U14140 (N_14140,N_13629,N_13265);
nor U14141 (N_14141,N_13204,N_13291);
or U14142 (N_14142,N_13253,N_13415);
or U14143 (N_14143,N_13239,N_13450);
or U14144 (N_14144,N_13281,N_13391);
or U14145 (N_14145,N_13439,N_13626);
nand U14146 (N_14146,N_13253,N_13631);
and U14147 (N_14147,N_13279,N_13660);
xor U14148 (N_14148,N_13270,N_13602);
xor U14149 (N_14149,N_13641,N_13767);
or U14150 (N_14150,N_13350,N_13406);
nor U14151 (N_14151,N_13689,N_13626);
nand U14152 (N_14152,N_13372,N_13326);
or U14153 (N_14153,N_13209,N_13295);
xnor U14154 (N_14154,N_13774,N_13655);
nor U14155 (N_14155,N_13272,N_13382);
and U14156 (N_14156,N_13685,N_13623);
nor U14157 (N_14157,N_13606,N_13322);
nand U14158 (N_14158,N_13581,N_13238);
nor U14159 (N_14159,N_13402,N_13661);
or U14160 (N_14160,N_13421,N_13392);
and U14161 (N_14161,N_13316,N_13768);
or U14162 (N_14162,N_13295,N_13678);
and U14163 (N_14163,N_13386,N_13300);
xor U14164 (N_14164,N_13351,N_13372);
or U14165 (N_14165,N_13240,N_13726);
or U14166 (N_14166,N_13256,N_13481);
xor U14167 (N_14167,N_13611,N_13693);
and U14168 (N_14168,N_13469,N_13776);
and U14169 (N_14169,N_13581,N_13322);
xnor U14170 (N_14170,N_13547,N_13251);
or U14171 (N_14171,N_13657,N_13318);
nand U14172 (N_14172,N_13415,N_13292);
nand U14173 (N_14173,N_13497,N_13601);
nand U14174 (N_14174,N_13786,N_13652);
nor U14175 (N_14175,N_13479,N_13691);
and U14176 (N_14176,N_13616,N_13639);
and U14177 (N_14177,N_13729,N_13217);
xnor U14178 (N_14178,N_13344,N_13633);
xnor U14179 (N_14179,N_13316,N_13743);
nand U14180 (N_14180,N_13327,N_13613);
nand U14181 (N_14181,N_13455,N_13646);
xor U14182 (N_14182,N_13494,N_13783);
nand U14183 (N_14183,N_13297,N_13500);
xor U14184 (N_14184,N_13492,N_13325);
xnor U14185 (N_14185,N_13595,N_13585);
or U14186 (N_14186,N_13595,N_13472);
xnor U14187 (N_14187,N_13203,N_13270);
nor U14188 (N_14188,N_13247,N_13266);
nor U14189 (N_14189,N_13403,N_13440);
nand U14190 (N_14190,N_13295,N_13623);
nand U14191 (N_14191,N_13298,N_13562);
or U14192 (N_14192,N_13609,N_13698);
or U14193 (N_14193,N_13738,N_13575);
xnor U14194 (N_14194,N_13536,N_13202);
nand U14195 (N_14195,N_13755,N_13203);
or U14196 (N_14196,N_13211,N_13246);
and U14197 (N_14197,N_13508,N_13407);
xor U14198 (N_14198,N_13265,N_13518);
nand U14199 (N_14199,N_13587,N_13676);
xor U14200 (N_14200,N_13556,N_13510);
nand U14201 (N_14201,N_13686,N_13445);
and U14202 (N_14202,N_13361,N_13752);
xnor U14203 (N_14203,N_13690,N_13361);
xor U14204 (N_14204,N_13292,N_13545);
xor U14205 (N_14205,N_13593,N_13317);
and U14206 (N_14206,N_13689,N_13359);
and U14207 (N_14207,N_13620,N_13789);
nand U14208 (N_14208,N_13269,N_13457);
xor U14209 (N_14209,N_13386,N_13299);
nor U14210 (N_14210,N_13282,N_13509);
or U14211 (N_14211,N_13307,N_13620);
nand U14212 (N_14212,N_13713,N_13448);
and U14213 (N_14213,N_13469,N_13772);
xnor U14214 (N_14214,N_13266,N_13407);
xor U14215 (N_14215,N_13568,N_13678);
or U14216 (N_14216,N_13384,N_13447);
or U14217 (N_14217,N_13615,N_13763);
nand U14218 (N_14218,N_13416,N_13592);
nor U14219 (N_14219,N_13308,N_13389);
xor U14220 (N_14220,N_13373,N_13776);
nand U14221 (N_14221,N_13210,N_13731);
nand U14222 (N_14222,N_13370,N_13346);
or U14223 (N_14223,N_13690,N_13572);
or U14224 (N_14224,N_13493,N_13788);
xor U14225 (N_14225,N_13237,N_13334);
nand U14226 (N_14226,N_13753,N_13388);
or U14227 (N_14227,N_13237,N_13671);
and U14228 (N_14228,N_13312,N_13706);
xnor U14229 (N_14229,N_13739,N_13444);
nor U14230 (N_14230,N_13627,N_13308);
xnor U14231 (N_14231,N_13324,N_13397);
or U14232 (N_14232,N_13282,N_13363);
and U14233 (N_14233,N_13540,N_13581);
nand U14234 (N_14234,N_13469,N_13639);
xnor U14235 (N_14235,N_13435,N_13527);
or U14236 (N_14236,N_13559,N_13716);
nor U14237 (N_14237,N_13336,N_13578);
or U14238 (N_14238,N_13702,N_13667);
xor U14239 (N_14239,N_13610,N_13331);
or U14240 (N_14240,N_13596,N_13558);
xnor U14241 (N_14241,N_13479,N_13248);
and U14242 (N_14242,N_13644,N_13275);
nor U14243 (N_14243,N_13524,N_13710);
nand U14244 (N_14244,N_13618,N_13572);
and U14245 (N_14245,N_13647,N_13503);
xor U14246 (N_14246,N_13288,N_13729);
or U14247 (N_14247,N_13241,N_13346);
nand U14248 (N_14248,N_13419,N_13495);
or U14249 (N_14249,N_13454,N_13220);
or U14250 (N_14250,N_13531,N_13685);
or U14251 (N_14251,N_13297,N_13713);
and U14252 (N_14252,N_13280,N_13272);
and U14253 (N_14253,N_13709,N_13347);
nand U14254 (N_14254,N_13468,N_13294);
or U14255 (N_14255,N_13798,N_13200);
xor U14256 (N_14256,N_13553,N_13786);
and U14257 (N_14257,N_13397,N_13225);
or U14258 (N_14258,N_13738,N_13268);
or U14259 (N_14259,N_13326,N_13712);
nor U14260 (N_14260,N_13510,N_13382);
and U14261 (N_14261,N_13671,N_13707);
xor U14262 (N_14262,N_13594,N_13412);
xnor U14263 (N_14263,N_13291,N_13394);
or U14264 (N_14264,N_13469,N_13320);
or U14265 (N_14265,N_13475,N_13255);
xnor U14266 (N_14266,N_13489,N_13249);
and U14267 (N_14267,N_13496,N_13350);
nor U14268 (N_14268,N_13214,N_13503);
or U14269 (N_14269,N_13743,N_13224);
xor U14270 (N_14270,N_13208,N_13757);
nor U14271 (N_14271,N_13740,N_13253);
and U14272 (N_14272,N_13551,N_13700);
nor U14273 (N_14273,N_13338,N_13451);
xor U14274 (N_14274,N_13522,N_13765);
nand U14275 (N_14275,N_13215,N_13664);
or U14276 (N_14276,N_13459,N_13533);
xor U14277 (N_14277,N_13308,N_13719);
or U14278 (N_14278,N_13762,N_13201);
or U14279 (N_14279,N_13720,N_13304);
xnor U14280 (N_14280,N_13530,N_13550);
or U14281 (N_14281,N_13241,N_13739);
nor U14282 (N_14282,N_13569,N_13762);
xnor U14283 (N_14283,N_13413,N_13454);
nand U14284 (N_14284,N_13695,N_13551);
nor U14285 (N_14285,N_13691,N_13776);
xnor U14286 (N_14286,N_13529,N_13278);
nor U14287 (N_14287,N_13357,N_13391);
or U14288 (N_14288,N_13372,N_13266);
or U14289 (N_14289,N_13660,N_13411);
or U14290 (N_14290,N_13310,N_13711);
and U14291 (N_14291,N_13581,N_13398);
nand U14292 (N_14292,N_13277,N_13477);
and U14293 (N_14293,N_13611,N_13689);
nor U14294 (N_14294,N_13673,N_13698);
nor U14295 (N_14295,N_13578,N_13700);
and U14296 (N_14296,N_13558,N_13234);
nor U14297 (N_14297,N_13458,N_13497);
nor U14298 (N_14298,N_13409,N_13298);
nor U14299 (N_14299,N_13362,N_13674);
and U14300 (N_14300,N_13403,N_13653);
nand U14301 (N_14301,N_13561,N_13339);
nand U14302 (N_14302,N_13374,N_13587);
and U14303 (N_14303,N_13669,N_13397);
nor U14304 (N_14304,N_13491,N_13547);
or U14305 (N_14305,N_13558,N_13522);
or U14306 (N_14306,N_13382,N_13700);
and U14307 (N_14307,N_13494,N_13798);
or U14308 (N_14308,N_13532,N_13270);
xor U14309 (N_14309,N_13736,N_13517);
and U14310 (N_14310,N_13649,N_13576);
nand U14311 (N_14311,N_13544,N_13768);
nand U14312 (N_14312,N_13614,N_13440);
nor U14313 (N_14313,N_13555,N_13238);
nand U14314 (N_14314,N_13714,N_13762);
and U14315 (N_14315,N_13782,N_13572);
nor U14316 (N_14316,N_13573,N_13351);
or U14317 (N_14317,N_13359,N_13371);
nand U14318 (N_14318,N_13215,N_13290);
nor U14319 (N_14319,N_13623,N_13699);
nor U14320 (N_14320,N_13221,N_13753);
xor U14321 (N_14321,N_13729,N_13493);
nand U14322 (N_14322,N_13702,N_13241);
nand U14323 (N_14323,N_13415,N_13781);
or U14324 (N_14324,N_13256,N_13335);
xnor U14325 (N_14325,N_13552,N_13330);
nand U14326 (N_14326,N_13370,N_13562);
xor U14327 (N_14327,N_13761,N_13646);
and U14328 (N_14328,N_13687,N_13648);
nor U14329 (N_14329,N_13403,N_13390);
xor U14330 (N_14330,N_13678,N_13770);
nor U14331 (N_14331,N_13684,N_13735);
nand U14332 (N_14332,N_13799,N_13397);
and U14333 (N_14333,N_13672,N_13281);
and U14334 (N_14334,N_13564,N_13366);
nand U14335 (N_14335,N_13366,N_13287);
nor U14336 (N_14336,N_13559,N_13262);
nor U14337 (N_14337,N_13620,N_13418);
nand U14338 (N_14338,N_13331,N_13712);
nand U14339 (N_14339,N_13764,N_13438);
xor U14340 (N_14340,N_13737,N_13407);
and U14341 (N_14341,N_13449,N_13766);
nor U14342 (N_14342,N_13528,N_13265);
and U14343 (N_14343,N_13371,N_13409);
nand U14344 (N_14344,N_13569,N_13650);
nor U14345 (N_14345,N_13227,N_13268);
xnor U14346 (N_14346,N_13256,N_13625);
nor U14347 (N_14347,N_13537,N_13630);
and U14348 (N_14348,N_13544,N_13556);
xor U14349 (N_14349,N_13358,N_13402);
or U14350 (N_14350,N_13567,N_13341);
nand U14351 (N_14351,N_13499,N_13372);
xor U14352 (N_14352,N_13380,N_13735);
or U14353 (N_14353,N_13723,N_13795);
xnor U14354 (N_14354,N_13236,N_13747);
or U14355 (N_14355,N_13456,N_13577);
nand U14356 (N_14356,N_13783,N_13754);
nand U14357 (N_14357,N_13578,N_13554);
nand U14358 (N_14358,N_13313,N_13322);
or U14359 (N_14359,N_13462,N_13791);
xnor U14360 (N_14360,N_13368,N_13265);
or U14361 (N_14361,N_13762,N_13407);
and U14362 (N_14362,N_13684,N_13633);
or U14363 (N_14363,N_13532,N_13205);
nor U14364 (N_14364,N_13697,N_13795);
and U14365 (N_14365,N_13713,N_13797);
nor U14366 (N_14366,N_13551,N_13515);
and U14367 (N_14367,N_13384,N_13593);
nor U14368 (N_14368,N_13645,N_13452);
xor U14369 (N_14369,N_13393,N_13288);
xnor U14370 (N_14370,N_13434,N_13460);
and U14371 (N_14371,N_13300,N_13669);
xor U14372 (N_14372,N_13286,N_13278);
nor U14373 (N_14373,N_13293,N_13284);
and U14374 (N_14374,N_13710,N_13292);
nand U14375 (N_14375,N_13599,N_13604);
nor U14376 (N_14376,N_13698,N_13439);
nand U14377 (N_14377,N_13768,N_13659);
nor U14378 (N_14378,N_13555,N_13233);
nand U14379 (N_14379,N_13769,N_13604);
nand U14380 (N_14380,N_13438,N_13246);
nand U14381 (N_14381,N_13371,N_13269);
nor U14382 (N_14382,N_13570,N_13671);
xor U14383 (N_14383,N_13701,N_13637);
or U14384 (N_14384,N_13219,N_13483);
and U14385 (N_14385,N_13228,N_13209);
or U14386 (N_14386,N_13657,N_13301);
nor U14387 (N_14387,N_13593,N_13718);
nor U14388 (N_14388,N_13469,N_13373);
xor U14389 (N_14389,N_13347,N_13656);
nand U14390 (N_14390,N_13520,N_13627);
nand U14391 (N_14391,N_13654,N_13783);
nand U14392 (N_14392,N_13575,N_13378);
or U14393 (N_14393,N_13767,N_13720);
or U14394 (N_14394,N_13357,N_13727);
or U14395 (N_14395,N_13264,N_13436);
or U14396 (N_14396,N_13645,N_13300);
nor U14397 (N_14397,N_13567,N_13761);
and U14398 (N_14398,N_13684,N_13228);
nand U14399 (N_14399,N_13286,N_13710);
xnor U14400 (N_14400,N_13864,N_14346);
or U14401 (N_14401,N_13879,N_14126);
and U14402 (N_14402,N_14107,N_14032);
nand U14403 (N_14403,N_14080,N_13935);
nand U14404 (N_14404,N_13900,N_14008);
nand U14405 (N_14405,N_14184,N_14097);
or U14406 (N_14406,N_14007,N_14054);
or U14407 (N_14407,N_13883,N_14254);
or U14408 (N_14408,N_14196,N_13819);
or U14409 (N_14409,N_14283,N_14015);
nor U14410 (N_14410,N_14278,N_14231);
nor U14411 (N_14411,N_14058,N_13895);
and U14412 (N_14412,N_14325,N_14379);
xnor U14413 (N_14413,N_13807,N_14153);
or U14414 (N_14414,N_14047,N_14089);
and U14415 (N_14415,N_14049,N_14189);
nor U14416 (N_14416,N_14033,N_14034);
nor U14417 (N_14417,N_13830,N_14030);
and U14418 (N_14418,N_14082,N_13832);
nor U14419 (N_14419,N_14165,N_14317);
xnor U14420 (N_14420,N_14155,N_13995);
nor U14421 (N_14421,N_14263,N_14255);
nand U14422 (N_14422,N_14182,N_14356);
or U14423 (N_14423,N_14077,N_14187);
nor U14424 (N_14424,N_14068,N_14177);
nand U14425 (N_14425,N_13925,N_14171);
nor U14426 (N_14426,N_14223,N_14136);
nor U14427 (N_14427,N_14198,N_14301);
and U14428 (N_14428,N_14072,N_13981);
xnor U14429 (N_14429,N_14133,N_13839);
or U14430 (N_14430,N_14370,N_14363);
or U14431 (N_14431,N_14134,N_13941);
nor U14432 (N_14432,N_14069,N_13814);
and U14433 (N_14433,N_14200,N_14152);
or U14434 (N_14434,N_14217,N_13805);
and U14435 (N_14435,N_13873,N_14002);
nand U14436 (N_14436,N_14391,N_14230);
or U14437 (N_14437,N_14161,N_14139);
and U14438 (N_14438,N_14237,N_14169);
or U14439 (N_14439,N_14327,N_14336);
nor U14440 (N_14440,N_14185,N_13823);
and U14441 (N_14441,N_14251,N_14326);
nor U14442 (N_14442,N_14113,N_13829);
nor U14443 (N_14443,N_14202,N_13937);
and U14444 (N_14444,N_14086,N_13970);
xnor U14445 (N_14445,N_14296,N_14221);
xnor U14446 (N_14446,N_14065,N_14112);
nor U14447 (N_14447,N_13847,N_13994);
nor U14448 (N_14448,N_14059,N_13863);
xnor U14449 (N_14449,N_13817,N_14249);
and U14450 (N_14450,N_14118,N_14061);
nand U14451 (N_14451,N_13905,N_14269);
and U14452 (N_14452,N_13802,N_14053);
or U14453 (N_14453,N_14273,N_14351);
nor U14454 (N_14454,N_13979,N_13950);
nand U14455 (N_14455,N_13841,N_14037);
nand U14456 (N_14456,N_14084,N_14384);
nor U14457 (N_14457,N_14124,N_14398);
nor U14458 (N_14458,N_14195,N_14312);
xnor U14459 (N_14459,N_13953,N_14019);
nand U14460 (N_14460,N_13877,N_13977);
nor U14461 (N_14461,N_13804,N_13811);
and U14462 (N_14462,N_13851,N_14151);
and U14463 (N_14463,N_13891,N_14274);
or U14464 (N_14464,N_13971,N_14396);
and U14465 (N_14465,N_13836,N_14399);
nand U14466 (N_14466,N_14244,N_14104);
nand U14467 (N_14467,N_14243,N_14388);
nor U14468 (N_14468,N_13958,N_13915);
nand U14469 (N_14469,N_13872,N_13813);
or U14470 (N_14470,N_14166,N_14102);
xnor U14471 (N_14471,N_14036,N_14295);
xor U14472 (N_14472,N_14150,N_14120);
xnor U14473 (N_14473,N_14383,N_13800);
xnor U14474 (N_14474,N_14309,N_13869);
and U14475 (N_14475,N_14228,N_14108);
or U14476 (N_14476,N_13985,N_14361);
nor U14477 (N_14477,N_14335,N_14375);
and U14478 (N_14478,N_14191,N_13833);
or U14479 (N_14479,N_13892,N_14143);
nor U14480 (N_14480,N_14313,N_14311);
and U14481 (N_14481,N_14055,N_13973);
nand U14482 (N_14482,N_14103,N_13907);
nor U14483 (N_14483,N_14329,N_13975);
or U14484 (N_14484,N_14376,N_14100);
or U14485 (N_14485,N_14048,N_13954);
and U14486 (N_14486,N_13936,N_14129);
or U14487 (N_14487,N_13947,N_13893);
nor U14488 (N_14488,N_14239,N_14178);
or U14489 (N_14489,N_14158,N_14145);
and U14490 (N_14490,N_13894,N_14302);
or U14491 (N_14491,N_13982,N_14211);
nand U14492 (N_14492,N_14156,N_13822);
xnor U14493 (N_14493,N_14157,N_14242);
nand U14494 (N_14494,N_14297,N_13920);
xor U14495 (N_14495,N_14234,N_14260);
nor U14496 (N_14496,N_14027,N_14079);
xnor U14497 (N_14497,N_13926,N_14052);
or U14498 (N_14498,N_14392,N_13992);
nor U14499 (N_14499,N_14083,N_13887);
and U14500 (N_14500,N_13824,N_14352);
and U14501 (N_14501,N_14378,N_14168);
or U14502 (N_14502,N_13838,N_14357);
or U14503 (N_14503,N_14341,N_14138);
nor U14504 (N_14504,N_14360,N_14374);
or U14505 (N_14505,N_14259,N_14394);
nand U14506 (N_14506,N_14170,N_13870);
and U14507 (N_14507,N_14250,N_13875);
nand U14508 (N_14508,N_14247,N_14095);
and U14509 (N_14509,N_14229,N_14193);
nand U14510 (N_14510,N_13845,N_13916);
and U14511 (N_14511,N_13998,N_14088);
xor U14512 (N_14512,N_14012,N_14021);
or U14513 (N_14513,N_14188,N_13943);
nand U14514 (N_14514,N_14010,N_14020);
and U14515 (N_14515,N_13986,N_14262);
nor U14516 (N_14516,N_14206,N_13889);
or U14517 (N_14517,N_14275,N_13821);
and U14518 (N_14518,N_14282,N_14330);
and U14519 (N_14519,N_13878,N_14213);
nand U14520 (N_14520,N_13853,N_13852);
xnor U14521 (N_14521,N_13918,N_13934);
xor U14522 (N_14522,N_14248,N_14321);
or U14523 (N_14523,N_14303,N_13865);
xnor U14524 (N_14524,N_13909,N_14026);
xnor U14525 (N_14525,N_14224,N_13960);
xnor U14526 (N_14526,N_14344,N_13993);
xor U14527 (N_14527,N_14253,N_13964);
nand U14528 (N_14528,N_13886,N_14245);
and U14529 (N_14529,N_14096,N_13850);
or U14530 (N_14530,N_14176,N_14160);
and U14531 (N_14531,N_14240,N_14289);
and U14532 (N_14532,N_14203,N_14114);
and U14533 (N_14533,N_13868,N_13988);
nor U14534 (N_14534,N_13898,N_14261);
xnor U14535 (N_14535,N_13965,N_14241);
nor U14536 (N_14536,N_14039,N_14132);
nor U14537 (N_14537,N_14219,N_14040);
and U14538 (N_14538,N_14149,N_13874);
and U14539 (N_14539,N_13882,N_14005);
xor U14540 (N_14540,N_13902,N_14397);
nand U14541 (N_14541,N_14041,N_13980);
and U14542 (N_14542,N_14286,N_14310);
nor U14543 (N_14543,N_13910,N_13952);
xnor U14544 (N_14544,N_13931,N_14382);
nand U14545 (N_14545,N_14071,N_13999);
xor U14546 (N_14546,N_14137,N_13911);
and U14547 (N_14547,N_13930,N_13978);
or U14548 (N_14548,N_14209,N_14135);
nand U14549 (N_14549,N_13949,N_14285);
nand U14550 (N_14550,N_14090,N_14372);
xnor U14551 (N_14551,N_14130,N_14038);
nor U14552 (N_14552,N_13904,N_14190);
nor U14553 (N_14553,N_14271,N_14226);
xor U14554 (N_14554,N_13884,N_14162);
and U14555 (N_14555,N_14050,N_14179);
nand U14556 (N_14556,N_13976,N_14011);
nand U14557 (N_14557,N_14390,N_14147);
nor U14558 (N_14558,N_14141,N_14081);
xnor U14559 (N_14559,N_14197,N_13932);
nor U14560 (N_14560,N_14334,N_13997);
xor U14561 (N_14561,N_14281,N_14345);
nor U14562 (N_14562,N_14280,N_13806);
or U14563 (N_14563,N_14385,N_13859);
or U14564 (N_14564,N_14101,N_13939);
nand U14565 (N_14565,N_14043,N_13858);
nand U14566 (N_14566,N_14279,N_13834);
xnor U14567 (N_14567,N_14098,N_13956);
and U14568 (N_14568,N_14354,N_14105);
or U14569 (N_14569,N_13974,N_14331);
nand U14570 (N_14570,N_14287,N_13913);
or U14571 (N_14571,N_14121,N_14056);
or U14572 (N_14572,N_14093,N_13854);
xor U14573 (N_14573,N_13843,N_14127);
nand U14574 (N_14574,N_14073,N_14268);
nand U14575 (N_14575,N_14210,N_13987);
xnor U14576 (N_14576,N_14208,N_14023);
nor U14577 (N_14577,N_14042,N_14001);
and U14578 (N_14578,N_13921,N_13996);
xnor U14579 (N_14579,N_14125,N_14235);
nor U14580 (N_14580,N_13881,N_14109);
nor U14581 (N_14581,N_14386,N_14094);
nand U14582 (N_14582,N_14115,N_14377);
nand U14583 (N_14583,N_13924,N_14288);
and U14584 (N_14584,N_14359,N_14045);
and U14585 (N_14585,N_13812,N_14131);
nand U14586 (N_14586,N_14233,N_14324);
xnor U14587 (N_14587,N_14075,N_14181);
nand U14588 (N_14588,N_14099,N_14290);
and U14589 (N_14589,N_14006,N_13951);
xnor U14590 (N_14590,N_14218,N_14348);
nor U14591 (N_14591,N_14332,N_14367);
xor U14592 (N_14592,N_14214,N_14294);
or U14593 (N_14593,N_14057,N_13808);
nor U14594 (N_14594,N_14174,N_13912);
nand U14595 (N_14595,N_14207,N_14364);
and U14596 (N_14596,N_14319,N_13831);
nor U14597 (N_14597,N_13914,N_13827);
nor U14598 (N_14598,N_13957,N_14186);
nand U14599 (N_14599,N_14172,N_14140);
nand U14600 (N_14600,N_14076,N_14175);
nor U14601 (N_14601,N_13967,N_14333);
xor U14602 (N_14602,N_14018,N_14365);
xnor U14603 (N_14603,N_14060,N_13903);
or U14604 (N_14604,N_14343,N_14236);
xnor U14605 (N_14605,N_14201,N_13842);
and U14606 (N_14606,N_13896,N_14142);
nand U14607 (N_14607,N_14117,N_14355);
nand U14608 (N_14608,N_14204,N_14066);
and U14609 (N_14609,N_13849,N_14291);
and U14610 (N_14610,N_13890,N_13933);
and U14611 (N_14611,N_14368,N_14315);
nand U14612 (N_14612,N_14087,N_14265);
xor U14613 (N_14613,N_14144,N_14024);
or U14614 (N_14614,N_13972,N_14222);
nand U14615 (N_14615,N_13908,N_13938);
xor U14616 (N_14616,N_14212,N_13871);
xnor U14617 (N_14617,N_13888,N_14225);
nand U14618 (N_14618,N_14277,N_14320);
xor U14619 (N_14619,N_14063,N_14122);
nor U14620 (N_14620,N_14092,N_14106);
nor U14621 (N_14621,N_14358,N_13917);
nor U14622 (N_14622,N_14276,N_14070);
nor U14623 (N_14623,N_13835,N_13815);
nand U14624 (N_14624,N_14267,N_14393);
xnor U14625 (N_14625,N_14322,N_14270);
xor U14626 (N_14626,N_14318,N_14167);
xnor U14627 (N_14627,N_13828,N_13929);
and U14628 (N_14628,N_14316,N_14299);
xor U14629 (N_14629,N_13848,N_14163);
nor U14630 (N_14630,N_13810,N_13948);
and U14631 (N_14631,N_14252,N_14389);
or U14632 (N_14632,N_14067,N_13899);
nand U14633 (N_14633,N_14028,N_13866);
nand U14634 (N_14634,N_14323,N_14340);
xnor U14635 (N_14635,N_14016,N_14022);
nand U14636 (N_14636,N_14159,N_14293);
and U14637 (N_14637,N_13861,N_14306);
or U14638 (N_14638,N_13968,N_14308);
xnor U14639 (N_14639,N_13818,N_14119);
or U14640 (N_14640,N_14300,N_14246);
nor U14641 (N_14641,N_14232,N_14074);
xor U14642 (N_14642,N_13955,N_14110);
or U14643 (N_14643,N_13961,N_13984);
nand U14644 (N_14644,N_13885,N_14272);
nand U14645 (N_14645,N_14305,N_13989);
xnor U14646 (N_14646,N_14284,N_14349);
or U14647 (N_14647,N_14381,N_14205);
or U14648 (N_14648,N_13857,N_14148);
or U14649 (N_14649,N_13944,N_14128);
nand U14650 (N_14650,N_13901,N_14003);
nor U14651 (N_14651,N_14017,N_14264);
nand U14652 (N_14652,N_13855,N_14258);
xnor U14653 (N_14653,N_14173,N_14000);
and U14654 (N_14654,N_14369,N_13816);
nand U14655 (N_14655,N_14338,N_13963);
nand U14656 (N_14656,N_14123,N_14078);
nand U14657 (N_14657,N_14009,N_13990);
nor U14658 (N_14658,N_13946,N_13801);
nor U14659 (N_14659,N_14371,N_14328);
xnor U14660 (N_14660,N_14292,N_14013);
nand U14661 (N_14661,N_14035,N_13942);
xnor U14662 (N_14662,N_14337,N_13940);
nand U14663 (N_14663,N_14307,N_14154);
xor U14664 (N_14664,N_13923,N_14350);
nor U14665 (N_14665,N_13927,N_13876);
and U14666 (N_14666,N_14192,N_14062);
nand U14667 (N_14667,N_13962,N_14238);
and U14668 (N_14668,N_14373,N_14085);
xor U14669 (N_14669,N_13856,N_14064);
nand U14670 (N_14670,N_14366,N_14347);
and U14671 (N_14671,N_14164,N_13846);
xor U14672 (N_14672,N_13844,N_13840);
nor U14673 (N_14673,N_14116,N_13966);
or U14674 (N_14674,N_14342,N_13862);
and U14675 (N_14675,N_14044,N_14031);
nor U14676 (N_14676,N_14146,N_13922);
nand U14677 (N_14677,N_13919,N_14298);
and U14678 (N_14678,N_14339,N_14199);
nand U14679 (N_14679,N_14362,N_14314);
nand U14680 (N_14680,N_14353,N_13880);
or U14681 (N_14681,N_13897,N_14220);
nor U14682 (N_14682,N_14266,N_14029);
or U14683 (N_14683,N_14046,N_14227);
xnor U14684 (N_14684,N_14215,N_13825);
and U14685 (N_14685,N_14216,N_13826);
nand U14686 (N_14686,N_14051,N_13983);
and U14687 (N_14687,N_14257,N_13860);
nand U14688 (N_14688,N_13837,N_14194);
nor U14689 (N_14689,N_14395,N_13803);
and U14690 (N_14690,N_14387,N_13959);
or U14691 (N_14691,N_13969,N_13991);
xor U14692 (N_14692,N_13820,N_14025);
nor U14693 (N_14693,N_14004,N_14380);
or U14694 (N_14694,N_14014,N_13867);
and U14695 (N_14695,N_13906,N_13928);
and U14696 (N_14696,N_14256,N_14180);
and U14697 (N_14697,N_14111,N_14304);
nand U14698 (N_14698,N_14183,N_13809);
nor U14699 (N_14699,N_13945,N_14091);
or U14700 (N_14700,N_14212,N_14135);
or U14701 (N_14701,N_13989,N_14107);
or U14702 (N_14702,N_13950,N_13956);
and U14703 (N_14703,N_14231,N_13900);
and U14704 (N_14704,N_14121,N_14217);
nor U14705 (N_14705,N_13858,N_14215);
nor U14706 (N_14706,N_14283,N_14148);
nand U14707 (N_14707,N_14005,N_13977);
nand U14708 (N_14708,N_14337,N_14142);
or U14709 (N_14709,N_14358,N_14334);
xnor U14710 (N_14710,N_14101,N_13921);
and U14711 (N_14711,N_14371,N_14049);
and U14712 (N_14712,N_14358,N_14333);
or U14713 (N_14713,N_14256,N_14287);
or U14714 (N_14714,N_14057,N_14346);
nand U14715 (N_14715,N_13815,N_14021);
nor U14716 (N_14716,N_14083,N_14103);
nor U14717 (N_14717,N_14220,N_13875);
nor U14718 (N_14718,N_14094,N_14053);
and U14719 (N_14719,N_13949,N_14138);
nand U14720 (N_14720,N_13854,N_14015);
nand U14721 (N_14721,N_14307,N_14109);
and U14722 (N_14722,N_13913,N_13827);
xor U14723 (N_14723,N_14135,N_13969);
nand U14724 (N_14724,N_13958,N_14232);
or U14725 (N_14725,N_14361,N_14000);
xor U14726 (N_14726,N_14339,N_14315);
and U14727 (N_14727,N_13966,N_14208);
xor U14728 (N_14728,N_14360,N_13980);
or U14729 (N_14729,N_14028,N_14291);
nand U14730 (N_14730,N_14313,N_14379);
and U14731 (N_14731,N_14207,N_13958);
and U14732 (N_14732,N_14240,N_13879);
nor U14733 (N_14733,N_14257,N_13911);
nand U14734 (N_14734,N_13960,N_14272);
nor U14735 (N_14735,N_13804,N_14158);
xnor U14736 (N_14736,N_14040,N_14342);
xor U14737 (N_14737,N_13863,N_13809);
and U14738 (N_14738,N_14314,N_14255);
nor U14739 (N_14739,N_13903,N_13815);
or U14740 (N_14740,N_14092,N_14385);
xnor U14741 (N_14741,N_13800,N_14205);
nor U14742 (N_14742,N_13817,N_14224);
or U14743 (N_14743,N_14018,N_14179);
xor U14744 (N_14744,N_14086,N_14330);
xor U14745 (N_14745,N_13902,N_14267);
xnor U14746 (N_14746,N_14012,N_14148);
or U14747 (N_14747,N_14127,N_14080);
nor U14748 (N_14748,N_14142,N_14182);
and U14749 (N_14749,N_13916,N_13921);
xor U14750 (N_14750,N_14045,N_14317);
and U14751 (N_14751,N_14163,N_14067);
nand U14752 (N_14752,N_14261,N_14232);
or U14753 (N_14753,N_14092,N_13936);
nor U14754 (N_14754,N_13895,N_14117);
or U14755 (N_14755,N_14346,N_14085);
or U14756 (N_14756,N_13918,N_13922);
or U14757 (N_14757,N_13910,N_14065);
nor U14758 (N_14758,N_14011,N_14042);
and U14759 (N_14759,N_13940,N_14236);
or U14760 (N_14760,N_13986,N_13809);
and U14761 (N_14761,N_14073,N_14213);
or U14762 (N_14762,N_14183,N_14284);
nor U14763 (N_14763,N_14049,N_13845);
xor U14764 (N_14764,N_14164,N_14202);
xor U14765 (N_14765,N_14268,N_13844);
nor U14766 (N_14766,N_14371,N_14022);
nand U14767 (N_14767,N_14157,N_14102);
xnor U14768 (N_14768,N_13829,N_14034);
nand U14769 (N_14769,N_13921,N_14274);
and U14770 (N_14770,N_13914,N_14027);
nand U14771 (N_14771,N_13913,N_14346);
or U14772 (N_14772,N_13997,N_14321);
nor U14773 (N_14773,N_13941,N_14095);
nand U14774 (N_14774,N_14228,N_14142);
or U14775 (N_14775,N_14104,N_14226);
and U14776 (N_14776,N_14312,N_14040);
nor U14777 (N_14777,N_13856,N_14316);
and U14778 (N_14778,N_14181,N_14305);
nand U14779 (N_14779,N_14382,N_14090);
nand U14780 (N_14780,N_14292,N_14050);
nor U14781 (N_14781,N_14383,N_14210);
nand U14782 (N_14782,N_13926,N_14085);
nand U14783 (N_14783,N_13863,N_13974);
or U14784 (N_14784,N_13984,N_14125);
xnor U14785 (N_14785,N_13954,N_13822);
xnor U14786 (N_14786,N_14045,N_13902);
or U14787 (N_14787,N_13957,N_14345);
nand U14788 (N_14788,N_13864,N_14292);
or U14789 (N_14789,N_14312,N_14355);
xor U14790 (N_14790,N_14313,N_13963);
nor U14791 (N_14791,N_14152,N_14360);
and U14792 (N_14792,N_14345,N_14095);
xor U14793 (N_14793,N_14341,N_14267);
and U14794 (N_14794,N_14235,N_14265);
nor U14795 (N_14795,N_14290,N_14101);
xnor U14796 (N_14796,N_13871,N_14215);
nor U14797 (N_14797,N_13963,N_14085);
or U14798 (N_14798,N_13817,N_13948);
or U14799 (N_14799,N_14288,N_13936);
xor U14800 (N_14800,N_14177,N_14269);
xor U14801 (N_14801,N_13860,N_13942);
and U14802 (N_14802,N_13921,N_13993);
xor U14803 (N_14803,N_14139,N_14291);
nand U14804 (N_14804,N_14365,N_14197);
and U14805 (N_14805,N_14226,N_14230);
and U14806 (N_14806,N_14133,N_14282);
and U14807 (N_14807,N_14121,N_13831);
nand U14808 (N_14808,N_13855,N_14043);
nand U14809 (N_14809,N_14066,N_14210);
nor U14810 (N_14810,N_13801,N_14036);
nand U14811 (N_14811,N_14093,N_14357);
nor U14812 (N_14812,N_14349,N_14044);
nor U14813 (N_14813,N_13906,N_13918);
and U14814 (N_14814,N_14307,N_14343);
xor U14815 (N_14815,N_13844,N_14146);
and U14816 (N_14816,N_14372,N_14263);
nor U14817 (N_14817,N_14087,N_13851);
and U14818 (N_14818,N_14246,N_13882);
nor U14819 (N_14819,N_13869,N_14378);
xor U14820 (N_14820,N_14091,N_14269);
nand U14821 (N_14821,N_14044,N_14067);
nor U14822 (N_14822,N_14393,N_14172);
nor U14823 (N_14823,N_14281,N_14227);
nand U14824 (N_14824,N_13906,N_14138);
nor U14825 (N_14825,N_14249,N_14327);
nand U14826 (N_14826,N_13837,N_14356);
and U14827 (N_14827,N_14100,N_13932);
xnor U14828 (N_14828,N_13935,N_13891);
or U14829 (N_14829,N_13856,N_14250);
or U14830 (N_14830,N_14116,N_14127);
nand U14831 (N_14831,N_14342,N_13857);
nor U14832 (N_14832,N_13980,N_14343);
and U14833 (N_14833,N_14054,N_14043);
nor U14834 (N_14834,N_13815,N_13988);
nor U14835 (N_14835,N_13860,N_14334);
nand U14836 (N_14836,N_14119,N_14100);
xnor U14837 (N_14837,N_14270,N_14089);
xnor U14838 (N_14838,N_14160,N_14057);
nand U14839 (N_14839,N_14014,N_14164);
or U14840 (N_14840,N_13897,N_14328);
and U14841 (N_14841,N_14291,N_14104);
or U14842 (N_14842,N_13900,N_14207);
xor U14843 (N_14843,N_14329,N_14382);
nor U14844 (N_14844,N_14176,N_14226);
and U14845 (N_14845,N_13894,N_13887);
and U14846 (N_14846,N_14021,N_14344);
nor U14847 (N_14847,N_14224,N_14357);
xor U14848 (N_14848,N_14066,N_13837);
or U14849 (N_14849,N_14355,N_14338);
nand U14850 (N_14850,N_14124,N_13995);
and U14851 (N_14851,N_14202,N_13819);
and U14852 (N_14852,N_14314,N_13952);
nand U14853 (N_14853,N_14201,N_14030);
nand U14854 (N_14854,N_13878,N_14120);
xor U14855 (N_14855,N_13904,N_13860);
nand U14856 (N_14856,N_14367,N_13964);
nor U14857 (N_14857,N_14139,N_14390);
nor U14858 (N_14858,N_14297,N_14162);
or U14859 (N_14859,N_14099,N_13990);
and U14860 (N_14860,N_14325,N_13881);
or U14861 (N_14861,N_14163,N_14320);
nand U14862 (N_14862,N_13879,N_13860);
nor U14863 (N_14863,N_14394,N_13974);
nand U14864 (N_14864,N_13924,N_14071);
or U14865 (N_14865,N_13926,N_13869);
and U14866 (N_14866,N_13851,N_14116);
xnor U14867 (N_14867,N_14060,N_13963);
nor U14868 (N_14868,N_14118,N_14037);
nand U14869 (N_14869,N_14186,N_14252);
and U14870 (N_14870,N_14259,N_14205);
or U14871 (N_14871,N_14012,N_14238);
and U14872 (N_14872,N_14064,N_14022);
or U14873 (N_14873,N_14088,N_14315);
xnor U14874 (N_14874,N_13905,N_14298);
and U14875 (N_14875,N_14022,N_13901);
and U14876 (N_14876,N_14081,N_14349);
and U14877 (N_14877,N_13853,N_13901);
nand U14878 (N_14878,N_13908,N_14157);
or U14879 (N_14879,N_14384,N_13901);
nand U14880 (N_14880,N_14307,N_14193);
nor U14881 (N_14881,N_14039,N_13934);
nor U14882 (N_14882,N_14154,N_14223);
xor U14883 (N_14883,N_14266,N_14337);
xnor U14884 (N_14884,N_14277,N_13859);
and U14885 (N_14885,N_13995,N_14207);
nor U14886 (N_14886,N_13838,N_13811);
or U14887 (N_14887,N_14044,N_13809);
or U14888 (N_14888,N_14089,N_14350);
xor U14889 (N_14889,N_14217,N_13994);
and U14890 (N_14890,N_14373,N_14017);
nand U14891 (N_14891,N_13879,N_14125);
or U14892 (N_14892,N_14232,N_14118);
or U14893 (N_14893,N_14084,N_13908);
nand U14894 (N_14894,N_14213,N_13865);
and U14895 (N_14895,N_13895,N_14391);
and U14896 (N_14896,N_14121,N_14375);
or U14897 (N_14897,N_14328,N_13956);
and U14898 (N_14898,N_14089,N_13926);
or U14899 (N_14899,N_13950,N_14191);
and U14900 (N_14900,N_14396,N_13909);
or U14901 (N_14901,N_14384,N_14119);
or U14902 (N_14902,N_14314,N_14087);
nand U14903 (N_14903,N_14361,N_14373);
and U14904 (N_14904,N_14063,N_14036);
xor U14905 (N_14905,N_13876,N_14053);
nand U14906 (N_14906,N_14116,N_14277);
or U14907 (N_14907,N_14228,N_13995);
xor U14908 (N_14908,N_14221,N_14120);
or U14909 (N_14909,N_14358,N_14082);
xnor U14910 (N_14910,N_13821,N_14255);
and U14911 (N_14911,N_13903,N_14394);
xor U14912 (N_14912,N_14358,N_14085);
nand U14913 (N_14913,N_13893,N_14025);
nand U14914 (N_14914,N_13964,N_14399);
or U14915 (N_14915,N_13950,N_14212);
nand U14916 (N_14916,N_14097,N_14356);
nand U14917 (N_14917,N_14241,N_14328);
and U14918 (N_14918,N_13800,N_14357);
xor U14919 (N_14919,N_13911,N_14037);
nor U14920 (N_14920,N_13992,N_13837);
or U14921 (N_14921,N_14028,N_14186);
and U14922 (N_14922,N_13941,N_14301);
or U14923 (N_14923,N_13819,N_14205);
or U14924 (N_14924,N_14157,N_13803);
and U14925 (N_14925,N_13914,N_14120);
or U14926 (N_14926,N_14152,N_14252);
nand U14927 (N_14927,N_14148,N_14356);
nand U14928 (N_14928,N_14023,N_14362);
and U14929 (N_14929,N_13912,N_14296);
nor U14930 (N_14930,N_14053,N_14272);
and U14931 (N_14931,N_14290,N_13983);
and U14932 (N_14932,N_13848,N_14059);
and U14933 (N_14933,N_13909,N_14022);
xor U14934 (N_14934,N_13975,N_14134);
or U14935 (N_14935,N_14237,N_14259);
or U14936 (N_14936,N_14109,N_14131);
or U14937 (N_14937,N_14320,N_14203);
or U14938 (N_14938,N_14211,N_14310);
nor U14939 (N_14939,N_13803,N_13836);
or U14940 (N_14940,N_14210,N_14001);
nand U14941 (N_14941,N_14046,N_14034);
or U14942 (N_14942,N_14031,N_13865);
and U14943 (N_14943,N_13874,N_14143);
nand U14944 (N_14944,N_14142,N_13972);
nor U14945 (N_14945,N_14253,N_13848);
xor U14946 (N_14946,N_14066,N_14235);
and U14947 (N_14947,N_14120,N_13947);
or U14948 (N_14948,N_13847,N_13838);
nand U14949 (N_14949,N_14063,N_13983);
xnor U14950 (N_14950,N_14341,N_14010);
nand U14951 (N_14951,N_13931,N_14248);
nand U14952 (N_14952,N_14235,N_14216);
and U14953 (N_14953,N_14195,N_14252);
nand U14954 (N_14954,N_14017,N_13884);
or U14955 (N_14955,N_14237,N_13976);
xor U14956 (N_14956,N_14173,N_14242);
and U14957 (N_14957,N_14391,N_13928);
or U14958 (N_14958,N_14256,N_13934);
nand U14959 (N_14959,N_13967,N_14237);
xor U14960 (N_14960,N_14173,N_14099);
xnor U14961 (N_14961,N_13840,N_14052);
or U14962 (N_14962,N_14079,N_14024);
or U14963 (N_14963,N_14041,N_13978);
nor U14964 (N_14964,N_14341,N_14332);
nand U14965 (N_14965,N_14342,N_13861);
or U14966 (N_14966,N_14307,N_14039);
nor U14967 (N_14967,N_13940,N_13893);
nor U14968 (N_14968,N_13895,N_14236);
nand U14969 (N_14969,N_14040,N_14153);
or U14970 (N_14970,N_13943,N_13830);
and U14971 (N_14971,N_14052,N_13844);
xor U14972 (N_14972,N_13875,N_14137);
and U14973 (N_14973,N_14359,N_14069);
or U14974 (N_14974,N_14180,N_14273);
nor U14975 (N_14975,N_14030,N_14075);
nand U14976 (N_14976,N_13962,N_13890);
nand U14977 (N_14977,N_14221,N_14008);
and U14978 (N_14978,N_14101,N_13844);
xnor U14979 (N_14979,N_13841,N_14085);
or U14980 (N_14980,N_14199,N_14066);
or U14981 (N_14981,N_14301,N_13864);
and U14982 (N_14982,N_13925,N_14113);
and U14983 (N_14983,N_13972,N_14306);
nand U14984 (N_14984,N_13966,N_14027);
or U14985 (N_14985,N_14312,N_14025);
and U14986 (N_14986,N_14188,N_14247);
and U14987 (N_14987,N_14381,N_13993);
nand U14988 (N_14988,N_14364,N_13939);
and U14989 (N_14989,N_14032,N_14123);
and U14990 (N_14990,N_14240,N_14213);
and U14991 (N_14991,N_13948,N_14034);
xor U14992 (N_14992,N_14195,N_13833);
nor U14993 (N_14993,N_14016,N_14027);
or U14994 (N_14994,N_14339,N_13914);
and U14995 (N_14995,N_14384,N_13892);
nor U14996 (N_14996,N_14150,N_14322);
nand U14997 (N_14997,N_13981,N_14004);
and U14998 (N_14998,N_13820,N_14124);
or U14999 (N_14999,N_13905,N_14124);
or U15000 (N_15000,N_14412,N_14549);
nor U15001 (N_15001,N_14806,N_14661);
and U15002 (N_15002,N_14708,N_14568);
nand U15003 (N_15003,N_14645,N_14490);
and U15004 (N_15004,N_14747,N_14590);
nor U15005 (N_15005,N_14581,N_14666);
nand U15006 (N_15006,N_14947,N_14693);
and U15007 (N_15007,N_14919,N_14959);
and U15008 (N_15008,N_14610,N_14470);
nor U15009 (N_15009,N_14658,N_14726);
nor U15010 (N_15010,N_14837,N_14773);
xor U15011 (N_15011,N_14636,N_14712);
or U15012 (N_15012,N_14824,N_14691);
xor U15013 (N_15013,N_14847,N_14879);
or U15014 (N_15014,N_14997,N_14598);
and U15015 (N_15015,N_14626,N_14809);
nor U15016 (N_15016,N_14755,N_14520);
nand U15017 (N_15017,N_14985,N_14438);
and U15018 (N_15018,N_14845,N_14701);
nor U15019 (N_15019,N_14830,N_14772);
or U15020 (N_15020,N_14484,N_14664);
or U15021 (N_15021,N_14776,N_14565);
nand U15022 (N_15022,N_14469,N_14711);
and U15023 (N_15023,N_14405,N_14494);
and U15024 (N_15024,N_14508,N_14482);
and U15025 (N_15025,N_14753,N_14514);
nor U15026 (N_15026,N_14991,N_14646);
or U15027 (N_15027,N_14870,N_14688);
nor U15028 (N_15028,N_14861,N_14439);
nand U15029 (N_15029,N_14450,N_14673);
or U15030 (N_15030,N_14987,N_14572);
nor U15031 (N_15031,N_14510,N_14551);
xor U15032 (N_15032,N_14805,N_14752);
nor U15033 (N_15033,N_14675,N_14952);
and U15034 (N_15034,N_14642,N_14634);
xnor U15035 (N_15035,N_14877,N_14523);
and U15036 (N_15036,N_14573,N_14721);
and U15037 (N_15037,N_14969,N_14769);
nand U15038 (N_15038,N_14791,N_14631);
and U15039 (N_15039,N_14865,N_14995);
or U15040 (N_15040,N_14818,N_14637);
xor U15041 (N_15041,N_14804,N_14859);
and U15042 (N_15042,N_14775,N_14992);
nand U15043 (N_15043,N_14671,N_14933);
nand U15044 (N_15044,N_14436,N_14623);
and U15045 (N_15045,N_14736,N_14846);
or U15046 (N_15046,N_14867,N_14717);
nor U15047 (N_15047,N_14541,N_14875);
and U15048 (N_15048,N_14702,N_14910);
xor U15049 (N_15049,N_14425,N_14593);
xor U15050 (N_15050,N_14869,N_14617);
or U15051 (N_15051,N_14902,N_14962);
nor U15052 (N_15052,N_14492,N_14827);
nand U15053 (N_15053,N_14421,N_14417);
xnor U15054 (N_15054,N_14912,N_14978);
and U15055 (N_15055,N_14588,N_14785);
nand U15056 (N_15056,N_14885,N_14532);
and U15057 (N_15057,N_14653,N_14457);
nand U15058 (N_15058,N_14624,N_14676);
and U15059 (N_15059,N_14918,N_14967);
or U15060 (N_15060,N_14871,N_14531);
xor U15061 (N_15061,N_14718,N_14451);
nand U15062 (N_15062,N_14850,N_14760);
and U15063 (N_15063,N_14665,N_14862);
or U15064 (N_15064,N_14955,N_14698);
nor U15065 (N_15065,N_14853,N_14834);
nand U15066 (N_15066,N_14468,N_14683);
or U15067 (N_15067,N_14836,N_14504);
nand U15068 (N_15068,N_14619,N_14560);
xnor U15069 (N_15069,N_14518,N_14731);
nand U15070 (N_15070,N_14603,N_14849);
or U15071 (N_15071,N_14414,N_14433);
or U15072 (N_15072,N_14872,N_14895);
and U15073 (N_15073,N_14897,N_14567);
nand U15074 (N_15074,N_14766,N_14607);
nor U15075 (N_15075,N_14722,N_14608);
xnor U15076 (N_15076,N_14855,N_14427);
and U15077 (N_15077,N_14898,N_14915);
and U15078 (N_15078,N_14822,N_14787);
and U15079 (N_15079,N_14615,N_14880);
nor U15080 (N_15080,N_14570,N_14444);
nand U15081 (N_15081,N_14876,N_14975);
nor U15082 (N_15082,N_14538,N_14627);
nand U15083 (N_15083,N_14957,N_14900);
nor U15084 (N_15084,N_14700,N_14909);
nand U15085 (N_15085,N_14908,N_14448);
and U15086 (N_15086,N_14467,N_14562);
xnor U15087 (N_15087,N_14556,N_14437);
nor U15088 (N_15088,N_14690,N_14651);
and U15089 (N_15089,N_14509,N_14486);
or U15090 (N_15090,N_14621,N_14481);
nand U15091 (N_15091,N_14612,N_14888);
and U15092 (N_15092,N_14783,N_14496);
and U15093 (N_15093,N_14793,N_14662);
and U15094 (N_15094,N_14543,N_14901);
and U15095 (N_15095,N_14819,N_14498);
xor U15096 (N_15096,N_14751,N_14817);
nand U15097 (N_15097,N_14782,N_14516);
and U15098 (N_15098,N_14848,N_14950);
xnor U15099 (N_15099,N_14931,N_14537);
xnor U15100 (N_15100,N_14887,N_14554);
or U15101 (N_15101,N_14935,N_14655);
xnor U15102 (N_15102,N_14595,N_14512);
or U15103 (N_15103,N_14811,N_14685);
and U15104 (N_15104,N_14944,N_14795);
nand U15105 (N_15105,N_14670,N_14695);
xnor U15106 (N_15106,N_14828,N_14426);
nand U15107 (N_15107,N_14737,N_14424);
or U15108 (N_15108,N_14639,N_14422);
xnor U15109 (N_15109,N_14728,N_14841);
nor U15110 (N_15110,N_14445,N_14899);
and U15111 (N_15111,N_14638,N_14896);
and U15112 (N_15112,N_14868,N_14584);
nor U15113 (N_15113,N_14812,N_14535);
or U15114 (N_15114,N_14792,N_14856);
xor U15115 (N_15115,N_14917,N_14883);
nor U15116 (N_15116,N_14943,N_14413);
and U15117 (N_15117,N_14613,N_14420);
and U15118 (N_15118,N_14526,N_14789);
nor U15119 (N_15119,N_14925,N_14431);
xnor U15120 (N_15120,N_14659,N_14720);
and U15121 (N_15121,N_14546,N_14432);
nor U15122 (N_15122,N_14843,N_14999);
xor U15123 (N_15123,N_14545,N_14493);
or U15124 (N_15124,N_14986,N_14694);
nand U15125 (N_15125,N_14686,N_14808);
or U15126 (N_15126,N_14790,N_14640);
nor U15127 (N_15127,N_14458,N_14566);
and U15128 (N_15128,N_14831,N_14744);
nor U15129 (N_15129,N_14650,N_14977);
nand U15130 (N_15130,N_14784,N_14973);
xnor U15131 (N_15131,N_14559,N_14480);
xor U15132 (N_15132,N_14697,N_14974);
xnor U15133 (N_15133,N_14982,N_14681);
xnor U15134 (N_15134,N_14501,N_14968);
xnor U15135 (N_15135,N_14716,N_14506);
or U15136 (N_15136,N_14852,N_14663);
nand U15137 (N_15137,N_14699,N_14878);
xnor U15138 (N_15138,N_14723,N_14507);
xor U15139 (N_15139,N_14739,N_14778);
and U15140 (N_15140,N_14522,N_14528);
nand U15141 (N_15141,N_14605,N_14553);
or U15142 (N_15142,N_14929,N_14600);
nor U15143 (N_15143,N_14732,N_14601);
nand U15144 (N_15144,N_14630,N_14561);
xnor U15145 (N_15145,N_14988,N_14569);
nor U15146 (N_15146,N_14749,N_14927);
xnor U15147 (N_15147,N_14799,N_14840);
xor U15148 (N_15148,N_14449,N_14548);
or U15149 (N_15149,N_14976,N_14625);
nand U15150 (N_15150,N_14611,N_14904);
nor U15151 (N_15151,N_14485,N_14923);
and U15152 (N_15152,N_14460,N_14418);
nand U15153 (N_15153,N_14403,N_14768);
nand U15154 (N_15154,N_14555,N_14402);
xor U15155 (N_15155,N_14594,N_14980);
or U15156 (N_15156,N_14415,N_14533);
and U15157 (N_15157,N_14668,N_14463);
or U15158 (N_15158,N_14550,N_14464);
nand U15159 (N_15159,N_14710,N_14972);
nand U15160 (N_15160,N_14802,N_14916);
nor U15161 (N_15161,N_14656,N_14680);
nand U15162 (N_15162,N_14609,N_14741);
xor U15163 (N_15163,N_14563,N_14578);
nand U15164 (N_15164,N_14735,N_14539);
nand U15165 (N_15165,N_14644,N_14410);
and U15166 (N_15166,N_14956,N_14993);
xor U15167 (N_15167,N_14928,N_14704);
xnor U15168 (N_15168,N_14602,N_14483);
and U15169 (N_15169,N_14527,N_14941);
xor U15170 (N_15170,N_14654,N_14443);
and U15171 (N_15171,N_14838,N_14798);
or U15172 (N_15172,N_14477,N_14459);
nor U15173 (N_15173,N_14961,N_14674);
xor U15174 (N_15174,N_14821,N_14715);
or U15175 (N_15175,N_14816,N_14796);
nand U15176 (N_15176,N_14954,N_14903);
xnor U15177 (N_15177,N_14404,N_14536);
or U15178 (N_15178,N_14564,N_14971);
or U15179 (N_15179,N_14970,N_14488);
nor U15180 (N_15180,N_14660,N_14814);
nand U15181 (N_15181,N_14779,N_14599);
and U15182 (N_15182,N_14505,N_14921);
nor U15183 (N_15183,N_14525,N_14589);
and U15184 (N_15184,N_14951,N_14489);
xor U15185 (N_15185,N_14705,N_14647);
xor U15186 (N_15186,N_14616,N_14765);
nor U15187 (N_15187,N_14430,N_14781);
nand U15188 (N_15188,N_14428,N_14472);
or U15189 (N_15189,N_14628,N_14979);
or U15190 (N_15190,N_14709,N_14677);
or U15191 (N_15191,N_14487,N_14960);
nor U15192 (N_15192,N_14983,N_14891);
nor U15193 (N_15193,N_14576,N_14825);
or U15194 (N_15194,N_14756,N_14416);
or U15195 (N_15195,N_14920,N_14586);
nand U15196 (N_15196,N_14771,N_14652);
xor U15197 (N_15197,N_14905,N_14641);
nand U15198 (N_15198,N_14734,N_14803);
and U15199 (N_15199,N_14930,N_14558);
xor U15200 (N_15200,N_14629,N_14913);
nand U15201 (N_15201,N_14863,N_14456);
and U15202 (N_15202,N_14733,N_14574);
xor U15203 (N_15203,N_14757,N_14953);
and U15204 (N_15204,N_14965,N_14884);
nand U15205 (N_15205,N_14810,N_14873);
nand U15206 (N_15206,N_14948,N_14860);
nand U15207 (N_15207,N_14832,N_14696);
and U15208 (N_15208,N_14529,N_14727);
or U15209 (N_15209,N_14936,N_14946);
xor U15210 (N_15210,N_14807,N_14742);
and U15211 (N_15211,N_14687,N_14743);
nand U15212 (N_15212,N_14465,N_14440);
nand U15213 (N_15213,N_14706,N_14764);
nor U15214 (N_15214,N_14497,N_14540);
nand U15215 (N_15215,N_14738,N_14866);
and U15216 (N_15216,N_14635,N_14940);
nand U15217 (N_15217,N_14874,N_14767);
or U15218 (N_15218,N_14893,N_14984);
or U15219 (N_15219,N_14761,N_14454);
and U15220 (N_15220,N_14906,N_14746);
or U15221 (N_15221,N_14689,N_14614);
and U15222 (N_15222,N_14476,N_14966);
xor U15223 (N_15223,N_14419,N_14990);
nor U15224 (N_15224,N_14473,N_14552);
or U15225 (N_15225,N_14446,N_14964);
and U15226 (N_15226,N_14981,N_14813);
nor U15227 (N_15227,N_14478,N_14754);
and U15228 (N_15228,N_14547,N_14544);
xor U15229 (N_15229,N_14892,N_14557);
xor U15230 (N_15230,N_14774,N_14713);
or U15231 (N_15231,N_14583,N_14500);
or U15232 (N_15232,N_14434,N_14643);
nand U15233 (N_15233,N_14491,N_14495);
or U15234 (N_15234,N_14934,N_14409);
xor U15235 (N_15235,N_14657,N_14423);
nand U15236 (N_15236,N_14667,N_14582);
or U15237 (N_15237,N_14839,N_14729);
nor U15238 (N_15238,N_14606,N_14442);
xnor U15239 (N_15239,N_14942,N_14530);
or U15240 (N_15240,N_14911,N_14407);
nor U15241 (N_15241,N_14592,N_14914);
nor U15242 (N_15242,N_14435,N_14844);
or U15243 (N_15243,N_14503,N_14447);
xnor U15244 (N_15244,N_14894,N_14429);
or U15245 (N_15245,N_14881,N_14949);
xor U15246 (N_15246,N_14826,N_14684);
nor U15247 (N_15247,N_14763,N_14864);
xnor U15248 (N_15248,N_14406,N_14725);
or U15249 (N_15249,N_14842,N_14703);
nand U15250 (N_15250,N_14998,N_14408);
or U15251 (N_15251,N_14672,N_14740);
nor U15252 (N_15252,N_14882,N_14730);
or U15253 (N_15253,N_14534,N_14829);
xor U15254 (N_15254,N_14707,N_14452);
nand U15255 (N_15255,N_14714,N_14800);
and U15256 (N_15256,N_14474,N_14835);
xor U15257 (N_15257,N_14462,N_14854);
or U15258 (N_15258,N_14937,N_14932);
nand U15259 (N_15259,N_14669,N_14519);
or U15260 (N_15260,N_14633,N_14511);
and U15261 (N_15261,N_14963,N_14939);
xnor U15262 (N_15262,N_14618,N_14945);
or U15263 (N_15263,N_14622,N_14889);
nor U15264 (N_15264,N_14788,N_14400);
or U15265 (N_15265,N_14679,N_14471);
or U15266 (N_15266,N_14801,N_14579);
xor U15267 (N_15267,N_14815,N_14938);
nor U15268 (N_15268,N_14886,N_14411);
nor U15269 (N_15269,N_14620,N_14502);
and U15270 (N_15270,N_14587,N_14648);
nor U15271 (N_15271,N_14571,N_14794);
xnor U15272 (N_15272,N_14907,N_14542);
xnor U15273 (N_15273,N_14748,N_14517);
and U15274 (N_15274,N_14524,N_14479);
nor U15275 (N_15275,N_14890,N_14466);
or U15276 (N_15276,N_14958,N_14575);
or U15277 (N_15277,N_14515,N_14926);
xnor U15278 (N_15278,N_14758,N_14759);
or U15279 (N_15279,N_14649,N_14604);
nand U15280 (N_15280,N_14521,N_14585);
or U15281 (N_15281,N_14989,N_14719);
and U15282 (N_15282,N_14833,N_14513);
or U15283 (N_15283,N_14632,N_14724);
or U15284 (N_15284,N_14692,N_14453);
xor U15285 (N_15285,N_14475,N_14762);
xnor U15286 (N_15286,N_14597,N_14455);
nand U15287 (N_15287,N_14858,N_14851);
xnor U15288 (N_15288,N_14591,N_14786);
and U15289 (N_15289,N_14596,N_14820);
nand U15290 (N_15290,N_14745,N_14797);
or U15291 (N_15291,N_14777,N_14922);
xnor U15292 (N_15292,N_14678,N_14401);
or U15293 (N_15293,N_14857,N_14770);
nor U15294 (N_15294,N_14499,N_14924);
xor U15295 (N_15295,N_14750,N_14994);
and U15296 (N_15296,N_14823,N_14461);
and U15297 (N_15297,N_14577,N_14682);
and U15298 (N_15298,N_14441,N_14580);
nor U15299 (N_15299,N_14996,N_14780);
and U15300 (N_15300,N_14508,N_14752);
xor U15301 (N_15301,N_14798,N_14702);
or U15302 (N_15302,N_14803,N_14460);
xor U15303 (N_15303,N_14782,N_14404);
nor U15304 (N_15304,N_14587,N_14820);
and U15305 (N_15305,N_14985,N_14654);
or U15306 (N_15306,N_14597,N_14939);
and U15307 (N_15307,N_14971,N_14520);
xnor U15308 (N_15308,N_14575,N_14540);
nand U15309 (N_15309,N_14910,N_14900);
xnor U15310 (N_15310,N_14951,N_14543);
or U15311 (N_15311,N_14485,N_14749);
nor U15312 (N_15312,N_14583,N_14906);
or U15313 (N_15313,N_14858,N_14978);
xor U15314 (N_15314,N_14945,N_14971);
and U15315 (N_15315,N_14836,N_14589);
and U15316 (N_15316,N_14836,N_14947);
or U15317 (N_15317,N_14441,N_14599);
or U15318 (N_15318,N_14752,N_14870);
and U15319 (N_15319,N_14757,N_14459);
nand U15320 (N_15320,N_14719,N_14421);
xnor U15321 (N_15321,N_14988,N_14643);
nor U15322 (N_15322,N_14971,N_14583);
and U15323 (N_15323,N_14763,N_14854);
xor U15324 (N_15324,N_14853,N_14790);
and U15325 (N_15325,N_14552,N_14880);
or U15326 (N_15326,N_14565,N_14498);
and U15327 (N_15327,N_14415,N_14508);
nand U15328 (N_15328,N_14913,N_14475);
nor U15329 (N_15329,N_14568,N_14718);
and U15330 (N_15330,N_14956,N_14481);
nand U15331 (N_15331,N_14626,N_14780);
nand U15332 (N_15332,N_14607,N_14947);
or U15333 (N_15333,N_14973,N_14967);
and U15334 (N_15334,N_14800,N_14546);
xor U15335 (N_15335,N_14458,N_14834);
nor U15336 (N_15336,N_14811,N_14495);
and U15337 (N_15337,N_14735,N_14723);
and U15338 (N_15338,N_14872,N_14544);
xor U15339 (N_15339,N_14917,N_14834);
or U15340 (N_15340,N_14922,N_14693);
xnor U15341 (N_15341,N_14470,N_14490);
nand U15342 (N_15342,N_14551,N_14879);
or U15343 (N_15343,N_14412,N_14595);
nand U15344 (N_15344,N_14658,N_14971);
or U15345 (N_15345,N_14409,N_14874);
or U15346 (N_15346,N_14706,N_14956);
and U15347 (N_15347,N_14693,N_14506);
or U15348 (N_15348,N_14895,N_14563);
nand U15349 (N_15349,N_14853,N_14703);
xor U15350 (N_15350,N_14658,N_14771);
or U15351 (N_15351,N_14675,N_14672);
or U15352 (N_15352,N_14452,N_14580);
nand U15353 (N_15353,N_14829,N_14970);
xor U15354 (N_15354,N_14944,N_14881);
xor U15355 (N_15355,N_14924,N_14811);
nor U15356 (N_15356,N_14846,N_14638);
xor U15357 (N_15357,N_14480,N_14992);
nand U15358 (N_15358,N_14933,N_14466);
nand U15359 (N_15359,N_14686,N_14451);
nand U15360 (N_15360,N_14802,N_14569);
nand U15361 (N_15361,N_14823,N_14922);
xnor U15362 (N_15362,N_14672,N_14797);
xor U15363 (N_15363,N_14428,N_14757);
and U15364 (N_15364,N_14777,N_14969);
or U15365 (N_15365,N_14438,N_14414);
nand U15366 (N_15366,N_14619,N_14792);
nand U15367 (N_15367,N_14415,N_14459);
xnor U15368 (N_15368,N_14743,N_14760);
nor U15369 (N_15369,N_14999,N_14892);
nand U15370 (N_15370,N_14951,N_14839);
nor U15371 (N_15371,N_14771,N_14559);
xor U15372 (N_15372,N_14782,N_14663);
nand U15373 (N_15373,N_14463,N_14785);
or U15374 (N_15374,N_14518,N_14467);
nor U15375 (N_15375,N_14593,N_14435);
nand U15376 (N_15376,N_14665,N_14473);
nand U15377 (N_15377,N_14770,N_14474);
or U15378 (N_15378,N_14500,N_14914);
nand U15379 (N_15379,N_14789,N_14978);
or U15380 (N_15380,N_14800,N_14678);
xor U15381 (N_15381,N_14459,N_14730);
and U15382 (N_15382,N_14985,N_14459);
xnor U15383 (N_15383,N_14690,N_14626);
or U15384 (N_15384,N_14605,N_14852);
and U15385 (N_15385,N_14419,N_14631);
nand U15386 (N_15386,N_14681,N_14573);
or U15387 (N_15387,N_14674,N_14663);
xor U15388 (N_15388,N_14726,N_14445);
xor U15389 (N_15389,N_14691,N_14986);
or U15390 (N_15390,N_14865,N_14828);
xor U15391 (N_15391,N_14402,N_14892);
nor U15392 (N_15392,N_14553,N_14407);
and U15393 (N_15393,N_14801,N_14676);
nand U15394 (N_15394,N_14459,N_14634);
nor U15395 (N_15395,N_14475,N_14889);
nor U15396 (N_15396,N_14678,N_14693);
or U15397 (N_15397,N_14727,N_14629);
xnor U15398 (N_15398,N_14410,N_14495);
xor U15399 (N_15399,N_14825,N_14625);
and U15400 (N_15400,N_14788,N_14791);
nor U15401 (N_15401,N_14945,N_14937);
nor U15402 (N_15402,N_14931,N_14892);
xnor U15403 (N_15403,N_14487,N_14498);
and U15404 (N_15404,N_14519,N_14805);
nand U15405 (N_15405,N_14676,N_14811);
xnor U15406 (N_15406,N_14889,N_14735);
xor U15407 (N_15407,N_14497,N_14478);
nand U15408 (N_15408,N_14554,N_14853);
xor U15409 (N_15409,N_14816,N_14422);
nand U15410 (N_15410,N_14606,N_14904);
and U15411 (N_15411,N_14647,N_14998);
xor U15412 (N_15412,N_14662,N_14454);
xnor U15413 (N_15413,N_14747,N_14970);
nor U15414 (N_15414,N_14725,N_14971);
nand U15415 (N_15415,N_14805,N_14759);
nor U15416 (N_15416,N_14634,N_14818);
and U15417 (N_15417,N_14940,N_14681);
xor U15418 (N_15418,N_14468,N_14878);
and U15419 (N_15419,N_14897,N_14453);
nand U15420 (N_15420,N_14576,N_14824);
or U15421 (N_15421,N_14535,N_14872);
nand U15422 (N_15422,N_14589,N_14651);
nand U15423 (N_15423,N_14929,N_14995);
or U15424 (N_15424,N_14961,N_14437);
nand U15425 (N_15425,N_14876,N_14830);
nor U15426 (N_15426,N_14688,N_14558);
nor U15427 (N_15427,N_14877,N_14927);
nor U15428 (N_15428,N_14576,N_14625);
and U15429 (N_15429,N_14774,N_14708);
nor U15430 (N_15430,N_14638,N_14479);
nor U15431 (N_15431,N_14765,N_14836);
xor U15432 (N_15432,N_14681,N_14856);
nand U15433 (N_15433,N_14552,N_14970);
nor U15434 (N_15434,N_14553,N_14618);
or U15435 (N_15435,N_14442,N_14844);
nor U15436 (N_15436,N_14891,N_14578);
or U15437 (N_15437,N_14784,N_14543);
or U15438 (N_15438,N_14510,N_14732);
nand U15439 (N_15439,N_14866,N_14695);
nor U15440 (N_15440,N_14550,N_14892);
xor U15441 (N_15441,N_14497,N_14469);
xnor U15442 (N_15442,N_14913,N_14632);
nor U15443 (N_15443,N_14860,N_14549);
nor U15444 (N_15444,N_14784,N_14923);
xor U15445 (N_15445,N_14767,N_14811);
nor U15446 (N_15446,N_14455,N_14936);
or U15447 (N_15447,N_14440,N_14663);
nand U15448 (N_15448,N_14768,N_14672);
xnor U15449 (N_15449,N_14553,N_14829);
and U15450 (N_15450,N_14532,N_14622);
or U15451 (N_15451,N_14719,N_14477);
nand U15452 (N_15452,N_14812,N_14741);
xor U15453 (N_15453,N_14626,N_14792);
nand U15454 (N_15454,N_14600,N_14616);
nor U15455 (N_15455,N_14709,N_14926);
and U15456 (N_15456,N_14634,N_14800);
and U15457 (N_15457,N_14669,N_14752);
nor U15458 (N_15458,N_14839,N_14766);
nand U15459 (N_15459,N_14725,N_14570);
nand U15460 (N_15460,N_14444,N_14842);
xor U15461 (N_15461,N_14602,N_14455);
or U15462 (N_15462,N_14585,N_14573);
or U15463 (N_15463,N_14807,N_14617);
and U15464 (N_15464,N_14517,N_14867);
and U15465 (N_15465,N_14630,N_14940);
and U15466 (N_15466,N_14841,N_14951);
xor U15467 (N_15467,N_14592,N_14974);
nor U15468 (N_15468,N_14735,N_14524);
and U15469 (N_15469,N_14993,N_14685);
or U15470 (N_15470,N_14646,N_14950);
nor U15471 (N_15471,N_14529,N_14793);
or U15472 (N_15472,N_14414,N_14507);
nand U15473 (N_15473,N_14815,N_14934);
or U15474 (N_15474,N_14600,N_14480);
nand U15475 (N_15475,N_14573,N_14424);
and U15476 (N_15476,N_14812,N_14539);
or U15477 (N_15477,N_14432,N_14783);
nor U15478 (N_15478,N_14975,N_14652);
xnor U15479 (N_15479,N_14926,N_14496);
or U15480 (N_15480,N_14534,N_14400);
xor U15481 (N_15481,N_14842,N_14592);
nand U15482 (N_15482,N_14414,N_14516);
nand U15483 (N_15483,N_14924,N_14705);
or U15484 (N_15484,N_14544,N_14500);
or U15485 (N_15485,N_14757,N_14776);
nand U15486 (N_15486,N_14914,N_14612);
xnor U15487 (N_15487,N_14706,N_14451);
or U15488 (N_15488,N_14779,N_14879);
or U15489 (N_15489,N_14515,N_14942);
and U15490 (N_15490,N_14907,N_14861);
xor U15491 (N_15491,N_14449,N_14628);
nor U15492 (N_15492,N_14802,N_14771);
nand U15493 (N_15493,N_14924,N_14527);
and U15494 (N_15494,N_14983,N_14604);
and U15495 (N_15495,N_14580,N_14895);
nor U15496 (N_15496,N_14829,N_14793);
nand U15497 (N_15497,N_14552,N_14542);
or U15498 (N_15498,N_14630,N_14936);
xor U15499 (N_15499,N_14893,N_14497);
nor U15500 (N_15500,N_14509,N_14888);
and U15501 (N_15501,N_14842,N_14445);
or U15502 (N_15502,N_14422,N_14546);
and U15503 (N_15503,N_14869,N_14720);
or U15504 (N_15504,N_14477,N_14505);
and U15505 (N_15505,N_14496,N_14467);
xor U15506 (N_15506,N_14940,N_14720);
and U15507 (N_15507,N_14522,N_14774);
nand U15508 (N_15508,N_14646,N_14887);
xor U15509 (N_15509,N_14534,N_14438);
nand U15510 (N_15510,N_14842,N_14455);
or U15511 (N_15511,N_14532,N_14421);
nand U15512 (N_15512,N_14572,N_14506);
and U15513 (N_15513,N_14976,N_14791);
or U15514 (N_15514,N_14648,N_14926);
or U15515 (N_15515,N_14546,N_14526);
nor U15516 (N_15516,N_14619,N_14848);
or U15517 (N_15517,N_14786,N_14477);
and U15518 (N_15518,N_14639,N_14516);
or U15519 (N_15519,N_14546,N_14999);
nand U15520 (N_15520,N_14700,N_14442);
xnor U15521 (N_15521,N_14996,N_14619);
xor U15522 (N_15522,N_14652,N_14628);
and U15523 (N_15523,N_14779,N_14526);
and U15524 (N_15524,N_14823,N_14633);
and U15525 (N_15525,N_14915,N_14412);
nand U15526 (N_15526,N_14545,N_14749);
or U15527 (N_15527,N_14730,N_14524);
xnor U15528 (N_15528,N_14647,N_14491);
xor U15529 (N_15529,N_14633,N_14466);
nor U15530 (N_15530,N_14604,N_14513);
xnor U15531 (N_15531,N_14989,N_14708);
nand U15532 (N_15532,N_14642,N_14637);
or U15533 (N_15533,N_14739,N_14688);
xor U15534 (N_15534,N_14470,N_14451);
or U15535 (N_15535,N_14790,N_14500);
and U15536 (N_15536,N_14733,N_14847);
xnor U15537 (N_15537,N_14809,N_14930);
nand U15538 (N_15538,N_14556,N_14831);
nand U15539 (N_15539,N_14844,N_14659);
nand U15540 (N_15540,N_14784,N_14546);
nand U15541 (N_15541,N_14906,N_14734);
nor U15542 (N_15542,N_14882,N_14963);
nand U15543 (N_15543,N_14945,N_14908);
xor U15544 (N_15544,N_14612,N_14902);
and U15545 (N_15545,N_14899,N_14520);
xor U15546 (N_15546,N_14412,N_14931);
nor U15547 (N_15547,N_14464,N_14825);
and U15548 (N_15548,N_14841,N_14420);
nor U15549 (N_15549,N_14515,N_14966);
nor U15550 (N_15550,N_14692,N_14814);
xor U15551 (N_15551,N_14885,N_14456);
and U15552 (N_15552,N_14446,N_14943);
or U15553 (N_15553,N_14875,N_14970);
nand U15554 (N_15554,N_14927,N_14816);
and U15555 (N_15555,N_14645,N_14728);
and U15556 (N_15556,N_14495,N_14730);
xor U15557 (N_15557,N_14703,N_14502);
or U15558 (N_15558,N_14447,N_14853);
and U15559 (N_15559,N_14834,N_14944);
or U15560 (N_15560,N_14685,N_14495);
xor U15561 (N_15561,N_14790,N_14467);
and U15562 (N_15562,N_14520,N_14668);
or U15563 (N_15563,N_14941,N_14721);
nor U15564 (N_15564,N_14920,N_14611);
nand U15565 (N_15565,N_14519,N_14473);
xnor U15566 (N_15566,N_14440,N_14520);
nor U15567 (N_15567,N_14960,N_14945);
nor U15568 (N_15568,N_14785,N_14952);
nand U15569 (N_15569,N_14589,N_14826);
nand U15570 (N_15570,N_14889,N_14821);
or U15571 (N_15571,N_14950,N_14865);
xnor U15572 (N_15572,N_14903,N_14848);
nand U15573 (N_15573,N_14436,N_14964);
nand U15574 (N_15574,N_14982,N_14590);
nand U15575 (N_15575,N_14798,N_14641);
or U15576 (N_15576,N_14621,N_14609);
nand U15577 (N_15577,N_14721,N_14715);
xor U15578 (N_15578,N_14919,N_14512);
nand U15579 (N_15579,N_14976,N_14631);
xor U15580 (N_15580,N_14594,N_14832);
xor U15581 (N_15581,N_14456,N_14585);
nor U15582 (N_15582,N_14524,N_14959);
nor U15583 (N_15583,N_14872,N_14905);
and U15584 (N_15584,N_14895,N_14618);
and U15585 (N_15585,N_14872,N_14545);
or U15586 (N_15586,N_14438,N_14720);
nand U15587 (N_15587,N_14636,N_14443);
nor U15588 (N_15588,N_14859,N_14436);
or U15589 (N_15589,N_14530,N_14828);
nor U15590 (N_15590,N_14764,N_14675);
and U15591 (N_15591,N_14912,N_14874);
nand U15592 (N_15592,N_14923,N_14593);
or U15593 (N_15593,N_14568,N_14624);
and U15594 (N_15594,N_14523,N_14448);
nor U15595 (N_15595,N_14867,N_14707);
or U15596 (N_15596,N_14691,N_14774);
xor U15597 (N_15597,N_14952,N_14730);
nand U15598 (N_15598,N_14474,N_14954);
and U15599 (N_15599,N_14790,N_14731);
nand U15600 (N_15600,N_15367,N_15317);
xnor U15601 (N_15601,N_15325,N_15228);
or U15602 (N_15602,N_15418,N_15191);
or U15603 (N_15603,N_15199,N_15296);
or U15604 (N_15604,N_15369,N_15545);
or U15605 (N_15605,N_15587,N_15091);
xor U15606 (N_15606,N_15313,N_15157);
or U15607 (N_15607,N_15424,N_15388);
nor U15608 (N_15608,N_15043,N_15022);
and U15609 (N_15609,N_15516,N_15336);
nor U15610 (N_15610,N_15229,N_15509);
xor U15611 (N_15611,N_15000,N_15289);
nand U15612 (N_15612,N_15205,N_15027);
or U15613 (N_15613,N_15494,N_15005);
or U15614 (N_15614,N_15534,N_15370);
or U15615 (N_15615,N_15459,N_15287);
nand U15616 (N_15616,N_15458,N_15446);
nor U15617 (N_15617,N_15498,N_15359);
nor U15618 (N_15618,N_15444,N_15206);
nor U15619 (N_15619,N_15442,N_15072);
or U15620 (N_15620,N_15169,N_15365);
nor U15621 (N_15621,N_15084,N_15501);
and U15622 (N_15622,N_15538,N_15330);
and U15623 (N_15623,N_15475,N_15593);
xor U15624 (N_15624,N_15343,N_15310);
nand U15625 (N_15625,N_15150,N_15140);
and U15626 (N_15626,N_15390,N_15009);
nor U15627 (N_15627,N_15536,N_15318);
or U15628 (N_15628,N_15300,N_15161);
or U15629 (N_15629,N_15360,N_15292);
xor U15630 (N_15630,N_15361,N_15294);
nor U15631 (N_15631,N_15013,N_15048);
and U15632 (N_15632,N_15101,N_15282);
or U15633 (N_15633,N_15414,N_15568);
and U15634 (N_15634,N_15519,N_15505);
xor U15635 (N_15635,N_15156,N_15577);
or U15636 (N_15636,N_15448,N_15065);
nand U15637 (N_15637,N_15098,N_15113);
and U15638 (N_15638,N_15123,N_15341);
or U15639 (N_15639,N_15306,N_15086);
or U15640 (N_15640,N_15307,N_15503);
and U15641 (N_15641,N_15014,N_15015);
xnor U15642 (N_15642,N_15346,N_15125);
and U15643 (N_15643,N_15426,N_15462);
nor U15644 (N_15644,N_15398,N_15399);
nand U15645 (N_15645,N_15429,N_15447);
and U15646 (N_15646,N_15251,N_15449);
and U15647 (N_15647,N_15511,N_15030);
or U15648 (N_15648,N_15338,N_15456);
nand U15649 (N_15649,N_15490,N_15514);
xor U15650 (N_15650,N_15384,N_15196);
nor U15651 (N_15651,N_15059,N_15147);
xnor U15652 (N_15652,N_15077,N_15097);
nor U15653 (N_15653,N_15152,N_15526);
or U15654 (N_15654,N_15576,N_15183);
or U15655 (N_15655,N_15172,N_15268);
or U15656 (N_15656,N_15102,N_15128);
nand U15657 (N_15657,N_15419,N_15401);
and U15658 (N_15658,N_15495,N_15181);
xor U15659 (N_15659,N_15254,N_15242);
or U15660 (N_15660,N_15345,N_15131);
or U15661 (N_15661,N_15510,N_15561);
nor U15662 (N_15662,N_15589,N_15432);
xor U15663 (N_15663,N_15539,N_15579);
xor U15664 (N_15664,N_15473,N_15303);
and U15665 (N_15665,N_15255,N_15542);
xnor U15666 (N_15666,N_15057,N_15350);
and U15667 (N_15667,N_15588,N_15258);
or U15668 (N_15668,N_15454,N_15198);
or U15669 (N_15669,N_15068,N_15468);
nand U15670 (N_15670,N_15524,N_15087);
and U15671 (N_15671,N_15415,N_15164);
nor U15672 (N_15672,N_15078,N_15315);
and U15673 (N_15673,N_15261,N_15063);
xnor U15674 (N_15674,N_15544,N_15266);
or U15675 (N_15675,N_15550,N_15331);
xor U15676 (N_15676,N_15353,N_15054);
nor U15677 (N_15677,N_15435,N_15582);
nor U15678 (N_15678,N_15194,N_15354);
nor U15679 (N_15679,N_15484,N_15549);
xor U15680 (N_15680,N_15061,N_15070);
or U15681 (N_15681,N_15520,N_15130);
nand U15682 (N_15682,N_15244,N_15402);
or U15683 (N_15683,N_15175,N_15221);
nand U15684 (N_15684,N_15437,N_15489);
and U15685 (N_15685,N_15339,N_15224);
nor U15686 (N_15686,N_15178,N_15347);
and U15687 (N_15687,N_15377,N_15075);
nand U15688 (N_15688,N_15197,N_15276);
nor U15689 (N_15689,N_15174,N_15450);
nor U15690 (N_15690,N_15136,N_15149);
xnor U15691 (N_15691,N_15485,N_15004);
and U15692 (N_15692,N_15522,N_15094);
nand U15693 (N_15693,N_15480,N_15222);
nor U15694 (N_15694,N_15529,N_15283);
nand U15695 (N_15695,N_15425,N_15492);
and U15696 (N_15696,N_15190,N_15141);
nand U15697 (N_15697,N_15559,N_15428);
or U15698 (N_15698,N_15278,N_15430);
and U15699 (N_15699,N_15036,N_15240);
nor U15700 (N_15700,N_15465,N_15556);
or U15701 (N_15701,N_15045,N_15560);
nor U15702 (N_15702,N_15396,N_15403);
xor U15703 (N_15703,N_15453,N_15200);
xor U15704 (N_15704,N_15460,N_15177);
nand U15705 (N_15705,N_15585,N_15400);
nand U15706 (N_15706,N_15351,N_15275);
nor U15707 (N_15707,N_15262,N_15575);
and U15708 (N_15708,N_15211,N_15017);
nor U15709 (N_15709,N_15451,N_15590);
and U15710 (N_15710,N_15231,N_15008);
nor U15711 (N_15711,N_15117,N_15021);
nor U15712 (N_15712,N_15387,N_15290);
nand U15713 (N_15713,N_15193,N_15328);
xnor U15714 (N_15714,N_15570,N_15090);
and U15715 (N_15715,N_15227,N_15481);
xnor U15716 (N_15716,N_15518,N_15154);
xnor U15717 (N_15717,N_15108,N_15105);
or U15718 (N_15718,N_15483,N_15597);
xor U15719 (N_15719,N_15270,N_15515);
xor U15720 (N_15720,N_15280,N_15376);
and U15721 (N_15721,N_15056,N_15566);
or U15722 (N_15722,N_15024,N_15368);
xnor U15723 (N_15723,N_15364,N_15411);
nor U15724 (N_15724,N_15394,N_15184);
or U15725 (N_15725,N_15159,N_15405);
and U15726 (N_15726,N_15257,N_15243);
nand U15727 (N_15727,N_15288,N_15037);
or U15728 (N_15728,N_15253,N_15120);
nand U15729 (N_15729,N_15115,N_15212);
and U15730 (N_15730,N_15019,N_15540);
or U15731 (N_15731,N_15069,N_15011);
nand U15732 (N_15732,N_15179,N_15274);
nand U15733 (N_15733,N_15273,N_15104);
and U15734 (N_15734,N_15391,N_15547);
xor U15735 (N_15735,N_15007,N_15295);
and U15736 (N_15736,N_15323,N_15153);
nand U15737 (N_15737,N_15578,N_15018);
xor U15738 (N_15738,N_15441,N_15472);
nor U15739 (N_15739,N_15423,N_15440);
and U15740 (N_15740,N_15305,N_15281);
nor U15741 (N_15741,N_15277,N_15041);
nor U15742 (N_15742,N_15286,N_15372);
nand U15743 (N_15743,N_15537,N_15562);
or U15744 (N_15744,N_15111,N_15026);
or U15745 (N_15745,N_15210,N_15312);
nand U15746 (N_15746,N_15223,N_15298);
nor U15747 (N_15747,N_15245,N_15554);
and U15748 (N_15748,N_15049,N_15548);
nor U15749 (N_15749,N_15046,N_15050);
and U15750 (N_15750,N_15192,N_15137);
xnor U15751 (N_15751,N_15010,N_15469);
nor U15752 (N_15752,N_15217,N_15003);
nand U15753 (N_15753,N_15521,N_15185);
nor U15754 (N_15754,N_15256,N_15076);
and U15755 (N_15755,N_15565,N_15166);
and U15756 (N_15756,N_15092,N_15356);
xnor U15757 (N_15757,N_15215,N_15119);
xor U15758 (N_15758,N_15241,N_15584);
nand U15759 (N_15759,N_15219,N_15297);
or U15760 (N_15760,N_15074,N_15265);
nor U15761 (N_15761,N_15332,N_15436);
or U15762 (N_15762,N_15006,N_15071);
nor U15763 (N_15763,N_15116,N_15064);
or U15764 (N_15764,N_15246,N_15082);
xnor U15765 (N_15765,N_15249,N_15322);
and U15766 (N_15766,N_15445,N_15513);
and U15767 (N_15767,N_15416,N_15103);
nand U15768 (N_15768,N_15118,N_15248);
xnor U15769 (N_15769,N_15263,N_15586);
xnor U15770 (N_15770,N_15126,N_15385);
and U15771 (N_15771,N_15525,N_15467);
and U15772 (N_15772,N_15477,N_15574);
or U15773 (N_15773,N_15327,N_15032);
nand U15774 (N_15774,N_15171,N_15496);
nor U15775 (N_15775,N_15357,N_15572);
and U15776 (N_15776,N_15393,N_15476);
nand U15777 (N_15777,N_15148,N_15583);
nor U15778 (N_15778,N_15500,N_15060);
nand U15779 (N_15779,N_15269,N_15417);
xnor U15780 (N_15780,N_15299,N_15382);
and U15781 (N_15781,N_15051,N_15052);
xor U15782 (N_15782,N_15029,N_15085);
xor U15783 (N_15783,N_15413,N_15238);
nor U15784 (N_15784,N_15404,N_15038);
nand U15785 (N_15785,N_15320,N_15284);
and U15786 (N_15786,N_15234,N_15134);
xnor U15787 (N_15787,N_15099,N_15167);
nor U15788 (N_15788,N_15095,N_15506);
xor U15789 (N_15789,N_15132,N_15230);
nand U15790 (N_15790,N_15507,N_15466);
xor U15791 (N_15791,N_15035,N_15016);
nand U15792 (N_15792,N_15067,N_15247);
or U15793 (N_15793,N_15220,N_15352);
nand U15794 (N_15794,N_15168,N_15378);
nand U15795 (N_15795,N_15573,N_15395);
or U15796 (N_15796,N_15478,N_15264);
xor U15797 (N_15797,N_15553,N_15366);
nor U15798 (N_15798,N_15319,N_15517);
xor U15799 (N_15799,N_15371,N_15493);
or U15800 (N_15800,N_15225,N_15055);
nor U15801 (N_15801,N_15488,N_15409);
nor U15802 (N_15802,N_15023,N_15564);
nand U15803 (N_15803,N_15552,N_15144);
nand U15804 (N_15804,N_15457,N_15421);
xor U15805 (N_15805,N_15358,N_15081);
nor U15806 (N_15806,N_15093,N_15592);
nand U15807 (N_15807,N_15129,N_15527);
and U15808 (N_15808,N_15233,N_15226);
nand U15809 (N_15809,N_15058,N_15504);
nand U15810 (N_15810,N_15541,N_15434);
and U15811 (N_15811,N_15362,N_15302);
xnor U15812 (N_15812,N_15232,N_15311);
nor U15813 (N_15813,N_15182,N_15380);
nor U15814 (N_15814,N_15237,N_15109);
nor U15815 (N_15815,N_15165,N_15598);
nand U15816 (N_15816,N_15452,N_15455);
and U15817 (N_15817,N_15073,N_15363);
nor U15818 (N_15818,N_15397,N_15107);
and U15819 (N_15819,N_15463,N_15293);
and U15820 (N_15820,N_15209,N_15112);
nand U15821 (N_15821,N_15508,N_15145);
xnor U15822 (N_15822,N_15591,N_15124);
nand U15823 (N_15823,N_15100,N_15188);
xnor U15824 (N_15824,N_15250,N_15431);
xnor U15825 (N_15825,N_15427,N_15146);
xnor U15826 (N_15826,N_15340,N_15208);
or U15827 (N_15827,N_15502,N_15532);
or U15828 (N_15828,N_15163,N_15180);
nor U15829 (N_15829,N_15580,N_15407);
or U15830 (N_15830,N_15487,N_15158);
nor U15831 (N_15831,N_15474,N_15213);
xnor U15832 (N_15832,N_15260,N_15321);
xor U15833 (N_15833,N_15558,N_15133);
nand U15834 (N_15834,N_15088,N_15412);
nor U15835 (N_15835,N_15309,N_15523);
xnor U15836 (N_15836,N_15408,N_15497);
xnor U15837 (N_15837,N_15594,N_15551);
nor U15838 (N_15838,N_15479,N_15595);
xor U15839 (N_15839,N_15034,N_15344);
nand U15840 (N_15840,N_15203,N_15151);
nor U15841 (N_15841,N_15002,N_15433);
or U15842 (N_15842,N_15316,N_15047);
or U15843 (N_15843,N_15216,N_15122);
nor U15844 (N_15844,N_15599,N_15569);
or U15845 (N_15845,N_15042,N_15271);
nand U15846 (N_15846,N_15439,N_15491);
or U15847 (N_15847,N_15044,N_15355);
or U15848 (N_15848,N_15186,N_15571);
nor U15849 (N_15849,N_15020,N_15386);
xnor U15850 (N_15850,N_15001,N_15348);
nand U15851 (N_15851,N_15555,N_15349);
nand U15852 (N_15852,N_15062,N_15443);
or U15853 (N_15853,N_15333,N_15272);
xnor U15854 (N_15854,N_15110,N_15025);
nor U15855 (N_15855,N_15499,N_15486);
nor U15856 (N_15856,N_15471,N_15202);
xor U15857 (N_15857,N_15581,N_15033);
nand U15858 (N_15858,N_15083,N_15531);
or U15859 (N_15859,N_15135,N_15383);
and U15860 (N_15860,N_15543,N_15329);
xnor U15861 (N_15861,N_15546,N_15381);
and U15862 (N_15862,N_15201,N_15374);
xor U15863 (N_15863,N_15334,N_15482);
or U15864 (N_15864,N_15337,N_15127);
nand U15865 (N_15865,N_15301,N_15342);
or U15866 (N_15866,N_15239,N_15031);
or U15867 (N_15867,N_15285,N_15187);
or U15868 (N_15868,N_15563,N_15533);
or U15869 (N_15869,N_15389,N_15039);
nor U15870 (N_15870,N_15096,N_15138);
nor U15871 (N_15871,N_15173,N_15596);
nor U15872 (N_15872,N_15304,N_15528);
nand U15873 (N_15873,N_15121,N_15259);
xor U15874 (N_15874,N_15160,N_15079);
or U15875 (N_15875,N_15512,N_15139);
nand U15876 (N_15876,N_15235,N_15207);
and U15877 (N_15877,N_15066,N_15218);
nor U15878 (N_15878,N_15214,N_15012);
nor U15879 (N_15879,N_15176,N_15308);
or U15880 (N_15880,N_15326,N_15530);
xor U15881 (N_15881,N_15314,N_15470);
nand U15882 (N_15882,N_15279,N_15162);
or U15883 (N_15883,N_15028,N_15379);
nor U15884 (N_15884,N_15438,N_15252);
or U15885 (N_15885,N_15189,N_15291);
or U15886 (N_15886,N_15114,N_15089);
or U15887 (N_15887,N_15267,N_15143);
and U15888 (N_15888,N_15406,N_15461);
or U15889 (N_15889,N_15236,N_15324);
and U15890 (N_15890,N_15040,N_15557);
and U15891 (N_15891,N_15335,N_15375);
and U15892 (N_15892,N_15106,N_15410);
nor U15893 (N_15893,N_15535,N_15373);
or U15894 (N_15894,N_15142,N_15195);
nor U15895 (N_15895,N_15170,N_15422);
or U15896 (N_15896,N_15567,N_15080);
nor U15897 (N_15897,N_15155,N_15392);
and U15898 (N_15898,N_15464,N_15420);
or U15899 (N_15899,N_15204,N_15053);
xor U15900 (N_15900,N_15196,N_15124);
xnor U15901 (N_15901,N_15219,N_15352);
nor U15902 (N_15902,N_15160,N_15025);
nand U15903 (N_15903,N_15278,N_15045);
or U15904 (N_15904,N_15405,N_15329);
or U15905 (N_15905,N_15188,N_15081);
and U15906 (N_15906,N_15069,N_15337);
xnor U15907 (N_15907,N_15088,N_15263);
nand U15908 (N_15908,N_15148,N_15578);
nor U15909 (N_15909,N_15266,N_15047);
nor U15910 (N_15910,N_15570,N_15457);
nor U15911 (N_15911,N_15362,N_15415);
nand U15912 (N_15912,N_15138,N_15560);
nor U15913 (N_15913,N_15475,N_15163);
or U15914 (N_15914,N_15431,N_15194);
and U15915 (N_15915,N_15451,N_15444);
and U15916 (N_15916,N_15034,N_15071);
nand U15917 (N_15917,N_15267,N_15531);
nor U15918 (N_15918,N_15020,N_15049);
nand U15919 (N_15919,N_15517,N_15516);
xnor U15920 (N_15920,N_15197,N_15000);
or U15921 (N_15921,N_15234,N_15419);
and U15922 (N_15922,N_15433,N_15250);
or U15923 (N_15923,N_15232,N_15354);
nand U15924 (N_15924,N_15520,N_15148);
nor U15925 (N_15925,N_15121,N_15145);
xor U15926 (N_15926,N_15196,N_15449);
or U15927 (N_15927,N_15255,N_15229);
or U15928 (N_15928,N_15406,N_15009);
xor U15929 (N_15929,N_15480,N_15251);
nor U15930 (N_15930,N_15395,N_15334);
xnor U15931 (N_15931,N_15425,N_15422);
nand U15932 (N_15932,N_15522,N_15150);
nor U15933 (N_15933,N_15278,N_15030);
xor U15934 (N_15934,N_15447,N_15504);
and U15935 (N_15935,N_15382,N_15401);
nor U15936 (N_15936,N_15509,N_15168);
and U15937 (N_15937,N_15545,N_15301);
and U15938 (N_15938,N_15563,N_15448);
nand U15939 (N_15939,N_15298,N_15397);
nand U15940 (N_15940,N_15057,N_15385);
nand U15941 (N_15941,N_15120,N_15484);
nand U15942 (N_15942,N_15175,N_15016);
nor U15943 (N_15943,N_15441,N_15079);
nand U15944 (N_15944,N_15563,N_15247);
or U15945 (N_15945,N_15178,N_15507);
nand U15946 (N_15946,N_15373,N_15498);
xor U15947 (N_15947,N_15064,N_15246);
nor U15948 (N_15948,N_15071,N_15395);
or U15949 (N_15949,N_15585,N_15011);
or U15950 (N_15950,N_15047,N_15282);
nor U15951 (N_15951,N_15277,N_15447);
xor U15952 (N_15952,N_15596,N_15302);
or U15953 (N_15953,N_15024,N_15406);
xnor U15954 (N_15954,N_15236,N_15396);
xnor U15955 (N_15955,N_15330,N_15364);
nand U15956 (N_15956,N_15224,N_15053);
xnor U15957 (N_15957,N_15297,N_15476);
xnor U15958 (N_15958,N_15516,N_15423);
xor U15959 (N_15959,N_15019,N_15130);
and U15960 (N_15960,N_15499,N_15439);
xnor U15961 (N_15961,N_15077,N_15058);
and U15962 (N_15962,N_15571,N_15372);
xnor U15963 (N_15963,N_15113,N_15273);
nor U15964 (N_15964,N_15153,N_15433);
xnor U15965 (N_15965,N_15235,N_15370);
nor U15966 (N_15966,N_15448,N_15455);
or U15967 (N_15967,N_15292,N_15230);
or U15968 (N_15968,N_15313,N_15533);
or U15969 (N_15969,N_15454,N_15116);
nor U15970 (N_15970,N_15279,N_15314);
nand U15971 (N_15971,N_15007,N_15037);
nand U15972 (N_15972,N_15206,N_15020);
xnor U15973 (N_15973,N_15359,N_15514);
nor U15974 (N_15974,N_15042,N_15132);
nor U15975 (N_15975,N_15006,N_15408);
and U15976 (N_15976,N_15266,N_15283);
nor U15977 (N_15977,N_15335,N_15523);
and U15978 (N_15978,N_15587,N_15358);
or U15979 (N_15979,N_15398,N_15505);
xor U15980 (N_15980,N_15538,N_15582);
xor U15981 (N_15981,N_15577,N_15276);
nor U15982 (N_15982,N_15444,N_15268);
or U15983 (N_15983,N_15483,N_15560);
or U15984 (N_15984,N_15156,N_15221);
or U15985 (N_15985,N_15597,N_15408);
or U15986 (N_15986,N_15504,N_15035);
and U15987 (N_15987,N_15233,N_15120);
xnor U15988 (N_15988,N_15391,N_15393);
or U15989 (N_15989,N_15588,N_15474);
xor U15990 (N_15990,N_15034,N_15284);
and U15991 (N_15991,N_15532,N_15128);
nand U15992 (N_15992,N_15406,N_15306);
or U15993 (N_15993,N_15505,N_15222);
nor U15994 (N_15994,N_15400,N_15560);
or U15995 (N_15995,N_15186,N_15356);
or U15996 (N_15996,N_15325,N_15161);
xnor U15997 (N_15997,N_15321,N_15265);
nand U15998 (N_15998,N_15331,N_15225);
nor U15999 (N_15999,N_15285,N_15055);
nor U16000 (N_16000,N_15595,N_15175);
nand U16001 (N_16001,N_15215,N_15518);
and U16002 (N_16002,N_15355,N_15175);
nor U16003 (N_16003,N_15485,N_15238);
and U16004 (N_16004,N_15444,N_15323);
xor U16005 (N_16005,N_15259,N_15187);
xnor U16006 (N_16006,N_15272,N_15229);
or U16007 (N_16007,N_15014,N_15087);
or U16008 (N_16008,N_15198,N_15217);
or U16009 (N_16009,N_15381,N_15309);
or U16010 (N_16010,N_15064,N_15120);
nor U16011 (N_16011,N_15408,N_15406);
xor U16012 (N_16012,N_15331,N_15251);
xor U16013 (N_16013,N_15258,N_15443);
nand U16014 (N_16014,N_15486,N_15237);
and U16015 (N_16015,N_15012,N_15366);
or U16016 (N_16016,N_15463,N_15575);
nor U16017 (N_16017,N_15080,N_15570);
or U16018 (N_16018,N_15460,N_15367);
nand U16019 (N_16019,N_15356,N_15034);
nor U16020 (N_16020,N_15346,N_15099);
or U16021 (N_16021,N_15154,N_15287);
and U16022 (N_16022,N_15143,N_15109);
or U16023 (N_16023,N_15183,N_15148);
xnor U16024 (N_16024,N_15448,N_15181);
or U16025 (N_16025,N_15302,N_15323);
nor U16026 (N_16026,N_15153,N_15592);
or U16027 (N_16027,N_15088,N_15440);
or U16028 (N_16028,N_15256,N_15107);
and U16029 (N_16029,N_15035,N_15499);
nor U16030 (N_16030,N_15353,N_15455);
and U16031 (N_16031,N_15080,N_15266);
nor U16032 (N_16032,N_15401,N_15345);
and U16033 (N_16033,N_15331,N_15139);
nand U16034 (N_16034,N_15401,N_15368);
nand U16035 (N_16035,N_15139,N_15551);
and U16036 (N_16036,N_15252,N_15420);
xnor U16037 (N_16037,N_15228,N_15217);
xor U16038 (N_16038,N_15179,N_15352);
or U16039 (N_16039,N_15077,N_15366);
and U16040 (N_16040,N_15338,N_15314);
xor U16041 (N_16041,N_15526,N_15599);
nand U16042 (N_16042,N_15219,N_15235);
xnor U16043 (N_16043,N_15479,N_15024);
nand U16044 (N_16044,N_15031,N_15417);
nor U16045 (N_16045,N_15067,N_15235);
nor U16046 (N_16046,N_15470,N_15054);
nor U16047 (N_16047,N_15081,N_15361);
nor U16048 (N_16048,N_15251,N_15298);
nor U16049 (N_16049,N_15574,N_15214);
nor U16050 (N_16050,N_15521,N_15008);
or U16051 (N_16051,N_15334,N_15254);
nor U16052 (N_16052,N_15428,N_15259);
nor U16053 (N_16053,N_15154,N_15478);
nor U16054 (N_16054,N_15099,N_15317);
nor U16055 (N_16055,N_15559,N_15591);
xor U16056 (N_16056,N_15214,N_15217);
nand U16057 (N_16057,N_15441,N_15322);
and U16058 (N_16058,N_15513,N_15175);
xor U16059 (N_16059,N_15312,N_15417);
nor U16060 (N_16060,N_15463,N_15020);
xor U16061 (N_16061,N_15254,N_15199);
nor U16062 (N_16062,N_15145,N_15348);
nand U16063 (N_16063,N_15497,N_15073);
and U16064 (N_16064,N_15109,N_15096);
and U16065 (N_16065,N_15201,N_15582);
nor U16066 (N_16066,N_15192,N_15493);
nand U16067 (N_16067,N_15113,N_15214);
or U16068 (N_16068,N_15152,N_15194);
or U16069 (N_16069,N_15556,N_15599);
nand U16070 (N_16070,N_15003,N_15450);
or U16071 (N_16071,N_15058,N_15477);
nor U16072 (N_16072,N_15561,N_15364);
nand U16073 (N_16073,N_15530,N_15132);
or U16074 (N_16074,N_15078,N_15174);
nand U16075 (N_16075,N_15299,N_15000);
or U16076 (N_16076,N_15389,N_15109);
xnor U16077 (N_16077,N_15122,N_15045);
xnor U16078 (N_16078,N_15057,N_15507);
xnor U16079 (N_16079,N_15260,N_15243);
xor U16080 (N_16080,N_15329,N_15060);
nor U16081 (N_16081,N_15016,N_15369);
nor U16082 (N_16082,N_15562,N_15016);
or U16083 (N_16083,N_15434,N_15014);
xor U16084 (N_16084,N_15502,N_15145);
and U16085 (N_16085,N_15065,N_15152);
nand U16086 (N_16086,N_15037,N_15407);
or U16087 (N_16087,N_15319,N_15132);
and U16088 (N_16088,N_15344,N_15576);
nand U16089 (N_16089,N_15429,N_15404);
or U16090 (N_16090,N_15220,N_15226);
xnor U16091 (N_16091,N_15284,N_15247);
xor U16092 (N_16092,N_15117,N_15193);
nor U16093 (N_16093,N_15257,N_15526);
nor U16094 (N_16094,N_15125,N_15270);
nand U16095 (N_16095,N_15567,N_15101);
and U16096 (N_16096,N_15253,N_15508);
and U16097 (N_16097,N_15345,N_15506);
nor U16098 (N_16098,N_15476,N_15511);
and U16099 (N_16099,N_15061,N_15109);
xnor U16100 (N_16100,N_15540,N_15568);
nor U16101 (N_16101,N_15244,N_15055);
xor U16102 (N_16102,N_15119,N_15181);
and U16103 (N_16103,N_15426,N_15227);
nand U16104 (N_16104,N_15329,N_15583);
nand U16105 (N_16105,N_15530,N_15508);
nand U16106 (N_16106,N_15351,N_15401);
xor U16107 (N_16107,N_15271,N_15166);
and U16108 (N_16108,N_15240,N_15372);
and U16109 (N_16109,N_15038,N_15023);
nor U16110 (N_16110,N_15360,N_15546);
and U16111 (N_16111,N_15128,N_15103);
xor U16112 (N_16112,N_15193,N_15308);
or U16113 (N_16113,N_15558,N_15116);
nor U16114 (N_16114,N_15427,N_15441);
nand U16115 (N_16115,N_15312,N_15187);
nand U16116 (N_16116,N_15555,N_15592);
nor U16117 (N_16117,N_15528,N_15427);
xnor U16118 (N_16118,N_15001,N_15273);
nor U16119 (N_16119,N_15402,N_15114);
xor U16120 (N_16120,N_15279,N_15125);
or U16121 (N_16121,N_15228,N_15270);
and U16122 (N_16122,N_15585,N_15290);
nor U16123 (N_16123,N_15329,N_15362);
or U16124 (N_16124,N_15328,N_15322);
or U16125 (N_16125,N_15204,N_15058);
or U16126 (N_16126,N_15511,N_15537);
nand U16127 (N_16127,N_15575,N_15332);
xnor U16128 (N_16128,N_15127,N_15249);
and U16129 (N_16129,N_15224,N_15225);
nor U16130 (N_16130,N_15326,N_15068);
xor U16131 (N_16131,N_15101,N_15109);
xor U16132 (N_16132,N_15376,N_15174);
nor U16133 (N_16133,N_15524,N_15513);
xor U16134 (N_16134,N_15024,N_15187);
or U16135 (N_16135,N_15067,N_15081);
xnor U16136 (N_16136,N_15400,N_15561);
xor U16137 (N_16137,N_15080,N_15572);
and U16138 (N_16138,N_15175,N_15458);
or U16139 (N_16139,N_15545,N_15582);
or U16140 (N_16140,N_15583,N_15479);
nand U16141 (N_16141,N_15349,N_15338);
xor U16142 (N_16142,N_15430,N_15464);
or U16143 (N_16143,N_15190,N_15083);
and U16144 (N_16144,N_15410,N_15464);
nor U16145 (N_16145,N_15270,N_15453);
or U16146 (N_16146,N_15147,N_15578);
or U16147 (N_16147,N_15366,N_15075);
and U16148 (N_16148,N_15351,N_15284);
and U16149 (N_16149,N_15211,N_15498);
or U16150 (N_16150,N_15186,N_15515);
nand U16151 (N_16151,N_15004,N_15225);
or U16152 (N_16152,N_15106,N_15315);
xor U16153 (N_16153,N_15398,N_15055);
and U16154 (N_16154,N_15153,N_15185);
or U16155 (N_16155,N_15163,N_15040);
nand U16156 (N_16156,N_15032,N_15363);
and U16157 (N_16157,N_15018,N_15408);
xor U16158 (N_16158,N_15501,N_15573);
nor U16159 (N_16159,N_15180,N_15196);
or U16160 (N_16160,N_15537,N_15174);
nor U16161 (N_16161,N_15237,N_15135);
nand U16162 (N_16162,N_15063,N_15379);
nand U16163 (N_16163,N_15533,N_15290);
xnor U16164 (N_16164,N_15110,N_15441);
nor U16165 (N_16165,N_15595,N_15150);
nor U16166 (N_16166,N_15077,N_15585);
and U16167 (N_16167,N_15230,N_15574);
xnor U16168 (N_16168,N_15237,N_15091);
xnor U16169 (N_16169,N_15460,N_15278);
nor U16170 (N_16170,N_15063,N_15068);
and U16171 (N_16171,N_15184,N_15019);
nand U16172 (N_16172,N_15297,N_15563);
nand U16173 (N_16173,N_15595,N_15519);
nor U16174 (N_16174,N_15431,N_15383);
nand U16175 (N_16175,N_15230,N_15387);
xor U16176 (N_16176,N_15292,N_15356);
and U16177 (N_16177,N_15017,N_15158);
nand U16178 (N_16178,N_15386,N_15327);
or U16179 (N_16179,N_15194,N_15523);
nand U16180 (N_16180,N_15403,N_15437);
xnor U16181 (N_16181,N_15261,N_15330);
xnor U16182 (N_16182,N_15399,N_15517);
nand U16183 (N_16183,N_15164,N_15351);
nor U16184 (N_16184,N_15170,N_15098);
or U16185 (N_16185,N_15111,N_15198);
xnor U16186 (N_16186,N_15513,N_15542);
and U16187 (N_16187,N_15201,N_15552);
xnor U16188 (N_16188,N_15280,N_15096);
xnor U16189 (N_16189,N_15259,N_15147);
nor U16190 (N_16190,N_15220,N_15574);
and U16191 (N_16191,N_15247,N_15066);
or U16192 (N_16192,N_15149,N_15584);
nand U16193 (N_16193,N_15127,N_15017);
and U16194 (N_16194,N_15126,N_15454);
or U16195 (N_16195,N_15057,N_15360);
and U16196 (N_16196,N_15086,N_15361);
or U16197 (N_16197,N_15045,N_15385);
nor U16198 (N_16198,N_15331,N_15071);
nor U16199 (N_16199,N_15445,N_15223);
nand U16200 (N_16200,N_15886,N_16115);
nand U16201 (N_16201,N_15853,N_15665);
or U16202 (N_16202,N_15661,N_15827);
xor U16203 (N_16203,N_15930,N_15650);
or U16204 (N_16204,N_15904,N_16069);
nor U16205 (N_16205,N_15803,N_16017);
xor U16206 (N_16206,N_15820,N_15859);
and U16207 (N_16207,N_15882,N_15828);
nand U16208 (N_16208,N_15795,N_16079);
nand U16209 (N_16209,N_15706,N_16065);
or U16210 (N_16210,N_15730,N_16000);
and U16211 (N_16211,N_15969,N_15919);
nor U16212 (N_16212,N_15658,N_15838);
and U16213 (N_16213,N_15979,N_15896);
xnor U16214 (N_16214,N_15961,N_15796);
and U16215 (N_16215,N_15681,N_15627);
or U16216 (N_16216,N_15967,N_15878);
nand U16217 (N_16217,N_16170,N_16198);
or U16218 (N_16218,N_15808,N_16083);
and U16219 (N_16219,N_15925,N_15909);
nand U16220 (N_16220,N_16076,N_15649);
nand U16221 (N_16221,N_16161,N_15678);
and U16222 (N_16222,N_15705,N_15943);
nand U16223 (N_16223,N_16106,N_15703);
and U16224 (N_16224,N_15867,N_16026);
nand U16225 (N_16225,N_15668,N_15852);
nand U16226 (N_16226,N_15955,N_15766);
nor U16227 (N_16227,N_15995,N_15986);
nor U16228 (N_16228,N_15667,N_15757);
nand U16229 (N_16229,N_15638,N_15713);
and U16230 (N_16230,N_15672,N_16098);
and U16231 (N_16231,N_15714,N_16038);
nand U16232 (N_16232,N_16158,N_15881);
nor U16233 (N_16233,N_15772,N_16027);
nor U16234 (N_16234,N_15855,N_15944);
nor U16235 (N_16235,N_15835,N_15850);
nand U16236 (N_16236,N_16007,N_16052);
or U16237 (N_16237,N_15611,N_15612);
and U16238 (N_16238,N_16041,N_15957);
or U16239 (N_16239,N_15809,N_15819);
or U16240 (N_16240,N_15785,N_16152);
and U16241 (N_16241,N_15916,N_15791);
nor U16242 (N_16242,N_15854,N_16105);
nand U16243 (N_16243,N_15635,N_15647);
nand U16244 (N_16244,N_15740,N_16133);
or U16245 (N_16245,N_16032,N_16188);
and U16246 (N_16246,N_15741,N_15839);
or U16247 (N_16247,N_16140,N_15604);
and U16248 (N_16248,N_16194,N_15966);
xnor U16249 (N_16249,N_15871,N_16103);
and U16250 (N_16250,N_16189,N_15920);
nand U16251 (N_16251,N_16139,N_16109);
and U16252 (N_16252,N_15862,N_15868);
nand U16253 (N_16253,N_16040,N_15847);
and U16254 (N_16254,N_15770,N_15712);
or U16255 (N_16255,N_15617,N_15794);
nand U16256 (N_16256,N_16055,N_16091);
nor U16257 (N_16257,N_16168,N_15998);
nor U16258 (N_16258,N_16048,N_16054);
and U16259 (N_16259,N_15980,N_16185);
nor U16260 (N_16260,N_16135,N_16180);
xnor U16261 (N_16261,N_15972,N_15620);
nand U16262 (N_16262,N_16049,N_15804);
xnor U16263 (N_16263,N_16031,N_15781);
or U16264 (N_16264,N_16111,N_15801);
and U16265 (N_16265,N_15610,N_15739);
and U16266 (N_16266,N_15737,N_16102);
xor U16267 (N_16267,N_15863,N_15716);
and U16268 (N_16268,N_15821,N_15824);
nand U16269 (N_16269,N_15945,N_16029);
nand U16270 (N_16270,N_15822,N_16149);
and U16271 (N_16271,N_16067,N_15630);
or U16272 (N_16272,N_15745,N_16124);
or U16273 (N_16273,N_15908,N_15616);
nor U16274 (N_16274,N_16036,N_16002);
nor U16275 (N_16275,N_16134,N_15790);
or U16276 (N_16276,N_15932,N_15768);
nand U16277 (N_16277,N_15985,N_15720);
xnor U16278 (N_16278,N_15990,N_16039);
nand U16279 (N_16279,N_15811,N_15989);
xnor U16280 (N_16280,N_16019,N_16119);
or U16281 (N_16281,N_15631,N_15776);
or U16282 (N_16282,N_15797,N_15732);
or U16283 (N_16283,N_15744,N_15912);
nor U16284 (N_16284,N_16154,N_15899);
xnor U16285 (N_16285,N_15701,N_15798);
nor U16286 (N_16286,N_15976,N_15700);
nor U16287 (N_16287,N_16128,N_15789);
xor U16288 (N_16288,N_16016,N_16130);
nor U16289 (N_16289,N_16051,N_15698);
xnor U16290 (N_16290,N_15775,N_15901);
xnor U16291 (N_16291,N_15953,N_15866);
nor U16292 (N_16292,N_16129,N_15949);
and U16293 (N_16293,N_16118,N_16110);
nor U16294 (N_16294,N_16196,N_15688);
xor U16295 (N_16295,N_15782,N_15763);
or U16296 (N_16296,N_15918,N_15632);
nand U16297 (N_16297,N_15929,N_16191);
nand U16298 (N_16298,N_16078,N_15625);
and U16299 (N_16299,N_15762,N_16075);
xor U16300 (N_16300,N_15940,N_15934);
nor U16301 (N_16301,N_16047,N_15893);
xor U16302 (N_16302,N_15876,N_16095);
or U16303 (N_16303,N_15965,N_16187);
nor U16304 (N_16304,N_15977,N_15885);
nand U16305 (N_16305,N_15687,N_15816);
and U16306 (N_16306,N_16126,N_15849);
and U16307 (N_16307,N_15845,N_15753);
nand U16308 (N_16308,N_16173,N_15606);
xor U16309 (N_16309,N_15880,N_16101);
nand U16310 (N_16310,N_15830,N_16160);
or U16311 (N_16311,N_16181,N_15749);
and U16312 (N_16312,N_16021,N_15659);
nor U16313 (N_16313,N_16023,N_16184);
xnor U16314 (N_16314,N_15778,N_16144);
and U16315 (N_16315,N_15890,N_16171);
xnor U16316 (N_16316,N_15626,N_15663);
nor U16317 (N_16317,N_16088,N_16192);
and U16318 (N_16318,N_16123,N_15993);
nor U16319 (N_16319,N_15767,N_16145);
and U16320 (N_16320,N_15842,N_15836);
or U16321 (N_16321,N_15709,N_15941);
or U16322 (N_16322,N_16070,N_15902);
and U16323 (N_16323,N_15914,N_16035);
xor U16324 (N_16324,N_15834,N_15846);
or U16325 (N_16325,N_15892,N_15900);
nor U16326 (N_16326,N_15642,N_15736);
nor U16327 (N_16327,N_15874,N_15906);
nor U16328 (N_16328,N_15897,N_16197);
or U16329 (N_16329,N_16193,N_15784);
nor U16330 (N_16330,N_15860,N_16009);
xor U16331 (N_16331,N_15946,N_15693);
or U16332 (N_16332,N_15725,N_15844);
nand U16333 (N_16333,N_16099,N_15677);
nand U16334 (N_16334,N_15652,N_16024);
and U16335 (N_16335,N_15910,N_16081);
nand U16336 (N_16336,N_15648,N_15869);
nor U16337 (N_16337,N_16082,N_15907);
nand U16338 (N_16338,N_15671,N_16072);
and U16339 (N_16339,N_16141,N_15666);
nand U16340 (N_16340,N_15807,N_15636);
and U16341 (N_16341,N_16094,N_15655);
xor U16342 (N_16342,N_15826,N_16014);
xnor U16343 (N_16343,N_15656,N_15779);
xnor U16344 (N_16344,N_15743,N_16068);
nor U16345 (N_16345,N_15856,N_15738);
and U16346 (N_16346,N_16142,N_15645);
or U16347 (N_16347,N_15673,N_15872);
and U16348 (N_16348,N_15702,N_15618);
xor U16349 (N_16349,N_15759,N_15686);
and U16350 (N_16350,N_15841,N_16008);
xor U16351 (N_16351,N_15723,N_15747);
nand U16352 (N_16352,N_15858,N_16074);
and U16353 (N_16353,N_15787,N_15950);
and U16354 (N_16354,N_15607,N_16003);
nand U16355 (N_16355,N_15697,N_15696);
xor U16356 (N_16356,N_15774,N_16195);
or U16357 (N_16357,N_16143,N_15734);
nand U16358 (N_16358,N_15963,N_15600);
nor U16359 (N_16359,N_16005,N_15613);
or U16360 (N_16360,N_15999,N_15962);
nor U16361 (N_16361,N_16136,N_15628);
and U16362 (N_16362,N_15857,N_15802);
nor U16363 (N_16363,N_15742,N_15621);
nand U16364 (N_16364,N_15889,N_16190);
or U16365 (N_16365,N_15695,N_15800);
nor U16366 (N_16366,N_15810,N_16004);
and U16367 (N_16367,N_15873,N_16182);
nand U16368 (N_16368,N_16117,N_15954);
nand U16369 (N_16369,N_16034,N_15923);
or U16370 (N_16370,N_16080,N_15711);
nand U16371 (N_16371,N_16179,N_15602);
nor U16372 (N_16372,N_16104,N_15691);
nor U16373 (N_16373,N_16097,N_15619);
xnor U16374 (N_16374,N_16122,N_15644);
or U16375 (N_16375,N_15765,N_16177);
or U16376 (N_16376,N_15664,N_15724);
xor U16377 (N_16377,N_16165,N_16164);
xnor U16378 (N_16378,N_16018,N_15973);
nor U16379 (N_16379,N_16107,N_16175);
xor U16380 (N_16380,N_15637,N_15833);
nand U16381 (N_16381,N_15913,N_15788);
and U16382 (N_16382,N_15817,N_16100);
or U16383 (N_16383,N_16157,N_15970);
xnor U16384 (N_16384,N_15684,N_15640);
and U16385 (N_16385,N_15984,N_15829);
or U16386 (N_16386,N_16132,N_15769);
or U16387 (N_16387,N_15639,N_16087);
or U16388 (N_16388,N_16011,N_16167);
and U16389 (N_16389,N_16178,N_15756);
nand U16390 (N_16390,N_16060,N_15722);
or U16391 (N_16391,N_16125,N_15771);
and U16392 (N_16392,N_16022,N_16147);
nand U16393 (N_16393,N_16153,N_15623);
and U16394 (N_16394,N_15605,N_15922);
or U16395 (N_16395,N_15685,N_16073);
and U16396 (N_16396,N_16174,N_15879);
nand U16397 (N_16397,N_15936,N_15812);
and U16398 (N_16398,N_15748,N_15773);
and U16399 (N_16399,N_16071,N_15641);
and U16400 (N_16400,N_15915,N_15996);
nand U16401 (N_16401,N_15964,N_15883);
and U16402 (N_16402,N_15680,N_16012);
nor U16403 (N_16403,N_15624,N_15894);
or U16404 (N_16404,N_15752,N_15926);
nand U16405 (N_16405,N_15699,N_16042);
and U16406 (N_16406,N_16062,N_16137);
xor U16407 (N_16407,N_16085,N_15848);
or U16408 (N_16408,N_15689,N_15662);
nor U16409 (N_16409,N_16030,N_15805);
and U16410 (N_16410,N_15751,N_15951);
or U16411 (N_16411,N_15608,N_15823);
nand U16412 (N_16412,N_15780,N_15750);
nand U16413 (N_16413,N_15861,N_15721);
nand U16414 (N_16414,N_15710,N_15622);
nor U16415 (N_16415,N_15733,N_16028);
and U16416 (N_16416,N_16176,N_16169);
and U16417 (N_16417,N_16058,N_16155);
xor U16418 (N_16418,N_15832,N_16172);
xor U16419 (N_16419,N_15992,N_16061);
nand U16420 (N_16420,N_15760,N_15674);
xnor U16421 (N_16421,N_15731,N_15937);
xor U16422 (N_16422,N_16001,N_15676);
nand U16423 (N_16423,N_15895,N_15755);
xor U16424 (N_16424,N_15994,N_15614);
nor U16425 (N_16425,N_15931,N_15707);
nor U16426 (N_16426,N_15870,N_15818);
xor U16427 (N_16427,N_15643,N_15975);
nand U16428 (N_16428,N_15669,N_16066);
nor U16429 (N_16429,N_16127,N_15657);
nor U16430 (N_16430,N_15793,N_15799);
and U16431 (N_16431,N_16020,N_16046);
nor U16432 (N_16432,N_15891,N_15815);
and U16433 (N_16433,N_15792,N_15983);
and U16434 (N_16434,N_15898,N_15921);
xnor U16435 (N_16435,N_15729,N_15903);
and U16436 (N_16436,N_15814,N_15806);
or U16437 (N_16437,N_15654,N_16092);
or U16438 (N_16438,N_15939,N_16156);
nand U16439 (N_16439,N_15646,N_15877);
or U16440 (N_16440,N_16120,N_16116);
or U16441 (N_16441,N_15968,N_15952);
xnor U16442 (N_16442,N_15997,N_15840);
and U16443 (N_16443,N_16146,N_15935);
xnor U16444 (N_16444,N_15813,N_15958);
xnor U16445 (N_16445,N_15679,N_15851);
nand U16446 (N_16446,N_16090,N_15735);
or U16447 (N_16447,N_15764,N_15991);
or U16448 (N_16448,N_15634,N_15708);
nand U16449 (N_16449,N_15988,N_15786);
and U16450 (N_16450,N_16093,N_16059);
and U16451 (N_16451,N_15948,N_16150);
nand U16452 (N_16452,N_15864,N_16186);
nor U16453 (N_16453,N_15746,N_16166);
or U16454 (N_16454,N_15758,N_15981);
or U16455 (N_16455,N_16084,N_15959);
and U16456 (N_16456,N_16089,N_15704);
xor U16457 (N_16457,N_15715,N_15629);
nor U16458 (N_16458,N_16025,N_15601);
and U16459 (N_16459,N_16138,N_15783);
and U16460 (N_16460,N_15942,N_15754);
or U16461 (N_16461,N_16056,N_16013);
xor U16462 (N_16462,N_15727,N_15887);
or U16463 (N_16463,N_15831,N_16112);
nand U16464 (N_16464,N_15938,N_16159);
or U16465 (N_16465,N_16010,N_15927);
nor U16466 (N_16466,N_16162,N_15683);
xnor U16467 (N_16467,N_15682,N_16053);
xnor U16468 (N_16468,N_16033,N_15777);
or U16469 (N_16469,N_16045,N_16006);
xnor U16470 (N_16470,N_15692,N_15651);
and U16471 (N_16471,N_15718,N_16163);
xnor U16472 (N_16472,N_15987,N_15843);
xor U16473 (N_16473,N_15960,N_15726);
or U16474 (N_16474,N_16183,N_15875);
nor U16475 (N_16475,N_15837,N_16096);
nor U16476 (N_16476,N_16151,N_15675);
xnor U16477 (N_16477,N_15888,N_15974);
nand U16478 (N_16478,N_15917,N_16086);
nor U16479 (N_16479,N_15905,N_15670);
nor U16480 (N_16480,N_16121,N_15947);
or U16481 (N_16481,N_15884,N_15694);
xor U16482 (N_16482,N_16113,N_15865);
or U16483 (N_16483,N_16114,N_16037);
and U16484 (N_16484,N_15933,N_16015);
nand U16485 (N_16485,N_15825,N_16057);
nand U16486 (N_16486,N_16199,N_16148);
or U16487 (N_16487,N_15633,N_15690);
and U16488 (N_16488,N_15761,N_16131);
nor U16489 (N_16489,N_15924,N_15609);
nand U16490 (N_16490,N_15603,N_15911);
and U16491 (N_16491,N_16044,N_15717);
nor U16492 (N_16492,N_15660,N_16063);
xnor U16493 (N_16493,N_16043,N_15978);
xnor U16494 (N_16494,N_16064,N_15728);
and U16495 (N_16495,N_16108,N_15956);
nand U16496 (N_16496,N_15982,N_15719);
nand U16497 (N_16497,N_16077,N_16050);
or U16498 (N_16498,N_15653,N_15615);
nand U16499 (N_16499,N_15971,N_15928);
or U16500 (N_16500,N_16167,N_15709);
xnor U16501 (N_16501,N_16133,N_15781);
nand U16502 (N_16502,N_15941,N_15963);
and U16503 (N_16503,N_15635,N_16008);
nor U16504 (N_16504,N_15842,N_15877);
and U16505 (N_16505,N_15716,N_15827);
xor U16506 (N_16506,N_15971,N_15879);
or U16507 (N_16507,N_15953,N_15932);
and U16508 (N_16508,N_15608,N_15602);
and U16509 (N_16509,N_15620,N_15796);
or U16510 (N_16510,N_15677,N_15929);
nor U16511 (N_16511,N_16009,N_16023);
nand U16512 (N_16512,N_15958,N_15617);
nor U16513 (N_16513,N_16040,N_15944);
nand U16514 (N_16514,N_16181,N_16083);
xor U16515 (N_16515,N_15848,N_16027);
nand U16516 (N_16516,N_15736,N_15800);
nand U16517 (N_16517,N_16014,N_15778);
or U16518 (N_16518,N_16165,N_15615);
nand U16519 (N_16519,N_15669,N_16083);
and U16520 (N_16520,N_15846,N_16005);
nand U16521 (N_16521,N_16196,N_15985);
nor U16522 (N_16522,N_16107,N_16187);
and U16523 (N_16523,N_15885,N_15832);
or U16524 (N_16524,N_15676,N_15958);
nor U16525 (N_16525,N_15880,N_16033);
nor U16526 (N_16526,N_15679,N_15685);
or U16527 (N_16527,N_16017,N_15782);
or U16528 (N_16528,N_15748,N_15994);
and U16529 (N_16529,N_16077,N_15714);
nand U16530 (N_16530,N_16187,N_16088);
or U16531 (N_16531,N_15675,N_15763);
or U16532 (N_16532,N_15746,N_16037);
and U16533 (N_16533,N_16189,N_15954);
nand U16534 (N_16534,N_15733,N_16081);
xnor U16535 (N_16535,N_15733,N_15888);
and U16536 (N_16536,N_16097,N_16139);
nor U16537 (N_16537,N_15849,N_15709);
nand U16538 (N_16538,N_15660,N_16031);
or U16539 (N_16539,N_15695,N_16053);
or U16540 (N_16540,N_15838,N_16008);
xor U16541 (N_16541,N_15636,N_15701);
xor U16542 (N_16542,N_16085,N_15675);
nor U16543 (N_16543,N_15739,N_16007);
nand U16544 (N_16544,N_16070,N_15997);
and U16545 (N_16545,N_16198,N_16179);
nand U16546 (N_16546,N_16189,N_15624);
and U16547 (N_16547,N_15954,N_16026);
and U16548 (N_16548,N_16048,N_16087);
nor U16549 (N_16549,N_15937,N_15941);
and U16550 (N_16550,N_15701,N_15869);
nor U16551 (N_16551,N_16104,N_15645);
or U16552 (N_16552,N_15759,N_15791);
or U16553 (N_16553,N_16141,N_16065);
and U16554 (N_16554,N_15644,N_15840);
nand U16555 (N_16555,N_15615,N_15797);
or U16556 (N_16556,N_15896,N_15985);
nand U16557 (N_16557,N_15890,N_16187);
or U16558 (N_16558,N_15737,N_15967);
or U16559 (N_16559,N_16146,N_15813);
and U16560 (N_16560,N_15691,N_16085);
and U16561 (N_16561,N_15809,N_16078);
and U16562 (N_16562,N_16015,N_16003);
nand U16563 (N_16563,N_16059,N_15922);
nor U16564 (N_16564,N_15870,N_16028);
or U16565 (N_16565,N_15931,N_15833);
and U16566 (N_16566,N_16161,N_16135);
nand U16567 (N_16567,N_15924,N_16014);
and U16568 (N_16568,N_15609,N_16194);
or U16569 (N_16569,N_16170,N_15881);
xnor U16570 (N_16570,N_15808,N_15944);
xnor U16571 (N_16571,N_15840,N_16199);
nand U16572 (N_16572,N_15957,N_15925);
xor U16573 (N_16573,N_15846,N_15702);
or U16574 (N_16574,N_16191,N_16062);
nor U16575 (N_16575,N_16181,N_16075);
or U16576 (N_16576,N_16145,N_15721);
nand U16577 (N_16577,N_15751,N_16069);
xnor U16578 (N_16578,N_16084,N_15907);
and U16579 (N_16579,N_15708,N_15859);
xor U16580 (N_16580,N_15670,N_16056);
and U16581 (N_16581,N_16083,N_15869);
nand U16582 (N_16582,N_15714,N_15601);
and U16583 (N_16583,N_16075,N_15953);
nor U16584 (N_16584,N_15704,N_16184);
nand U16585 (N_16585,N_16048,N_16181);
xor U16586 (N_16586,N_15752,N_15750);
nand U16587 (N_16587,N_15778,N_16094);
nor U16588 (N_16588,N_15728,N_16166);
or U16589 (N_16589,N_15776,N_15897);
nor U16590 (N_16590,N_15742,N_15757);
nand U16591 (N_16591,N_16082,N_15889);
xnor U16592 (N_16592,N_15979,N_15834);
or U16593 (N_16593,N_15702,N_15696);
or U16594 (N_16594,N_16088,N_15627);
or U16595 (N_16595,N_16091,N_15661);
nor U16596 (N_16596,N_15832,N_16082);
xor U16597 (N_16597,N_15888,N_15993);
or U16598 (N_16598,N_16121,N_15778);
nor U16599 (N_16599,N_16101,N_15993);
xor U16600 (N_16600,N_15638,N_16072);
nor U16601 (N_16601,N_16088,N_15602);
and U16602 (N_16602,N_15633,N_16182);
nor U16603 (N_16603,N_16022,N_16143);
or U16604 (N_16604,N_15882,N_15682);
xnor U16605 (N_16605,N_15928,N_16166);
xor U16606 (N_16606,N_16141,N_15811);
nor U16607 (N_16607,N_16159,N_15880);
nand U16608 (N_16608,N_16155,N_15673);
nand U16609 (N_16609,N_15881,N_16131);
nor U16610 (N_16610,N_16123,N_16185);
xnor U16611 (N_16611,N_15637,N_15771);
xor U16612 (N_16612,N_16163,N_16061);
and U16613 (N_16613,N_15621,N_16102);
or U16614 (N_16614,N_15772,N_15712);
nor U16615 (N_16615,N_15846,N_16011);
and U16616 (N_16616,N_16182,N_16157);
nand U16617 (N_16617,N_16067,N_15684);
nand U16618 (N_16618,N_16047,N_16038);
and U16619 (N_16619,N_15671,N_15789);
nand U16620 (N_16620,N_15737,N_15727);
nand U16621 (N_16621,N_15741,N_15613);
and U16622 (N_16622,N_15752,N_16090);
or U16623 (N_16623,N_15642,N_16114);
or U16624 (N_16624,N_15780,N_16128);
xor U16625 (N_16625,N_16132,N_16146);
and U16626 (N_16626,N_15957,N_15955);
and U16627 (N_16627,N_15805,N_16096);
nor U16628 (N_16628,N_15663,N_15965);
xnor U16629 (N_16629,N_16045,N_15788);
xor U16630 (N_16630,N_15717,N_15658);
nand U16631 (N_16631,N_15930,N_15702);
nand U16632 (N_16632,N_15617,N_16182);
nand U16633 (N_16633,N_16193,N_16113);
nand U16634 (N_16634,N_15908,N_15935);
xnor U16635 (N_16635,N_16084,N_15826);
nand U16636 (N_16636,N_15867,N_15974);
and U16637 (N_16637,N_15633,N_15924);
nor U16638 (N_16638,N_15943,N_15888);
nor U16639 (N_16639,N_15606,N_15791);
nor U16640 (N_16640,N_15925,N_15740);
xnor U16641 (N_16641,N_15709,N_16007);
and U16642 (N_16642,N_16096,N_15766);
xor U16643 (N_16643,N_15943,N_15804);
nand U16644 (N_16644,N_15854,N_15921);
and U16645 (N_16645,N_15663,N_15985);
or U16646 (N_16646,N_15869,N_15850);
and U16647 (N_16647,N_15600,N_15930);
or U16648 (N_16648,N_15624,N_15949);
and U16649 (N_16649,N_15894,N_15627);
nand U16650 (N_16650,N_15748,N_15665);
or U16651 (N_16651,N_15699,N_15869);
nand U16652 (N_16652,N_15615,N_15946);
xor U16653 (N_16653,N_15924,N_15988);
nand U16654 (N_16654,N_16055,N_15791);
xor U16655 (N_16655,N_15723,N_15801);
or U16656 (N_16656,N_16144,N_16189);
or U16657 (N_16657,N_15679,N_15683);
or U16658 (N_16658,N_15632,N_15806);
nor U16659 (N_16659,N_16165,N_16190);
nand U16660 (N_16660,N_15879,N_16020);
nor U16661 (N_16661,N_15632,N_15830);
nor U16662 (N_16662,N_16020,N_15695);
and U16663 (N_16663,N_15609,N_16131);
nand U16664 (N_16664,N_15795,N_15749);
xnor U16665 (N_16665,N_15923,N_15786);
nand U16666 (N_16666,N_16192,N_15813);
nor U16667 (N_16667,N_16090,N_15999);
nand U16668 (N_16668,N_15959,N_16082);
nor U16669 (N_16669,N_15848,N_16035);
or U16670 (N_16670,N_15934,N_15649);
nand U16671 (N_16671,N_16103,N_16164);
nor U16672 (N_16672,N_15811,N_15781);
xnor U16673 (N_16673,N_15882,N_15878);
nand U16674 (N_16674,N_16104,N_15897);
nor U16675 (N_16675,N_15824,N_16031);
nand U16676 (N_16676,N_15727,N_15977);
xnor U16677 (N_16677,N_16162,N_16111);
nand U16678 (N_16678,N_16098,N_15880);
nand U16679 (N_16679,N_16049,N_15826);
xor U16680 (N_16680,N_16075,N_15611);
nor U16681 (N_16681,N_16183,N_15706);
xnor U16682 (N_16682,N_15690,N_15785);
xnor U16683 (N_16683,N_15974,N_15902);
nand U16684 (N_16684,N_15722,N_15816);
and U16685 (N_16685,N_16124,N_15785);
nand U16686 (N_16686,N_16180,N_16032);
and U16687 (N_16687,N_15667,N_16150);
nor U16688 (N_16688,N_15888,N_15668);
xnor U16689 (N_16689,N_15687,N_15808);
nor U16690 (N_16690,N_15857,N_15687);
and U16691 (N_16691,N_15917,N_15709);
nor U16692 (N_16692,N_15873,N_15647);
nand U16693 (N_16693,N_16123,N_15870);
nand U16694 (N_16694,N_15622,N_15895);
nor U16695 (N_16695,N_15826,N_16092);
and U16696 (N_16696,N_15724,N_15881);
xor U16697 (N_16697,N_16099,N_15803);
nand U16698 (N_16698,N_16165,N_16070);
nor U16699 (N_16699,N_16198,N_16071);
nand U16700 (N_16700,N_15751,N_15638);
nand U16701 (N_16701,N_15716,N_15814);
xor U16702 (N_16702,N_15722,N_16186);
xor U16703 (N_16703,N_16087,N_15983);
xnor U16704 (N_16704,N_15867,N_15923);
nand U16705 (N_16705,N_16179,N_15876);
nor U16706 (N_16706,N_15840,N_15955);
nand U16707 (N_16707,N_16152,N_16094);
nand U16708 (N_16708,N_15995,N_16118);
xnor U16709 (N_16709,N_15690,N_16159);
xnor U16710 (N_16710,N_15732,N_16038);
or U16711 (N_16711,N_15618,N_16168);
and U16712 (N_16712,N_15927,N_16062);
nand U16713 (N_16713,N_15612,N_15670);
nor U16714 (N_16714,N_15639,N_15725);
or U16715 (N_16715,N_16064,N_15822);
or U16716 (N_16716,N_15663,N_15970);
and U16717 (N_16717,N_16093,N_15680);
nor U16718 (N_16718,N_15683,N_15640);
or U16719 (N_16719,N_16172,N_15744);
or U16720 (N_16720,N_15802,N_15882);
xnor U16721 (N_16721,N_16029,N_15912);
or U16722 (N_16722,N_15780,N_16190);
nor U16723 (N_16723,N_15693,N_16131);
xor U16724 (N_16724,N_15686,N_15914);
and U16725 (N_16725,N_15694,N_15741);
xor U16726 (N_16726,N_16023,N_15881);
xor U16727 (N_16727,N_15853,N_15760);
and U16728 (N_16728,N_15632,N_16134);
nor U16729 (N_16729,N_16094,N_15967);
xnor U16730 (N_16730,N_15676,N_16016);
nand U16731 (N_16731,N_15883,N_15758);
xor U16732 (N_16732,N_15637,N_16034);
xor U16733 (N_16733,N_15958,N_15914);
or U16734 (N_16734,N_16045,N_15629);
nand U16735 (N_16735,N_16082,N_15915);
or U16736 (N_16736,N_15651,N_15799);
and U16737 (N_16737,N_15848,N_15692);
xnor U16738 (N_16738,N_15624,N_15976);
nor U16739 (N_16739,N_15612,N_15938);
or U16740 (N_16740,N_15681,N_15672);
nor U16741 (N_16741,N_15900,N_15634);
or U16742 (N_16742,N_15601,N_15837);
nor U16743 (N_16743,N_15948,N_15910);
and U16744 (N_16744,N_15861,N_15639);
or U16745 (N_16745,N_15739,N_16128);
nor U16746 (N_16746,N_16160,N_15913);
or U16747 (N_16747,N_16056,N_16173);
xnor U16748 (N_16748,N_16042,N_16109);
and U16749 (N_16749,N_15690,N_15612);
or U16750 (N_16750,N_15608,N_15724);
xnor U16751 (N_16751,N_16006,N_15631);
and U16752 (N_16752,N_16006,N_15648);
nor U16753 (N_16753,N_15624,N_16126);
nor U16754 (N_16754,N_15904,N_16066);
nor U16755 (N_16755,N_15679,N_16025);
and U16756 (N_16756,N_16147,N_15890);
nand U16757 (N_16757,N_15841,N_15728);
xnor U16758 (N_16758,N_15790,N_16047);
nor U16759 (N_16759,N_15858,N_15688);
or U16760 (N_16760,N_16192,N_15795);
xor U16761 (N_16761,N_15930,N_15943);
xor U16762 (N_16762,N_16079,N_15982);
and U16763 (N_16763,N_16185,N_16057);
nand U16764 (N_16764,N_15807,N_15798);
or U16765 (N_16765,N_16199,N_16147);
and U16766 (N_16766,N_15999,N_16116);
or U16767 (N_16767,N_15997,N_16016);
nand U16768 (N_16768,N_16155,N_16153);
nand U16769 (N_16769,N_16187,N_16117);
and U16770 (N_16770,N_15626,N_16074);
or U16771 (N_16771,N_15648,N_15763);
or U16772 (N_16772,N_15803,N_15789);
or U16773 (N_16773,N_15606,N_15607);
or U16774 (N_16774,N_16141,N_15799);
xor U16775 (N_16775,N_15820,N_15608);
nand U16776 (N_16776,N_16049,N_16160);
xnor U16777 (N_16777,N_16178,N_15914);
xor U16778 (N_16778,N_15794,N_15775);
and U16779 (N_16779,N_15661,N_16083);
xnor U16780 (N_16780,N_16011,N_15837);
xnor U16781 (N_16781,N_15993,N_15655);
and U16782 (N_16782,N_16189,N_16024);
and U16783 (N_16783,N_15814,N_16160);
nand U16784 (N_16784,N_15744,N_15980);
xnor U16785 (N_16785,N_15777,N_15972);
and U16786 (N_16786,N_15925,N_15883);
nand U16787 (N_16787,N_15617,N_15777);
nand U16788 (N_16788,N_16062,N_15658);
nor U16789 (N_16789,N_15636,N_15669);
xnor U16790 (N_16790,N_15973,N_15746);
nand U16791 (N_16791,N_15860,N_16035);
and U16792 (N_16792,N_15948,N_15794);
and U16793 (N_16793,N_16152,N_15916);
nand U16794 (N_16794,N_16100,N_15643);
xor U16795 (N_16795,N_16092,N_16171);
xor U16796 (N_16796,N_15720,N_15668);
nor U16797 (N_16797,N_15766,N_15917);
and U16798 (N_16798,N_15935,N_15639);
nand U16799 (N_16799,N_15688,N_16133);
nand U16800 (N_16800,N_16733,N_16253);
and U16801 (N_16801,N_16554,N_16405);
nor U16802 (N_16802,N_16383,N_16746);
and U16803 (N_16803,N_16755,N_16664);
nand U16804 (N_16804,N_16787,N_16744);
or U16805 (N_16805,N_16718,N_16707);
xnor U16806 (N_16806,N_16201,N_16630);
nand U16807 (N_16807,N_16551,N_16501);
or U16808 (N_16808,N_16596,N_16628);
xnor U16809 (N_16809,N_16672,N_16452);
xor U16810 (N_16810,N_16447,N_16429);
nand U16811 (N_16811,N_16430,N_16298);
xor U16812 (N_16812,N_16602,N_16606);
or U16813 (N_16813,N_16682,N_16562);
xor U16814 (N_16814,N_16489,N_16417);
or U16815 (N_16815,N_16775,N_16369);
or U16816 (N_16816,N_16327,N_16764);
or U16817 (N_16817,N_16293,N_16490);
and U16818 (N_16818,N_16530,N_16565);
nor U16819 (N_16819,N_16559,N_16712);
nand U16820 (N_16820,N_16622,N_16593);
nor U16821 (N_16821,N_16415,N_16462);
nor U16822 (N_16822,N_16423,N_16548);
xor U16823 (N_16823,N_16739,N_16276);
or U16824 (N_16824,N_16458,N_16419);
or U16825 (N_16825,N_16643,N_16541);
and U16826 (N_16826,N_16629,N_16491);
xnor U16827 (N_16827,N_16334,N_16705);
nand U16828 (N_16828,N_16400,N_16307);
and U16829 (N_16829,N_16588,N_16403);
xor U16830 (N_16830,N_16555,N_16756);
nand U16831 (N_16831,N_16326,N_16219);
nand U16832 (N_16832,N_16519,N_16473);
nor U16833 (N_16833,N_16757,N_16557);
and U16834 (N_16834,N_16401,N_16552);
or U16835 (N_16835,N_16432,N_16494);
or U16836 (N_16836,N_16485,N_16679);
or U16837 (N_16837,N_16619,N_16671);
nor U16838 (N_16838,N_16260,N_16259);
xnor U16839 (N_16839,N_16637,N_16795);
nor U16840 (N_16840,N_16304,N_16624);
and U16841 (N_16841,N_16478,N_16623);
and U16842 (N_16842,N_16512,N_16526);
and U16843 (N_16843,N_16498,N_16355);
nor U16844 (N_16844,N_16675,N_16697);
and U16845 (N_16845,N_16218,N_16451);
nor U16846 (N_16846,N_16251,N_16231);
nand U16847 (N_16847,N_16751,N_16314);
nor U16848 (N_16848,N_16514,N_16324);
xor U16849 (N_16849,N_16250,N_16439);
or U16850 (N_16850,N_16564,N_16266);
nand U16851 (N_16851,N_16377,N_16550);
or U16852 (N_16852,N_16396,N_16418);
nand U16853 (N_16853,N_16684,N_16468);
or U16854 (N_16854,N_16654,N_16657);
xor U16855 (N_16855,N_16496,N_16653);
or U16856 (N_16856,N_16603,N_16566);
nand U16857 (N_16857,N_16204,N_16502);
xor U16858 (N_16858,N_16380,N_16706);
xor U16859 (N_16859,N_16763,N_16299);
and U16860 (N_16860,N_16661,N_16291);
and U16861 (N_16861,N_16558,N_16772);
nand U16862 (N_16862,N_16736,N_16782);
xnor U16863 (N_16863,N_16513,N_16210);
nor U16864 (N_16864,N_16337,N_16495);
and U16865 (N_16865,N_16248,N_16649);
nor U16866 (N_16866,N_16776,N_16670);
nand U16867 (N_16867,N_16261,N_16793);
xnor U16868 (N_16868,N_16389,N_16446);
nor U16869 (N_16869,N_16797,N_16209);
or U16870 (N_16870,N_16683,N_16594);
xor U16871 (N_16871,N_16711,N_16433);
or U16872 (N_16872,N_16573,N_16268);
nand U16873 (N_16873,N_16504,N_16421);
nor U16874 (N_16874,N_16295,N_16642);
xor U16875 (N_16875,N_16262,N_16243);
nand U16876 (N_16876,N_16408,N_16282);
xor U16877 (N_16877,N_16246,N_16450);
or U16878 (N_16878,N_16445,N_16789);
nor U16879 (N_16879,N_16686,N_16488);
xnor U16880 (N_16880,N_16778,N_16680);
nor U16881 (N_16881,N_16639,N_16455);
xnor U16882 (N_16882,N_16788,N_16272);
or U16883 (N_16883,N_16374,N_16339);
nand U16884 (N_16884,N_16545,N_16375);
and U16885 (N_16885,N_16576,N_16613);
nand U16886 (N_16886,N_16297,N_16636);
or U16887 (N_16887,N_16715,N_16615);
xnor U16888 (N_16888,N_16581,N_16748);
or U16889 (N_16889,N_16437,N_16651);
or U16890 (N_16890,N_16505,N_16652);
nand U16891 (N_16891,N_16730,N_16540);
xnor U16892 (N_16892,N_16691,N_16200);
nor U16893 (N_16893,N_16372,N_16704);
xnor U16894 (N_16894,N_16290,N_16416);
nor U16895 (N_16895,N_16471,N_16463);
xor U16896 (N_16896,N_16567,N_16318);
nand U16897 (N_16897,N_16647,N_16743);
or U16898 (N_16898,N_16228,N_16348);
nor U16899 (N_16899,N_16402,N_16759);
nor U16900 (N_16900,N_16393,N_16523);
or U16901 (N_16901,N_16745,N_16331);
or U16902 (N_16902,N_16710,N_16328);
and U16903 (N_16903,N_16235,N_16784);
nand U16904 (N_16904,N_16359,N_16525);
nor U16905 (N_16905,N_16645,N_16760);
nand U16906 (N_16906,N_16330,N_16363);
nand U16907 (N_16907,N_16611,N_16758);
and U16908 (N_16908,N_16285,N_16256);
nor U16909 (N_16909,N_16294,N_16798);
or U16910 (N_16910,N_16738,N_16434);
nand U16911 (N_16911,N_16280,N_16750);
nor U16912 (N_16912,N_16522,N_16510);
nor U16913 (N_16913,N_16729,N_16720);
nor U16914 (N_16914,N_16224,N_16534);
nor U16915 (N_16915,N_16366,N_16741);
and U16916 (N_16916,N_16516,N_16234);
nor U16917 (N_16917,N_16215,N_16395);
or U16918 (N_16918,N_16466,N_16258);
xnor U16919 (N_16919,N_16783,N_16308);
and U16920 (N_16920,N_16589,N_16579);
nand U16921 (N_16921,N_16518,N_16221);
and U16922 (N_16922,N_16665,N_16600);
or U16923 (N_16923,N_16352,N_16353);
or U16924 (N_16924,N_16226,N_16765);
and U16925 (N_16925,N_16538,N_16317);
nand U16926 (N_16926,N_16799,N_16791);
and U16927 (N_16927,N_16220,N_16693);
nor U16928 (N_16928,N_16336,N_16321);
nor U16929 (N_16929,N_16217,N_16278);
xor U16930 (N_16930,N_16539,N_16263);
xnor U16931 (N_16931,N_16205,N_16371);
nand U16932 (N_16932,N_16794,N_16486);
nand U16933 (N_16933,N_16482,N_16406);
nand U16934 (N_16934,N_16203,N_16271);
nor U16935 (N_16935,N_16673,N_16236);
nand U16936 (N_16936,N_16460,N_16781);
nor U16937 (N_16937,N_16747,N_16277);
or U16938 (N_16938,N_16472,N_16364);
nor U16939 (N_16939,N_16431,N_16244);
xor U16940 (N_16940,N_16598,N_16583);
nor U16941 (N_16941,N_16255,N_16230);
nor U16942 (N_16942,N_16238,N_16681);
nand U16943 (N_16943,N_16560,N_16289);
xor U16944 (N_16944,N_16597,N_16785);
or U16945 (N_16945,N_16279,N_16790);
xor U16946 (N_16946,N_16695,N_16608);
nor U16947 (N_16947,N_16356,N_16737);
or U16948 (N_16948,N_16570,N_16265);
and U16949 (N_16949,N_16254,N_16225);
or U16950 (N_16950,N_16283,N_16604);
nand U16951 (N_16951,N_16329,N_16731);
xnor U16952 (N_16952,N_16634,N_16520);
and U16953 (N_16953,N_16216,N_16240);
nor U16954 (N_16954,N_16275,N_16666);
xnor U16955 (N_16955,N_16378,N_16753);
nor U16956 (N_16956,N_16724,N_16392);
or U16957 (N_16957,N_16614,N_16655);
nor U16958 (N_16958,N_16477,N_16590);
xnor U16959 (N_16959,N_16341,N_16620);
or U16960 (N_16960,N_16333,N_16273);
nor U16961 (N_16961,N_16346,N_16792);
xor U16962 (N_16962,N_16373,N_16440);
and U16963 (N_16963,N_16311,N_16553);
nand U16964 (N_16964,N_16397,N_16700);
or U16965 (N_16965,N_16459,N_16556);
nor U16966 (N_16966,N_16752,N_16726);
nand U16967 (N_16967,N_16441,N_16703);
nand U16968 (N_16968,N_16281,N_16420);
nor U16969 (N_16969,N_16245,N_16270);
or U16970 (N_16970,N_16368,N_16702);
xor U16971 (N_16971,N_16587,N_16667);
xnor U16972 (N_16972,N_16233,N_16592);
xor U16973 (N_16973,N_16500,N_16696);
nor U16974 (N_16974,N_16528,N_16508);
or U16975 (N_16975,N_16610,N_16476);
and U16976 (N_16976,N_16762,N_16475);
nor U16977 (N_16977,N_16379,N_16487);
nand U16978 (N_16978,N_16668,N_16537);
nor U16979 (N_16979,N_16529,N_16612);
xor U16980 (N_16980,N_16267,N_16777);
xnor U16981 (N_16981,N_16444,N_16319);
or U16982 (N_16982,N_16521,N_16780);
xor U16983 (N_16983,N_16467,N_16524);
xnor U16984 (N_16984,N_16428,N_16320);
or U16985 (N_16985,N_16584,N_16699);
nand U16986 (N_16986,N_16338,N_16728);
and U16987 (N_16987,N_16347,N_16438);
or U16988 (N_16988,N_16384,N_16616);
nor U16989 (N_16989,N_16771,N_16207);
xnor U16990 (N_16990,N_16701,N_16399);
nand U16991 (N_16991,N_16309,N_16786);
nand U16992 (N_16992,N_16342,N_16621);
and U16993 (N_16993,N_16345,N_16507);
xnor U16994 (N_16994,N_16527,N_16465);
and U16995 (N_16995,N_16768,N_16533);
and U16996 (N_16996,N_16544,N_16674);
or U16997 (N_16997,N_16698,N_16411);
and U16998 (N_16998,N_16350,N_16692);
xor U16999 (N_16999,N_16663,N_16386);
nand U17000 (N_17000,N_16409,N_16761);
nor U17001 (N_17001,N_16381,N_16274);
nor U17002 (N_17002,N_16727,N_16766);
and U17003 (N_17003,N_16300,N_16424);
nor U17004 (N_17004,N_16625,N_16388);
nor U17005 (N_17005,N_16484,N_16288);
nand U17006 (N_17006,N_16769,N_16713);
nor U17007 (N_17007,N_16313,N_16492);
nand U17008 (N_17008,N_16626,N_16227);
nor U17009 (N_17009,N_16499,N_16332);
or U17010 (N_17010,N_16515,N_16725);
nor U17011 (N_17011,N_16264,N_16578);
and U17012 (N_17012,N_16365,N_16412);
and U17013 (N_17013,N_16607,N_16532);
nand U17014 (N_17014,N_16662,N_16571);
and U17015 (N_17015,N_16493,N_16360);
or U17016 (N_17016,N_16208,N_16456);
xnor U17017 (N_17017,N_16362,N_16249);
nor U17018 (N_17018,N_16586,N_16640);
and U17019 (N_17019,N_16676,N_16394);
nor U17020 (N_17020,N_16660,N_16453);
and U17021 (N_17021,N_16252,N_16301);
xnor U17022 (N_17022,N_16382,N_16410);
or U17023 (N_17023,N_16497,N_16591);
or U17024 (N_17024,N_16483,N_16694);
nand U17025 (N_17025,N_16237,N_16580);
or U17026 (N_17026,N_16464,N_16722);
and U17027 (N_17027,N_16442,N_16425);
nor U17028 (N_17028,N_16214,N_16656);
and U17029 (N_17029,N_16443,N_16582);
nor U17030 (N_17030,N_16323,N_16632);
and U17031 (N_17031,N_16511,N_16517);
nor U17032 (N_17032,N_16232,N_16469);
xnor U17033 (N_17033,N_16689,N_16367);
or U17034 (N_17034,N_16646,N_16796);
nor U17035 (N_17035,N_16561,N_16357);
nand U17036 (N_17036,N_16316,N_16312);
nor U17037 (N_17037,N_16688,N_16742);
xor U17038 (N_17038,N_16480,N_16638);
nand U17039 (N_17039,N_16569,N_16413);
and U17040 (N_17040,N_16286,N_16422);
nor U17041 (N_17041,N_16754,N_16644);
xnor U17042 (N_17042,N_16773,N_16574);
xnor U17043 (N_17043,N_16229,N_16770);
or U17044 (N_17044,N_16322,N_16457);
or U17045 (N_17045,N_16641,N_16242);
and U17046 (N_17046,N_16648,N_16387);
xnor U17047 (N_17047,N_16536,N_16677);
nor U17048 (N_17048,N_16376,N_16354);
nor U17049 (N_17049,N_16284,N_16474);
nand U17050 (N_17050,N_16454,N_16351);
or U17051 (N_17051,N_16325,N_16358);
xnor U17052 (N_17052,N_16734,N_16721);
and U17053 (N_17053,N_16202,N_16749);
xor U17054 (N_17054,N_16257,N_16435);
nor U17055 (N_17055,N_16658,N_16310);
or U17056 (N_17056,N_16585,N_16206);
xor U17057 (N_17057,N_16735,N_16449);
and U17058 (N_17058,N_16344,N_16343);
nor U17059 (N_17059,N_16407,N_16549);
nor U17060 (N_17060,N_16223,N_16635);
xnor U17061 (N_17061,N_16740,N_16709);
or U17062 (N_17062,N_16631,N_16687);
and U17063 (N_17063,N_16398,N_16774);
or U17064 (N_17064,N_16575,N_16685);
or U17065 (N_17065,N_16404,N_16213);
nand U17066 (N_17066,N_16426,N_16296);
and U17067 (N_17067,N_16436,N_16601);
and U17068 (N_17068,N_16577,N_16335);
and U17069 (N_17069,N_16719,N_16650);
nand U17070 (N_17070,N_16292,N_16595);
xor U17071 (N_17071,N_16678,N_16531);
and U17072 (N_17072,N_16627,N_16535);
nor U17073 (N_17073,N_16563,N_16287);
and U17074 (N_17074,N_16470,N_16509);
nand U17075 (N_17075,N_16659,N_16302);
nand U17076 (N_17076,N_16546,N_16361);
nor U17077 (N_17077,N_16506,N_16716);
and U17078 (N_17078,N_16690,N_16222);
or U17079 (N_17079,N_16212,N_16385);
or U17080 (N_17080,N_16211,N_16247);
nor U17081 (N_17081,N_16568,N_16479);
nor U17082 (N_17082,N_16414,N_16303);
xor U17083 (N_17083,N_16708,N_16779);
nand U17084 (N_17084,N_16547,N_16269);
or U17085 (N_17085,N_16241,N_16448);
nand U17086 (N_17086,N_16461,N_16370);
or U17087 (N_17087,N_16239,N_16315);
nor U17088 (N_17088,N_16767,N_16717);
xnor U17089 (N_17089,N_16714,N_16669);
and U17090 (N_17090,N_16391,N_16599);
or U17091 (N_17091,N_16349,N_16732);
and U17092 (N_17092,N_16427,N_16503);
nor U17093 (N_17093,N_16390,N_16617);
nand U17094 (N_17094,N_16340,N_16605);
nor U17095 (N_17095,N_16618,N_16572);
xor U17096 (N_17096,N_16542,N_16609);
nand U17097 (N_17097,N_16723,N_16481);
nor U17098 (N_17098,N_16305,N_16543);
xor U17099 (N_17099,N_16306,N_16633);
nand U17100 (N_17100,N_16353,N_16201);
or U17101 (N_17101,N_16277,N_16316);
nor U17102 (N_17102,N_16720,N_16382);
nand U17103 (N_17103,N_16479,N_16263);
or U17104 (N_17104,N_16383,N_16391);
xnor U17105 (N_17105,N_16291,N_16735);
nor U17106 (N_17106,N_16690,N_16781);
nor U17107 (N_17107,N_16581,N_16269);
nor U17108 (N_17108,N_16675,N_16469);
xnor U17109 (N_17109,N_16342,N_16280);
or U17110 (N_17110,N_16296,N_16535);
nor U17111 (N_17111,N_16220,N_16685);
nand U17112 (N_17112,N_16395,N_16234);
or U17113 (N_17113,N_16657,N_16313);
nand U17114 (N_17114,N_16667,N_16419);
xor U17115 (N_17115,N_16767,N_16630);
nor U17116 (N_17116,N_16346,N_16370);
nand U17117 (N_17117,N_16788,N_16450);
nand U17118 (N_17118,N_16456,N_16424);
nand U17119 (N_17119,N_16438,N_16788);
and U17120 (N_17120,N_16591,N_16477);
xnor U17121 (N_17121,N_16514,N_16626);
or U17122 (N_17122,N_16426,N_16739);
nor U17123 (N_17123,N_16267,N_16729);
and U17124 (N_17124,N_16424,N_16219);
nand U17125 (N_17125,N_16396,N_16224);
nor U17126 (N_17126,N_16237,N_16568);
nand U17127 (N_17127,N_16336,N_16305);
nor U17128 (N_17128,N_16604,N_16475);
and U17129 (N_17129,N_16311,N_16624);
nand U17130 (N_17130,N_16586,N_16261);
nand U17131 (N_17131,N_16287,N_16250);
nand U17132 (N_17132,N_16771,N_16244);
nand U17133 (N_17133,N_16564,N_16756);
nor U17134 (N_17134,N_16758,N_16368);
nand U17135 (N_17135,N_16707,N_16410);
nor U17136 (N_17136,N_16539,N_16789);
nand U17137 (N_17137,N_16604,N_16598);
xnor U17138 (N_17138,N_16330,N_16774);
nand U17139 (N_17139,N_16225,N_16701);
nand U17140 (N_17140,N_16247,N_16795);
nand U17141 (N_17141,N_16575,N_16310);
and U17142 (N_17142,N_16443,N_16744);
or U17143 (N_17143,N_16672,N_16505);
xnor U17144 (N_17144,N_16750,N_16778);
and U17145 (N_17145,N_16614,N_16682);
xor U17146 (N_17146,N_16778,N_16404);
nand U17147 (N_17147,N_16769,N_16784);
xor U17148 (N_17148,N_16321,N_16729);
xnor U17149 (N_17149,N_16365,N_16557);
or U17150 (N_17150,N_16747,N_16675);
nand U17151 (N_17151,N_16447,N_16240);
nand U17152 (N_17152,N_16277,N_16552);
or U17153 (N_17153,N_16694,N_16552);
or U17154 (N_17154,N_16748,N_16710);
and U17155 (N_17155,N_16334,N_16282);
or U17156 (N_17156,N_16711,N_16674);
xor U17157 (N_17157,N_16512,N_16529);
nand U17158 (N_17158,N_16626,N_16332);
nand U17159 (N_17159,N_16617,N_16531);
nor U17160 (N_17160,N_16293,N_16202);
nand U17161 (N_17161,N_16295,N_16286);
or U17162 (N_17162,N_16458,N_16404);
or U17163 (N_17163,N_16475,N_16415);
and U17164 (N_17164,N_16695,N_16770);
and U17165 (N_17165,N_16626,N_16516);
nor U17166 (N_17166,N_16348,N_16257);
xnor U17167 (N_17167,N_16411,N_16797);
and U17168 (N_17168,N_16587,N_16213);
or U17169 (N_17169,N_16325,N_16772);
or U17170 (N_17170,N_16327,N_16638);
xor U17171 (N_17171,N_16530,N_16321);
or U17172 (N_17172,N_16584,N_16590);
nand U17173 (N_17173,N_16759,N_16655);
nand U17174 (N_17174,N_16203,N_16277);
nor U17175 (N_17175,N_16322,N_16666);
xor U17176 (N_17176,N_16463,N_16420);
nor U17177 (N_17177,N_16220,N_16526);
nor U17178 (N_17178,N_16489,N_16552);
or U17179 (N_17179,N_16282,N_16385);
xnor U17180 (N_17180,N_16267,N_16228);
and U17181 (N_17181,N_16582,N_16713);
and U17182 (N_17182,N_16306,N_16624);
nor U17183 (N_17183,N_16316,N_16275);
nor U17184 (N_17184,N_16267,N_16345);
and U17185 (N_17185,N_16485,N_16576);
nand U17186 (N_17186,N_16259,N_16676);
or U17187 (N_17187,N_16763,N_16557);
nand U17188 (N_17188,N_16641,N_16528);
nor U17189 (N_17189,N_16422,N_16298);
nand U17190 (N_17190,N_16514,N_16448);
or U17191 (N_17191,N_16409,N_16364);
nor U17192 (N_17192,N_16657,N_16612);
xnor U17193 (N_17193,N_16752,N_16585);
or U17194 (N_17194,N_16320,N_16227);
nand U17195 (N_17195,N_16598,N_16661);
and U17196 (N_17196,N_16689,N_16686);
or U17197 (N_17197,N_16435,N_16313);
or U17198 (N_17198,N_16303,N_16431);
or U17199 (N_17199,N_16584,N_16620);
nor U17200 (N_17200,N_16716,N_16201);
and U17201 (N_17201,N_16344,N_16488);
xnor U17202 (N_17202,N_16457,N_16795);
xor U17203 (N_17203,N_16238,N_16563);
nor U17204 (N_17204,N_16787,N_16758);
nor U17205 (N_17205,N_16395,N_16525);
and U17206 (N_17206,N_16734,N_16209);
and U17207 (N_17207,N_16504,N_16404);
nand U17208 (N_17208,N_16667,N_16462);
nand U17209 (N_17209,N_16766,N_16280);
nand U17210 (N_17210,N_16748,N_16785);
or U17211 (N_17211,N_16491,N_16369);
nor U17212 (N_17212,N_16358,N_16376);
or U17213 (N_17213,N_16530,N_16624);
or U17214 (N_17214,N_16703,N_16780);
or U17215 (N_17215,N_16340,N_16613);
nor U17216 (N_17216,N_16652,N_16709);
or U17217 (N_17217,N_16593,N_16710);
or U17218 (N_17218,N_16588,N_16732);
xnor U17219 (N_17219,N_16501,N_16202);
xnor U17220 (N_17220,N_16792,N_16332);
or U17221 (N_17221,N_16686,N_16266);
nand U17222 (N_17222,N_16477,N_16704);
or U17223 (N_17223,N_16485,N_16791);
xnor U17224 (N_17224,N_16642,N_16275);
nor U17225 (N_17225,N_16222,N_16305);
nor U17226 (N_17226,N_16326,N_16465);
or U17227 (N_17227,N_16612,N_16203);
and U17228 (N_17228,N_16466,N_16430);
xor U17229 (N_17229,N_16300,N_16543);
xnor U17230 (N_17230,N_16296,N_16357);
nand U17231 (N_17231,N_16516,N_16433);
nor U17232 (N_17232,N_16608,N_16516);
or U17233 (N_17233,N_16768,N_16614);
or U17234 (N_17234,N_16441,N_16492);
nor U17235 (N_17235,N_16633,N_16347);
or U17236 (N_17236,N_16764,N_16796);
or U17237 (N_17237,N_16567,N_16484);
nand U17238 (N_17238,N_16626,N_16476);
nand U17239 (N_17239,N_16727,N_16238);
nand U17240 (N_17240,N_16605,N_16727);
nand U17241 (N_17241,N_16641,N_16211);
and U17242 (N_17242,N_16688,N_16565);
nand U17243 (N_17243,N_16541,N_16692);
nor U17244 (N_17244,N_16688,N_16484);
nand U17245 (N_17245,N_16481,N_16781);
xor U17246 (N_17246,N_16245,N_16773);
nand U17247 (N_17247,N_16317,N_16439);
and U17248 (N_17248,N_16785,N_16431);
nand U17249 (N_17249,N_16460,N_16677);
nor U17250 (N_17250,N_16650,N_16407);
and U17251 (N_17251,N_16621,N_16631);
xnor U17252 (N_17252,N_16301,N_16287);
nor U17253 (N_17253,N_16499,N_16732);
and U17254 (N_17254,N_16560,N_16346);
and U17255 (N_17255,N_16493,N_16374);
and U17256 (N_17256,N_16479,N_16316);
or U17257 (N_17257,N_16348,N_16411);
and U17258 (N_17258,N_16684,N_16409);
nand U17259 (N_17259,N_16603,N_16753);
or U17260 (N_17260,N_16232,N_16298);
or U17261 (N_17261,N_16280,N_16637);
or U17262 (N_17262,N_16745,N_16627);
nor U17263 (N_17263,N_16686,N_16653);
and U17264 (N_17264,N_16497,N_16502);
xnor U17265 (N_17265,N_16452,N_16269);
nor U17266 (N_17266,N_16359,N_16351);
nand U17267 (N_17267,N_16311,N_16797);
or U17268 (N_17268,N_16654,N_16798);
nor U17269 (N_17269,N_16436,N_16236);
nor U17270 (N_17270,N_16485,N_16553);
nand U17271 (N_17271,N_16573,N_16385);
xor U17272 (N_17272,N_16628,N_16575);
and U17273 (N_17273,N_16369,N_16225);
and U17274 (N_17274,N_16275,N_16451);
or U17275 (N_17275,N_16669,N_16361);
nor U17276 (N_17276,N_16510,N_16660);
or U17277 (N_17277,N_16282,N_16515);
nand U17278 (N_17278,N_16265,N_16737);
or U17279 (N_17279,N_16463,N_16349);
xor U17280 (N_17280,N_16208,N_16674);
and U17281 (N_17281,N_16582,N_16480);
and U17282 (N_17282,N_16612,N_16509);
nand U17283 (N_17283,N_16203,N_16629);
or U17284 (N_17284,N_16764,N_16436);
nor U17285 (N_17285,N_16383,N_16647);
or U17286 (N_17286,N_16574,N_16604);
nor U17287 (N_17287,N_16652,N_16380);
nand U17288 (N_17288,N_16678,N_16612);
or U17289 (N_17289,N_16607,N_16300);
or U17290 (N_17290,N_16508,N_16548);
xnor U17291 (N_17291,N_16375,N_16705);
nor U17292 (N_17292,N_16664,N_16712);
or U17293 (N_17293,N_16655,N_16362);
or U17294 (N_17294,N_16491,N_16514);
or U17295 (N_17295,N_16287,N_16321);
and U17296 (N_17296,N_16638,N_16411);
or U17297 (N_17297,N_16440,N_16200);
xor U17298 (N_17298,N_16264,N_16761);
nand U17299 (N_17299,N_16678,N_16445);
nand U17300 (N_17300,N_16204,N_16430);
xor U17301 (N_17301,N_16585,N_16576);
nand U17302 (N_17302,N_16553,N_16250);
or U17303 (N_17303,N_16620,N_16411);
and U17304 (N_17304,N_16688,N_16569);
or U17305 (N_17305,N_16539,N_16428);
xnor U17306 (N_17306,N_16752,N_16666);
and U17307 (N_17307,N_16781,N_16479);
nor U17308 (N_17308,N_16200,N_16270);
nor U17309 (N_17309,N_16383,N_16768);
xor U17310 (N_17310,N_16755,N_16347);
nor U17311 (N_17311,N_16250,N_16234);
or U17312 (N_17312,N_16271,N_16566);
xor U17313 (N_17313,N_16705,N_16759);
nor U17314 (N_17314,N_16695,N_16283);
and U17315 (N_17315,N_16768,N_16776);
nand U17316 (N_17316,N_16314,N_16453);
and U17317 (N_17317,N_16519,N_16542);
nand U17318 (N_17318,N_16663,N_16686);
and U17319 (N_17319,N_16424,N_16340);
or U17320 (N_17320,N_16749,N_16434);
and U17321 (N_17321,N_16210,N_16374);
nor U17322 (N_17322,N_16362,N_16522);
or U17323 (N_17323,N_16249,N_16276);
nand U17324 (N_17324,N_16776,N_16550);
or U17325 (N_17325,N_16683,N_16714);
and U17326 (N_17326,N_16364,N_16459);
and U17327 (N_17327,N_16249,N_16211);
nor U17328 (N_17328,N_16467,N_16209);
nor U17329 (N_17329,N_16585,N_16674);
or U17330 (N_17330,N_16465,N_16588);
xnor U17331 (N_17331,N_16682,N_16673);
nor U17332 (N_17332,N_16517,N_16651);
nand U17333 (N_17333,N_16576,N_16674);
nand U17334 (N_17334,N_16353,N_16468);
xnor U17335 (N_17335,N_16662,N_16517);
nand U17336 (N_17336,N_16359,N_16694);
xnor U17337 (N_17337,N_16695,N_16615);
or U17338 (N_17338,N_16268,N_16281);
or U17339 (N_17339,N_16697,N_16502);
nor U17340 (N_17340,N_16302,N_16649);
xnor U17341 (N_17341,N_16764,N_16777);
and U17342 (N_17342,N_16541,N_16674);
xor U17343 (N_17343,N_16218,N_16337);
nand U17344 (N_17344,N_16293,N_16352);
nor U17345 (N_17345,N_16390,N_16612);
and U17346 (N_17346,N_16210,N_16782);
nand U17347 (N_17347,N_16798,N_16459);
xor U17348 (N_17348,N_16374,N_16658);
xnor U17349 (N_17349,N_16274,N_16463);
nand U17350 (N_17350,N_16446,N_16229);
xnor U17351 (N_17351,N_16296,N_16609);
nand U17352 (N_17352,N_16384,N_16542);
nor U17353 (N_17353,N_16428,N_16371);
nand U17354 (N_17354,N_16713,N_16783);
nor U17355 (N_17355,N_16309,N_16771);
or U17356 (N_17356,N_16516,N_16277);
or U17357 (N_17357,N_16223,N_16245);
xor U17358 (N_17358,N_16712,N_16679);
nand U17359 (N_17359,N_16591,N_16582);
nand U17360 (N_17360,N_16749,N_16659);
nand U17361 (N_17361,N_16710,N_16266);
or U17362 (N_17362,N_16412,N_16741);
xor U17363 (N_17363,N_16423,N_16303);
nand U17364 (N_17364,N_16686,N_16779);
and U17365 (N_17365,N_16206,N_16473);
or U17366 (N_17366,N_16423,N_16669);
and U17367 (N_17367,N_16506,N_16501);
nor U17368 (N_17368,N_16761,N_16295);
or U17369 (N_17369,N_16575,N_16261);
or U17370 (N_17370,N_16674,N_16275);
or U17371 (N_17371,N_16650,N_16347);
nand U17372 (N_17372,N_16290,N_16366);
nand U17373 (N_17373,N_16797,N_16379);
or U17374 (N_17374,N_16575,N_16779);
nand U17375 (N_17375,N_16594,N_16454);
xor U17376 (N_17376,N_16695,N_16558);
nand U17377 (N_17377,N_16562,N_16432);
xor U17378 (N_17378,N_16550,N_16792);
nand U17379 (N_17379,N_16529,N_16604);
or U17380 (N_17380,N_16501,N_16773);
nor U17381 (N_17381,N_16210,N_16327);
and U17382 (N_17382,N_16668,N_16529);
xor U17383 (N_17383,N_16264,N_16627);
or U17384 (N_17384,N_16558,N_16764);
nand U17385 (N_17385,N_16680,N_16667);
nand U17386 (N_17386,N_16752,N_16646);
and U17387 (N_17387,N_16525,N_16526);
nor U17388 (N_17388,N_16681,N_16269);
xnor U17389 (N_17389,N_16787,N_16736);
and U17390 (N_17390,N_16299,N_16480);
or U17391 (N_17391,N_16265,N_16451);
xor U17392 (N_17392,N_16487,N_16317);
nand U17393 (N_17393,N_16453,N_16458);
nor U17394 (N_17394,N_16222,N_16757);
xnor U17395 (N_17395,N_16244,N_16677);
or U17396 (N_17396,N_16563,N_16565);
xnor U17397 (N_17397,N_16783,N_16344);
or U17398 (N_17398,N_16679,N_16249);
nor U17399 (N_17399,N_16796,N_16439);
nor U17400 (N_17400,N_16899,N_17234);
xnor U17401 (N_17401,N_17317,N_17299);
nand U17402 (N_17402,N_17241,N_17075);
xnor U17403 (N_17403,N_17045,N_17322);
nor U17404 (N_17404,N_17292,N_17202);
and U17405 (N_17405,N_17186,N_17362);
and U17406 (N_17406,N_17331,N_17065);
xor U17407 (N_17407,N_17313,N_17129);
nor U17408 (N_17408,N_17181,N_17268);
nor U17409 (N_17409,N_17219,N_17354);
nor U17410 (N_17410,N_17191,N_17023);
nor U17411 (N_17411,N_16819,N_17260);
nor U17412 (N_17412,N_16845,N_16816);
nand U17413 (N_17413,N_17270,N_16924);
nor U17414 (N_17414,N_17022,N_17286);
nor U17415 (N_17415,N_16846,N_17300);
xor U17416 (N_17416,N_17176,N_17247);
and U17417 (N_17417,N_17013,N_16946);
or U17418 (N_17418,N_17112,N_16910);
nand U17419 (N_17419,N_16891,N_17388);
or U17420 (N_17420,N_17215,N_17337);
nor U17421 (N_17421,N_17303,N_17040);
or U17422 (N_17422,N_16893,N_16979);
or U17423 (N_17423,N_17077,N_17352);
or U17424 (N_17424,N_17068,N_16943);
and U17425 (N_17425,N_17096,N_16894);
xnor U17426 (N_17426,N_17309,N_17204);
nor U17427 (N_17427,N_17055,N_17175);
nand U17428 (N_17428,N_17277,N_17381);
xnor U17429 (N_17429,N_16855,N_17335);
xor U17430 (N_17430,N_17320,N_17248);
nand U17431 (N_17431,N_17285,N_16942);
nand U17432 (N_17432,N_17069,N_16962);
or U17433 (N_17433,N_17377,N_16945);
or U17434 (N_17434,N_16853,N_16976);
and U17435 (N_17435,N_17090,N_16960);
xnor U17436 (N_17436,N_17095,N_17177);
nor U17437 (N_17437,N_17263,N_17258);
nand U17438 (N_17438,N_16867,N_17036);
xnor U17439 (N_17439,N_17029,N_16836);
xnor U17440 (N_17440,N_17272,N_17019);
nand U17441 (N_17441,N_17012,N_17153);
and U17442 (N_17442,N_17238,N_17025);
nand U17443 (N_17443,N_16869,N_17171);
or U17444 (N_17444,N_17061,N_16915);
nor U17445 (N_17445,N_17017,N_16801);
xnor U17446 (N_17446,N_17127,N_16827);
or U17447 (N_17447,N_17318,N_17372);
nand U17448 (N_17448,N_17330,N_16844);
nor U17449 (N_17449,N_16951,N_17106);
and U17450 (N_17450,N_17146,N_16849);
nor U17451 (N_17451,N_16829,N_17102);
and U17452 (N_17452,N_17060,N_17047);
xnor U17453 (N_17453,N_16858,N_17133);
nand U17454 (N_17454,N_17305,N_17071);
or U17455 (N_17455,N_16848,N_17244);
and U17456 (N_17456,N_17150,N_17130);
and U17457 (N_17457,N_17093,N_17000);
xor U17458 (N_17458,N_17342,N_17197);
xor U17459 (N_17459,N_16825,N_17304);
nor U17460 (N_17460,N_16980,N_17203);
nand U17461 (N_17461,N_17020,N_17345);
nor U17462 (N_17462,N_17135,N_17218);
and U17463 (N_17463,N_17076,N_17373);
nor U17464 (N_17464,N_17233,N_17333);
or U17465 (N_17465,N_17161,N_16870);
xor U17466 (N_17466,N_17306,N_16922);
xnor U17467 (N_17467,N_17144,N_17166);
xnor U17468 (N_17468,N_17289,N_17028);
and U17469 (N_17469,N_16935,N_16938);
and U17470 (N_17470,N_17397,N_16807);
and U17471 (N_17471,N_17230,N_17113);
or U17472 (N_17472,N_17010,N_17399);
and U17473 (N_17473,N_17240,N_16859);
nand U17474 (N_17474,N_16874,N_16991);
nor U17475 (N_17475,N_16931,N_16965);
and U17476 (N_17476,N_17126,N_17201);
and U17477 (N_17477,N_16863,N_16914);
nand U17478 (N_17478,N_17349,N_17274);
nor U17479 (N_17479,N_17250,N_17243);
xnor U17480 (N_17480,N_16852,N_16964);
nand U17481 (N_17481,N_17251,N_17190);
or U17482 (N_17482,N_16972,N_17207);
xnor U17483 (N_17483,N_17189,N_17236);
xnor U17484 (N_17484,N_17004,N_17284);
or U17485 (N_17485,N_17375,N_17343);
nand U17486 (N_17486,N_16973,N_17001);
xor U17487 (N_17487,N_17136,N_16838);
and U17488 (N_17488,N_16895,N_17363);
or U17489 (N_17489,N_17054,N_16969);
and U17490 (N_17490,N_17092,N_17152);
nor U17491 (N_17491,N_17174,N_17114);
nor U17492 (N_17492,N_16947,N_17137);
nand U17493 (N_17493,N_17097,N_17057);
or U17494 (N_17494,N_17315,N_17051);
and U17495 (N_17495,N_17367,N_16865);
or U17496 (N_17496,N_17160,N_17027);
nand U17497 (N_17497,N_17334,N_17101);
nand U17498 (N_17498,N_16934,N_16984);
nor U17499 (N_17499,N_16996,N_17366);
and U17500 (N_17500,N_16989,N_16916);
nand U17501 (N_17501,N_16927,N_17246);
or U17502 (N_17502,N_17182,N_16957);
nor U17503 (N_17503,N_16904,N_17231);
nand U17504 (N_17504,N_17262,N_16820);
nor U17505 (N_17505,N_17086,N_16803);
nor U17506 (N_17506,N_16955,N_17346);
or U17507 (N_17507,N_17326,N_17217);
nor U17508 (N_17508,N_17016,N_16993);
or U17509 (N_17509,N_17259,N_17257);
xnor U17510 (N_17510,N_17100,N_17026);
and U17511 (N_17511,N_17111,N_17383);
or U17512 (N_17512,N_17324,N_17206);
xnor U17513 (N_17513,N_16982,N_17142);
and U17514 (N_17514,N_17216,N_16908);
xnor U17515 (N_17515,N_17145,N_16889);
and U17516 (N_17516,N_17103,N_16890);
xnor U17517 (N_17517,N_16990,N_17371);
or U17518 (N_17518,N_17037,N_16995);
nand U17519 (N_17519,N_16886,N_16833);
xor U17520 (N_17520,N_17296,N_16831);
xor U17521 (N_17521,N_17155,N_16949);
and U17522 (N_17522,N_17063,N_16911);
nor U17523 (N_17523,N_16987,N_16923);
and U17524 (N_17524,N_16876,N_16808);
and U17525 (N_17525,N_17364,N_16902);
or U17526 (N_17526,N_17167,N_17163);
nand U17527 (N_17527,N_16861,N_17173);
nor U17528 (N_17528,N_16907,N_17098);
xor U17529 (N_17529,N_17214,N_17070);
or U17530 (N_17530,N_17120,N_17325);
or U17531 (N_17531,N_16868,N_16818);
nor U17532 (N_17532,N_17183,N_16978);
xor U17533 (N_17533,N_17121,N_17083);
nand U17534 (N_17534,N_17254,N_16887);
nand U17535 (N_17535,N_17132,N_17165);
and U17536 (N_17536,N_16856,N_17297);
xnor U17537 (N_17537,N_17269,N_17385);
or U17538 (N_17538,N_17172,N_17099);
or U17539 (N_17539,N_17221,N_16847);
nand U17540 (N_17540,N_16968,N_17006);
and U17541 (N_17541,N_17396,N_17356);
xor U17542 (N_17542,N_17311,N_16805);
xnor U17543 (N_17543,N_16954,N_17185);
and U17544 (N_17544,N_17290,N_17389);
nor U17545 (N_17545,N_17082,N_17359);
and U17546 (N_17546,N_17050,N_17323);
or U17547 (N_17547,N_17107,N_16871);
and U17548 (N_17548,N_17156,N_17351);
and U17549 (N_17549,N_16961,N_17344);
nand U17550 (N_17550,N_16999,N_17105);
nand U17551 (N_17551,N_17229,N_17079);
nand U17552 (N_17552,N_16997,N_16941);
nor U17553 (N_17553,N_17162,N_17225);
or U17554 (N_17554,N_17141,N_16842);
nand U17555 (N_17555,N_16953,N_16821);
or U17556 (N_17556,N_17316,N_17275);
nor U17557 (N_17557,N_17108,N_16885);
and U17558 (N_17558,N_17222,N_17123);
and U17559 (N_17559,N_16906,N_16981);
nor U17560 (N_17560,N_17003,N_17252);
nand U17561 (N_17561,N_17031,N_17293);
nand U17562 (N_17562,N_17287,N_17194);
nand U17563 (N_17563,N_17291,N_17208);
nand U17564 (N_17564,N_17005,N_17384);
nor U17565 (N_17565,N_17188,N_16988);
nand U17566 (N_17566,N_16860,N_17298);
nor U17567 (N_17567,N_16880,N_16937);
xnor U17568 (N_17568,N_17209,N_17224);
or U17569 (N_17569,N_17310,N_17210);
nor U17570 (N_17570,N_17347,N_17376);
nand U17571 (N_17571,N_16840,N_16862);
and U17572 (N_17572,N_17053,N_17007);
or U17573 (N_17573,N_16888,N_16866);
nand U17574 (N_17574,N_16878,N_16854);
and U17575 (N_17575,N_16851,N_16948);
nor U17576 (N_17576,N_17339,N_17294);
nand U17577 (N_17577,N_16919,N_17187);
and U17578 (N_17578,N_17237,N_16921);
and U17579 (N_17579,N_16814,N_16966);
and U17580 (N_17580,N_17281,N_17276);
and U17581 (N_17581,N_17308,N_16971);
and U17582 (N_17582,N_16909,N_17193);
nor U17583 (N_17583,N_17211,N_17340);
and U17584 (N_17584,N_17391,N_17213);
xnor U17585 (N_17585,N_17115,N_17032);
and U17586 (N_17586,N_17264,N_16959);
nor U17587 (N_17587,N_17018,N_17169);
and U17588 (N_17588,N_17128,N_16952);
xnor U17589 (N_17589,N_17052,N_17361);
or U17590 (N_17590,N_16802,N_17242);
and U17591 (N_17591,N_16932,N_16837);
nand U17592 (N_17592,N_16839,N_16967);
nor U17593 (N_17593,N_17282,N_16832);
nand U17594 (N_17594,N_17073,N_16817);
and U17595 (N_17595,N_16898,N_16873);
or U17596 (N_17596,N_16857,N_16929);
nand U17597 (N_17597,N_17280,N_17048);
and U17598 (N_17598,N_17042,N_17198);
nand U17599 (N_17599,N_16926,N_16963);
or U17600 (N_17600,N_16811,N_16815);
or U17601 (N_17601,N_16994,N_17200);
and U17602 (N_17602,N_16970,N_17398);
xor U17603 (N_17603,N_17085,N_16804);
xor U17604 (N_17604,N_17283,N_17255);
xnor U17605 (N_17605,N_17266,N_17245);
and U17606 (N_17606,N_17149,N_16822);
xor U17607 (N_17607,N_17271,N_17196);
and U17608 (N_17608,N_17232,N_17002);
and U17609 (N_17609,N_17332,N_16944);
and U17610 (N_17610,N_17253,N_16974);
nor U17611 (N_17611,N_17064,N_17011);
nand U17612 (N_17612,N_16826,N_17386);
or U17613 (N_17613,N_17038,N_17009);
nor U17614 (N_17614,N_17109,N_17394);
nand U17615 (N_17615,N_16875,N_17159);
and U17616 (N_17616,N_17091,N_17360);
or U17617 (N_17617,N_17140,N_17044);
or U17618 (N_17618,N_16913,N_17072);
nand U17619 (N_17619,N_17279,N_16998);
and U17620 (N_17620,N_17139,N_17131);
and U17621 (N_17621,N_17393,N_16975);
and U17622 (N_17622,N_16879,N_17365);
and U17623 (N_17623,N_16896,N_17235);
nor U17624 (N_17624,N_17049,N_16939);
or U17625 (N_17625,N_16930,N_17226);
nor U17626 (N_17626,N_17273,N_17212);
or U17627 (N_17627,N_17164,N_17327);
nor U17628 (N_17628,N_17261,N_16956);
xnor U17629 (N_17629,N_16892,N_16950);
xor U17630 (N_17630,N_17369,N_17094);
or U17631 (N_17631,N_16936,N_16872);
nor U17632 (N_17632,N_16983,N_16823);
and U17633 (N_17633,N_17307,N_17024);
xnor U17634 (N_17634,N_17014,N_16809);
or U17635 (N_17635,N_17195,N_16810);
or U17636 (N_17636,N_17265,N_17056);
and U17637 (N_17637,N_17059,N_16918);
or U17638 (N_17638,N_17074,N_16806);
and U17639 (N_17639,N_16812,N_17084);
or U17640 (N_17640,N_16977,N_17089);
xor U17641 (N_17641,N_16830,N_16813);
nand U17642 (N_17642,N_17033,N_17312);
nand U17643 (N_17643,N_17179,N_16843);
and U17644 (N_17644,N_17302,N_17267);
nand U17645 (N_17645,N_17184,N_17104);
xnor U17646 (N_17646,N_17041,N_16881);
nand U17647 (N_17647,N_17157,N_17021);
and U17648 (N_17648,N_17087,N_16985);
and U17649 (N_17649,N_17321,N_17116);
nand U17650 (N_17650,N_17088,N_17357);
or U17651 (N_17651,N_17078,N_17081);
nor U17652 (N_17652,N_17125,N_17119);
or U17653 (N_17653,N_16883,N_17353);
nand U17654 (N_17654,N_17301,N_17046);
nand U17655 (N_17655,N_17338,N_16835);
nand U17656 (N_17656,N_17341,N_16958);
and U17657 (N_17657,N_17035,N_17328);
xor U17658 (N_17658,N_17058,N_16824);
and U17659 (N_17659,N_17066,N_17178);
and U17660 (N_17660,N_16834,N_16900);
nand U17661 (N_17661,N_17249,N_16992);
nand U17662 (N_17662,N_17374,N_16800);
or U17663 (N_17663,N_17180,N_17239);
nand U17664 (N_17664,N_17392,N_16884);
and U17665 (N_17665,N_16905,N_17329);
nor U17666 (N_17666,N_17158,N_17370);
xor U17667 (N_17667,N_17143,N_17387);
nand U17668 (N_17668,N_17034,N_17278);
nand U17669 (N_17669,N_17015,N_17220);
nor U17670 (N_17670,N_17199,N_17350);
or U17671 (N_17671,N_16928,N_17043);
and U17672 (N_17672,N_17080,N_16917);
or U17673 (N_17673,N_17039,N_17228);
and U17674 (N_17674,N_16877,N_17348);
or U17675 (N_17675,N_16901,N_17168);
nand U17676 (N_17676,N_16986,N_17008);
nand U17677 (N_17677,N_16940,N_17223);
or U17678 (N_17678,N_17336,N_17288);
nor U17679 (N_17679,N_16912,N_17117);
or U17680 (N_17680,N_16933,N_16828);
and U17681 (N_17681,N_17170,N_17147);
and U17682 (N_17682,N_17382,N_17368);
xnor U17683 (N_17683,N_17030,N_17355);
nor U17684 (N_17684,N_17314,N_17295);
or U17685 (N_17685,N_16841,N_17118);
and U17686 (N_17686,N_17067,N_17138);
xor U17687 (N_17687,N_17380,N_17062);
nor U17688 (N_17688,N_17390,N_17192);
nor U17689 (N_17689,N_17256,N_16903);
or U17690 (N_17690,N_17205,N_17319);
nor U17691 (N_17691,N_16897,N_16882);
and U17692 (N_17692,N_17151,N_17395);
nand U17693 (N_17693,N_16920,N_17110);
nor U17694 (N_17694,N_17154,N_16850);
xor U17695 (N_17695,N_17378,N_17122);
or U17696 (N_17696,N_17134,N_17124);
nor U17697 (N_17697,N_17358,N_17227);
nor U17698 (N_17698,N_16925,N_17379);
or U17699 (N_17699,N_17148,N_16864);
and U17700 (N_17700,N_16919,N_17189);
xor U17701 (N_17701,N_17054,N_16843);
nor U17702 (N_17702,N_17277,N_17114);
nor U17703 (N_17703,N_17020,N_16820);
nand U17704 (N_17704,N_17086,N_17105);
xnor U17705 (N_17705,N_17327,N_17236);
xnor U17706 (N_17706,N_16841,N_17061);
nor U17707 (N_17707,N_17109,N_16991);
nand U17708 (N_17708,N_17055,N_16823);
or U17709 (N_17709,N_16912,N_17366);
and U17710 (N_17710,N_16938,N_17218);
or U17711 (N_17711,N_17225,N_17222);
and U17712 (N_17712,N_16849,N_16893);
nand U17713 (N_17713,N_16958,N_17183);
nor U17714 (N_17714,N_17035,N_17001);
nand U17715 (N_17715,N_17287,N_17215);
nor U17716 (N_17716,N_16883,N_17365);
and U17717 (N_17717,N_16862,N_17053);
and U17718 (N_17718,N_17294,N_17089);
and U17719 (N_17719,N_17232,N_17301);
xnor U17720 (N_17720,N_16920,N_17286);
nand U17721 (N_17721,N_16935,N_16801);
xnor U17722 (N_17722,N_16818,N_17302);
nand U17723 (N_17723,N_17148,N_16930);
or U17724 (N_17724,N_17150,N_16937);
and U17725 (N_17725,N_16871,N_16818);
nor U17726 (N_17726,N_16938,N_17253);
nand U17727 (N_17727,N_17309,N_16949);
nor U17728 (N_17728,N_17055,N_17340);
xnor U17729 (N_17729,N_17139,N_17391);
or U17730 (N_17730,N_17119,N_16936);
nor U17731 (N_17731,N_17175,N_17122);
or U17732 (N_17732,N_17178,N_17047);
nand U17733 (N_17733,N_16829,N_17223);
xnor U17734 (N_17734,N_17021,N_16886);
or U17735 (N_17735,N_17252,N_17054);
nor U17736 (N_17736,N_16845,N_16988);
nor U17737 (N_17737,N_17248,N_16806);
nand U17738 (N_17738,N_16969,N_17273);
nor U17739 (N_17739,N_16883,N_17144);
nor U17740 (N_17740,N_17144,N_17390);
nor U17741 (N_17741,N_16912,N_16985);
or U17742 (N_17742,N_17126,N_17221);
nor U17743 (N_17743,N_17354,N_17043);
and U17744 (N_17744,N_17205,N_17391);
and U17745 (N_17745,N_17240,N_17007);
nand U17746 (N_17746,N_16910,N_17100);
nor U17747 (N_17747,N_16931,N_17320);
xnor U17748 (N_17748,N_16953,N_17074);
nand U17749 (N_17749,N_17126,N_17058);
and U17750 (N_17750,N_16817,N_16852);
nand U17751 (N_17751,N_16895,N_17308);
nor U17752 (N_17752,N_17155,N_16826);
xor U17753 (N_17753,N_17355,N_17295);
nor U17754 (N_17754,N_17374,N_16882);
and U17755 (N_17755,N_17354,N_17134);
nor U17756 (N_17756,N_16833,N_16813);
xnor U17757 (N_17757,N_17375,N_16835);
and U17758 (N_17758,N_17275,N_16885);
xor U17759 (N_17759,N_17353,N_17025);
nor U17760 (N_17760,N_17246,N_17381);
or U17761 (N_17761,N_17282,N_17328);
nor U17762 (N_17762,N_17159,N_16959);
nand U17763 (N_17763,N_17337,N_17213);
nand U17764 (N_17764,N_17245,N_17134);
xnor U17765 (N_17765,N_17214,N_17080);
and U17766 (N_17766,N_17271,N_17217);
and U17767 (N_17767,N_17209,N_17274);
and U17768 (N_17768,N_16932,N_17028);
or U17769 (N_17769,N_17221,N_16850);
nand U17770 (N_17770,N_16800,N_17362);
xor U17771 (N_17771,N_17353,N_17244);
nand U17772 (N_17772,N_16990,N_17025);
or U17773 (N_17773,N_16934,N_16861);
xnor U17774 (N_17774,N_17254,N_17146);
nand U17775 (N_17775,N_17339,N_17303);
and U17776 (N_17776,N_17149,N_17362);
and U17777 (N_17777,N_17239,N_16997);
nand U17778 (N_17778,N_16950,N_16885);
nand U17779 (N_17779,N_17095,N_17329);
nor U17780 (N_17780,N_17339,N_17176);
and U17781 (N_17781,N_16913,N_17365);
or U17782 (N_17782,N_17278,N_17358);
or U17783 (N_17783,N_16991,N_17033);
and U17784 (N_17784,N_17363,N_17046);
and U17785 (N_17785,N_17390,N_16890);
nand U17786 (N_17786,N_17135,N_17025);
nor U17787 (N_17787,N_16857,N_17365);
or U17788 (N_17788,N_16986,N_17056);
or U17789 (N_17789,N_17276,N_16920);
and U17790 (N_17790,N_16872,N_17181);
nand U17791 (N_17791,N_17197,N_16886);
or U17792 (N_17792,N_17026,N_17372);
xnor U17793 (N_17793,N_16826,N_16946);
nand U17794 (N_17794,N_17107,N_17364);
nor U17795 (N_17795,N_17179,N_17270);
nor U17796 (N_17796,N_17335,N_16871);
and U17797 (N_17797,N_17230,N_16888);
nor U17798 (N_17798,N_17159,N_16889);
nor U17799 (N_17799,N_17094,N_17321);
xnor U17800 (N_17800,N_17175,N_17216);
xnor U17801 (N_17801,N_17213,N_17016);
nor U17802 (N_17802,N_17012,N_17347);
nor U17803 (N_17803,N_17186,N_17066);
or U17804 (N_17804,N_17258,N_17199);
and U17805 (N_17805,N_17351,N_17071);
nand U17806 (N_17806,N_16978,N_16915);
and U17807 (N_17807,N_16836,N_16828);
and U17808 (N_17808,N_17133,N_17364);
xnor U17809 (N_17809,N_16890,N_17199);
xor U17810 (N_17810,N_17200,N_17178);
nor U17811 (N_17811,N_17250,N_17019);
nand U17812 (N_17812,N_16954,N_17064);
nand U17813 (N_17813,N_17149,N_17390);
or U17814 (N_17814,N_17390,N_16834);
nand U17815 (N_17815,N_16885,N_17252);
xnor U17816 (N_17816,N_16835,N_16874);
or U17817 (N_17817,N_17194,N_17351);
nor U17818 (N_17818,N_17105,N_16969);
xnor U17819 (N_17819,N_17030,N_16982);
and U17820 (N_17820,N_17030,N_16896);
xnor U17821 (N_17821,N_17106,N_17314);
nor U17822 (N_17822,N_17395,N_17160);
and U17823 (N_17823,N_16836,N_17040);
nor U17824 (N_17824,N_16991,N_16811);
nor U17825 (N_17825,N_17329,N_17325);
and U17826 (N_17826,N_16954,N_16965);
nand U17827 (N_17827,N_17152,N_16960);
or U17828 (N_17828,N_17017,N_17178);
and U17829 (N_17829,N_16962,N_17372);
and U17830 (N_17830,N_16940,N_17369);
nor U17831 (N_17831,N_17230,N_17348);
xnor U17832 (N_17832,N_17220,N_16998);
xnor U17833 (N_17833,N_17313,N_17230);
and U17834 (N_17834,N_17287,N_16832);
and U17835 (N_17835,N_17380,N_17089);
xor U17836 (N_17836,N_17369,N_17232);
xor U17837 (N_17837,N_17119,N_17305);
xor U17838 (N_17838,N_17012,N_17229);
nor U17839 (N_17839,N_17029,N_17014);
nand U17840 (N_17840,N_16987,N_17083);
nand U17841 (N_17841,N_17214,N_17282);
or U17842 (N_17842,N_16958,N_17063);
and U17843 (N_17843,N_17367,N_17241);
nor U17844 (N_17844,N_17291,N_16941);
and U17845 (N_17845,N_17309,N_17008);
nand U17846 (N_17846,N_17008,N_17001);
or U17847 (N_17847,N_17355,N_17185);
xor U17848 (N_17848,N_17068,N_17072);
nand U17849 (N_17849,N_17082,N_16842);
nor U17850 (N_17850,N_17168,N_17275);
nand U17851 (N_17851,N_17086,N_17144);
nand U17852 (N_17852,N_16863,N_17226);
xnor U17853 (N_17853,N_17038,N_17013);
or U17854 (N_17854,N_17376,N_17137);
and U17855 (N_17855,N_17180,N_17108);
or U17856 (N_17856,N_17163,N_17340);
nor U17857 (N_17857,N_17192,N_17395);
nand U17858 (N_17858,N_16886,N_17188);
nor U17859 (N_17859,N_16814,N_17044);
nor U17860 (N_17860,N_17153,N_17203);
and U17861 (N_17861,N_17163,N_17074);
or U17862 (N_17862,N_17132,N_17006);
nand U17863 (N_17863,N_17030,N_17371);
xnor U17864 (N_17864,N_17335,N_17050);
nand U17865 (N_17865,N_17237,N_17329);
or U17866 (N_17866,N_17045,N_16843);
nand U17867 (N_17867,N_17162,N_16975);
xnor U17868 (N_17868,N_16923,N_17121);
nand U17869 (N_17869,N_17144,N_16944);
or U17870 (N_17870,N_16895,N_16932);
or U17871 (N_17871,N_17240,N_17326);
nand U17872 (N_17872,N_17327,N_16906);
and U17873 (N_17873,N_17214,N_17272);
nand U17874 (N_17874,N_17349,N_17172);
nand U17875 (N_17875,N_17198,N_17364);
or U17876 (N_17876,N_16852,N_17375);
nor U17877 (N_17877,N_16891,N_17119);
xnor U17878 (N_17878,N_17255,N_17170);
nor U17879 (N_17879,N_16854,N_17028);
or U17880 (N_17880,N_17104,N_17335);
nor U17881 (N_17881,N_16843,N_16893);
xor U17882 (N_17882,N_17218,N_17199);
and U17883 (N_17883,N_16945,N_17223);
nor U17884 (N_17884,N_16969,N_17347);
nand U17885 (N_17885,N_17284,N_17002);
xnor U17886 (N_17886,N_17171,N_16845);
xnor U17887 (N_17887,N_16915,N_17220);
or U17888 (N_17888,N_17232,N_17293);
nor U17889 (N_17889,N_16997,N_17307);
nand U17890 (N_17890,N_17332,N_17106);
xor U17891 (N_17891,N_17002,N_17335);
nand U17892 (N_17892,N_16917,N_17275);
or U17893 (N_17893,N_17103,N_17107);
and U17894 (N_17894,N_17137,N_16803);
xor U17895 (N_17895,N_17358,N_17157);
nor U17896 (N_17896,N_17327,N_16801);
or U17897 (N_17897,N_17209,N_17233);
nor U17898 (N_17898,N_17380,N_16903);
xor U17899 (N_17899,N_16800,N_16817);
nand U17900 (N_17900,N_17333,N_17099);
nand U17901 (N_17901,N_17235,N_17227);
or U17902 (N_17902,N_17205,N_16847);
nand U17903 (N_17903,N_16906,N_17365);
nand U17904 (N_17904,N_17347,N_17391);
nor U17905 (N_17905,N_17011,N_16920);
xnor U17906 (N_17906,N_17008,N_16871);
nor U17907 (N_17907,N_17030,N_16950);
and U17908 (N_17908,N_17102,N_16813);
and U17909 (N_17909,N_16954,N_17256);
nand U17910 (N_17910,N_17164,N_17100);
nor U17911 (N_17911,N_16833,N_17019);
nand U17912 (N_17912,N_17137,N_17164);
or U17913 (N_17913,N_17158,N_17226);
xor U17914 (N_17914,N_16833,N_16937);
or U17915 (N_17915,N_16856,N_17204);
nand U17916 (N_17916,N_17392,N_17238);
or U17917 (N_17917,N_17071,N_17213);
nand U17918 (N_17918,N_17103,N_16898);
and U17919 (N_17919,N_17186,N_16890);
or U17920 (N_17920,N_17268,N_16858);
xor U17921 (N_17921,N_17172,N_17304);
or U17922 (N_17922,N_16972,N_16968);
or U17923 (N_17923,N_16906,N_16823);
nor U17924 (N_17924,N_17121,N_17250);
nand U17925 (N_17925,N_17069,N_17392);
xor U17926 (N_17926,N_17374,N_17116);
and U17927 (N_17927,N_16819,N_16874);
nand U17928 (N_17928,N_17052,N_16983);
and U17929 (N_17929,N_17249,N_16862);
or U17930 (N_17930,N_17330,N_17140);
xor U17931 (N_17931,N_17280,N_17263);
nand U17932 (N_17932,N_16833,N_17205);
and U17933 (N_17933,N_17040,N_16966);
nor U17934 (N_17934,N_17147,N_17080);
nor U17935 (N_17935,N_17303,N_16902);
nand U17936 (N_17936,N_17100,N_16948);
or U17937 (N_17937,N_16933,N_16979);
nand U17938 (N_17938,N_17301,N_16829);
nor U17939 (N_17939,N_16805,N_17376);
nand U17940 (N_17940,N_16804,N_17260);
xnor U17941 (N_17941,N_17343,N_17048);
and U17942 (N_17942,N_16978,N_17246);
or U17943 (N_17943,N_17041,N_17256);
or U17944 (N_17944,N_16906,N_17345);
nand U17945 (N_17945,N_16955,N_17069);
or U17946 (N_17946,N_16982,N_17042);
nor U17947 (N_17947,N_17057,N_17083);
xnor U17948 (N_17948,N_16887,N_17361);
nor U17949 (N_17949,N_17378,N_17101);
nand U17950 (N_17950,N_16990,N_17228);
nor U17951 (N_17951,N_17155,N_17365);
nor U17952 (N_17952,N_16838,N_16923);
or U17953 (N_17953,N_17381,N_17217);
xnor U17954 (N_17954,N_17047,N_17265);
nand U17955 (N_17955,N_17123,N_17007);
nand U17956 (N_17956,N_17052,N_16851);
nand U17957 (N_17957,N_17304,N_17131);
or U17958 (N_17958,N_17051,N_17159);
xnor U17959 (N_17959,N_17135,N_17294);
or U17960 (N_17960,N_16920,N_16913);
or U17961 (N_17961,N_16952,N_17027);
and U17962 (N_17962,N_17227,N_16929);
xnor U17963 (N_17963,N_16837,N_17096);
nand U17964 (N_17964,N_16905,N_17035);
xor U17965 (N_17965,N_17199,N_16838);
or U17966 (N_17966,N_17117,N_16864);
or U17967 (N_17967,N_17271,N_16810);
xor U17968 (N_17968,N_16881,N_17192);
and U17969 (N_17969,N_16893,N_16956);
and U17970 (N_17970,N_17174,N_17098);
nor U17971 (N_17971,N_17193,N_17272);
or U17972 (N_17972,N_16923,N_17235);
or U17973 (N_17973,N_17332,N_16816);
and U17974 (N_17974,N_16943,N_16985);
xnor U17975 (N_17975,N_17025,N_16996);
and U17976 (N_17976,N_16965,N_17211);
nand U17977 (N_17977,N_17308,N_17168);
xor U17978 (N_17978,N_17018,N_17369);
nor U17979 (N_17979,N_17084,N_16883);
or U17980 (N_17980,N_16826,N_16843);
and U17981 (N_17981,N_16924,N_17218);
or U17982 (N_17982,N_16811,N_17180);
and U17983 (N_17983,N_16972,N_17061);
xnor U17984 (N_17984,N_17133,N_16946);
xnor U17985 (N_17985,N_17087,N_17294);
nor U17986 (N_17986,N_17368,N_17274);
or U17987 (N_17987,N_17159,N_16861);
xnor U17988 (N_17988,N_17192,N_17016);
xor U17989 (N_17989,N_17365,N_17309);
and U17990 (N_17990,N_17395,N_16864);
nand U17991 (N_17991,N_17030,N_16856);
or U17992 (N_17992,N_17118,N_16829);
and U17993 (N_17993,N_16847,N_17098);
or U17994 (N_17994,N_16864,N_17174);
xor U17995 (N_17995,N_16834,N_16850);
and U17996 (N_17996,N_16943,N_17147);
nor U17997 (N_17997,N_16925,N_16971);
or U17998 (N_17998,N_16974,N_17359);
and U17999 (N_17999,N_17226,N_17054);
and U18000 (N_18000,N_17563,N_17538);
and U18001 (N_18001,N_17557,N_17794);
xor U18002 (N_18002,N_17659,N_17592);
xnor U18003 (N_18003,N_17919,N_17930);
and U18004 (N_18004,N_17999,N_17738);
and U18005 (N_18005,N_17616,N_17631);
nand U18006 (N_18006,N_17945,N_17526);
nand U18007 (N_18007,N_17862,N_17825);
and U18008 (N_18008,N_17402,N_17879);
and U18009 (N_18009,N_17482,N_17904);
and U18010 (N_18010,N_17823,N_17928);
xnor U18011 (N_18011,N_17706,N_17605);
or U18012 (N_18012,N_17829,N_17649);
and U18013 (N_18013,N_17552,N_17872);
nand U18014 (N_18014,N_17536,N_17780);
and U18015 (N_18015,N_17735,N_17569);
xor U18016 (N_18016,N_17502,N_17845);
nor U18017 (N_18017,N_17586,N_17763);
nor U18018 (N_18018,N_17899,N_17516);
nand U18019 (N_18019,N_17967,N_17558);
nor U18020 (N_18020,N_17579,N_17956);
or U18021 (N_18021,N_17600,N_17454);
xor U18022 (N_18022,N_17878,N_17813);
nand U18023 (N_18023,N_17988,N_17820);
and U18024 (N_18024,N_17549,N_17651);
and U18025 (N_18025,N_17689,N_17602);
xnor U18026 (N_18026,N_17641,N_17461);
xor U18027 (N_18027,N_17800,N_17556);
nor U18028 (N_18028,N_17969,N_17575);
xnor U18029 (N_18029,N_17601,N_17484);
nand U18030 (N_18030,N_17861,N_17693);
nand U18031 (N_18031,N_17968,N_17889);
xnor U18032 (N_18032,N_17867,N_17405);
xnor U18033 (N_18033,N_17456,N_17417);
and U18034 (N_18034,N_17920,N_17459);
nor U18035 (N_18035,N_17610,N_17770);
xor U18036 (N_18036,N_17773,N_17535);
or U18037 (N_18037,N_17871,N_17550);
xnor U18038 (N_18038,N_17881,N_17636);
and U18039 (N_18039,N_17477,N_17795);
or U18040 (N_18040,N_17804,N_17755);
or U18041 (N_18041,N_17962,N_17759);
and U18042 (N_18042,N_17849,N_17769);
nor U18043 (N_18043,N_17474,N_17634);
xnor U18044 (N_18044,N_17437,N_17814);
and U18045 (N_18045,N_17966,N_17974);
xnor U18046 (N_18046,N_17577,N_17705);
nand U18047 (N_18047,N_17870,N_17790);
or U18048 (N_18048,N_17765,N_17426);
nand U18049 (N_18049,N_17589,N_17810);
or U18050 (N_18050,N_17597,N_17985);
or U18051 (N_18051,N_17553,N_17677);
or U18052 (N_18052,N_17472,N_17764);
or U18053 (N_18053,N_17653,N_17485);
xor U18054 (N_18054,N_17448,N_17725);
and U18055 (N_18055,N_17704,N_17785);
or U18056 (N_18056,N_17548,N_17740);
or U18057 (N_18057,N_17991,N_17528);
nor U18058 (N_18058,N_17750,N_17446);
xor U18059 (N_18059,N_17913,N_17987);
xnor U18060 (N_18060,N_17938,N_17873);
xnor U18061 (N_18061,N_17854,N_17565);
nor U18062 (N_18062,N_17645,N_17452);
xnor U18063 (N_18063,N_17860,N_17890);
nor U18064 (N_18064,N_17953,N_17627);
and U18065 (N_18065,N_17533,N_17604);
and U18066 (N_18066,N_17975,N_17468);
and U18067 (N_18067,N_17445,N_17572);
and U18068 (N_18068,N_17828,N_17692);
nand U18069 (N_18069,N_17841,N_17929);
xnor U18070 (N_18070,N_17529,N_17674);
nor U18071 (N_18071,N_17582,N_17696);
xnor U18072 (N_18072,N_17722,N_17744);
xnor U18073 (N_18073,N_17702,N_17793);
xor U18074 (N_18074,N_17686,N_17590);
xor U18075 (N_18075,N_17884,N_17671);
and U18076 (N_18076,N_17858,N_17918);
or U18077 (N_18077,N_17957,N_17493);
xnor U18078 (N_18078,N_17835,N_17670);
nor U18079 (N_18079,N_17460,N_17925);
xnor U18080 (N_18080,N_17635,N_17897);
nor U18081 (N_18081,N_17965,N_17580);
xor U18082 (N_18082,N_17784,N_17505);
xor U18083 (N_18083,N_17863,N_17584);
nor U18084 (N_18084,N_17833,N_17506);
nand U18085 (N_18085,N_17831,N_17638);
nand U18086 (N_18086,N_17665,N_17737);
or U18087 (N_18087,N_17788,N_17591);
xnor U18088 (N_18088,N_17660,N_17412);
nand U18089 (N_18089,N_17707,N_17611);
or U18090 (N_18090,N_17514,N_17490);
xor U18091 (N_18091,N_17643,N_17926);
and U18092 (N_18092,N_17416,N_17699);
nor U18093 (N_18093,N_17522,N_17973);
nand U18094 (N_18094,N_17840,N_17666);
nand U18095 (N_18095,N_17779,N_17747);
nand U18096 (N_18096,N_17503,N_17910);
and U18097 (N_18097,N_17714,N_17441);
and U18098 (N_18098,N_17802,N_17466);
or U18099 (N_18099,N_17475,N_17687);
and U18100 (N_18100,N_17573,N_17719);
nand U18101 (N_18101,N_17859,N_17527);
and U18102 (N_18102,N_17422,N_17762);
nand U18103 (N_18103,N_17685,N_17712);
or U18104 (N_18104,N_17922,N_17510);
and U18105 (N_18105,N_17612,N_17663);
nor U18106 (N_18106,N_17621,N_17874);
nand U18107 (N_18107,N_17458,N_17727);
nor U18108 (N_18108,N_17546,N_17941);
nor U18109 (N_18109,N_17512,N_17955);
xnor U18110 (N_18110,N_17495,N_17467);
nand U18111 (N_18111,N_17811,N_17471);
nand U18112 (N_18112,N_17561,N_17620);
xnor U18113 (N_18113,N_17921,N_17430);
and U18114 (N_18114,N_17574,N_17530);
or U18115 (N_18115,N_17406,N_17979);
or U18116 (N_18116,N_17887,N_17730);
nor U18117 (N_18117,N_17915,N_17888);
and U18118 (N_18118,N_17568,N_17715);
xor U18119 (N_18119,N_17734,N_17494);
nor U18120 (N_18120,N_17669,N_17786);
xor U18121 (N_18121,N_17992,N_17838);
nand U18122 (N_18122,N_17729,N_17892);
nor U18123 (N_18123,N_17500,N_17542);
and U18124 (N_18124,N_17772,N_17718);
or U18125 (N_18125,N_17951,N_17853);
and U18126 (N_18126,N_17544,N_17521);
or U18127 (N_18127,N_17710,N_17809);
and U18128 (N_18128,N_17907,N_17639);
nand U18129 (N_18129,N_17632,N_17499);
or U18130 (N_18130,N_17511,N_17864);
or U18131 (N_18131,N_17935,N_17541);
nand U18132 (N_18132,N_17743,N_17911);
and U18133 (N_18133,N_17619,N_17876);
xnor U18134 (N_18134,N_17713,N_17900);
nand U18135 (N_18135,N_17761,N_17792);
or U18136 (N_18136,N_17599,N_17443);
nor U18137 (N_18137,N_17656,N_17491);
nand U18138 (N_18138,N_17637,N_17432);
nor U18139 (N_18139,N_17421,N_17807);
or U18140 (N_18140,N_17882,N_17749);
nor U18141 (N_18141,N_17944,N_17723);
xor U18142 (N_18142,N_17428,N_17980);
and U18143 (N_18143,N_17983,N_17594);
nor U18144 (N_18144,N_17690,N_17554);
or U18145 (N_18145,N_17768,N_17676);
nor U18146 (N_18146,N_17856,N_17400);
nor U18147 (N_18147,N_17698,N_17532);
nor U18148 (N_18148,N_17497,N_17865);
and U18149 (N_18149,N_17425,N_17531);
nand U18150 (N_18150,N_17776,N_17647);
and U18151 (N_18151,N_17834,N_17731);
nand U18152 (N_18152,N_17836,N_17478);
xor U18153 (N_18153,N_17682,N_17995);
nor U18154 (N_18154,N_17439,N_17673);
xnor U18155 (N_18155,N_17797,N_17436);
nor U18156 (N_18156,N_17444,N_17457);
nand U18157 (N_18157,N_17701,N_17739);
and U18158 (N_18158,N_17778,N_17893);
or U18159 (N_18159,N_17520,N_17427);
xnor U18160 (N_18160,N_17709,N_17816);
or U18161 (N_18161,N_17424,N_17782);
or U18162 (N_18162,N_17756,N_17912);
nand U18163 (N_18163,N_17751,N_17447);
and U18164 (N_18164,N_17555,N_17675);
nor U18165 (N_18165,N_17453,N_17805);
and U18166 (N_18166,N_17821,N_17423);
nand U18167 (N_18167,N_17700,N_17667);
or U18168 (N_18168,N_17551,N_17851);
nand U18169 (N_18169,N_17746,N_17917);
nand U18170 (N_18170,N_17508,N_17817);
and U18171 (N_18171,N_17924,N_17905);
xor U18172 (N_18172,N_17661,N_17517);
xnor U18173 (N_18173,N_17545,N_17684);
nor U18174 (N_18174,N_17766,N_17679);
or U18175 (N_18175,N_17562,N_17409);
or U18176 (N_18176,N_17564,N_17672);
or U18177 (N_18177,N_17606,N_17624);
xor U18178 (N_18178,N_17411,N_17964);
nand U18179 (N_18179,N_17614,N_17775);
and U18180 (N_18180,N_17808,N_17540);
nor U18181 (N_18181,N_17767,N_17509);
xnor U18182 (N_18182,N_17914,N_17681);
nand U18183 (N_18183,N_17644,N_17431);
nor U18184 (N_18184,N_17483,N_17933);
nor U18185 (N_18185,N_17523,N_17803);
or U18186 (N_18186,N_17830,N_17465);
or U18187 (N_18187,N_17891,N_17613);
or U18188 (N_18188,N_17648,N_17943);
and U18189 (N_18189,N_17642,N_17916);
or U18190 (N_18190,N_17998,N_17615);
or U18191 (N_18191,N_17986,N_17844);
xnor U18192 (N_18192,N_17691,N_17539);
or U18193 (N_18193,N_17826,N_17408);
nand U18194 (N_18194,N_17880,N_17513);
and U18195 (N_18195,N_17434,N_17440);
nand U18196 (N_18196,N_17728,N_17489);
xor U18197 (N_18197,N_17418,N_17741);
or U18198 (N_18198,N_17753,N_17822);
nand U18199 (N_18199,N_17629,N_17946);
xor U18200 (N_18200,N_17559,N_17617);
xnor U18201 (N_18201,N_17855,N_17625);
nand U18202 (N_18202,N_17976,N_17404);
nand U18203 (N_18203,N_17717,N_17898);
nor U18204 (N_18204,N_17593,N_17984);
nand U18205 (N_18205,N_17463,N_17507);
nor U18206 (N_18206,N_17479,N_17664);
nand U18207 (N_18207,N_17566,N_17748);
nand U18208 (N_18208,N_17680,N_17850);
xnor U18209 (N_18209,N_17451,N_17950);
nand U18210 (N_18210,N_17678,N_17487);
or U18211 (N_18211,N_17783,N_17996);
xor U18212 (N_18212,N_17947,N_17757);
xnor U18213 (N_18213,N_17796,N_17583);
nand U18214 (N_18214,N_17640,N_17752);
or U18215 (N_18215,N_17852,N_17883);
and U18216 (N_18216,N_17571,N_17812);
nand U18217 (N_18217,N_17997,N_17449);
nand U18218 (N_18218,N_17407,N_17414);
and U18219 (N_18219,N_17628,N_17901);
and U18220 (N_18220,N_17630,N_17952);
and U18221 (N_18221,N_17442,N_17958);
and U18222 (N_18222,N_17504,N_17476);
xor U18223 (N_18223,N_17760,N_17972);
xor U18224 (N_18224,N_17618,N_17857);
or U18225 (N_18225,N_17654,N_17724);
nand U18226 (N_18226,N_17726,N_17837);
nor U18227 (N_18227,N_17931,N_17403);
nand U18228 (N_18228,N_17819,N_17470);
xnor U18229 (N_18229,N_17877,N_17588);
nand U18230 (N_18230,N_17515,N_17971);
nor U18231 (N_18231,N_17695,N_17842);
xor U18232 (N_18232,N_17438,N_17771);
or U18233 (N_18233,N_17435,N_17906);
or U18234 (N_18234,N_17462,N_17721);
nor U18235 (N_18235,N_17868,N_17662);
nor U18236 (N_18236,N_17658,N_17777);
xor U18237 (N_18237,N_17492,N_17733);
or U18238 (N_18238,N_17596,N_17498);
xnor U18239 (N_18239,N_17801,N_17758);
xor U18240 (N_18240,N_17818,N_17622);
nor U18241 (N_18241,N_17464,N_17543);
or U18242 (N_18242,N_17708,N_17978);
xor U18243 (N_18243,N_17909,N_17537);
xnor U18244 (N_18244,N_17433,N_17595);
or U18245 (N_18245,N_17961,N_17940);
or U18246 (N_18246,N_17450,N_17413);
nand U18247 (N_18247,N_17732,N_17827);
nor U18248 (N_18248,N_17419,N_17866);
and U18249 (N_18249,N_17903,N_17895);
xor U18250 (N_18250,N_17989,N_17902);
nand U18251 (N_18251,N_17960,N_17486);
or U18252 (N_18252,N_17480,N_17815);
xnor U18253 (N_18253,N_17623,N_17798);
and U18254 (N_18254,N_17609,N_17525);
and U18255 (N_18255,N_17547,N_17993);
nor U18256 (N_18256,N_17608,N_17626);
nor U18257 (N_18257,N_17469,N_17652);
or U18258 (N_18258,N_17481,N_17774);
or U18259 (N_18259,N_17963,N_17789);
nor U18260 (N_18260,N_17455,N_17703);
nand U18261 (N_18261,N_17832,N_17581);
nor U18262 (N_18262,N_17496,N_17839);
nand U18263 (N_18263,N_17754,N_17429);
xor U18264 (N_18264,N_17587,N_17646);
and U18265 (N_18265,N_17657,N_17846);
nor U18266 (N_18266,N_17720,N_17994);
nor U18267 (N_18267,N_17875,N_17745);
nand U18268 (N_18268,N_17534,N_17942);
or U18269 (N_18269,N_17959,N_17415);
xnor U18270 (N_18270,N_17650,N_17473);
and U18271 (N_18271,N_17791,N_17567);
nand U18272 (N_18272,N_17711,N_17990);
nand U18273 (N_18273,N_17948,N_17633);
xnor U18274 (N_18274,N_17697,N_17410);
or U18275 (N_18275,N_17518,N_17716);
xor U18276 (N_18276,N_17932,N_17420);
nand U18277 (N_18277,N_17781,N_17488);
and U18278 (N_18278,N_17806,N_17578);
nor U18279 (N_18279,N_17937,N_17896);
xor U18280 (N_18280,N_17576,N_17970);
xnor U18281 (N_18281,N_17894,N_17401);
and U18282 (N_18282,N_17799,N_17570);
nand U18283 (N_18283,N_17908,N_17787);
nor U18284 (N_18284,N_17688,N_17598);
or U18285 (N_18285,N_17847,N_17923);
xor U18286 (N_18286,N_17655,N_17949);
nand U18287 (N_18287,N_17736,N_17585);
and U18288 (N_18288,N_17843,N_17560);
or U18289 (N_18289,N_17982,N_17603);
nand U18290 (N_18290,N_17977,N_17668);
nor U18291 (N_18291,N_17927,N_17848);
xnor U18292 (N_18292,N_17981,N_17869);
xnor U18293 (N_18293,N_17519,N_17501);
xnor U18294 (N_18294,N_17934,N_17683);
or U18295 (N_18295,N_17742,N_17936);
nor U18296 (N_18296,N_17954,N_17885);
or U18297 (N_18297,N_17939,N_17824);
xnor U18298 (N_18298,N_17694,N_17524);
nor U18299 (N_18299,N_17886,N_17607);
nand U18300 (N_18300,N_17817,N_17990);
and U18301 (N_18301,N_17622,N_17929);
nor U18302 (N_18302,N_17446,N_17706);
nand U18303 (N_18303,N_17955,N_17830);
or U18304 (N_18304,N_17658,N_17776);
nand U18305 (N_18305,N_17841,N_17838);
nor U18306 (N_18306,N_17440,N_17978);
xor U18307 (N_18307,N_17519,N_17537);
or U18308 (N_18308,N_17567,N_17886);
nor U18309 (N_18309,N_17523,N_17647);
or U18310 (N_18310,N_17854,N_17842);
or U18311 (N_18311,N_17598,N_17946);
nand U18312 (N_18312,N_17807,N_17411);
xor U18313 (N_18313,N_17524,N_17560);
xnor U18314 (N_18314,N_17581,N_17566);
xor U18315 (N_18315,N_17503,N_17944);
or U18316 (N_18316,N_17491,N_17838);
xor U18317 (N_18317,N_17583,N_17757);
nand U18318 (N_18318,N_17831,N_17677);
or U18319 (N_18319,N_17921,N_17547);
nor U18320 (N_18320,N_17949,N_17815);
and U18321 (N_18321,N_17406,N_17776);
nor U18322 (N_18322,N_17721,N_17522);
or U18323 (N_18323,N_17952,N_17729);
xnor U18324 (N_18324,N_17744,N_17491);
nor U18325 (N_18325,N_17430,N_17939);
nand U18326 (N_18326,N_17443,N_17999);
xnor U18327 (N_18327,N_17432,N_17931);
or U18328 (N_18328,N_17454,N_17744);
nand U18329 (N_18329,N_17656,N_17562);
xnor U18330 (N_18330,N_17651,N_17672);
nand U18331 (N_18331,N_17830,N_17404);
and U18332 (N_18332,N_17613,N_17580);
xnor U18333 (N_18333,N_17413,N_17666);
nand U18334 (N_18334,N_17787,N_17845);
xor U18335 (N_18335,N_17458,N_17438);
or U18336 (N_18336,N_17907,N_17723);
or U18337 (N_18337,N_17686,N_17841);
and U18338 (N_18338,N_17805,N_17932);
nor U18339 (N_18339,N_17504,N_17846);
or U18340 (N_18340,N_17419,N_17591);
nor U18341 (N_18341,N_17619,N_17408);
nand U18342 (N_18342,N_17630,N_17830);
nand U18343 (N_18343,N_17680,N_17507);
nand U18344 (N_18344,N_17784,N_17772);
xnor U18345 (N_18345,N_17541,N_17422);
nor U18346 (N_18346,N_17610,N_17775);
or U18347 (N_18347,N_17791,N_17608);
and U18348 (N_18348,N_17856,N_17922);
nand U18349 (N_18349,N_17511,N_17749);
and U18350 (N_18350,N_17887,N_17521);
xnor U18351 (N_18351,N_17749,N_17617);
and U18352 (N_18352,N_17552,N_17845);
xnor U18353 (N_18353,N_17495,N_17402);
xnor U18354 (N_18354,N_17498,N_17706);
nand U18355 (N_18355,N_17797,N_17734);
or U18356 (N_18356,N_17570,N_17870);
nor U18357 (N_18357,N_17945,N_17895);
or U18358 (N_18358,N_17680,N_17415);
nor U18359 (N_18359,N_17819,N_17708);
nor U18360 (N_18360,N_17866,N_17987);
and U18361 (N_18361,N_17542,N_17623);
or U18362 (N_18362,N_17692,N_17631);
xnor U18363 (N_18363,N_17694,N_17902);
and U18364 (N_18364,N_17491,N_17812);
nand U18365 (N_18365,N_17748,N_17467);
or U18366 (N_18366,N_17632,N_17740);
nand U18367 (N_18367,N_17587,N_17936);
nor U18368 (N_18368,N_17516,N_17495);
xor U18369 (N_18369,N_17781,N_17715);
nand U18370 (N_18370,N_17506,N_17515);
xor U18371 (N_18371,N_17973,N_17839);
nand U18372 (N_18372,N_17915,N_17627);
nand U18373 (N_18373,N_17652,N_17665);
xnor U18374 (N_18374,N_17850,N_17552);
and U18375 (N_18375,N_17730,N_17590);
nor U18376 (N_18376,N_17663,N_17593);
or U18377 (N_18377,N_17877,N_17828);
or U18378 (N_18378,N_17966,N_17991);
nand U18379 (N_18379,N_17665,N_17405);
nor U18380 (N_18380,N_17610,N_17763);
or U18381 (N_18381,N_17537,N_17695);
nand U18382 (N_18382,N_17957,N_17582);
nor U18383 (N_18383,N_17660,N_17434);
or U18384 (N_18384,N_17749,N_17744);
nor U18385 (N_18385,N_17595,N_17547);
or U18386 (N_18386,N_17546,N_17489);
or U18387 (N_18387,N_17987,N_17686);
and U18388 (N_18388,N_17751,N_17752);
nor U18389 (N_18389,N_17571,N_17703);
nor U18390 (N_18390,N_17593,N_17837);
xor U18391 (N_18391,N_17785,N_17939);
nor U18392 (N_18392,N_17787,N_17808);
xor U18393 (N_18393,N_17557,N_17811);
nor U18394 (N_18394,N_17722,N_17925);
nor U18395 (N_18395,N_17852,N_17592);
nand U18396 (N_18396,N_17510,N_17874);
or U18397 (N_18397,N_17541,N_17463);
and U18398 (N_18398,N_17405,N_17795);
or U18399 (N_18399,N_17563,N_17723);
nor U18400 (N_18400,N_17403,N_17632);
and U18401 (N_18401,N_17458,N_17695);
and U18402 (N_18402,N_17993,N_17567);
nand U18403 (N_18403,N_17914,N_17563);
xor U18404 (N_18404,N_17443,N_17981);
nor U18405 (N_18405,N_17796,N_17911);
nand U18406 (N_18406,N_17515,N_17445);
and U18407 (N_18407,N_17640,N_17408);
nand U18408 (N_18408,N_17964,N_17896);
nand U18409 (N_18409,N_17660,N_17568);
or U18410 (N_18410,N_17603,N_17434);
xnor U18411 (N_18411,N_17857,N_17486);
and U18412 (N_18412,N_17787,N_17900);
or U18413 (N_18413,N_17516,N_17504);
nor U18414 (N_18414,N_17488,N_17596);
nor U18415 (N_18415,N_17519,N_17893);
nor U18416 (N_18416,N_17812,N_17901);
or U18417 (N_18417,N_17844,N_17678);
or U18418 (N_18418,N_17471,N_17795);
nor U18419 (N_18419,N_17730,N_17579);
and U18420 (N_18420,N_17980,N_17786);
nor U18421 (N_18421,N_17780,N_17875);
or U18422 (N_18422,N_17975,N_17826);
nand U18423 (N_18423,N_17473,N_17907);
nor U18424 (N_18424,N_17891,N_17636);
and U18425 (N_18425,N_17860,N_17420);
xnor U18426 (N_18426,N_17620,N_17455);
xnor U18427 (N_18427,N_17816,N_17972);
or U18428 (N_18428,N_17480,N_17508);
or U18429 (N_18429,N_17518,N_17713);
xor U18430 (N_18430,N_17718,N_17871);
xnor U18431 (N_18431,N_17723,N_17955);
and U18432 (N_18432,N_17751,N_17849);
and U18433 (N_18433,N_17496,N_17581);
and U18434 (N_18434,N_17671,N_17559);
xor U18435 (N_18435,N_17877,N_17505);
nor U18436 (N_18436,N_17736,N_17806);
nand U18437 (N_18437,N_17719,N_17679);
or U18438 (N_18438,N_17611,N_17879);
and U18439 (N_18439,N_17431,N_17781);
or U18440 (N_18440,N_17547,N_17898);
xor U18441 (N_18441,N_17752,N_17714);
and U18442 (N_18442,N_17882,N_17837);
xnor U18443 (N_18443,N_17501,N_17944);
or U18444 (N_18444,N_17599,N_17863);
nor U18445 (N_18445,N_17621,N_17726);
nor U18446 (N_18446,N_17911,N_17477);
or U18447 (N_18447,N_17893,N_17818);
nor U18448 (N_18448,N_17776,N_17564);
nand U18449 (N_18449,N_17440,N_17548);
or U18450 (N_18450,N_17692,N_17696);
or U18451 (N_18451,N_17639,N_17568);
or U18452 (N_18452,N_17412,N_17538);
nor U18453 (N_18453,N_17685,N_17953);
and U18454 (N_18454,N_17440,N_17932);
nand U18455 (N_18455,N_17907,N_17809);
nand U18456 (N_18456,N_17567,N_17643);
and U18457 (N_18457,N_17606,N_17684);
and U18458 (N_18458,N_17530,N_17611);
and U18459 (N_18459,N_17824,N_17680);
or U18460 (N_18460,N_17760,N_17812);
and U18461 (N_18461,N_17631,N_17652);
nor U18462 (N_18462,N_17937,N_17873);
nor U18463 (N_18463,N_17478,N_17807);
nand U18464 (N_18464,N_17968,N_17825);
nand U18465 (N_18465,N_17935,N_17945);
and U18466 (N_18466,N_17858,N_17635);
nand U18467 (N_18467,N_17524,N_17984);
or U18468 (N_18468,N_17535,N_17599);
nor U18469 (N_18469,N_17434,N_17905);
nor U18470 (N_18470,N_17912,N_17904);
or U18471 (N_18471,N_17619,N_17674);
or U18472 (N_18472,N_17550,N_17413);
xnor U18473 (N_18473,N_17423,N_17530);
nand U18474 (N_18474,N_17550,N_17487);
xor U18475 (N_18475,N_17504,N_17485);
or U18476 (N_18476,N_17445,N_17411);
nand U18477 (N_18477,N_17929,N_17437);
nor U18478 (N_18478,N_17779,N_17566);
xor U18479 (N_18479,N_17826,N_17715);
nand U18480 (N_18480,N_17942,N_17754);
or U18481 (N_18481,N_17762,N_17503);
or U18482 (N_18482,N_17582,N_17872);
and U18483 (N_18483,N_17416,N_17991);
nor U18484 (N_18484,N_17950,N_17729);
xor U18485 (N_18485,N_17434,N_17795);
nand U18486 (N_18486,N_17466,N_17493);
and U18487 (N_18487,N_17520,N_17452);
and U18488 (N_18488,N_17661,N_17899);
nand U18489 (N_18489,N_17976,N_17442);
or U18490 (N_18490,N_17454,N_17625);
nand U18491 (N_18491,N_17999,N_17590);
or U18492 (N_18492,N_17449,N_17746);
nor U18493 (N_18493,N_17992,N_17882);
or U18494 (N_18494,N_17894,N_17875);
xnor U18495 (N_18495,N_17609,N_17844);
nor U18496 (N_18496,N_17973,N_17906);
xor U18497 (N_18497,N_17660,N_17686);
xnor U18498 (N_18498,N_17536,N_17852);
or U18499 (N_18499,N_17649,N_17786);
nor U18500 (N_18500,N_17700,N_17790);
xor U18501 (N_18501,N_17548,N_17582);
and U18502 (N_18502,N_17624,N_17912);
or U18503 (N_18503,N_17684,N_17907);
or U18504 (N_18504,N_17681,N_17954);
or U18505 (N_18505,N_17663,N_17894);
xor U18506 (N_18506,N_17653,N_17788);
or U18507 (N_18507,N_17689,N_17614);
nor U18508 (N_18508,N_17919,N_17644);
and U18509 (N_18509,N_17491,N_17792);
xor U18510 (N_18510,N_17700,N_17794);
and U18511 (N_18511,N_17878,N_17764);
or U18512 (N_18512,N_17545,N_17517);
and U18513 (N_18513,N_17836,N_17703);
xnor U18514 (N_18514,N_17824,N_17541);
nand U18515 (N_18515,N_17484,N_17875);
or U18516 (N_18516,N_17588,N_17768);
or U18517 (N_18517,N_17760,N_17433);
nor U18518 (N_18518,N_17791,N_17776);
or U18519 (N_18519,N_17973,N_17892);
or U18520 (N_18520,N_17505,N_17612);
nor U18521 (N_18521,N_17881,N_17976);
or U18522 (N_18522,N_17515,N_17464);
and U18523 (N_18523,N_17929,N_17750);
or U18524 (N_18524,N_17778,N_17552);
xnor U18525 (N_18525,N_17722,N_17875);
nor U18526 (N_18526,N_17504,N_17413);
or U18527 (N_18527,N_17842,N_17606);
and U18528 (N_18528,N_17583,N_17606);
nand U18529 (N_18529,N_17989,N_17526);
nand U18530 (N_18530,N_17945,N_17462);
and U18531 (N_18531,N_17518,N_17895);
and U18532 (N_18532,N_17578,N_17781);
nand U18533 (N_18533,N_17661,N_17604);
xor U18534 (N_18534,N_17647,N_17887);
or U18535 (N_18535,N_17836,N_17681);
xor U18536 (N_18536,N_17797,N_17518);
nand U18537 (N_18537,N_17481,N_17702);
xnor U18538 (N_18538,N_17595,N_17995);
nor U18539 (N_18539,N_17448,N_17447);
or U18540 (N_18540,N_17556,N_17451);
nand U18541 (N_18541,N_17481,N_17740);
nand U18542 (N_18542,N_17963,N_17756);
and U18543 (N_18543,N_17661,N_17420);
nor U18544 (N_18544,N_17515,N_17946);
nand U18545 (N_18545,N_17821,N_17778);
xnor U18546 (N_18546,N_17745,N_17860);
nand U18547 (N_18547,N_17557,N_17958);
nor U18548 (N_18548,N_17571,N_17429);
or U18549 (N_18549,N_17624,N_17520);
and U18550 (N_18550,N_17664,N_17743);
nand U18551 (N_18551,N_17514,N_17865);
nor U18552 (N_18552,N_17933,N_17925);
nand U18553 (N_18553,N_17943,N_17897);
and U18554 (N_18554,N_17803,N_17606);
nor U18555 (N_18555,N_17929,N_17980);
and U18556 (N_18556,N_17639,N_17602);
nor U18557 (N_18557,N_17841,N_17867);
and U18558 (N_18558,N_17562,N_17747);
and U18559 (N_18559,N_17972,N_17618);
nor U18560 (N_18560,N_17718,N_17674);
xnor U18561 (N_18561,N_17489,N_17517);
xnor U18562 (N_18562,N_17489,N_17463);
nor U18563 (N_18563,N_17958,N_17996);
and U18564 (N_18564,N_17928,N_17571);
nand U18565 (N_18565,N_17514,N_17807);
and U18566 (N_18566,N_17555,N_17845);
or U18567 (N_18567,N_17549,N_17448);
nor U18568 (N_18568,N_17647,N_17495);
or U18569 (N_18569,N_17966,N_17447);
nand U18570 (N_18570,N_17467,N_17595);
or U18571 (N_18571,N_17650,N_17993);
or U18572 (N_18572,N_17524,N_17896);
nor U18573 (N_18573,N_17619,N_17897);
nor U18574 (N_18574,N_17733,N_17746);
xor U18575 (N_18575,N_17507,N_17833);
xor U18576 (N_18576,N_17867,N_17949);
or U18577 (N_18577,N_17453,N_17488);
nand U18578 (N_18578,N_17921,N_17490);
or U18579 (N_18579,N_17588,N_17911);
or U18580 (N_18580,N_17702,N_17639);
xnor U18581 (N_18581,N_17437,N_17874);
and U18582 (N_18582,N_17677,N_17697);
nand U18583 (N_18583,N_17858,N_17713);
and U18584 (N_18584,N_17460,N_17836);
or U18585 (N_18585,N_17452,N_17590);
xnor U18586 (N_18586,N_17868,N_17798);
and U18587 (N_18587,N_17730,N_17962);
nor U18588 (N_18588,N_17708,N_17925);
and U18589 (N_18589,N_17802,N_17856);
xor U18590 (N_18590,N_17714,N_17777);
or U18591 (N_18591,N_17651,N_17907);
xnor U18592 (N_18592,N_17924,N_17411);
or U18593 (N_18593,N_17655,N_17474);
nor U18594 (N_18594,N_17557,N_17708);
xor U18595 (N_18595,N_17867,N_17901);
nand U18596 (N_18596,N_17568,N_17493);
or U18597 (N_18597,N_17675,N_17601);
or U18598 (N_18598,N_17613,N_17423);
and U18599 (N_18599,N_17583,N_17898);
nand U18600 (N_18600,N_18033,N_18449);
and U18601 (N_18601,N_18163,N_18122);
nand U18602 (N_18602,N_18203,N_18521);
nand U18603 (N_18603,N_18080,N_18433);
and U18604 (N_18604,N_18061,N_18001);
nor U18605 (N_18605,N_18127,N_18015);
xor U18606 (N_18606,N_18024,N_18316);
xor U18607 (N_18607,N_18327,N_18329);
or U18608 (N_18608,N_18592,N_18397);
and U18609 (N_18609,N_18356,N_18538);
nand U18610 (N_18610,N_18292,N_18256);
xnor U18611 (N_18611,N_18290,N_18109);
nor U18612 (N_18612,N_18529,N_18310);
nand U18613 (N_18613,N_18276,N_18293);
or U18614 (N_18614,N_18126,N_18539);
and U18615 (N_18615,N_18145,N_18053);
nand U18616 (N_18616,N_18365,N_18467);
or U18617 (N_18617,N_18005,N_18055);
and U18618 (N_18618,N_18060,N_18373);
and U18619 (N_18619,N_18110,N_18338);
and U18620 (N_18620,N_18194,N_18560);
xnor U18621 (N_18621,N_18452,N_18037);
nor U18622 (N_18622,N_18413,N_18102);
xnor U18623 (N_18623,N_18531,N_18380);
xnor U18624 (N_18624,N_18130,N_18266);
xor U18625 (N_18625,N_18402,N_18583);
nand U18626 (N_18626,N_18525,N_18099);
or U18627 (N_18627,N_18408,N_18161);
or U18628 (N_18628,N_18075,N_18275);
xnor U18629 (N_18629,N_18143,N_18027);
or U18630 (N_18630,N_18104,N_18279);
nor U18631 (N_18631,N_18546,N_18453);
xor U18632 (N_18632,N_18091,N_18299);
nand U18633 (N_18633,N_18242,N_18481);
xor U18634 (N_18634,N_18580,N_18065);
nor U18635 (N_18635,N_18274,N_18471);
and U18636 (N_18636,N_18074,N_18359);
or U18637 (N_18637,N_18556,N_18483);
xnor U18638 (N_18638,N_18106,N_18170);
and U18639 (N_18639,N_18462,N_18358);
nand U18640 (N_18640,N_18526,N_18271);
nor U18641 (N_18641,N_18087,N_18188);
and U18642 (N_18642,N_18388,N_18378);
nand U18643 (N_18643,N_18506,N_18206);
xor U18644 (N_18644,N_18247,N_18222);
or U18645 (N_18645,N_18202,N_18432);
or U18646 (N_18646,N_18362,N_18458);
xnor U18647 (N_18647,N_18002,N_18094);
or U18648 (N_18648,N_18208,N_18485);
xnor U18649 (N_18649,N_18025,N_18323);
and U18650 (N_18650,N_18023,N_18566);
xnor U18651 (N_18651,N_18088,N_18153);
nand U18652 (N_18652,N_18335,N_18003);
and U18653 (N_18653,N_18595,N_18520);
and U18654 (N_18654,N_18315,N_18178);
nand U18655 (N_18655,N_18246,N_18594);
or U18656 (N_18656,N_18308,N_18541);
and U18657 (N_18657,N_18496,N_18532);
and U18658 (N_18658,N_18133,N_18076);
and U18659 (N_18659,N_18499,N_18112);
xnor U18660 (N_18660,N_18424,N_18486);
nand U18661 (N_18661,N_18459,N_18547);
xnor U18662 (N_18662,N_18277,N_18225);
xnor U18663 (N_18663,N_18140,N_18346);
nand U18664 (N_18664,N_18073,N_18047);
or U18665 (N_18665,N_18548,N_18298);
or U18666 (N_18666,N_18146,N_18302);
nand U18667 (N_18667,N_18405,N_18326);
xor U18668 (N_18668,N_18063,N_18129);
nand U18669 (N_18669,N_18534,N_18447);
or U18670 (N_18670,N_18183,N_18192);
and U18671 (N_18671,N_18445,N_18217);
or U18672 (N_18672,N_18084,N_18083);
nand U18673 (N_18673,N_18134,N_18454);
nand U18674 (N_18674,N_18043,N_18269);
nand U18675 (N_18675,N_18333,N_18392);
nor U18676 (N_18676,N_18197,N_18281);
and U18677 (N_18677,N_18530,N_18219);
nand U18678 (N_18678,N_18574,N_18240);
nor U18679 (N_18679,N_18550,N_18351);
xnor U18680 (N_18680,N_18105,N_18597);
xor U18681 (N_18681,N_18353,N_18250);
and U18682 (N_18682,N_18064,N_18441);
and U18683 (N_18683,N_18108,N_18168);
nor U18684 (N_18684,N_18502,N_18020);
nand U18685 (N_18685,N_18051,N_18077);
or U18686 (N_18686,N_18022,N_18350);
and U18687 (N_18687,N_18295,N_18561);
xnor U18688 (N_18688,N_18337,N_18185);
or U18689 (N_18689,N_18554,N_18514);
nor U18690 (N_18690,N_18120,N_18210);
or U18691 (N_18691,N_18066,N_18165);
xnor U18692 (N_18692,N_18370,N_18488);
nand U18693 (N_18693,N_18111,N_18317);
and U18694 (N_18694,N_18420,N_18227);
nand U18695 (N_18695,N_18189,N_18142);
and U18696 (N_18696,N_18552,N_18577);
xnor U18697 (N_18697,N_18427,N_18513);
nand U18698 (N_18698,N_18394,N_18330);
xnor U18699 (N_18699,N_18576,N_18557);
or U18700 (N_18700,N_18196,N_18450);
xor U18701 (N_18701,N_18131,N_18558);
nand U18702 (N_18702,N_18321,N_18389);
and U18703 (N_18703,N_18118,N_18205);
nand U18704 (N_18704,N_18280,N_18259);
and U18705 (N_18705,N_18411,N_18400);
or U18706 (N_18706,N_18218,N_18490);
xnor U18707 (N_18707,N_18528,N_18430);
and U18708 (N_18708,N_18584,N_18429);
nor U18709 (N_18709,N_18287,N_18226);
or U18710 (N_18710,N_18573,N_18031);
nand U18711 (N_18711,N_18575,N_18213);
and U18712 (N_18712,N_18439,N_18230);
nor U18713 (N_18713,N_18193,N_18187);
xnor U18714 (N_18714,N_18119,N_18207);
xnor U18715 (N_18715,N_18423,N_18349);
nand U18716 (N_18716,N_18121,N_18578);
xnor U18717 (N_18717,N_18086,N_18512);
nor U18718 (N_18718,N_18369,N_18224);
or U18719 (N_18719,N_18428,N_18314);
nand U18720 (N_18720,N_18387,N_18419);
or U18721 (N_18721,N_18048,N_18100);
nor U18722 (N_18722,N_18278,N_18232);
nand U18723 (N_18723,N_18549,N_18085);
nand U18724 (N_18724,N_18007,N_18363);
nor U18725 (N_18725,N_18136,N_18443);
or U18726 (N_18726,N_18406,N_18044);
and U18727 (N_18727,N_18017,N_18233);
and U18728 (N_18728,N_18565,N_18011);
nor U18729 (N_18729,N_18057,N_18253);
and U18730 (N_18730,N_18303,N_18431);
nor U18731 (N_18731,N_18404,N_18535);
xor U18732 (N_18732,N_18115,N_18537);
nor U18733 (N_18733,N_18035,N_18474);
or U18734 (N_18734,N_18176,N_18154);
or U18735 (N_18735,N_18463,N_18036);
nand U18736 (N_18736,N_18200,N_18465);
nor U18737 (N_18737,N_18039,N_18345);
xor U18738 (N_18738,N_18503,N_18270);
or U18739 (N_18739,N_18562,N_18236);
or U18740 (N_18740,N_18248,N_18067);
nor U18741 (N_18741,N_18152,N_18306);
nor U18742 (N_18742,N_18181,N_18368);
or U18743 (N_18743,N_18050,N_18480);
nor U18744 (N_18744,N_18078,N_18596);
nor U18745 (N_18745,N_18089,N_18384);
nor U18746 (N_18746,N_18383,N_18564);
nand U18747 (N_18747,N_18286,N_18245);
nand U18748 (N_18748,N_18093,N_18343);
nor U18749 (N_18749,N_18010,N_18508);
nor U18750 (N_18750,N_18204,N_18177);
nand U18751 (N_18751,N_18101,N_18434);
xor U18752 (N_18752,N_18173,N_18150);
xor U18753 (N_18753,N_18252,N_18588);
nand U18754 (N_18754,N_18147,N_18386);
and U18755 (N_18755,N_18294,N_18418);
xnor U18756 (N_18756,N_18518,N_18396);
nor U18757 (N_18757,N_18331,N_18062);
xor U18758 (N_18758,N_18341,N_18399);
nand U18759 (N_18759,N_18340,N_18301);
xor U18760 (N_18760,N_18071,N_18265);
xnor U18761 (N_18761,N_18510,N_18135);
or U18762 (N_18762,N_18437,N_18385);
or U18763 (N_18763,N_18367,N_18460);
xnor U18764 (N_18764,N_18032,N_18410);
nand U18765 (N_18765,N_18466,N_18325);
or U18766 (N_18766,N_18046,N_18482);
nand U18767 (N_18767,N_18231,N_18026);
nor U18768 (N_18768,N_18138,N_18328);
and U18769 (N_18769,N_18190,N_18374);
xnor U18770 (N_18770,N_18360,N_18267);
nand U18771 (N_18771,N_18228,N_18096);
and U18772 (N_18772,N_18097,N_18004);
xor U18773 (N_18773,N_18167,N_18169);
or U18774 (N_18774,N_18174,N_18257);
and U18775 (N_18775,N_18162,N_18254);
nor U18776 (N_18776,N_18379,N_18018);
or U18777 (N_18777,N_18516,N_18235);
or U18778 (N_18778,N_18195,N_18124);
xor U18779 (N_18779,N_18484,N_18300);
xnor U18780 (N_18780,N_18008,N_18056);
nand U18781 (N_18781,N_18422,N_18555);
nor U18782 (N_18782,N_18139,N_18068);
and U18783 (N_18783,N_18371,N_18426);
nor U18784 (N_18784,N_18209,N_18241);
nand U18785 (N_18785,N_18357,N_18533);
nand U18786 (N_18786,N_18262,N_18421);
xnor U18787 (N_18787,N_18296,N_18336);
nor U18788 (N_18788,N_18137,N_18155);
or U18789 (N_18789,N_18390,N_18021);
nand U18790 (N_18790,N_18081,N_18568);
xnor U18791 (N_18791,N_18473,N_18401);
xnor U18792 (N_18792,N_18461,N_18334);
and U18793 (N_18793,N_18457,N_18570);
and U18794 (N_18794,N_18304,N_18216);
nand U18795 (N_18795,N_18059,N_18113);
and U18796 (N_18796,N_18128,N_18545);
nand U18797 (N_18797,N_18182,N_18435);
and U18798 (N_18798,N_18090,N_18523);
nand U18799 (N_18799,N_18487,N_18030);
nor U18800 (N_18800,N_18214,N_18519);
nand U18801 (N_18801,N_18491,N_18536);
or U18802 (N_18802,N_18442,N_18000);
or U18803 (N_18803,N_18366,N_18072);
nand U18804 (N_18804,N_18284,N_18238);
and U18805 (N_18805,N_18395,N_18186);
nand U18806 (N_18806,N_18464,N_18599);
nand U18807 (N_18807,N_18489,N_18339);
xnor U18808 (N_18808,N_18288,N_18220);
xnor U18809 (N_18809,N_18377,N_18261);
nand U18810 (N_18810,N_18544,N_18095);
and U18811 (N_18811,N_18103,N_18159);
xnor U18812 (N_18812,N_18149,N_18019);
and U18813 (N_18813,N_18114,N_18372);
xor U18814 (N_18814,N_18470,N_18148);
xnor U18815 (N_18815,N_18285,N_18014);
and U18816 (N_18816,N_18477,N_18311);
and U18817 (N_18817,N_18237,N_18376);
nand U18818 (N_18818,N_18313,N_18352);
or U18819 (N_18819,N_18239,N_18478);
nand U18820 (N_18820,N_18132,N_18590);
nand U18821 (N_18821,N_18157,N_18527);
and U18822 (N_18822,N_18361,N_18009);
xnor U18823 (N_18823,N_18391,N_18472);
and U18824 (N_18824,N_18319,N_18543);
nand U18825 (N_18825,N_18469,N_18409);
or U18826 (N_18826,N_18013,N_18354);
nor U18827 (N_18827,N_18006,N_18318);
nand U18828 (N_18828,N_18123,N_18289);
or U18829 (N_18829,N_18572,N_18273);
nand U18830 (N_18830,N_18492,N_18414);
nand U18831 (N_18831,N_18342,N_18455);
nor U18832 (N_18832,N_18184,N_18559);
or U18833 (N_18833,N_18355,N_18515);
nand U18834 (N_18834,N_18524,N_18542);
nor U18835 (N_18835,N_18028,N_18320);
nor U18836 (N_18836,N_18309,N_18223);
nor U18837 (N_18837,N_18347,N_18551);
nand U18838 (N_18838,N_18175,N_18272);
and U18839 (N_18839,N_18212,N_18012);
and U18840 (N_18840,N_18479,N_18511);
xnor U18841 (N_18841,N_18215,N_18540);
nor U18842 (N_18842,N_18312,N_18569);
nand U18843 (N_18843,N_18264,N_18079);
or U18844 (N_18844,N_18507,N_18070);
nand U18845 (N_18845,N_18307,N_18591);
nand U18846 (N_18846,N_18581,N_18451);
xnor U18847 (N_18847,N_18497,N_18417);
xnor U18848 (N_18848,N_18322,N_18283);
or U18849 (N_18849,N_18438,N_18058);
nor U18850 (N_18850,N_18522,N_18156);
or U18851 (N_18851,N_18517,N_18116);
xnor U18852 (N_18852,N_18416,N_18587);
xnor U18853 (N_18853,N_18364,N_18260);
nor U18854 (N_18854,N_18016,N_18598);
nand U18855 (N_18855,N_18029,N_18034);
nand U18856 (N_18856,N_18268,N_18348);
or U18857 (N_18857,N_18038,N_18191);
or U18858 (N_18858,N_18381,N_18172);
or U18859 (N_18859,N_18468,N_18049);
and U18860 (N_18860,N_18082,N_18504);
or U18861 (N_18861,N_18456,N_18098);
nor U18862 (N_18862,N_18158,N_18553);
nor U18863 (N_18863,N_18042,N_18412);
or U18864 (N_18864,N_18164,N_18249);
and U18865 (N_18865,N_18305,N_18475);
nor U18866 (N_18866,N_18052,N_18436);
nor U18867 (N_18867,N_18446,N_18344);
nand U18868 (N_18868,N_18476,N_18054);
nor U18869 (N_18869,N_18179,N_18107);
or U18870 (N_18870,N_18444,N_18493);
and U18871 (N_18871,N_18415,N_18582);
nand U18872 (N_18872,N_18234,N_18045);
or U18873 (N_18873,N_18198,N_18201);
nor U18874 (N_18874,N_18407,N_18375);
and U18875 (N_18875,N_18495,N_18180);
xnor U18876 (N_18876,N_18291,N_18498);
or U18877 (N_18877,N_18332,N_18500);
xor U18878 (N_18878,N_18282,N_18141);
xor U18879 (N_18879,N_18092,N_18398);
nand U18880 (N_18880,N_18509,N_18589);
xnor U18881 (N_18881,N_18585,N_18382);
or U18882 (N_18882,N_18501,N_18393);
or U18883 (N_18883,N_18160,N_18171);
and U18884 (N_18884,N_18505,N_18579);
and U18885 (N_18885,N_18403,N_18243);
or U18886 (N_18886,N_18151,N_18425);
nor U18887 (N_18887,N_18117,N_18586);
or U18888 (N_18888,N_18567,N_18263);
xor U18889 (N_18889,N_18563,N_18221);
nor U18890 (N_18890,N_18125,N_18324);
and U18891 (N_18891,N_18571,N_18144);
or U18892 (N_18892,N_18244,N_18041);
and U18893 (N_18893,N_18593,N_18069);
nor U18894 (N_18894,N_18211,N_18494);
nand U18895 (N_18895,N_18251,N_18258);
or U18896 (N_18896,N_18297,N_18199);
xor U18897 (N_18897,N_18166,N_18440);
nor U18898 (N_18898,N_18255,N_18448);
xnor U18899 (N_18899,N_18229,N_18040);
nand U18900 (N_18900,N_18364,N_18325);
or U18901 (N_18901,N_18460,N_18414);
nand U18902 (N_18902,N_18056,N_18593);
and U18903 (N_18903,N_18532,N_18037);
nor U18904 (N_18904,N_18592,N_18386);
nor U18905 (N_18905,N_18271,N_18277);
nor U18906 (N_18906,N_18499,N_18392);
nand U18907 (N_18907,N_18334,N_18200);
nor U18908 (N_18908,N_18333,N_18109);
and U18909 (N_18909,N_18423,N_18140);
and U18910 (N_18910,N_18150,N_18144);
and U18911 (N_18911,N_18049,N_18160);
or U18912 (N_18912,N_18218,N_18305);
nand U18913 (N_18913,N_18398,N_18107);
or U18914 (N_18914,N_18363,N_18304);
and U18915 (N_18915,N_18276,N_18058);
nor U18916 (N_18916,N_18382,N_18551);
nor U18917 (N_18917,N_18442,N_18561);
nor U18918 (N_18918,N_18575,N_18252);
or U18919 (N_18919,N_18506,N_18096);
xor U18920 (N_18920,N_18594,N_18436);
or U18921 (N_18921,N_18002,N_18013);
xnor U18922 (N_18922,N_18401,N_18115);
xor U18923 (N_18923,N_18198,N_18408);
or U18924 (N_18924,N_18026,N_18269);
or U18925 (N_18925,N_18072,N_18385);
and U18926 (N_18926,N_18048,N_18174);
or U18927 (N_18927,N_18569,N_18449);
nor U18928 (N_18928,N_18069,N_18013);
nor U18929 (N_18929,N_18053,N_18202);
nand U18930 (N_18930,N_18538,N_18474);
or U18931 (N_18931,N_18530,N_18501);
nand U18932 (N_18932,N_18035,N_18417);
nor U18933 (N_18933,N_18455,N_18294);
nand U18934 (N_18934,N_18559,N_18577);
xnor U18935 (N_18935,N_18523,N_18195);
nor U18936 (N_18936,N_18118,N_18296);
xnor U18937 (N_18937,N_18354,N_18031);
and U18938 (N_18938,N_18541,N_18591);
nor U18939 (N_18939,N_18096,N_18443);
or U18940 (N_18940,N_18327,N_18239);
nor U18941 (N_18941,N_18365,N_18039);
and U18942 (N_18942,N_18194,N_18033);
or U18943 (N_18943,N_18127,N_18513);
and U18944 (N_18944,N_18508,N_18140);
xnor U18945 (N_18945,N_18104,N_18004);
nor U18946 (N_18946,N_18346,N_18093);
nand U18947 (N_18947,N_18020,N_18368);
nor U18948 (N_18948,N_18397,N_18229);
nand U18949 (N_18949,N_18141,N_18026);
or U18950 (N_18950,N_18175,N_18007);
or U18951 (N_18951,N_18538,N_18162);
xnor U18952 (N_18952,N_18227,N_18349);
nand U18953 (N_18953,N_18466,N_18107);
nand U18954 (N_18954,N_18554,N_18337);
and U18955 (N_18955,N_18018,N_18440);
and U18956 (N_18956,N_18406,N_18242);
and U18957 (N_18957,N_18004,N_18381);
and U18958 (N_18958,N_18157,N_18023);
nand U18959 (N_18959,N_18537,N_18418);
nand U18960 (N_18960,N_18242,N_18139);
nor U18961 (N_18961,N_18317,N_18499);
nand U18962 (N_18962,N_18099,N_18022);
or U18963 (N_18963,N_18174,N_18200);
or U18964 (N_18964,N_18435,N_18084);
nand U18965 (N_18965,N_18096,N_18333);
or U18966 (N_18966,N_18422,N_18264);
and U18967 (N_18967,N_18458,N_18512);
nor U18968 (N_18968,N_18101,N_18401);
xor U18969 (N_18969,N_18345,N_18021);
nor U18970 (N_18970,N_18508,N_18087);
nor U18971 (N_18971,N_18398,N_18291);
or U18972 (N_18972,N_18201,N_18568);
or U18973 (N_18973,N_18311,N_18190);
or U18974 (N_18974,N_18118,N_18011);
xnor U18975 (N_18975,N_18572,N_18425);
nand U18976 (N_18976,N_18561,N_18006);
nand U18977 (N_18977,N_18442,N_18104);
and U18978 (N_18978,N_18419,N_18141);
xnor U18979 (N_18979,N_18270,N_18291);
nand U18980 (N_18980,N_18061,N_18136);
xnor U18981 (N_18981,N_18555,N_18278);
nand U18982 (N_18982,N_18313,N_18102);
nor U18983 (N_18983,N_18022,N_18202);
xnor U18984 (N_18984,N_18422,N_18369);
nor U18985 (N_18985,N_18095,N_18184);
or U18986 (N_18986,N_18289,N_18175);
nand U18987 (N_18987,N_18581,N_18561);
or U18988 (N_18988,N_18138,N_18063);
xor U18989 (N_18989,N_18244,N_18555);
and U18990 (N_18990,N_18024,N_18574);
and U18991 (N_18991,N_18562,N_18130);
and U18992 (N_18992,N_18351,N_18262);
xor U18993 (N_18993,N_18523,N_18251);
nand U18994 (N_18994,N_18537,N_18267);
and U18995 (N_18995,N_18061,N_18417);
nor U18996 (N_18996,N_18365,N_18242);
xor U18997 (N_18997,N_18588,N_18259);
and U18998 (N_18998,N_18091,N_18282);
or U18999 (N_18999,N_18496,N_18401);
or U19000 (N_19000,N_18070,N_18082);
or U19001 (N_19001,N_18014,N_18189);
or U19002 (N_19002,N_18544,N_18192);
nand U19003 (N_19003,N_18204,N_18327);
nand U19004 (N_19004,N_18044,N_18200);
nand U19005 (N_19005,N_18479,N_18219);
and U19006 (N_19006,N_18035,N_18299);
or U19007 (N_19007,N_18390,N_18407);
nand U19008 (N_19008,N_18369,N_18278);
nor U19009 (N_19009,N_18181,N_18358);
nand U19010 (N_19010,N_18489,N_18524);
or U19011 (N_19011,N_18379,N_18278);
or U19012 (N_19012,N_18329,N_18480);
nor U19013 (N_19013,N_18012,N_18360);
xnor U19014 (N_19014,N_18385,N_18223);
nand U19015 (N_19015,N_18109,N_18083);
nor U19016 (N_19016,N_18480,N_18063);
and U19017 (N_19017,N_18085,N_18420);
nand U19018 (N_19018,N_18080,N_18565);
nand U19019 (N_19019,N_18573,N_18478);
nand U19020 (N_19020,N_18185,N_18452);
or U19021 (N_19021,N_18175,N_18232);
nand U19022 (N_19022,N_18533,N_18405);
and U19023 (N_19023,N_18433,N_18465);
or U19024 (N_19024,N_18157,N_18014);
or U19025 (N_19025,N_18113,N_18348);
and U19026 (N_19026,N_18474,N_18055);
nor U19027 (N_19027,N_18331,N_18129);
xor U19028 (N_19028,N_18190,N_18136);
and U19029 (N_19029,N_18496,N_18403);
xor U19030 (N_19030,N_18097,N_18343);
nor U19031 (N_19031,N_18338,N_18041);
and U19032 (N_19032,N_18520,N_18139);
and U19033 (N_19033,N_18025,N_18585);
nor U19034 (N_19034,N_18237,N_18261);
nand U19035 (N_19035,N_18131,N_18185);
nor U19036 (N_19036,N_18598,N_18269);
and U19037 (N_19037,N_18196,N_18528);
nand U19038 (N_19038,N_18507,N_18251);
or U19039 (N_19039,N_18468,N_18149);
nand U19040 (N_19040,N_18340,N_18379);
nand U19041 (N_19041,N_18048,N_18073);
nand U19042 (N_19042,N_18124,N_18469);
xnor U19043 (N_19043,N_18595,N_18229);
or U19044 (N_19044,N_18256,N_18105);
and U19045 (N_19045,N_18145,N_18508);
nand U19046 (N_19046,N_18578,N_18417);
and U19047 (N_19047,N_18328,N_18473);
xor U19048 (N_19048,N_18492,N_18109);
and U19049 (N_19049,N_18016,N_18436);
xor U19050 (N_19050,N_18470,N_18522);
nand U19051 (N_19051,N_18160,N_18002);
nand U19052 (N_19052,N_18398,N_18082);
xnor U19053 (N_19053,N_18018,N_18217);
or U19054 (N_19054,N_18314,N_18223);
or U19055 (N_19055,N_18237,N_18005);
nand U19056 (N_19056,N_18349,N_18002);
and U19057 (N_19057,N_18193,N_18498);
xor U19058 (N_19058,N_18001,N_18313);
or U19059 (N_19059,N_18511,N_18173);
nor U19060 (N_19060,N_18180,N_18139);
and U19061 (N_19061,N_18277,N_18197);
nor U19062 (N_19062,N_18160,N_18211);
nand U19063 (N_19063,N_18467,N_18190);
or U19064 (N_19064,N_18184,N_18313);
and U19065 (N_19065,N_18589,N_18086);
or U19066 (N_19066,N_18349,N_18248);
nor U19067 (N_19067,N_18288,N_18517);
and U19068 (N_19068,N_18283,N_18160);
or U19069 (N_19069,N_18155,N_18563);
or U19070 (N_19070,N_18442,N_18006);
and U19071 (N_19071,N_18325,N_18223);
nand U19072 (N_19072,N_18561,N_18411);
and U19073 (N_19073,N_18477,N_18564);
or U19074 (N_19074,N_18290,N_18299);
or U19075 (N_19075,N_18057,N_18583);
and U19076 (N_19076,N_18157,N_18589);
xnor U19077 (N_19077,N_18241,N_18036);
xnor U19078 (N_19078,N_18598,N_18039);
nand U19079 (N_19079,N_18055,N_18108);
xnor U19080 (N_19080,N_18104,N_18182);
or U19081 (N_19081,N_18324,N_18020);
and U19082 (N_19082,N_18392,N_18409);
and U19083 (N_19083,N_18347,N_18198);
xor U19084 (N_19084,N_18244,N_18266);
and U19085 (N_19085,N_18160,N_18185);
or U19086 (N_19086,N_18387,N_18015);
xor U19087 (N_19087,N_18395,N_18088);
nor U19088 (N_19088,N_18116,N_18555);
nor U19089 (N_19089,N_18491,N_18473);
xnor U19090 (N_19090,N_18420,N_18465);
or U19091 (N_19091,N_18209,N_18029);
nand U19092 (N_19092,N_18195,N_18232);
and U19093 (N_19093,N_18195,N_18236);
or U19094 (N_19094,N_18006,N_18544);
or U19095 (N_19095,N_18133,N_18405);
xor U19096 (N_19096,N_18207,N_18532);
and U19097 (N_19097,N_18264,N_18491);
nor U19098 (N_19098,N_18246,N_18344);
and U19099 (N_19099,N_18384,N_18034);
nand U19100 (N_19100,N_18272,N_18123);
or U19101 (N_19101,N_18592,N_18567);
or U19102 (N_19102,N_18569,N_18069);
nand U19103 (N_19103,N_18500,N_18505);
nand U19104 (N_19104,N_18254,N_18127);
nand U19105 (N_19105,N_18287,N_18501);
nor U19106 (N_19106,N_18443,N_18467);
or U19107 (N_19107,N_18032,N_18522);
and U19108 (N_19108,N_18472,N_18580);
xor U19109 (N_19109,N_18070,N_18561);
nor U19110 (N_19110,N_18439,N_18585);
xor U19111 (N_19111,N_18497,N_18102);
nor U19112 (N_19112,N_18061,N_18159);
xnor U19113 (N_19113,N_18595,N_18581);
or U19114 (N_19114,N_18268,N_18330);
nand U19115 (N_19115,N_18395,N_18193);
nor U19116 (N_19116,N_18210,N_18246);
nand U19117 (N_19117,N_18427,N_18419);
xnor U19118 (N_19118,N_18481,N_18187);
and U19119 (N_19119,N_18300,N_18156);
nand U19120 (N_19120,N_18022,N_18514);
xor U19121 (N_19121,N_18470,N_18350);
or U19122 (N_19122,N_18420,N_18525);
nand U19123 (N_19123,N_18537,N_18257);
and U19124 (N_19124,N_18319,N_18344);
xnor U19125 (N_19125,N_18206,N_18578);
and U19126 (N_19126,N_18089,N_18319);
nor U19127 (N_19127,N_18408,N_18288);
nor U19128 (N_19128,N_18450,N_18499);
xnor U19129 (N_19129,N_18177,N_18088);
and U19130 (N_19130,N_18090,N_18047);
nor U19131 (N_19131,N_18123,N_18222);
and U19132 (N_19132,N_18113,N_18207);
and U19133 (N_19133,N_18317,N_18455);
xnor U19134 (N_19134,N_18138,N_18398);
xnor U19135 (N_19135,N_18438,N_18138);
nand U19136 (N_19136,N_18261,N_18370);
and U19137 (N_19137,N_18137,N_18340);
or U19138 (N_19138,N_18476,N_18008);
xor U19139 (N_19139,N_18444,N_18437);
or U19140 (N_19140,N_18156,N_18577);
xor U19141 (N_19141,N_18400,N_18237);
xor U19142 (N_19142,N_18455,N_18393);
nand U19143 (N_19143,N_18304,N_18116);
nor U19144 (N_19144,N_18014,N_18294);
or U19145 (N_19145,N_18440,N_18349);
xnor U19146 (N_19146,N_18023,N_18285);
and U19147 (N_19147,N_18579,N_18512);
nand U19148 (N_19148,N_18559,N_18509);
or U19149 (N_19149,N_18344,N_18407);
xor U19150 (N_19150,N_18473,N_18194);
or U19151 (N_19151,N_18331,N_18535);
nor U19152 (N_19152,N_18229,N_18059);
and U19153 (N_19153,N_18361,N_18232);
nor U19154 (N_19154,N_18209,N_18149);
xnor U19155 (N_19155,N_18065,N_18082);
xor U19156 (N_19156,N_18325,N_18509);
nor U19157 (N_19157,N_18350,N_18192);
and U19158 (N_19158,N_18325,N_18280);
nand U19159 (N_19159,N_18558,N_18000);
nand U19160 (N_19160,N_18340,N_18147);
nand U19161 (N_19161,N_18584,N_18035);
or U19162 (N_19162,N_18424,N_18173);
or U19163 (N_19163,N_18485,N_18476);
nand U19164 (N_19164,N_18119,N_18226);
nor U19165 (N_19165,N_18557,N_18519);
nor U19166 (N_19166,N_18045,N_18028);
nand U19167 (N_19167,N_18156,N_18003);
or U19168 (N_19168,N_18068,N_18318);
xnor U19169 (N_19169,N_18154,N_18271);
nor U19170 (N_19170,N_18526,N_18336);
or U19171 (N_19171,N_18023,N_18308);
xor U19172 (N_19172,N_18404,N_18491);
xor U19173 (N_19173,N_18249,N_18327);
nor U19174 (N_19174,N_18361,N_18095);
xor U19175 (N_19175,N_18115,N_18456);
or U19176 (N_19176,N_18177,N_18588);
and U19177 (N_19177,N_18045,N_18178);
nand U19178 (N_19178,N_18020,N_18342);
and U19179 (N_19179,N_18283,N_18399);
xor U19180 (N_19180,N_18569,N_18144);
nor U19181 (N_19181,N_18234,N_18512);
xor U19182 (N_19182,N_18468,N_18109);
nor U19183 (N_19183,N_18291,N_18080);
xnor U19184 (N_19184,N_18175,N_18000);
and U19185 (N_19185,N_18317,N_18585);
xnor U19186 (N_19186,N_18491,N_18416);
nand U19187 (N_19187,N_18569,N_18542);
nor U19188 (N_19188,N_18381,N_18280);
xor U19189 (N_19189,N_18369,N_18556);
nor U19190 (N_19190,N_18218,N_18452);
and U19191 (N_19191,N_18289,N_18572);
nand U19192 (N_19192,N_18044,N_18221);
or U19193 (N_19193,N_18116,N_18004);
and U19194 (N_19194,N_18223,N_18273);
xor U19195 (N_19195,N_18549,N_18080);
or U19196 (N_19196,N_18495,N_18515);
nor U19197 (N_19197,N_18458,N_18529);
nor U19198 (N_19198,N_18219,N_18164);
nor U19199 (N_19199,N_18453,N_18146);
xor U19200 (N_19200,N_19022,N_18986);
xnor U19201 (N_19201,N_18926,N_18960);
xnor U19202 (N_19202,N_19107,N_19117);
and U19203 (N_19203,N_18938,N_18876);
nand U19204 (N_19204,N_18625,N_18601);
nand U19205 (N_19205,N_18877,N_18615);
nand U19206 (N_19206,N_19021,N_18880);
xor U19207 (N_19207,N_18609,N_19180);
and U19208 (N_19208,N_18672,N_18712);
and U19209 (N_19209,N_18622,N_18697);
xor U19210 (N_19210,N_18851,N_18873);
nor U19211 (N_19211,N_19056,N_18774);
xnor U19212 (N_19212,N_19085,N_18935);
nand U19213 (N_19213,N_18908,N_19181);
or U19214 (N_19214,N_19146,N_19149);
nand U19215 (N_19215,N_18909,N_18958);
nand U19216 (N_19216,N_18830,N_19089);
xnor U19217 (N_19217,N_19077,N_18725);
and U19218 (N_19218,N_19175,N_18603);
and U19219 (N_19219,N_18997,N_18947);
xnor U19220 (N_19220,N_18983,N_19179);
nand U19221 (N_19221,N_19122,N_18741);
nor U19222 (N_19222,N_18764,N_18722);
and U19223 (N_19223,N_18789,N_18688);
xnor U19224 (N_19224,N_18889,N_19119);
nand U19225 (N_19225,N_18825,N_18927);
or U19226 (N_19226,N_19116,N_19031);
nand U19227 (N_19227,N_18823,N_19010);
nand U19228 (N_19228,N_18612,N_19118);
xnor U19229 (N_19229,N_18755,N_19113);
or U19230 (N_19230,N_18716,N_18932);
or U19231 (N_19231,N_18901,N_19019);
and U19232 (N_19232,N_18750,N_18727);
and U19233 (N_19233,N_18813,N_18811);
nand U19234 (N_19234,N_18638,N_19040);
xor U19235 (N_19235,N_19055,N_19093);
xnor U19236 (N_19236,N_18659,N_18629);
xnor U19237 (N_19237,N_18772,N_18840);
nand U19238 (N_19238,N_19133,N_19170);
and U19239 (N_19239,N_18635,N_19076);
or U19240 (N_19240,N_19034,N_19100);
nor U19241 (N_19241,N_19017,N_18858);
xnor U19242 (N_19242,N_19191,N_18956);
and U19243 (N_19243,N_18865,N_18718);
nor U19244 (N_19244,N_19008,N_18883);
xnor U19245 (N_19245,N_18757,N_18841);
xnor U19246 (N_19246,N_18870,N_18864);
nor U19247 (N_19247,N_18894,N_18801);
nand U19248 (N_19248,N_19199,N_18949);
xnor U19249 (N_19249,N_18826,N_19197);
xnor U19250 (N_19250,N_18814,N_18940);
or U19251 (N_19251,N_19104,N_19114);
xor U19252 (N_19252,N_19005,N_19079);
nor U19253 (N_19253,N_19038,N_19153);
xnor U19254 (N_19254,N_18608,N_18753);
or U19255 (N_19255,N_18793,N_18892);
nor U19256 (N_19256,N_18703,N_19087);
and U19257 (N_19257,N_18842,N_18861);
and U19258 (N_19258,N_18905,N_18992);
nor U19259 (N_19259,N_19108,N_18925);
nor U19260 (N_19260,N_19063,N_18762);
and U19261 (N_19261,N_18745,N_19189);
nor U19262 (N_19262,N_19044,N_18669);
nand U19263 (N_19263,N_18975,N_18969);
or U19264 (N_19264,N_18668,N_18748);
nand U19265 (N_19265,N_19131,N_18933);
xnor U19266 (N_19266,N_18845,N_18868);
or U19267 (N_19267,N_19082,N_19120);
nor U19268 (N_19268,N_18637,N_18856);
xnor U19269 (N_19269,N_18673,N_18756);
and U19270 (N_19270,N_18844,N_19178);
nand U19271 (N_19271,N_18639,N_18783);
nand U19272 (N_19272,N_18624,N_18995);
or U19273 (N_19273,N_19042,N_18939);
or U19274 (N_19274,N_18738,N_18924);
xor U19275 (N_19275,N_19150,N_18828);
and U19276 (N_19276,N_18666,N_19025);
xor U19277 (N_19277,N_19046,N_18963);
and U19278 (N_19278,N_19186,N_19035);
xor U19279 (N_19279,N_18994,N_19002);
xnor U19280 (N_19280,N_19177,N_18633);
xnor U19281 (N_19281,N_19184,N_18979);
xor U19282 (N_19282,N_18693,N_18686);
and U19283 (N_19283,N_19051,N_18962);
xnor U19284 (N_19284,N_19066,N_18759);
and U19285 (N_19285,N_18965,N_19103);
nand U19286 (N_19286,N_19083,N_19037);
xnor U19287 (N_19287,N_18808,N_18974);
nand U19288 (N_19288,N_18912,N_18807);
nand U19289 (N_19289,N_18928,N_18884);
or U19290 (N_19290,N_18736,N_18675);
nand U19291 (N_19291,N_18867,N_19050);
or U19292 (N_19292,N_18679,N_19172);
and U19293 (N_19293,N_18729,N_18849);
or U19294 (N_19294,N_18695,N_19090);
nor U19295 (N_19295,N_19070,N_18782);
or U19296 (N_19296,N_18677,N_19139);
nor U19297 (N_19297,N_18984,N_18667);
nor U19298 (N_19298,N_19169,N_18838);
xnor U19299 (N_19299,N_19043,N_19032);
xor U19300 (N_19300,N_18882,N_19136);
or U19301 (N_19301,N_18663,N_18816);
or U19302 (N_19302,N_18752,N_18737);
nor U19303 (N_19303,N_18735,N_18797);
xor U19304 (N_19304,N_18893,N_18773);
and U19305 (N_19305,N_18714,N_18812);
or U19306 (N_19306,N_18871,N_18904);
and U19307 (N_19307,N_18929,N_18839);
nand U19308 (N_19308,N_18780,N_18758);
xnor U19309 (N_19309,N_18690,N_18617);
nand U19310 (N_19310,N_18796,N_18670);
xnor U19311 (N_19311,N_19135,N_18618);
or U19312 (N_19312,N_18645,N_18990);
or U19313 (N_19313,N_19049,N_18616);
and U19314 (N_19314,N_18721,N_18863);
or U19315 (N_19315,N_18798,N_19143);
nor U19316 (N_19316,N_19166,N_18818);
nor U19317 (N_19317,N_19111,N_18692);
xnor U19318 (N_19318,N_18746,N_18656);
and U19319 (N_19319,N_19001,N_18785);
xor U19320 (N_19320,N_18799,N_19020);
nand U19321 (N_19321,N_19156,N_18862);
or U19322 (N_19322,N_19075,N_19144);
and U19323 (N_19323,N_19013,N_18902);
and U19324 (N_19324,N_19047,N_18857);
nand U19325 (N_19325,N_19165,N_18606);
nand U19326 (N_19326,N_18946,N_19157);
or U19327 (N_19327,N_18985,N_18600);
and U19328 (N_19328,N_18761,N_19062);
nand U19329 (N_19329,N_18848,N_18936);
and U19330 (N_19330,N_18906,N_18850);
nand U19331 (N_19331,N_18919,N_18691);
nand U19332 (N_19332,N_18653,N_18836);
nor U19333 (N_19333,N_19173,N_19195);
or U19334 (N_19334,N_19036,N_19029);
xor U19335 (N_19335,N_19171,N_19067);
and U19336 (N_19336,N_18895,N_18771);
nor U19337 (N_19337,N_19094,N_19162);
nand U19338 (N_19338,N_18847,N_18943);
xnor U19339 (N_19339,N_18972,N_18760);
xor U19340 (N_19340,N_19026,N_18646);
nand U19341 (N_19341,N_19092,N_18739);
nand U19342 (N_19342,N_18800,N_18875);
and U19343 (N_19343,N_19060,N_18696);
nand U19344 (N_19344,N_18731,N_18790);
xnor U19345 (N_19345,N_19128,N_18820);
nor U19346 (N_19346,N_19007,N_18910);
or U19347 (N_19347,N_18705,N_18605);
and U19348 (N_19348,N_19065,N_18855);
nand U19349 (N_19349,N_19106,N_19190);
xor U19350 (N_19350,N_18611,N_18959);
xor U19351 (N_19351,N_18887,N_18640);
xor U19352 (N_19352,N_18824,N_19000);
and U19353 (N_19353,N_18689,N_18993);
and U19354 (N_19354,N_18623,N_18702);
xnor U19355 (N_19355,N_18767,N_18809);
nand U19356 (N_19356,N_19145,N_18953);
xnor U19357 (N_19357,N_18632,N_19187);
nand U19358 (N_19358,N_18794,N_18636);
xor U19359 (N_19359,N_18966,N_19155);
nor U19360 (N_19360,N_19099,N_18768);
xor U19361 (N_19361,N_18916,N_18982);
xnor U19362 (N_19362,N_18957,N_19142);
or U19363 (N_19363,N_18724,N_18723);
or U19364 (N_19364,N_18896,N_18701);
nor U19365 (N_19365,N_18680,N_18879);
nor U19366 (N_19366,N_18743,N_18749);
nand U19367 (N_19367,N_18643,N_18776);
nor U19368 (N_19368,N_18674,N_18747);
or U19369 (N_19369,N_18810,N_18687);
xnor U19370 (N_19370,N_18922,N_19101);
and U19371 (N_19371,N_18654,N_18918);
nand U19372 (N_19372,N_19152,N_19112);
nor U19373 (N_19373,N_18941,N_18866);
and U19374 (N_19374,N_18833,N_18775);
and U19375 (N_19375,N_18715,N_18859);
xnor U19376 (N_19376,N_18898,N_18655);
xor U19377 (N_19377,N_19052,N_18961);
xor U19378 (N_19378,N_18754,N_18710);
nand U19379 (N_19379,N_18602,N_18971);
and U19380 (N_19380,N_18897,N_19130);
and U19381 (N_19381,N_19048,N_18977);
nand U19382 (N_19382,N_19069,N_18996);
or U19383 (N_19383,N_19097,N_18620);
xor U19384 (N_19384,N_18628,N_18931);
nor U19385 (N_19385,N_19161,N_19160);
xnor U19386 (N_19386,N_19126,N_18950);
and U19387 (N_19387,N_19059,N_18683);
and U19388 (N_19388,N_18763,N_19057);
nor U19389 (N_19389,N_19159,N_19138);
xor U19390 (N_19390,N_18854,N_18917);
and U19391 (N_19391,N_18846,N_18651);
nand U19392 (N_19392,N_18676,N_18937);
nand U19393 (N_19393,N_18817,N_19054);
nand U19394 (N_19394,N_18967,N_19086);
xor U19395 (N_19395,N_18821,N_18795);
xor U19396 (N_19396,N_18698,N_19096);
nor U19397 (N_19397,N_18834,N_18803);
and U19398 (N_19398,N_19154,N_18694);
and U19399 (N_19399,N_18742,N_18709);
xnor U19400 (N_19400,N_18744,N_19127);
or U19401 (N_19401,N_19183,N_18664);
nand U19402 (N_19402,N_18829,N_18734);
nand U19403 (N_19403,N_19023,N_18610);
or U19404 (N_19404,N_18991,N_18835);
or U19405 (N_19405,N_18787,N_18740);
and U19406 (N_19406,N_19185,N_18831);
nand U19407 (N_19407,N_18649,N_18613);
nor U19408 (N_19408,N_19098,N_18779);
nand U19409 (N_19409,N_18978,N_19061);
nor U19410 (N_19410,N_19045,N_19003);
and U19411 (N_19411,N_18976,N_19095);
nor U19412 (N_19412,N_18852,N_19134);
xnor U19413 (N_19413,N_19176,N_18837);
and U19414 (N_19414,N_18955,N_19105);
nor U19415 (N_19415,N_19132,N_19091);
nand U19416 (N_19416,N_18899,N_18678);
and U19417 (N_19417,N_18988,N_18766);
or U19418 (N_19418,N_18970,N_19004);
xnor U19419 (N_19419,N_19168,N_18815);
or U19420 (N_19420,N_19073,N_18832);
nor U19421 (N_19421,N_18660,N_18682);
and U19422 (N_19422,N_18888,N_19071);
xnor U19423 (N_19423,N_19018,N_18998);
nand U19424 (N_19424,N_18999,N_18989);
nor U19425 (N_19425,N_18920,N_18711);
nand U19426 (N_19426,N_18719,N_18923);
xor U19427 (N_19427,N_19115,N_18619);
nor U19428 (N_19428,N_18872,N_19198);
nand U19429 (N_19429,N_19121,N_18614);
xnor U19430 (N_19430,N_18650,N_18641);
xnor U19431 (N_19431,N_18886,N_18732);
nand U19432 (N_19432,N_18822,N_18630);
xnor U19433 (N_19433,N_19009,N_18942);
xnor U19434 (N_19434,N_18903,N_18805);
nor U19435 (N_19435,N_18874,N_18642);
and U19436 (N_19436,N_18827,N_19006);
and U19437 (N_19437,N_18981,N_18900);
and U19438 (N_19438,N_19078,N_19058);
nor U19439 (N_19439,N_18802,N_19102);
nand U19440 (N_19440,N_18778,N_18913);
and U19441 (N_19441,N_19072,N_18707);
nor U19442 (N_19442,N_19147,N_18648);
nand U19443 (N_19443,N_18765,N_18791);
and U19444 (N_19444,N_18915,N_19140);
xnor U19445 (N_19445,N_18708,N_18786);
xnor U19446 (N_19446,N_18968,N_18973);
nand U19447 (N_19447,N_19033,N_19081);
nor U19448 (N_19448,N_18885,N_19027);
nand U19449 (N_19449,N_18964,N_19163);
nor U19450 (N_19450,N_18730,N_18784);
or U19451 (N_19451,N_18781,N_19011);
xnor U19452 (N_19452,N_18626,N_19164);
or U19453 (N_19453,N_18921,N_19012);
and U19454 (N_19454,N_18671,N_19039);
xor U19455 (N_19455,N_18860,N_19014);
or U19456 (N_19456,N_18788,N_19110);
xor U19457 (N_19457,N_18945,N_18804);
and U19458 (N_19458,N_19196,N_18881);
nand U19459 (N_19459,N_18607,N_18728);
xnor U19460 (N_19460,N_18685,N_19041);
nor U19461 (N_19461,N_18770,N_18713);
nor U19462 (N_19462,N_19030,N_18657);
nor U19463 (N_19463,N_19174,N_18684);
and U19464 (N_19464,N_19024,N_18658);
and U19465 (N_19465,N_18751,N_19151);
and U19466 (N_19466,N_19123,N_18891);
and U19467 (N_19467,N_19028,N_19016);
and U19468 (N_19468,N_18644,N_19141);
nor U19469 (N_19469,N_19148,N_18726);
nand U19470 (N_19470,N_18717,N_19158);
nand U19471 (N_19471,N_18954,N_19124);
xor U19472 (N_19472,N_18720,N_19192);
xor U19473 (N_19473,N_18733,N_18634);
nor U19474 (N_19474,N_19088,N_18952);
nand U19475 (N_19475,N_18853,N_19080);
xnor U19476 (N_19476,N_18914,N_18647);
or U19477 (N_19477,N_18911,N_18951);
nand U19478 (N_19478,N_18890,N_19137);
xnor U19479 (N_19479,N_18604,N_18878);
xor U19480 (N_19480,N_18652,N_18792);
xor U19481 (N_19481,N_19074,N_18699);
xnor U19482 (N_19482,N_18944,N_18627);
xnor U19483 (N_19483,N_18930,N_19188);
xnor U19484 (N_19484,N_19182,N_18706);
and U19485 (N_19485,N_18704,N_18662);
or U19486 (N_19486,N_18806,N_19015);
xor U19487 (N_19487,N_18769,N_19167);
or U19488 (N_19488,N_19125,N_18700);
nor U19489 (N_19489,N_18843,N_19193);
xnor U19490 (N_19490,N_19129,N_18681);
nand U19491 (N_19491,N_18631,N_18987);
and U19492 (N_19492,N_19109,N_18907);
nand U19493 (N_19493,N_18665,N_18819);
nand U19494 (N_19494,N_18661,N_18777);
or U19495 (N_19495,N_18621,N_18980);
nand U19496 (N_19496,N_18948,N_18934);
and U19497 (N_19497,N_19084,N_19064);
nor U19498 (N_19498,N_19194,N_19068);
or U19499 (N_19499,N_18869,N_19053);
nor U19500 (N_19500,N_18928,N_18780);
nor U19501 (N_19501,N_18935,N_18721);
and U19502 (N_19502,N_18894,N_19013);
and U19503 (N_19503,N_18948,N_18737);
or U19504 (N_19504,N_18754,N_19141);
xnor U19505 (N_19505,N_18831,N_19120);
xnor U19506 (N_19506,N_18616,N_18940);
or U19507 (N_19507,N_18913,N_19154);
nor U19508 (N_19508,N_19115,N_19094);
and U19509 (N_19509,N_18726,N_18661);
nand U19510 (N_19510,N_18718,N_18710);
or U19511 (N_19511,N_18959,N_19023);
and U19512 (N_19512,N_19061,N_18878);
and U19513 (N_19513,N_18962,N_18874);
or U19514 (N_19514,N_18860,N_18853);
nand U19515 (N_19515,N_18960,N_19049);
nand U19516 (N_19516,N_19092,N_18870);
and U19517 (N_19517,N_19012,N_18897);
or U19518 (N_19518,N_19053,N_18743);
or U19519 (N_19519,N_19139,N_18903);
xor U19520 (N_19520,N_18673,N_19055);
and U19521 (N_19521,N_18981,N_18809);
xnor U19522 (N_19522,N_18992,N_18851);
xnor U19523 (N_19523,N_19119,N_18784);
or U19524 (N_19524,N_18845,N_19076);
and U19525 (N_19525,N_18919,N_19011);
and U19526 (N_19526,N_19004,N_19151);
or U19527 (N_19527,N_18641,N_18613);
or U19528 (N_19528,N_19039,N_19062);
or U19529 (N_19529,N_19164,N_19141);
nand U19530 (N_19530,N_18967,N_19143);
xnor U19531 (N_19531,N_19024,N_19003);
nor U19532 (N_19532,N_19030,N_19129);
or U19533 (N_19533,N_19080,N_18810);
nand U19534 (N_19534,N_18769,N_19076);
nor U19535 (N_19535,N_18926,N_18733);
or U19536 (N_19536,N_19082,N_18968);
or U19537 (N_19537,N_18912,N_18628);
nand U19538 (N_19538,N_18813,N_18885);
xnor U19539 (N_19539,N_18909,N_18697);
xnor U19540 (N_19540,N_18916,N_18867);
or U19541 (N_19541,N_18819,N_18611);
and U19542 (N_19542,N_19160,N_18727);
nand U19543 (N_19543,N_18851,N_18779);
nand U19544 (N_19544,N_19118,N_18809);
xnor U19545 (N_19545,N_18925,N_18997);
xor U19546 (N_19546,N_19185,N_18799);
or U19547 (N_19547,N_18989,N_18722);
nand U19548 (N_19548,N_18627,N_19152);
nand U19549 (N_19549,N_18910,N_18773);
and U19550 (N_19550,N_18952,N_18656);
nand U19551 (N_19551,N_18682,N_19019);
xnor U19552 (N_19552,N_18700,N_18783);
and U19553 (N_19553,N_18980,N_18958);
or U19554 (N_19554,N_19002,N_18843);
and U19555 (N_19555,N_19106,N_18629);
or U19556 (N_19556,N_18835,N_18914);
nand U19557 (N_19557,N_18841,N_18801);
xor U19558 (N_19558,N_19032,N_18613);
xor U19559 (N_19559,N_18884,N_18860);
and U19560 (N_19560,N_19138,N_19130);
nand U19561 (N_19561,N_18859,N_19045);
xor U19562 (N_19562,N_19150,N_18926);
xnor U19563 (N_19563,N_18689,N_19053);
nor U19564 (N_19564,N_18688,N_18650);
nand U19565 (N_19565,N_19055,N_18826);
nand U19566 (N_19566,N_18985,N_19137);
and U19567 (N_19567,N_19165,N_18984);
xor U19568 (N_19568,N_19148,N_19196);
xor U19569 (N_19569,N_18942,N_18754);
xnor U19570 (N_19570,N_19101,N_19151);
nand U19571 (N_19571,N_18789,N_19065);
xor U19572 (N_19572,N_19039,N_18902);
and U19573 (N_19573,N_18633,N_18654);
or U19574 (N_19574,N_18626,N_18789);
and U19575 (N_19575,N_18728,N_18729);
xor U19576 (N_19576,N_19012,N_18987);
xor U19577 (N_19577,N_18672,N_18863);
xor U19578 (N_19578,N_18737,N_19168);
xnor U19579 (N_19579,N_19142,N_19131);
nand U19580 (N_19580,N_19065,N_18602);
nor U19581 (N_19581,N_18868,N_18830);
nor U19582 (N_19582,N_18975,N_18652);
nand U19583 (N_19583,N_18659,N_18669);
and U19584 (N_19584,N_18716,N_18788);
xnor U19585 (N_19585,N_19021,N_19181);
or U19586 (N_19586,N_18730,N_18937);
nand U19587 (N_19587,N_19064,N_19059);
and U19588 (N_19588,N_19141,N_18890);
nand U19589 (N_19589,N_18728,N_18805);
and U19590 (N_19590,N_19009,N_18906);
or U19591 (N_19591,N_18633,N_19180);
nor U19592 (N_19592,N_18974,N_19178);
and U19593 (N_19593,N_19064,N_19024);
nand U19594 (N_19594,N_18861,N_18884);
or U19595 (N_19595,N_18626,N_18641);
or U19596 (N_19596,N_18696,N_19103);
and U19597 (N_19597,N_18808,N_18908);
xor U19598 (N_19598,N_19149,N_18734);
xnor U19599 (N_19599,N_18652,N_19130);
or U19600 (N_19600,N_18617,N_19195);
xnor U19601 (N_19601,N_18637,N_18730);
xor U19602 (N_19602,N_19074,N_18872);
nand U19603 (N_19603,N_19009,N_18797);
or U19604 (N_19604,N_18794,N_18840);
and U19605 (N_19605,N_18623,N_19082);
nand U19606 (N_19606,N_19028,N_18777);
xnor U19607 (N_19607,N_18701,N_18852);
nand U19608 (N_19608,N_18871,N_18761);
nor U19609 (N_19609,N_19164,N_18618);
nor U19610 (N_19610,N_19037,N_18924);
nor U19611 (N_19611,N_19059,N_18947);
and U19612 (N_19612,N_19124,N_18981);
nand U19613 (N_19613,N_18785,N_18936);
nor U19614 (N_19614,N_19132,N_18658);
or U19615 (N_19615,N_18668,N_18604);
and U19616 (N_19616,N_18855,N_18609);
nand U19617 (N_19617,N_18770,N_19108);
xnor U19618 (N_19618,N_18933,N_19096);
or U19619 (N_19619,N_19187,N_18615);
nor U19620 (N_19620,N_18800,N_19182);
nor U19621 (N_19621,N_18850,N_19035);
and U19622 (N_19622,N_19166,N_18938);
xor U19623 (N_19623,N_18957,N_18834);
or U19624 (N_19624,N_18995,N_18938);
and U19625 (N_19625,N_18873,N_19130);
and U19626 (N_19626,N_19006,N_18658);
nor U19627 (N_19627,N_18881,N_18670);
nand U19628 (N_19628,N_18613,N_19019);
and U19629 (N_19629,N_18745,N_18646);
nor U19630 (N_19630,N_18637,N_18862);
or U19631 (N_19631,N_19079,N_18763);
xor U19632 (N_19632,N_19123,N_18911);
nor U19633 (N_19633,N_18957,N_19176);
or U19634 (N_19634,N_19145,N_18632);
and U19635 (N_19635,N_18798,N_18877);
xnor U19636 (N_19636,N_18876,N_19188);
nor U19637 (N_19637,N_19061,N_18667);
and U19638 (N_19638,N_18817,N_18757);
and U19639 (N_19639,N_19126,N_18665);
nand U19640 (N_19640,N_18931,N_18721);
or U19641 (N_19641,N_18674,N_19041);
or U19642 (N_19642,N_18971,N_18681);
nand U19643 (N_19643,N_19120,N_18667);
nand U19644 (N_19644,N_18642,N_18821);
nor U19645 (N_19645,N_19111,N_19151);
and U19646 (N_19646,N_19009,N_19158);
or U19647 (N_19647,N_19182,N_18837);
nand U19648 (N_19648,N_19099,N_18657);
xnor U19649 (N_19649,N_18949,N_19196);
or U19650 (N_19650,N_18691,N_18840);
nand U19651 (N_19651,N_18970,N_19100);
and U19652 (N_19652,N_19081,N_19068);
or U19653 (N_19653,N_18769,N_18800);
xnor U19654 (N_19654,N_19031,N_18979);
or U19655 (N_19655,N_19136,N_18778);
or U19656 (N_19656,N_18641,N_18700);
nor U19657 (N_19657,N_19170,N_18678);
and U19658 (N_19658,N_19183,N_18815);
xor U19659 (N_19659,N_19158,N_18975);
and U19660 (N_19660,N_18698,N_18998);
nand U19661 (N_19661,N_18929,N_19149);
xnor U19662 (N_19662,N_18824,N_18696);
or U19663 (N_19663,N_18863,N_18626);
or U19664 (N_19664,N_18820,N_18638);
nand U19665 (N_19665,N_19063,N_19026);
xnor U19666 (N_19666,N_18632,N_19136);
nand U19667 (N_19667,N_18874,N_18992);
and U19668 (N_19668,N_18817,N_18919);
xnor U19669 (N_19669,N_19004,N_19080);
or U19670 (N_19670,N_18898,N_18658);
and U19671 (N_19671,N_18694,N_18990);
nor U19672 (N_19672,N_19129,N_19152);
nor U19673 (N_19673,N_18688,N_18868);
and U19674 (N_19674,N_18844,N_19125);
and U19675 (N_19675,N_19002,N_18744);
nor U19676 (N_19676,N_18840,N_18722);
nand U19677 (N_19677,N_19015,N_18814);
or U19678 (N_19678,N_19000,N_19086);
nand U19679 (N_19679,N_19090,N_18751);
and U19680 (N_19680,N_19031,N_19106);
nand U19681 (N_19681,N_19157,N_19056);
nand U19682 (N_19682,N_19189,N_19120);
xnor U19683 (N_19683,N_18866,N_19011);
and U19684 (N_19684,N_18844,N_18750);
nand U19685 (N_19685,N_18909,N_18946);
nand U19686 (N_19686,N_18959,N_18659);
or U19687 (N_19687,N_18686,N_18903);
xor U19688 (N_19688,N_18781,N_18768);
xnor U19689 (N_19689,N_19123,N_18688);
nor U19690 (N_19690,N_18753,N_18748);
nor U19691 (N_19691,N_18673,N_18946);
nor U19692 (N_19692,N_18890,N_18916);
xor U19693 (N_19693,N_18882,N_18724);
and U19694 (N_19694,N_18895,N_19188);
or U19695 (N_19695,N_18924,N_19043);
or U19696 (N_19696,N_18989,N_18788);
xor U19697 (N_19697,N_18671,N_19162);
nor U19698 (N_19698,N_18658,N_19000);
nand U19699 (N_19699,N_19129,N_18737);
and U19700 (N_19700,N_18846,N_19074);
nor U19701 (N_19701,N_18740,N_18614);
nand U19702 (N_19702,N_18882,N_18966);
nor U19703 (N_19703,N_19004,N_18824);
nand U19704 (N_19704,N_18864,N_18732);
nand U19705 (N_19705,N_19189,N_18947);
xor U19706 (N_19706,N_19007,N_18688);
xor U19707 (N_19707,N_19189,N_18964);
nand U19708 (N_19708,N_19103,N_19169);
or U19709 (N_19709,N_19031,N_18920);
and U19710 (N_19710,N_18810,N_18625);
nor U19711 (N_19711,N_18956,N_19156);
and U19712 (N_19712,N_18866,N_18769);
or U19713 (N_19713,N_19006,N_19063);
or U19714 (N_19714,N_19137,N_18970);
or U19715 (N_19715,N_19051,N_18990);
nor U19716 (N_19716,N_18732,N_18776);
xor U19717 (N_19717,N_18688,N_19058);
xnor U19718 (N_19718,N_19015,N_18970);
nand U19719 (N_19719,N_19056,N_19184);
nor U19720 (N_19720,N_19159,N_18874);
or U19721 (N_19721,N_19196,N_18973);
or U19722 (N_19722,N_19129,N_18768);
and U19723 (N_19723,N_19139,N_18806);
xnor U19724 (N_19724,N_18884,N_18612);
or U19725 (N_19725,N_18733,N_18809);
or U19726 (N_19726,N_18606,N_18882);
xnor U19727 (N_19727,N_19039,N_18874);
nor U19728 (N_19728,N_19192,N_19037);
xnor U19729 (N_19729,N_19140,N_18757);
xnor U19730 (N_19730,N_18663,N_18640);
xnor U19731 (N_19731,N_19064,N_19134);
and U19732 (N_19732,N_18697,N_18961);
nor U19733 (N_19733,N_18883,N_18705);
nor U19734 (N_19734,N_18730,N_18815);
nor U19735 (N_19735,N_18816,N_19183);
or U19736 (N_19736,N_18970,N_19169);
or U19737 (N_19737,N_19190,N_18927);
nor U19738 (N_19738,N_18993,N_19159);
or U19739 (N_19739,N_18602,N_18720);
nor U19740 (N_19740,N_18885,N_19192);
nor U19741 (N_19741,N_18648,N_18884);
nand U19742 (N_19742,N_18912,N_19078);
and U19743 (N_19743,N_18678,N_18636);
nand U19744 (N_19744,N_19128,N_19126);
nor U19745 (N_19745,N_18745,N_18960);
nor U19746 (N_19746,N_18605,N_18855);
nor U19747 (N_19747,N_18937,N_18819);
nand U19748 (N_19748,N_19151,N_18681);
nor U19749 (N_19749,N_18649,N_18779);
or U19750 (N_19750,N_19038,N_19059);
nand U19751 (N_19751,N_18912,N_18865);
nor U19752 (N_19752,N_18960,N_19105);
nor U19753 (N_19753,N_19102,N_18784);
and U19754 (N_19754,N_19005,N_18938);
and U19755 (N_19755,N_19046,N_18848);
or U19756 (N_19756,N_19055,N_19185);
nand U19757 (N_19757,N_18875,N_18950);
xor U19758 (N_19758,N_19081,N_19182);
xor U19759 (N_19759,N_18610,N_18735);
nor U19760 (N_19760,N_19046,N_19189);
and U19761 (N_19761,N_19023,N_19033);
nor U19762 (N_19762,N_19183,N_19039);
or U19763 (N_19763,N_18763,N_19002);
or U19764 (N_19764,N_18738,N_19137);
nor U19765 (N_19765,N_18699,N_19126);
nor U19766 (N_19766,N_19004,N_19026);
or U19767 (N_19767,N_19179,N_18749);
and U19768 (N_19768,N_18684,N_18835);
and U19769 (N_19769,N_18801,N_18674);
or U19770 (N_19770,N_19007,N_18917);
nand U19771 (N_19771,N_18992,N_19063);
nand U19772 (N_19772,N_18787,N_18763);
or U19773 (N_19773,N_18882,N_18609);
nor U19774 (N_19774,N_19016,N_19092);
nand U19775 (N_19775,N_19120,N_18782);
and U19776 (N_19776,N_19061,N_19054);
nand U19777 (N_19777,N_18971,N_18911);
nor U19778 (N_19778,N_19154,N_19146);
xnor U19779 (N_19779,N_19005,N_18788);
and U19780 (N_19780,N_18803,N_18680);
nand U19781 (N_19781,N_18659,N_18887);
and U19782 (N_19782,N_18896,N_18923);
nand U19783 (N_19783,N_19097,N_19150);
nand U19784 (N_19784,N_18918,N_18639);
or U19785 (N_19785,N_18714,N_18752);
xor U19786 (N_19786,N_18693,N_19059);
or U19787 (N_19787,N_19080,N_18619);
nand U19788 (N_19788,N_18790,N_18810);
nand U19789 (N_19789,N_19057,N_18874);
and U19790 (N_19790,N_18692,N_18755);
and U19791 (N_19791,N_18686,N_19157);
nand U19792 (N_19792,N_18976,N_18988);
and U19793 (N_19793,N_19149,N_19166);
nor U19794 (N_19794,N_19138,N_18794);
nand U19795 (N_19795,N_18620,N_19174);
nand U19796 (N_19796,N_18695,N_18832);
xor U19797 (N_19797,N_18974,N_18809);
nand U19798 (N_19798,N_18914,N_18859);
or U19799 (N_19799,N_18859,N_18875);
or U19800 (N_19800,N_19267,N_19674);
nor U19801 (N_19801,N_19422,N_19552);
or U19802 (N_19802,N_19771,N_19598);
nand U19803 (N_19803,N_19283,N_19512);
or U19804 (N_19804,N_19276,N_19209);
nand U19805 (N_19805,N_19466,N_19420);
or U19806 (N_19806,N_19444,N_19502);
or U19807 (N_19807,N_19590,N_19456);
or U19808 (N_19808,N_19718,N_19449);
xor U19809 (N_19809,N_19204,N_19599);
nor U19810 (N_19810,N_19462,N_19404);
nor U19811 (N_19811,N_19406,N_19323);
nand U19812 (N_19812,N_19364,N_19604);
or U19813 (N_19813,N_19287,N_19421);
and U19814 (N_19814,N_19366,N_19586);
xnor U19815 (N_19815,N_19705,N_19752);
and U19816 (N_19816,N_19577,N_19378);
or U19817 (N_19817,N_19351,N_19787);
or U19818 (N_19818,N_19260,N_19355);
nor U19819 (N_19819,N_19201,N_19247);
nand U19820 (N_19820,N_19435,N_19282);
xnor U19821 (N_19821,N_19682,N_19678);
nand U19822 (N_19822,N_19263,N_19239);
nand U19823 (N_19823,N_19333,N_19438);
nor U19824 (N_19824,N_19491,N_19337);
nand U19825 (N_19825,N_19311,N_19402);
or U19826 (N_19826,N_19521,N_19547);
nand U19827 (N_19827,N_19386,N_19341);
nor U19828 (N_19828,N_19332,N_19517);
nor U19829 (N_19829,N_19373,N_19579);
xnor U19830 (N_19830,N_19660,N_19764);
and U19831 (N_19831,N_19496,N_19472);
or U19832 (N_19832,N_19501,N_19321);
and U19833 (N_19833,N_19785,N_19264);
and U19834 (N_19834,N_19725,N_19277);
xor U19835 (N_19835,N_19707,N_19289);
nand U19836 (N_19836,N_19451,N_19743);
nor U19837 (N_19837,N_19668,N_19279);
xor U19838 (N_19838,N_19687,N_19303);
and U19839 (N_19839,N_19436,N_19683);
or U19840 (N_19840,N_19256,N_19470);
and U19841 (N_19841,N_19381,N_19253);
and U19842 (N_19842,N_19508,N_19412);
nand U19843 (N_19843,N_19790,N_19442);
nand U19844 (N_19844,N_19214,N_19680);
or U19845 (N_19845,N_19701,N_19588);
and U19846 (N_19846,N_19222,N_19580);
nand U19847 (N_19847,N_19739,N_19597);
nor U19848 (N_19848,N_19249,N_19748);
or U19849 (N_19849,N_19257,N_19477);
nand U19850 (N_19850,N_19629,N_19644);
nor U19851 (N_19851,N_19592,N_19403);
or U19852 (N_19852,N_19711,N_19266);
xor U19853 (N_19853,N_19713,N_19318);
nor U19854 (N_19854,N_19285,N_19493);
nand U19855 (N_19855,N_19657,N_19555);
nand U19856 (N_19856,N_19231,N_19347);
or U19857 (N_19857,N_19626,N_19760);
nor U19858 (N_19858,N_19419,N_19716);
or U19859 (N_19859,N_19518,N_19464);
nand U19860 (N_19860,N_19797,N_19335);
and U19861 (N_19861,N_19269,N_19542);
or U19862 (N_19862,N_19226,N_19227);
nor U19863 (N_19863,N_19389,N_19284);
xnor U19864 (N_19864,N_19609,N_19791);
and U19865 (N_19865,N_19394,N_19677);
nand U19866 (N_19866,N_19543,N_19712);
nor U19867 (N_19867,N_19538,N_19476);
nand U19868 (N_19868,N_19544,N_19516);
xnor U19869 (N_19869,N_19327,N_19439);
nand U19870 (N_19870,N_19654,N_19245);
nor U19871 (N_19871,N_19407,N_19241);
xnor U19872 (N_19872,N_19563,N_19324);
nand U19873 (N_19873,N_19640,N_19693);
or U19874 (N_19874,N_19726,N_19280);
and U19875 (N_19875,N_19469,N_19221);
nor U19876 (N_19876,N_19423,N_19430);
and U19877 (N_19877,N_19288,N_19583);
nor U19878 (N_19878,N_19417,N_19489);
xnor U19879 (N_19879,N_19755,N_19754);
nand U19880 (N_19880,N_19229,N_19663);
nand U19881 (N_19881,N_19425,N_19675);
and U19882 (N_19882,N_19672,N_19584);
and U19883 (N_19883,N_19702,N_19409);
or U19884 (N_19884,N_19769,N_19643);
xor U19885 (N_19885,N_19623,N_19782);
and U19886 (N_19886,N_19740,N_19559);
xor U19887 (N_19887,N_19673,N_19789);
nand U19888 (N_19888,N_19238,N_19618);
nor U19889 (N_19889,N_19515,N_19714);
xor U19890 (N_19890,N_19399,N_19310);
or U19891 (N_19891,N_19520,N_19569);
or U19892 (N_19892,N_19688,N_19433);
nor U19893 (N_19893,N_19639,N_19459);
and U19894 (N_19894,N_19709,N_19322);
nor U19895 (N_19895,N_19610,N_19786);
and U19896 (N_19896,N_19776,N_19465);
xnor U19897 (N_19897,N_19453,N_19727);
nor U19898 (N_19898,N_19205,N_19655);
xnor U19899 (N_19899,N_19628,N_19642);
nand U19900 (N_19900,N_19443,N_19391);
and U19901 (N_19901,N_19374,N_19645);
nand U19902 (N_19902,N_19360,N_19292);
or U19903 (N_19903,N_19703,N_19486);
and U19904 (N_19904,N_19262,N_19593);
xnor U19905 (N_19905,N_19298,N_19418);
nand U19906 (N_19906,N_19715,N_19622);
nor U19907 (N_19907,N_19634,N_19594);
or U19908 (N_19908,N_19549,N_19211);
and U19909 (N_19909,N_19525,N_19281);
and U19910 (N_19910,N_19777,N_19255);
xor U19911 (N_19911,N_19363,N_19385);
nor U19912 (N_19912,N_19788,N_19390);
and U19913 (N_19913,N_19568,N_19710);
or U19914 (N_19914,N_19372,N_19499);
and U19915 (N_19915,N_19473,N_19601);
xor U19916 (N_19916,N_19218,N_19296);
and U19917 (N_19917,N_19684,N_19573);
and U19918 (N_19918,N_19796,N_19766);
xor U19919 (N_19919,N_19414,N_19763);
nor U19920 (N_19920,N_19638,N_19736);
xnor U19921 (N_19921,N_19582,N_19474);
or U19922 (N_19922,N_19536,N_19234);
and U19923 (N_19923,N_19210,N_19509);
and U19924 (N_19924,N_19306,N_19745);
nand U19925 (N_19925,N_19550,N_19452);
nor U19926 (N_19926,N_19546,N_19614);
or U19927 (N_19927,N_19700,N_19557);
nor U19928 (N_19928,N_19564,N_19494);
xor U19929 (N_19929,N_19387,N_19367);
nand U19930 (N_19930,N_19503,N_19375);
nor U19931 (N_19931,N_19571,N_19778);
xor U19932 (N_19932,N_19230,N_19772);
or U19933 (N_19933,N_19649,N_19779);
nand U19934 (N_19934,N_19336,N_19307);
xor U19935 (N_19935,N_19428,N_19242);
nand U19936 (N_19936,N_19291,N_19780);
nor U19937 (N_19937,N_19762,N_19290);
xor U19938 (N_19938,N_19728,N_19250);
xor U19939 (N_19939,N_19723,N_19319);
and U19940 (N_19940,N_19330,N_19765);
nor U19941 (N_19941,N_19699,N_19434);
nand U19942 (N_19942,N_19671,N_19349);
xnor U19943 (N_19943,N_19431,N_19560);
or U19944 (N_19944,N_19539,N_19455);
nor U19945 (N_19945,N_19795,N_19567);
xnor U19946 (N_19946,N_19395,N_19696);
and U19947 (N_19947,N_19488,N_19630);
and U19948 (N_19948,N_19596,N_19408);
xor U19949 (N_19949,N_19342,N_19405);
or U19950 (N_19950,N_19468,N_19556);
or U19951 (N_19951,N_19708,N_19565);
and U19952 (N_19952,N_19737,N_19799);
and U19953 (N_19953,N_19270,N_19664);
and U19954 (N_19954,N_19382,N_19357);
and U19955 (N_19955,N_19460,N_19656);
or U19956 (N_19956,N_19490,N_19295);
nor U19957 (N_19957,N_19398,N_19265);
or U19958 (N_19958,N_19792,N_19527);
nand U19959 (N_19959,N_19294,N_19676);
and U19960 (N_19960,N_19691,N_19775);
and U19961 (N_19961,N_19717,N_19602);
and U19962 (N_19962,N_19302,N_19314);
nor U19963 (N_19963,N_19293,N_19695);
nand U19964 (N_19964,N_19299,N_19457);
and U19965 (N_19965,N_19767,N_19220);
or U19966 (N_19966,N_19570,N_19346);
and U19967 (N_19967,N_19356,N_19219);
nor U19968 (N_19968,N_19659,N_19781);
nor U19969 (N_19969,N_19376,N_19396);
xnor U19970 (N_19970,N_19612,N_19733);
nand U19971 (N_19971,N_19523,N_19320);
or U19972 (N_19972,N_19305,N_19756);
or U19973 (N_19973,N_19237,N_19608);
xor U19974 (N_19974,N_19437,N_19344);
and U19975 (N_19975,N_19441,N_19729);
or U19976 (N_19976,N_19576,N_19794);
xor U19977 (N_19977,N_19424,N_19768);
nor U19978 (N_19978,N_19345,N_19625);
nor U19979 (N_19979,N_19361,N_19400);
and U19980 (N_19980,N_19783,N_19617);
and U19981 (N_19981,N_19531,N_19741);
or U19982 (N_19982,N_19524,N_19721);
and U19983 (N_19983,N_19275,N_19665);
nor U19984 (N_19984,N_19522,N_19313);
nand U19985 (N_19985,N_19749,N_19316);
xnor U19986 (N_19986,N_19545,N_19471);
or U19987 (N_19987,N_19510,N_19575);
or U19988 (N_19988,N_19500,N_19235);
xor U19989 (N_19989,N_19246,N_19377);
and U19990 (N_19990,N_19480,N_19497);
or U19991 (N_19991,N_19233,N_19798);
or U19992 (N_19992,N_19591,N_19653);
or U19993 (N_19993,N_19268,N_19690);
xor U19994 (N_19994,N_19300,N_19482);
xor U19995 (N_19995,N_19720,N_19208);
xor U19996 (N_19996,N_19706,N_19483);
nor U19997 (N_19997,N_19621,N_19526);
nand U19998 (N_19998,N_19669,N_19587);
nand U19999 (N_19999,N_19380,N_19605);
xor U20000 (N_20000,N_19606,N_19384);
nand U20001 (N_20001,N_19758,N_19379);
or U20002 (N_20002,N_19304,N_19388);
and U20003 (N_20003,N_19365,N_19475);
nand U20004 (N_20004,N_19742,N_19325);
or U20005 (N_20005,N_19426,N_19532);
nor U20006 (N_20006,N_19370,N_19259);
or U20007 (N_20007,N_19506,N_19589);
nor U20008 (N_20008,N_19228,N_19784);
xor U20009 (N_20009,N_19603,N_19392);
nand U20010 (N_20010,N_19574,N_19734);
and U20011 (N_20011,N_19272,N_19697);
and U20012 (N_20012,N_19338,N_19362);
or U20013 (N_20013,N_19761,N_19467);
nor U20014 (N_20014,N_19636,N_19410);
nor U20015 (N_20015,N_19411,N_19751);
xnor U20016 (N_20016,N_19679,N_19600);
and U20017 (N_20017,N_19251,N_19463);
nand U20018 (N_20018,N_19732,N_19243);
or U20019 (N_20019,N_19206,N_19507);
nor U20020 (N_20020,N_19561,N_19413);
nand U20021 (N_20021,N_19286,N_19719);
or U20022 (N_20022,N_19492,N_19607);
and U20023 (N_20023,N_19746,N_19624);
and U20024 (N_20024,N_19334,N_19773);
and U20025 (N_20025,N_19658,N_19694);
nor U20026 (N_20026,N_19498,N_19529);
and U20027 (N_20027,N_19535,N_19692);
nor U20028 (N_20028,N_19511,N_19340);
and U20029 (N_20029,N_19551,N_19301);
or U20030 (N_20030,N_19458,N_19248);
and U20031 (N_20031,N_19200,N_19533);
nand U20032 (N_20032,N_19258,N_19454);
nand U20033 (N_20033,N_19440,N_19528);
and U20034 (N_20034,N_19401,N_19757);
or U20035 (N_20035,N_19328,N_19650);
and U20036 (N_20036,N_19633,N_19641);
xor U20037 (N_20037,N_19213,N_19530);
and U20038 (N_20038,N_19447,N_19317);
xnor U20039 (N_20039,N_19487,N_19566);
xor U20040 (N_20040,N_19730,N_19724);
nor U20041 (N_20041,N_19747,N_19353);
or U20042 (N_20042,N_19297,N_19274);
nand U20043 (N_20043,N_19358,N_19354);
nand U20044 (N_20044,N_19369,N_19651);
xnor U20045 (N_20045,N_19308,N_19236);
nand U20046 (N_20046,N_19461,N_19661);
nor U20047 (N_20047,N_19666,N_19273);
xnor U20048 (N_20048,N_19212,N_19232);
xor U20049 (N_20049,N_19331,N_19478);
xnor U20050 (N_20050,N_19685,N_19240);
nand U20051 (N_20051,N_19548,N_19359);
or U20052 (N_20052,N_19514,N_19271);
or U20053 (N_20053,N_19744,N_19371);
nand U20054 (N_20054,N_19224,N_19627);
or U20055 (N_20055,N_19585,N_19479);
and U20056 (N_20056,N_19735,N_19445);
nand U20057 (N_20057,N_19611,N_19541);
and U20058 (N_20058,N_19632,N_19667);
nand U20059 (N_20059,N_19558,N_19495);
nand U20060 (N_20060,N_19202,N_19770);
and U20061 (N_20061,N_19753,N_19537);
or U20062 (N_20062,N_19254,N_19670);
nand U20063 (N_20063,N_19689,N_19484);
xnor U20064 (N_20064,N_19505,N_19432);
nand U20065 (N_20065,N_19217,N_19513);
xnor U20066 (N_20066,N_19793,N_19450);
and U20067 (N_20067,N_19315,N_19646);
xor U20068 (N_20068,N_19415,N_19774);
xor U20069 (N_20069,N_19416,N_19309);
nand U20070 (N_20070,N_19704,N_19343);
nor U20071 (N_20071,N_19759,N_19722);
and U20072 (N_20072,N_19613,N_19648);
xor U20073 (N_20073,N_19225,N_19207);
nand U20074 (N_20074,N_19244,N_19326);
and U20075 (N_20075,N_19393,N_19348);
and U20076 (N_20076,N_19686,N_19572);
nor U20077 (N_20077,N_19637,N_19339);
or U20078 (N_20078,N_19698,N_19554);
nand U20079 (N_20079,N_19681,N_19616);
nand U20080 (N_20080,N_19578,N_19352);
or U20081 (N_20081,N_19731,N_19562);
xnor U20082 (N_20082,N_19620,N_19540);
or U20083 (N_20083,N_19397,N_19662);
xnor U20084 (N_20084,N_19252,N_19615);
nand U20085 (N_20085,N_19429,N_19446);
xor U20086 (N_20086,N_19595,N_19485);
nor U20087 (N_20087,N_19553,N_19278);
nand U20088 (N_20088,N_19519,N_19223);
or U20089 (N_20089,N_19427,N_19448);
nor U20090 (N_20090,N_19350,N_19619);
or U20091 (N_20091,N_19481,N_19750);
nand U20092 (N_20092,N_19631,N_19216);
nor U20093 (N_20093,N_19368,N_19215);
xnor U20094 (N_20094,N_19312,N_19261);
nor U20095 (N_20095,N_19383,N_19329);
nor U20096 (N_20096,N_19738,N_19504);
xor U20097 (N_20097,N_19652,N_19534);
nand U20098 (N_20098,N_19203,N_19635);
nor U20099 (N_20099,N_19581,N_19647);
or U20100 (N_20100,N_19426,N_19672);
or U20101 (N_20101,N_19750,N_19249);
nand U20102 (N_20102,N_19505,N_19277);
nand U20103 (N_20103,N_19332,N_19333);
nand U20104 (N_20104,N_19585,N_19756);
nand U20105 (N_20105,N_19219,N_19689);
xor U20106 (N_20106,N_19417,N_19768);
xnor U20107 (N_20107,N_19421,N_19769);
and U20108 (N_20108,N_19724,N_19791);
or U20109 (N_20109,N_19226,N_19517);
and U20110 (N_20110,N_19721,N_19301);
nor U20111 (N_20111,N_19648,N_19686);
nand U20112 (N_20112,N_19688,N_19700);
xnor U20113 (N_20113,N_19790,N_19709);
xnor U20114 (N_20114,N_19702,N_19579);
nand U20115 (N_20115,N_19772,N_19322);
xor U20116 (N_20116,N_19569,N_19677);
or U20117 (N_20117,N_19273,N_19252);
or U20118 (N_20118,N_19420,N_19495);
nand U20119 (N_20119,N_19668,N_19722);
and U20120 (N_20120,N_19707,N_19554);
or U20121 (N_20121,N_19469,N_19466);
and U20122 (N_20122,N_19663,N_19428);
and U20123 (N_20123,N_19443,N_19247);
or U20124 (N_20124,N_19397,N_19702);
xnor U20125 (N_20125,N_19502,N_19233);
and U20126 (N_20126,N_19468,N_19507);
or U20127 (N_20127,N_19371,N_19300);
nor U20128 (N_20128,N_19786,N_19752);
or U20129 (N_20129,N_19593,N_19789);
nor U20130 (N_20130,N_19668,N_19231);
nor U20131 (N_20131,N_19207,N_19662);
and U20132 (N_20132,N_19223,N_19617);
and U20133 (N_20133,N_19437,N_19553);
nand U20134 (N_20134,N_19428,N_19246);
xnor U20135 (N_20135,N_19640,N_19477);
xor U20136 (N_20136,N_19384,N_19567);
nand U20137 (N_20137,N_19718,N_19238);
or U20138 (N_20138,N_19660,N_19401);
nor U20139 (N_20139,N_19457,N_19318);
and U20140 (N_20140,N_19686,N_19237);
or U20141 (N_20141,N_19365,N_19395);
or U20142 (N_20142,N_19293,N_19385);
nor U20143 (N_20143,N_19523,N_19785);
nand U20144 (N_20144,N_19666,N_19792);
nand U20145 (N_20145,N_19560,N_19452);
or U20146 (N_20146,N_19250,N_19754);
and U20147 (N_20147,N_19513,N_19731);
nor U20148 (N_20148,N_19251,N_19536);
xnor U20149 (N_20149,N_19361,N_19258);
xor U20150 (N_20150,N_19797,N_19476);
or U20151 (N_20151,N_19721,N_19327);
and U20152 (N_20152,N_19759,N_19251);
nand U20153 (N_20153,N_19587,N_19382);
nor U20154 (N_20154,N_19278,N_19510);
xnor U20155 (N_20155,N_19617,N_19488);
nor U20156 (N_20156,N_19623,N_19602);
nor U20157 (N_20157,N_19273,N_19570);
or U20158 (N_20158,N_19508,N_19334);
and U20159 (N_20159,N_19417,N_19215);
nor U20160 (N_20160,N_19668,N_19762);
nor U20161 (N_20161,N_19300,N_19739);
or U20162 (N_20162,N_19475,N_19538);
xnor U20163 (N_20163,N_19317,N_19500);
or U20164 (N_20164,N_19207,N_19712);
nor U20165 (N_20165,N_19766,N_19382);
nor U20166 (N_20166,N_19478,N_19519);
xor U20167 (N_20167,N_19449,N_19565);
or U20168 (N_20168,N_19791,N_19377);
and U20169 (N_20169,N_19328,N_19797);
or U20170 (N_20170,N_19312,N_19744);
nand U20171 (N_20171,N_19502,N_19384);
nor U20172 (N_20172,N_19262,N_19751);
nand U20173 (N_20173,N_19521,N_19536);
or U20174 (N_20174,N_19443,N_19753);
nor U20175 (N_20175,N_19544,N_19298);
nand U20176 (N_20176,N_19359,N_19676);
xor U20177 (N_20177,N_19514,N_19541);
xnor U20178 (N_20178,N_19618,N_19387);
nor U20179 (N_20179,N_19280,N_19559);
nor U20180 (N_20180,N_19211,N_19483);
nor U20181 (N_20181,N_19622,N_19539);
or U20182 (N_20182,N_19642,N_19587);
and U20183 (N_20183,N_19451,N_19330);
or U20184 (N_20184,N_19364,N_19617);
xor U20185 (N_20185,N_19270,N_19677);
xor U20186 (N_20186,N_19624,N_19231);
and U20187 (N_20187,N_19705,N_19742);
xnor U20188 (N_20188,N_19692,N_19371);
nor U20189 (N_20189,N_19589,N_19630);
and U20190 (N_20190,N_19321,N_19309);
nand U20191 (N_20191,N_19294,N_19240);
and U20192 (N_20192,N_19273,N_19243);
nand U20193 (N_20193,N_19644,N_19216);
xor U20194 (N_20194,N_19458,N_19609);
nor U20195 (N_20195,N_19605,N_19270);
and U20196 (N_20196,N_19555,N_19708);
nor U20197 (N_20197,N_19420,N_19709);
and U20198 (N_20198,N_19520,N_19284);
nor U20199 (N_20199,N_19467,N_19417);
and U20200 (N_20200,N_19550,N_19242);
or U20201 (N_20201,N_19225,N_19476);
nor U20202 (N_20202,N_19740,N_19604);
nand U20203 (N_20203,N_19228,N_19641);
xor U20204 (N_20204,N_19462,N_19248);
xnor U20205 (N_20205,N_19697,N_19344);
nor U20206 (N_20206,N_19287,N_19564);
xnor U20207 (N_20207,N_19371,N_19785);
or U20208 (N_20208,N_19628,N_19206);
or U20209 (N_20209,N_19272,N_19322);
xor U20210 (N_20210,N_19690,N_19759);
nand U20211 (N_20211,N_19726,N_19764);
or U20212 (N_20212,N_19251,N_19656);
or U20213 (N_20213,N_19535,N_19430);
and U20214 (N_20214,N_19260,N_19619);
or U20215 (N_20215,N_19498,N_19613);
or U20216 (N_20216,N_19692,N_19609);
xnor U20217 (N_20217,N_19640,N_19654);
nand U20218 (N_20218,N_19504,N_19326);
and U20219 (N_20219,N_19531,N_19410);
nand U20220 (N_20220,N_19519,N_19798);
or U20221 (N_20221,N_19774,N_19285);
nor U20222 (N_20222,N_19391,N_19264);
or U20223 (N_20223,N_19735,N_19301);
and U20224 (N_20224,N_19692,N_19590);
xor U20225 (N_20225,N_19471,N_19337);
nor U20226 (N_20226,N_19526,N_19306);
xor U20227 (N_20227,N_19640,N_19296);
or U20228 (N_20228,N_19444,N_19783);
nand U20229 (N_20229,N_19698,N_19293);
nand U20230 (N_20230,N_19661,N_19326);
xor U20231 (N_20231,N_19497,N_19215);
xor U20232 (N_20232,N_19235,N_19372);
and U20233 (N_20233,N_19450,N_19602);
nor U20234 (N_20234,N_19390,N_19267);
or U20235 (N_20235,N_19487,N_19207);
nor U20236 (N_20236,N_19629,N_19445);
and U20237 (N_20237,N_19353,N_19313);
and U20238 (N_20238,N_19455,N_19573);
or U20239 (N_20239,N_19308,N_19729);
and U20240 (N_20240,N_19724,N_19554);
and U20241 (N_20241,N_19560,N_19727);
xor U20242 (N_20242,N_19262,N_19527);
and U20243 (N_20243,N_19444,N_19411);
nor U20244 (N_20244,N_19570,N_19241);
xor U20245 (N_20245,N_19334,N_19323);
and U20246 (N_20246,N_19659,N_19359);
nand U20247 (N_20247,N_19328,N_19492);
and U20248 (N_20248,N_19611,N_19467);
and U20249 (N_20249,N_19713,N_19429);
or U20250 (N_20250,N_19379,N_19663);
nor U20251 (N_20251,N_19406,N_19560);
nand U20252 (N_20252,N_19537,N_19564);
nand U20253 (N_20253,N_19208,N_19713);
nand U20254 (N_20254,N_19402,N_19713);
nor U20255 (N_20255,N_19315,N_19771);
nand U20256 (N_20256,N_19670,N_19631);
nor U20257 (N_20257,N_19751,N_19332);
or U20258 (N_20258,N_19615,N_19651);
xnor U20259 (N_20259,N_19568,N_19685);
or U20260 (N_20260,N_19551,N_19206);
and U20261 (N_20261,N_19696,N_19711);
nand U20262 (N_20262,N_19465,N_19361);
or U20263 (N_20263,N_19464,N_19305);
and U20264 (N_20264,N_19484,N_19619);
nor U20265 (N_20265,N_19323,N_19399);
nand U20266 (N_20266,N_19233,N_19545);
or U20267 (N_20267,N_19331,N_19448);
and U20268 (N_20268,N_19556,N_19566);
or U20269 (N_20269,N_19590,N_19714);
nand U20270 (N_20270,N_19491,N_19732);
and U20271 (N_20271,N_19486,N_19723);
or U20272 (N_20272,N_19222,N_19552);
and U20273 (N_20273,N_19701,N_19797);
or U20274 (N_20274,N_19614,N_19785);
nor U20275 (N_20275,N_19318,N_19370);
xnor U20276 (N_20276,N_19714,N_19704);
xor U20277 (N_20277,N_19708,N_19246);
or U20278 (N_20278,N_19427,N_19777);
and U20279 (N_20279,N_19391,N_19660);
nor U20280 (N_20280,N_19451,N_19272);
nor U20281 (N_20281,N_19582,N_19298);
and U20282 (N_20282,N_19296,N_19490);
nand U20283 (N_20283,N_19698,N_19446);
or U20284 (N_20284,N_19416,N_19533);
and U20285 (N_20285,N_19746,N_19663);
nand U20286 (N_20286,N_19721,N_19470);
and U20287 (N_20287,N_19541,N_19694);
or U20288 (N_20288,N_19522,N_19576);
xnor U20289 (N_20289,N_19734,N_19730);
nor U20290 (N_20290,N_19609,N_19699);
or U20291 (N_20291,N_19262,N_19455);
and U20292 (N_20292,N_19255,N_19458);
xor U20293 (N_20293,N_19296,N_19417);
or U20294 (N_20294,N_19568,N_19657);
and U20295 (N_20295,N_19559,N_19651);
or U20296 (N_20296,N_19214,N_19533);
nand U20297 (N_20297,N_19386,N_19294);
nand U20298 (N_20298,N_19382,N_19412);
nor U20299 (N_20299,N_19501,N_19473);
and U20300 (N_20300,N_19355,N_19621);
and U20301 (N_20301,N_19497,N_19273);
nor U20302 (N_20302,N_19636,N_19530);
nor U20303 (N_20303,N_19584,N_19573);
xor U20304 (N_20304,N_19738,N_19599);
nor U20305 (N_20305,N_19391,N_19256);
or U20306 (N_20306,N_19437,N_19652);
nand U20307 (N_20307,N_19770,N_19311);
nand U20308 (N_20308,N_19516,N_19460);
nand U20309 (N_20309,N_19504,N_19312);
nor U20310 (N_20310,N_19664,N_19587);
or U20311 (N_20311,N_19642,N_19679);
and U20312 (N_20312,N_19663,N_19478);
or U20313 (N_20313,N_19251,N_19572);
and U20314 (N_20314,N_19231,N_19213);
xnor U20315 (N_20315,N_19591,N_19679);
nand U20316 (N_20316,N_19358,N_19673);
nand U20317 (N_20317,N_19399,N_19266);
xnor U20318 (N_20318,N_19293,N_19557);
nor U20319 (N_20319,N_19296,N_19779);
and U20320 (N_20320,N_19263,N_19743);
xnor U20321 (N_20321,N_19356,N_19226);
nand U20322 (N_20322,N_19711,N_19417);
xor U20323 (N_20323,N_19497,N_19749);
or U20324 (N_20324,N_19661,N_19440);
and U20325 (N_20325,N_19220,N_19504);
xnor U20326 (N_20326,N_19292,N_19388);
nand U20327 (N_20327,N_19527,N_19276);
and U20328 (N_20328,N_19453,N_19784);
nor U20329 (N_20329,N_19771,N_19685);
and U20330 (N_20330,N_19477,N_19550);
xor U20331 (N_20331,N_19497,N_19411);
or U20332 (N_20332,N_19671,N_19428);
or U20333 (N_20333,N_19666,N_19614);
nand U20334 (N_20334,N_19320,N_19475);
or U20335 (N_20335,N_19670,N_19713);
or U20336 (N_20336,N_19284,N_19665);
or U20337 (N_20337,N_19366,N_19205);
xor U20338 (N_20338,N_19647,N_19570);
or U20339 (N_20339,N_19285,N_19310);
nor U20340 (N_20340,N_19717,N_19257);
nor U20341 (N_20341,N_19621,N_19280);
xor U20342 (N_20342,N_19209,N_19710);
nor U20343 (N_20343,N_19261,N_19604);
xnor U20344 (N_20344,N_19724,N_19717);
nor U20345 (N_20345,N_19257,N_19531);
xor U20346 (N_20346,N_19734,N_19552);
nand U20347 (N_20347,N_19773,N_19411);
nor U20348 (N_20348,N_19731,N_19616);
xnor U20349 (N_20349,N_19654,N_19785);
nor U20350 (N_20350,N_19788,N_19227);
nand U20351 (N_20351,N_19650,N_19795);
nand U20352 (N_20352,N_19776,N_19230);
nand U20353 (N_20353,N_19442,N_19511);
and U20354 (N_20354,N_19539,N_19619);
and U20355 (N_20355,N_19370,N_19275);
or U20356 (N_20356,N_19383,N_19271);
nor U20357 (N_20357,N_19566,N_19752);
nand U20358 (N_20358,N_19659,N_19521);
or U20359 (N_20359,N_19521,N_19594);
nand U20360 (N_20360,N_19688,N_19333);
xnor U20361 (N_20361,N_19780,N_19217);
or U20362 (N_20362,N_19709,N_19524);
nand U20363 (N_20363,N_19407,N_19549);
and U20364 (N_20364,N_19568,N_19409);
or U20365 (N_20365,N_19463,N_19470);
and U20366 (N_20366,N_19561,N_19338);
or U20367 (N_20367,N_19533,N_19419);
nand U20368 (N_20368,N_19747,N_19787);
and U20369 (N_20369,N_19626,N_19539);
xnor U20370 (N_20370,N_19594,N_19290);
xnor U20371 (N_20371,N_19213,N_19511);
and U20372 (N_20372,N_19672,N_19336);
nand U20373 (N_20373,N_19792,N_19318);
nor U20374 (N_20374,N_19773,N_19573);
or U20375 (N_20375,N_19286,N_19480);
nor U20376 (N_20376,N_19398,N_19576);
nand U20377 (N_20377,N_19658,N_19486);
or U20378 (N_20378,N_19665,N_19516);
or U20379 (N_20379,N_19216,N_19502);
nand U20380 (N_20380,N_19547,N_19596);
or U20381 (N_20381,N_19476,N_19286);
or U20382 (N_20382,N_19756,N_19268);
or U20383 (N_20383,N_19623,N_19505);
or U20384 (N_20384,N_19342,N_19359);
nor U20385 (N_20385,N_19644,N_19488);
or U20386 (N_20386,N_19653,N_19719);
xnor U20387 (N_20387,N_19622,N_19690);
and U20388 (N_20388,N_19662,N_19499);
nor U20389 (N_20389,N_19430,N_19339);
or U20390 (N_20390,N_19422,N_19698);
xnor U20391 (N_20391,N_19435,N_19399);
nor U20392 (N_20392,N_19458,N_19624);
xor U20393 (N_20393,N_19404,N_19709);
or U20394 (N_20394,N_19687,N_19788);
nor U20395 (N_20395,N_19667,N_19767);
and U20396 (N_20396,N_19451,N_19523);
nor U20397 (N_20397,N_19481,N_19657);
and U20398 (N_20398,N_19230,N_19327);
xor U20399 (N_20399,N_19554,N_19656);
or U20400 (N_20400,N_20371,N_20189);
or U20401 (N_20401,N_20070,N_20042);
nand U20402 (N_20402,N_20011,N_20229);
nand U20403 (N_20403,N_20050,N_19878);
xnor U20404 (N_20404,N_20372,N_20194);
xnor U20405 (N_20405,N_20224,N_20043);
or U20406 (N_20406,N_20370,N_19944);
nor U20407 (N_20407,N_20089,N_20246);
nand U20408 (N_20408,N_20395,N_19937);
or U20409 (N_20409,N_19911,N_19931);
nand U20410 (N_20410,N_19820,N_20082);
nor U20411 (N_20411,N_20083,N_20167);
nor U20412 (N_20412,N_20090,N_20381);
nor U20413 (N_20413,N_19901,N_20084);
and U20414 (N_20414,N_20054,N_19929);
or U20415 (N_20415,N_20029,N_20225);
xnor U20416 (N_20416,N_19905,N_19885);
nor U20417 (N_20417,N_20285,N_20305);
and U20418 (N_20418,N_20284,N_20234);
and U20419 (N_20419,N_19818,N_20109);
nand U20420 (N_20420,N_19889,N_20261);
nand U20421 (N_20421,N_20205,N_20272);
nor U20422 (N_20422,N_19817,N_19861);
xnor U20423 (N_20423,N_20368,N_20119);
nor U20424 (N_20424,N_19830,N_19962);
xnor U20425 (N_20425,N_20377,N_20046);
nor U20426 (N_20426,N_20072,N_20062);
nand U20427 (N_20427,N_20282,N_19974);
and U20428 (N_20428,N_20164,N_20220);
and U20429 (N_20429,N_20100,N_19829);
and U20430 (N_20430,N_19886,N_20186);
nand U20431 (N_20431,N_20346,N_20379);
or U20432 (N_20432,N_19916,N_19907);
or U20433 (N_20433,N_19834,N_20324);
or U20434 (N_20434,N_19959,N_20095);
xnor U20435 (N_20435,N_20107,N_20006);
nand U20436 (N_20436,N_20059,N_20034);
or U20437 (N_20437,N_19847,N_20061);
nand U20438 (N_20438,N_20303,N_19897);
xor U20439 (N_20439,N_19917,N_20389);
nor U20440 (N_20440,N_20003,N_19971);
nor U20441 (N_20441,N_20295,N_20274);
or U20442 (N_20442,N_20240,N_20217);
nand U20443 (N_20443,N_20360,N_20275);
and U20444 (N_20444,N_19855,N_19992);
nand U20445 (N_20445,N_20338,N_20198);
or U20446 (N_20446,N_20355,N_20088);
or U20447 (N_20447,N_19835,N_20258);
xnor U20448 (N_20448,N_19895,N_20004);
and U20449 (N_20449,N_20316,N_20383);
nand U20450 (N_20450,N_19894,N_19947);
nor U20451 (N_20451,N_19921,N_20040);
nor U20452 (N_20452,N_19819,N_20369);
nand U20453 (N_20453,N_20388,N_20163);
xnor U20454 (N_20454,N_20300,N_19823);
xnor U20455 (N_20455,N_19942,N_20067);
and U20456 (N_20456,N_19859,N_20124);
and U20457 (N_20457,N_20208,N_20000);
nand U20458 (N_20458,N_20178,N_20045);
and U20459 (N_20459,N_20253,N_19953);
and U20460 (N_20460,N_20126,N_19881);
and U20461 (N_20461,N_20273,N_20117);
or U20462 (N_20462,N_20157,N_19803);
xor U20463 (N_20463,N_19925,N_19913);
nand U20464 (N_20464,N_19966,N_19806);
or U20465 (N_20465,N_19918,N_20140);
and U20466 (N_20466,N_19903,N_20196);
nand U20467 (N_20467,N_20064,N_20356);
or U20468 (N_20468,N_20147,N_19909);
and U20469 (N_20469,N_19970,N_20152);
and U20470 (N_20470,N_20214,N_20121);
and U20471 (N_20471,N_20182,N_20023);
or U20472 (N_20472,N_20375,N_20218);
and U20473 (N_20473,N_19956,N_20221);
xor U20474 (N_20474,N_20212,N_20028);
nor U20475 (N_20475,N_20291,N_20238);
or U20476 (N_20476,N_20048,N_20123);
nand U20477 (N_20477,N_20181,N_20122);
xor U20478 (N_20478,N_20174,N_20236);
xnor U20479 (N_20479,N_20330,N_20038);
or U20480 (N_20480,N_20166,N_20199);
and U20481 (N_20481,N_19828,N_19968);
and U20482 (N_20482,N_20076,N_19896);
xor U20483 (N_20483,N_20318,N_20037);
xnor U20484 (N_20484,N_20103,N_20021);
nand U20485 (N_20485,N_20333,N_20365);
nand U20486 (N_20486,N_20227,N_20080);
nor U20487 (N_20487,N_20005,N_19813);
or U20488 (N_20488,N_20130,N_19833);
nor U20489 (N_20489,N_20287,N_19914);
or U20490 (N_20490,N_20058,N_19910);
and U20491 (N_20491,N_20108,N_20328);
nand U20492 (N_20492,N_20215,N_20289);
nand U20493 (N_20493,N_20331,N_19994);
xor U20494 (N_20494,N_19809,N_20110);
or U20495 (N_20495,N_20216,N_20133);
nand U20496 (N_20496,N_20161,N_20051);
nand U20497 (N_20497,N_20184,N_20337);
and U20498 (N_20498,N_20128,N_20294);
nor U20499 (N_20499,N_20177,N_20343);
nor U20500 (N_20500,N_20116,N_20024);
or U20501 (N_20501,N_20226,N_20081);
nand U20502 (N_20502,N_19812,N_20304);
nor U20503 (N_20503,N_20271,N_19890);
xor U20504 (N_20504,N_19906,N_20131);
nor U20505 (N_20505,N_20270,N_20269);
nor U20506 (N_20506,N_20078,N_19998);
nand U20507 (N_20507,N_19802,N_20094);
or U20508 (N_20508,N_20044,N_19816);
or U20509 (N_20509,N_19986,N_20314);
nand U20510 (N_20510,N_20086,N_20142);
nand U20511 (N_20511,N_20035,N_20339);
xor U20512 (N_20512,N_20120,N_19837);
nor U20513 (N_20513,N_19843,N_20286);
and U20514 (N_20514,N_19972,N_20247);
or U20515 (N_20515,N_20266,N_20113);
nand U20516 (N_20516,N_20341,N_19934);
xor U20517 (N_20517,N_20149,N_19943);
xor U20518 (N_20518,N_20380,N_19995);
nor U20519 (N_20519,N_19892,N_20327);
nand U20520 (N_20520,N_20168,N_20374);
nor U20521 (N_20521,N_20001,N_20392);
and U20522 (N_20522,N_20399,N_20071);
or U20523 (N_20523,N_19811,N_20345);
xor U20524 (N_20524,N_19955,N_19988);
nand U20525 (N_20525,N_20326,N_19872);
xnor U20526 (N_20526,N_19854,N_20039);
and U20527 (N_20527,N_20280,N_20159);
nor U20528 (N_20528,N_20052,N_20311);
nand U20529 (N_20529,N_20230,N_20022);
and U20530 (N_20530,N_20079,N_19853);
nor U20531 (N_20531,N_20008,N_20183);
and U20532 (N_20532,N_19825,N_19891);
xnor U20533 (N_20533,N_20077,N_19844);
and U20534 (N_20534,N_20252,N_20222);
or U20535 (N_20535,N_20397,N_19923);
xor U20536 (N_20536,N_20055,N_20127);
and U20537 (N_20537,N_20138,N_20144);
xnor U20538 (N_20538,N_20170,N_20201);
or U20539 (N_20539,N_19801,N_19873);
nor U20540 (N_20540,N_19800,N_19804);
or U20541 (N_20541,N_20002,N_20366);
xnor U20542 (N_20542,N_19877,N_20364);
xnor U20543 (N_20543,N_20066,N_20193);
and U20544 (N_20544,N_19983,N_20036);
nand U20545 (N_20545,N_19805,N_19849);
and U20546 (N_20546,N_20332,N_20114);
nand U20547 (N_20547,N_20171,N_20267);
nor U20548 (N_20548,N_19946,N_20394);
or U20549 (N_20549,N_20185,N_20146);
nor U20550 (N_20550,N_19935,N_19848);
nand U20551 (N_20551,N_20243,N_19883);
nor U20552 (N_20552,N_20101,N_19884);
or U20553 (N_20553,N_20309,N_20030);
nand U20554 (N_20554,N_20298,N_20145);
or U20555 (N_20555,N_19824,N_19845);
and U20556 (N_20556,N_19990,N_20386);
nand U20557 (N_20557,N_19926,N_20192);
xnor U20558 (N_20558,N_20250,N_19887);
nor U20559 (N_20559,N_20065,N_20219);
nor U20560 (N_20560,N_19924,N_20228);
xor U20561 (N_20561,N_19950,N_20376);
xor U20562 (N_20562,N_20204,N_20092);
and U20563 (N_20563,N_20281,N_20031);
and U20564 (N_20564,N_20085,N_19997);
and U20565 (N_20565,N_19930,N_20262);
and U20566 (N_20566,N_19960,N_20319);
and U20567 (N_20567,N_20047,N_19987);
xor U20568 (N_20568,N_20249,N_19939);
and U20569 (N_20569,N_19826,N_19836);
xor U20570 (N_20570,N_20179,N_19832);
xor U20571 (N_20571,N_19871,N_19949);
nor U20572 (N_20572,N_20137,N_19821);
nand U20573 (N_20573,N_20359,N_19899);
and U20574 (N_20574,N_20393,N_20165);
or U20575 (N_20575,N_19838,N_20302);
nand U20576 (N_20576,N_20074,N_19948);
nand U20577 (N_20577,N_19951,N_20025);
and U20578 (N_20578,N_20202,N_20248);
nand U20579 (N_20579,N_20132,N_20254);
xor U20580 (N_20580,N_20136,N_20172);
nor U20581 (N_20581,N_20329,N_20239);
or U20582 (N_20582,N_20325,N_19851);
nor U20583 (N_20583,N_19973,N_20334);
or U20584 (N_20584,N_20060,N_20241);
nand U20585 (N_20585,N_20197,N_20322);
nand U20586 (N_20586,N_20056,N_20310);
nor U20587 (N_20587,N_19866,N_20347);
or U20588 (N_20588,N_20187,N_20232);
nor U20589 (N_20589,N_19940,N_20188);
nor U20590 (N_20590,N_20200,N_20158);
and U20591 (N_20591,N_20351,N_20169);
nand U20592 (N_20592,N_20278,N_20154);
and U20593 (N_20593,N_20073,N_19952);
nand U20594 (N_20594,N_20032,N_19984);
and U20595 (N_20595,N_20190,N_19868);
and U20596 (N_20596,N_19898,N_20155);
nor U20597 (N_20597,N_19870,N_20012);
nor U20598 (N_20598,N_20357,N_19864);
and U20599 (N_20599,N_20010,N_19912);
or U20600 (N_20600,N_19981,N_20026);
nor U20601 (N_20601,N_20277,N_20087);
nor U20602 (N_20602,N_20283,N_20013);
or U20603 (N_20603,N_20098,N_19865);
or U20604 (N_20604,N_20191,N_19882);
xor U20605 (N_20605,N_20244,N_19976);
and U20606 (N_20606,N_20141,N_20276);
nor U20607 (N_20607,N_20139,N_20290);
or U20608 (N_20608,N_20350,N_19858);
nor U20609 (N_20609,N_20057,N_20260);
xnor U20610 (N_20610,N_20068,N_20344);
or U20611 (N_20611,N_20148,N_19856);
or U20612 (N_20612,N_20175,N_20207);
nand U20613 (N_20613,N_19900,N_20162);
nand U20614 (N_20614,N_20323,N_20361);
xnor U20615 (N_20615,N_19827,N_19985);
xor U20616 (N_20616,N_20112,N_19941);
xnor U20617 (N_20617,N_19852,N_19999);
or U20618 (N_20618,N_19979,N_19965);
nor U20619 (N_20619,N_20069,N_20315);
nor U20620 (N_20620,N_19857,N_20237);
nor U20621 (N_20621,N_19915,N_20293);
nand U20622 (N_20622,N_19869,N_19982);
nor U20623 (N_20623,N_20210,N_20180);
and U20624 (N_20624,N_20296,N_19977);
nor U20625 (N_20625,N_20041,N_20385);
and U20626 (N_20626,N_20173,N_20213);
and U20627 (N_20627,N_19945,N_20367);
nor U20628 (N_20628,N_19815,N_19928);
nand U20629 (N_20629,N_20053,N_20349);
and U20630 (N_20630,N_20125,N_20352);
nor U20631 (N_20631,N_19860,N_19822);
xor U20632 (N_20632,N_20105,N_19936);
or U20633 (N_20633,N_20019,N_20129);
nor U20634 (N_20634,N_20396,N_20049);
nor U20635 (N_20635,N_20242,N_19902);
nand U20636 (N_20636,N_20176,N_20231);
xor U20637 (N_20637,N_19876,N_19927);
xor U20638 (N_20638,N_19933,N_20382);
nand U20639 (N_20639,N_20104,N_19922);
nor U20640 (N_20640,N_20308,N_20209);
and U20641 (N_20641,N_19879,N_20292);
xnor U20642 (N_20642,N_20143,N_19808);
and U20643 (N_20643,N_19810,N_20135);
xor U20644 (N_20644,N_19893,N_20363);
and U20645 (N_20645,N_20263,N_20235);
and U20646 (N_20646,N_20195,N_19814);
and U20647 (N_20647,N_20317,N_19888);
nand U20648 (N_20648,N_19842,N_20373);
nor U20649 (N_20649,N_20009,N_20153);
xnor U20650 (N_20650,N_19920,N_20378);
xor U20651 (N_20651,N_19996,N_20288);
nand U20652 (N_20652,N_20097,N_20340);
or U20653 (N_20653,N_19967,N_20398);
or U20654 (N_20654,N_19993,N_20279);
nor U20655 (N_20655,N_19954,N_20233);
and U20656 (N_20656,N_20075,N_20342);
or U20657 (N_20657,N_20299,N_20151);
xnor U20658 (N_20658,N_20307,N_19964);
nand U20659 (N_20659,N_20245,N_20020);
nand U20660 (N_20660,N_19919,N_20102);
xor U20661 (N_20661,N_20391,N_19980);
and U20662 (N_20662,N_20063,N_20268);
nand U20663 (N_20663,N_20321,N_20312);
or U20664 (N_20664,N_20096,N_19961);
and U20665 (N_20665,N_20256,N_20206);
and U20666 (N_20666,N_19841,N_20306);
or U20667 (N_20667,N_20093,N_20118);
or U20668 (N_20668,N_19862,N_19904);
and U20669 (N_20669,N_20016,N_19839);
and U20670 (N_20670,N_19850,N_20259);
nor U20671 (N_20671,N_20255,N_19807);
nor U20672 (N_20672,N_20160,N_19978);
nand U20673 (N_20673,N_20384,N_20027);
or U20674 (N_20674,N_20320,N_20264);
nor U20675 (N_20675,N_20211,N_19880);
nand U20676 (N_20676,N_20297,N_19957);
nor U20677 (N_20677,N_20348,N_20150);
or U20678 (N_20678,N_20203,N_20015);
xnor U20679 (N_20679,N_20223,N_19932);
nor U20680 (N_20680,N_20156,N_19867);
xnor U20681 (N_20681,N_20134,N_20106);
nand U20682 (N_20682,N_20362,N_20033);
or U20683 (N_20683,N_19969,N_20335);
and U20684 (N_20684,N_20387,N_20099);
xor U20685 (N_20685,N_19875,N_19846);
xor U20686 (N_20686,N_20301,N_19958);
nand U20687 (N_20687,N_20390,N_20313);
and U20688 (N_20688,N_19863,N_20336);
nor U20689 (N_20689,N_19908,N_19831);
xnor U20690 (N_20690,N_20014,N_19963);
or U20691 (N_20691,N_20115,N_19991);
nor U20692 (N_20692,N_20265,N_20111);
nor U20693 (N_20693,N_20251,N_20017);
and U20694 (N_20694,N_19989,N_20354);
xor U20695 (N_20695,N_20007,N_20358);
xor U20696 (N_20696,N_19975,N_20018);
or U20697 (N_20697,N_20091,N_20353);
xnor U20698 (N_20698,N_19938,N_20257);
xor U20699 (N_20699,N_19840,N_19874);
nand U20700 (N_20700,N_20224,N_19945);
and U20701 (N_20701,N_19847,N_19864);
or U20702 (N_20702,N_19837,N_20111);
and U20703 (N_20703,N_20125,N_19964);
nand U20704 (N_20704,N_20071,N_19855);
nor U20705 (N_20705,N_20325,N_19884);
xnor U20706 (N_20706,N_20299,N_19838);
nand U20707 (N_20707,N_19875,N_20399);
xor U20708 (N_20708,N_20262,N_20109);
nor U20709 (N_20709,N_19955,N_20126);
nand U20710 (N_20710,N_20101,N_19936);
or U20711 (N_20711,N_20256,N_20386);
or U20712 (N_20712,N_20273,N_20026);
xor U20713 (N_20713,N_20205,N_20298);
nor U20714 (N_20714,N_20131,N_19909);
nand U20715 (N_20715,N_20368,N_19921);
nor U20716 (N_20716,N_19903,N_20076);
nor U20717 (N_20717,N_20015,N_20098);
and U20718 (N_20718,N_20389,N_19909);
xor U20719 (N_20719,N_19925,N_19888);
nand U20720 (N_20720,N_20206,N_20042);
nand U20721 (N_20721,N_20116,N_19999);
or U20722 (N_20722,N_19955,N_19832);
and U20723 (N_20723,N_20083,N_20234);
and U20724 (N_20724,N_20384,N_20037);
xnor U20725 (N_20725,N_19854,N_20136);
and U20726 (N_20726,N_20079,N_19951);
nor U20727 (N_20727,N_19925,N_19939);
xnor U20728 (N_20728,N_20151,N_20377);
nor U20729 (N_20729,N_19832,N_19878);
and U20730 (N_20730,N_19911,N_20160);
nor U20731 (N_20731,N_19945,N_20147);
xor U20732 (N_20732,N_20123,N_20247);
and U20733 (N_20733,N_20350,N_20059);
and U20734 (N_20734,N_20149,N_20287);
or U20735 (N_20735,N_20267,N_20012);
or U20736 (N_20736,N_20289,N_19843);
and U20737 (N_20737,N_19930,N_20153);
nand U20738 (N_20738,N_20053,N_20010);
and U20739 (N_20739,N_20255,N_20133);
and U20740 (N_20740,N_20315,N_20048);
xnor U20741 (N_20741,N_20010,N_19902);
and U20742 (N_20742,N_20123,N_20069);
nor U20743 (N_20743,N_20205,N_20121);
nor U20744 (N_20744,N_20321,N_19875);
nor U20745 (N_20745,N_20053,N_20140);
xnor U20746 (N_20746,N_20036,N_20242);
and U20747 (N_20747,N_20089,N_19811);
nand U20748 (N_20748,N_20378,N_20088);
or U20749 (N_20749,N_20342,N_19850);
and U20750 (N_20750,N_20352,N_19929);
nor U20751 (N_20751,N_20340,N_20016);
or U20752 (N_20752,N_19995,N_20211);
xor U20753 (N_20753,N_19925,N_20000);
and U20754 (N_20754,N_20187,N_20047);
nor U20755 (N_20755,N_20073,N_20046);
nand U20756 (N_20756,N_20265,N_20177);
nor U20757 (N_20757,N_19862,N_19856);
or U20758 (N_20758,N_20099,N_20329);
or U20759 (N_20759,N_19801,N_19892);
xnor U20760 (N_20760,N_20293,N_20047);
nand U20761 (N_20761,N_20181,N_19821);
and U20762 (N_20762,N_19904,N_19872);
nor U20763 (N_20763,N_19906,N_19895);
nand U20764 (N_20764,N_20346,N_19960);
or U20765 (N_20765,N_19804,N_20274);
and U20766 (N_20766,N_20159,N_20142);
xnor U20767 (N_20767,N_19815,N_20376);
nand U20768 (N_20768,N_20178,N_20374);
nor U20769 (N_20769,N_20389,N_20290);
nand U20770 (N_20770,N_20340,N_19935);
nor U20771 (N_20771,N_19858,N_19945);
and U20772 (N_20772,N_20102,N_20234);
and U20773 (N_20773,N_19830,N_20313);
nor U20774 (N_20774,N_20195,N_20273);
and U20775 (N_20775,N_20141,N_20033);
xor U20776 (N_20776,N_20119,N_20009);
xnor U20777 (N_20777,N_20038,N_19809);
or U20778 (N_20778,N_20076,N_19804);
and U20779 (N_20779,N_20295,N_20230);
nand U20780 (N_20780,N_19849,N_20326);
xor U20781 (N_20781,N_20213,N_19878);
nand U20782 (N_20782,N_20026,N_19816);
xnor U20783 (N_20783,N_19869,N_20352);
and U20784 (N_20784,N_20080,N_20258);
xor U20785 (N_20785,N_20240,N_20244);
nand U20786 (N_20786,N_19957,N_20036);
and U20787 (N_20787,N_20294,N_20352);
xnor U20788 (N_20788,N_20318,N_19956);
nor U20789 (N_20789,N_20202,N_19994);
and U20790 (N_20790,N_20132,N_19909);
nor U20791 (N_20791,N_19950,N_20394);
nor U20792 (N_20792,N_20045,N_19982);
or U20793 (N_20793,N_20327,N_19893);
nor U20794 (N_20794,N_19982,N_19919);
nor U20795 (N_20795,N_20267,N_20336);
xnor U20796 (N_20796,N_20029,N_20059);
nand U20797 (N_20797,N_20237,N_20172);
and U20798 (N_20798,N_20043,N_20034);
nand U20799 (N_20799,N_20024,N_20285);
xor U20800 (N_20800,N_20016,N_20113);
nor U20801 (N_20801,N_20013,N_19946);
or U20802 (N_20802,N_20310,N_20080);
xnor U20803 (N_20803,N_20295,N_19834);
xnor U20804 (N_20804,N_19857,N_20114);
nor U20805 (N_20805,N_20237,N_20340);
and U20806 (N_20806,N_20319,N_19983);
or U20807 (N_20807,N_20391,N_20058);
nand U20808 (N_20808,N_19848,N_19914);
nor U20809 (N_20809,N_20060,N_20360);
and U20810 (N_20810,N_20273,N_20353);
nand U20811 (N_20811,N_20314,N_20158);
nand U20812 (N_20812,N_20190,N_20047);
xor U20813 (N_20813,N_20383,N_20240);
nor U20814 (N_20814,N_20396,N_20029);
and U20815 (N_20815,N_19803,N_19833);
or U20816 (N_20816,N_20093,N_19851);
nor U20817 (N_20817,N_19945,N_19919);
or U20818 (N_20818,N_20094,N_20063);
xnor U20819 (N_20819,N_20187,N_20264);
xor U20820 (N_20820,N_20330,N_20104);
or U20821 (N_20821,N_19990,N_20143);
xor U20822 (N_20822,N_19934,N_20334);
nor U20823 (N_20823,N_20115,N_19818);
nand U20824 (N_20824,N_20087,N_19987);
xnor U20825 (N_20825,N_20302,N_19966);
and U20826 (N_20826,N_19891,N_20269);
or U20827 (N_20827,N_20045,N_20084);
nand U20828 (N_20828,N_20133,N_20035);
nor U20829 (N_20829,N_20012,N_20235);
or U20830 (N_20830,N_19986,N_19868);
or U20831 (N_20831,N_20102,N_20185);
and U20832 (N_20832,N_20135,N_19906);
nor U20833 (N_20833,N_19913,N_20080);
xor U20834 (N_20834,N_20036,N_19830);
nand U20835 (N_20835,N_20029,N_19880);
and U20836 (N_20836,N_20303,N_19890);
nand U20837 (N_20837,N_20308,N_20030);
or U20838 (N_20838,N_20305,N_20367);
or U20839 (N_20839,N_20140,N_20001);
nand U20840 (N_20840,N_20314,N_19903);
and U20841 (N_20841,N_20245,N_20189);
nor U20842 (N_20842,N_20331,N_20289);
nor U20843 (N_20843,N_19841,N_19854);
nand U20844 (N_20844,N_19995,N_19951);
nand U20845 (N_20845,N_19877,N_20273);
nand U20846 (N_20846,N_20163,N_20009);
xnor U20847 (N_20847,N_19865,N_20180);
nor U20848 (N_20848,N_19868,N_20025);
xor U20849 (N_20849,N_20302,N_20393);
and U20850 (N_20850,N_19840,N_19888);
xnor U20851 (N_20851,N_20291,N_20246);
nand U20852 (N_20852,N_19941,N_20070);
xnor U20853 (N_20853,N_20126,N_20008);
xnor U20854 (N_20854,N_20052,N_20249);
or U20855 (N_20855,N_20201,N_19947);
and U20856 (N_20856,N_20140,N_19971);
and U20857 (N_20857,N_20093,N_20040);
xor U20858 (N_20858,N_20370,N_20078);
nor U20859 (N_20859,N_19890,N_19967);
nor U20860 (N_20860,N_20004,N_20009);
nand U20861 (N_20861,N_20159,N_20036);
xor U20862 (N_20862,N_20284,N_19826);
nand U20863 (N_20863,N_19945,N_19835);
nor U20864 (N_20864,N_20249,N_20384);
nand U20865 (N_20865,N_20267,N_19989);
or U20866 (N_20866,N_20089,N_19803);
nor U20867 (N_20867,N_20075,N_20244);
and U20868 (N_20868,N_20304,N_19971);
nand U20869 (N_20869,N_20149,N_20337);
and U20870 (N_20870,N_20076,N_20031);
nand U20871 (N_20871,N_19938,N_19854);
nand U20872 (N_20872,N_19930,N_20394);
nand U20873 (N_20873,N_20002,N_20065);
nor U20874 (N_20874,N_19917,N_20033);
xor U20875 (N_20875,N_20269,N_20219);
and U20876 (N_20876,N_19835,N_20304);
xor U20877 (N_20877,N_19910,N_20395);
xnor U20878 (N_20878,N_19864,N_20260);
xnor U20879 (N_20879,N_19956,N_20331);
nor U20880 (N_20880,N_19965,N_20234);
nand U20881 (N_20881,N_19874,N_19914);
nor U20882 (N_20882,N_19981,N_20257);
or U20883 (N_20883,N_20177,N_20278);
xor U20884 (N_20884,N_20177,N_19953);
nand U20885 (N_20885,N_19894,N_20239);
or U20886 (N_20886,N_20000,N_20304);
nand U20887 (N_20887,N_20390,N_20334);
and U20888 (N_20888,N_20327,N_20258);
and U20889 (N_20889,N_20085,N_20256);
or U20890 (N_20890,N_19877,N_20222);
xor U20891 (N_20891,N_20020,N_20129);
and U20892 (N_20892,N_20308,N_20304);
or U20893 (N_20893,N_19840,N_20122);
or U20894 (N_20894,N_20287,N_20061);
nand U20895 (N_20895,N_20293,N_20140);
xor U20896 (N_20896,N_19816,N_20237);
or U20897 (N_20897,N_20193,N_20079);
and U20898 (N_20898,N_20366,N_19908);
nor U20899 (N_20899,N_20214,N_20051);
or U20900 (N_20900,N_20107,N_19936);
nor U20901 (N_20901,N_20020,N_19802);
and U20902 (N_20902,N_20362,N_20245);
and U20903 (N_20903,N_20034,N_20112);
nor U20904 (N_20904,N_20069,N_19994);
and U20905 (N_20905,N_20135,N_19900);
nand U20906 (N_20906,N_19993,N_19933);
or U20907 (N_20907,N_20214,N_19822);
nor U20908 (N_20908,N_20016,N_19860);
and U20909 (N_20909,N_20174,N_20010);
or U20910 (N_20910,N_19979,N_20062);
nand U20911 (N_20911,N_20241,N_20264);
and U20912 (N_20912,N_20163,N_20186);
xnor U20913 (N_20913,N_20235,N_19933);
and U20914 (N_20914,N_20038,N_20375);
xnor U20915 (N_20915,N_19882,N_19875);
nand U20916 (N_20916,N_20218,N_19810);
nor U20917 (N_20917,N_20223,N_19950);
nor U20918 (N_20918,N_19977,N_20264);
or U20919 (N_20919,N_20168,N_20196);
nor U20920 (N_20920,N_20309,N_20362);
nand U20921 (N_20921,N_19923,N_19961);
and U20922 (N_20922,N_19928,N_20342);
nor U20923 (N_20923,N_20397,N_20162);
or U20924 (N_20924,N_19950,N_19940);
nand U20925 (N_20925,N_20279,N_19854);
or U20926 (N_20926,N_20263,N_20117);
or U20927 (N_20927,N_20306,N_20097);
or U20928 (N_20928,N_19850,N_19992);
nand U20929 (N_20929,N_19880,N_20390);
or U20930 (N_20930,N_19907,N_20012);
nor U20931 (N_20931,N_19803,N_19974);
and U20932 (N_20932,N_20372,N_20141);
or U20933 (N_20933,N_20350,N_20313);
nand U20934 (N_20934,N_20227,N_20374);
or U20935 (N_20935,N_19824,N_20180);
or U20936 (N_20936,N_20291,N_20178);
and U20937 (N_20937,N_20134,N_20207);
nor U20938 (N_20938,N_20338,N_20178);
nor U20939 (N_20939,N_20116,N_20195);
and U20940 (N_20940,N_20263,N_20349);
nor U20941 (N_20941,N_20039,N_19984);
or U20942 (N_20942,N_20085,N_20218);
or U20943 (N_20943,N_20294,N_20361);
xor U20944 (N_20944,N_19843,N_19978);
and U20945 (N_20945,N_19840,N_20216);
xor U20946 (N_20946,N_20345,N_20185);
nor U20947 (N_20947,N_20032,N_19952);
nor U20948 (N_20948,N_20200,N_20238);
and U20949 (N_20949,N_19831,N_20001);
nand U20950 (N_20950,N_20136,N_19952);
nor U20951 (N_20951,N_20177,N_20395);
or U20952 (N_20952,N_19875,N_19999);
nand U20953 (N_20953,N_20154,N_20217);
xor U20954 (N_20954,N_20116,N_20124);
or U20955 (N_20955,N_20014,N_19869);
nand U20956 (N_20956,N_19843,N_19865);
nand U20957 (N_20957,N_20211,N_20208);
nand U20958 (N_20958,N_19831,N_19964);
and U20959 (N_20959,N_20055,N_20156);
and U20960 (N_20960,N_20157,N_19984);
or U20961 (N_20961,N_20252,N_20286);
xnor U20962 (N_20962,N_19991,N_20054);
nand U20963 (N_20963,N_20274,N_20319);
nand U20964 (N_20964,N_20198,N_19939);
xor U20965 (N_20965,N_20001,N_20044);
xor U20966 (N_20966,N_19944,N_20190);
nor U20967 (N_20967,N_20124,N_20242);
or U20968 (N_20968,N_20151,N_20378);
and U20969 (N_20969,N_20155,N_20168);
or U20970 (N_20970,N_20345,N_19803);
and U20971 (N_20971,N_20364,N_20314);
nor U20972 (N_20972,N_19800,N_20383);
xnor U20973 (N_20973,N_19900,N_20103);
and U20974 (N_20974,N_20266,N_19861);
nand U20975 (N_20975,N_19800,N_19853);
and U20976 (N_20976,N_19965,N_19919);
nor U20977 (N_20977,N_20380,N_20118);
xor U20978 (N_20978,N_19838,N_20159);
nand U20979 (N_20979,N_20369,N_20015);
or U20980 (N_20980,N_20114,N_20006);
xnor U20981 (N_20981,N_19854,N_19830);
or U20982 (N_20982,N_20359,N_20397);
nand U20983 (N_20983,N_20145,N_20374);
or U20984 (N_20984,N_20084,N_20276);
xnor U20985 (N_20985,N_19969,N_20297);
and U20986 (N_20986,N_19823,N_20147);
nor U20987 (N_20987,N_20153,N_20365);
xor U20988 (N_20988,N_20018,N_19865);
or U20989 (N_20989,N_19891,N_20353);
or U20990 (N_20990,N_20081,N_20177);
or U20991 (N_20991,N_19853,N_20184);
xnor U20992 (N_20992,N_20355,N_19926);
and U20993 (N_20993,N_20343,N_19922);
nand U20994 (N_20994,N_20223,N_20169);
xor U20995 (N_20995,N_20159,N_20249);
or U20996 (N_20996,N_20266,N_19911);
and U20997 (N_20997,N_20362,N_20046);
and U20998 (N_20998,N_19913,N_20396);
nor U20999 (N_20999,N_20304,N_19958);
and U21000 (N_21000,N_20823,N_20784);
xnor U21001 (N_21001,N_20890,N_20456);
xor U21002 (N_21002,N_20941,N_20982);
or U21003 (N_21003,N_20606,N_20408);
and U21004 (N_21004,N_20762,N_20731);
nor U21005 (N_21005,N_20805,N_20786);
xnor U21006 (N_21006,N_20788,N_20780);
or U21007 (N_21007,N_20492,N_20778);
nand U21008 (N_21008,N_20645,N_20730);
or U21009 (N_21009,N_20697,N_20848);
xor U21010 (N_21010,N_20517,N_20845);
nand U21011 (N_21011,N_20956,N_20815);
xnor U21012 (N_21012,N_20767,N_20495);
xor U21013 (N_21013,N_20553,N_20842);
nand U21014 (N_21014,N_20400,N_20875);
and U21015 (N_21015,N_20558,N_20938);
nor U21016 (N_21016,N_20959,N_20807);
or U21017 (N_21017,N_20855,N_20640);
xor U21018 (N_21018,N_20797,N_20853);
or U21019 (N_21019,N_20970,N_20917);
xnor U21020 (N_21020,N_20421,N_20943);
xnor U21021 (N_21021,N_20979,N_20490);
nand U21022 (N_21022,N_20465,N_20446);
or U21023 (N_21023,N_20605,N_20967);
and U21024 (N_21024,N_20876,N_20448);
or U21025 (N_21025,N_20552,N_20531);
or U21026 (N_21026,N_20779,N_20856);
nand U21027 (N_21027,N_20945,N_20427);
nor U21028 (N_21028,N_20568,N_20739);
nand U21029 (N_21029,N_20885,N_20700);
and U21030 (N_21030,N_20732,N_20570);
nor U21031 (N_21031,N_20756,N_20992);
and U21032 (N_21032,N_20476,N_20707);
or U21033 (N_21033,N_20668,N_20954);
nand U21034 (N_21034,N_20961,N_20701);
nor U21035 (N_21035,N_20630,N_20991);
or U21036 (N_21036,N_20453,N_20463);
xor U21037 (N_21037,N_20716,N_20912);
and U21038 (N_21038,N_20884,N_20703);
nor U21039 (N_21039,N_20549,N_20627);
xor U21040 (N_21040,N_20693,N_20502);
xnor U21041 (N_21041,N_20550,N_20541);
nor U21042 (N_21042,N_20804,N_20574);
and U21043 (N_21043,N_20470,N_20987);
nor U21044 (N_21044,N_20749,N_20994);
nor U21045 (N_21045,N_20443,N_20567);
or U21046 (N_21046,N_20530,N_20711);
or U21047 (N_21047,N_20418,N_20824);
nor U21048 (N_21048,N_20903,N_20653);
or U21049 (N_21049,N_20820,N_20763);
nand U21050 (N_21050,N_20911,N_20491);
or U21051 (N_21051,N_20699,N_20962);
nor U21052 (N_21052,N_20920,N_20859);
or U21053 (N_21053,N_20978,N_20602);
nand U21054 (N_21054,N_20737,N_20613);
or U21055 (N_21055,N_20863,N_20615);
and U21056 (N_21056,N_20719,N_20721);
xnor U21057 (N_21057,N_20433,N_20772);
nor U21058 (N_21058,N_20940,N_20520);
nor U21059 (N_21059,N_20586,N_20841);
and U21060 (N_21060,N_20585,N_20907);
and U21061 (N_21061,N_20617,N_20647);
nor U21062 (N_21062,N_20838,N_20872);
or U21063 (N_21063,N_20489,N_20769);
nand U21064 (N_21064,N_20434,N_20458);
xnor U21065 (N_21065,N_20877,N_20633);
nand U21066 (N_21066,N_20901,N_20487);
and U21067 (N_21067,N_20404,N_20592);
or U21068 (N_21068,N_20768,N_20524);
or U21069 (N_21069,N_20459,N_20514);
nor U21070 (N_21070,N_20904,N_20965);
or U21071 (N_21071,N_20663,N_20950);
and U21072 (N_21072,N_20858,N_20790);
xnor U21073 (N_21073,N_20773,N_20411);
nor U21074 (N_21074,N_20847,N_20683);
nand U21075 (N_21075,N_20713,N_20942);
xor U21076 (N_21076,N_20747,N_20547);
or U21077 (N_21077,N_20641,N_20832);
and U21078 (N_21078,N_20679,N_20626);
nor U21079 (N_21079,N_20803,N_20622);
xor U21080 (N_21080,N_20422,N_20808);
xor U21081 (N_21081,N_20480,N_20720);
nor U21082 (N_21082,N_20589,N_20474);
or U21083 (N_21083,N_20637,N_20826);
nand U21084 (N_21084,N_20948,N_20793);
nor U21085 (N_21085,N_20406,N_20734);
xor U21086 (N_21086,N_20706,N_20416);
or U21087 (N_21087,N_20436,N_20523);
and U21088 (N_21088,N_20946,N_20695);
xor U21089 (N_21089,N_20728,N_20817);
nor U21090 (N_21090,N_20423,N_20795);
and U21091 (N_21091,N_20849,N_20594);
xnor U21092 (N_21092,N_20764,N_20934);
xor U21093 (N_21093,N_20914,N_20560);
nor U21094 (N_21094,N_20766,N_20441);
nor U21095 (N_21095,N_20506,N_20437);
or U21096 (N_21096,N_20902,N_20512);
and U21097 (N_21097,N_20454,N_20789);
nor U21098 (N_21098,N_20401,N_20887);
xnor U21099 (N_21099,N_20787,N_20684);
xor U21100 (N_21100,N_20481,N_20566);
and U21101 (N_21101,N_20559,N_20922);
and U21102 (N_21102,N_20968,N_20515);
or U21103 (N_21103,N_20781,N_20582);
or U21104 (N_21104,N_20714,N_20442);
and U21105 (N_21105,N_20993,N_20844);
nand U21106 (N_21106,N_20745,N_20634);
nor U21107 (N_21107,N_20818,N_20879);
nor U21108 (N_21108,N_20727,N_20537);
and U21109 (N_21109,N_20871,N_20625);
nand U21110 (N_21110,N_20715,N_20510);
or U21111 (N_21111,N_20462,N_20403);
xor U21112 (N_21112,N_20452,N_20986);
nand U21113 (N_21113,N_20483,N_20659);
nor U21114 (N_21114,N_20665,N_20616);
and U21115 (N_21115,N_20735,N_20931);
nand U21116 (N_21116,N_20681,N_20581);
xor U21117 (N_21117,N_20464,N_20973);
nor U21118 (N_21118,N_20981,N_20729);
and U21119 (N_21119,N_20833,N_20525);
nand U21120 (N_21120,N_20930,N_20866);
xnor U21121 (N_21121,N_20542,N_20526);
xor U21122 (N_21122,N_20504,N_20688);
nand U21123 (N_21123,N_20676,N_20445);
or U21124 (N_21124,N_20989,N_20527);
nor U21125 (N_21125,N_20825,N_20646);
and U21126 (N_21126,N_20494,N_20674);
nor U21127 (N_21127,N_20428,N_20460);
nand U21128 (N_21128,N_20748,N_20852);
and U21129 (N_21129,N_20759,N_20596);
or U21130 (N_21130,N_20750,N_20412);
nor U21131 (N_21131,N_20984,N_20758);
or U21132 (N_21132,N_20738,N_20600);
xnor U21133 (N_21133,N_20425,N_20998);
xor U21134 (N_21134,N_20892,N_20806);
nand U21135 (N_21135,N_20794,N_20846);
or U21136 (N_21136,N_20587,N_20621);
xor U21137 (N_21137,N_20839,N_20821);
nor U21138 (N_21138,N_20644,N_20840);
nor U21139 (N_21139,N_20649,N_20429);
and U21140 (N_21140,N_20664,N_20573);
xnor U21141 (N_21141,N_20761,N_20609);
xnor U21142 (N_21142,N_20447,N_20635);
nor U21143 (N_21143,N_20535,N_20862);
and U21144 (N_21144,N_20742,N_20673);
xnor U21145 (N_21145,N_20897,N_20886);
xnor U21146 (N_21146,N_20643,N_20963);
or U21147 (N_21147,N_20791,N_20977);
nor U21148 (N_21148,N_20623,N_20424);
nand U21149 (N_21149,N_20869,N_20819);
nor U21150 (N_21150,N_20562,N_20975);
nor U21151 (N_21151,N_20451,N_20677);
nand U21152 (N_21152,N_20572,N_20528);
or U21153 (N_21153,N_20686,N_20509);
nand U21154 (N_21154,N_20996,N_20583);
and U21155 (N_21155,N_20976,N_20657);
xor U21156 (N_21156,N_20532,N_20880);
xnor U21157 (N_21157,N_20420,N_20933);
nand U21158 (N_21158,N_20417,N_20923);
nand U21159 (N_21159,N_20682,N_20540);
xnor U21160 (N_21160,N_20698,N_20811);
or U21161 (N_21161,N_20926,N_20444);
and U21162 (N_21162,N_20680,N_20958);
and U21163 (N_21163,N_20857,N_20607);
or U21164 (N_21164,N_20836,N_20571);
nand U21165 (N_21165,N_20783,N_20801);
xor U21166 (N_21166,N_20538,N_20947);
nand U21167 (N_21167,N_20472,N_20776);
and U21168 (N_21168,N_20752,N_20936);
or U21169 (N_21169,N_20753,N_20988);
xor U21170 (N_21170,N_20900,N_20899);
nand U21171 (N_21171,N_20705,N_20757);
and U21172 (N_21172,N_20662,N_20685);
and U21173 (N_21173,N_20642,N_20419);
nand U21174 (N_21174,N_20765,N_20499);
nand U21175 (N_21175,N_20407,N_20928);
xor U21176 (N_21176,N_20505,N_20544);
nor U21177 (N_21177,N_20500,N_20733);
xor U21178 (N_21178,N_20726,N_20496);
nor U21179 (N_21179,N_20850,N_20593);
nand U21180 (N_21180,N_20628,N_20614);
xor U21181 (N_21181,N_20955,N_20966);
and U21182 (N_21182,N_20438,N_20932);
or U21183 (N_21183,N_20529,N_20744);
nand U21184 (N_21184,N_20835,N_20409);
nor U21185 (N_21185,N_20898,N_20830);
or U21186 (N_21186,N_20503,N_20608);
xor U21187 (N_21187,N_20953,N_20485);
or U21188 (N_21188,N_20770,N_20837);
nand U21189 (N_21189,N_20557,N_20771);
nand U21190 (N_21190,N_20522,N_20618);
nor U21191 (N_21191,N_20812,N_20478);
or U21192 (N_21192,N_20908,N_20473);
xor U21193 (N_21193,N_20661,N_20980);
nor U21194 (N_21194,N_20648,N_20997);
nor U21195 (N_21195,N_20906,N_20450);
xnor U21196 (N_21196,N_20736,N_20760);
nor U21197 (N_21197,N_20482,N_20577);
nor U21198 (N_21198,N_20533,N_20691);
nor U21199 (N_21199,N_20655,N_20591);
nor U21200 (N_21200,N_20689,N_20569);
and U21201 (N_21201,N_20939,N_20822);
xor U21202 (N_21202,N_20548,N_20414);
xor U21203 (N_21203,N_20894,N_20410);
or U21204 (N_21204,N_20670,N_20755);
and U21205 (N_21205,N_20814,N_20435);
and U21206 (N_21206,N_20519,N_20488);
nand U21207 (N_21207,N_20666,N_20829);
or U21208 (N_21208,N_20584,N_20580);
and U21209 (N_21209,N_20590,N_20893);
nor U21210 (N_21210,N_20651,N_20467);
and U21211 (N_21211,N_20466,N_20426);
xnor U21212 (N_21212,N_20831,N_20656);
or U21213 (N_21213,N_20694,N_20619);
and U21214 (N_21214,N_20985,N_20971);
nor U21215 (N_21215,N_20710,N_20889);
and U21216 (N_21216,N_20951,N_20579);
xnor U21217 (N_21217,N_20484,N_20798);
or U21218 (N_21218,N_20565,N_20782);
xor U21219 (N_21219,N_20743,N_20775);
or U21220 (N_21220,N_20690,N_20927);
nand U21221 (N_21221,N_20874,N_20652);
nor U21222 (N_21222,N_20539,N_20905);
xnor U21223 (N_21223,N_20999,N_20702);
and U21224 (N_21224,N_20654,N_20888);
nor U21225 (N_21225,N_20861,N_20974);
and U21226 (N_21226,N_20471,N_20631);
nor U21227 (N_21227,N_20810,N_20561);
or U21228 (N_21228,N_20599,N_20595);
nand U21229 (N_21229,N_20816,N_20669);
nand U21230 (N_21230,N_20671,N_20722);
or U21231 (N_21231,N_20604,N_20545);
nor U21232 (N_21232,N_20878,N_20827);
xor U21233 (N_21233,N_20612,N_20774);
or U21234 (N_21234,N_20475,N_20461);
nor U21235 (N_21235,N_20834,N_20439);
or U21236 (N_21236,N_20915,N_20629);
xor U21237 (N_21237,N_20972,N_20498);
nand U21238 (N_21238,N_20588,N_20518);
nand U21239 (N_21239,N_20477,N_20723);
nor U21240 (N_21240,N_20546,N_20575);
nor U21241 (N_21241,N_20620,N_20983);
xor U21242 (N_21242,N_20611,N_20860);
nand U21243 (N_21243,N_20740,N_20431);
or U21244 (N_21244,N_20990,N_20724);
or U21245 (N_21245,N_20712,N_20828);
nand U21246 (N_21246,N_20457,N_20658);
and U21247 (N_21247,N_20455,N_20678);
nor U21248 (N_21248,N_20598,N_20718);
nand U21249 (N_21249,N_20469,N_20868);
or U21250 (N_21250,N_20513,N_20957);
and U21251 (N_21251,N_20796,N_20430);
xor U21252 (N_21252,N_20964,N_20809);
nand U21253 (N_21253,N_20751,N_20925);
xnor U21254 (N_21254,N_20479,N_20675);
xnor U21255 (N_21255,N_20864,N_20854);
and U21256 (N_21256,N_20660,N_20883);
nor U21257 (N_21257,N_20534,N_20777);
nand U21258 (N_21258,N_20725,N_20536);
and U21259 (N_21259,N_20937,N_20687);
or U21260 (N_21260,N_20468,N_20555);
or U21261 (N_21261,N_20597,N_20891);
xnor U21262 (N_21262,N_20717,N_20402);
nor U21263 (N_21263,N_20919,N_20944);
or U21264 (N_21264,N_20449,N_20501);
nand U21265 (N_21265,N_20610,N_20754);
or U21266 (N_21266,N_20521,N_20516);
or U21267 (N_21267,N_20918,N_20667);
or U21268 (N_21268,N_20709,N_20865);
nor U21269 (N_21269,N_20867,N_20881);
xnor U21270 (N_21270,N_20909,N_20799);
or U21271 (N_21271,N_20916,N_20636);
or U21272 (N_21272,N_20802,N_20440);
nor U21273 (N_21273,N_20493,N_20708);
nand U21274 (N_21274,N_20813,N_20639);
and U21275 (N_21275,N_20935,N_20969);
nor U21276 (N_21276,N_20696,N_20895);
nor U21277 (N_21277,N_20432,N_20870);
nor U21278 (N_21278,N_20910,N_20413);
and U21279 (N_21279,N_20929,N_20624);
and U21280 (N_21280,N_20896,N_20672);
and U21281 (N_21281,N_20960,N_20564);
or U21282 (N_21282,N_20603,N_20704);
and U21283 (N_21283,N_20785,N_20995);
nor U21284 (N_21284,N_20952,N_20873);
or U21285 (N_21285,N_20405,N_20792);
nand U21286 (N_21286,N_20508,N_20576);
nand U21287 (N_21287,N_20563,N_20551);
nor U21288 (N_21288,N_20924,N_20415);
and U21289 (N_21289,N_20632,N_20556);
nand U21290 (N_21290,N_20843,N_20851);
and U21291 (N_21291,N_20741,N_20746);
xor U21292 (N_21292,N_20650,N_20882);
nand U21293 (N_21293,N_20601,N_20543);
nor U21294 (N_21294,N_20507,N_20921);
and U21295 (N_21295,N_20800,N_20486);
xor U21296 (N_21296,N_20511,N_20554);
nor U21297 (N_21297,N_20913,N_20578);
nand U21298 (N_21298,N_20497,N_20638);
and U21299 (N_21299,N_20949,N_20692);
nand U21300 (N_21300,N_20536,N_20991);
nand U21301 (N_21301,N_20986,N_20727);
nor U21302 (N_21302,N_20444,N_20578);
nor U21303 (N_21303,N_20683,N_20436);
nand U21304 (N_21304,N_20499,N_20813);
and U21305 (N_21305,N_20922,N_20990);
nor U21306 (N_21306,N_20546,N_20852);
nor U21307 (N_21307,N_20881,N_20704);
xnor U21308 (N_21308,N_20760,N_20752);
nand U21309 (N_21309,N_20738,N_20401);
and U21310 (N_21310,N_20846,N_20875);
xor U21311 (N_21311,N_20739,N_20907);
nand U21312 (N_21312,N_20588,N_20932);
nand U21313 (N_21313,N_20495,N_20521);
nor U21314 (N_21314,N_20869,N_20921);
or U21315 (N_21315,N_20964,N_20607);
nor U21316 (N_21316,N_20914,N_20869);
and U21317 (N_21317,N_20748,N_20724);
or U21318 (N_21318,N_20866,N_20758);
and U21319 (N_21319,N_20839,N_20877);
nor U21320 (N_21320,N_20669,N_20735);
nor U21321 (N_21321,N_20756,N_20786);
nand U21322 (N_21322,N_20620,N_20907);
nand U21323 (N_21323,N_20553,N_20869);
nand U21324 (N_21324,N_20664,N_20725);
nand U21325 (N_21325,N_20469,N_20979);
or U21326 (N_21326,N_20821,N_20408);
xor U21327 (N_21327,N_20570,N_20995);
or U21328 (N_21328,N_20629,N_20982);
nand U21329 (N_21329,N_20985,N_20572);
and U21330 (N_21330,N_20640,N_20616);
xnor U21331 (N_21331,N_20771,N_20474);
or U21332 (N_21332,N_20728,N_20476);
nor U21333 (N_21333,N_20499,N_20418);
xnor U21334 (N_21334,N_20850,N_20685);
and U21335 (N_21335,N_20794,N_20442);
or U21336 (N_21336,N_20987,N_20754);
or U21337 (N_21337,N_20670,N_20489);
or U21338 (N_21338,N_20450,N_20742);
xor U21339 (N_21339,N_20995,N_20588);
or U21340 (N_21340,N_20906,N_20444);
xor U21341 (N_21341,N_20928,N_20587);
or U21342 (N_21342,N_20419,N_20576);
or U21343 (N_21343,N_20700,N_20866);
xor U21344 (N_21344,N_20472,N_20415);
and U21345 (N_21345,N_20897,N_20651);
nand U21346 (N_21346,N_20850,N_20616);
nor U21347 (N_21347,N_20507,N_20660);
nand U21348 (N_21348,N_20993,N_20765);
xnor U21349 (N_21349,N_20911,N_20853);
nand U21350 (N_21350,N_20469,N_20583);
nor U21351 (N_21351,N_20549,N_20755);
or U21352 (N_21352,N_20667,N_20441);
nand U21353 (N_21353,N_20726,N_20930);
nand U21354 (N_21354,N_20545,N_20898);
nand U21355 (N_21355,N_20875,N_20799);
xor U21356 (N_21356,N_20524,N_20913);
or U21357 (N_21357,N_20579,N_20949);
xor U21358 (N_21358,N_20655,N_20978);
xnor U21359 (N_21359,N_20950,N_20486);
nor U21360 (N_21360,N_20759,N_20882);
nor U21361 (N_21361,N_20426,N_20520);
or U21362 (N_21362,N_20943,N_20770);
or U21363 (N_21363,N_20963,N_20618);
and U21364 (N_21364,N_20635,N_20541);
or U21365 (N_21365,N_20656,N_20768);
or U21366 (N_21366,N_20485,N_20408);
nand U21367 (N_21367,N_20430,N_20637);
xor U21368 (N_21368,N_20451,N_20968);
and U21369 (N_21369,N_20470,N_20575);
and U21370 (N_21370,N_20407,N_20708);
or U21371 (N_21371,N_20406,N_20900);
xnor U21372 (N_21372,N_20865,N_20544);
nand U21373 (N_21373,N_20896,N_20789);
nor U21374 (N_21374,N_20560,N_20452);
nand U21375 (N_21375,N_20458,N_20681);
nand U21376 (N_21376,N_20999,N_20825);
and U21377 (N_21377,N_20932,N_20765);
and U21378 (N_21378,N_20759,N_20838);
and U21379 (N_21379,N_20540,N_20908);
nor U21380 (N_21380,N_20969,N_20581);
or U21381 (N_21381,N_20882,N_20981);
nor U21382 (N_21382,N_20832,N_20820);
or U21383 (N_21383,N_20533,N_20526);
nor U21384 (N_21384,N_20934,N_20869);
or U21385 (N_21385,N_20431,N_20547);
xor U21386 (N_21386,N_20625,N_20763);
xnor U21387 (N_21387,N_20744,N_20667);
xnor U21388 (N_21388,N_20886,N_20772);
xor U21389 (N_21389,N_20794,N_20515);
and U21390 (N_21390,N_20763,N_20771);
nand U21391 (N_21391,N_20511,N_20876);
nor U21392 (N_21392,N_20678,N_20900);
nand U21393 (N_21393,N_20498,N_20820);
or U21394 (N_21394,N_20896,N_20507);
xnor U21395 (N_21395,N_20974,N_20789);
nor U21396 (N_21396,N_20612,N_20469);
xor U21397 (N_21397,N_20585,N_20435);
nand U21398 (N_21398,N_20444,N_20952);
and U21399 (N_21399,N_20902,N_20730);
nor U21400 (N_21400,N_20603,N_20497);
and U21401 (N_21401,N_20817,N_20612);
nand U21402 (N_21402,N_20924,N_20897);
nand U21403 (N_21403,N_20852,N_20948);
nand U21404 (N_21404,N_20732,N_20659);
and U21405 (N_21405,N_20428,N_20553);
or U21406 (N_21406,N_20947,N_20882);
nor U21407 (N_21407,N_20920,N_20849);
xor U21408 (N_21408,N_20811,N_20683);
xor U21409 (N_21409,N_20973,N_20663);
nor U21410 (N_21410,N_20651,N_20682);
nand U21411 (N_21411,N_20925,N_20710);
or U21412 (N_21412,N_20791,N_20792);
xnor U21413 (N_21413,N_20993,N_20430);
or U21414 (N_21414,N_20568,N_20430);
xor U21415 (N_21415,N_20756,N_20508);
xnor U21416 (N_21416,N_20421,N_20467);
nand U21417 (N_21417,N_20634,N_20717);
nor U21418 (N_21418,N_20980,N_20625);
and U21419 (N_21419,N_20474,N_20927);
and U21420 (N_21420,N_20633,N_20834);
nor U21421 (N_21421,N_20412,N_20589);
nor U21422 (N_21422,N_20658,N_20943);
nand U21423 (N_21423,N_20873,N_20499);
xnor U21424 (N_21424,N_20513,N_20583);
and U21425 (N_21425,N_20874,N_20905);
xnor U21426 (N_21426,N_20913,N_20671);
or U21427 (N_21427,N_20898,N_20578);
xor U21428 (N_21428,N_20582,N_20602);
nand U21429 (N_21429,N_20949,N_20403);
xnor U21430 (N_21430,N_20630,N_20497);
nor U21431 (N_21431,N_20737,N_20412);
nand U21432 (N_21432,N_20547,N_20963);
xor U21433 (N_21433,N_20869,N_20707);
nor U21434 (N_21434,N_20402,N_20417);
xnor U21435 (N_21435,N_20926,N_20910);
nand U21436 (N_21436,N_20674,N_20565);
and U21437 (N_21437,N_20666,N_20632);
and U21438 (N_21438,N_20592,N_20573);
nand U21439 (N_21439,N_20580,N_20779);
xor U21440 (N_21440,N_20703,N_20697);
or U21441 (N_21441,N_20459,N_20903);
nand U21442 (N_21442,N_20565,N_20473);
nor U21443 (N_21443,N_20995,N_20625);
xnor U21444 (N_21444,N_20996,N_20531);
nor U21445 (N_21445,N_20426,N_20623);
and U21446 (N_21446,N_20634,N_20789);
or U21447 (N_21447,N_20979,N_20887);
nand U21448 (N_21448,N_20592,N_20752);
and U21449 (N_21449,N_20524,N_20823);
or U21450 (N_21450,N_20649,N_20761);
or U21451 (N_21451,N_20421,N_20744);
and U21452 (N_21452,N_20431,N_20942);
or U21453 (N_21453,N_20648,N_20743);
nand U21454 (N_21454,N_20867,N_20857);
xor U21455 (N_21455,N_20425,N_20571);
nand U21456 (N_21456,N_20982,N_20661);
or U21457 (N_21457,N_20456,N_20554);
nand U21458 (N_21458,N_20471,N_20585);
nand U21459 (N_21459,N_20774,N_20849);
nor U21460 (N_21460,N_20470,N_20431);
nor U21461 (N_21461,N_20588,N_20658);
nor U21462 (N_21462,N_20638,N_20514);
or U21463 (N_21463,N_20661,N_20669);
nor U21464 (N_21464,N_20722,N_20988);
or U21465 (N_21465,N_20544,N_20901);
nor U21466 (N_21466,N_20705,N_20746);
and U21467 (N_21467,N_20813,N_20657);
xor U21468 (N_21468,N_20610,N_20681);
nand U21469 (N_21469,N_20853,N_20903);
nor U21470 (N_21470,N_20588,N_20645);
nand U21471 (N_21471,N_20690,N_20704);
nor U21472 (N_21472,N_20774,N_20567);
nor U21473 (N_21473,N_20968,N_20853);
xnor U21474 (N_21474,N_20629,N_20810);
nor U21475 (N_21475,N_20816,N_20780);
nor U21476 (N_21476,N_20755,N_20690);
or U21477 (N_21477,N_20511,N_20947);
or U21478 (N_21478,N_20866,N_20515);
and U21479 (N_21479,N_20790,N_20730);
nor U21480 (N_21480,N_20581,N_20724);
or U21481 (N_21481,N_20526,N_20771);
nand U21482 (N_21482,N_20794,N_20718);
or U21483 (N_21483,N_20922,N_20944);
xnor U21484 (N_21484,N_20535,N_20409);
nor U21485 (N_21485,N_20775,N_20946);
xor U21486 (N_21486,N_20832,N_20478);
and U21487 (N_21487,N_20790,N_20664);
xor U21488 (N_21488,N_20435,N_20721);
nand U21489 (N_21489,N_20552,N_20666);
xor U21490 (N_21490,N_20818,N_20820);
nor U21491 (N_21491,N_20431,N_20419);
nor U21492 (N_21492,N_20431,N_20465);
nand U21493 (N_21493,N_20718,N_20553);
or U21494 (N_21494,N_20793,N_20769);
xor U21495 (N_21495,N_20689,N_20755);
nand U21496 (N_21496,N_20580,N_20924);
and U21497 (N_21497,N_20983,N_20473);
nand U21498 (N_21498,N_20551,N_20935);
nand U21499 (N_21499,N_20536,N_20949);
xnor U21500 (N_21500,N_20684,N_20694);
xor U21501 (N_21501,N_20599,N_20822);
nand U21502 (N_21502,N_20407,N_20427);
or U21503 (N_21503,N_20996,N_20645);
nand U21504 (N_21504,N_20664,N_20749);
xor U21505 (N_21505,N_20485,N_20990);
nor U21506 (N_21506,N_20679,N_20771);
nand U21507 (N_21507,N_20764,N_20562);
or U21508 (N_21508,N_20902,N_20992);
nand U21509 (N_21509,N_20426,N_20787);
nor U21510 (N_21510,N_20432,N_20645);
nor U21511 (N_21511,N_20719,N_20838);
or U21512 (N_21512,N_20929,N_20599);
nor U21513 (N_21513,N_20653,N_20998);
xnor U21514 (N_21514,N_20630,N_20978);
or U21515 (N_21515,N_20704,N_20662);
nor U21516 (N_21516,N_20984,N_20833);
xor U21517 (N_21517,N_20733,N_20860);
or U21518 (N_21518,N_20616,N_20976);
xor U21519 (N_21519,N_20965,N_20542);
nand U21520 (N_21520,N_20449,N_20627);
or U21521 (N_21521,N_20835,N_20401);
or U21522 (N_21522,N_20866,N_20864);
nor U21523 (N_21523,N_20578,N_20738);
or U21524 (N_21524,N_20961,N_20521);
and U21525 (N_21525,N_20732,N_20683);
nor U21526 (N_21526,N_20449,N_20417);
nor U21527 (N_21527,N_20797,N_20870);
nand U21528 (N_21528,N_20977,N_20897);
nand U21529 (N_21529,N_20826,N_20747);
xor U21530 (N_21530,N_20756,N_20472);
or U21531 (N_21531,N_20403,N_20474);
or U21532 (N_21532,N_20436,N_20655);
xnor U21533 (N_21533,N_20644,N_20509);
or U21534 (N_21534,N_20640,N_20530);
xnor U21535 (N_21535,N_20436,N_20819);
nor U21536 (N_21536,N_20642,N_20579);
nand U21537 (N_21537,N_20851,N_20653);
xor U21538 (N_21538,N_20449,N_20569);
nand U21539 (N_21539,N_20814,N_20481);
nor U21540 (N_21540,N_20699,N_20909);
nand U21541 (N_21541,N_20950,N_20588);
xor U21542 (N_21542,N_20653,N_20787);
xnor U21543 (N_21543,N_20990,N_20596);
nand U21544 (N_21544,N_20844,N_20821);
nand U21545 (N_21545,N_20782,N_20898);
nand U21546 (N_21546,N_20506,N_20945);
or U21547 (N_21547,N_20776,N_20970);
nand U21548 (N_21548,N_20785,N_20840);
nor U21549 (N_21549,N_20621,N_20862);
nor U21550 (N_21550,N_20863,N_20881);
or U21551 (N_21551,N_20829,N_20816);
and U21552 (N_21552,N_20939,N_20482);
nand U21553 (N_21553,N_20806,N_20414);
nor U21554 (N_21554,N_20711,N_20583);
xnor U21555 (N_21555,N_20841,N_20964);
and U21556 (N_21556,N_20911,N_20607);
nor U21557 (N_21557,N_20799,N_20920);
nor U21558 (N_21558,N_20621,N_20994);
nor U21559 (N_21559,N_20898,N_20918);
nand U21560 (N_21560,N_20841,N_20761);
nor U21561 (N_21561,N_20522,N_20951);
nand U21562 (N_21562,N_20576,N_20561);
nand U21563 (N_21563,N_20702,N_20807);
and U21564 (N_21564,N_20769,N_20986);
nor U21565 (N_21565,N_20683,N_20669);
nor U21566 (N_21566,N_20597,N_20835);
nand U21567 (N_21567,N_20463,N_20930);
or U21568 (N_21568,N_20452,N_20421);
xnor U21569 (N_21569,N_20858,N_20625);
and U21570 (N_21570,N_20625,N_20760);
and U21571 (N_21571,N_20447,N_20665);
and U21572 (N_21572,N_20880,N_20757);
nor U21573 (N_21573,N_20911,N_20650);
and U21574 (N_21574,N_20921,N_20772);
nand U21575 (N_21575,N_20997,N_20728);
xor U21576 (N_21576,N_20707,N_20848);
nor U21577 (N_21577,N_20625,N_20682);
and U21578 (N_21578,N_20824,N_20950);
xor U21579 (N_21579,N_20778,N_20819);
and U21580 (N_21580,N_20899,N_20961);
or U21581 (N_21581,N_20425,N_20583);
nor U21582 (N_21582,N_20723,N_20559);
nand U21583 (N_21583,N_20941,N_20551);
and U21584 (N_21584,N_20666,N_20826);
nand U21585 (N_21585,N_20654,N_20515);
nand U21586 (N_21586,N_20850,N_20949);
and U21587 (N_21587,N_20976,N_20556);
nand U21588 (N_21588,N_20870,N_20590);
and U21589 (N_21589,N_20646,N_20851);
nor U21590 (N_21590,N_20673,N_20986);
and U21591 (N_21591,N_20622,N_20832);
and U21592 (N_21592,N_20672,N_20527);
nand U21593 (N_21593,N_20443,N_20956);
nor U21594 (N_21594,N_20977,N_20532);
or U21595 (N_21595,N_20429,N_20749);
nand U21596 (N_21596,N_20711,N_20400);
or U21597 (N_21597,N_20470,N_20631);
nand U21598 (N_21598,N_20698,N_20910);
nor U21599 (N_21599,N_20910,N_20909);
xor U21600 (N_21600,N_21466,N_21400);
or U21601 (N_21601,N_21195,N_21096);
xnor U21602 (N_21602,N_21463,N_21072);
or U21603 (N_21603,N_21217,N_21546);
and U21604 (N_21604,N_21022,N_21432);
nor U21605 (N_21605,N_21447,N_21272);
nand U21606 (N_21606,N_21364,N_21251);
xor U21607 (N_21607,N_21495,N_21549);
or U21608 (N_21608,N_21352,N_21468);
or U21609 (N_21609,N_21535,N_21425);
or U21610 (N_21610,N_21524,N_21006);
nor U21611 (N_21611,N_21194,N_21223);
xor U21612 (N_21612,N_21051,N_21299);
xnor U21613 (N_21613,N_21274,N_21211);
xnor U21614 (N_21614,N_21530,N_21550);
and U21615 (N_21615,N_21474,N_21513);
and U21616 (N_21616,N_21316,N_21357);
or U21617 (N_21617,N_21556,N_21236);
or U21618 (N_21618,N_21449,N_21067);
or U21619 (N_21619,N_21553,N_21087);
nand U21620 (N_21620,N_21141,N_21255);
nor U21621 (N_21621,N_21328,N_21406);
or U21622 (N_21622,N_21142,N_21075);
xor U21623 (N_21623,N_21534,N_21107);
and U21624 (N_21624,N_21089,N_21128);
nand U21625 (N_21625,N_21370,N_21247);
xor U21626 (N_21626,N_21060,N_21069);
or U21627 (N_21627,N_21053,N_21371);
xor U21628 (N_21628,N_21309,N_21202);
and U21629 (N_21629,N_21266,N_21313);
and U21630 (N_21630,N_21506,N_21099);
nand U21631 (N_21631,N_21333,N_21153);
nor U21632 (N_21632,N_21215,N_21189);
or U21633 (N_21633,N_21441,N_21058);
xor U21634 (N_21634,N_21159,N_21030);
and U21635 (N_21635,N_21175,N_21212);
nand U21636 (N_21636,N_21348,N_21482);
or U21637 (N_21637,N_21599,N_21054);
or U21638 (N_21638,N_21293,N_21584);
nand U21639 (N_21639,N_21042,N_21041);
xor U21640 (N_21640,N_21507,N_21283);
xor U21641 (N_21641,N_21487,N_21170);
and U21642 (N_21642,N_21484,N_21164);
or U21643 (N_21643,N_21095,N_21509);
nand U21644 (N_21644,N_21214,N_21291);
nand U21645 (N_21645,N_21252,N_21290);
xnor U21646 (N_21646,N_21376,N_21210);
xor U21647 (N_21647,N_21322,N_21169);
nor U21648 (N_21648,N_21512,N_21500);
or U21649 (N_21649,N_21080,N_21472);
or U21650 (N_21650,N_21485,N_21174);
and U21651 (N_21651,N_21342,N_21124);
or U21652 (N_21652,N_21511,N_21008);
nand U21653 (N_21653,N_21039,N_21454);
nor U21654 (N_21654,N_21043,N_21200);
xnor U21655 (N_21655,N_21122,N_21372);
nand U21656 (N_21656,N_21577,N_21455);
and U21657 (N_21657,N_21418,N_21315);
and U21658 (N_21658,N_21413,N_21559);
nor U21659 (N_21659,N_21350,N_21477);
nand U21660 (N_21660,N_21542,N_21243);
and U21661 (N_21661,N_21388,N_21088);
xnor U21662 (N_21662,N_21526,N_21579);
nor U21663 (N_21663,N_21057,N_21445);
or U21664 (N_21664,N_21369,N_21392);
xor U21665 (N_21665,N_21156,N_21135);
nand U21666 (N_21666,N_21544,N_21408);
nand U21667 (N_21667,N_21181,N_21327);
xor U21668 (N_21668,N_21358,N_21363);
nor U21669 (N_21669,N_21049,N_21384);
or U21670 (N_21670,N_21160,N_21325);
or U21671 (N_21671,N_21578,N_21233);
xor U21672 (N_21672,N_21422,N_21476);
or U21673 (N_21673,N_21587,N_21027);
nand U21674 (N_21674,N_21197,N_21586);
xnor U21675 (N_21675,N_21411,N_21521);
nand U21676 (N_21676,N_21321,N_21176);
and U21677 (N_21677,N_21032,N_21136);
nand U21678 (N_21678,N_21115,N_21345);
or U21679 (N_21679,N_21204,N_21470);
and U21680 (N_21680,N_21209,N_21462);
nand U21681 (N_21681,N_21101,N_21368);
nor U21682 (N_21682,N_21227,N_21131);
or U21683 (N_21683,N_21488,N_21551);
xor U21684 (N_21684,N_21589,N_21028);
nand U21685 (N_21685,N_21344,N_21149);
nand U21686 (N_21686,N_21306,N_21230);
or U21687 (N_21687,N_21162,N_21527);
and U21688 (N_21688,N_21003,N_21073);
nor U21689 (N_21689,N_21178,N_21410);
or U21690 (N_21690,N_21292,N_21140);
and U21691 (N_21691,N_21055,N_21168);
or U21692 (N_21692,N_21415,N_21013);
nand U21693 (N_21693,N_21186,N_21496);
nand U21694 (N_21694,N_21451,N_21307);
nor U21695 (N_21695,N_21575,N_21064);
and U21696 (N_21696,N_21098,N_21375);
nand U21697 (N_21697,N_21450,N_21320);
nand U21698 (N_21698,N_21420,N_21297);
nor U21699 (N_21699,N_21112,N_21289);
and U21700 (N_21700,N_21383,N_21199);
or U21701 (N_21701,N_21574,N_21172);
nor U21702 (N_21702,N_21385,N_21021);
nand U21703 (N_21703,N_21009,N_21590);
or U21704 (N_21704,N_21024,N_21148);
xnor U21705 (N_21705,N_21597,N_21235);
nor U21706 (N_21706,N_21117,N_21409);
or U21707 (N_21707,N_21120,N_21395);
xor U21708 (N_21708,N_21015,N_21092);
and U21709 (N_21709,N_21503,N_21276);
or U21710 (N_21710,N_21097,N_21545);
or U21711 (N_21711,N_21341,N_21104);
or U21712 (N_21712,N_21185,N_21537);
nand U21713 (N_21713,N_21020,N_21007);
nor U21714 (N_21714,N_21330,N_21173);
nand U21715 (N_21715,N_21271,N_21225);
nand U21716 (N_21716,N_21340,N_21491);
nand U21717 (N_21717,N_21403,N_21563);
nor U21718 (N_21718,N_21048,N_21267);
xor U21719 (N_21719,N_21184,N_21257);
or U21720 (N_21720,N_21571,N_21314);
or U21721 (N_21721,N_21347,N_21430);
and U21722 (N_21722,N_21434,N_21253);
nand U21723 (N_21723,N_21045,N_21224);
xor U21724 (N_21724,N_21473,N_21331);
nand U21725 (N_21725,N_21146,N_21285);
or U21726 (N_21726,N_21499,N_21443);
nor U21727 (N_21727,N_21300,N_21324);
xnor U21728 (N_21728,N_21558,N_21061);
xnor U21729 (N_21729,N_21259,N_21256);
or U21730 (N_21730,N_21222,N_21019);
or U21731 (N_21731,N_21431,N_21298);
nor U21732 (N_21732,N_21111,N_21529);
or U21733 (N_21733,N_21165,N_21326);
or U21734 (N_21734,N_21226,N_21479);
nor U21735 (N_21735,N_21158,N_21244);
nor U21736 (N_21736,N_21594,N_21317);
xor U21737 (N_21737,N_21573,N_21126);
xnor U21738 (N_21738,N_21490,N_21448);
xor U21739 (N_21739,N_21481,N_21068);
nand U21740 (N_21740,N_21467,N_21002);
xnor U21741 (N_21741,N_21062,N_21572);
nor U21742 (N_21742,N_21220,N_21429);
nor U21743 (N_21743,N_21277,N_21036);
nand U21744 (N_21744,N_21242,N_21005);
and U21745 (N_21745,N_21396,N_21241);
nand U21746 (N_21746,N_21338,N_21110);
xor U21747 (N_21747,N_21380,N_21303);
nor U21748 (N_21748,N_21504,N_21090);
nor U21749 (N_21749,N_21123,N_21493);
and U21750 (N_21750,N_21401,N_21436);
nor U21751 (N_21751,N_21171,N_21052);
and U21752 (N_21752,N_21564,N_21519);
nand U21753 (N_21753,N_21163,N_21311);
or U21754 (N_21754,N_21078,N_21494);
and U21755 (N_21755,N_21555,N_21355);
and U21756 (N_21756,N_21382,N_21044);
nand U21757 (N_21757,N_21492,N_21213);
nand U21758 (N_21758,N_21407,N_21386);
nand U21759 (N_21759,N_21151,N_21025);
xnor U21760 (N_21760,N_21446,N_21261);
or U21761 (N_21761,N_21514,N_21000);
and U21762 (N_21762,N_21296,N_21014);
nor U21763 (N_21763,N_21423,N_21294);
nor U21764 (N_21764,N_21460,N_21387);
xor U21765 (N_21765,N_21077,N_21510);
and U21766 (N_21766,N_21568,N_21031);
or U21767 (N_21767,N_21456,N_21428);
or U21768 (N_21768,N_21084,N_21483);
and U21769 (N_21769,N_21581,N_21398);
nor U21770 (N_21770,N_21312,N_21001);
nor U21771 (N_21771,N_21541,N_21308);
xor U21772 (N_21772,N_21304,N_21548);
nor U21773 (N_21773,N_21121,N_21130);
xnor U21774 (N_21774,N_21240,N_21017);
and U21775 (N_21775,N_21576,N_21250);
or U21776 (N_21776,N_21502,N_21177);
nand U21777 (N_21777,N_21232,N_21295);
nand U21778 (N_21778,N_21405,N_21360);
and U21779 (N_21779,N_21248,N_21166);
or U21780 (N_21780,N_21154,N_21543);
nor U21781 (N_21781,N_21547,N_21245);
and U21782 (N_21782,N_21318,N_21183);
xor U21783 (N_21783,N_21016,N_21161);
xor U21784 (N_21784,N_21560,N_21012);
and U21785 (N_21785,N_21249,N_21262);
nor U21786 (N_21786,N_21378,N_21066);
nor U21787 (N_21787,N_21440,N_21349);
or U21788 (N_21788,N_21287,N_21516);
and U21789 (N_21789,N_21139,N_21343);
xor U21790 (N_21790,N_21365,N_21505);
nor U21791 (N_21791,N_21182,N_21528);
xnor U21792 (N_21792,N_21145,N_21419);
nand U21793 (N_21793,N_21480,N_21010);
nor U21794 (N_21794,N_21023,N_21539);
xnor U21795 (N_21795,N_21498,N_21206);
or U21796 (N_21796,N_21187,N_21034);
or U21797 (N_21797,N_21421,N_21532);
nand U21798 (N_21798,N_21583,N_21147);
or U21799 (N_21799,N_21246,N_21118);
xnor U21800 (N_21800,N_21391,N_21438);
nor U21801 (N_21801,N_21582,N_21439);
or U21802 (N_21802,N_21336,N_21278);
and U21803 (N_21803,N_21208,N_21337);
or U21804 (N_21804,N_21339,N_21374);
and U21805 (N_21805,N_21114,N_21414);
or U21806 (N_21806,N_21557,N_21093);
nor U21807 (N_21807,N_21508,N_21091);
nand U21808 (N_21808,N_21113,N_21228);
nand U21809 (N_21809,N_21458,N_21155);
xor U21810 (N_21810,N_21279,N_21038);
nand U21811 (N_21811,N_21486,N_21323);
xor U21812 (N_21812,N_21302,N_21533);
xor U21813 (N_21813,N_21191,N_21301);
or U21814 (N_21814,N_21471,N_21196);
nand U21815 (N_21815,N_21437,N_21305);
nand U21816 (N_21816,N_21346,N_21353);
nor U21817 (N_21817,N_21237,N_21083);
nand U21818 (N_21818,N_21134,N_21426);
xnor U21819 (N_21819,N_21379,N_21065);
or U21820 (N_21820,N_21591,N_21469);
nand U21821 (N_21821,N_21457,N_21116);
xor U21822 (N_21822,N_21452,N_21517);
xor U21823 (N_21823,N_21050,N_21442);
nor U21824 (N_21824,N_21100,N_21074);
or U21825 (N_21825,N_21231,N_21404);
and U21826 (N_21826,N_21063,N_21465);
and U21827 (N_21827,N_21361,N_21179);
and U21828 (N_21828,N_21076,N_21565);
or U21829 (N_21829,N_21129,N_21596);
nor U21830 (N_21830,N_21004,N_21201);
xor U21831 (N_21831,N_21359,N_21035);
and U21832 (N_21832,N_21132,N_21523);
and U21833 (N_21833,N_21399,N_21585);
or U21834 (N_21834,N_21354,N_21566);
nor U21835 (N_21835,N_21263,N_21188);
and U21836 (N_21836,N_21453,N_21275);
or U21837 (N_21837,N_21103,N_21515);
nor U21838 (N_21838,N_21540,N_21310);
and U21839 (N_21839,N_21234,N_21280);
nor U21840 (N_21840,N_21086,N_21193);
nor U21841 (N_21841,N_21552,N_21071);
xnor U21842 (N_21842,N_21150,N_21152);
xor U21843 (N_21843,N_21269,N_21033);
nor U21844 (N_21844,N_21284,N_21127);
nand U21845 (N_21845,N_21580,N_21264);
nand U21846 (N_21846,N_21288,N_21203);
nand U21847 (N_21847,N_21070,N_21367);
and U21848 (N_21848,N_21109,N_21377);
or U21849 (N_21849,N_21037,N_21133);
nor U21850 (N_21850,N_21018,N_21417);
nor U21851 (N_21851,N_21167,N_21459);
and U21852 (N_21852,N_21282,N_21381);
and U21853 (N_21853,N_21119,N_21082);
xnor U21854 (N_21854,N_21281,N_21531);
nand U21855 (N_21855,N_21595,N_21536);
or U21856 (N_21856,N_21047,N_21598);
xnor U21857 (N_21857,N_21356,N_21416);
or U21858 (N_21858,N_21489,N_21319);
xnor U21859 (N_21859,N_21567,N_21138);
or U21860 (N_21860,N_21258,N_21094);
xnor U21861 (N_21861,N_21366,N_21273);
or U21862 (N_21862,N_21334,N_21040);
nand U21863 (N_21863,N_21570,N_21229);
nand U21864 (N_21864,N_21569,N_21046);
xor U21865 (N_21865,N_21444,N_21079);
nor U21866 (N_21866,N_21335,N_21497);
nor U21867 (N_21867,N_21389,N_21554);
nand U21868 (N_21868,N_21518,N_21106);
or U21869 (N_21869,N_21265,N_21190);
and U21870 (N_21870,N_21105,N_21221);
xnor U21871 (N_21871,N_21143,N_21268);
xnor U21872 (N_21872,N_21435,N_21538);
nand U21873 (N_21873,N_21219,N_21397);
and U21874 (N_21874,N_21085,N_21056);
or U21875 (N_21875,N_21286,N_21205);
xor U21876 (N_21876,N_21393,N_21402);
nor U21877 (N_21877,N_21412,N_21522);
and U21878 (N_21878,N_21207,N_21260);
xnor U21879 (N_21879,N_21593,N_21520);
nand U21880 (N_21880,N_21218,N_21464);
nand U21881 (N_21881,N_21137,N_21592);
nand U21882 (N_21882,N_21029,N_21157);
and U21883 (N_21883,N_21059,N_21332);
nor U21884 (N_21884,N_21198,N_21394);
nor U21885 (N_21885,N_21026,N_21108);
or U21886 (N_21886,N_21424,N_21390);
nand U21887 (N_21887,N_21125,N_21427);
and U21888 (N_21888,N_21238,N_21192);
xor U21889 (N_21889,N_21081,N_21270);
nand U21890 (N_21890,N_21239,N_21254);
nor U21891 (N_21891,N_21180,N_21362);
and U21892 (N_21892,N_21525,N_21433);
xor U21893 (N_21893,N_21216,N_21011);
nand U21894 (N_21894,N_21329,N_21478);
nor U21895 (N_21895,N_21461,N_21102);
or U21896 (N_21896,N_21144,N_21562);
xor U21897 (N_21897,N_21373,N_21501);
nand U21898 (N_21898,N_21351,N_21588);
nand U21899 (N_21899,N_21475,N_21561);
xnor U21900 (N_21900,N_21206,N_21329);
or U21901 (N_21901,N_21099,N_21217);
or U21902 (N_21902,N_21421,N_21086);
or U21903 (N_21903,N_21421,N_21471);
or U21904 (N_21904,N_21114,N_21177);
nor U21905 (N_21905,N_21507,N_21035);
xnor U21906 (N_21906,N_21154,N_21189);
or U21907 (N_21907,N_21467,N_21478);
nor U21908 (N_21908,N_21558,N_21442);
xor U21909 (N_21909,N_21262,N_21358);
and U21910 (N_21910,N_21441,N_21039);
xor U21911 (N_21911,N_21262,N_21467);
nor U21912 (N_21912,N_21596,N_21239);
or U21913 (N_21913,N_21181,N_21105);
nor U21914 (N_21914,N_21133,N_21129);
nor U21915 (N_21915,N_21515,N_21460);
nand U21916 (N_21916,N_21367,N_21170);
and U21917 (N_21917,N_21569,N_21329);
nand U21918 (N_21918,N_21453,N_21244);
xor U21919 (N_21919,N_21405,N_21341);
or U21920 (N_21920,N_21496,N_21165);
nand U21921 (N_21921,N_21334,N_21095);
nor U21922 (N_21922,N_21480,N_21503);
or U21923 (N_21923,N_21541,N_21217);
or U21924 (N_21924,N_21547,N_21584);
xor U21925 (N_21925,N_21122,N_21127);
nand U21926 (N_21926,N_21203,N_21222);
nand U21927 (N_21927,N_21555,N_21458);
nand U21928 (N_21928,N_21382,N_21140);
or U21929 (N_21929,N_21167,N_21242);
and U21930 (N_21930,N_21260,N_21474);
or U21931 (N_21931,N_21325,N_21169);
xnor U21932 (N_21932,N_21452,N_21401);
or U21933 (N_21933,N_21276,N_21100);
nor U21934 (N_21934,N_21219,N_21468);
nor U21935 (N_21935,N_21525,N_21524);
and U21936 (N_21936,N_21505,N_21005);
nor U21937 (N_21937,N_21581,N_21228);
xnor U21938 (N_21938,N_21383,N_21499);
or U21939 (N_21939,N_21562,N_21006);
or U21940 (N_21940,N_21500,N_21009);
nand U21941 (N_21941,N_21394,N_21056);
nor U21942 (N_21942,N_21401,N_21065);
nand U21943 (N_21943,N_21545,N_21222);
nand U21944 (N_21944,N_21511,N_21102);
nand U21945 (N_21945,N_21341,N_21365);
or U21946 (N_21946,N_21223,N_21451);
nand U21947 (N_21947,N_21502,N_21058);
or U21948 (N_21948,N_21209,N_21001);
xor U21949 (N_21949,N_21061,N_21044);
or U21950 (N_21950,N_21574,N_21039);
nand U21951 (N_21951,N_21583,N_21102);
and U21952 (N_21952,N_21469,N_21252);
nand U21953 (N_21953,N_21068,N_21331);
xor U21954 (N_21954,N_21314,N_21187);
nand U21955 (N_21955,N_21267,N_21178);
and U21956 (N_21956,N_21264,N_21144);
and U21957 (N_21957,N_21039,N_21489);
nand U21958 (N_21958,N_21092,N_21473);
and U21959 (N_21959,N_21378,N_21295);
xnor U21960 (N_21960,N_21221,N_21347);
nand U21961 (N_21961,N_21189,N_21166);
nand U21962 (N_21962,N_21350,N_21496);
xnor U21963 (N_21963,N_21191,N_21562);
or U21964 (N_21964,N_21348,N_21552);
nand U21965 (N_21965,N_21595,N_21309);
or U21966 (N_21966,N_21518,N_21001);
nor U21967 (N_21967,N_21222,N_21445);
nor U21968 (N_21968,N_21381,N_21437);
nor U21969 (N_21969,N_21051,N_21491);
nand U21970 (N_21970,N_21490,N_21583);
or U21971 (N_21971,N_21544,N_21139);
nand U21972 (N_21972,N_21238,N_21206);
or U21973 (N_21973,N_21494,N_21235);
or U21974 (N_21974,N_21358,N_21053);
xor U21975 (N_21975,N_21557,N_21213);
xor U21976 (N_21976,N_21337,N_21433);
nor U21977 (N_21977,N_21219,N_21531);
or U21978 (N_21978,N_21304,N_21148);
or U21979 (N_21979,N_21035,N_21054);
or U21980 (N_21980,N_21171,N_21188);
nand U21981 (N_21981,N_21233,N_21515);
nand U21982 (N_21982,N_21426,N_21110);
xor U21983 (N_21983,N_21551,N_21074);
and U21984 (N_21984,N_21198,N_21038);
nor U21985 (N_21985,N_21429,N_21033);
xor U21986 (N_21986,N_21025,N_21083);
or U21987 (N_21987,N_21504,N_21391);
or U21988 (N_21988,N_21265,N_21254);
or U21989 (N_21989,N_21244,N_21181);
nor U21990 (N_21990,N_21400,N_21412);
or U21991 (N_21991,N_21582,N_21346);
nand U21992 (N_21992,N_21304,N_21456);
nand U21993 (N_21993,N_21442,N_21216);
nand U21994 (N_21994,N_21281,N_21529);
xnor U21995 (N_21995,N_21400,N_21322);
nor U21996 (N_21996,N_21566,N_21307);
xor U21997 (N_21997,N_21235,N_21095);
or U21998 (N_21998,N_21406,N_21028);
and U21999 (N_21999,N_21313,N_21558);
and U22000 (N_22000,N_21154,N_21517);
nand U22001 (N_22001,N_21006,N_21252);
and U22002 (N_22002,N_21149,N_21506);
nor U22003 (N_22003,N_21559,N_21500);
xor U22004 (N_22004,N_21377,N_21598);
and U22005 (N_22005,N_21180,N_21482);
nand U22006 (N_22006,N_21393,N_21345);
and U22007 (N_22007,N_21061,N_21489);
xor U22008 (N_22008,N_21254,N_21436);
and U22009 (N_22009,N_21148,N_21598);
nand U22010 (N_22010,N_21016,N_21227);
or U22011 (N_22011,N_21589,N_21375);
nor U22012 (N_22012,N_21219,N_21476);
and U22013 (N_22013,N_21296,N_21270);
xnor U22014 (N_22014,N_21219,N_21071);
or U22015 (N_22015,N_21439,N_21318);
xor U22016 (N_22016,N_21016,N_21081);
nand U22017 (N_22017,N_21071,N_21111);
nand U22018 (N_22018,N_21355,N_21069);
xnor U22019 (N_22019,N_21191,N_21178);
nand U22020 (N_22020,N_21099,N_21115);
nand U22021 (N_22021,N_21371,N_21160);
nor U22022 (N_22022,N_21424,N_21498);
and U22023 (N_22023,N_21251,N_21086);
or U22024 (N_22024,N_21344,N_21514);
nor U22025 (N_22025,N_21370,N_21537);
xor U22026 (N_22026,N_21474,N_21512);
nor U22027 (N_22027,N_21527,N_21279);
xor U22028 (N_22028,N_21561,N_21195);
nand U22029 (N_22029,N_21490,N_21047);
nor U22030 (N_22030,N_21490,N_21596);
nand U22031 (N_22031,N_21202,N_21197);
and U22032 (N_22032,N_21065,N_21597);
or U22033 (N_22033,N_21490,N_21250);
nor U22034 (N_22034,N_21115,N_21294);
nor U22035 (N_22035,N_21511,N_21201);
xnor U22036 (N_22036,N_21285,N_21042);
or U22037 (N_22037,N_21522,N_21405);
nand U22038 (N_22038,N_21490,N_21366);
or U22039 (N_22039,N_21446,N_21310);
nor U22040 (N_22040,N_21212,N_21051);
or U22041 (N_22041,N_21477,N_21393);
and U22042 (N_22042,N_21395,N_21407);
and U22043 (N_22043,N_21267,N_21086);
nor U22044 (N_22044,N_21161,N_21403);
xor U22045 (N_22045,N_21466,N_21396);
nand U22046 (N_22046,N_21119,N_21316);
nand U22047 (N_22047,N_21308,N_21504);
nand U22048 (N_22048,N_21238,N_21392);
nand U22049 (N_22049,N_21558,N_21148);
nand U22050 (N_22050,N_21005,N_21307);
nand U22051 (N_22051,N_21555,N_21168);
nor U22052 (N_22052,N_21359,N_21403);
or U22053 (N_22053,N_21446,N_21540);
xor U22054 (N_22054,N_21082,N_21231);
and U22055 (N_22055,N_21271,N_21422);
and U22056 (N_22056,N_21175,N_21075);
nand U22057 (N_22057,N_21560,N_21312);
and U22058 (N_22058,N_21152,N_21116);
and U22059 (N_22059,N_21330,N_21586);
or U22060 (N_22060,N_21156,N_21325);
xnor U22061 (N_22061,N_21013,N_21438);
or U22062 (N_22062,N_21090,N_21480);
nor U22063 (N_22063,N_21110,N_21262);
and U22064 (N_22064,N_21329,N_21200);
or U22065 (N_22065,N_21460,N_21419);
and U22066 (N_22066,N_21008,N_21505);
xor U22067 (N_22067,N_21118,N_21334);
nor U22068 (N_22068,N_21521,N_21055);
nor U22069 (N_22069,N_21475,N_21263);
or U22070 (N_22070,N_21250,N_21523);
nand U22071 (N_22071,N_21256,N_21401);
nand U22072 (N_22072,N_21400,N_21495);
nand U22073 (N_22073,N_21416,N_21305);
or U22074 (N_22074,N_21044,N_21040);
xnor U22075 (N_22075,N_21507,N_21180);
nand U22076 (N_22076,N_21028,N_21521);
xnor U22077 (N_22077,N_21044,N_21558);
xor U22078 (N_22078,N_21138,N_21324);
xor U22079 (N_22079,N_21239,N_21494);
nor U22080 (N_22080,N_21351,N_21251);
or U22081 (N_22081,N_21415,N_21381);
nand U22082 (N_22082,N_21487,N_21097);
nand U22083 (N_22083,N_21000,N_21446);
xnor U22084 (N_22084,N_21489,N_21238);
nor U22085 (N_22085,N_21407,N_21126);
nand U22086 (N_22086,N_21065,N_21212);
nand U22087 (N_22087,N_21293,N_21276);
and U22088 (N_22088,N_21227,N_21189);
nor U22089 (N_22089,N_21524,N_21272);
or U22090 (N_22090,N_21277,N_21070);
nand U22091 (N_22091,N_21478,N_21385);
nand U22092 (N_22092,N_21138,N_21449);
nor U22093 (N_22093,N_21482,N_21509);
nand U22094 (N_22094,N_21530,N_21023);
or U22095 (N_22095,N_21416,N_21119);
nor U22096 (N_22096,N_21356,N_21086);
and U22097 (N_22097,N_21227,N_21304);
or U22098 (N_22098,N_21416,N_21143);
xnor U22099 (N_22099,N_21432,N_21421);
or U22100 (N_22100,N_21472,N_21072);
nand U22101 (N_22101,N_21469,N_21416);
xor U22102 (N_22102,N_21563,N_21169);
or U22103 (N_22103,N_21149,N_21461);
nand U22104 (N_22104,N_21423,N_21235);
and U22105 (N_22105,N_21349,N_21463);
xnor U22106 (N_22106,N_21548,N_21388);
or U22107 (N_22107,N_21054,N_21130);
or U22108 (N_22108,N_21311,N_21074);
xnor U22109 (N_22109,N_21106,N_21324);
xnor U22110 (N_22110,N_21484,N_21201);
nand U22111 (N_22111,N_21128,N_21104);
nand U22112 (N_22112,N_21548,N_21576);
or U22113 (N_22113,N_21032,N_21030);
or U22114 (N_22114,N_21247,N_21432);
and U22115 (N_22115,N_21006,N_21320);
nor U22116 (N_22116,N_21225,N_21081);
or U22117 (N_22117,N_21333,N_21095);
or U22118 (N_22118,N_21521,N_21248);
xor U22119 (N_22119,N_21406,N_21576);
and U22120 (N_22120,N_21303,N_21058);
xor U22121 (N_22121,N_21073,N_21040);
nand U22122 (N_22122,N_21314,N_21393);
xor U22123 (N_22123,N_21296,N_21482);
nor U22124 (N_22124,N_21556,N_21121);
nor U22125 (N_22125,N_21393,N_21059);
nor U22126 (N_22126,N_21241,N_21049);
nor U22127 (N_22127,N_21429,N_21062);
or U22128 (N_22128,N_21251,N_21158);
and U22129 (N_22129,N_21535,N_21021);
xor U22130 (N_22130,N_21349,N_21536);
or U22131 (N_22131,N_21292,N_21109);
and U22132 (N_22132,N_21484,N_21020);
or U22133 (N_22133,N_21037,N_21497);
nand U22134 (N_22134,N_21086,N_21572);
nor U22135 (N_22135,N_21396,N_21424);
xnor U22136 (N_22136,N_21233,N_21374);
nand U22137 (N_22137,N_21126,N_21278);
and U22138 (N_22138,N_21176,N_21402);
nand U22139 (N_22139,N_21299,N_21091);
or U22140 (N_22140,N_21444,N_21513);
nand U22141 (N_22141,N_21327,N_21238);
or U22142 (N_22142,N_21116,N_21167);
and U22143 (N_22143,N_21117,N_21555);
xnor U22144 (N_22144,N_21307,N_21311);
nand U22145 (N_22145,N_21230,N_21202);
or U22146 (N_22146,N_21383,N_21227);
or U22147 (N_22147,N_21377,N_21083);
or U22148 (N_22148,N_21316,N_21071);
or U22149 (N_22149,N_21308,N_21497);
and U22150 (N_22150,N_21538,N_21187);
and U22151 (N_22151,N_21253,N_21575);
nand U22152 (N_22152,N_21083,N_21440);
nand U22153 (N_22153,N_21036,N_21057);
and U22154 (N_22154,N_21319,N_21369);
or U22155 (N_22155,N_21424,N_21399);
or U22156 (N_22156,N_21352,N_21236);
nor U22157 (N_22157,N_21145,N_21026);
xor U22158 (N_22158,N_21530,N_21270);
or U22159 (N_22159,N_21510,N_21150);
nor U22160 (N_22160,N_21583,N_21409);
nor U22161 (N_22161,N_21209,N_21338);
xnor U22162 (N_22162,N_21495,N_21313);
nand U22163 (N_22163,N_21181,N_21095);
nand U22164 (N_22164,N_21378,N_21257);
xor U22165 (N_22165,N_21006,N_21497);
or U22166 (N_22166,N_21188,N_21013);
or U22167 (N_22167,N_21536,N_21529);
nand U22168 (N_22168,N_21511,N_21532);
nor U22169 (N_22169,N_21593,N_21363);
nand U22170 (N_22170,N_21245,N_21225);
nand U22171 (N_22171,N_21178,N_21033);
nand U22172 (N_22172,N_21504,N_21560);
nor U22173 (N_22173,N_21531,N_21113);
or U22174 (N_22174,N_21013,N_21387);
nand U22175 (N_22175,N_21369,N_21047);
and U22176 (N_22176,N_21342,N_21063);
nand U22177 (N_22177,N_21067,N_21018);
nor U22178 (N_22178,N_21539,N_21279);
xnor U22179 (N_22179,N_21085,N_21223);
xor U22180 (N_22180,N_21586,N_21149);
nor U22181 (N_22181,N_21551,N_21201);
nor U22182 (N_22182,N_21165,N_21440);
xnor U22183 (N_22183,N_21521,N_21067);
nand U22184 (N_22184,N_21268,N_21397);
nand U22185 (N_22185,N_21337,N_21202);
nor U22186 (N_22186,N_21102,N_21331);
or U22187 (N_22187,N_21153,N_21276);
or U22188 (N_22188,N_21024,N_21129);
and U22189 (N_22189,N_21364,N_21055);
and U22190 (N_22190,N_21112,N_21045);
xor U22191 (N_22191,N_21465,N_21594);
and U22192 (N_22192,N_21129,N_21583);
nand U22193 (N_22193,N_21569,N_21518);
and U22194 (N_22194,N_21317,N_21212);
xor U22195 (N_22195,N_21324,N_21402);
and U22196 (N_22196,N_21477,N_21123);
xor U22197 (N_22197,N_21001,N_21447);
or U22198 (N_22198,N_21124,N_21220);
xnor U22199 (N_22199,N_21008,N_21262);
nor U22200 (N_22200,N_21820,N_21635);
nor U22201 (N_22201,N_22056,N_21710);
nor U22202 (N_22202,N_22191,N_21948);
and U22203 (N_22203,N_21881,N_22142);
xnor U22204 (N_22204,N_22045,N_21852);
nor U22205 (N_22205,N_21691,N_21883);
and U22206 (N_22206,N_22013,N_22090);
nor U22207 (N_22207,N_21799,N_21938);
and U22208 (N_22208,N_21681,N_21798);
and U22209 (N_22209,N_21833,N_21665);
xor U22210 (N_22210,N_22131,N_21625);
nand U22211 (N_22211,N_21991,N_21807);
and U22212 (N_22212,N_21687,N_22148);
nor U22213 (N_22213,N_22019,N_21740);
nor U22214 (N_22214,N_21651,N_21742);
or U22215 (N_22215,N_21673,N_21850);
nand U22216 (N_22216,N_21660,N_21616);
or U22217 (N_22217,N_21677,N_22101);
nand U22218 (N_22218,N_21893,N_21679);
nand U22219 (N_22219,N_21809,N_21849);
or U22220 (N_22220,N_21769,N_22020);
nor U22221 (N_22221,N_21767,N_22181);
xnor U22222 (N_22222,N_22168,N_21810);
nand U22223 (N_22223,N_21964,N_22034);
or U22224 (N_22224,N_21856,N_22081);
nand U22225 (N_22225,N_21613,N_21689);
xnor U22226 (N_22226,N_22152,N_22102);
nor U22227 (N_22227,N_22130,N_21996);
xor U22228 (N_22228,N_21933,N_22033);
or U22229 (N_22229,N_21756,N_21955);
and U22230 (N_22230,N_21664,N_22193);
nand U22231 (N_22231,N_21715,N_21828);
xnor U22232 (N_22232,N_22080,N_21984);
nor U22233 (N_22233,N_21792,N_22150);
xnor U22234 (N_22234,N_21618,N_21992);
nand U22235 (N_22235,N_21790,N_22064);
and U22236 (N_22236,N_21644,N_21844);
nand U22237 (N_22237,N_21789,N_21954);
and U22238 (N_22238,N_21752,N_21650);
and U22239 (N_22239,N_21877,N_21979);
and U22240 (N_22240,N_22057,N_22071);
nor U22241 (N_22241,N_21997,N_21903);
nor U22242 (N_22242,N_21732,N_21894);
nand U22243 (N_22243,N_21880,N_21686);
nand U22244 (N_22244,N_22001,N_22067);
xor U22245 (N_22245,N_21939,N_21861);
nor U22246 (N_22246,N_21629,N_21912);
nor U22247 (N_22247,N_21859,N_21985);
and U22248 (N_22248,N_21796,N_21794);
or U22249 (N_22249,N_22197,N_21649);
or U22250 (N_22250,N_21653,N_21899);
xnor U22251 (N_22251,N_21693,N_21608);
xor U22252 (N_22252,N_22109,N_21908);
or U22253 (N_22253,N_21842,N_21812);
or U22254 (N_22254,N_21944,N_21662);
xnor U22255 (N_22255,N_22117,N_22156);
or U22256 (N_22256,N_21940,N_21659);
nand U22257 (N_22257,N_21895,N_21970);
nor U22258 (N_22258,N_22073,N_21669);
xor U22259 (N_22259,N_21619,N_21860);
nor U22260 (N_22260,N_21879,N_21995);
and U22261 (N_22261,N_21676,N_21874);
xnor U22262 (N_22262,N_21834,N_21617);
or U22263 (N_22263,N_21943,N_21823);
nor U22264 (N_22264,N_21962,N_21734);
or U22265 (N_22265,N_21873,N_21657);
or U22266 (N_22266,N_21921,N_22084);
or U22267 (N_22267,N_21890,N_21813);
nor U22268 (N_22268,N_22118,N_21675);
xor U22269 (N_22269,N_21994,N_21902);
or U22270 (N_22270,N_22079,N_21897);
nor U22271 (N_22271,N_21727,N_21785);
nand U22272 (N_22272,N_22059,N_21947);
nand U22273 (N_22273,N_21671,N_21911);
nand U22274 (N_22274,N_21950,N_22053);
xor U22275 (N_22275,N_22078,N_22014);
nor U22276 (N_22276,N_21696,N_21806);
nor U22277 (N_22277,N_22027,N_22082);
or U22278 (N_22278,N_21942,N_21776);
nor U22279 (N_22279,N_21631,N_22002);
nor U22280 (N_22280,N_21999,N_21854);
nand U22281 (N_22281,N_22055,N_21763);
and U22282 (N_22282,N_21887,N_21885);
xnor U22283 (N_22283,N_21772,N_21712);
nor U22284 (N_22284,N_21723,N_21827);
xor U22285 (N_22285,N_22198,N_21980);
nand U22286 (N_22286,N_22030,N_21698);
xor U22287 (N_22287,N_22098,N_21972);
xor U22288 (N_22288,N_21878,N_21977);
and U22289 (N_22289,N_21661,N_22041);
and U22290 (N_22290,N_22010,N_21602);
and U22291 (N_22291,N_22087,N_21843);
and U22292 (N_22292,N_22186,N_21835);
nand U22293 (N_22293,N_22077,N_21803);
nand U22294 (N_22294,N_21620,N_22112);
nor U22295 (N_22295,N_21937,N_22066);
nand U22296 (N_22296,N_22173,N_22177);
or U22297 (N_22297,N_22011,N_22089);
and U22298 (N_22298,N_21925,N_21765);
xor U22299 (N_22299,N_22012,N_21853);
xnor U22300 (N_22300,N_21837,N_21869);
xnor U22301 (N_22301,N_21986,N_21720);
and U22302 (N_22302,N_21845,N_21915);
and U22303 (N_22303,N_21703,N_21728);
xnor U22304 (N_22304,N_21857,N_22110);
or U22305 (N_22305,N_22021,N_22141);
nor U22306 (N_22306,N_21634,N_21805);
xnor U22307 (N_22307,N_21927,N_22192);
nor U22308 (N_22308,N_21919,N_22037);
xnor U22309 (N_22309,N_21808,N_21697);
xor U22310 (N_22310,N_21655,N_21847);
and U22311 (N_22311,N_21797,N_22040);
and U22312 (N_22312,N_22175,N_22017);
or U22313 (N_22313,N_22190,N_21988);
and U22314 (N_22314,N_21678,N_21882);
xor U22315 (N_22315,N_21910,N_21817);
nor U22316 (N_22316,N_22157,N_21858);
xor U22317 (N_22317,N_21783,N_21735);
and U22318 (N_22318,N_21707,N_21758);
or U22319 (N_22319,N_21876,N_22094);
nand U22320 (N_22320,N_22184,N_21917);
xnor U22321 (N_22321,N_21802,N_22196);
nand U22322 (N_22322,N_21747,N_22035);
nand U22323 (N_22323,N_22006,N_21738);
and U22324 (N_22324,N_22129,N_22183);
nand U22325 (N_22325,N_22029,N_21666);
and U22326 (N_22326,N_22144,N_21609);
or U22327 (N_22327,N_22049,N_21941);
and U22328 (N_22328,N_21682,N_21952);
nor U22329 (N_22329,N_21801,N_21713);
xor U22330 (N_22330,N_21726,N_22063);
nand U22331 (N_22331,N_22091,N_22106);
xor U22332 (N_22332,N_21993,N_22151);
xor U22333 (N_22333,N_21832,N_22111);
nor U22334 (N_22334,N_21654,N_21975);
nor U22335 (N_22335,N_22194,N_22172);
and U22336 (N_22336,N_21711,N_22134);
or U22337 (N_22337,N_22188,N_22054);
or U22338 (N_22338,N_22036,N_22031);
nor U22339 (N_22339,N_21643,N_21777);
xnor U22340 (N_22340,N_21848,N_22108);
nor U22341 (N_22341,N_21766,N_21830);
or U22342 (N_22342,N_21888,N_21702);
xnor U22343 (N_22343,N_22143,N_22114);
nand U22344 (N_22344,N_22161,N_21709);
nor U22345 (N_22345,N_21627,N_21958);
nand U22346 (N_22346,N_21974,N_21824);
nor U22347 (N_22347,N_22179,N_21749);
nor U22348 (N_22348,N_22024,N_21928);
nor U22349 (N_22349,N_21865,N_21733);
or U22350 (N_22350,N_21829,N_22145);
xnor U22351 (N_22351,N_21922,N_21953);
and U22352 (N_22352,N_21670,N_21804);
nand U22353 (N_22353,N_21757,N_22138);
xnor U22354 (N_22354,N_21648,N_21626);
nor U22355 (N_22355,N_21640,N_21725);
nor U22356 (N_22356,N_21612,N_21998);
nand U22357 (N_22357,N_21892,N_21889);
or U22358 (N_22358,N_22120,N_22003);
nor U22359 (N_22359,N_21755,N_22178);
nand U22360 (N_22360,N_21760,N_21633);
and U22361 (N_22361,N_22038,N_22164);
nand U22362 (N_22362,N_21656,N_21768);
nor U22363 (N_22363,N_21764,N_22126);
xor U22364 (N_22364,N_21621,N_22007);
xor U22365 (N_22365,N_21690,N_21729);
xor U22366 (N_22366,N_22050,N_21864);
and U22367 (N_22367,N_21784,N_21700);
and U22368 (N_22368,N_21736,N_21795);
and U22369 (N_22369,N_21791,N_21632);
or U22370 (N_22370,N_21731,N_21699);
xnor U22371 (N_22371,N_21818,N_21701);
or U22372 (N_22372,N_22018,N_22189);
or U22373 (N_22373,N_21906,N_22122);
nand U22374 (N_22374,N_21914,N_22005);
and U22375 (N_22375,N_22096,N_21672);
nand U22376 (N_22376,N_22076,N_21787);
or U22377 (N_22377,N_22008,N_22167);
or U22378 (N_22378,N_21737,N_22028);
and U22379 (N_22379,N_22169,N_21774);
nand U22380 (N_22380,N_21907,N_21949);
or U22381 (N_22381,N_21923,N_22133);
xor U22382 (N_22382,N_22158,N_21793);
nor U22383 (N_22383,N_21905,N_21788);
and U22384 (N_22384,N_22051,N_22116);
nor U22385 (N_22385,N_21825,N_21770);
nor U22386 (N_22386,N_21934,N_21645);
nand U22387 (N_22387,N_21628,N_21642);
nor U22388 (N_22388,N_21786,N_22100);
or U22389 (N_22389,N_21875,N_21782);
xor U22390 (N_22390,N_21607,N_21983);
xnor U22391 (N_22391,N_21936,N_21603);
or U22392 (N_22392,N_21606,N_22032);
nor U22393 (N_22393,N_21722,N_22170);
xor U22394 (N_22394,N_21694,N_22163);
nor U22395 (N_22395,N_22039,N_21840);
and U22396 (N_22396,N_21667,N_21932);
and U22397 (N_22397,N_21663,N_21615);
nor U22398 (N_22398,N_21967,N_22153);
xor U22399 (N_22399,N_21904,N_21773);
or U22400 (N_22400,N_21704,N_21614);
nand U22401 (N_22401,N_21730,N_22159);
and U22402 (N_22402,N_22058,N_22136);
nor U22403 (N_22403,N_21610,N_22187);
xor U22404 (N_22404,N_22199,N_21945);
nor U22405 (N_22405,N_22155,N_21744);
xnor U22406 (N_22406,N_21674,N_22074);
nor U22407 (N_22407,N_22185,N_22160);
xnor U22408 (N_22408,N_22119,N_21688);
xor U22409 (N_22409,N_22016,N_21990);
or U22410 (N_22410,N_22000,N_21721);
or U22411 (N_22411,N_21963,N_22149);
xnor U22412 (N_22412,N_22086,N_21819);
or U22413 (N_22413,N_21898,N_22061);
nor U22414 (N_22414,N_21901,N_22182);
xor U22415 (N_22415,N_21753,N_21821);
or U22416 (N_22416,N_22171,N_21623);
xnor U22417 (N_22417,N_22115,N_22128);
or U22418 (N_22418,N_21814,N_21826);
xor U22419 (N_22419,N_21636,N_21630);
nand U22420 (N_22420,N_22105,N_21961);
xnor U22421 (N_22421,N_21822,N_21708);
and U22422 (N_22422,N_21855,N_21965);
or U22423 (N_22423,N_21931,N_21868);
nand U22424 (N_22424,N_22047,N_21746);
or U22425 (N_22425,N_21639,N_21761);
xor U22426 (N_22426,N_21989,N_21683);
nor U22427 (N_22427,N_22140,N_21695);
nor U22428 (N_22428,N_22113,N_21692);
nand U22429 (N_22429,N_21816,N_22180);
xor U22430 (N_22430,N_21846,N_21867);
or U22431 (N_22431,N_21982,N_22048);
or U22432 (N_22432,N_21987,N_22043);
and U22433 (N_22433,N_22104,N_21706);
nand U22434 (N_22434,N_21759,N_21771);
nand U22435 (N_22435,N_22022,N_21638);
and U22436 (N_22436,N_21637,N_22097);
nand U22437 (N_22437,N_22135,N_21924);
or U22438 (N_22438,N_21811,N_22068);
and U22439 (N_22439,N_22125,N_22195);
nand U22440 (N_22440,N_21871,N_21971);
and U22441 (N_22441,N_22065,N_22075);
nand U22442 (N_22442,N_21929,N_22015);
nor U22443 (N_22443,N_22044,N_21739);
nand U22444 (N_22444,N_22025,N_21870);
and U22445 (N_22445,N_22103,N_22121);
and U22446 (N_22446,N_21622,N_22004);
nor U22447 (N_22447,N_21668,N_21900);
nor U22448 (N_22448,N_21951,N_21916);
nor U22449 (N_22449,N_22124,N_21946);
nor U22450 (N_22450,N_21745,N_22072);
and U22451 (N_22451,N_22070,N_22099);
nor U22452 (N_22452,N_21913,N_22009);
or U22453 (N_22453,N_21719,N_21762);
or U22454 (N_22454,N_21718,N_21600);
nor U22455 (N_22455,N_22166,N_21641);
or U22456 (N_22456,N_21750,N_22023);
nand U22457 (N_22457,N_21743,N_22042);
nor U22458 (N_22458,N_21866,N_21851);
xor U22459 (N_22459,N_22139,N_22083);
nand U22460 (N_22460,N_21604,N_21935);
and U22461 (N_22461,N_21896,N_22107);
nand U22462 (N_22462,N_22162,N_21966);
or U22463 (N_22463,N_21779,N_21884);
xnor U22464 (N_22464,N_21960,N_21969);
or U22465 (N_22465,N_21716,N_21705);
xnor U22466 (N_22466,N_21959,N_21754);
xor U22467 (N_22467,N_21841,N_21839);
nand U22468 (N_22468,N_21981,N_22092);
nand U22469 (N_22469,N_22060,N_21831);
and U22470 (N_22470,N_21624,N_21973);
nand U22471 (N_22471,N_21714,N_21780);
and U22472 (N_22472,N_22165,N_21930);
nand U22473 (N_22473,N_21976,N_22026);
and U22474 (N_22474,N_21647,N_21652);
and U22475 (N_22475,N_21920,N_21838);
or U22476 (N_22476,N_21800,N_21978);
and U22477 (N_22477,N_21926,N_22046);
and U22478 (N_22478,N_21605,N_22132);
xnor U22479 (N_22479,N_22062,N_22085);
nand U22480 (N_22480,N_22154,N_22174);
and U22481 (N_22481,N_21680,N_22069);
nand U22482 (N_22482,N_21778,N_21601);
and U22483 (N_22483,N_22147,N_21957);
or U22484 (N_22484,N_21751,N_21748);
nand U22485 (N_22485,N_22146,N_22052);
and U22486 (N_22486,N_21836,N_22127);
nor U22487 (N_22487,N_21886,N_21968);
or U22488 (N_22488,N_21684,N_21611);
xnor U22489 (N_22489,N_21918,N_21862);
xnor U22490 (N_22490,N_21724,N_22137);
nor U22491 (N_22491,N_21891,N_21685);
nand U22492 (N_22492,N_21741,N_21775);
or U22493 (N_22493,N_21909,N_21815);
xnor U22494 (N_22494,N_21863,N_22123);
or U22495 (N_22495,N_21872,N_21781);
xor U22496 (N_22496,N_22095,N_22088);
nor U22497 (N_22497,N_21658,N_21646);
nor U22498 (N_22498,N_21717,N_22093);
and U22499 (N_22499,N_22176,N_21956);
and U22500 (N_22500,N_21742,N_22008);
and U22501 (N_22501,N_21955,N_21674);
and U22502 (N_22502,N_21994,N_21638);
xnor U22503 (N_22503,N_22114,N_22082);
nand U22504 (N_22504,N_21673,N_21694);
or U22505 (N_22505,N_22008,N_21642);
nor U22506 (N_22506,N_21732,N_21914);
xnor U22507 (N_22507,N_22051,N_22180);
nand U22508 (N_22508,N_22192,N_22024);
nand U22509 (N_22509,N_22077,N_21723);
nor U22510 (N_22510,N_22148,N_22048);
nor U22511 (N_22511,N_22029,N_21927);
nand U22512 (N_22512,N_21998,N_21680);
and U22513 (N_22513,N_21885,N_22112);
xnor U22514 (N_22514,N_22150,N_21771);
or U22515 (N_22515,N_21736,N_21623);
and U22516 (N_22516,N_21959,N_22191);
nor U22517 (N_22517,N_21650,N_21700);
nand U22518 (N_22518,N_22112,N_22135);
or U22519 (N_22519,N_21889,N_21791);
and U22520 (N_22520,N_21994,N_22014);
or U22521 (N_22521,N_21757,N_21647);
nand U22522 (N_22522,N_21695,N_21895);
nand U22523 (N_22523,N_21699,N_22142);
nand U22524 (N_22524,N_22126,N_21604);
and U22525 (N_22525,N_22185,N_21835);
nor U22526 (N_22526,N_21942,N_22090);
or U22527 (N_22527,N_22000,N_21724);
or U22528 (N_22528,N_21933,N_21819);
xnor U22529 (N_22529,N_21753,N_21954);
nand U22530 (N_22530,N_21879,N_21867);
and U22531 (N_22531,N_22127,N_22097);
and U22532 (N_22532,N_21602,N_21832);
or U22533 (N_22533,N_22127,N_22089);
nor U22534 (N_22534,N_21848,N_21778);
xor U22535 (N_22535,N_22070,N_22114);
or U22536 (N_22536,N_21934,N_21677);
and U22537 (N_22537,N_22159,N_22137);
and U22538 (N_22538,N_21994,N_21926);
nor U22539 (N_22539,N_22198,N_21689);
xnor U22540 (N_22540,N_21926,N_21931);
nor U22541 (N_22541,N_21893,N_21947);
nor U22542 (N_22542,N_21892,N_21776);
xor U22543 (N_22543,N_21704,N_21993);
xnor U22544 (N_22544,N_21788,N_21928);
nand U22545 (N_22545,N_21892,N_22159);
or U22546 (N_22546,N_22167,N_21739);
xnor U22547 (N_22547,N_22047,N_21762);
xnor U22548 (N_22548,N_21848,N_22106);
and U22549 (N_22549,N_22140,N_21799);
and U22550 (N_22550,N_21927,N_21715);
xor U22551 (N_22551,N_21987,N_21602);
nand U22552 (N_22552,N_21762,N_21656);
nor U22553 (N_22553,N_21610,N_22010);
xnor U22554 (N_22554,N_21757,N_22163);
nand U22555 (N_22555,N_21742,N_22065);
xnor U22556 (N_22556,N_21686,N_22066);
xor U22557 (N_22557,N_21772,N_21935);
xor U22558 (N_22558,N_22177,N_21727);
xnor U22559 (N_22559,N_21823,N_22010);
xnor U22560 (N_22560,N_21777,N_21868);
nor U22561 (N_22561,N_21817,N_21781);
and U22562 (N_22562,N_22122,N_21675);
nand U22563 (N_22563,N_22164,N_21936);
nor U22564 (N_22564,N_21947,N_21642);
or U22565 (N_22565,N_21964,N_22074);
nor U22566 (N_22566,N_22141,N_21770);
xnor U22567 (N_22567,N_22076,N_21633);
xor U22568 (N_22568,N_22061,N_22143);
and U22569 (N_22569,N_21896,N_22135);
nor U22570 (N_22570,N_22048,N_22195);
nor U22571 (N_22571,N_21979,N_22133);
or U22572 (N_22572,N_22005,N_21689);
or U22573 (N_22573,N_22041,N_21990);
xnor U22574 (N_22574,N_21622,N_21697);
nand U22575 (N_22575,N_21738,N_21982);
nand U22576 (N_22576,N_21990,N_21660);
nand U22577 (N_22577,N_21689,N_22141);
and U22578 (N_22578,N_22066,N_21638);
or U22579 (N_22579,N_21944,N_21693);
nor U22580 (N_22580,N_21716,N_21740);
nor U22581 (N_22581,N_21759,N_21828);
or U22582 (N_22582,N_21897,N_21704);
or U22583 (N_22583,N_22040,N_22131);
and U22584 (N_22584,N_21856,N_21823);
or U22585 (N_22585,N_21610,N_22164);
and U22586 (N_22586,N_22195,N_22056);
and U22587 (N_22587,N_21738,N_21933);
nand U22588 (N_22588,N_21623,N_22044);
or U22589 (N_22589,N_21692,N_21982);
xor U22590 (N_22590,N_21882,N_22145);
xor U22591 (N_22591,N_21671,N_22164);
or U22592 (N_22592,N_21647,N_21783);
nand U22593 (N_22593,N_21968,N_21779);
or U22594 (N_22594,N_22066,N_22013);
xnor U22595 (N_22595,N_21742,N_22197);
nand U22596 (N_22596,N_21729,N_21657);
and U22597 (N_22597,N_21759,N_22050);
nand U22598 (N_22598,N_21627,N_22127);
nand U22599 (N_22599,N_21862,N_21929);
xnor U22600 (N_22600,N_21716,N_21612);
nor U22601 (N_22601,N_21931,N_21659);
nor U22602 (N_22602,N_21904,N_21628);
nor U22603 (N_22603,N_22075,N_22076);
nor U22604 (N_22604,N_22136,N_21649);
nand U22605 (N_22605,N_21966,N_21883);
nor U22606 (N_22606,N_21733,N_21945);
nand U22607 (N_22607,N_22176,N_22059);
xor U22608 (N_22608,N_22159,N_21847);
nand U22609 (N_22609,N_22091,N_21976);
or U22610 (N_22610,N_21848,N_22105);
nor U22611 (N_22611,N_21828,N_21657);
nand U22612 (N_22612,N_21877,N_21755);
nor U22613 (N_22613,N_21953,N_22010);
nand U22614 (N_22614,N_21723,N_21925);
or U22615 (N_22615,N_22037,N_22159);
or U22616 (N_22616,N_21991,N_21935);
nand U22617 (N_22617,N_21995,N_21627);
or U22618 (N_22618,N_21723,N_21880);
or U22619 (N_22619,N_21948,N_21645);
nand U22620 (N_22620,N_21892,N_21749);
or U22621 (N_22621,N_21984,N_21960);
xor U22622 (N_22622,N_22191,N_22174);
xor U22623 (N_22623,N_22089,N_21652);
or U22624 (N_22624,N_21933,N_21694);
or U22625 (N_22625,N_21621,N_22028);
xor U22626 (N_22626,N_21720,N_21602);
or U22627 (N_22627,N_22189,N_21618);
xor U22628 (N_22628,N_22051,N_22198);
nor U22629 (N_22629,N_21689,N_21777);
nor U22630 (N_22630,N_22171,N_22085);
nor U22631 (N_22631,N_22116,N_22019);
nand U22632 (N_22632,N_22127,N_21673);
nand U22633 (N_22633,N_21915,N_22191);
xor U22634 (N_22634,N_21652,N_21865);
or U22635 (N_22635,N_22112,N_21935);
and U22636 (N_22636,N_21847,N_22177);
and U22637 (N_22637,N_21660,N_22019);
or U22638 (N_22638,N_21863,N_22198);
nand U22639 (N_22639,N_21992,N_21611);
and U22640 (N_22640,N_22035,N_21901);
and U22641 (N_22641,N_22182,N_22177);
xor U22642 (N_22642,N_22012,N_22135);
nand U22643 (N_22643,N_21636,N_21930);
nor U22644 (N_22644,N_22133,N_21745);
nor U22645 (N_22645,N_21727,N_21954);
or U22646 (N_22646,N_22145,N_21903);
xnor U22647 (N_22647,N_21805,N_21654);
nor U22648 (N_22648,N_21681,N_21795);
and U22649 (N_22649,N_21759,N_21946);
or U22650 (N_22650,N_21630,N_21752);
nand U22651 (N_22651,N_21778,N_21926);
nor U22652 (N_22652,N_21800,N_21675);
nor U22653 (N_22653,N_22162,N_21620);
or U22654 (N_22654,N_21985,N_22077);
or U22655 (N_22655,N_22079,N_21856);
nand U22656 (N_22656,N_21999,N_21985);
and U22657 (N_22657,N_21995,N_21826);
or U22658 (N_22658,N_21902,N_22034);
xor U22659 (N_22659,N_21890,N_22059);
nand U22660 (N_22660,N_21838,N_21966);
nand U22661 (N_22661,N_21904,N_22060);
nor U22662 (N_22662,N_21975,N_21871);
and U22663 (N_22663,N_22175,N_21807);
or U22664 (N_22664,N_21907,N_21743);
or U22665 (N_22665,N_22182,N_21854);
nor U22666 (N_22666,N_21736,N_21810);
and U22667 (N_22667,N_22028,N_22127);
or U22668 (N_22668,N_22098,N_21856);
and U22669 (N_22669,N_22010,N_21729);
nor U22670 (N_22670,N_21613,N_22150);
and U22671 (N_22671,N_22118,N_22046);
or U22672 (N_22672,N_21691,N_21698);
or U22673 (N_22673,N_21987,N_21804);
or U22674 (N_22674,N_21675,N_21657);
nand U22675 (N_22675,N_21630,N_22057);
nand U22676 (N_22676,N_21747,N_21692);
nand U22677 (N_22677,N_21713,N_21872);
and U22678 (N_22678,N_22090,N_21691);
xor U22679 (N_22679,N_21759,N_21676);
xnor U22680 (N_22680,N_21708,N_22024);
and U22681 (N_22681,N_21960,N_22060);
nor U22682 (N_22682,N_22096,N_21719);
xor U22683 (N_22683,N_21890,N_21800);
nand U22684 (N_22684,N_21633,N_22000);
nor U22685 (N_22685,N_21732,N_21731);
or U22686 (N_22686,N_21736,N_21678);
xor U22687 (N_22687,N_21856,N_22143);
nor U22688 (N_22688,N_21610,N_21679);
xor U22689 (N_22689,N_21708,N_21610);
and U22690 (N_22690,N_21846,N_21984);
nand U22691 (N_22691,N_21738,N_21820);
or U22692 (N_22692,N_22077,N_22015);
nand U22693 (N_22693,N_22144,N_21726);
and U22694 (N_22694,N_21910,N_22144);
nor U22695 (N_22695,N_21936,N_21666);
nand U22696 (N_22696,N_21668,N_22181);
and U22697 (N_22697,N_21628,N_22159);
xor U22698 (N_22698,N_21765,N_21885);
xor U22699 (N_22699,N_21775,N_21767);
xor U22700 (N_22700,N_22004,N_21858);
nand U22701 (N_22701,N_22157,N_21777);
nor U22702 (N_22702,N_22153,N_22064);
nand U22703 (N_22703,N_22169,N_22052);
or U22704 (N_22704,N_21954,N_21911);
or U22705 (N_22705,N_21646,N_21707);
xor U22706 (N_22706,N_22170,N_21713);
and U22707 (N_22707,N_22116,N_22008);
xor U22708 (N_22708,N_21685,N_22168);
xnor U22709 (N_22709,N_21744,N_21906);
and U22710 (N_22710,N_21650,N_21975);
nor U22711 (N_22711,N_21698,N_21763);
and U22712 (N_22712,N_21964,N_21685);
nor U22713 (N_22713,N_21773,N_21670);
xor U22714 (N_22714,N_21801,N_22120);
nand U22715 (N_22715,N_21883,N_21909);
nand U22716 (N_22716,N_21689,N_22083);
nand U22717 (N_22717,N_21835,N_21976);
and U22718 (N_22718,N_21723,N_22188);
xor U22719 (N_22719,N_21820,N_21772);
nor U22720 (N_22720,N_21884,N_22154);
or U22721 (N_22721,N_22021,N_22128);
and U22722 (N_22722,N_21764,N_21659);
or U22723 (N_22723,N_21989,N_22011);
nor U22724 (N_22724,N_22061,N_22174);
nand U22725 (N_22725,N_21993,N_21904);
and U22726 (N_22726,N_22131,N_22190);
nand U22727 (N_22727,N_21857,N_21648);
xor U22728 (N_22728,N_21792,N_21953);
nor U22729 (N_22729,N_21815,N_22153);
nand U22730 (N_22730,N_22003,N_21745);
and U22731 (N_22731,N_22157,N_21986);
nor U22732 (N_22732,N_22100,N_21627);
and U22733 (N_22733,N_22030,N_21678);
or U22734 (N_22734,N_22032,N_21956);
nor U22735 (N_22735,N_21829,N_21807);
and U22736 (N_22736,N_21832,N_21833);
and U22737 (N_22737,N_22139,N_22065);
and U22738 (N_22738,N_22118,N_21987);
or U22739 (N_22739,N_21821,N_21949);
or U22740 (N_22740,N_21610,N_21663);
or U22741 (N_22741,N_21632,N_21872);
nand U22742 (N_22742,N_21926,N_21645);
nand U22743 (N_22743,N_22018,N_21721);
nand U22744 (N_22744,N_21614,N_21740);
xnor U22745 (N_22745,N_21610,N_22053);
nand U22746 (N_22746,N_22158,N_21808);
nand U22747 (N_22747,N_22103,N_21726);
xnor U22748 (N_22748,N_21855,N_21958);
nand U22749 (N_22749,N_21727,N_21847);
nand U22750 (N_22750,N_21771,N_22112);
and U22751 (N_22751,N_21904,N_21785);
nand U22752 (N_22752,N_22068,N_21825);
nor U22753 (N_22753,N_21724,N_21620);
nand U22754 (N_22754,N_21765,N_21615);
nand U22755 (N_22755,N_21893,N_21877);
nand U22756 (N_22756,N_22087,N_22044);
nor U22757 (N_22757,N_21722,N_21862);
or U22758 (N_22758,N_21902,N_21964);
and U22759 (N_22759,N_21818,N_22180);
nor U22760 (N_22760,N_21995,N_22049);
nor U22761 (N_22761,N_21787,N_21631);
nand U22762 (N_22762,N_22197,N_21936);
nor U22763 (N_22763,N_21927,N_22007);
and U22764 (N_22764,N_22088,N_21800);
or U22765 (N_22765,N_21973,N_21623);
nor U22766 (N_22766,N_21730,N_22019);
and U22767 (N_22767,N_21762,N_22159);
nand U22768 (N_22768,N_22023,N_22167);
xor U22769 (N_22769,N_22088,N_22038);
and U22770 (N_22770,N_21851,N_21952);
xnor U22771 (N_22771,N_22034,N_21863);
and U22772 (N_22772,N_22145,N_22062);
xor U22773 (N_22773,N_21922,N_21734);
and U22774 (N_22774,N_22130,N_21679);
xor U22775 (N_22775,N_21872,N_21942);
nor U22776 (N_22776,N_21962,N_21633);
nand U22777 (N_22777,N_21744,N_21937);
nand U22778 (N_22778,N_21716,N_21850);
nor U22779 (N_22779,N_22049,N_21998);
nand U22780 (N_22780,N_21790,N_21913);
nor U22781 (N_22781,N_21870,N_22056);
xnor U22782 (N_22782,N_21826,N_22178);
and U22783 (N_22783,N_21868,N_21830);
nand U22784 (N_22784,N_21608,N_21743);
or U22785 (N_22785,N_21693,N_22098);
or U22786 (N_22786,N_22192,N_22088);
xnor U22787 (N_22787,N_21893,N_22144);
and U22788 (N_22788,N_21850,N_21672);
nand U22789 (N_22789,N_21998,N_22055);
or U22790 (N_22790,N_21889,N_21608);
nand U22791 (N_22791,N_21881,N_21636);
nor U22792 (N_22792,N_21793,N_22007);
nor U22793 (N_22793,N_22024,N_21656);
xor U22794 (N_22794,N_21858,N_21947);
and U22795 (N_22795,N_21834,N_22022);
or U22796 (N_22796,N_21670,N_22116);
xor U22797 (N_22797,N_22027,N_22140);
and U22798 (N_22798,N_21939,N_21774);
and U22799 (N_22799,N_21687,N_21886);
xor U22800 (N_22800,N_22458,N_22487);
or U22801 (N_22801,N_22402,N_22386);
or U22802 (N_22802,N_22395,N_22226);
or U22803 (N_22803,N_22296,N_22283);
nor U22804 (N_22804,N_22549,N_22624);
xor U22805 (N_22805,N_22761,N_22780);
or U22806 (N_22806,N_22332,N_22443);
nor U22807 (N_22807,N_22415,N_22744);
and U22808 (N_22808,N_22499,N_22786);
nor U22809 (N_22809,N_22542,N_22733);
nor U22810 (N_22810,N_22298,N_22412);
and U22811 (N_22811,N_22358,N_22235);
nand U22812 (N_22812,N_22306,N_22436);
xor U22813 (N_22813,N_22615,N_22308);
and U22814 (N_22814,N_22480,N_22746);
and U22815 (N_22815,N_22470,N_22548);
nor U22816 (N_22816,N_22385,N_22252);
nor U22817 (N_22817,N_22679,N_22785);
nand U22818 (N_22818,N_22322,N_22769);
or U22819 (N_22819,N_22753,N_22242);
nand U22820 (N_22820,N_22715,N_22245);
nor U22821 (N_22821,N_22772,N_22247);
nor U22822 (N_22822,N_22418,N_22609);
xor U22823 (N_22823,N_22474,N_22647);
and U22824 (N_22824,N_22241,N_22616);
xor U22825 (N_22825,N_22633,N_22424);
nand U22826 (N_22826,N_22486,N_22434);
xnor U22827 (N_22827,N_22595,N_22762);
nor U22828 (N_22828,N_22573,N_22777);
nor U22829 (N_22829,N_22462,N_22526);
xor U22830 (N_22830,N_22690,N_22745);
or U22831 (N_22831,N_22676,N_22782);
and U22832 (N_22832,N_22560,N_22380);
or U22833 (N_22833,N_22407,N_22400);
nand U22834 (N_22834,N_22445,N_22209);
xor U22835 (N_22835,N_22796,N_22278);
xnor U22836 (N_22836,N_22569,N_22401);
or U22837 (N_22837,N_22604,N_22637);
or U22838 (N_22838,N_22764,N_22629);
xnor U22839 (N_22839,N_22712,N_22513);
nand U22840 (N_22840,N_22249,N_22288);
nand U22841 (N_22841,N_22724,N_22767);
xnor U22842 (N_22842,N_22580,N_22389);
or U22843 (N_22843,N_22508,N_22422);
and U22844 (N_22844,N_22261,N_22708);
nand U22845 (N_22845,N_22481,N_22693);
nor U22846 (N_22846,N_22632,N_22545);
and U22847 (N_22847,N_22363,N_22246);
nand U22848 (N_22848,N_22509,N_22416);
nand U22849 (N_22849,N_22338,N_22790);
and U22850 (N_22850,N_22641,N_22357);
or U22851 (N_22851,N_22515,N_22531);
nor U22852 (N_22852,N_22506,N_22553);
nand U22853 (N_22853,N_22223,N_22277);
or U22854 (N_22854,N_22546,N_22671);
xor U22855 (N_22855,N_22463,N_22765);
and U22856 (N_22856,N_22397,N_22228);
nand U22857 (N_22857,N_22353,N_22653);
and U22858 (N_22858,N_22367,N_22496);
xor U22859 (N_22859,N_22409,N_22294);
xnor U22860 (N_22860,N_22634,N_22362);
nor U22861 (N_22861,N_22584,N_22649);
xnor U22862 (N_22862,N_22608,N_22378);
or U22863 (N_22863,N_22621,N_22221);
and U22864 (N_22864,N_22320,N_22758);
nand U22865 (N_22865,N_22342,N_22628);
xnor U22866 (N_22866,N_22562,N_22302);
nor U22867 (N_22867,N_22272,N_22340);
or U22868 (N_22868,N_22222,N_22295);
nor U22869 (N_22869,N_22410,N_22469);
or U22870 (N_22870,N_22799,N_22476);
and U22871 (N_22871,N_22328,N_22722);
nand U22872 (N_22872,N_22452,N_22307);
xor U22873 (N_22873,N_22251,N_22279);
and U22874 (N_22874,N_22681,N_22669);
and U22875 (N_22875,N_22258,N_22368);
and U22876 (N_22876,N_22711,N_22344);
and U22877 (N_22877,N_22356,N_22626);
nor U22878 (N_22878,N_22444,N_22601);
nand U22879 (N_22879,N_22593,N_22347);
nand U22880 (N_22880,N_22774,N_22795);
nor U22881 (N_22881,N_22694,N_22420);
nand U22882 (N_22882,N_22285,N_22525);
nor U22883 (N_22883,N_22738,N_22740);
nand U22884 (N_22884,N_22300,N_22218);
nand U22885 (N_22885,N_22527,N_22440);
or U22886 (N_22886,N_22393,N_22668);
xnor U22887 (N_22887,N_22396,N_22243);
nor U22888 (N_22888,N_22642,N_22316);
and U22889 (N_22889,N_22696,N_22464);
or U22890 (N_22890,N_22346,N_22568);
xnor U22891 (N_22891,N_22592,N_22382);
or U22892 (N_22892,N_22327,N_22490);
nand U22893 (N_22893,N_22333,N_22299);
or U22894 (N_22894,N_22489,N_22651);
or U22895 (N_22895,N_22234,N_22384);
and U22896 (N_22896,N_22747,N_22714);
and U22897 (N_22897,N_22534,N_22229);
and U22898 (N_22898,N_22349,N_22250);
xnor U22899 (N_22899,N_22706,N_22427);
and U22900 (N_22900,N_22787,N_22485);
nor U22901 (N_22901,N_22541,N_22459);
xnor U22902 (N_22902,N_22257,N_22329);
nand U22903 (N_22903,N_22672,N_22304);
nand U22904 (N_22904,N_22454,N_22719);
nor U22905 (N_22905,N_22465,N_22766);
nor U22906 (N_22906,N_22430,N_22212);
nor U22907 (N_22907,N_22594,N_22543);
nor U22908 (N_22908,N_22754,N_22544);
or U22909 (N_22909,N_22207,N_22611);
xor U22910 (N_22910,N_22551,N_22652);
and U22911 (N_22911,N_22301,N_22627);
or U22912 (N_22912,N_22704,N_22742);
nand U22913 (N_22913,N_22664,N_22540);
xor U22914 (N_22914,N_22596,N_22453);
and U22915 (N_22915,N_22578,N_22330);
nor U22916 (N_22916,N_22220,N_22703);
nand U22917 (N_22917,N_22381,N_22311);
nand U22918 (N_22918,N_22720,N_22488);
nand U22919 (N_22919,N_22203,N_22336);
nor U22920 (N_22920,N_22210,N_22361);
xor U22921 (N_22921,N_22403,N_22326);
nand U22922 (N_22922,N_22590,N_22586);
nor U22923 (N_22923,N_22518,N_22289);
or U22924 (N_22924,N_22314,N_22734);
or U22925 (N_22925,N_22282,N_22791);
nand U22926 (N_22926,N_22709,N_22648);
nor U22927 (N_22927,N_22530,N_22645);
xor U22928 (N_22928,N_22717,N_22446);
or U22929 (N_22929,N_22600,N_22661);
nand U22930 (N_22930,N_22755,N_22437);
nand U22931 (N_22931,N_22484,N_22723);
nand U22932 (N_22932,N_22639,N_22570);
nand U22933 (N_22933,N_22268,N_22211);
nor U22934 (N_22934,N_22267,N_22576);
nor U22935 (N_22935,N_22319,N_22448);
nor U22936 (N_22936,N_22575,N_22275);
or U22937 (N_22937,N_22726,N_22483);
nor U22938 (N_22938,N_22201,N_22659);
nand U22939 (N_22939,N_22773,N_22497);
and U22940 (N_22940,N_22309,N_22689);
xor U22941 (N_22941,N_22438,N_22219);
or U22942 (N_22942,N_22582,N_22524);
and U22943 (N_22943,N_22398,N_22725);
xnor U22944 (N_22944,N_22479,N_22574);
or U22945 (N_22945,N_22529,N_22699);
xor U22946 (N_22946,N_22665,N_22371);
nor U22947 (N_22947,N_22768,N_22502);
nand U22948 (N_22948,N_22345,N_22388);
or U22949 (N_22949,N_22650,N_22646);
and U22950 (N_22950,N_22365,N_22292);
or U22951 (N_22951,N_22577,N_22442);
nor U22952 (N_22952,N_22376,N_22230);
or U22953 (N_22953,N_22682,N_22431);
or U22954 (N_22954,N_22225,N_22516);
xnor U22955 (N_22955,N_22325,N_22493);
nor U22956 (N_22956,N_22503,N_22213);
and U22957 (N_22957,N_22591,N_22291);
nor U22958 (N_22958,N_22775,N_22697);
nor U22959 (N_22959,N_22798,N_22663);
and U22960 (N_22960,N_22735,N_22750);
xnor U22961 (N_22961,N_22264,N_22716);
nand U22962 (N_22962,N_22731,N_22414);
or U22963 (N_22963,N_22495,N_22788);
nand U22964 (N_22964,N_22475,N_22451);
and U22965 (N_22965,N_22227,N_22687);
or U22966 (N_22966,N_22290,N_22238);
xnor U22967 (N_22967,N_22334,N_22460);
nor U22968 (N_22968,N_22449,N_22472);
and U22969 (N_22969,N_22635,N_22439);
or U22970 (N_22970,N_22539,N_22394);
xor U22971 (N_22971,N_22538,N_22331);
and U22972 (N_22972,N_22339,N_22482);
xnor U22973 (N_22973,N_22204,N_22528);
and U22974 (N_22974,N_22217,N_22287);
xnor U22975 (N_22975,N_22589,N_22613);
or U22976 (N_22976,N_22321,N_22739);
nand U22977 (N_22977,N_22718,N_22721);
or U22978 (N_22978,N_22441,N_22748);
xor U22979 (N_22979,N_22760,N_22364);
nand U22980 (N_22980,N_22793,N_22473);
nor U22981 (N_22981,N_22749,N_22552);
or U22982 (N_22982,N_22224,N_22683);
nand U22983 (N_22983,N_22781,N_22677);
nand U22984 (N_22984,N_22547,N_22667);
nor U22985 (N_22985,N_22567,N_22236);
nand U22986 (N_22986,N_22432,N_22566);
xor U22987 (N_22987,N_22359,N_22656);
nor U22988 (N_22988,N_22205,N_22390);
nor U22989 (N_22989,N_22455,N_22408);
xnor U22990 (N_22990,N_22315,N_22644);
and U22991 (N_22991,N_22572,N_22550);
and U22992 (N_22992,N_22305,N_22603);
xor U22993 (N_22993,N_22216,N_22523);
and U22994 (N_22994,N_22280,N_22532);
nand U22995 (N_22995,N_22266,N_22310);
or U22996 (N_22996,N_22244,N_22779);
or U22997 (N_22997,N_22728,N_22654);
nand U22998 (N_22998,N_22752,N_22684);
nor U22999 (N_22999,N_22743,N_22265);
or U23000 (N_23000,N_22662,N_22500);
nand U23001 (N_23001,N_22466,N_22680);
or U23002 (N_23002,N_22686,N_22501);
nand U23003 (N_23003,N_22617,N_22607);
or U23004 (N_23004,N_22701,N_22324);
nand U23005 (N_23005,N_22563,N_22232);
nor U23006 (N_23006,N_22597,N_22433);
xnor U23007 (N_23007,N_22254,N_22271);
nor U23008 (N_23008,N_22556,N_22504);
xnor U23009 (N_23009,N_22666,N_22710);
xor U23010 (N_23010,N_22751,N_22429);
or U23011 (N_23011,N_22564,N_22623);
nor U23012 (N_23012,N_22625,N_22519);
nor U23013 (N_23013,N_22581,N_22571);
or U23014 (N_23014,N_22215,N_22618);
xor U23015 (N_23015,N_22730,N_22557);
nand U23016 (N_23016,N_22352,N_22757);
and U23017 (N_23017,N_22741,N_22660);
nand U23018 (N_23018,N_22348,N_22383);
or U23019 (N_23019,N_22237,N_22643);
xor U23020 (N_23020,N_22377,N_22756);
xnor U23021 (N_23021,N_22565,N_22610);
nor U23022 (N_23022,N_22771,N_22256);
nand U23023 (N_23023,N_22792,N_22354);
xnor U23024 (N_23024,N_22554,N_22417);
or U23025 (N_23025,N_22387,N_22558);
and U23026 (N_23026,N_22640,N_22369);
xnor U23027 (N_23027,N_22521,N_22281);
nor U23028 (N_23028,N_22262,N_22318);
nand U23029 (N_23029,N_22794,N_22702);
xnor U23030 (N_23030,N_22612,N_22248);
nand U23031 (N_23031,N_22507,N_22413);
xor U23032 (N_23032,N_22655,N_22456);
or U23033 (N_23033,N_22355,N_22657);
and U23034 (N_23034,N_22675,N_22263);
nand U23035 (N_23035,N_22269,N_22270);
nand U23036 (N_23036,N_22535,N_22555);
and U23037 (N_23037,N_22457,N_22517);
xnor U23038 (N_23038,N_22411,N_22259);
nand U23039 (N_23039,N_22208,N_22477);
nand U23040 (N_23040,N_22511,N_22685);
nor U23041 (N_23041,N_22428,N_22537);
nand U23042 (N_23042,N_22425,N_22729);
and U23043 (N_23043,N_22695,N_22678);
nor U23044 (N_23044,N_22405,N_22491);
and U23045 (N_23045,N_22622,N_22605);
and U23046 (N_23046,N_22323,N_22406);
nor U23047 (N_23047,N_22494,N_22233);
nand U23048 (N_23048,N_22467,N_22688);
or U23049 (N_23049,N_22636,N_22276);
nor U23050 (N_23050,N_22736,N_22674);
xor U23051 (N_23051,N_22274,N_22602);
or U23052 (N_23052,N_22468,N_22588);
nand U23053 (N_23053,N_22587,N_22505);
or U23054 (N_23054,N_22692,N_22404);
and U23055 (N_23055,N_22375,N_22200);
xnor U23056 (N_23056,N_22317,N_22343);
and U23057 (N_23057,N_22392,N_22732);
xnor U23058 (N_23058,N_22670,N_22421);
xnor U23059 (N_23059,N_22559,N_22260);
xor U23060 (N_23060,N_22391,N_22770);
and U23061 (N_23061,N_22658,N_22520);
xnor U23062 (N_23062,N_22673,N_22514);
nand U23063 (N_23063,N_22313,N_22579);
nor U23064 (N_23064,N_22630,N_22797);
nand U23065 (N_23065,N_22585,N_22737);
or U23066 (N_23066,N_22776,N_22379);
nand U23067 (N_23067,N_22471,N_22435);
xor U23068 (N_23068,N_22373,N_22303);
xnor U23069 (N_23069,N_22286,N_22599);
and U23070 (N_23070,N_22705,N_22450);
nand U23071 (N_23071,N_22447,N_22536);
nand U23072 (N_23072,N_22360,N_22284);
and U23073 (N_23073,N_22510,N_22202);
nand U23074 (N_23074,N_22240,N_22231);
nand U23075 (N_23075,N_22366,N_22583);
xnor U23076 (N_23076,N_22727,N_22698);
and U23077 (N_23077,N_22700,N_22619);
or U23078 (N_23078,N_22492,N_22426);
xor U23079 (N_23079,N_22691,N_22423);
and U23080 (N_23080,N_22351,N_22374);
xnor U23081 (N_23081,N_22783,N_22399);
nand U23082 (N_23082,N_22335,N_22631);
xor U23083 (N_23083,N_22522,N_22255);
and U23084 (N_23084,N_22370,N_22713);
and U23085 (N_23085,N_22759,N_22461);
nand U23086 (N_23086,N_22273,N_22614);
and U23087 (N_23087,N_22533,N_22606);
xnor U23088 (N_23088,N_22239,N_22341);
and U23089 (N_23089,N_22512,N_22214);
or U23090 (N_23090,N_22561,N_22419);
nand U23091 (N_23091,N_22784,N_22206);
and U23092 (N_23092,N_22293,N_22789);
and U23093 (N_23093,N_22372,N_22778);
nand U23094 (N_23094,N_22253,N_22312);
or U23095 (N_23095,N_22350,N_22598);
nand U23096 (N_23096,N_22297,N_22763);
xnor U23097 (N_23097,N_22638,N_22620);
and U23098 (N_23098,N_22498,N_22478);
or U23099 (N_23099,N_22707,N_22337);
and U23100 (N_23100,N_22282,N_22632);
or U23101 (N_23101,N_22410,N_22758);
and U23102 (N_23102,N_22515,N_22407);
xnor U23103 (N_23103,N_22306,N_22790);
or U23104 (N_23104,N_22435,N_22714);
nor U23105 (N_23105,N_22299,N_22284);
and U23106 (N_23106,N_22512,N_22798);
and U23107 (N_23107,N_22385,N_22586);
xnor U23108 (N_23108,N_22285,N_22517);
or U23109 (N_23109,N_22722,N_22703);
nor U23110 (N_23110,N_22502,N_22345);
or U23111 (N_23111,N_22680,N_22229);
xnor U23112 (N_23112,N_22736,N_22276);
or U23113 (N_23113,N_22683,N_22350);
or U23114 (N_23114,N_22405,N_22641);
and U23115 (N_23115,N_22320,N_22601);
and U23116 (N_23116,N_22323,N_22336);
nor U23117 (N_23117,N_22567,N_22425);
nand U23118 (N_23118,N_22474,N_22379);
nand U23119 (N_23119,N_22328,N_22255);
and U23120 (N_23120,N_22788,N_22781);
nand U23121 (N_23121,N_22492,N_22799);
and U23122 (N_23122,N_22316,N_22632);
nand U23123 (N_23123,N_22686,N_22447);
and U23124 (N_23124,N_22271,N_22794);
nor U23125 (N_23125,N_22386,N_22480);
xnor U23126 (N_23126,N_22335,N_22617);
or U23127 (N_23127,N_22736,N_22364);
nor U23128 (N_23128,N_22265,N_22674);
xnor U23129 (N_23129,N_22248,N_22753);
nand U23130 (N_23130,N_22680,N_22598);
or U23131 (N_23131,N_22398,N_22393);
or U23132 (N_23132,N_22309,N_22225);
or U23133 (N_23133,N_22564,N_22335);
and U23134 (N_23134,N_22588,N_22585);
and U23135 (N_23135,N_22405,N_22544);
and U23136 (N_23136,N_22574,N_22355);
nand U23137 (N_23137,N_22732,N_22782);
nand U23138 (N_23138,N_22521,N_22374);
xnor U23139 (N_23139,N_22705,N_22531);
xor U23140 (N_23140,N_22663,N_22749);
nand U23141 (N_23141,N_22770,N_22787);
nand U23142 (N_23142,N_22242,N_22302);
nor U23143 (N_23143,N_22731,N_22697);
or U23144 (N_23144,N_22758,N_22767);
nand U23145 (N_23145,N_22693,N_22261);
nand U23146 (N_23146,N_22390,N_22742);
and U23147 (N_23147,N_22726,N_22241);
nand U23148 (N_23148,N_22511,N_22480);
or U23149 (N_23149,N_22490,N_22379);
nand U23150 (N_23150,N_22248,N_22628);
or U23151 (N_23151,N_22452,N_22783);
nand U23152 (N_23152,N_22374,N_22347);
and U23153 (N_23153,N_22626,N_22224);
nand U23154 (N_23154,N_22438,N_22762);
or U23155 (N_23155,N_22210,N_22341);
nand U23156 (N_23156,N_22213,N_22692);
and U23157 (N_23157,N_22723,N_22394);
nor U23158 (N_23158,N_22268,N_22212);
or U23159 (N_23159,N_22245,N_22788);
xor U23160 (N_23160,N_22510,N_22361);
and U23161 (N_23161,N_22292,N_22203);
nor U23162 (N_23162,N_22741,N_22269);
and U23163 (N_23163,N_22623,N_22541);
and U23164 (N_23164,N_22275,N_22629);
xnor U23165 (N_23165,N_22363,N_22585);
xnor U23166 (N_23166,N_22640,N_22606);
xor U23167 (N_23167,N_22225,N_22315);
nor U23168 (N_23168,N_22551,N_22614);
and U23169 (N_23169,N_22770,N_22340);
and U23170 (N_23170,N_22287,N_22798);
nor U23171 (N_23171,N_22672,N_22500);
nor U23172 (N_23172,N_22738,N_22519);
or U23173 (N_23173,N_22583,N_22409);
and U23174 (N_23174,N_22569,N_22412);
nor U23175 (N_23175,N_22436,N_22778);
nor U23176 (N_23176,N_22258,N_22631);
or U23177 (N_23177,N_22645,N_22424);
xor U23178 (N_23178,N_22366,N_22762);
xor U23179 (N_23179,N_22266,N_22574);
or U23180 (N_23180,N_22346,N_22766);
nand U23181 (N_23181,N_22679,N_22481);
xnor U23182 (N_23182,N_22350,N_22346);
nor U23183 (N_23183,N_22665,N_22254);
xor U23184 (N_23184,N_22480,N_22732);
nor U23185 (N_23185,N_22205,N_22652);
and U23186 (N_23186,N_22778,N_22441);
nor U23187 (N_23187,N_22331,N_22772);
xnor U23188 (N_23188,N_22649,N_22690);
nand U23189 (N_23189,N_22362,N_22744);
and U23190 (N_23190,N_22226,N_22718);
nor U23191 (N_23191,N_22349,N_22516);
nor U23192 (N_23192,N_22253,N_22266);
and U23193 (N_23193,N_22330,N_22411);
or U23194 (N_23194,N_22522,N_22631);
nand U23195 (N_23195,N_22504,N_22414);
nor U23196 (N_23196,N_22724,N_22283);
or U23197 (N_23197,N_22740,N_22543);
and U23198 (N_23198,N_22384,N_22203);
nand U23199 (N_23199,N_22671,N_22612);
nand U23200 (N_23200,N_22340,N_22207);
xor U23201 (N_23201,N_22347,N_22362);
xor U23202 (N_23202,N_22671,N_22267);
or U23203 (N_23203,N_22772,N_22457);
xor U23204 (N_23204,N_22584,N_22459);
and U23205 (N_23205,N_22509,N_22618);
nor U23206 (N_23206,N_22335,N_22346);
or U23207 (N_23207,N_22513,N_22319);
nor U23208 (N_23208,N_22739,N_22650);
xor U23209 (N_23209,N_22731,N_22448);
nor U23210 (N_23210,N_22624,N_22289);
and U23211 (N_23211,N_22464,N_22234);
or U23212 (N_23212,N_22234,N_22460);
nor U23213 (N_23213,N_22761,N_22579);
nand U23214 (N_23214,N_22577,N_22607);
xor U23215 (N_23215,N_22453,N_22661);
nor U23216 (N_23216,N_22416,N_22263);
and U23217 (N_23217,N_22716,N_22548);
nor U23218 (N_23218,N_22328,N_22573);
nor U23219 (N_23219,N_22629,N_22363);
nor U23220 (N_23220,N_22669,N_22672);
nor U23221 (N_23221,N_22539,N_22321);
nor U23222 (N_23222,N_22348,N_22664);
nand U23223 (N_23223,N_22266,N_22763);
nand U23224 (N_23224,N_22207,N_22683);
or U23225 (N_23225,N_22538,N_22675);
nor U23226 (N_23226,N_22419,N_22650);
xnor U23227 (N_23227,N_22444,N_22284);
nand U23228 (N_23228,N_22201,N_22522);
and U23229 (N_23229,N_22222,N_22462);
nor U23230 (N_23230,N_22251,N_22582);
nand U23231 (N_23231,N_22623,N_22659);
nand U23232 (N_23232,N_22256,N_22606);
nor U23233 (N_23233,N_22455,N_22606);
and U23234 (N_23234,N_22724,N_22713);
and U23235 (N_23235,N_22227,N_22303);
xor U23236 (N_23236,N_22426,N_22306);
xor U23237 (N_23237,N_22473,N_22667);
or U23238 (N_23238,N_22436,N_22288);
and U23239 (N_23239,N_22269,N_22214);
xor U23240 (N_23240,N_22692,N_22425);
and U23241 (N_23241,N_22338,N_22318);
or U23242 (N_23242,N_22275,N_22485);
xnor U23243 (N_23243,N_22771,N_22297);
or U23244 (N_23244,N_22639,N_22295);
nor U23245 (N_23245,N_22520,N_22276);
or U23246 (N_23246,N_22265,N_22518);
nand U23247 (N_23247,N_22201,N_22251);
nand U23248 (N_23248,N_22747,N_22649);
and U23249 (N_23249,N_22594,N_22637);
and U23250 (N_23250,N_22244,N_22733);
xnor U23251 (N_23251,N_22729,N_22726);
nor U23252 (N_23252,N_22345,N_22649);
nand U23253 (N_23253,N_22330,N_22389);
xor U23254 (N_23254,N_22336,N_22319);
xor U23255 (N_23255,N_22523,N_22635);
and U23256 (N_23256,N_22320,N_22360);
and U23257 (N_23257,N_22247,N_22701);
and U23258 (N_23258,N_22672,N_22718);
or U23259 (N_23259,N_22788,N_22338);
and U23260 (N_23260,N_22687,N_22220);
or U23261 (N_23261,N_22468,N_22476);
or U23262 (N_23262,N_22685,N_22778);
and U23263 (N_23263,N_22719,N_22308);
or U23264 (N_23264,N_22496,N_22696);
and U23265 (N_23265,N_22252,N_22676);
xnor U23266 (N_23266,N_22528,N_22464);
or U23267 (N_23267,N_22504,N_22459);
nor U23268 (N_23268,N_22694,N_22275);
or U23269 (N_23269,N_22498,N_22439);
and U23270 (N_23270,N_22491,N_22271);
nand U23271 (N_23271,N_22779,N_22462);
nor U23272 (N_23272,N_22739,N_22745);
nand U23273 (N_23273,N_22324,N_22202);
nand U23274 (N_23274,N_22483,N_22440);
nand U23275 (N_23275,N_22450,N_22392);
nand U23276 (N_23276,N_22537,N_22758);
or U23277 (N_23277,N_22410,N_22699);
and U23278 (N_23278,N_22425,N_22549);
or U23279 (N_23279,N_22793,N_22273);
xor U23280 (N_23280,N_22535,N_22407);
nand U23281 (N_23281,N_22304,N_22443);
xor U23282 (N_23282,N_22200,N_22653);
nand U23283 (N_23283,N_22212,N_22281);
or U23284 (N_23284,N_22390,N_22372);
or U23285 (N_23285,N_22492,N_22644);
nor U23286 (N_23286,N_22550,N_22280);
xnor U23287 (N_23287,N_22573,N_22302);
and U23288 (N_23288,N_22379,N_22551);
nand U23289 (N_23289,N_22755,N_22244);
xor U23290 (N_23290,N_22544,N_22680);
or U23291 (N_23291,N_22785,N_22560);
nor U23292 (N_23292,N_22228,N_22404);
nor U23293 (N_23293,N_22427,N_22790);
nor U23294 (N_23294,N_22686,N_22482);
nand U23295 (N_23295,N_22350,N_22747);
and U23296 (N_23296,N_22449,N_22784);
and U23297 (N_23297,N_22309,N_22442);
nor U23298 (N_23298,N_22516,N_22357);
or U23299 (N_23299,N_22312,N_22412);
or U23300 (N_23300,N_22391,N_22269);
or U23301 (N_23301,N_22412,N_22590);
nand U23302 (N_23302,N_22409,N_22268);
or U23303 (N_23303,N_22455,N_22503);
or U23304 (N_23304,N_22535,N_22306);
or U23305 (N_23305,N_22652,N_22680);
xor U23306 (N_23306,N_22588,N_22318);
nand U23307 (N_23307,N_22616,N_22216);
nand U23308 (N_23308,N_22455,N_22483);
nor U23309 (N_23309,N_22759,N_22230);
xor U23310 (N_23310,N_22346,N_22204);
xnor U23311 (N_23311,N_22733,N_22650);
and U23312 (N_23312,N_22356,N_22448);
nor U23313 (N_23313,N_22414,N_22445);
or U23314 (N_23314,N_22418,N_22590);
and U23315 (N_23315,N_22387,N_22308);
nor U23316 (N_23316,N_22786,N_22403);
or U23317 (N_23317,N_22595,N_22652);
nor U23318 (N_23318,N_22629,N_22396);
or U23319 (N_23319,N_22378,N_22230);
or U23320 (N_23320,N_22312,N_22564);
xnor U23321 (N_23321,N_22318,N_22668);
or U23322 (N_23322,N_22579,N_22715);
nand U23323 (N_23323,N_22545,N_22601);
xor U23324 (N_23324,N_22241,N_22606);
nand U23325 (N_23325,N_22322,N_22733);
xnor U23326 (N_23326,N_22704,N_22275);
xor U23327 (N_23327,N_22386,N_22242);
and U23328 (N_23328,N_22387,N_22351);
nor U23329 (N_23329,N_22784,N_22594);
xor U23330 (N_23330,N_22669,N_22719);
nor U23331 (N_23331,N_22656,N_22251);
or U23332 (N_23332,N_22315,N_22304);
or U23333 (N_23333,N_22758,N_22527);
nor U23334 (N_23334,N_22492,N_22402);
nor U23335 (N_23335,N_22616,N_22458);
or U23336 (N_23336,N_22244,N_22690);
nor U23337 (N_23337,N_22637,N_22267);
nand U23338 (N_23338,N_22286,N_22716);
xnor U23339 (N_23339,N_22711,N_22721);
nor U23340 (N_23340,N_22306,N_22352);
nand U23341 (N_23341,N_22529,N_22298);
xor U23342 (N_23342,N_22256,N_22324);
nand U23343 (N_23343,N_22367,N_22498);
nor U23344 (N_23344,N_22548,N_22502);
xor U23345 (N_23345,N_22669,N_22627);
nor U23346 (N_23346,N_22724,N_22256);
nand U23347 (N_23347,N_22519,N_22413);
nor U23348 (N_23348,N_22333,N_22276);
nand U23349 (N_23349,N_22488,N_22621);
and U23350 (N_23350,N_22358,N_22222);
or U23351 (N_23351,N_22554,N_22522);
and U23352 (N_23352,N_22420,N_22283);
xnor U23353 (N_23353,N_22265,N_22207);
and U23354 (N_23354,N_22566,N_22519);
xnor U23355 (N_23355,N_22390,N_22233);
and U23356 (N_23356,N_22430,N_22521);
xnor U23357 (N_23357,N_22770,N_22630);
and U23358 (N_23358,N_22610,N_22644);
nand U23359 (N_23359,N_22581,N_22444);
nand U23360 (N_23360,N_22220,N_22295);
nand U23361 (N_23361,N_22405,N_22682);
nand U23362 (N_23362,N_22247,N_22617);
xor U23363 (N_23363,N_22241,N_22383);
nand U23364 (N_23364,N_22588,N_22553);
xor U23365 (N_23365,N_22550,N_22478);
and U23366 (N_23366,N_22533,N_22333);
or U23367 (N_23367,N_22708,N_22461);
or U23368 (N_23368,N_22513,N_22734);
nand U23369 (N_23369,N_22370,N_22431);
nor U23370 (N_23370,N_22232,N_22528);
nand U23371 (N_23371,N_22459,N_22727);
nor U23372 (N_23372,N_22777,N_22601);
nand U23373 (N_23373,N_22209,N_22577);
nor U23374 (N_23374,N_22650,N_22277);
nand U23375 (N_23375,N_22586,N_22458);
nor U23376 (N_23376,N_22327,N_22733);
nand U23377 (N_23377,N_22687,N_22360);
nand U23378 (N_23378,N_22432,N_22474);
and U23379 (N_23379,N_22301,N_22349);
and U23380 (N_23380,N_22273,N_22291);
and U23381 (N_23381,N_22720,N_22338);
xor U23382 (N_23382,N_22407,N_22409);
and U23383 (N_23383,N_22362,N_22205);
nor U23384 (N_23384,N_22480,N_22462);
and U23385 (N_23385,N_22604,N_22636);
or U23386 (N_23386,N_22341,N_22255);
nor U23387 (N_23387,N_22602,N_22754);
or U23388 (N_23388,N_22565,N_22209);
and U23389 (N_23389,N_22259,N_22352);
nor U23390 (N_23390,N_22257,N_22622);
nor U23391 (N_23391,N_22366,N_22632);
xnor U23392 (N_23392,N_22670,N_22611);
or U23393 (N_23393,N_22348,N_22576);
or U23394 (N_23394,N_22219,N_22779);
nor U23395 (N_23395,N_22438,N_22573);
xor U23396 (N_23396,N_22653,N_22400);
nand U23397 (N_23397,N_22719,N_22721);
nand U23398 (N_23398,N_22611,N_22386);
nor U23399 (N_23399,N_22427,N_22390);
xnor U23400 (N_23400,N_23171,N_23352);
or U23401 (N_23401,N_23027,N_23244);
or U23402 (N_23402,N_22949,N_22822);
or U23403 (N_23403,N_22928,N_23219);
nand U23404 (N_23404,N_23231,N_23012);
or U23405 (N_23405,N_23025,N_23347);
nand U23406 (N_23406,N_23216,N_23143);
and U23407 (N_23407,N_22923,N_23030);
nor U23408 (N_23408,N_23134,N_23001);
xor U23409 (N_23409,N_23234,N_22953);
nand U23410 (N_23410,N_22944,N_23304);
and U23411 (N_23411,N_23239,N_23059);
or U23412 (N_23412,N_23049,N_23034);
nand U23413 (N_23413,N_22937,N_23100);
nor U23414 (N_23414,N_22968,N_23033);
xnor U23415 (N_23415,N_22935,N_23380);
nand U23416 (N_23416,N_23179,N_23266);
nor U23417 (N_23417,N_22877,N_23357);
nor U23418 (N_23418,N_23312,N_23305);
nand U23419 (N_23419,N_22894,N_22800);
nor U23420 (N_23420,N_23285,N_23036);
and U23421 (N_23421,N_23140,N_22857);
nand U23422 (N_23422,N_23210,N_23293);
nand U23423 (N_23423,N_22985,N_23350);
xnor U23424 (N_23424,N_23105,N_23342);
and U23425 (N_23425,N_23302,N_23270);
xor U23426 (N_23426,N_22890,N_22999);
nor U23427 (N_23427,N_22836,N_23102);
or U23428 (N_23428,N_22841,N_22812);
xor U23429 (N_23429,N_23117,N_23050);
and U23430 (N_23430,N_23386,N_23055);
xor U23431 (N_23431,N_22811,N_23323);
and U23432 (N_23432,N_23104,N_23024);
and U23433 (N_23433,N_23045,N_22843);
and U23434 (N_23434,N_23156,N_23046);
xor U23435 (N_23435,N_22964,N_23068);
and U23436 (N_23436,N_23113,N_22952);
and U23437 (N_23437,N_22895,N_23004);
nand U23438 (N_23438,N_23295,N_23203);
xor U23439 (N_23439,N_23209,N_23009);
xnor U23440 (N_23440,N_23311,N_23136);
and U23441 (N_23441,N_23262,N_22902);
nand U23442 (N_23442,N_23016,N_23353);
nand U23443 (N_23443,N_23044,N_23280);
xnor U23444 (N_23444,N_22929,N_23324);
and U23445 (N_23445,N_23196,N_22927);
and U23446 (N_23446,N_23251,N_22962);
and U23447 (N_23447,N_23273,N_22912);
nand U23448 (N_23448,N_23056,N_23088);
nor U23449 (N_23449,N_22819,N_22904);
nor U23450 (N_23450,N_22974,N_22861);
xnor U23451 (N_23451,N_23072,N_22809);
or U23452 (N_23452,N_22879,N_23213);
xnor U23453 (N_23453,N_22860,N_23131);
and U23454 (N_23454,N_23083,N_23002);
and U23455 (N_23455,N_22804,N_22853);
xnor U23456 (N_23456,N_23278,N_23167);
and U23457 (N_23457,N_23346,N_22901);
nand U23458 (N_23458,N_23189,N_22854);
nor U23459 (N_23459,N_23249,N_23343);
nand U23460 (N_23460,N_23335,N_23398);
nor U23461 (N_23461,N_23162,N_22963);
xor U23462 (N_23462,N_23397,N_22858);
nor U23463 (N_23463,N_22940,N_23381);
nor U23464 (N_23464,N_23076,N_22961);
xor U23465 (N_23465,N_23388,N_23145);
or U23466 (N_23466,N_23023,N_23298);
or U23467 (N_23467,N_22889,N_22862);
or U23468 (N_23468,N_22820,N_23374);
nor U23469 (N_23469,N_23057,N_23396);
nor U23470 (N_23470,N_23301,N_23325);
and U23471 (N_23471,N_22917,N_23132);
nor U23472 (N_23472,N_22826,N_23263);
or U23473 (N_23473,N_22876,N_22914);
nand U23474 (N_23474,N_23190,N_23297);
and U23475 (N_23475,N_23256,N_23199);
and U23476 (N_23476,N_22838,N_23067);
nand U23477 (N_23477,N_23037,N_23365);
nor U23478 (N_23478,N_22806,N_22840);
nor U23479 (N_23479,N_23317,N_23092);
nand U23480 (N_23480,N_23390,N_22971);
and U23481 (N_23481,N_22907,N_23385);
nand U23482 (N_23482,N_22808,N_22849);
and U23483 (N_23483,N_23032,N_23071);
and U23484 (N_23484,N_23279,N_23316);
and U23485 (N_23485,N_23207,N_22810);
or U23486 (N_23486,N_23334,N_23308);
nand U23487 (N_23487,N_23159,N_23269);
and U23488 (N_23488,N_22918,N_22863);
xor U23489 (N_23489,N_23178,N_23303);
and U23490 (N_23490,N_23310,N_23114);
or U23491 (N_23491,N_23369,N_23064);
or U23492 (N_23492,N_23202,N_23022);
or U23493 (N_23493,N_23370,N_22855);
xnor U23494 (N_23494,N_23363,N_23326);
nand U23495 (N_23495,N_23031,N_23255);
nor U23496 (N_23496,N_23361,N_23395);
or U23497 (N_23497,N_22994,N_23226);
nand U23498 (N_23498,N_23364,N_23052);
nand U23499 (N_23499,N_23081,N_23164);
nor U23500 (N_23500,N_22969,N_23250);
or U23501 (N_23501,N_22977,N_23082);
xnor U23502 (N_23502,N_22903,N_23201);
nor U23503 (N_23503,N_22831,N_22837);
nor U23504 (N_23504,N_23391,N_22955);
nor U23505 (N_23505,N_23314,N_22815);
or U23506 (N_23506,N_23135,N_23260);
nor U23507 (N_23507,N_23166,N_23247);
nand U23508 (N_23508,N_23393,N_22991);
xnor U23509 (N_23509,N_22960,N_22818);
and U23510 (N_23510,N_23130,N_23264);
nor U23511 (N_23511,N_23122,N_23101);
and U23512 (N_23512,N_22970,N_22941);
or U23513 (N_23513,N_23149,N_22998);
and U23514 (N_23514,N_23174,N_22930);
nor U23515 (N_23515,N_23133,N_23095);
nor U23516 (N_23516,N_22984,N_23351);
xor U23517 (N_23517,N_22906,N_22922);
xnor U23518 (N_23518,N_22992,N_23268);
nand U23519 (N_23519,N_22946,N_23319);
or U23520 (N_23520,N_22884,N_23309);
nand U23521 (N_23521,N_23080,N_22911);
and U23522 (N_23522,N_22891,N_22945);
nor U23523 (N_23523,N_23169,N_23233);
nand U23524 (N_23524,N_22867,N_23187);
nor U23525 (N_23525,N_23139,N_23220);
nand U23526 (N_23526,N_22919,N_22823);
and U23527 (N_23527,N_23123,N_23377);
or U23528 (N_23528,N_23315,N_23204);
and U23529 (N_23529,N_23253,N_23153);
nand U23530 (N_23530,N_23090,N_23359);
and U23531 (N_23531,N_23007,N_23089);
nor U23532 (N_23532,N_23106,N_23194);
nand U23533 (N_23533,N_22878,N_23107);
nor U23534 (N_23534,N_23079,N_22896);
nand U23535 (N_23535,N_23154,N_23112);
nor U23536 (N_23536,N_23110,N_23281);
and U23537 (N_23537,N_23307,N_23096);
xnor U23538 (N_23538,N_22830,N_22886);
xor U23539 (N_23539,N_22954,N_22926);
or U23540 (N_23540,N_23138,N_22873);
nor U23541 (N_23541,N_23184,N_23177);
or U23542 (N_23542,N_23318,N_23185);
xor U23543 (N_23543,N_23217,N_23331);
nor U23544 (N_23544,N_23000,N_22980);
nor U23545 (N_23545,N_23294,N_22909);
nor U23546 (N_23546,N_23108,N_22990);
or U23547 (N_23547,N_22978,N_23376);
nor U23548 (N_23548,N_23077,N_23116);
xnor U23549 (N_23549,N_23332,N_23274);
xor U23550 (N_23550,N_23075,N_23005);
or U23551 (N_23551,N_23236,N_22859);
nand U23552 (N_23552,N_23243,N_22829);
nand U23553 (N_23553,N_23257,N_22936);
or U23554 (N_23554,N_22865,N_23214);
xnor U23555 (N_23555,N_22915,N_23337);
nand U23556 (N_23556,N_22844,N_23040);
or U23557 (N_23557,N_22932,N_23222);
nand U23558 (N_23558,N_22973,N_22824);
or U23559 (N_23559,N_23086,N_22847);
or U23560 (N_23560,N_23259,N_23211);
xor U23561 (N_23561,N_23235,N_23028);
nand U23562 (N_23562,N_23212,N_23065);
xnor U23563 (N_23563,N_23392,N_23091);
nand U23564 (N_23564,N_23223,N_22835);
xnor U23565 (N_23565,N_22864,N_23356);
xnor U23566 (N_23566,N_23277,N_23158);
xnor U23567 (N_23567,N_23058,N_23144);
or U23568 (N_23568,N_22979,N_22875);
xor U23569 (N_23569,N_22976,N_22816);
nand U23570 (N_23570,N_23328,N_23163);
nand U23571 (N_23571,N_23017,N_22933);
xnor U23572 (N_23572,N_23284,N_22845);
and U23573 (N_23573,N_23366,N_23373);
or U23574 (N_23574,N_23029,N_23271);
nand U23575 (N_23575,N_22869,N_23120);
nand U23576 (N_23576,N_23013,N_23188);
nor U23577 (N_23577,N_22996,N_23286);
nor U23578 (N_23578,N_23399,N_23349);
nor U23579 (N_23579,N_23043,N_23230);
xor U23580 (N_23580,N_23197,N_23125);
xnor U23581 (N_23581,N_23141,N_23109);
and U23582 (N_23582,N_23282,N_23206);
or U23583 (N_23583,N_22948,N_23047);
nor U23584 (N_23584,N_23367,N_23183);
or U23585 (N_23585,N_22870,N_23321);
or U23586 (N_23586,N_22951,N_23192);
or U23587 (N_23587,N_23290,N_23333);
nor U23588 (N_23588,N_22986,N_23176);
nor U23589 (N_23589,N_23362,N_23340);
nor U23590 (N_23590,N_22898,N_23245);
nor U23591 (N_23591,N_22967,N_23003);
nand U23592 (N_23592,N_22839,N_23011);
xnor U23593 (N_23593,N_23287,N_23119);
nand U23594 (N_23594,N_23146,N_23066);
xnor U23595 (N_23595,N_23165,N_23168);
nor U23596 (N_23596,N_22817,N_23306);
xnor U23597 (N_23597,N_23339,N_23389);
xor U23598 (N_23598,N_23205,N_23097);
nand U23599 (N_23599,N_23111,N_23085);
nand U23600 (N_23600,N_23228,N_23267);
and U23601 (N_23601,N_23008,N_23193);
and U23602 (N_23602,N_23289,N_23103);
nor U23603 (N_23603,N_23338,N_23252);
or U23604 (N_23604,N_23148,N_22943);
xor U23605 (N_23605,N_23379,N_23227);
nor U23606 (N_23606,N_23300,N_22834);
and U23607 (N_23607,N_23355,N_22874);
nor U23608 (N_23608,N_23142,N_22942);
and U23609 (N_23609,N_23387,N_22931);
xnor U23610 (N_23610,N_23010,N_23382);
and U23611 (N_23611,N_23137,N_23225);
nand U23612 (N_23612,N_23344,N_22920);
or U23613 (N_23613,N_23191,N_22805);
or U23614 (N_23614,N_23151,N_22851);
and U23615 (N_23615,N_22908,N_23313);
xor U23616 (N_23616,N_23147,N_22913);
xor U23617 (N_23617,N_22958,N_23006);
xor U23618 (N_23618,N_22885,N_23152);
and U23619 (N_23619,N_23014,N_22965);
xor U23620 (N_23620,N_23128,N_23261);
nor U23621 (N_23621,N_23232,N_23053);
xor U23622 (N_23622,N_23384,N_22868);
nor U23623 (N_23623,N_23341,N_22925);
xor U23624 (N_23624,N_22850,N_22956);
nor U23625 (N_23625,N_22957,N_23129);
or U23626 (N_23626,N_23296,N_23336);
xor U23627 (N_23627,N_23265,N_22813);
nor U23628 (N_23628,N_23394,N_23354);
and U23629 (N_23629,N_23242,N_22916);
nand U23630 (N_23630,N_23020,N_22934);
or U23631 (N_23631,N_22872,N_23299);
nor U23632 (N_23632,N_22848,N_22881);
and U23633 (N_23633,N_22892,N_23358);
or U23634 (N_23634,N_23093,N_23062);
nand U23635 (N_23635,N_23155,N_22814);
or U23636 (N_23636,N_23371,N_22825);
nor U23637 (N_23637,N_23060,N_22947);
xnor U23638 (N_23638,N_23378,N_23215);
nand U23639 (N_23639,N_23198,N_23375);
nand U23640 (N_23640,N_22972,N_22866);
or U23641 (N_23641,N_23070,N_23115);
nand U23642 (N_23642,N_22993,N_23322);
and U23643 (N_23643,N_22989,N_22921);
and U23644 (N_23644,N_22871,N_23078);
nand U23645 (N_23645,N_22924,N_23084);
xor U23646 (N_23646,N_22883,N_22888);
nor U23647 (N_23647,N_22887,N_23283);
nor U23648 (N_23648,N_22846,N_23041);
nand U23649 (N_23649,N_23195,N_23021);
or U23650 (N_23650,N_22959,N_23157);
and U23651 (N_23651,N_23348,N_23087);
and U23652 (N_23652,N_23238,N_23063);
and U23653 (N_23653,N_23237,N_22987);
nor U23654 (N_23654,N_23200,N_22802);
nand U23655 (N_23655,N_23015,N_23254);
xnor U23656 (N_23656,N_23330,N_22950);
xor U23657 (N_23657,N_23276,N_23019);
or U23658 (N_23658,N_22852,N_23170);
or U23659 (N_23659,N_23288,N_23275);
and U23660 (N_23660,N_23186,N_23069);
or U23661 (N_23661,N_23042,N_22966);
or U23662 (N_23662,N_23291,N_22981);
nor U23663 (N_23663,N_22899,N_23221);
or U23664 (N_23664,N_23182,N_22897);
xnor U23665 (N_23665,N_22938,N_23048);
or U23666 (N_23666,N_23118,N_23051);
xor U23667 (N_23667,N_22856,N_22905);
nand U23668 (N_23668,N_22827,N_22975);
nor U23669 (N_23669,N_23180,N_23208);
and U23670 (N_23670,N_23320,N_23368);
nor U23671 (N_23671,N_22939,N_22821);
and U23672 (N_23672,N_23218,N_23241);
nor U23673 (N_23673,N_23150,N_23372);
nand U23674 (N_23674,N_23248,N_23181);
or U23675 (N_23675,N_22995,N_23099);
and U23676 (N_23676,N_23074,N_23038);
or U23677 (N_23677,N_22832,N_22988);
or U23678 (N_23678,N_23172,N_23035);
nand U23679 (N_23679,N_23054,N_22807);
and U23680 (N_23680,N_22900,N_22910);
and U23681 (N_23681,N_23292,N_23121);
nand U23682 (N_23682,N_23360,N_22893);
nand U23683 (N_23683,N_23175,N_23383);
nand U23684 (N_23684,N_23127,N_23124);
or U23685 (N_23685,N_23039,N_22828);
xnor U23686 (N_23686,N_22982,N_22803);
xnor U23687 (N_23687,N_23160,N_23224);
nand U23688 (N_23688,N_23327,N_23258);
and U23689 (N_23689,N_22983,N_22833);
nand U23690 (N_23690,N_23073,N_23229);
and U23691 (N_23691,N_22882,N_23161);
nor U23692 (N_23692,N_23345,N_23173);
nor U23693 (N_23693,N_23272,N_22880);
or U23694 (N_23694,N_22801,N_23094);
xor U23695 (N_23695,N_23246,N_23126);
and U23696 (N_23696,N_23018,N_23098);
or U23697 (N_23697,N_22842,N_22997);
nand U23698 (N_23698,N_23061,N_23026);
nor U23699 (N_23699,N_23240,N_23329);
and U23700 (N_23700,N_22885,N_23115);
nand U23701 (N_23701,N_23156,N_23186);
nor U23702 (N_23702,N_23051,N_23053);
xnor U23703 (N_23703,N_22922,N_23267);
nand U23704 (N_23704,N_23341,N_23236);
xor U23705 (N_23705,N_23158,N_22852);
xor U23706 (N_23706,N_23302,N_23015);
nor U23707 (N_23707,N_22909,N_23347);
and U23708 (N_23708,N_23195,N_23309);
and U23709 (N_23709,N_23219,N_23177);
and U23710 (N_23710,N_23372,N_22832);
xor U23711 (N_23711,N_22832,N_23338);
or U23712 (N_23712,N_23133,N_22949);
and U23713 (N_23713,N_23348,N_23132);
or U23714 (N_23714,N_22962,N_23248);
or U23715 (N_23715,N_23269,N_23051);
and U23716 (N_23716,N_22861,N_22903);
nor U23717 (N_23717,N_23038,N_22937);
or U23718 (N_23718,N_23196,N_23147);
or U23719 (N_23719,N_22989,N_23115);
nor U23720 (N_23720,N_22809,N_22922);
nor U23721 (N_23721,N_23182,N_23191);
xor U23722 (N_23722,N_23038,N_23151);
nor U23723 (N_23723,N_22835,N_23106);
nand U23724 (N_23724,N_23019,N_23094);
and U23725 (N_23725,N_23037,N_23284);
xnor U23726 (N_23726,N_22832,N_23124);
xor U23727 (N_23727,N_22864,N_23340);
and U23728 (N_23728,N_23329,N_23292);
nand U23729 (N_23729,N_23156,N_23066);
xnor U23730 (N_23730,N_23011,N_23050);
nor U23731 (N_23731,N_23210,N_23310);
nand U23732 (N_23732,N_23335,N_22828);
nand U23733 (N_23733,N_22927,N_23181);
xnor U23734 (N_23734,N_23287,N_22858);
or U23735 (N_23735,N_23331,N_23238);
and U23736 (N_23736,N_23071,N_22820);
or U23737 (N_23737,N_23346,N_23396);
nor U23738 (N_23738,N_23154,N_23290);
nor U23739 (N_23739,N_23339,N_22852);
and U23740 (N_23740,N_23193,N_22998);
and U23741 (N_23741,N_23333,N_23394);
xor U23742 (N_23742,N_23341,N_23181);
nand U23743 (N_23743,N_22833,N_23309);
xnor U23744 (N_23744,N_23070,N_23254);
and U23745 (N_23745,N_22809,N_22814);
xnor U23746 (N_23746,N_22803,N_23236);
and U23747 (N_23747,N_22977,N_23329);
nand U23748 (N_23748,N_23135,N_22962);
and U23749 (N_23749,N_23089,N_22904);
nand U23750 (N_23750,N_22930,N_22966);
nand U23751 (N_23751,N_22942,N_23349);
nor U23752 (N_23752,N_23245,N_23201);
xor U23753 (N_23753,N_23353,N_23094);
or U23754 (N_23754,N_23015,N_23244);
or U23755 (N_23755,N_22927,N_23363);
xor U23756 (N_23756,N_23155,N_22943);
nand U23757 (N_23757,N_23289,N_22986);
nor U23758 (N_23758,N_23206,N_23355);
nand U23759 (N_23759,N_22979,N_23013);
nor U23760 (N_23760,N_22902,N_23211);
and U23761 (N_23761,N_23101,N_23234);
and U23762 (N_23762,N_22931,N_23378);
xnor U23763 (N_23763,N_22963,N_23312);
nor U23764 (N_23764,N_23282,N_23176);
nand U23765 (N_23765,N_23339,N_22870);
nor U23766 (N_23766,N_23049,N_23251);
and U23767 (N_23767,N_23159,N_22887);
nand U23768 (N_23768,N_23113,N_23114);
or U23769 (N_23769,N_23048,N_23221);
nor U23770 (N_23770,N_23336,N_23111);
and U23771 (N_23771,N_22845,N_23146);
nand U23772 (N_23772,N_23290,N_23274);
nand U23773 (N_23773,N_23141,N_23261);
or U23774 (N_23774,N_23278,N_23105);
or U23775 (N_23775,N_23287,N_22918);
xor U23776 (N_23776,N_22882,N_23208);
xor U23777 (N_23777,N_23339,N_23029);
nand U23778 (N_23778,N_23030,N_22963);
nor U23779 (N_23779,N_23143,N_22999);
nor U23780 (N_23780,N_23064,N_23071);
and U23781 (N_23781,N_23123,N_23342);
nor U23782 (N_23782,N_22890,N_23077);
xor U23783 (N_23783,N_23297,N_23076);
xnor U23784 (N_23784,N_23293,N_23009);
or U23785 (N_23785,N_23265,N_22862);
nand U23786 (N_23786,N_23005,N_23344);
or U23787 (N_23787,N_23217,N_23258);
nand U23788 (N_23788,N_23185,N_23396);
and U23789 (N_23789,N_23381,N_22968);
or U23790 (N_23790,N_23015,N_22804);
nand U23791 (N_23791,N_22841,N_23341);
and U23792 (N_23792,N_22892,N_22974);
nand U23793 (N_23793,N_23296,N_23239);
or U23794 (N_23794,N_23381,N_23280);
xnor U23795 (N_23795,N_22857,N_22849);
nand U23796 (N_23796,N_22981,N_23037);
nor U23797 (N_23797,N_22895,N_23031);
xnor U23798 (N_23798,N_23031,N_23150);
or U23799 (N_23799,N_23212,N_23329);
and U23800 (N_23800,N_22889,N_22983);
xnor U23801 (N_23801,N_22979,N_23340);
nand U23802 (N_23802,N_23126,N_22948);
or U23803 (N_23803,N_23152,N_22985);
or U23804 (N_23804,N_23008,N_23161);
xor U23805 (N_23805,N_23004,N_23007);
nand U23806 (N_23806,N_23143,N_23028);
nand U23807 (N_23807,N_23268,N_23264);
nor U23808 (N_23808,N_23062,N_23350);
or U23809 (N_23809,N_23171,N_22921);
nand U23810 (N_23810,N_23050,N_23350);
xor U23811 (N_23811,N_22846,N_23299);
nand U23812 (N_23812,N_23010,N_23109);
or U23813 (N_23813,N_22970,N_23020);
nand U23814 (N_23814,N_22817,N_23321);
and U23815 (N_23815,N_22806,N_23156);
or U23816 (N_23816,N_22911,N_22967);
xor U23817 (N_23817,N_23213,N_23384);
and U23818 (N_23818,N_23045,N_23353);
nand U23819 (N_23819,N_23051,N_22986);
nor U23820 (N_23820,N_23348,N_22919);
nand U23821 (N_23821,N_23295,N_23284);
xor U23822 (N_23822,N_23121,N_23380);
or U23823 (N_23823,N_23094,N_23335);
and U23824 (N_23824,N_23226,N_22838);
xnor U23825 (N_23825,N_22829,N_22866);
or U23826 (N_23826,N_23095,N_23260);
or U23827 (N_23827,N_22837,N_23170);
or U23828 (N_23828,N_23011,N_23369);
nand U23829 (N_23829,N_23112,N_23295);
and U23830 (N_23830,N_23137,N_23145);
xor U23831 (N_23831,N_22854,N_23335);
xor U23832 (N_23832,N_22867,N_23397);
xnor U23833 (N_23833,N_22932,N_22935);
and U23834 (N_23834,N_23317,N_22889);
xnor U23835 (N_23835,N_23161,N_23094);
and U23836 (N_23836,N_23123,N_23168);
xor U23837 (N_23837,N_23333,N_23358);
and U23838 (N_23838,N_23027,N_22802);
nand U23839 (N_23839,N_22974,N_22829);
xnor U23840 (N_23840,N_23027,N_23390);
and U23841 (N_23841,N_23275,N_23207);
or U23842 (N_23842,N_22838,N_23033);
xnor U23843 (N_23843,N_22848,N_22927);
and U23844 (N_23844,N_23176,N_22946);
nand U23845 (N_23845,N_23095,N_22894);
xnor U23846 (N_23846,N_23340,N_23048);
or U23847 (N_23847,N_23063,N_22848);
and U23848 (N_23848,N_22915,N_23126);
or U23849 (N_23849,N_23339,N_22895);
or U23850 (N_23850,N_23076,N_22891);
nor U23851 (N_23851,N_23121,N_22806);
xor U23852 (N_23852,N_22873,N_23121);
or U23853 (N_23853,N_23160,N_22800);
xnor U23854 (N_23854,N_22847,N_23074);
xnor U23855 (N_23855,N_23220,N_23356);
nor U23856 (N_23856,N_22950,N_23047);
xor U23857 (N_23857,N_23185,N_23389);
xor U23858 (N_23858,N_23274,N_23054);
nor U23859 (N_23859,N_23015,N_22916);
nand U23860 (N_23860,N_22957,N_23197);
or U23861 (N_23861,N_23398,N_22909);
nor U23862 (N_23862,N_23086,N_22827);
nand U23863 (N_23863,N_23164,N_23090);
and U23864 (N_23864,N_22957,N_22882);
nor U23865 (N_23865,N_22917,N_23108);
and U23866 (N_23866,N_23144,N_23214);
or U23867 (N_23867,N_23077,N_23214);
or U23868 (N_23868,N_23023,N_22894);
xor U23869 (N_23869,N_22816,N_23166);
nand U23870 (N_23870,N_23074,N_23370);
and U23871 (N_23871,N_23238,N_23219);
or U23872 (N_23872,N_23358,N_23212);
or U23873 (N_23873,N_23030,N_23009);
and U23874 (N_23874,N_22826,N_23217);
nand U23875 (N_23875,N_23363,N_23330);
nand U23876 (N_23876,N_22953,N_23017);
nor U23877 (N_23877,N_23167,N_22986);
or U23878 (N_23878,N_23147,N_22860);
nand U23879 (N_23879,N_23195,N_23347);
nand U23880 (N_23880,N_22974,N_23106);
and U23881 (N_23881,N_23286,N_22952);
and U23882 (N_23882,N_23347,N_23242);
nand U23883 (N_23883,N_23303,N_23093);
xor U23884 (N_23884,N_23353,N_22910);
nand U23885 (N_23885,N_23373,N_23272);
xnor U23886 (N_23886,N_23062,N_23363);
nor U23887 (N_23887,N_23266,N_23027);
xor U23888 (N_23888,N_23236,N_23376);
nor U23889 (N_23889,N_23295,N_23267);
and U23890 (N_23890,N_23043,N_23109);
nor U23891 (N_23891,N_23306,N_23377);
and U23892 (N_23892,N_22993,N_22933);
nand U23893 (N_23893,N_22882,N_23195);
and U23894 (N_23894,N_23290,N_23121);
and U23895 (N_23895,N_22847,N_23220);
nand U23896 (N_23896,N_22903,N_23225);
xor U23897 (N_23897,N_22987,N_23178);
or U23898 (N_23898,N_23214,N_23211);
nand U23899 (N_23899,N_23022,N_22991);
or U23900 (N_23900,N_23195,N_23132);
nor U23901 (N_23901,N_22954,N_23244);
xor U23902 (N_23902,N_23254,N_23136);
nand U23903 (N_23903,N_23266,N_22994);
and U23904 (N_23904,N_23354,N_23181);
xor U23905 (N_23905,N_22974,N_23204);
or U23906 (N_23906,N_23363,N_23356);
or U23907 (N_23907,N_22914,N_23263);
xor U23908 (N_23908,N_22858,N_23333);
xnor U23909 (N_23909,N_23255,N_22936);
nor U23910 (N_23910,N_23128,N_23222);
and U23911 (N_23911,N_22961,N_22931);
xnor U23912 (N_23912,N_23232,N_22837);
nor U23913 (N_23913,N_22892,N_23060);
nor U23914 (N_23914,N_23210,N_23279);
nand U23915 (N_23915,N_22920,N_23323);
xnor U23916 (N_23916,N_23246,N_22850);
and U23917 (N_23917,N_23042,N_23178);
or U23918 (N_23918,N_22955,N_23159);
nor U23919 (N_23919,N_23016,N_22894);
xnor U23920 (N_23920,N_23035,N_23127);
nor U23921 (N_23921,N_23266,N_22942);
nor U23922 (N_23922,N_23187,N_22981);
or U23923 (N_23923,N_22939,N_22953);
or U23924 (N_23924,N_22987,N_23093);
xor U23925 (N_23925,N_23106,N_23332);
nand U23926 (N_23926,N_23187,N_22988);
nand U23927 (N_23927,N_23288,N_22996);
nand U23928 (N_23928,N_23258,N_23114);
or U23929 (N_23929,N_22915,N_23033);
nand U23930 (N_23930,N_22826,N_23376);
xnor U23931 (N_23931,N_22819,N_23373);
nand U23932 (N_23932,N_23191,N_22834);
nor U23933 (N_23933,N_23156,N_22829);
or U23934 (N_23934,N_23034,N_22839);
nor U23935 (N_23935,N_23319,N_22846);
or U23936 (N_23936,N_23368,N_22862);
nor U23937 (N_23937,N_23211,N_23293);
nand U23938 (N_23938,N_23101,N_23206);
nor U23939 (N_23939,N_22972,N_23196);
nor U23940 (N_23940,N_22954,N_22917);
nand U23941 (N_23941,N_22920,N_22885);
and U23942 (N_23942,N_23197,N_23272);
and U23943 (N_23943,N_23040,N_22846);
or U23944 (N_23944,N_22980,N_23295);
nand U23945 (N_23945,N_23317,N_23260);
xor U23946 (N_23946,N_23155,N_22817);
or U23947 (N_23947,N_23055,N_23392);
and U23948 (N_23948,N_23192,N_23004);
or U23949 (N_23949,N_23286,N_22824);
nor U23950 (N_23950,N_23071,N_22848);
or U23951 (N_23951,N_23349,N_22986);
or U23952 (N_23952,N_22858,N_22909);
and U23953 (N_23953,N_23079,N_23213);
or U23954 (N_23954,N_23330,N_22994);
nor U23955 (N_23955,N_23249,N_22818);
nor U23956 (N_23956,N_23193,N_23317);
or U23957 (N_23957,N_23068,N_23366);
xor U23958 (N_23958,N_23170,N_22965);
nor U23959 (N_23959,N_23366,N_23355);
or U23960 (N_23960,N_23353,N_22842);
or U23961 (N_23961,N_23081,N_23048);
nor U23962 (N_23962,N_23282,N_23088);
nor U23963 (N_23963,N_23221,N_23348);
nand U23964 (N_23964,N_22829,N_23109);
nor U23965 (N_23965,N_23269,N_23240);
nand U23966 (N_23966,N_23172,N_23361);
xor U23967 (N_23967,N_23351,N_22893);
xnor U23968 (N_23968,N_23120,N_22830);
or U23969 (N_23969,N_23244,N_23066);
and U23970 (N_23970,N_22970,N_22813);
nand U23971 (N_23971,N_23393,N_22997);
or U23972 (N_23972,N_23158,N_23357);
xor U23973 (N_23973,N_22833,N_22987);
or U23974 (N_23974,N_22961,N_23046);
or U23975 (N_23975,N_23349,N_22958);
or U23976 (N_23976,N_23105,N_23024);
nand U23977 (N_23977,N_23220,N_23072);
nand U23978 (N_23978,N_22825,N_22837);
xor U23979 (N_23979,N_23021,N_22954);
xor U23980 (N_23980,N_23209,N_23384);
nor U23981 (N_23981,N_23117,N_22864);
or U23982 (N_23982,N_23228,N_22838);
xnor U23983 (N_23983,N_23054,N_23201);
xor U23984 (N_23984,N_23396,N_23359);
xor U23985 (N_23985,N_22867,N_23221);
nor U23986 (N_23986,N_22973,N_22957);
xor U23987 (N_23987,N_23334,N_23186);
nand U23988 (N_23988,N_22865,N_23160);
or U23989 (N_23989,N_23100,N_23046);
nand U23990 (N_23990,N_23252,N_22876);
xnor U23991 (N_23991,N_23319,N_22865);
or U23992 (N_23992,N_23020,N_22974);
or U23993 (N_23993,N_23307,N_22805);
nand U23994 (N_23994,N_22841,N_23302);
nand U23995 (N_23995,N_23214,N_22967);
xor U23996 (N_23996,N_23360,N_23151);
nor U23997 (N_23997,N_23258,N_23190);
nor U23998 (N_23998,N_23329,N_22859);
and U23999 (N_23999,N_23313,N_22854);
nor U24000 (N_24000,N_23833,N_23596);
and U24001 (N_24001,N_23904,N_23960);
xor U24002 (N_24002,N_23923,N_23490);
xnor U24003 (N_24003,N_23853,N_23629);
nor U24004 (N_24004,N_23901,N_23911);
or U24005 (N_24005,N_23869,N_23501);
xnor U24006 (N_24006,N_23761,N_23829);
xnor U24007 (N_24007,N_23456,N_23788);
nand U24008 (N_24008,N_23451,N_23733);
or U24009 (N_24009,N_23509,N_23540);
xnor U24010 (N_24010,N_23422,N_23500);
xor U24011 (N_24011,N_23618,N_23494);
nand U24012 (N_24012,N_23408,N_23903);
nand U24013 (N_24013,N_23782,N_23493);
xor U24014 (N_24014,N_23866,N_23816);
nand U24015 (N_24015,N_23675,N_23971);
and U24016 (N_24016,N_23663,N_23569);
and U24017 (N_24017,N_23822,N_23699);
and U24018 (N_24018,N_23900,N_23760);
nand U24019 (N_24019,N_23450,N_23842);
and U24020 (N_24020,N_23909,N_23514);
nand U24021 (N_24021,N_23669,N_23639);
nor U24022 (N_24022,N_23885,N_23849);
nand U24023 (N_24023,N_23735,N_23654);
and U24024 (N_24024,N_23440,N_23640);
nand U24025 (N_24025,N_23883,N_23870);
or U24026 (N_24026,N_23465,N_23492);
xor U24027 (N_24027,N_23448,N_23820);
nand U24028 (N_24028,N_23527,N_23600);
or U24029 (N_24029,N_23779,N_23617);
and U24030 (N_24030,N_23928,N_23586);
nand U24031 (N_24031,N_23996,N_23589);
and U24032 (N_24032,N_23466,N_23786);
and U24033 (N_24033,N_23957,N_23576);
and U24034 (N_24034,N_23970,N_23848);
or U24035 (N_24035,N_23799,N_23687);
and U24036 (N_24036,N_23955,N_23621);
nand U24037 (N_24037,N_23886,N_23910);
or U24038 (N_24038,N_23716,N_23784);
or U24039 (N_24039,N_23562,N_23858);
or U24040 (N_24040,N_23752,N_23495);
or U24041 (N_24041,N_23993,N_23859);
or U24042 (N_24042,N_23845,N_23682);
xor U24043 (N_24043,N_23704,N_23726);
nor U24044 (N_24044,N_23579,N_23933);
nand U24045 (N_24045,N_23830,N_23964);
or U24046 (N_24046,N_23718,N_23815);
nor U24047 (N_24047,N_23470,N_23624);
or U24048 (N_24048,N_23953,N_23647);
nand U24049 (N_24049,N_23787,N_23980);
xor U24050 (N_24050,N_23918,N_23432);
nand U24051 (N_24051,N_23839,N_23413);
or U24052 (N_24052,N_23539,N_23550);
xor U24053 (N_24053,N_23890,N_23502);
or U24054 (N_24054,N_23537,N_23952);
nor U24055 (N_24055,N_23747,N_23671);
or U24056 (N_24056,N_23659,N_23513);
or U24057 (N_24057,N_23604,N_23685);
nand U24058 (N_24058,N_23677,N_23414);
nor U24059 (N_24059,N_23504,N_23857);
nor U24060 (N_24060,N_23731,N_23547);
nor U24061 (N_24061,N_23407,N_23945);
nor U24062 (N_24062,N_23692,N_23518);
and U24063 (N_24063,N_23622,N_23558);
xor U24064 (N_24064,N_23744,N_23442);
xor U24065 (N_24065,N_23931,N_23420);
xor U24066 (N_24066,N_23631,N_23989);
and U24067 (N_24067,N_23568,N_23723);
xor U24068 (N_24068,N_23976,N_23482);
nand U24069 (N_24069,N_23906,N_23444);
nand U24070 (N_24070,N_23905,N_23535);
and U24071 (N_24071,N_23472,N_23481);
xnor U24072 (N_24072,N_23628,N_23423);
nand U24073 (N_24073,N_23690,N_23561);
and U24074 (N_24074,N_23917,N_23710);
or U24075 (N_24075,N_23524,N_23860);
and U24076 (N_24076,N_23555,N_23646);
xnor U24077 (N_24077,N_23552,N_23814);
nor U24078 (N_24078,N_23889,N_23963);
xor U24079 (N_24079,N_23874,N_23881);
nand U24080 (N_24080,N_23431,N_23656);
and U24081 (N_24081,N_23892,N_23672);
xnor U24082 (N_24082,N_23427,N_23824);
nand U24083 (N_24083,N_23651,N_23843);
or U24084 (N_24084,N_23770,N_23975);
nand U24085 (N_24085,N_23566,N_23584);
nand U24086 (N_24086,N_23678,N_23499);
or U24087 (N_24087,N_23532,N_23411);
nor U24088 (N_24088,N_23581,N_23673);
nand U24089 (N_24089,N_23962,N_23400);
nand U24090 (N_24090,N_23523,N_23762);
and U24091 (N_24091,N_23878,N_23734);
and U24092 (N_24092,N_23553,N_23438);
nand U24093 (N_24093,N_23441,N_23832);
nor U24094 (N_24094,N_23597,N_23412);
nand U24095 (N_24095,N_23825,N_23759);
nand U24096 (N_24096,N_23608,N_23999);
xor U24097 (N_24097,N_23473,N_23491);
nor U24098 (N_24098,N_23961,N_23425);
xnor U24099 (N_24099,N_23912,N_23577);
and U24100 (N_24100,N_23988,N_23769);
and U24101 (N_24101,N_23697,N_23609);
xor U24102 (N_24102,N_23560,N_23474);
xnor U24103 (N_24103,N_23968,N_23781);
and U24104 (N_24104,N_23700,N_23691);
xor U24105 (N_24105,N_23614,N_23969);
and U24106 (N_24106,N_23611,N_23635);
nand U24107 (N_24107,N_23668,N_23938);
nor U24108 (N_24108,N_23409,N_23876);
and U24109 (N_24109,N_23997,N_23974);
or U24110 (N_24110,N_23467,N_23879);
and U24111 (N_24111,N_23517,N_23670);
and U24112 (N_24112,N_23947,N_23741);
xnor U24113 (N_24113,N_23793,N_23606);
nor U24114 (N_24114,N_23913,N_23926);
nor U24115 (N_24115,N_23486,N_23683);
or U24116 (N_24116,N_23521,N_23994);
or U24117 (N_24117,N_23462,N_23454);
nor U24118 (N_24118,N_23705,N_23840);
nor U24119 (N_24119,N_23607,N_23772);
xnor U24120 (N_24120,N_23959,N_23534);
nand U24121 (N_24121,N_23636,N_23895);
nand U24122 (N_24122,N_23946,N_23686);
and U24123 (N_24123,N_23455,N_23437);
or U24124 (N_24124,N_23661,N_23585);
nand U24125 (N_24125,N_23823,N_23739);
nor U24126 (N_24126,N_23632,N_23755);
and U24127 (N_24127,N_23757,N_23542);
and U24128 (N_24128,N_23593,N_23696);
nand U24129 (N_24129,N_23520,N_23819);
xnor U24130 (N_24130,N_23867,N_23863);
nor U24131 (N_24131,N_23873,N_23754);
or U24132 (N_24132,N_23446,N_23736);
nand U24133 (N_24133,N_23851,N_23655);
xnor U24134 (N_24134,N_23844,N_23806);
and U24135 (N_24135,N_23557,N_23526);
nor U24136 (N_24136,N_23775,N_23485);
nor U24137 (N_24137,N_23469,N_23573);
nor U24138 (N_24138,N_23914,N_23496);
or U24139 (N_24139,N_23554,N_23835);
and U24140 (N_24140,N_23460,N_23740);
xnor U24141 (N_24141,N_23801,N_23538);
nand U24142 (N_24142,N_23694,N_23642);
xnor U24143 (N_24143,N_23689,N_23464);
or U24144 (N_24144,N_23737,N_23877);
nor U24145 (N_24145,N_23443,N_23613);
and U24146 (N_24146,N_23765,N_23846);
nor U24147 (N_24147,N_23748,N_23461);
or U24148 (N_24148,N_23983,N_23891);
or U24149 (N_24149,N_23536,N_23567);
xnor U24150 (N_24150,N_23986,N_23813);
and U24151 (N_24151,N_23602,N_23447);
and U24152 (N_24152,N_23476,N_23459);
xnor U24153 (N_24153,N_23920,N_23641);
or U24154 (N_24154,N_23954,N_23809);
nor U24155 (N_24155,N_23803,N_23882);
and U24156 (N_24156,N_23528,N_23591);
xor U24157 (N_24157,N_23750,N_23771);
nor U24158 (N_24158,N_23410,N_23800);
or U24159 (N_24159,N_23942,N_23712);
nor U24160 (N_24160,N_23990,N_23966);
xor U24161 (N_24161,N_23559,N_23680);
xor U24162 (N_24162,N_23565,N_23574);
nand U24163 (N_24163,N_23834,N_23403);
nor U24164 (N_24164,N_23479,N_23643);
and U24165 (N_24165,N_23615,N_23753);
nor U24166 (N_24166,N_23714,N_23637);
nor U24167 (N_24167,N_23548,N_23807);
nor U24168 (N_24168,N_23648,N_23727);
nand U24169 (N_24169,N_23850,N_23977);
nor U24170 (N_24170,N_23506,N_23545);
nor U24171 (N_24171,N_23929,N_23452);
nor U24172 (N_24172,N_23595,N_23907);
nand U24173 (N_24173,N_23480,N_23941);
or U24174 (N_24174,N_23798,N_23664);
nor U24175 (N_24175,N_23838,N_23688);
and U24176 (N_24176,N_23575,N_23507);
xor U24177 (N_24177,N_23415,N_23984);
nand U24178 (N_24178,N_23828,N_23936);
xor U24179 (N_24179,N_23871,N_23603);
nor U24180 (N_24180,N_23525,N_23489);
nand U24181 (N_24181,N_23533,N_23658);
and U24182 (N_24182,N_23570,N_23638);
nand U24183 (N_24183,N_23665,N_23483);
or U24184 (N_24184,N_23797,N_23921);
and U24185 (N_24185,N_23973,N_23836);
nor U24186 (N_24186,N_23949,N_23939);
nor U24187 (N_24187,N_23572,N_23995);
nor U24188 (N_24188,N_23660,N_23657);
or U24189 (N_24189,N_23897,N_23987);
and U24190 (N_24190,N_23630,N_23457);
xnor U24191 (N_24191,N_23601,N_23783);
nand U24192 (N_24192,N_23743,N_23551);
nor U24193 (N_24193,N_23676,N_23512);
and U24194 (N_24194,N_23543,N_23580);
and U24195 (N_24195,N_23854,N_23826);
and U24196 (N_24196,N_23777,N_23544);
nand U24197 (N_24197,N_23531,N_23902);
nand U24198 (N_24198,N_23426,N_23667);
xnor U24199 (N_24199,N_23571,N_23898);
xnor U24200 (N_24200,N_23713,N_23893);
nor U24201 (N_24201,N_23767,N_23896);
and U24202 (N_24202,N_23421,N_23841);
and U24203 (N_24203,N_23721,N_23702);
nand U24204 (N_24204,N_23818,N_23888);
and U24205 (N_24205,N_23563,N_23796);
nand U24206 (N_24206,N_23430,N_23649);
and U24207 (N_24207,N_23695,N_23619);
or U24208 (N_24208,N_23717,N_23416);
nor U24209 (N_24209,N_23445,N_23868);
or U24210 (N_24210,N_23471,N_23666);
nand U24211 (N_24211,N_23634,N_23530);
nand U24212 (N_24212,N_23653,N_23745);
xor U24213 (N_24213,N_23763,N_23728);
nand U24214 (N_24214,N_23764,N_23645);
and U24215 (N_24215,N_23436,N_23674);
or U24216 (N_24216,N_23458,N_23556);
xnor U24217 (N_24217,N_23505,N_23402);
or U24218 (N_24218,N_23852,N_23616);
or U24219 (N_24219,N_23605,N_23729);
nor U24220 (N_24220,N_23428,N_23419);
nand U24221 (N_24221,N_23434,N_23488);
xnor U24222 (N_24222,N_23880,N_23698);
nand U24223 (N_24223,N_23644,N_23623);
xnor U24224 (N_24224,N_23406,N_23522);
or U24225 (N_24225,N_23679,N_23681);
nand U24226 (N_24226,N_23915,N_23706);
xnor U24227 (N_24227,N_23684,N_23855);
or U24228 (N_24228,N_23732,N_23497);
xnor U24229 (N_24229,N_23780,N_23992);
nor U24230 (N_24230,N_23956,N_23592);
nand U24231 (N_24231,N_23773,N_23404);
and U24232 (N_24232,N_23435,N_23894);
nand U24233 (N_24233,N_23982,N_23919);
xnor U24234 (N_24234,N_23872,N_23937);
nand U24235 (N_24235,N_23429,N_23967);
xnor U24236 (N_24236,N_23758,N_23564);
and U24237 (N_24237,N_23932,N_23707);
or U24238 (N_24238,N_23711,N_23943);
and U24239 (N_24239,N_23519,N_23865);
nand U24240 (N_24240,N_23701,N_23503);
nor U24241 (N_24241,N_23862,N_23417);
and U24242 (N_24242,N_23720,N_23985);
xnor U24243 (N_24243,N_23940,N_23484);
nand U24244 (N_24244,N_23511,N_23510);
nand U24245 (N_24245,N_23612,N_23626);
or U24246 (N_24246,N_23908,N_23746);
xnor U24247 (N_24247,N_23722,N_23715);
nor U24248 (N_24248,N_23463,N_23590);
and U24249 (N_24249,N_23810,N_23925);
and U24250 (N_24250,N_23477,N_23978);
xor U24251 (N_24251,N_23756,N_23792);
and U24252 (N_24252,N_23927,N_23709);
or U24253 (N_24253,N_23725,N_23821);
nand U24254 (N_24254,N_23487,N_23981);
and U24255 (N_24255,N_23625,N_23508);
nand U24256 (N_24256,N_23827,N_23899);
and U24257 (N_24257,N_23478,N_23738);
nor U24258 (N_24258,N_23847,N_23944);
nand U24259 (N_24259,N_23778,N_23498);
and U24260 (N_24260,N_23774,N_23516);
nand U24261 (N_24261,N_23439,N_23998);
or U24262 (N_24262,N_23965,N_23875);
nor U24263 (N_24263,N_23768,N_23587);
xnor U24264 (N_24264,N_23627,N_23958);
nor U24265 (N_24265,N_23703,N_23856);
or U24266 (N_24266,N_23529,N_23749);
xor U24267 (N_24267,N_23950,N_23449);
nand U24268 (N_24268,N_23433,N_23650);
xnor U24269 (N_24269,N_23837,N_23594);
nor U24270 (N_24270,N_23812,N_23418);
nand U24271 (N_24271,N_23951,N_23453);
and U24272 (N_24272,N_23405,N_23401);
and U24273 (N_24273,N_23934,N_23662);
or U24274 (N_24274,N_23817,N_23766);
or U24275 (N_24275,N_23719,N_23884);
or U24276 (N_24276,N_23610,N_23794);
nor U24277 (N_24277,N_23991,N_23808);
xnor U24278 (N_24278,N_23541,N_23811);
nand U24279 (N_24279,N_23930,N_23652);
or U24280 (N_24280,N_23582,N_23924);
nand U24281 (N_24281,N_23588,N_23795);
and U24282 (N_24282,N_23776,N_23751);
xnor U24283 (N_24283,N_23546,N_23549);
nand U24284 (N_24284,N_23598,N_23935);
nor U24285 (N_24285,N_23468,N_23831);
or U24286 (N_24286,N_23633,N_23789);
nand U24287 (N_24287,N_23424,N_23979);
nand U24288 (N_24288,N_23864,N_23730);
xor U24289 (N_24289,N_23620,N_23922);
xnor U24290 (N_24290,N_23475,N_23578);
or U24291 (N_24291,N_23861,N_23708);
nand U24292 (N_24292,N_23804,N_23805);
and U24293 (N_24293,N_23790,N_23515);
and U24294 (N_24294,N_23948,N_23802);
and U24295 (N_24295,N_23785,N_23972);
nor U24296 (N_24296,N_23742,N_23791);
nor U24297 (N_24297,N_23583,N_23887);
or U24298 (N_24298,N_23693,N_23599);
or U24299 (N_24299,N_23916,N_23724);
nand U24300 (N_24300,N_23825,N_23532);
or U24301 (N_24301,N_23832,N_23901);
xnor U24302 (N_24302,N_23998,N_23415);
nand U24303 (N_24303,N_23519,N_23607);
nor U24304 (N_24304,N_23778,N_23533);
or U24305 (N_24305,N_23444,N_23828);
nand U24306 (N_24306,N_23619,N_23649);
xor U24307 (N_24307,N_23448,N_23618);
nor U24308 (N_24308,N_23811,N_23823);
and U24309 (N_24309,N_23638,N_23725);
or U24310 (N_24310,N_23791,N_23836);
or U24311 (N_24311,N_23776,N_23810);
and U24312 (N_24312,N_23664,N_23890);
and U24313 (N_24313,N_23824,N_23648);
nand U24314 (N_24314,N_23612,N_23971);
nand U24315 (N_24315,N_23710,N_23568);
or U24316 (N_24316,N_23760,N_23775);
and U24317 (N_24317,N_23481,N_23498);
xor U24318 (N_24318,N_23883,N_23765);
nor U24319 (N_24319,N_23677,N_23568);
nor U24320 (N_24320,N_23836,N_23970);
and U24321 (N_24321,N_23966,N_23985);
nor U24322 (N_24322,N_23883,N_23588);
or U24323 (N_24323,N_23902,N_23416);
nand U24324 (N_24324,N_23564,N_23739);
nor U24325 (N_24325,N_23414,N_23783);
nand U24326 (N_24326,N_23622,N_23544);
xor U24327 (N_24327,N_23994,N_23409);
and U24328 (N_24328,N_23925,N_23411);
and U24329 (N_24329,N_23994,N_23661);
and U24330 (N_24330,N_23517,N_23989);
xnor U24331 (N_24331,N_23996,N_23656);
xor U24332 (N_24332,N_23952,N_23780);
xor U24333 (N_24333,N_23442,N_23580);
nand U24334 (N_24334,N_23984,N_23440);
and U24335 (N_24335,N_23650,N_23916);
or U24336 (N_24336,N_23836,N_23642);
xnor U24337 (N_24337,N_23979,N_23433);
and U24338 (N_24338,N_23806,N_23837);
nand U24339 (N_24339,N_23550,N_23893);
nor U24340 (N_24340,N_23474,N_23615);
or U24341 (N_24341,N_23497,N_23702);
nor U24342 (N_24342,N_23989,N_23429);
nand U24343 (N_24343,N_23831,N_23408);
nor U24344 (N_24344,N_23537,N_23652);
xnor U24345 (N_24345,N_23613,N_23441);
or U24346 (N_24346,N_23905,N_23835);
xor U24347 (N_24347,N_23778,N_23806);
nand U24348 (N_24348,N_23904,N_23528);
nor U24349 (N_24349,N_23689,N_23613);
or U24350 (N_24350,N_23599,N_23898);
xnor U24351 (N_24351,N_23895,N_23453);
and U24352 (N_24352,N_23836,N_23852);
or U24353 (N_24353,N_23437,N_23484);
or U24354 (N_24354,N_23860,N_23439);
xnor U24355 (N_24355,N_23778,N_23528);
xor U24356 (N_24356,N_23693,N_23602);
nor U24357 (N_24357,N_23944,N_23430);
or U24358 (N_24358,N_23889,N_23555);
nor U24359 (N_24359,N_23600,N_23846);
xor U24360 (N_24360,N_23834,N_23860);
nand U24361 (N_24361,N_23668,N_23450);
nand U24362 (N_24362,N_23493,N_23873);
nand U24363 (N_24363,N_23761,N_23741);
nand U24364 (N_24364,N_23704,N_23801);
xnor U24365 (N_24365,N_23993,N_23935);
and U24366 (N_24366,N_23606,N_23730);
xor U24367 (N_24367,N_23462,N_23900);
or U24368 (N_24368,N_23478,N_23525);
nor U24369 (N_24369,N_23921,N_23927);
or U24370 (N_24370,N_23479,N_23533);
nand U24371 (N_24371,N_23670,N_23594);
nand U24372 (N_24372,N_23625,N_23759);
nand U24373 (N_24373,N_23887,N_23510);
xor U24374 (N_24374,N_23476,N_23811);
and U24375 (N_24375,N_23883,N_23988);
nand U24376 (N_24376,N_23446,N_23943);
and U24377 (N_24377,N_23429,N_23530);
or U24378 (N_24378,N_23536,N_23967);
xnor U24379 (N_24379,N_23679,N_23939);
or U24380 (N_24380,N_23726,N_23660);
or U24381 (N_24381,N_23738,N_23498);
or U24382 (N_24382,N_23442,N_23718);
and U24383 (N_24383,N_23792,N_23438);
nor U24384 (N_24384,N_23460,N_23759);
and U24385 (N_24385,N_23520,N_23730);
or U24386 (N_24386,N_23620,N_23400);
nand U24387 (N_24387,N_23630,N_23623);
xnor U24388 (N_24388,N_23979,N_23451);
nor U24389 (N_24389,N_23766,N_23472);
and U24390 (N_24390,N_23642,N_23594);
or U24391 (N_24391,N_23770,N_23634);
and U24392 (N_24392,N_23586,N_23860);
nor U24393 (N_24393,N_23406,N_23401);
xnor U24394 (N_24394,N_23799,N_23959);
xor U24395 (N_24395,N_23619,N_23852);
nor U24396 (N_24396,N_23543,N_23820);
xnor U24397 (N_24397,N_23498,N_23560);
nand U24398 (N_24398,N_23735,N_23782);
and U24399 (N_24399,N_23898,N_23855);
nor U24400 (N_24400,N_23466,N_23455);
xnor U24401 (N_24401,N_23599,N_23757);
xnor U24402 (N_24402,N_23773,N_23721);
nor U24403 (N_24403,N_23933,N_23723);
nand U24404 (N_24404,N_23725,N_23610);
nor U24405 (N_24405,N_23983,N_23459);
nand U24406 (N_24406,N_23643,N_23707);
nor U24407 (N_24407,N_23503,N_23843);
nor U24408 (N_24408,N_23671,N_23907);
nor U24409 (N_24409,N_23687,N_23727);
nand U24410 (N_24410,N_23515,N_23902);
or U24411 (N_24411,N_23703,N_23999);
or U24412 (N_24412,N_23863,N_23745);
nand U24413 (N_24413,N_23454,N_23595);
nand U24414 (N_24414,N_23680,N_23492);
nand U24415 (N_24415,N_23486,N_23405);
nand U24416 (N_24416,N_23882,N_23726);
nor U24417 (N_24417,N_23791,N_23723);
and U24418 (N_24418,N_23861,N_23958);
and U24419 (N_24419,N_23872,N_23569);
or U24420 (N_24420,N_23571,N_23590);
xnor U24421 (N_24421,N_23965,N_23872);
and U24422 (N_24422,N_23805,N_23824);
or U24423 (N_24423,N_23612,N_23584);
xor U24424 (N_24424,N_23617,N_23515);
xor U24425 (N_24425,N_23702,N_23424);
nand U24426 (N_24426,N_23610,N_23550);
xor U24427 (N_24427,N_23722,N_23757);
xnor U24428 (N_24428,N_23418,N_23798);
xnor U24429 (N_24429,N_23676,N_23535);
xor U24430 (N_24430,N_23887,N_23702);
nand U24431 (N_24431,N_23610,N_23468);
xor U24432 (N_24432,N_23413,N_23708);
nor U24433 (N_24433,N_23825,N_23726);
or U24434 (N_24434,N_23852,N_23467);
or U24435 (N_24435,N_23560,N_23857);
nand U24436 (N_24436,N_23931,N_23886);
xor U24437 (N_24437,N_23468,N_23908);
nor U24438 (N_24438,N_23784,N_23898);
nand U24439 (N_24439,N_23755,N_23894);
nand U24440 (N_24440,N_23591,N_23861);
and U24441 (N_24441,N_23826,N_23427);
xnor U24442 (N_24442,N_23775,N_23790);
xor U24443 (N_24443,N_23851,N_23481);
or U24444 (N_24444,N_23485,N_23606);
xnor U24445 (N_24445,N_23901,N_23409);
and U24446 (N_24446,N_23749,N_23573);
nor U24447 (N_24447,N_23923,N_23631);
or U24448 (N_24448,N_23678,N_23636);
nor U24449 (N_24449,N_23722,N_23915);
xnor U24450 (N_24450,N_23647,N_23771);
nor U24451 (N_24451,N_23678,N_23719);
nor U24452 (N_24452,N_23598,N_23918);
and U24453 (N_24453,N_23923,N_23594);
nor U24454 (N_24454,N_23469,N_23904);
or U24455 (N_24455,N_23891,N_23772);
xor U24456 (N_24456,N_23594,N_23858);
and U24457 (N_24457,N_23623,N_23429);
or U24458 (N_24458,N_23508,N_23556);
or U24459 (N_24459,N_23913,N_23464);
nor U24460 (N_24460,N_23919,N_23426);
xor U24461 (N_24461,N_23789,N_23770);
xnor U24462 (N_24462,N_23423,N_23405);
or U24463 (N_24463,N_23871,N_23797);
nand U24464 (N_24464,N_23931,N_23512);
nor U24465 (N_24465,N_23987,N_23992);
or U24466 (N_24466,N_23594,N_23471);
nor U24467 (N_24467,N_23523,N_23908);
and U24468 (N_24468,N_23946,N_23563);
nand U24469 (N_24469,N_23821,N_23426);
or U24470 (N_24470,N_23854,N_23526);
nand U24471 (N_24471,N_23482,N_23546);
nor U24472 (N_24472,N_23535,N_23677);
nor U24473 (N_24473,N_23970,N_23743);
nor U24474 (N_24474,N_23895,N_23833);
xor U24475 (N_24475,N_23980,N_23627);
and U24476 (N_24476,N_23804,N_23452);
xnor U24477 (N_24477,N_23748,N_23754);
nand U24478 (N_24478,N_23673,N_23634);
nand U24479 (N_24479,N_23735,N_23976);
nor U24480 (N_24480,N_23895,N_23981);
or U24481 (N_24481,N_23418,N_23851);
nor U24482 (N_24482,N_23950,N_23418);
or U24483 (N_24483,N_23705,N_23409);
and U24484 (N_24484,N_23987,N_23686);
nand U24485 (N_24485,N_23876,N_23993);
or U24486 (N_24486,N_23713,N_23507);
nand U24487 (N_24487,N_23998,N_23979);
and U24488 (N_24488,N_23901,N_23615);
nand U24489 (N_24489,N_23672,N_23650);
and U24490 (N_24490,N_23750,N_23859);
nor U24491 (N_24491,N_23822,N_23970);
nor U24492 (N_24492,N_23551,N_23936);
nand U24493 (N_24493,N_23942,N_23964);
and U24494 (N_24494,N_23552,N_23599);
or U24495 (N_24495,N_23606,N_23779);
xnor U24496 (N_24496,N_23864,N_23935);
or U24497 (N_24497,N_23865,N_23993);
nor U24498 (N_24498,N_23665,N_23670);
or U24499 (N_24499,N_23987,N_23700);
or U24500 (N_24500,N_23471,N_23675);
nand U24501 (N_24501,N_23673,N_23436);
nor U24502 (N_24502,N_23934,N_23821);
or U24503 (N_24503,N_23759,N_23863);
or U24504 (N_24504,N_23442,N_23850);
nor U24505 (N_24505,N_23699,N_23756);
nor U24506 (N_24506,N_23807,N_23965);
and U24507 (N_24507,N_23860,N_23667);
nand U24508 (N_24508,N_23497,N_23635);
nor U24509 (N_24509,N_23760,N_23592);
and U24510 (N_24510,N_23951,N_23431);
and U24511 (N_24511,N_23869,N_23970);
xnor U24512 (N_24512,N_23989,N_23635);
nor U24513 (N_24513,N_23478,N_23836);
or U24514 (N_24514,N_23457,N_23576);
nand U24515 (N_24515,N_23932,N_23716);
and U24516 (N_24516,N_23826,N_23718);
nor U24517 (N_24517,N_23448,N_23794);
or U24518 (N_24518,N_23680,N_23738);
nor U24519 (N_24519,N_23684,N_23596);
and U24520 (N_24520,N_23589,N_23795);
or U24521 (N_24521,N_23680,N_23521);
and U24522 (N_24522,N_23633,N_23700);
nand U24523 (N_24523,N_23428,N_23466);
nor U24524 (N_24524,N_23865,N_23794);
or U24525 (N_24525,N_23840,N_23644);
and U24526 (N_24526,N_23852,N_23709);
xor U24527 (N_24527,N_23649,N_23861);
nor U24528 (N_24528,N_23430,N_23404);
and U24529 (N_24529,N_23513,N_23900);
or U24530 (N_24530,N_23991,N_23618);
and U24531 (N_24531,N_23941,N_23491);
nor U24532 (N_24532,N_23764,N_23894);
and U24533 (N_24533,N_23777,N_23479);
nor U24534 (N_24534,N_23834,N_23535);
xnor U24535 (N_24535,N_23560,N_23482);
xnor U24536 (N_24536,N_23776,N_23719);
nand U24537 (N_24537,N_23937,N_23705);
nand U24538 (N_24538,N_23843,N_23552);
and U24539 (N_24539,N_23862,N_23600);
and U24540 (N_24540,N_23572,N_23605);
xnor U24541 (N_24541,N_23872,N_23839);
and U24542 (N_24542,N_23824,N_23943);
and U24543 (N_24543,N_23596,N_23980);
nor U24544 (N_24544,N_23919,N_23804);
or U24545 (N_24545,N_23970,N_23610);
nor U24546 (N_24546,N_23619,N_23467);
or U24547 (N_24547,N_23667,N_23862);
xnor U24548 (N_24548,N_23665,N_23503);
xor U24549 (N_24549,N_23482,N_23821);
xnor U24550 (N_24550,N_23868,N_23783);
xnor U24551 (N_24551,N_23575,N_23614);
xnor U24552 (N_24552,N_23837,N_23911);
and U24553 (N_24553,N_23853,N_23511);
nor U24554 (N_24554,N_23464,N_23789);
or U24555 (N_24555,N_23456,N_23583);
xnor U24556 (N_24556,N_23795,N_23524);
nor U24557 (N_24557,N_23440,N_23835);
xnor U24558 (N_24558,N_23892,N_23717);
xor U24559 (N_24559,N_23516,N_23454);
or U24560 (N_24560,N_23890,N_23409);
xor U24561 (N_24561,N_23741,N_23817);
and U24562 (N_24562,N_23556,N_23945);
xor U24563 (N_24563,N_23686,N_23643);
or U24564 (N_24564,N_23840,N_23516);
nand U24565 (N_24565,N_23943,N_23952);
or U24566 (N_24566,N_23487,N_23753);
and U24567 (N_24567,N_23519,N_23994);
and U24568 (N_24568,N_23777,N_23994);
nand U24569 (N_24569,N_23577,N_23855);
or U24570 (N_24570,N_23824,N_23632);
or U24571 (N_24571,N_23774,N_23722);
nor U24572 (N_24572,N_23888,N_23808);
xor U24573 (N_24573,N_23507,N_23599);
or U24574 (N_24574,N_23631,N_23560);
and U24575 (N_24575,N_23476,N_23513);
nor U24576 (N_24576,N_23718,N_23429);
xnor U24577 (N_24577,N_23859,N_23628);
xor U24578 (N_24578,N_23492,N_23775);
or U24579 (N_24579,N_23847,N_23867);
or U24580 (N_24580,N_23843,N_23462);
xnor U24581 (N_24581,N_23436,N_23464);
and U24582 (N_24582,N_23710,N_23890);
nor U24583 (N_24583,N_23686,N_23824);
xor U24584 (N_24584,N_23762,N_23608);
or U24585 (N_24585,N_23711,N_23506);
nand U24586 (N_24586,N_23727,N_23772);
and U24587 (N_24587,N_23660,N_23528);
or U24588 (N_24588,N_23813,N_23835);
xor U24589 (N_24589,N_23477,N_23855);
nand U24590 (N_24590,N_23574,N_23774);
or U24591 (N_24591,N_23803,N_23444);
xnor U24592 (N_24592,N_23985,N_23736);
xor U24593 (N_24593,N_23976,N_23773);
or U24594 (N_24594,N_23565,N_23606);
or U24595 (N_24595,N_23600,N_23958);
and U24596 (N_24596,N_23937,N_23631);
or U24597 (N_24597,N_23714,N_23789);
and U24598 (N_24598,N_23473,N_23438);
nor U24599 (N_24599,N_23468,N_23921);
nor U24600 (N_24600,N_24266,N_24554);
nor U24601 (N_24601,N_24041,N_24337);
nor U24602 (N_24602,N_24191,N_24067);
nand U24603 (N_24603,N_24079,N_24034);
xnor U24604 (N_24604,N_24003,N_24358);
and U24605 (N_24605,N_24472,N_24414);
or U24606 (N_24606,N_24298,N_24528);
nand U24607 (N_24607,N_24381,N_24286);
or U24608 (N_24608,N_24170,N_24301);
xnor U24609 (N_24609,N_24408,N_24084);
xnor U24610 (N_24610,N_24299,N_24468);
or U24611 (N_24611,N_24407,N_24123);
and U24612 (N_24612,N_24546,N_24105);
nor U24613 (N_24613,N_24163,N_24184);
or U24614 (N_24614,N_24587,N_24101);
and U24615 (N_24615,N_24194,N_24265);
and U24616 (N_24616,N_24596,N_24553);
nor U24617 (N_24617,N_24389,N_24280);
or U24618 (N_24618,N_24519,N_24518);
nand U24619 (N_24619,N_24134,N_24157);
nor U24620 (N_24620,N_24489,N_24429);
nor U24621 (N_24621,N_24565,N_24169);
nand U24622 (N_24622,N_24181,N_24568);
nand U24623 (N_24623,N_24237,N_24219);
xor U24624 (N_24624,N_24193,N_24108);
xnor U24625 (N_24625,N_24345,N_24051);
and U24626 (N_24626,N_24448,N_24016);
nand U24627 (N_24627,N_24391,N_24413);
nand U24628 (N_24628,N_24200,N_24333);
and U24629 (N_24629,N_24271,N_24483);
and U24630 (N_24630,N_24324,N_24251);
and U24631 (N_24631,N_24201,N_24461);
nor U24632 (N_24632,N_24007,N_24015);
nor U24633 (N_24633,N_24187,N_24115);
or U24634 (N_24634,N_24186,N_24061);
or U24635 (N_24635,N_24427,N_24372);
and U24636 (N_24636,N_24014,N_24527);
or U24637 (N_24637,N_24475,N_24444);
and U24638 (N_24638,N_24539,N_24496);
xor U24639 (N_24639,N_24326,N_24292);
nor U24640 (N_24640,N_24270,N_24420);
nand U24641 (N_24641,N_24070,N_24315);
nand U24642 (N_24642,N_24150,N_24208);
and U24643 (N_24643,N_24428,N_24177);
nor U24644 (N_24644,N_24396,N_24185);
nand U24645 (N_24645,N_24558,N_24154);
and U24646 (N_24646,N_24031,N_24118);
nor U24647 (N_24647,N_24453,N_24144);
and U24648 (N_24648,N_24231,N_24235);
and U24649 (N_24649,N_24090,N_24196);
and U24650 (N_24650,N_24497,N_24121);
or U24651 (N_24651,N_24591,N_24319);
and U24652 (N_24652,N_24164,N_24367);
nor U24653 (N_24653,N_24113,N_24149);
xor U24654 (N_24654,N_24541,N_24452);
nand U24655 (N_24655,N_24279,N_24143);
and U24656 (N_24656,N_24024,N_24523);
and U24657 (N_24657,N_24435,N_24330);
or U24658 (N_24658,N_24290,N_24147);
xor U24659 (N_24659,N_24403,N_24455);
and U24660 (N_24660,N_24569,N_24387);
or U24661 (N_24661,N_24006,N_24543);
and U24662 (N_24662,N_24487,N_24263);
xnor U24663 (N_24663,N_24348,N_24599);
or U24664 (N_24664,N_24027,N_24042);
nor U24665 (N_24665,N_24556,N_24465);
xnor U24666 (N_24666,N_24514,N_24437);
and U24667 (N_24667,N_24040,N_24313);
nor U24668 (N_24668,N_24431,N_24555);
nand U24669 (N_24669,N_24028,N_24230);
nand U24670 (N_24670,N_24321,N_24269);
or U24671 (N_24671,N_24512,N_24272);
and U24672 (N_24672,N_24233,N_24060);
or U24673 (N_24673,N_24171,N_24240);
and U24674 (N_24674,N_24103,N_24495);
or U24675 (N_24675,N_24498,N_24480);
and U24676 (N_24676,N_24305,N_24393);
nor U24677 (N_24677,N_24352,N_24579);
nand U24678 (N_24678,N_24582,N_24140);
or U24679 (N_24679,N_24559,N_24173);
or U24680 (N_24680,N_24493,N_24283);
nand U24681 (N_24681,N_24394,N_24013);
nor U24682 (N_24682,N_24276,N_24373);
nand U24683 (N_24683,N_24309,N_24092);
xor U24684 (N_24684,N_24530,N_24334);
and U24685 (N_24685,N_24471,N_24343);
nand U24686 (N_24686,N_24259,N_24162);
nand U24687 (N_24687,N_24397,N_24088);
nand U24688 (N_24688,N_24360,N_24368);
or U24689 (N_24689,N_24202,N_24390);
nor U24690 (N_24690,N_24277,N_24404);
and U24691 (N_24691,N_24438,N_24083);
xor U24692 (N_24692,N_24106,N_24222);
nor U24693 (N_24693,N_24048,N_24111);
and U24694 (N_24694,N_24398,N_24338);
and U24695 (N_24695,N_24211,N_24241);
and U24696 (N_24696,N_24535,N_24047);
and U24697 (N_24697,N_24578,N_24310);
nor U24698 (N_24698,N_24346,N_24341);
or U24699 (N_24699,N_24257,N_24043);
or U24700 (N_24700,N_24570,N_24126);
or U24701 (N_24701,N_24087,N_24536);
nand U24702 (N_24702,N_24250,N_24490);
nand U24703 (N_24703,N_24418,N_24306);
nor U24704 (N_24704,N_24089,N_24593);
or U24705 (N_24705,N_24562,N_24260);
nand U24706 (N_24706,N_24076,N_24441);
nor U24707 (N_24707,N_24145,N_24449);
nor U24708 (N_24708,N_24316,N_24405);
xnor U24709 (N_24709,N_24561,N_24255);
nor U24710 (N_24710,N_24017,N_24062);
or U24711 (N_24711,N_24248,N_24294);
nor U24712 (N_24712,N_24133,N_24500);
nor U24713 (N_24713,N_24071,N_24095);
nand U24714 (N_24714,N_24479,N_24585);
or U24715 (N_24715,N_24226,N_24592);
nor U24716 (N_24716,N_24151,N_24029);
or U24717 (N_24717,N_24597,N_24058);
or U24718 (N_24718,N_24085,N_24586);
or U24719 (N_24719,N_24188,N_24399);
and U24720 (N_24720,N_24142,N_24424);
and U24721 (N_24721,N_24363,N_24366);
nand U24722 (N_24722,N_24550,N_24533);
and U24723 (N_24723,N_24478,N_24351);
and U24724 (N_24724,N_24100,N_24353);
nor U24725 (N_24725,N_24529,N_24349);
nand U24726 (N_24726,N_24544,N_24331);
nor U24727 (N_24727,N_24332,N_24386);
nor U24728 (N_24728,N_24462,N_24112);
xor U24729 (N_24729,N_24282,N_24234);
or U24730 (N_24730,N_24093,N_24510);
xor U24731 (N_24731,N_24409,N_24155);
xnor U24732 (N_24732,N_24137,N_24267);
xor U24733 (N_24733,N_24127,N_24156);
nor U24734 (N_24734,N_24488,N_24012);
and U24735 (N_24735,N_24339,N_24476);
nand U24736 (N_24736,N_24295,N_24022);
nand U24737 (N_24737,N_24246,N_24551);
and U24738 (N_24738,N_24590,N_24074);
nand U24739 (N_24739,N_24576,N_24454);
or U24740 (N_24740,N_24581,N_24102);
nor U24741 (N_24741,N_24521,N_24412);
xnor U24742 (N_24742,N_24508,N_24355);
nand U24743 (N_24743,N_24384,N_24362);
or U24744 (N_24744,N_24046,N_24274);
and U24745 (N_24745,N_24470,N_24442);
nand U24746 (N_24746,N_24460,N_24538);
nor U24747 (N_24747,N_24050,N_24011);
and U24748 (N_24748,N_24481,N_24008);
and U24749 (N_24749,N_24244,N_24039);
and U24750 (N_24750,N_24467,N_24161);
nand U24751 (N_24751,N_24209,N_24053);
xor U24752 (N_24752,N_24261,N_24411);
nand U24753 (N_24753,N_24018,N_24369);
xor U24754 (N_24754,N_24594,N_24165);
or U24755 (N_24755,N_24374,N_24342);
nand U24756 (N_24756,N_24192,N_24128);
nor U24757 (N_24757,N_24542,N_24421);
nand U24758 (N_24758,N_24433,N_24588);
or U24759 (N_24759,N_24117,N_24549);
nand U24760 (N_24760,N_24078,N_24371);
nor U24761 (N_24761,N_24002,N_24522);
and U24762 (N_24762,N_24253,N_24439);
nand U24763 (N_24763,N_24347,N_24158);
nor U24764 (N_24764,N_24504,N_24395);
nand U24765 (N_24765,N_24328,N_24059);
and U24766 (N_24766,N_24056,N_24135);
or U24767 (N_24767,N_24232,N_24213);
nand U24768 (N_24768,N_24236,N_24167);
and U24769 (N_24769,N_24318,N_24010);
nor U24770 (N_24770,N_24036,N_24216);
xnor U24771 (N_24771,N_24447,N_24136);
and U24772 (N_24772,N_24224,N_24443);
or U24773 (N_24773,N_24254,N_24350);
nor U24774 (N_24774,N_24598,N_24515);
nor U24775 (N_24775,N_24107,N_24206);
or U24776 (N_24776,N_24491,N_24289);
nand U24777 (N_24777,N_24320,N_24297);
and U24778 (N_24778,N_24375,N_24300);
or U24779 (N_24779,N_24327,N_24466);
or U24780 (N_24780,N_24264,N_24178);
nand U24781 (N_24781,N_24073,N_24198);
and U24782 (N_24782,N_24473,N_24425);
or U24783 (N_24783,N_24445,N_24189);
or U24784 (N_24784,N_24220,N_24066);
xor U24785 (N_24785,N_24218,N_24068);
nor U24786 (N_24786,N_24458,N_24000);
nand U24787 (N_24787,N_24037,N_24552);
nand U24788 (N_24788,N_24122,N_24560);
xnor U24789 (N_24789,N_24492,N_24456);
nand U24790 (N_24790,N_24446,N_24019);
or U24791 (N_24791,N_24580,N_24055);
nand U24792 (N_24792,N_24168,N_24451);
and U24793 (N_24793,N_24459,N_24436);
nand U24794 (N_24794,N_24025,N_24104);
and U24795 (N_24795,N_24214,N_24566);
and U24796 (N_24796,N_24422,N_24584);
nor U24797 (N_24797,N_24091,N_24457);
or U24798 (N_24798,N_24575,N_24540);
and U24799 (N_24799,N_24082,N_24287);
xor U24800 (N_24800,N_24365,N_24534);
or U24801 (N_24801,N_24573,N_24440);
or U24802 (N_24802,N_24146,N_24335);
xnor U24803 (N_24803,N_24172,N_24505);
nand U24804 (N_24804,N_24314,N_24020);
nand U24805 (N_24805,N_24217,N_24243);
and U24806 (N_24806,N_24033,N_24098);
and U24807 (N_24807,N_24506,N_24406);
and U24808 (N_24808,N_24049,N_24524);
nand U24809 (N_24809,N_24469,N_24494);
xnor U24810 (N_24810,N_24148,N_24129);
nand U24811 (N_24811,N_24038,N_24563);
or U24812 (N_24812,N_24160,N_24474);
or U24813 (N_24813,N_24400,N_24197);
xor U24814 (N_24814,N_24052,N_24380);
xnor U24815 (N_24815,N_24205,N_24419);
xor U24816 (N_24816,N_24225,N_24388);
nor U24817 (N_24817,N_24005,N_24531);
and U24818 (N_24818,N_24284,N_24159);
or U24819 (N_24819,N_24166,N_24340);
nand U24820 (N_24820,N_24401,N_24153);
or U24821 (N_24821,N_24141,N_24081);
nand U24822 (N_24822,N_24080,N_24545);
nand U24823 (N_24823,N_24293,N_24557);
and U24824 (N_24824,N_24110,N_24238);
or U24825 (N_24825,N_24572,N_24450);
or U24826 (N_24826,N_24434,N_24072);
xor U24827 (N_24827,N_24589,N_24507);
and U24828 (N_24828,N_24262,N_24215);
or U24829 (N_24829,N_24207,N_24138);
nor U24830 (N_24830,N_24464,N_24595);
or U24831 (N_24831,N_24120,N_24004);
nor U24832 (N_24832,N_24247,N_24516);
and U24833 (N_24833,N_24376,N_24275);
nand U24834 (N_24834,N_24245,N_24385);
nand U24835 (N_24835,N_24482,N_24329);
or U24836 (N_24836,N_24182,N_24021);
nand U24837 (N_24837,N_24520,N_24484);
or U24838 (N_24838,N_24063,N_24526);
nand U24839 (N_24839,N_24203,N_24502);
nand U24840 (N_24840,N_24547,N_24370);
xnor U24841 (N_24841,N_24116,N_24139);
nand U24842 (N_24842,N_24190,N_24023);
nand U24843 (N_24843,N_24291,N_24288);
or U24844 (N_24844,N_24307,N_24513);
nor U24845 (N_24845,N_24035,N_24285);
or U24846 (N_24846,N_24077,N_24410);
and U24847 (N_24847,N_24125,N_24183);
and U24848 (N_24848,N_24097,N_24179);
or U24849 (N_24849,N_24322,N_24009);
nor U24850 (N_24850,N_24030,N_24571);
nand U24851 (N_24851,N_24308,N_24477);
nor U24852 (N_24852,N_24426,N_24383);
xor U24853 (N_24853,N_24278,N_24537);
xor U24854 (N_24854,N_24336,N_24296);
nand U24855 (N_24855,N_24130,N_24174);
nor U24856 (N_24856,N_24548,N_24054);
xnor U24857 (N_24857,N_24415,N_24044);
nor U24858 (N_24858,N_24281,N_24486);
xnor U24859 (N_24859,N_24199,N_24354);
or U24860 (N_24860,N_24119,N_24302);
xnor U24861 (N_24861,N_24176,N_24463);
xor U24862 (N_24862,N_24430,N_24499);
nor U24863 (N_24863,N_24323,N_24432);
nand U24864 (N_24864,N_24382,N_24525);
or U24865 (N_24865,N_24228,N_24256);
xnor U24866 (N_24866,N_24364,N_24511);
xnor U24867 (N_24867,N_24221,N_24075);
nand U24868 (N_24868,N_24096,N_24045);
and U24869 (N_24869,N_24032,N_24239);
nor U24870 (N_24870,N_24212,N_24423);
and U24871 (N_24871,N_24574,N_24359);
and U24872 (N_24872,N_24273,N_24583);
nor U24873 (N_24873,N_24064,N_24099);
nor U24874 (N_24874,N_24258,N_24311);
xnor U24875 (N_24875,N_24210,N_24249);
or U24876 (N_24876,N_24325,N_24001);
xor U24877 (N_24877,N_24057,N_24356);
and U24878 (N_24878,N_24361,N_24564);
or U24879 (N_24879,N_24252,N_24303);
nand U24880 (N_24880,N_24417,N_24065);
nand U24881 (N_24881,N_24195,N_24131);
xnor U24882 (N_24882,N_24485,N_24567);
or U24883 (N_24883,N_24124,N_24069);
nand U24884 (N_24884,N_24204,N_24094);
xor U24885 (N_24885,N_24509,N_24268);
nand U24886 (N_24886,N_24114,N_24517);
or U24887 (N_24887,N_24180,N_24577);
and U24888 (N_24888,N_24086,N_24109);
nor U24889 (N_24889,N_24304,N_24501);
or U24890 (N_24890,N_24402,N_24312);
or U24891 (N_24891,N_24229,N_24175);
nor U24892 (N_24892,N_24132,N_24223);
or U24893 (N_24893,N_24378,N_24242);
xor U24894 (N_24894,N_24227,N_24532);
nand U24895 (N_24895,N_24379,N_24377);
or U24896 (N_24896,N_24317,N_24344);
xnor U24897 (N_24897,N_24357,N_24392);
nand U24898 (N_24898,N_24026,N_24416);
xor U24899 (N_24899,N_24152,N_24503);
and U24900 (N_24900,N_24283,N_24242);
xor U24901 (N_24901,N_24375,N_24554);
nand U24902 (N_24902,N_24035,N_24151);
and U24903 (N_24903,N_24412,N_24187);
or U24904 (N_24904,N_24165,N_24589);
or U24905 (N_24905,N_24573,N_24304);
nor U24906 (N_24906,N_24168,N_24145);
and U24907 (N_24907,N_24194,N_24584);
xnor U24908 (N_24908,N_24424,N_24186);
or U24909 (N_24909,N_24547,N_24218);
nand U24910 (N_24910,N_24484,N_24527);
or U24911 (N_24911,N_24399,N_24314);
nor U24912 (N_24912,N_24103,N_24524);
xnor U24913 (N_24913,N_24091,N_24024);
or U24914 (N_24914,N_24480,N_24223);
and U24915 (N_24915,N_24563,N_24128);
or U24916 (N_24916,N_24209,N_24355);
and U24917 (N_24917,N_24038,N_24170);
or U24918 (N_24918,N_24565,N_24339);
and U24919 (N_24919,N_24024,N_24033);
nand U24920 (N_24920,N_24473,N_24073);
xnor U24921 (N_24921,N_24199,N_24493);
or U24922 (N_24922,N_24094,N_24552);
or U24923 (N_24923,N_24426,N_24287);
nand U24924 (N_24924,N_24231,N_24119);
nor U24925 (N_24925,N_24543,N_24104);
or U24926 (N_24926,N_24372,N_24373);
xor U24927 (N_24927,N_24111,N_24267);
nand U24928 (N_24928,N_24418,N_24428);
nand U24929 (N_24929,N_24520,N_24202);
or U24930 (N_24930,N_24276,N_24423);
nand U24931 (N_24931,N_24333,N_24168);
nand U24932 (N_24932,N_24050,N_24136);
nor U24933 (N_24933,N_24390,N_24510);
xnor U24934 (N_24934,N_24397,N_24531);
and U24935 (N_24935,N_24575,N_24339);
nor U24936 (N_24936,N_24390,N_24349);
nor U24937 (N_24937,N_24195,N_24434);
nand U24938 (N_24938,N_24598,N_24062);
xnor U24939 (N_24939,N_24487,N_24450);
nor U24940 (N_24940,N_24332,N_24231);
and U24941 (N_24941,N_24229,N_24323);
or U24942 (N_24942,N_24373,N_24486);
and U24943 (N_24943,N_24470,N_24207);
nand U24944 (N_24944,N_24585,N_24554);
xnor U24945 (N_24945,N_24380,N_24342);
xor U24946 (N_24946,N_24198,N_24425);
or U24947 (N_24947,N_24417,N_24329);
xor U24948 (N_24948,N_24497,N_24219);
or U24949 (N_24949,N_24451,N_24425);
nand U24950 (N_24950,N_24037,N_24545);
and U24951 (N_24951,N_24080,N_24308);
or U24952 (N_24952,N_24573,N_24550);
and U24953 (N_24953,N_24296,N_24335);
nand U24954 (N_24954,N_24322,N_24223);
xor U24955 (N_24955,N_24303,N_24132);
xor U24956 (N_24956,N_24561,N_24593);
xnor U24957 (N_24957,N_24011,N_24238);
or U24958 (N_24958,N_24276,N_24195);
xnor U24959 (N_24959,N_24079,N_24481);
and U24960 (N_24960,N_24085,N_24338);
nor U24961 (N_24961,N_24531,N_24568);
xnor U24962 (N_24962,N_24115,N_24379);
or U24963 (N_24963,N_24315,N_24472);
and U24964 (N_24964,N_24546,N_24351);
nand U24965 (N_24965,N_24189,N_24002);
xor U24966 (N_24966,N_24463,N_24349);
nand U24967 (N_24967,N_24119,N_24441);
or U24968 (N_24968,N_24096,N_24537);
and U24969 (N_24969,N_24110,N_24547);
xor U24970 (N_24970,N_24302,N_24107);
nand U24971 (N_24971,N_24407,N_24432);
or U24972 (N_24972,N_24542,N_24534);
and U24973 (N_24973,N_24201,N_24314);
xnor U24974 (N_24974,N_24438,N_24565);
or U24975 (N_24975,N_24087,N_24301);
and U24976 (N_24976,N_24494,N_24331);
and U24977 (N_24977,N_24119,N_24174);
and U24978 (N_24978,N_24343,N_24208);
nand U24979 (N_24979,N_24542,N_24226);
or U24980 (N_24980,N_24255,N_24060);
xor U24981 (N_24981,N_24129,N_24305);
nand U24982 (N_24982,N_24357,N_24295);
nor U24983 (N_24983,N_24495,N_24385);
nand U24984 (N_24984,N_24385,N_24339);
or U24985 (N_24985,N_24354,N_24506);
nor U24986 (N_24986,N_24573,N_24125);
nor U24987 (N_24987,N_24041,N_24344);
xor U24988 (N_24988,N_24368,N_24269);
or U24989 (N_24989,N_24490,N_24089);
xor U24990 (N_24990,N_24217,N_24213);
or U24991 (N_24991,N_24574,N_24266);
and U24992 (N_24992,N_24566,N_24476);
and U24993 (N_24993,N_24235,N_24138);
nor U24994 (N_24994,N_24052,N_24506);
or U24995 (N_24995,N_24055,N_24226);
and U24996 (N_24996,N_24503,N_24468);
or U24997 (N_24997,N_24344,N_24334);
xnor U24998 (N_24998,N_24387,N_24374);
nor U24999 (N_24999,N_24371,N_24225);
and U25000 (N_25000,N_24197,N_24373);
nand U25001 (N_25001,N_24519,N_24145);
or U25002 (N_25002,N_24165,N_24392);
or U25003 (N_25003,N_24145,N_24408);
or U25004 (N_25004,N_24024,N_24346);
nor U25005 (N_25005,N_24306,N_24127);
or U25006 (N_25006,N_24035,N_24484);
and U25007 (N_25007,N_24524,N_24257);
xor U25008 (N_25008,N_24066,N_24251);
nor U25009 (N_25009,N_24210,N_24116);
nor U25010 (N_25010,N_24525,N_24515);
or U25011 (N_25011,N_24317,N_24134);
and U25012 (N_25012,N_24079,N_24433);
xor U25013 (N_25013,N_24089,N_24206);
or U25014 (N_25014,N_24579,N_24325);
xor U25015 (N_25015,N_24288,N_24575);
and U25016 (N_25016,N_24347,N_24517);
nor U25017 (N_25017,N_24585,N_24113);
nor U25018 (N_25018,N_24340,N_24463);
or U25019 (N_25019,N_24416,N_24071);
nand U25020 (N_25020,N_24370,N_24056);
or U25021 (N_25021,N_24001,N_24077);
and U25022 (N_25022,N_24581,N_24509);
xnor U25023 (N_25023,N_24161,N_24529);
nor U25024 (N_25024,N_24463,N_24450);
nand U25025 (N_25025,N_24205,N_24041);
nand U25026 (N_25026,N_24325,N_24258);
nor U25027 (N_25027,N_24247,N_24483);
nand U25028 (N_25028,N_24255,N_24357);
nand U25029 (N_25029,N_24340,N_24338);
xor U25030 (N_25030,N_24552,N_24522);
xor U25031 (N_25031,N_24262,N_24063);
and U25032 (N_25032,N_24493,N_24033);
nor U25033 (N_25033,N_24072,N_24402);
nand U25034 (N_25034,N_24377,N_24134);
xnor U25035 (N_25035,N_24502,N_24019);
or U25036 (N_25036,N_24522,N_24105);
nand U25037 (N_25037,N_24536,N_24224);
nand U25038 (N_25038,N_24340,N_24369);
and U25039 (N_25039,N_24102,N_24049);
nor U25040 (N_25040,N_24071,N_24339);
and U25041 (N_25041,N_24523,N_24199);
and U25042 (N_25042,N_24431,N_24387);
nor U25043 (N_25043,N_24156,N_24417);
and U25044 (N_25044,N_24215,N_24538);
nand U25045 (N_25045,N_24313,N_24582);
nand U25046 (N_25046,N_24211,N_24175);
nand U25047 (N_25047,N_24370,N_24010);
nand U25048 (N_25048,N_24146,N_24126);
xnor U25049 (N_25049,N_24134,N_24473);
nor U25050 (N_25050,N_24417,N_24224);
xor U25051 (N_25051,N_24004,N_24028);
nor U25052 (N_25052,N_24199,N_24564);
nand U25053 (N_25053,N_24552,N_24223);
xor U25054 (N_25054,N_24021,N_24070);
xor U25055 (N_25055,N_24554,N_24125);
nand U25056 (N_25056,N_24025,N_24008);
or U25057 (N_25057,N_24373,N_24344);
xnor U25058 (N_25058,N_24187,N_24398);
and U25059 (N_25059,N_24533,N_24333);
and U25060 (N_25060,N_24130,N_24542);
or U25061 (N_25061,N_24298,N_24410);
xor U25062 (N_25062,N_24359,N_24554);
xnor U25063 (N_25063,N_24310,N_24195);
xnor U25064 (N_25064,N_24295,N_24434);
and U25065 (N_25065,N_24022,N_24558);
nand U25066 (N_25066,N_24243,N_24137);
xor U25067 (N_25067,N_24547,N_24571);
or U25068 (N_25068,N_24517,N_24575);
or U25069 (N_25069,N_24577,N_24375);
or U25070 (N_25070,N_24478,N_24363);
and U25071 (N_25071,N_24556,N_24213);
nand U25072 (N_25072,N_24265,N_24174);
nor U25073 (N_25073,N_24186,N_24201);
nor U25074 (N_25074,N_24075,N_24465);
or U25075 (N_25075,N_24332,N_24398);
nand U25076 (N_25076,N_24059,N_24178);
xor U25077 (N_25077,N_24431,N_24195);
xor U25078 (N_25078,N_24507,N_24320);
and U25079 (N_25079,N_24023,N_24337);
and U25080 (N_25080,N_24233,N_24208);
xor U25081 (N_25081,N_24070,N_24411);
and U25082 (N_25082,N_24366,N_24044);
nor U25083 (N_25083,N_24210,N_24422);
nand U25084 (N_25084,N_24464,N_24072);
and U25085 (N_25085,N_24214,N_24302);
nor U25086 (N_25086,N_24300,N_24380);
nand U25087 (N_25087,N_24431,N_24108);
or U25088 (N_25088,N_24016,N_24469);
nor U25089 (N_25089,N_24143,N_24368);
nand U25090 (N_25090,N_24065,N_24469);
and U25091 (N_25091,N_24300,N_24225);
xnor U25092 (N_25092,N_24399,N_24233);
or U25093 (N_25093,N_24181,N_24029);
nand U25094 (N_25094,N_24395,N_24439);
xor U25095 (N_25095,N_24144,N_24437);
nor U25096 (N_25096,N_24345,N_24187);
and U25097 (N_25097,N_24070,N_24359);
xnor U25098 (N_25098,N_24255,N_24103);
nor U25099 (N_25099,N_24254,N_24487);
xnor U25100 (N_25100,N_24431,N_24441);
nand U25101 (N_25101,N_24556,N_24153);
nand U25102 (N_25102,N_24366,N_24041);
nor U25103 (N_25103,N_24179,N_24452);
nand U25104 (N_25104,N_24058,N_24261);
xor U25105 (N_25105,N_24274,N_24155);
or U25106 (N_25106,N_24208,N_24561);
and U25107 (N_25107,N_24340,N_24064);
nor U25108 (N_25108,N_24383,N_24022);
and U25109 (N_25109,N_24157,N_24103);
xnor U25110 (N_25110,N_24444,N_24203);
xnor U25111 (N_25111,N_24239,N_24392);
nor U25112 (N_25112,N_24072,N_24107);
nor U25113 (N_25113,N_24369,N_24327);
and U25114 (N_25114,N_24347,N_24257);
xor U25115 (N_25115,N_24202,N_24156);
xor U25116 (N_25116,N_24040,N_24414);
xnor U25117 (N_25117,N_24382,N_24017);
xor U25118 (N_25118,N_24129,N_24543);
nand U25119 (N_25119,N_24343,N_24083);
xnor U25120 (N_25120,N_24323,N_24403);
nor U25121 (N_25121,N_24580,N_24321);
xnor U25122 (N_25122,N_24568,N_24528);
or U25123 (N_25123,N_24228,N_24110);
or U25124 (N_25124,N_24291,N_24061);
nor U25125 (N_25125,N_24263,N_24474);
nor U25126 (N_25126,N_24224,N_24033);
and U25127 (N_25127,N_24400,N_24095);
nand U25128 (N_25128,N_24022,N_24097);
nor U25129 (N_25129,N_24228,N_24470);
and U25130 (N_25130,N_24134,N_24131);
xor U25131 (N_25131,N_24129,N_24252);
or U25132 (N_25132,N_24428,N_24116);
or U25133 (N_25133,N_24144,N_24455);
nand U25134 (N_25134,N_24096,N_24031);
and U25135 (N_25135,N_24591,N_24239);
nor U25136 (N_25136,N_24591,N_24143);
nand U25137 (N_25137,N_24175,N_24486);
xor U25138 (N_25138,N_24554,N_24485);
or U25139 (N_25139,N_24164,N_24477);
or U25140 (N_25140,N_24333,N_24588);
xor U25141 (N_25141,N_24497,N_24365);
or U25142 (N_25142,N_24151,N_24373);
and U25143 (N_25143,N_24290,N_24203);
nor U25144 (N_25144,N_24024,N_24400);
nor U25145 (N_25145,N_24093,N_24123);
xor U25146 (N_25146,N_24373,N_24448);
or U25147 (N_25147,N_24411,N_24317);
xor U25148 (N_25148,N_24121,N_24492);
nor U25149 (N_25149,N_24273,N_24346);
xnor U25150 (N_25150,N_24480,N_24027);
or U25151 (N_25151,N_24560,N_24087);
xnor U25152 (N_25152,N_24334,N_24314);
xor U25153 (N_25153,N_24101,N_24449);
xnor U25154 (N_25154,N_24411,N_24500);
and U25155 (N_25155,N_24591,N_24526);
xor U25156 (N_25156,N_24338,N_24027);
nand U25157 (N_25157,N_24424,N_24383);
xnor U25158 (N_25158,N_24179,N_24456);
and U25159 (N_25159,N_24303,N_24466);
and U25160 (N_25160,N_24237,N_24548);
or U25161 (N_25161,N_24265,N_24497);
nand U25162 (N_25162,N_24409,N_24090);
nand U25163 (N_25163,N_24467,N_24466);
xor U25164 (N_25164,N_24563,N_24183);
nor U25165 (N_25165,N_24561,N_24250);
or U25166 (N_25166,N_24304,N_24381);
or U25167 (N_25167,N_24118,N_24262);
xor U25168 (N_25168,N_24559,N_24511);
nand U25169 (N_25169,N_24507,N_24063);
nor U25170 (N_25170,N_24571,N_24302);
or U25171 (N_25171,N_24494,N_24308);
xor U25172 (N_25172,N_24491,N_24498);
xor U25173 (N_25173,N_24537,N_24473);
or U25174 (N_25174,N_24262,N_24319);
or U25175 (N_25175,N_24400,N_24440);
nor U25176 (N_25176,N_24235,N_24397);
nor U25177 (N_25177,N_24179,N_24430);
xor U25178 (N_25178,N_24089,N_24398);
nand U25179 (N_25179,N_24053,N_24591);
and U25180 (N_25180,N_24153,N_24307);
nor U25181 (N_25181,N_24049,N_24075);
and U25182 (N_25182,N_24382,N_24136);
or U25183 (N_25183,N_24484,N_24055);
nor U25184 (N_25184,N_24199,N_24063);
and U25185 (N_25185,N_24340,N_24356);
xor U25186 (N_25186,N_24003,N_24550);
nor U25187 (N_25187,N_24241,N_24171);
xnor U25188 (N_25188,N_24544,N_24333);
nand U25189 (N_25189,N_24215,N_24119);
xor U25190 (N_25190,N_24498,N_24252);
xor U25191 (N_25191,N_24382,N_24537);
or U25192 (N_25192,N_24138,N_24335);
xor U25193 (N_25193,N_24131,N_24106);
or U25194 (N_25194,N_24036,N_24590);
nand U25195 (N_25195,N_24586,N_24469);
and U25196 (N_25196,N_24026,N_24436);
nor U25197 (N_25197,N_24366,N_24167);
or U25198 (N_25198,N_24417,N_24112);
or U25199 (N_25199,N_24517,N_24195);
or U25200 (N_25200,N_24880,N_24785);
or U25201 (N_25201,N_24713,N_25190);
and U25202 (N_25202,N_24951,N_25150);
nand U25203 (N_25203,N_24729,N_24975);
xor U25204 (N_25204,N_24775,N_24631);
nand U25205 (N_25205,N_24963,N_24640);
nor U25206 (N_25206,N_24994,N_24978);
nor U25207 (N_25207,N_24600,N_25107);
or U25208 (N_25208,N_25096,N_24678);
or U25209 (N_25209,N_24894,N_25126);
or U25210 (N_25210,N_24816,N_24998);
and U25211 (N_25211,N_24666,N_25199);
nand U25212 (N_25212,N_24723,N_25066);
nand U25213 (N_25213,N_24934,N_24956);
and U25214 (N_25214,N_25075,N_24626);
or U25215 (N_25215,N_24703,N_25164);
nor U25216 (N_25216,N_25191,N_24862);
or U25217 (N_25217,N_25026,N_24759);
xnor U25218 (N_25218,N_24728,N_25175);
nor U25219 (N_25219,N_24846,N_25024);
nor U25220 (N_25220,N_24909,N_24753);
nand U25221 (N_25221,N_25056,N_25020);
nor U25222 (N_25222,N_25114,N_24930);
xor U25223 (N_25223,N_25122,N_24700);
xor U25224 (N_25224,N_25072,N_24986);
xnor U25225 (N_25225,N_24739,N_24848);
xnor U25226 (N_25226,N_24830,N_25166);
nand U25227 (N_25227,N_25161,N_24622);
xnor U25228 (N_25228,N_24896,N_24853);
xnor U25229 (N_25229,N_25111,N_24709);
nand U25230 (N_25230,N_24945,N_24714);
nand U25231 (N_25231,N_25094,N_24991);
and U25232 (N_25232,N_24919,N_24607);
nor U25233 (N_25233,N_24800,N_25037);
nand U25234 (N_25234,N_24958,N_24618);
nand U25235 (N_25235,N_24653,N_24855);
nor U25236 (N_25236,N_24736,N_25062);
nand U25237 (N_25237,N_24903,N_24658);
nand U25238 (N_25238,N_25130,N_24886);
xnor U25239 (N_25239,N_24645,N_24946);
nor U25240 (N_25240,N_24665,N_25137);
or U25241 (N_25241,N_24677,N_25148);
xnor U25242 (N_25242,N_24927,N_24811);
and U25243 (N_25243,N_24773,N_25180);
nor U25244 (N_25244,N_24711,N_24831);
nor U25245 (N_25245,N_24905,N_24720);
nand U25246 (N_25246,N_24871,N_24791);
or U25247 (N_25247,N_25140,N_24808);
nand U25248 (N_25248,N_25116,N_25165);
nand U25249 (N_25249,N_24629,N_25045);
xnor U25250 (N_25250,N_24997,N_24619);
nand U25251 (N_25251,N_25173,N_24803);
nand U25252 (N_25252,N_24628,N_24688);
or U25253 (N_25253,N_24922,N_24962);
or U25254 (N_25254,N_25077,N_24699);
or U25255 (N_25255,N_25174,N_24790);
nor U25256 (N_25256,N_24959,N_25055);
nor U25257 (N_25257,N_25101,N_24877);
nand U25258 (N_25258,N_25134,N_24737);
xnor U25259 (N_25259,N_24606,N_25186);
nand U25260 (N_25260,N_24719,N_24957);
nor U25261 (N_25261,N_25038,N_24879);
or U25262 (N_25262,N_24671,N_24679);
and U25263 (N_25263,N_24863,N_25043);
nor U25264 (N_25264,N_25001,N_24970);
and U25265 (N_25265,N_24837,N_24797);
nand U25266 (N_25266,N_25095,N_24832);
or U25267 (N_25267,N_25171,N_25083);
or U25268 (N_25268,N_24721,N_24984);
and U25269 (N_25269,N_25081,N_25048);
nand U25270 (N_25270,N_24647,N_24814);
nor U25271 (N_25271,N_24899,N_24869);
nand U25272 (N_25272,N_24710,N_25103);
nand U25273 (N_25273,N_25160,N_24870);
nand U25274 (N_25274,N_24605,N_25109);
nor U25275 (N_25275,N_24952,N_24937);
nor U25276 (N_25276,N_25181,N_24972);
or U25277 (N_25277,N_24692,N_24732);
or U25278 (N_25278,N_24741,N_24602);
and U25279 (N_25279,N_25000,N_24722);
nand U25280 (N_25280,N_24954,N_25155);
nor U25281 (N_25281,N_24988,N_25098);
nand U25282 (N_25282,N_24992,N_25035);
and U25283 (N_25283,N_24941,N_25058);
nand U25284 (N_25284,N_25074,N_24915);
xnor U25285 (N_25285,N_24778,N_25105);
nor U25286 (N_25286,N_24769,N_24825);
xnor U25287 (N_25287,N_25082,N_24616);
and U25288 (N_25288,N_24743,N_25011);
xnor U25289 (N_25289,N_24895,N_25071);
xnor U25290 (N_25290,N_24891,N_24780);
and U25291 (N_25291,N_25015,N_24921);
and U25292 (N_25292,N_24772,N_25167);
nand U25293 (N_25293,N_24718,N_24652);
and U25294 (N_25294,N_24748,N_24768);
xnor U25295 (N_25295,N_24627,N_25127);
and U25296 (N_25296,N_24795,N_24980);
nor U25297 (N_25297,N_24751,N_24900);
nand U25298 (N_25298,N_24784,N_24985);
or U25299 (N_25299,N_25016,N_24668);
nand U25300 (N_25300,N_24839,N_25121);
nand U25301 (N_25301,N_24644,N_24686);
xor U25302 (N_25302,N_24684,N_24966);
or U25303 (N_25303,N_24939,N_24872);
and U25304 (N_25304,N_24757,N_24824);
or U25305 (N_25305,N_25002,N_25009);
or U25306 (N_25306,N_24804,N_25034);
xor U25307 (N_25307,N_25070,N_24614);
nand U25308 (N_25308,N_25168,N_25032);
xnor U25309 (N_25309,N_24819,N_25040);
xnor U25310 (N_25310,N_25143,N_25136);
and U25311 (N_25311,N_25019,N_24885);
or U25312 (N_25312,N_25133,N_24747);
and U25313 (N_25313,N_24641,N_24866);
and U25314 (N_25314,N_24776,N_24989);
nand U25315 (N_25315,N_24760,N_24620);
or U25316 (N_25316,N_24664,N_24977);
nor U25317 (N_25317,N_24655,N_24925);
nor U25318 (N_25318,N_24648,N_24758);
and U25319 (N_25319,N_24706,N_24812);
nor U25320 (N_25320,N_24782,N_25087);
or U25321 (N_25321,N_25146,N_24821);
or U25322 (N_25322,N_25147,N_25142);
nor U25323 (N_25323,N_24673,N_24796);
nor U25324 (N_25324,N_24828,N_25088);
nor U25325 (N_25325,N_24983,N_25196);
xnor U25326 (N_25326,N_25036,N_24923);
nor U25327 (N_25327,N_25198,N_24765);
nor U25328 (N_25328,N_24738,N_24726);
nor U25329 (N_25329,N_25139,N_25172);
nand U25330 (N_25330,N_24623,N_24624);
or U25331 (N_25331,N_24842,N_25120);
and U25332 (N_25332,N_24806,N_24663);
nand U25333 (N_25333,N_24897,N_24702);
or U25334 (N_25334,N_25159,N_24734);
nor U25335 (N_25335,N_25068,N_24854);
xnor U25336 (N_25336,N_24889,N_24874);
or U25337 (N_25337,N_24860,N_24676);
xnor U25338 (N_25338,N_25162,N_25033);
nand U25339 (N_25339,N_24745,N_25086);
nor U25340 (N_25340,N_25017,N_25061);
or U25341 (N_25341,N_24650,N_25169);
xnor U25342 (N_25342,N_24730,N_25102);
xnor U25343 (N_25343,N_25010,N_25118);
and U25344 (N_25344,N_24693,N_24820);
xnor U25345 (N_25345,N_24953,N_24932);
nand U25346 (N_25346,N_24928,N_25065);
and U25347 (N_25347,N_24987,N_24906);
nand U25348 (N_25348,N_24783,N_24960);
xor U25349 (N_25349,N_25123,N_24681);
nor U25350 (N_25350,N_24731,N_24834);
xnor U25351 (N_25351,N_24973,N_24637);
or U25352 (N_25352,N_24868,N_25021);
and U25353 (N_25353,N_24733,N_24704);
or U25354 (N_25354,N_25158,N_25022);
or U25355 (N_25355,N_25135,N_24892);
and U25356 (N_25356,N_25131,N_25063);
xnor U25357 (N_25357,N_25025,N_25193);
nand U25358 (N_25358,N_24969,N_24849);
xnor U25359 (N_25359,N_24770,N_25084);
or U25360 (N_25360,N_24815,N_25047);
xor U25361 (N_25361,N_24764,N_24852);
nor U25362 (N_25362,N_25151,N_24695);
nor U25363 (N_25363,N_24917,N_24636);
or U25364 (N_25364,N_24993,N_24774);
nor U25365 (N_25365,N_24755,N_25046);
nor U25366 (N_25366,N_24883,N_24807);
nor U25367 (N_25367,N_24818,N_24938);
and U25368 (N_25368,N_24944,N_25124);
or U25369 (N_25369,N_25141,N_25092);
nor U25370 (N_25370,N_24982,N_25106);
nor U25371 (N_25371,N_24777,N_24675);
or U25372 (N_25372,N_24792,N_24754);
or U25373 (N_25373,N_24875,N_25197);
nor U25374 (N_25374,N_24904,N_24621);
nor U25375 (N_25375,N_24836,N_25089);
nor U25376 (N_25376,N_24639,N_24810);
or U25377 (N_25377,N_24697,N_24685);
or U25378 (N_25378,N_24793,N_24746);
or U25379 (N_25379,N_24826,N_25179);
nor U25380 (N_25380,N_24612,N_24943);
nand U25381 (N_25381,N_24601,N_25182);
nor U25382 (N_25382,N_25064,N_24916);
nor U25383 (N_25383,N_24630,N_24833);
and U25384 (N_25384,N_24691,N_25187);
xor U25385 (N_25385,N_24799,N_25156);
xor U25386 (N_25386,N_24656,N_24705);
nand U25387 (N_25387,N_24657,N_25079);
xor U25388 (N_25388,N_25041,N_25049);
xor U25389 (N_25389,N_24634,N_25090);
nor U25390 (N_25390,N_24841,N_24786);
nand U25391 (N_25391,N_25195,N_24749);
xnor U25392 (N_25392,N_24838,N_25080);
or U25393 (N_25393,N_24843,N_25053);
nand U25394 (N_25394,N_24756,N_24609);
or U25395 (N_25395,N_25091,N_25144);
nand U25396 (N_25396,N_24981,N_24861);
or U25397 (N_25397,N_24682,N_25117);
nor U25398 (N_25398,N_24873,N_24935);
xnor U25399 (N_25399,N_24781,N_25054);
nor U25400 (N_25400,N_24767,N_25192);
nand U25401 (N_25401,N_24742,N_25113);
nand U25402 (N_25402,N_24926,N_24914);
nor U25403 (N_25403,N_24787,N_24701);
and U25404 (N_25404,N_24893,N_24670);
nand U25405 (N_25405,N_24689,N_24662);
xnor U25406 (N_25406,N_25154,N_24632);
nand U25407 (N_25407,N_24865,N_25078);
and U25408 (N_25408,N_25050,N_25030);
nor U25409 (N_25409,N_25145,N_24835);
or U25410 (N_25410,N_24851,N_25119);
nand U25411 (N_25411,N_24635,N_25051);
or U25412 (N_25412,N_25183,N_24968);
or U25413 (N_25413,N_24822,N_24912);
xnor U25414 (N_25414,N_24603,N_25004);
or U25415 (N_25415,N_24680,N_25153);
xnor U25416 (N_25416,N_24976,N_24876);
nor U25417 (N_25417,N_24687,N_25012);
and U25418 (N_25418,N_25194,N_25044);
or U25419 (N_25419,N_24651,N_24918);
nand U25420 (N_25420,N_24694,N_24887);
nand U25421 (N_25421,N_25129,N_25176);
nor U25422 (N_25422,N_24890,N_24999);
nand U25423 (N_25423,N_24660,N_24990);
xor U25424 (N_25424,N_24613,N_24844);
or U25425 (N_25425,N_24805,N_24744);
nor U25426 (N_25426,N_24610,N_24750);
xnor U25427 (N_25427,N_25112,N_24717);
and U25428 (N_25428,N_24789,N_25073);
and U25429 (N_25429,N_25149,N_24654);
nand U25430 (N_25430,N_24633,N_24642);
nor U25431 (N_25431,N_25067,N_24817);
or U25432 (N_25432,N_24667,N_25029);
nor U25433 (N_25433,N_24942,N_24672);
nand U25434 (N_25434,N_24617,N_24604);
and U25435 (N_25435,N_24995,N_24931);
or U25436 (N_25436,N_24625,N_24878);
or U25437 (N_25437,N_24974,N_25006);
and U25438 (N_25438,N_24725,N_25099);
nand U25439 (N_25439,N_25076,N_25185);
xnor U25440 (N_25440,N_24615,N_25184);
and U25441 (N_25441,N_24809,N_25132);
nand U25442 (N_25442,N_24924,N_24882);
nand U25443 (N_25443,N_25005,N_24898);
nand U25444 (N_25444,N_24936,N_24902);
or U25445 (N_25445,N_24727,N_25039);
nor U25446 (N_25446,N_25028,N_25189);
nand U25447 (N_25447,N_25093,N_24961);
nor U25448 (N_25448,N_24971,N_24850);
and U25449 (N_25449,N_25152,N_24771);
nor U25450 (N_25450,N_24801,N_24696);
nand U25451 (N_25451,N_24901,N_24856);
nand U25452 (N_25452,N_24779,N_25027);
and U25453 (N_25453,N_24683,N_24920);
nand U25454 (N_25454,N_24712,N_24929);
or U25455 (N_25455,N_24823,N_24967);
and U25456 (N_25456,N_24669,N_24661);
nand U25457 (N_25457,N_24798,N_25108);
xnor U25458 (N_25458,N_25008,N_24707);
nand U25459 (N_25459,N_25014,N_24888);
nor U25460 (N_25460,N_24735,N_24761);
nand U25461 (N_25461,N_25115,N_24864);
xnor U25462 (N_25462,N_24867,N_25125);
nor U25463 (N_25463,N_24950,N_25069);
and U25464 (N_25464,N_25188,N_24911);
xor U25465 (N_25465,N_25097,N_24716);
nand U25466 (N_25466,N_25042,N_24740);
and U25467 (N_25467,N_24884,N_24847);
nor U25468 (N_25468,N_24674,N_25128);
or U25469 (N_25469,N_24708,N_25163);
xor U25470 (N_25470,N_25177,N_24788);
nor U25471 (N_25471,N_24643,N_25104);
nor U25472 (N_25472,N_24840,N_24827);
or U25473 (N_25473,N_24940,N_25059);
xnor U25474 (N_25474,N_24845,N_24763);
nand U25475 (N_25475,N_24859,N_25018);
nor U25476 (N_25476,N_24724,N_25170);
and U25477 (N_25477,N_25007,N_24690);
and U25478 (N_25478,N_24802,N_24813);
nor U25479 (N_25479,N_24762,N_25085);
nor U25480 (N_25480,N_25003,N_24933);
xor U25481 (N_25481,N_24948,N_24965);
and U25482 (N_25482,N_24910,N_24955);
nor U25483 (N_25483,N_24766,N_25157);
or U25484 (N_25484,N_25023,N_24964);
nor U25485 (N_25485,N_25057,N_24947);
nand U25486 (N_25486,N_25100,N_25110);
or U25487 (N_25487,N_25138,N_25052);
nor U25488 (N_25488,N_24979,N_24611);
or U25489 (N_25489,N_24881,N_24698);
and U25490 (N_25490,N_24858,N_24715);
nand U25491 (N_25491,N_24908,N_24913);
nor U25492 (N_25492,N_24794,N_24638);
nand U25493 (N_25493,N_24829,N_24996);
or U25494 (N_25494,N_24907,N_24646);
nor U25495 (N_25495,N_24608,N_25031);
nand U25496 (N_25496,N_24857,N_24752);
and U25497 (N_25497,N_24649,N_25178);
nor U25498 (N_25498,N_25060,N_24949);
nand U25499 (N_25499,N_25013,N_24659);
and U25500 (N_25500,N_25074,N_24615);
xnor U25501 (N_25501,N_25185,N_24734);
or U25502 (N_25502,N_24862,N_24765);
xor U25503 (N_25503,N_24923,N_24938);
and U25504 (N_25504,N_24770,N_25169);
nor U25505 (N_25505,N_24717,N_24832);
or U25506 (N_25506,N_24962,N_24733);
and U25507 (N_25507,N_25158,N_25166);
nand U25508 (N_25508,N_25009,N_25110);
xor U25509 (N_25509,N_24693,N_24959);
xor U25510 (N_25510,N_24792,N_24961);
xnor U25511 (N_25511,N_24806,N_24966);
nand U25512 (N_25512,N_25020,N_24745);
or U25513 (N_25513,N_24689,N_24986);
or U25514 (N_25514,N_24913,N_24755);
xor U25515 (N_25515,N_25151,N_24937);
xor U25516 (N_25516,N_24734,N_24855);
nand U25517 (N_25517,N_24831,N_24818);
nand U25518 (N_25518,N_25011,N_24923);
and U25519 (N_25519,N_25100,N_24846);
and U25520 (N_25520,N_24903,N_24795);
nor U25521 (N_25521,N_25054,N_24725);
xor U25522 (N_25522,N_24851,N_25107);
xnor U25523 (N_25523,N_25083,N_24634);
nor U25524 (N_25524,N_24724,N_24662);
nand U25525 (N_25525,N_24711,N_24958);
nor U25526 (N_25526,N_24931,N_24711);
nand U25527 (N_25527,N_24927,N_24727);
or U25528 (N_25528,N_25002,N_24866);
and U25529 (N_25529,N_25050,N_24809);
nand U25530 (N_25530,N_24891,N_25008);
and U25531 (N_25531,N_24742,N_24964);
nor U25532 (N_25532,N_24620,N_24787);
nor U25533 (N_25533,N_25044,N_25008);
or U25534 (N_25534,N_24695,N_25087);
nand U25535 (N_25535,N_24847,N_24903);
and U25536 (N_25536,N_24758,N_25037);
nand U25537 (N_25537,N_25087,N_24868);
xor U25538 (N_25538,N_24764,N_25136);
xor U25539 (N_25539,N_24899,N_25090);
or U25540 (N_25540,N_24987,N_25113);
or U25541 (N_25541,N_25095,N_24772);
and U25542 (N_25542,N_25109,N_24710);
nor U25543 (N_25543,N_24866,N_24949);
or U25544 (N_25544,N_24856,N_24828);
or U25545 (N_25545,N_24609,N_24713);
nor U25546 (N_25546,N_24729,N_25156);
nor U25547 (N_25547,N_24680,N_25147);
nand U25548 (N_25548,N_25042,N_25019);
or U25549 (N_25549,N_25064,N_25172);
nor U25550 (N_25550,N_24739,N_24744);
xor U25551 (N_25551,N_24674,N_24734);
nand U25552 (N_25552,N_25105,N_24824);
or U25553 (N_25553,N_24713,N_24818);
and U25554 (N_25554,N_24864,N_24947);
xor U25555 (N_25555,N_25019,N_24875);
xor U25556 (N_25556,N_25072,N_24805);
xor U25557 (N_25557,N_24935,N_24844);
and U25558 (N_25558,N_24676,N_24939);
nor U25559 (N_25559,N_24865,N_25034);
nor U25560 (N_25560,N_24968,N_24631);
or U25561 (N_25561,N_24650,N_24990);
xnor U25562 (N_25562,N_24691,N_24623);
or U25563 (N_25563,N_25005,N_24945);
nor U25564 (N_25564,N_24865,N_25046);
or U25565 (N_25565,N_25084,N_24873);
and U25566 (N_25566,N_25065,N_24980);
or U25567 (N_25567,N_24846,N_24817);
xor U25568 (N_25568,N_25062,N_25141);
nor U25569 (N_25569,N_24613,N_24879);
and U25570 (N_25570,N_24601,N_24745);
nor U25571 (N_25571,N_25180,N_25102);
nor U25572 (N_25572,N_24944,N_24625);
nand U25573 (N_25573,N_24732,N_25015);
nand U25574 (N_25574,N_25043,N_24756);
xnor U25575 (N_25575,N_25195,N_25078);
nand U25576 (N_25576,N_24679,N_25188);
and U25577 (N_25577,N_24657,N_24942);
or U25578 (N_25578,N_24836,N_24724);
nor U25579 (N_25579,N_24978,N_24657);
or U25580 (N_25580,N_24620,N_24753);
xnor U25581 (N_25581,N_24664,N_24829);
or U25582 (N_25582,N_24615,N_25058);
or U25583 (N_25583,N_25020,N_25122);
nand U25584 (N_25584,N_24967,N_24963);
or U25585 (N_25585,N_24856,N_25024);
and U25586 (N_25586,N_24724,N_25091);
xor U25587 (N_25587,N_24691,N_25167);
or U25588 (N_25588,N_24968,N_24634);
xnor U25589 (N_25589,N_25067,N_24664);
nor U25590 (N_25590,N_24804,N_25198);
and U25591 (N_25591,N_24608,N_25187);
nor U25592 (N_25592,N_24833,N_24814);
nor U25593 (N_25593,N_25024,N_24731);
or U25594 (N_25594,N_24710,N_24794);
and U25595 (N_25595,N_24710,N_25004);
nand U25596 (N_25596,N_25008,N_25072);
nand U25597 (N_25597,N_24777,N_24990);
and U25598 (N_25598,N_24669,N_24813);
nor U25599 (N_25599,N_24927,N_25037);
or U25600 (N_25600,N_24795,N_25108);
nand U25601 (N_25601,N_24922,N_24985);
nand U25602 (N_25602,N_24930,N_25179);
nor U25603 (N_25603,N_24763,N_25057);
xnor U25604 (N_25604,N_24841,N_24621);
and U25605 (N_25605,N_24954,N_24855);
nor U25606 (N_25606,N_25196,N_24617);
nor U25607 (N_25607,N_24960,N_24601);
nor U25608 (N_25608,N_24926,N_25088);
and U25609 (N_25609,N_24707,N_24710);
or U25610 (N_25610,N_25005,N_24705);
xor U25611 (N_25611,N_25188,N_24809);
xnor U25612 (N_25612,N_25028,N_25014);
xor U25613 (N_25613,N_24985,N_24773);
nand U25614 (N_25614,N_25084,N_25033);
xor U25615 (N_25615,N_24835,N_24853);
xor U25616 (N_25616,N_24618,N_25037);
nand U25617 (N_25617,N_25017,N_24962);
or U25618 (N_25618,N_24654,N_24772);
or U25619 (N_25619,N_24673,N_24658);
and U25620 (N_25620,N_24842,N_25067);
or U25621 (N_25621,N_24942,N_25118);
and U25622 (N_25622,N_25150,N_24607);
xor U25623 (N_25623,N_25046,N_24753);
xnor U25624 (N_25624,N_24958,N_25196);
nor U25625 (N_25625,N_24847,N_25133);
nor U25626 (N_25626,N_24687,N_24936);
nor U25627 (N_25627,N_25134,N_25163);
nor U25628 (N_25628,N_24890,N_24661);
nor U25629 (N_25629,N_24857,N_24662);
and U25630 (N_25630,N_24662,N_24628);
nand U25631 (N_25631,N_25006,N_24697);
and U25632 (N_25632,N_24971,N_25135);
nor U25633 (N_25633,N_25012,N_24850);
and U25634 (N_25634,N_25003,N_24606);
and U25635 (N_25635,N_24777,N_24848);
and U25636 (N_25636,N_24828,N_24691);
or U25637 (N_25637,N_25076,N_24873);
nor U25638 (N_25638,N_24834,N_25066);
and U25639 (N_25639,N_24732,N_25157);
nand U25640 (N_25640,N_24812,N_25143);
nand U25641 (N_25641,N_24618,N_24990);
nand U25642 (N_25642,N_24969,N_25170);
or U25643 (N_25643,N_24780,N_24896);
and U25644 (N_25644,N_25117,N_24970);
nand U25645 (N_25645,N_24693,N_25101);
and U25646 (N_25646,N_24906,N_24623);
or U25647 (N_25647,N_24789,N_24944);
xnor U25648 (N_25648,N_24629,N_24765);
and U25649 (N_25649,N_25095,N_24623);
and U25650 (N_25650,N_24873,N_25031);
and U25651 (N_25651,N_24658,N_24779);
xor U25652 (N_25652,N_24762,N_24735);
xnor U25653 (N_25653,N_25107,N_24879);
xnor U25654 (N_25654,N_24885,N_24934);
nand U25655 (N_25655,N_25061,N_24801);
nor U25656 (N_25656,N_24791,N_25030);
and U25657 (N_25657,N_24643,N_25097);
nor U25658 (N_25658,N_25076,N_24711);
nand U25659 (N_25659,N_24660,N_25162);
or U25660 (N_25660,N_24781,N_25115);
nor U25661 (N_25661,N_24934,N_25191);
or U25662 (N_25662,N_24720,N_24994);
or U25663 (N_25663,N_24742,N_25082);
and U25664 (N_25664,N_24862,N_24658);
nand U25665 (N_25665,N_24808,N_25024);
and U25666 (N_25666,N_25068,N_25008);
nor U25667 (N_25667,N_24715,N_24761);
or U25668 (N_25668,N_25053,N_24835);
and U25669 (N_25669,N_25094,N_24951);
xor U25670 (N_25670,N_24846,N_24865);
or U25671 (N_25671,N_24667,N_24966);
nand U25672 (N_25672,N_24736,N_24682);
nand U25673 (N_25673,N_25100,N_24896);
or U25674 (N_25674,N_25078,N_24726);
or U25675 (N_25675,N_25139,N_24603);
and U25676 (N_25676,N_24716,N_24620);
or U25677 (N_25677,N_25162,N_25042);
xor U25678 (N_25678,N_25045,N_25144);
or U25679 (N_25679,N_24996,N_24770);
nor U25680 (N_25680,N_24918,N_25181);
nor U25681 (N_25681,N_25094,N_24990);
xnor U25682 (N_25682,N_24780,N_25180);
nand U25683 (N_25683,N_25021,N_25055);
nor U25684 (N_25684,N_24603,N_24698);
and U25685 (N_25685,N_24773,N_24847);
nand U25686 (N_25686,N_24654,N_24745);
xor U25687 (N_25687,N_24919,N_24647);
nor U25688 (N_25688,N_24885,N_24648);
xor U25689 (N_25689,N_24780,N_24695);
nor U25690 (N_25690,N_25015,N_24906);
nor U25691 (N_25691,N_25042,N_24945);
xnor U25692 (N_25692,N_24897,N_25064);
or U25693 (N_25693,N_24929,N_24657);
and U25694 (N_25694,N_24758,N_24642);
and U25695 (N_25695,N_24909,N_24923);
or U25696 (N_25696,N_24849,N_24797);
or U25697 (N_25697,N_24693,N_24751);
nand U25698 (N_25698,N_24644,N_24749);
or U25699 (N_25699,N_25024,N_24834);
and U25700 (N_25700,N_24933,N_24667);
xnor U25701 (N_25701,N_24687,N_24974);
or U25702 (N_25702,N_24702,N_25173);
and U25703 (N_25703,N_24712,N_24753);
and U25704 (N_25704,N_24734,N_24800);
xnor U25705 (N_25705,N_24932,N_24646);
and U25706 (N_25706,N_25165,N_25162);
and U25707 (N_25707,N_24713,N_24980);
and U25708 (N_25708,N_25183,N_24710);
nand U25709 (N_25709,N_24711,N_24617);
nand U25710 (N_25710,N_25144,N_25041);
nor U25711 (N_25711,N_25195,N_24774);
xor U25712 (N_25712,N_25103,N_25147);
xor U25713 (N_25713,N_25195,N_25143);
nand U25714 (N_25714,N_25180,N_24776);
xnor U25715 (N_25715,N_24810,N_24831);
nor U25716 (N_25716,N_25032,N_25143);
xnor U25717 (N_25717,N_24764,N_24668);
xor U25718 (N_25718,N_24983,N_25163);
and U25719 (N_25719,N_24998,N_24601);
or U25720 (N_25720,N_24938,N_24865);
nand U25721 (N_25721,N_25063,N_24789);
or U25722 (N_25722,N_25092,N_24656);
xor U25723 (N_25723,N_25007,N_24696);
xor U25724 (N_25724,N_24690,N_24822);
xor U25725 (N_25725,N_24698,N_24719);
xnor U25726 (N_25726,N_25101,N_24930);
or U25727 (N_25727,N_25077,N_24645);
and U25728 (N_25728,N_25108,N_25045);
and U25729 (N_25729,N_25019,N_24668);
nand U25730 (N_25730,N_25088,N_24734);
and U25731 (N_25731,N_24613,N_24797);
nor U25732 (N_25732,N_24902,N_25094);
and U25733 (N_25733,N_24670,N_25182);
and U25734 (N_25734,N_24864,N_24844);
xor U25735 (N_25735,N_24819,N_24621);
xor U25736 (N_25736,N_24800,N_25049);
or U25737 (N_25737,N_24610,N_24739);
xnor U25738 (N_25738,N_24995,N_24751);
and U25739 (N_25739,N_25073,N_25016);
nand U25740 (N_25740,N_25143,N_24619);
nand U25741 (N_25741,N_24767,N_24890);
or U25742 (N_25742,N_24726,N_25189);
and U25743 (N_25743,N_24978,N_24697);
nor U25744 (N_25744,N_24808,N_25096);
nor U25745 (N_25745,N_25004,N_24696);
xor U25746 (N_25746,N_25010,N_25068);
or U25747 (N_25747,N_24629,N_24953);
nand U25748 (N_25748,N_24734,N_24835);
xor U25749 (N_25749,N_24761,N_24970);
and U25750 (N_25750,N_24636,N_24640);
or U25751 (N_25751,N_24727,N_24896);
xor U25752 (N_25752,N_24699,N_24919);
xnor U25753 (N_25753,N_24720,N_25107);
nor U25754 (N_25754,N_24708,N_24707);
nor U25755 (N_25755,N_24749,N_24934);
or U25756 (N_25756,N_24677,N_24629);
nor U25757 (N_25757,N_25047,N_25066);
xor U25758 (N_25758,N_24634,N_24652);
or U25759 (N_25759,N_24920,N_25063);
nor U25760 (N_25760,N_25134,N_24788);
and U25761 (N_25761,N_24707,N_25074);
xor U25762 (N_25762,N_25028,N_25143);
and U25763 (N_25763,N_25184,N_24684);
or U25764 (N_25764,N_24967,N_24797);
nand U25765 (N_25765,N_24786,N_25116);
nand U25766 (N_25766,N_25189,N_24687);
nor U25767 (N_25767,N_24724,N_24717);
and U25768 (N_25768,N_24769,N_25138);
nor U25769 (N_25769,N_25168,N_25145);
and U25770 (N_25770,N_24752,N_24617);
xor U25771 (N_25771,N_24803,N_24614);
xnor U25772 (N_25772,N_24790,N_24968);
and U25773 (N_25773,N_24757,N_24685);
or U25774 (N_25774,N_24870,N_25057);
nor U25775 (N_25775,N_25008,N_24912);
nor U25776 (N_25776,N_24893,N_24964);
or U25777 (N_25777,N_24678,N_24982);
and U25778 (N_25778,N_24764,N_24989);
or U25779 (N_25779,N_24685,N_25067);
or U25780 (N_25780,N_25042,N_24651);
and U25781 (N_25781,N_24996,N_24836);
and U25782 (N_25782,N_25066,N_25068);
and U25783 (N_25783,N_25096,N_24972);
or U25784 (N_25784,N_24633,N_24644);
and U25785 (N_25785,N_24755,N_24884);
or U25786 (N_25786,N_25034,N_24740);
nand U25787 (N_25787,N_24702,N_24748);
xnor U25788 (N_25788,N_25168,N_25167);
or U25789 (N_25789,N_24849,N_24958);
xnor U25790 (N_25790,N_25065,N_24919);
nand U25791 (N_25791,N_24623,N_24800);
and U25792 (N_25792,N_24745,N_24698);
nand U25793 (N_25793,N_24612,N_24606);
nor U25794 (N_25794,N_24840,N_24980);
or U25795 (N_25795,N_24824,N_24615);
or U25796 (N_25796,N_24663,N_25107);
xnor U25797 (N_25797,N_25114,N_24948);
or U25798 (N_25798,N_25008,N_24722);
xnor U25799 (N_25799,N_24634,N_25137);
nand U25800 (N_25800,N_25278,N_25654);
xnor U25801 (N_25801,N_25304,N_25318);
nor U25802 (N_25802,N_25424,N_25390);
nor U25803 (N_25803,N_25410,N_25203);
xnor U25804 (N_25804,N_25350,N_25411);
nand U25805 (N_25805,N_25574,N_25566);
or U25806 (N_25806,N_25261,N_25564);
or U25807 (N_25807,N_25495,N_25699);
xnor U25808 (N_25808,N_25263,N_25353);
nor U25809 (N_25809,N_25751,N_25641);
nand U25810 (N_25810,N_25563,N_25334);
and U25811 (N_25811,N_25493,N_25282);
and U25812 (N_25812,N_25218,N_25775);
or U25813 (N_25813,N_25548,N_25670);
or U25814 (N_25814,N_25719,N_25594);
and U25815 (N_25815,N_25302,N_25447);
or U25816 (N_25816,N_25403,N_25718);
and U25817 (N_25817,N_25363,N_25264);
xnor U25818 (N_25818,N_25409,N_25682);
or U25819 (N_25819,N_25680,N_25454);
nand U25820 (N_25820,N_25287,N_25288);
nor U25821 (N_25821,N_25477,N_25676);
or U25822 (N_25822,N_25590,N_25244);
nand U25823 (N_25823,N_25637,N_25734);
and U25824 (N_25824,N_25300,N_25456);
nor U25825 (N_25825,N_25484,N_25588);
nand U25826 (N_25826,N_25402,N_25742);
nor U25827 (N_25827,N_25233,N_25247);
or U25828 (N_25828,N_25679,N_25219);
nor U25829 (N_25829,N_25327,N_25643);
nor U25830 (N_25830,N_25416,N_25313);
nand U25831 (N_25831,N_25202,N_25509);
or U25832 (N_25832,N_25686,N_25624);
or U25833 (N_25833,N_25413,N_25607);
xnor U25834 (N_25834,N_25284,N_25489);
or U25835 (N_25835,N_25796,N_25614);
nor U25836 (N_25836,N_25726,N_25227);
nand U25837 (N_25837,N_25464,N_25246);
or U25838 (N_25838,N_25364,N_25746);
xnor U25839 (N_25839,N_25513,N_25757);
or U25840 (N_25840,N_25440,N_25492);
xor U25841 (N_25841,N_25605,N_25298);
nor U25842 (N_25842,N_25538,N_25581);
and U25843 (N_25843,N_25703,N_25226);
nor U25844 (N_25844,N_25317,N_25683);
or U25845 (N_25845,N_25595,N_25729);
and U25846 (N_25846,N_25740,N_25367);
and U25847 (N_25847,N_25618,N_25391);
and U25848 (N_25848,N_25475,N_25270);
and U25849 (N_25849,N_25356,N_25379);
nor U25850 (N_25850,N_25268,N_25530);
nand U25851 (N_25851,N_25343,N_25553);
xor U25852 (N_25852,N_25617,N_25250);
xnor U25853 (N_25853,N_25591,N_25400);
nor U25854 (N_25854,N_25764,N_25319);
nand U25855 (N_25855,N_25545,N_25612);
nor U25856 (N_25856,N_25584,N_25488);
xor U25857 (N_25857,N_25421,N_25442);
or U25858 (N_25858,N_25779,N_25474);
xor U25859 (N_25859,N_25639,N_25341);
nand U25860 (N_25860,N_25205,N_25648);
nand U25861 (N_25861,N_25370,N_25234);
and U25862 (N_25862,N_25557,N_25646);
nor U25863 (N_25863,N_25321,N_25256);
or U25864 (N_25864,N_25510,N_25295);
or U25865 (N_25865,N_25453,N_25254);
nor U25866 (N_25866,N_25542,N_25497);
nand U25867 (N_25867,N_25312,N_25438);
xor U25868 (N_25868,N_25737,N_25422);
nor U25869 (N_25869,N_25677,N_25231);
nand U25870 (N_25870,N_25655,N_25745);
nand U25871 (N_25871,N_25790,N_25396);
and U25872 (N_25872,N_25596,N_25361);
or U25873 (N_25873,N_25266,N_25522);
nand U25874 (N_25874,N_25487,N_25665);
nand U25875 (N_25875,N_25499,N_25380);
and U25876 (N_25876,N_25210,N_25385);
nand U25877 (N_25877,N_25782,N_25406);
or U25878 (N_25878,N_25441,N_25430);
and U25879 (N_25879,N_25723,N_25393);
nor U25880 (N_25880,N_25613,N_25537);
xnor U25881 (N_25881,N_25412,N_25242);
nand U25882 (N_25882,N_25223,N_25759);
nand U25883 (N_25883,N_25708,N_25389);
nor U25884 (N_25884,N_25797,N_25352);
xnor U25885 (N_25885,N_25539,N_25299);
xor U25886 (N_25886,N_25705,N_25798);
or U25887 (N_25887,N_25372,N_25650);
nand U25888 (N_25888,N_25669,N_25518);
and U25889 (N_25889,N_25238,N_25761);
nor U25890 (N_25890,N_25448,N_25692);
nand U25891 (N_25891,N_25360,N_25490);
xnor U25892 (N_25892,N_25371,N_25307);
nor U25893 (N_25893,N_25633,N_25551);
or U25894 (N_25894,N_25444,N_25659);
nand U25895 (N_25895,N_25697,N_25662);
nand U25896 (N_25896,N_25600,N_25204);
nor U25897 (N_25897,N_25672,N_25582);
nand U25898 (N_25898,N_25407,N_25735);
nand U25899 (N_25899,N_25731,N_25359);
and U25900 (N_25900,N_25273,N_25554);
or U25901 (N_25901,N_25575,N_25434);
nor U25902 (N_25902,N_25674,N_25373);
nor U25903 (N_25903,N_25652,N_25713);
xnor U25904 (N_25904,N_25435,N_25230);
nand U25905 (N_25905,N_25215,N_25388);
nand U25906 (N_25906,N_25336,N_25636);
or U25907 (N_25907,N_25786,N_25675);
or U25908 (N_25908,N_25211,N_25512);
nor U25909 (N_25909,N_25747,N_25251);
nor U25910 (N_25910,N_25606,N_25766);
or U25911 (N_25911,N_25452,N_25774);
xnor U25912 (N_25912,N_25329,N_25239);
or U25913 (N_25913,N_25698,N_25781);
or U25914 (N_25914,N_25339,N_25638);
nor U25915 (N_25915,N_25561,N_25365);
xnor U25916 (N_25916,N_25583,N_25736);
xor U25917 (N_25917,N_25503,N_25611);
and U25918 (N_25918,N_25622,N_25756);
nor U25919 (N_25919,N_25661,N_25232);
xor U25920 (N_25920,N_25292,N_25324);
and U25921 (N_25921,N_25303,N_25501);
nor U25922 (N_25922,N_25533,N_25541);
nand U25923 (N_25923,N_25506,N_25269);
nand U25924 (N_25924,N_25525,N_25604);
or U25925 (N_25925,N_25763,N_25465);
and U25926 (N_25926,N_25634,N_25463);
or U25927 (N_25927,N_25549,N_25651);
nor U25928 (N_25928,N_25445,N_25241);
xnor U25929 (N_25929,N_25631,N_25340);
nor U25930 (N_25930,N_25476,N_25658);
nand U25931 (N_25931,N_25788,N_25418);
and U25932 (N_25932,N_25656,N_25310);
nor U25933 (N_25933,N_25296,N_25647);
and U25934 (N_25934,N_25458,N_25570);
nand U25935 (N_25935,N_25377,N_25381);
nor U25936 (N_25936,N_25259,N_25758);
xor U25937 (N_25937,N_25320,N_25220);
and U25938 (N_25938,N_25291,N_25635);
and U25939 (N_25939,N_25593,N_25265);
xor U25940 (N_25940,N_25369,N_25399);
and U25941 (N_25941,N_25335,N_25481);
or U25942 (N_25942,N_25550,N_25450);
or U25943 (N_25943,N_25212,N_25527);
xor U25944 (N_25944,N_25768,N_25696);
xnor U25945 (N_25945,N_25619,N_25540);
or U25946 (N_25946,N_25602,N_25201);
nand U25947 (N_25947,N_25744,N_25383);
nor U25948 (N_25948,N_25678,N_25290);
nand U25949 (N_25949,N_25494,N_25671);
nand U25950 (N_25950,N_25355,N_25689);
xor U25951 (N_25951,N_25260,N_25394);
and U25952 (N_25952,N_25565,N_25289);
xnor U25953 (N_25953,N_25623,N_25701);
or U25954 (N_25954,N_25741,N_25576);
and U25955 (N_25955,N_25280,N_25514);
and U25956 (N_25956,N_25274,N_25459);
xor U25957 (N_25957,N_25249,N_25547);
and U25958 (N_25958,N_25610,N_25222);
nand U25959 (N_25959,N_25479,N_25237);
xnor U25960 (N_25960,N_25668,N_25235);
and U25961 (N_25961,N_25787,N_25657);
nand U25962 (N_25962,N_25748,N_25532);
and U25963 (N_25963,N_25560,N_25630);
and U25964 (N_25964,N_25586,N_25415);
and U25965 (N_25965,N_25375,N_25649);
or U25966 (N_25966,N_25534,N_25704);
nor U25967 (N_25967,N_25626,N_25221);
and U25968 (N_25968,N_25520,N_25414);
and U25969 (N_25969,N_25694,N_25608);
nand U25970 (N_25970,N_25653,N_25301);
xnor U25971 (N_25971,N_25433,N_25598);
or U25972 (N_25972,N_25519,N_25555);
or U25973 (N_25973,N_25710,N_25257);
or U25974 (N_25974,N_25378,N_25286);
nor U25975 (N_25975,N_25240,N_25620);
and U25976 (N_25976,N_25724,N_25754);
and U25977 (N_25977,N_25208,N_25449);
or U25978 (N_25978,N_25755,N_25770);
or U25979 (N_25979,N_25516,N_25603);
and U25980 (N_25980,N_25358,N_25794);
and U25981 (N_25981,N_25673,N_25248);
nand U25982 (N_25982,N_25599,N_25423);
nand U25983 (N_25983,N_25792,N_25640);
and U25984 (N_25984,N_25521,N_25386);
xor U25985 (N_25985,N_25368,N_25200);
xor U25986 (N_25986,N_25773,N_25348);
nor U25987 (N_25987,N_25795,N_25294);
or U25988 (N_25988,N_25285,N_25397);
nor U25989 (N_25989,N_25228,N_25702);
and U25990 (N_25990,N_25486,N_25332);
nand U25991 (N_25991,N_25799,N_25727);
nand U25992 (N_25992,N_25712,N_25217);
and U25993 (N_25993,N_25467,N_25717);
xnor U25994 (N_25994,N_25739,N_25419);
nand U25995 (N_25995,N_25515,N_25535);
xor U25996 (N_25996,N_25362,N_25722);
xnor U25997 (N_25997,N_25482,N_25688);
nor U25998 (N_25998,N_25589,N_25609);
nand U25999 (N_25999,N_25711,N_25427);
nand U26000 (N_26000,N_25568,N_25667);
nor U26001 (N_26001,N_25436,N_25483);
nand U26002 (N_26002,N_25432,N_25354);
and U26003 (N_26003,N_25730,N_25267);
and U26004 (N_26004,N_25376,N_25750);
nor U26005 (N_26005,N_25401,N_25245);
and U26006 (N_26006,N_25460,N_25780);
and U26007 (N_26007,N_25272,N_25349);
xor U26008 (N_26008,N_25491,N_25695);
nand U26009 (N_26009,N_25597,N_25209);
nand U26010 (N_26010,N_25255,N_25714);
or U26011 (N_26011,N_25243,N_25429);
and U26012 (N_26012,N_25338,N_25342);
or U26013 (N_26013,N_25536,N_25225);
xnor U26014 (N_26014,N_25398,N_25733);
xnor U26015 (N_26015,N_25732,N_25496);
or U26016 (N_26016,N_25507,N_25504);
or U26017 (N_26017,N_25451,N_25687);
nand U26018 (N_26018,N_25666,N_25559);
or U26019 (N_26019,N_25743,N_25505);
or U26020 (N_26020,N_25431,N_25769);
nor U26021 (N_26021,N_25544,N_25439);
xor U26022 (N_26022,N_25425,N_25328);
nor U26023 (N_26023,N_25587,N_25366);
or U26024 (N_26024,N_25715,N_25793);
nor U26025 (N_26025,N_25615,N_25738);
and U26026 (N_26026,N_25473,N_25275);
xor U26027 (N_26027,N_25592,N_25469);
or U26028 (N_26028,N_25405,N_25783);
or U26029 (N_26029,N_25660,N_25420);
nor U26030 (N_26030,N_25480,N_25567);
or U26031 (N_26031,N_25572,N_25772);
or U26032 (N_26032,N_25236,N_25784);
nor U26033 (N_26033,N_25778,N_25326);
nor U26034 (N_26034,N_25214,N_25485);
nor U26035 (N_26035,N_25315,N_25752);
and U26036 (N_26036,N_25767,N_25771);
nand U26037 (N_26037,N_25791,N_25314);
or U26038 (N_26038,N_25322,N_25279);
xnor U26039 (N_26039,N_25466,N_25345);
or U26040 (N_26040,N_25517,N_25691);
nand U26041 (N_26041,N_25252,N_25580);
nand U26042 (N_26042,N_25585,N_25281);
xor U26043 (N_26043,N_25663,N_25681);
nand U26044 (N_26044,N_25706,N_25543);
or U26045 (N_26045,N_25344,N_25556);
xor U26046 (N_26046,N_25297,N_25625);
or U26047 (N_26047,N_25524,N_25229);
nor U26048 (N_26048,N_25558,N_25627);
xor U26049 (N_26049,N_25428,N_25351);
xor U26050 (N_26050,N_25309,N_25392);
and U26051 (N_26051,N_25569,N_25621);
and U26052 (N_26052,N_25404,N_25562);
or U26053 (N_26053,N_25446,N_25725);
nor U26054 (N_26054,N_25276,N_25628);
xnor U26055 (N_26055,N_25461,N_25789);
or U26056 (N_26056,N_25721,N_25395);
and U26057 (N_26057,N_25258,N_25384);
xnor U26058 (N_26058,N_25206,N_25762);
nor U26059 (N_26059,N_25426,N_25508);
nand U26060 (N_26060,N_25293,N_25776);
and U26061 (N_26061,N_25213,N_25330);
nand U26062 (N_26062,N_25523,N_25316);
nand U26063 (N_26063,N_25632,N_25308);
and U26064 (N_26064,N_25707,N_25601);
and U26065 (N_26065,N_25526,N_25577);
or U26066 (N_26066,N_25765,N_25437);
or U26067 (N_26067,N_25224,N_25753);
nand U26068 (N_26068,N_25374,N_25690);
nand U26069 (N_26069,N_25785,N_25531);
nand U26070 (N_26070,N_25271,N_25529);
nand U26071 (N_26071,N_25500,N_25664);
nand U26072 (N_26072,N_25498,N_25457);
and U26073 (N_26073,N_25305,N_25471);
and U26074 (N_26074,N_25337,N_25262);
nor U26075 (N_26075,N_25684,N_25645);
nand U26076 (N_26076,N_25579,N_25616);
nand U26077 (N_26077,N_25323,N_25777);
or U26078 (N_26078,N_25760,N_25216);
nor U26079 (N_26079,N_25387,N_25716);
xnor U26080 (N_26080,N_25573,N_25642);
nor U26081 (N_26081,N_25685,N_25478);
and U26082 (N_26082,N_25472,N_25720);
nand U26083 (N_26083,N_25700,N_25283);
or U26084 (N_26084,N_25306,N_25357);
xnor U26085 (N_26085,N_25644,N_25207);
nor U26086 (N_26086,N_25408,N_25511);
and U26087 (N_26087,N_25528,N_25325);
xor U26088 (N_26088,N_25693,N_25253);
xor U26089 (N_26089,N_25470,N_25749);
xnor U26090 (N_26090,N_25502,N_25331);
or U26091 (N_26091,N_25462,N_25277);
or U26092 (N_26092,N_25311,N_25629);
or U26093 (N_26093,N_25443,N_25455);
xor U26094 (N_26094,N_25347,N_25709);
xor U26095 (N_26095,N_25382,N_25578);
nor U26096 (N_26096,N_25552,N_25346);
and U26097 (N_26097,N_25546,N_25333);
or U26098 (N_26098,N_25468,N_25571);
nand U26099 (N_26099,N_25417,N_25728);
nand U26100 (N_26100,N_25652,N_25752);
and U26101 (N_26101,N_25230,N_25495);
and U26102 (N_26102,N_25298,N_25375);
nor U26103 (N_26103,N_25471,N_25539);
nand U26104 (N_26104,N_25248,N_25312);
nor U26105 (N_26105,N_25698,N_25612);
nand U26106 (N_26106,N_25738,N_25314);
or U26107 (N_26107,N_25243,N_25632);
or U26108 (N_26108,N_25589,N_25359);
nand U26109 (N_26109,N_25245,N_25302);
or U26110 (N_26110,N_25645,N_25509);
xnor U26111 (N_26111,N_25760,N_25609);
and U26112 (N_26112,N_25709,N_25647);
or U26113 (N_26113,N_25763,N_25742);
nor U26114 (N_26114,N_25216,N_25787);
and U26115 (N_26115,N_25498,N_25494);
nand U26116 (N_26116,N_25424,N_25308);
xor U26117 (N_26117,N_25303,N_25449);
nor U26118 (N_26118,N_25275,N_25589);
nand U26119 (N_26119,N_25276,N_25226);
nand U26120 (N_26120,N_25309,N_25717);
nand U26121 (N_26121,N_25497,N_25330);
and U26122 (N_26122,N_25710,N_25672);
or U26123 (N_26123,N_25401,N_25248);
or U26124 (N_26124,N_25637,N_25755);
or U26125 (N_26125,N_25380,N_25590);
or U26126 (N_26126,N_25403,N_25746);
and U26127 (N_26127,N_25562,N_25784);
nor U26128 (N_26128,N_25312,N_25693);
nand U26129 (N_26129,N_25442,N_25629);
or U26130 (N_26130,N_25612,N_25594);
nand U26131 (N_26131,N_25310,N_25683);
nor U26132 (N_26132,N_25269,N_25708);
and U26133 (N_26133,N_25745,N_25444);
nor U26134 (N_26134,N_25393,N_25239);
and U26135 (N_26135,N_25381,N_25492);
xnor U26136 (N_26136,N_25543,N_25386);
nor U26137 (N_26137,N_25324,N_25540);
nor U26138 (N_26138,N_25401,N_25442);
or U26139 (N_26139,N_25420,N_25765);
nand U26140 (N_26140,N_25339,N_25791);
nor U26141 (N_26141,N_25374,N_25425);
or U26142 (N_26142,N_25632,N_25515);
or U26143 (N_26143,N_25392,N_25235);
nor U26144 (N_26144,N_25486,N_25387);
and U26145 (N_26145,N_25546,N_25578);
nand U26146 (N_26146,N_25372,N_25623);
nor U26147 (N_26147,N_25226,N_25566);
xor U26148 (N_26148,N_25258,N_25296);
xnor U26149 (N_26149,N_25402,N_25709);
nor U26150 (N_26150,N_25369,N_25245);
and U26151 (N_26151,N_25332,N_25447);
nand U26152 (N_26152,N_25407,N_25435);
nand U26153 (N_26153,N_25388,N_25337);
nand U26154 (N_26154,N_25352,N_25588);
nor U26155 (N_26155,N_25290,N_25336);
nand U26156 (N_26156,N_25554,N_25583);
or U26157 (N_26157,N_25602,N_25504);
nor U26158 (N_26158,N_25381,N_25658);
nand U26159 (N_26159,N_25601,N_25201);
xor U26160 (N_26160,N_25511,N_25554);
or U26161 (N_26161,N_25673,N_25334);
nand U26162 (N_26162,N_25532,N_25757);
nand U26163 (N_26163,N_25201,N_25382);
or U26164 (N_26164,N_25346,N_25440);
and U26165 (N_26165,N_25770,N_25273);
and U26166 (N_26166,N_25752,N_25230);
nand U26167 (N_26167,N_25472,N_25698);
and U26168 (N_26168,N_25621,N_25600);
nor U26169 (N_26169,N_25509,N_25583);
xnor U26170 (N_26170,N_25328,N_25212);
nor U26171 (N_26171,N_25780,N_25561);
nor U26172 (N_26172,N_25424,N_25480);
xor U26173 (N_26173,N_25701,N_25225);
xnor U26174 (N_26174,N_25219,N_25413);
or U26175 (N_26175,N_25531,N_25463);
nor U26176 (N_26176,N_25388,N_25698);
nor U26177 (N_26177,N_25473,N_25403);
and U26178 (N_26178,N_25699,N_25394);
nand U26179 (N_26179,N_25452,N_25548);
xor U26180 (N_26180,N_25320,N_25245);
and U26181 (N_26181,N_25717,N_25294);
nand U26182 (N_26182,N_25202,N_25589);
and U26183 (N_26183,N_25218,N_25314);
or U26184 (N_26184,N_25260,N_25712);
xor U26185 (N_26185,N_25435,N_25381);
nor U26186 (N_26186,N_25402,N_25652);
nor U26187 (N_26187,N_25471,N_25311);
xnor U26188 (N_26188,N_25528,N_25784);
or U26189 (N_26189,N_25396,N_25710);
or U26190 (N_26190,N_25598,N_25204);
or U26191 (N_26191,N_25239,N_25509);
nor U26192 (N_26192,N_25364,N_25301);
nand U26193 (N_26193,N_25746,N_25672);
nor U26194 (N_26194,N_25742,N_25218);
nor U26195 (N_26195,N_25537,N_25680);
and U26196 (N_26196,N_25512,N_25254);
xnor U26197 (N_26197,N_25427,N_25714);
nand U26198 (N_26198,N_25521,N_25739);
and U26199 (N_26199,N_25218,N_25431);
nand U26200 (N_26200,N_25604,N_25770);
or U26201 (N_26201,N_25561,N_25472);
nand U26202 (N_26202,N_25736,N_25252);
nand U26203 (N_26203,N_25565,N_25473);
and U26204 (N_26204,N_25547,N_25622);
and U26205 (N_26205,N_25310,N_25603);
nor U26206 (N_26206,N_25295,N_25205);
nor U26207 (N_26207,N_25699,N_25632);
nor U26208 (N_26208,N_25238,N_25774);
and U26209 (N_26209,N_25288,N_25319);
nor U26210 (N_26210,N_25243,N_25444);
or U26211 (N_26211,N_25645,N_25228);
nor U26212 (N_26212,N_25570,N_25432);
or U26213 (N_26213,N_25437,N_25561);
or U26214 (N_26214,N_25712,N_25206);
and U26215 (N_26215,N_25480,N_25404);
xor U26216 (N_26216,N_25376,N_25549);
or U26217 (N_26217,N_25440,N_25364);
nand U26218 (N_26218,N_25290,N_25667);
or U26219 (N_26219,N_25371,N_25389);
or U26220 (N_26220,N_25492,N_25628);
or U26221 (N_26221,N_25698,N_25799);
and U26222 (N_26222,N_25799,N_25524);
xnor U26223 (N_26223,N_25455,N_25641);
or U26224 (N_26224,N_25506,N_25519);
xor U26225 (N_26225,N_25656,N_25248);
nor U26226 (N_26226,N_25485,N_25361);
or U26227 (N_26227,N_25502,N_25421);
xor U26228 (N_26228,N_25213,N_25491);
and U26229 (N_26229,N_25652,N_25591);
nand U26230 (N_26230,N_25636,N_25730);
and U26231 (N_26231,N_25370,N_25206);
nand U26232 (N_26232,N_25512,N_25228);
nor U26233 (N_26233,N_25500,N_25326);
nor U26234 (N_26234,N_25483,N_25529);
nand U26235 (N_26235,N_25515,N_25503);
nand U26236 (N_26236,N_25722,N_25226);
xor U26237 (N_26237,N_25590,N_25658);
and U26238 (N_26238,N_25342,N_25273);
nand U26239 (N_26239,N_25321,N_25352);
nand U26240 (N_26240,N_25678,N_25216);
and U26241 (N_26241,N_25774,N_25466);
nor U26242 (N_26242,N_25427,N_25456);
or U26243 (N_26243,N_25228,N_25341);
xnor U26244 (N_26244,N_25360,N_25313);
and U26245 (N_26245,N_25616,N_25420);
xor U26246 (N_26246,N_25783,N_25359);
nor U26247 (N_26247,N_25671,N_25782);
nor U26248 (N_26248,N_25242,N_25711);
or U26249 (N_26249,N_25350,N_25517);
xor U26250 (N_26250,N_25678,N_25269);
or U26251 (N_26251,N_25290,N_25537);
xnor U26252 (N_26252,N_25249,N_25369);
and U26253 (N_26253,N_25254,N_25403);
xnor U26254 (N_26254,N_25785,N_25706);
xor U26255 (N_26255,N_25677,N_25405);
nand U26256 (N_26256,N_25469,N_25331);
xor U26257 (N_26257,N_25498,N_25493);
nor U26258 (N_26258,N_25771,N_25210);
xnor U26259 (N_26259,N_25436,N_25592);
and U26260 (N_26260,N_25696,N_25481);
or U26261 (N_26261,N_25486,N_25396);
nand U26262 (N_26262,N_25476,N_25779);
xnor U26263 (N_26263,N_25502,N_25637);
and U26264 (N_26264,N_25576,N_25233);
or U26265 (N_26265,N_25567,N_25745);
nand U26266 (N_26266,N_25527,N_25294);
nand U26267 (N_26267,N_25341,N_25324);
or U26268 (N_26268,N_25752,N_25607);
nor U26269 (N_26269,N_25628,N_25262);
and U26270 (N_26270,N_25681,N_25453);
nor U26271 (N_26271,N_25755,N_25533);
and U26272 (N_26272,N_25713,N_25458);
nand U26273 (N_26273,N_25348,N_25212);
nand U26274 (N_26274,N_25476,N_25250);
nor U26275 (N_26275,N_25665,N_25258);
and U26276 (N_26276,N_25494,N_25645);
nor U26277 (N_26277,N_25591,N_25752);
nor U26278 (N_26278,N_25660,N_25419);
or U26279 (N_26279,N_25582,N_25522);
xor U26280 (N_26280,N_25251,N_25658);
nor U26281 (N_26281,N_25224,N_25675);
nor U26282 (N_26282,N_25465,N_25559);
nor U26283 (N_26283,N_25257,N_25585);
or U26284 (N_26284,N_25651,N_25717);
xor U26285 (N_26285,N_25523,N_25735);
and U26286 (N_26286,N_25572,N_25214);
xor U26287 (N_26287,N_25420,N_25363);
nand U26288 (N_26288,N_25387,N_25728);
and U26289 (N_26289,N_25515,N_25438);
nor U26290 (N_26290,N_25260,N_25651);
xor U26291 (N_26291,N_25297,N_25270);
or U26292 (N_26292,N_25606,N_25707);
nor U26293 (N_26293,N_25363,N_25536);
nor U26294 (N_26294,N_25675,N_25338);
nand U26295 (N_26295,N_25242,N_25209);
nor U26296 (N_26296,N_25642,N_25406);
and U26297 (N_26297,N_25798,N_25653);
and U26298 (N_26298,N_25577,N_25214);
nand U26299 (N_26299,N_25406,N_25216);
nor U26300 (N_26300,N_25636,N_25776);
or U26301 (N_26301,N_25321,N_25450);
xor U26302 (N_26302,N_25414,N_25441);
or U26303 (N_26303,N_25263,N_25201);
and U26304 (N_26304,N_25578,N_25235);
or U26305 (N_26305,N_25348,N_25699);
and U26306 (N_26306,N_25745,N_25637);
xnor U26307 (N_26307,N_25795,N_25494);
xor U26308 (N_26308,N_25596,N_25594);
and U26309 (N_26309,N_25533,N_25766);
nand U26310 (N_26310,N_25457,N_25329);
or U26311 (N_26311,N_25205,N_25751);
and U26312 (N_26312,N_25484,N_25513);
nor U26313 (N_26313,N_25337,N_25257);
nand U26314 (N_26314,N_25613,N_25752);
xnor U26315 (N_26315,N_25751,N_25535);
and U26316 (N_26316,N_25484,N_25606);
or U26317 (N_26317,N_25253,N_25785);
xnor U26318 (N_26318,N_25760,N_25366);
or U26319 (N_26319,N_25733,N_25530);
nor U26320 (N_26320,N_25287,N_25578);
and U26321 (N_26321,N_25460,N_25787);
and U26322 (N_26322,N_25780,N_25655);
xnor U26323 (N_26323,N_25660,N_25782);
and U26324 (N_26324,N_25384,N_25666);
nor U26325 (N_26325,N_25765,N_25722);
or U26326 (N_26326,N_25747,N_25603);
and U26327 (N_26327,N_25354,N_25495);
xor U26328 (N_26328,N_25558,N_25418);
nor U26329 (N_26329,N_25457,N_25558);
xnor U26330 (N_26330,N_25374,N_25239);
nor U26331 (N_26331,N_25480,N_25592);
and U26332 (N_26332,N_25274,N_25777);
or U26333 (N_26333,N_25429,N_25687);
or U26334 (N_26334,N_25226,N_25538);
and U26335 (N_26335,N_25686,N_25266);
xnor U26336 (N_26336,N_25709,N_25540);
or U26337 (N_26337,N_25454,N_25399);
nor U26338 (N_26338,N_25709,N_25358);
nor U26339 (N_26339,N_25698,N_25420);
and U26340 (N_26340,N_25250,N_25421);
xor U26341 (N_26341,N_25409,N_25248);
xnor U26342 (N_26342,N_25633,N_25488);
or U26343 (N_26343,N_25739,N_25334);
nor U26344 (N_26344,N_25737,N_25426);
nand U26345 (N_26345,N_25363,N_25217);
or U26346 (N_26346,N_25250,N_25530);
xor U26347 (N_26347,N_25247,N_25282);
nand U26348 (N_26348,N_25388,N_25486);
or U26349 (N_26349,N_25701,N_25777);
and U26350 (N_26350,N_25761,N_25514);
and U26351 (N_26351,N_25297,N_25435);
and U26352 (N_26352,N_25526,N_25402);
nor U26353 (N_26353,N_25412,N_25201);
nor U26354 (N_26354,N_25293,N_25638);
and U26355 (N_26355,N_25312,N_25436);
or U26356 (N_26356,N_25433,N_25450);
nor U26357 (N_26357,N_25683,N_25741);
and U26358 (N_26358,N_25793,N_25475);
nand U26359 (N_26359,N_25290,N_25541);
nand U26360 (N_26360,N_25735,N_25559);
or U26361 (N_26361,N_25756,N_25719);
and U26362 (N_26362,N_25442,N_25439);
nor U26363 (N_26363,N_25758,N_25511);
and U26364 (N_26364,N_25568,N_25534);
or U26365 (N_26365,N_25655,N_25335);
and U26366 (N_26366,N_25255,N_25766);
nand U26367 (N_26367,N_25440,N_25632);
and U26368 (N_26368,N_25215,N_25281);
or U26369 (N_26369,N_25710,N_25442);
nand U26370 (N_26370,N_25790,N_25217);
xor U26371 (N_26371,N_25243,N_25322);
and U26372 (N_26372,N_25310,N_25441);
nor U26373 (N_26373,N_25792,N_25553);
nand U26374 (N_26374,N_25445,N_25240);
nor U26375 (N_26375,N_25711,N_25441);
or U26376 (N_26376,N_25242,N_25797);
or U26377 (N_26377,N_25650,N_25287);
or U26378 (N_26378,N_25468,N_25528);
or U26379 (N_26379,N_25771,N_25681);
xnor U26380 (N_26380,N_25361,N_25547);
xnor U26381 (N_26381,N_25668,N_25702);
nand U26382 (N_26382,N_25478,N_25428);
xor U26383 (N_26383,N_25478,N_25730);
nand U26384 (N_26384,N_25219,N_25618);
nor U26385 (N_26385,N_25435,N_25348);
nand U26386 (N_26386,N_25559,N_25509);
xor U26387 (N_26387,N_25616,N_25416);
or U26388 (N_26388,N_25322,N_25493);
nand U26389 (N_26389,N_25480,N_25732);
and U26390 (N_26390,N_25316,N_25650);
nand U26391 (N_26391,N_25670,N_25241);
xnor U26392 (N_26392,N_25619,N_25529);
and U26393 (N_26393,N_25622,N_25421);
xor U26394 (N_26394,N_25602,N_25580);
and U26395 (N_26395,N_25567,N_25689);
xnor U26396 (N_26396,N_25687,N_25301);
and U26397 (N_26397,N_25347,N_25769);
and U26398 (N_26398,N_25538,N_25671);
or U26399 (N_26399,N_25303,N_25342);
nor U26400 (N_26400,N_26075,N_26035);
and U26401 (N_26401,N_25850,N_25967);
nand U26402 (N_26402,N_26117,N_26334);
nand U26403 (N_26403,N_26219,N_25863);
nand U26404 (N_26404,N_26056,N_26032);
xor U26405 (N_26405,N_26010,N_25973);
nand U26406 (N_26406,N_26108,N_26224);
nand U26407 (N_26407,N_26202,N_26366);
nor U26408 (N_26408,N_26335,N_26367);
xnor U26409 (N_26409,N_26391,N_25872);
xor U26410 (N_26410,N_26231,N_25836);
nand U26411 (N_26411,N_25827,N_26396);
nand U26412 (N_26412,N_26167,N_25875);
nand U26413 (N_26413,N_26354,N_26174);
xor U26414 (N_26414,N_25886,N_26166);
and U26415 (N_26415,N_26001,N_26381);
and U26416 (N_26416,N_26038,N_26230);
or U26417 (N_26417,N_26223,N_26241);
nand U26418 (N_26418,N_25834,N_26042);
or U26419 (N_26419,N_26346,N_25940);
or U26420 (N_26420,N_26024,N_26143);
or U26421 (N_26421,N_25873,N_26287);
nand U26422 (N_26422,N_26064,N_26158);
nand U26423 (N_26423,N_26220,N_26003);
or U26424 (N_26424,N_26159,N_25825);
nand U26425 (N_26425,N_25982,N_25903);
nor U26426 (N_26426,N_25972,N_26097);
xor U26427 (N_26427,N_26157,N_25930);
xnor U26428 (N_26428,N_25812,N_26155);
and U26429 (N_26429,N_26000,N_26209);
nor U26430 (N_26430,N_26070,N_26237);
and U26431 (N_26431,N_26076,N_25829);
nand U26432 (N_26432,N_25810,N_26074);
nand U26433 (N_26433,N_25889,N_26058);
nor U26434 (N_26434,N_26011,N_26292);
and U26435 (N_26435,N_26306,N_26265);
or U26436 (N_26436,N_25820,N_25879);
and U26437 (N_26437,N_26267,N_26029);
nor U26438 (N_26438,N_26393,N_26025);
or U26439 (N_26439,N_25946,N_26204);
or U26440 (N_26440,N_26194,N_25932);
xor U26441 (N_26441,N_25884,N_26066);
or U26442 (N_26442,N_26006,N_26180);
or U26443 (N_26443,N_25987,N_26004);
xor U26444 (N_26444,N_26144,N_26007);
nor U26445 (N_26445,N_26200,N_25839);
nor U26446 (N_26446,N_26090,N_26085);
xor U26447 (N_26447,N_25821,N_26197);
nand U26448 (N_26448,N_26254,N_26274);
nor U26449 (N_26449,N_26095,N_25920);
nor U26450 (N_26450,N_26271,N_25801);
nand U26451 (N_26451,N_25811,N_26278);
or U26452 (N_26452,N_26017,N_25990);
xor U26453 (N_26453,N_26033,N_26169);
nand U26454 (N_26454,N_25885,N_26141);
xor U26455 (N_26455,N_26380,N_26350);
and U26456 (N_26456,N_26039,N_26146);
xor U26457 (N_26457,N_26047,N_26187);
or U26458 (N_26458,N_26084,N_26283);
nor U26459 (N_26459,N_26318,N_26092);
nor U26460 (N_26460,N_25916,N_26020);
nor U26461 (N_26461,N_26236,N_26094);
and U26462 (N_26462,N_26082,N_25809);
nor U26463 (N_26463,N_26168,N_26215);
and U26464 (N_26464,N_26028,N_26255);
or U26465 (N_26465,N_26360,N_26014);
and U26466 (N_26466,N_25806,N_25960);
nor U26467 (N_26467,N_25866,N_25907);
and U26468 (N_26468,N_25911,N_26100);
xnor U26469 (N_26469,N_26282,N_25881);
xnor U26470 (N_26470,N_26170,N_25924);
or U26471 (N_26471,N_26310,N_25837);
and U26472 (N_26472,N_25853,N_26218);
xor U26473 (N_26473,N_25888,N_25800);
and U26474 (N_26474,N_25852,N_25986);
nor U26475 (N_26475,N_26044,N_25962);
xnor U26476 (N_26476,N_26379,N_26121);
nor U26477 (N_26477,N_26342,N_26387);
nor U26478 (N_26478,N_26289,N_26164);
nand U26479 (N_26479,N_25926,N_26286);
nand U26480 (N_26480,N_26273,N_25943);
xor U26481 (N_26481,N_26071,N_25938);
or U26482 (N_26482,N_25859,N_25965);
xnor U26483 (N_26483,N_26134,N_26009);
and U26484 (N_26484,N_26152,N_26019);
and U26485 (N_26485,N_25896,N_26055);
or U26486 (N_26486,N_25913,N_25945);
and U26487 (N_26487,N_25985,N_26221);
nor U26488 (N_26488,N_25871,N_26323);
xnor U26489 (N_26489,N_26299,N_25925);
or U26490 (N_26490,N_26199,N_26160);
or U26491 (N_26491,N_25988,N_25909);
nand U26492 (N_26492,N_26312,N_26198);
or U26493 (N_26493,N_25966,N_26002);
or U26494 (N_26494,N_26129,N_25858);
nand U26495 (N_26495,N_26284,N_26301);
xnor U26496 (N_26496,N_26300,N_25844);
xnor U26497 (N_26497,N_25931,N_26295);
xnor U26498 (N_26498,N_25832,N_26232);
xnor U26499 (N_26499,N_25890,N_25848);
xnor U26500 (N_26500,N_26319,N_26131);
nand U26501 (N_26501,N_25833,N_26345);
nand U26502 (N_26502,N_26057,N_26238);
or U26503 (N_26503,N_25955,N_26089);
xor U26504 (N_26504,N_26302,N_26389);
and U26505 (N_26505,N_25906,N_25995);
nor U26506 (N_26506,N_25803,N_25997);
and U26507 (N_26507,N_25808,N_25894);
nor U26508 (N_26508,N_25855,N_25892);
xnor U26509 (N_26509,N_25977,N_26321);
or U26510 (N_26510,N_26244,N_25813);
xnor U26511 (N_26511,N_25893,N_25961);
nor U26512 (N_26512,N_25915,N_26153);
nor U26513 (N_26513,N_26245,N_26373);
nor U26514 (N_26514,N_25921,N_26296);
xor U26515 (N_26515,N_26397,N_26112);
nand U26516 (N_26516,N_25935,N_26163);
or U26517 (N_26517,N_25948,N_26041);
and U26518 (N_26518,N_26088,N_26133);
nor U26519 (N_26519,N_26105,N_25895);
xor U26520 (N_26520,N_26030,N_25878);
nor U26521 (N_26521,N_26316,N_25983);
or U26522 (N_26522,N_26247,N_26288);
xnor U26523 (N_26523,N_26149,N_26102);
nand U26524 (N_26524,N_26322,N_25950);
nand U26525 (N_26525,N_26239,N_25994);
xnor U26526 (N_26526,N_25956,N_26226);
and U26527 (N_26527,N_25814,N_26252);
and U26528 (N_26528,N_26214,N_26353);
nor U26529 (N_26529,N_26190,N_26291);
xor U26530 (N_26530,N_26183,N_26059);
xor U26531 (N_26531,N_25993,N_26358);
nor U26532 (N_26532,N_26383,N_26336);
and U26533 (N_26533,N_25937,N_26398);
or U26534 (N_26534,N_26069,N_26313);
xnor U26535 (N_26535,N_25914,N_26080);
nand U26536 (N_26536,N_26065,N_26176);
and U26537 (N_26537,N_25816,N_25975);
or U26538 (N_26538,N_26052,N_26150);
xor U26539 (N_26539,N_25870,N_26242);
and U26540 (N_26540,N_26365,N_25949);
nor U26541 (N_26541,N_25835,N_26091);
or U26542 (N_26542,N_26258,N_26051);
and U26543 (N_26543,N_26324,N_25992);
xor U26544 (N_26544,N_26061,N_26063);
and U26545 (N_26545,N_26332,N_26196);
and U26546 (N_26546,N_26227,N_26340);
nand U26547 (N_26547,N_26369,N_26062);
nand U26548 (N_26548,N_25849,N_25802);
nor U26549 (N_26549,N_26096,N_26251);
nand U26550 (N_26550,N_25954,N_26048);
nor U26551 (N_26551,N_26109,N_25826);
nand U26552 (N_26552,N_26027,N_26375);
or U26553 (N_26553,N_25856,N_26378);
nand U26554 (N_26554,N_25868,N_25851);
xor U26555 (N_26555,N_26266,N_26103);
and U26556 (N_26556,N_25981,N_26377);
xnor U26557 (N_26557,N_26040,N_26270);
nor U26558 (N_26558,N_26165,N_26280);
xnor U26559 (N_26559,N_26186,N_25807);
nor U26560 (N_26560,N_25928,N_26349);
or U26561 (N_26561,N_26344,N_26297);
nor U26562 (N_26562,N_26113,N_25840);
xor U26563 (N_26563,N_25822,N_26264);
or U26564 (N_26564,N_26077,N_26026);
and U26565 (N_26565,N_26116,N_26118);
xor U26566 (N_26566,N_25865,N_26399);
xnor U26567 (N_26567,N_26339,N_26012);
nand U26568 (N_26568,N_26293,N_26177);
nand U26569 (N_26569,N_25912,N_25980);
nor U26570 (N_26570,N_26384,N_26357);
or U26571 (N_26571,N_26225,N_26326);
or U26572 (N_26572,N_26120,N_26162);
or U26573 (N_26573,N_26208,N_26263);
or U26574 (N_26574,N_26181,N_26317);
or U26575 (N_26575,N_25991,N_25902);
and U26576 (N_26576,N_26046,N_25952);
xor U26577 (N_26577,N_26207,N_26104);
nand U26578 (N_26578,N_26217,N_26151);
or U26579 (N_26579,N_26098,N_26175);
xor U26580 (N_26580,N_25815,N_26193);
xor U26581 (N_26581,N_25819,N_25908);
xor U26582 (N_26582,N_26385,N_26277);
and U26583 (N_26583,N_26216,N_26364);
or U26584 (N_26584,N_26363,N_25976);
and U26585 (N_26585,N_26172,N_26184);
xor U26586 (N_26586,N_25939,N_25867);
xor U26587 (N_26587,N_25984,N_26272);
and U26588 (N_26588,N_25934,N_26171);
nor U26589 (N_26589,N_25963,N_26078);
nand U26590 (N_26590,N_25880,N_26308);
nand U26591 (N_26591,N_26348,N_25971);
xnor U26592 (N_26592,N_25970,N_26081);
xnor U26593 (N_26593,N_25904,N_26212);
nor U26594 (N_26594,N_26083,N_25933);
or U26595 (N_26595,N_26182,N_26362);
and U26596 (N_26596,N_25927,N_25883);
xnor U26597 (N_26597,N_26234,N_25989);
and U26598 (N_26598,N_26013,N_26005);
nand U26599 (N_26599,N_26213,N_26110);
and U26600 (N_26600,N_26136,N_26201);
and U26601 (N_26601,N_26137,N_26205);
nand U26602 (N_26602,N_26068,N_25887);
nand U26603 (N_26603,N_25996,N_26371);
nand U26604 (N_26604,N_26262,N_26229);
xor U26605 (N_26605,N_26279,N_26079);
or U26606 (N_26606,N_25864,N_26388);
and U26607 (N_26607,N_26053,N_25953);
xnor U26608 (N_26608,N_26338,N_26276);
nand U26609 (N_26609,N_26222,N_25917);
xnor U26610 (N_26610,N_26018,N_26359);
or U26611 (N_26611,N_25900,N_26145);
nor U26612 (N_26612,N_26154,N_25830);
nor U26613 (N_26613,N_25823,N_26337);
or U26614 (N_26614,N_26320,N_25899);
or U26615 (N_26615,N_26243,N_25999);
nand U26616 (N_26616,N_26124,N_26086);
nor U26617 (N_26617,N_26132,N_26185);
or U26618 (N_26618,N_26043,N_26123);
and U26619 (N_26619,N_26073,N_26138);
xnor U26620 (N_26620,N_26307,N_25957);
nor U26621 (N_26621,N_26161,N_26303);
or U26622 (N_26622,N_26034,N_26341);
nand U26623 (N_26623,N_26119,N_26093);
xor U26624 (N_26624,N_25824,N_26233);
and U26625 (N_26625,N_26250,N_25862);
nor U26626 (N_26626,N_26189,N_26395);
or U26627 (N_26627,N_26370,N_26260);
xor U26628 (N_26628,N_26268,N_26015);
xnor U26629 (N_26629,N_26281,N_25891);
xnor U26630 (N_26630,N_25874,N_26256);
nor U26631 (N_26631,N_26122,N_25846);
nand U26632 (N_26632,N_26173,N_25882);
and U26633 (N_26633,N_25942,N_26022);
or U26634 (N_26634,N_26101,N_26135);
or U26635 (N_26635,N_25919,N_26178);
and U26636 (N_26636,N_25922,N_25929);
xnor U26637 (N_26637,N_25828,N_26099);
and U26638 (N_26638,N_26253,N_26275);
xnor U26639 (N_26639,N_26188,N_26106);
xor U26640 (N_26640,N_26111,N_25869);
xnor U26641 (N_26641,N_26191,N_26305);
or U26642 (N_26642,N_26021,N_26328);
and U26643 (N_26643,N_26107,N_25818);
and U26644 (N_26644,N_26228,N_25898);
xnor U26645 (N_26645,N_26060,N_26050);
and U26646 (N_26646,N_26142,N_25817);
and U26647 (N_26647,N_26240,N_25843);
or U26648 (N_26648,N_25805,N_26148);
xnor U26649 (N_26649,N_26368,N_26246);
xnor U26650 (N_26650,N_26206,N_26023);
xnor U26651 (N_26651,N_26298,N_25845);
and U26652 (N_26652,N_26072,N_26374);
nand U26653 (N_26653,N_26347,N_25969);
nor U26654 (N_26654,N_25905,N_25831);
and U26655 (N_26655,N_25918,N_26325);
nor U26656 (N_26656,N_26128,N_25841);
nor U26657 (N_26657,N_26248,N_26372);
nand U26658 (N_26658,N_26016,N_26127);
nor U26659 (N_26659,N_25897,N_26343);
xnor U26660 (N_26660,N_26285,N_26294);
nor U26661 (N_26661,N_25910,N_25959);
nand U26662 (N_26662,N_25958,N_26327);
nor U26663 (N_26663,N_25941,N_26195);
nor U26664 (N_26664,N_25842,N_26114);
xnor U26665 (N_26665,N_26179,N_26259);
nand U26666 (N_26666,N_25936,N_25861);
nand U26667 (N_26667,N_26394,N_25944);
nand U26668 (N_26668,N_26355,N_26130);
and U26669 (N_26669,N_25854,N_26356);
or U26670 (N_26670,N_26352,N_26139);
and U26671 (N_26671,N_25947,N_26147);
nand U26672 (N_26672,N_26376,N_25876);
nor U26673 (N_26673,N_25951,N_26304);
or U26674 (N_26674,N_25877,N_26054);
or U26675 (N_26675,N_25838,N_25847);
nand U26676 (N_26676,N_26125,N_25978);
and U26677 (N_26677,N_26192,N_26037);
nor U26678 (N_26678,N_26203,N_26008);
nand U26679 (N_26679,N_26311,N_26036);
nor U26680 (N_26680,N_26210,N_26049);
and U26681 (N_26681,N_26126,N_26390);
or U26682 (N_26682,N_26257,N_25901);
or U26683 (N_26683,N_25860,N_26290);
xor U26684 (N_26684,N_26330,N_25968);
nor U26685 (N_26685,N_26333,N_26156);
nor U26686 (N_26686,N_26261,N_26115);
xnor U26687 (N_26687,N_26329,N_26031);
xnor U26688 (N_26688,N_26211,N_25964);
nor U26689 (N_26689,N_26140,N_26314);
and U26690 (N_26690,N_25923,N_25979);
or U26691 (N_26691,N_26331,N_26351);
or U26692 (N_26692,N_26235,N_25974);
nand U26693 (N_26693,N_25998,N_26315);
nand U26694 (N_26694,N_26249,N_25804);
and U26695 (N_26695,N_26361,N_26045);
nand U26696 (N_26696,N_26269,N_26386);
or U26697 (N_26697,N_26309,N_25857);
xnor U26698 (N_26698,N_26382,N_26087);
and U26699 (N_26699,N_26067,N_26392);
nor U26700 (N_26700,N_25836,N_25970);
and U26701 (N_26701,N_26228,N_26290);
or U26702 (N_26702,N_26157,N_26314);
nand U26703 (N_26703,N_26147,N_26178);
nand U26704 (N_26704,N_26190,N_26146);
xor U26705 (N_26705,N_25887,N_26057);
xor U26706 (N_26706,N_26165,N_25939);
nand U26707 (N_26707,N_26319,N_26191);
nor U26708 (N_26708,N_26165,N_26339);
or U26709 (N_26709,N_26326,N_26167);
nor U26710 (N_26710,N_26208,N_25935);
and U26711 (N_26711,N_26281,N_26133);
and U26712 (N_26712,N_26330,N_26037);
nor U26713 (N_26713,N_26027,N_25849);
and U26714 (N_26714,N_26037,N_26297);
nand U26715 (N_26715,N_26127,N_26013);
xnor U26716 (N_26716,N_26016,N_26148);
nor U26717 (N_26717,N_26311,N_26023);
and U26718 (N_26718,N_26215,N_25975);
xnor U26719 (N_26719,N_26397,N_25894);
or U26720 (N_26720,N_25898,N_25982);
xnor U26721 (N_26721,N_26142,N_26014);
nor U26722 (N_26722,N_26026,N_26216);
nand U26723 (N_26723,N_26387,N_26167);
nand U26724 (N_26724,N_25856,N_25896);
and U26725 (N_26725,N_26163,N_26296);
or U26726 (N_26726,N_26055,N_25939);
or U26727 (N_26727,N_25874,N_26006);
and U26728 (N_26728,N_25895,N_26208);
or U26729 (N_26729,N_26144,N_26026);
nor U26730 (N_26730,N_26073,N_26382);
xor U26731 (N_26731,N_26006,N_25919);
xor U26732 (N_26732,N_26139,N_26060);
or U26733 (N_26733,N_25902,N_25970);
or U26734 (N_26734,N_26093,N_25887);
xnor U26735 (N_26735,N_26349,N_25906);
nand U26736 (N_26736,N_26372,N_26064);
and U26737 (N_26737,N_26013,N_26253);
nor U26738 (N_26738,N_26161,N_26209);
nor U26739 (N_26739,N_26092,N_26185);
nor U26740 (N_26740,N_25944,N_25868);
nand U26741 (N_26741,N_26060,N_26131);
or U26742 (N_26742,N_26219,N_26084);
or U26743 (N_26743,N_26115,N_26228);
or U26744 (N_26744,N_26029,N_26212);
xnor U26745 (N_26745,N_25827,N_26035);
and U26746 (N_26746,N_26147,N_26298);
xor U26747 (N_26747,N_26089,N_26190);
and U26748 (N_26748,N_26273,N_26175);
nor U26749 (N_26749,N_26379,N_26126);
or U26750 (N_26750,N_26249,N_26174);
xor U26751 (N_26751,N_26372,N_26158);
or U26752 (N_26752,N_26132,N_26367);
or U26753 (N_26753,N_25815,N_26029);
xor U26754 (N_26754,N_25926,N_25876);
nor U26755 (N_26755,N_26269,N_26280);
or U26756 (N_26756,N_26132,N_26167);
nor U26757 (N_26757,N_26163,N_26351);
or U26758 (N_26758,N_26117,N_25957);
nor U26759 (N_26759,N_25952,N_25920);
and U26760 (N_26760,N_25959,N_26249);
and U26761 (N_26761,N_26144,N_25849);
nor U26762 (N_26762,N_25980,N_26223);
and U26763 (N_26763,N_26149,N_25870);
nand U26764 (N_26764,N_26272,N_26328);
and U26765 (N_26765,N_26369,N_25986);
xnor U26766 (N_26766,N_26349,N_26027);
nand U26767 (N_26767,N_26362,N_26045);
and U26768 (N_26768,N_26043,N_26098);
or U26769 (N_26769,N_26183,N_25851);
xor U26770 (N_26770,N_26382,N_25968);
xnor U26771 (N_26771,N_26168,N_26338);
or U26772 (N_26772,N_25867,N_25945);
and U26773 (N_26773,N_26333,N_26312);
nor U26774 (N_26774,N_26110,N_26371);
and U26775 (N_26775,N_25863,N_25840);
xor U26776 (N_26776,N_25866,N_25820);
xor U26777 (N_26777,N_25970,N_25914);
xnor U26778 (N_26778,N_25919,N_26094);
nor U26779 (N_26779,N_25970,N_25807);
xnor U26780 (N_26780,N_26370,N_26240);
nor U26781 (N_26781,N_25903,N_26301);
nor U26782 (N_26782,N_26365,N_25841);
nor U26783 (N_26783,N_26106,N_25824);
xnor U26784 (N_26784,N_25897,N_26244);
nor U26785 (N_26785,N_25955,N_25959);
or U26786 (N_26786,N_25964,N_26231);
nand U26787 (N_26787,N_25873,N_25877);
nand U26788 (N_26788,N_26065,N_26025);
or U26789 (N_26789,N_26315,N_25892);
nor U26790 (N_26790,N_26221,N_26029);
or U26791 (N_26791,N_26344,N_26369);
or U26792 (N_26792,N_26190,N_25973);
nor U26793 (N_26793,N_26151,N_25974);
or U26794 (N_26794,N_26176,N_26129);
nand U26795 (N_26795,N_25840,N_26317);
and U26796 (N_26796,N_25923,N_26039);
nor U26797 (N_26797,N_26263,N_26242);
nor U26798 (N_26798,N_25908,N_26380);
or U26799 (N_26799,N_26236,N_25809);
or U26800 (N_26800,N_26288,N_26238);
xor U26801 (N_26801,N_26037,N_26240);
nor U26802 (N_26802,N_26394,N_26135);
nand U26803 (N_26803,N_26056,N_25931);
and U26804 (N_26804,N_26123,N_26347);
nor U26805 (N_26805,N_25920,N_26309);
nor U26806 (N_26806,N_26285,N_26073);
and U26807 (N_26807,N_26335,N_25801);
xor U26808 (N_26808,N_25837,N_26156);
or U26809 (N_26809,N_25949,N_25884);
and U26810 (N_26810,N_26077,N_25829);
nor U26811 (N_26811,N_26220,N_26060);
nand U26812 (N_26812,N_26230,N_26153);
and U26813 (N_26813,N_25904,N_26048);
or U26814 (N_26814,N_26132,N_26260);
xnor U26815 (N_26815,N_26098,N_25837);
or U26816 (N_26816,N_25814,N_25892);
xnor U26817 (N_26817,N_26122,N_26297);
xnor U26818 (N_26818,N_25860,N_26150);
nand U26819 (N_26819,N_25971,N_25967);
and U26820 (N_26820,N_26143,N_26282);
and U26821 (N_26821,N_26283,N_26256);
xnor U26822 (N_26822,N_26107,N_26354);
nand U26823 (N_26823,N_26334,N_25806);
xor U26824 (N_26824,N_25926,N_25875);
nand U26825 (N_26825,N_26263,N_26093);
nor U26826 (N_26826,N_26179,N_26244);
nor U26827 (N_26827,N_26353,N_26013);
xnor U26828 (N_26828,N_26128,N_26296);
xnor U26829 (N_26829,N_25915,N_26190);
nor U26830 (N_26830,N_25814,N_26192);
nor U26831 (N_26831,N_26227,N_26089);
nor U26832 (N_26832,N_25888,N_25898);
and U26833 (N_26833,N_26150,N_26311);
and U26834 (N_26834,N_26296,N_26338);
xnor U26835 (N_26835,N_26296,N_26347);
nor U26836 (N_26836,N_26006,N_26195);
xnor U26837 (N_26837,N_26312,N_25925);
nand U26838 (N_26838,N_26266,N_26205);
and U26839 (N_26839,N_25806,N_26142);
or U26840 (N_26840,N_26333,N_26373);
and U26841 (N_26841,N_25948,N_26205);
and U26842 (N_26842,N_26086,N_26173);
and U26843 (N_26843,N_25928,N_26263);
nand U26844 (N_26844,N_26098,N_25962);
nand U26845 (N_26845,N_26036,N_25859);
and U26846 (N_26846,N_26027,N_25883);
or U26847 (N_26847,N_26396,N_26255);
and U26848 (N_26848,N_26196,N_26117);
and U26849 (N_26849,N_25997,N_25824);
or U26850 (N_26850,N_26233,N_26081);
or U26851 (N_26851,N_26025,N_26163);
xnor U26852 (N_26852,N_26253,N_26012);
nand U26853 (N_26853,N_25988,N_26300);
and U26854 (N_26854,N_26397,N_25844);
nor U26855 (N_26855,N_25975,N_26151);
xnor U26856 (N_26856,N_26104,N_26348);
nor U26857 (N_26857,N_26174,N_26160);
nor U26858 (N_26858,N_25961,N_25878);
nor U26859 (N_26859,N_26015,N_26042);
nand U26860 (N_26860,N_26022,N_26051);
nor U26861 (N_26861,N_26018,N_25894);
and U26862 (N_26862,N_26304,N_25891);
or U26863 (N_26863,N_26283,N_25810);
and U26864 (N_26864,N_26204,N_25965);
or U26865 (N_26865,N_26264,N_26101);
nand U26866 (N_26866,N_26377,N_26072);
and U26867 (N_26867,N_26290,N_26385);
nand U26868 (N_26868,N_25987,N_26380);
xnor U26869 (N_26869,N_26142,N_26076);
and U26870 (N_26870,N_25853,N_26080);
nand U26871 (N_26871,N_26127,N_25949);
nor U26872 (N_26872,N_26234,N_25830);
xnor U26873 (N_26873,N_25832,N_26274);
and U26874 (N_26874,N_26058,N_26170);
nand U26875 (N_26875,N_25892,N_26257);
nor U26876 (N_26876,N_26265,N_25986);
or U26877 (N_26877,N_26200,N_26106);
nand U26878 (N_26878,N_26285,N_25876);
and U26879 (N_26879,N_26076,N_26389);
or U26880 (N_26880,N_26111,N_26326);
xnor U26881 (N_26881,N_25926,N_26350);
nor U26882 (N_26882,N_25877,N_25837);
nor U26883 (N_26883,N_26212,N_25988);
and U26884 (N_26884,N_26032,N_25821);
and U26885 (N_26885,N_26395,N_26204);
xor U26886 (N_26886,N_25825,N_26290);
xor U26887 (N_26887,N_26091,N_25860);
nor U26888 (N_26888,N_25882,N_25979);
and U26889 (N_26889,N_26172,N_26035);
nand U26890 (N_26890,N_26285,N_26350);
and U26891 (N_26891,N_25819,N_26161);
nor U26892 (N_26892,N_26246,N_26365);
nor U26893 (N_26893,N_26098,N_26106);
nor U26894 (N_26894,N_25815,N_26241);
or U26895 (N_26895,N_26018,N_26153);
and U26896 (N_26896,N_26107,N_26382);
nor U26897 (N_26897,N_26317,N_26006);
or U26898 (N_26898,N_25898,N_26365);
or U26899 (N_26899,N_25815,N_26342);
or U26900 (N_26900,N_25872,N_25879);
xnor U26901 (N_26901,N_26271,N_25926);
xnor U26902 (N_26902,N_26012,N_26257);
nand U26903 (N_26903,N_25894,N_25874);
nor U26904 (N_26904,N_25832,N_25971);
xnor U26905 (N_26905,N_26022,N_26371);
and U26906 (N_26906,N_26243,N_25884);
xnor U26907 (N_26907,N_25980,N_26007);
nor U26908 (N_26908,N_26197,N_25909);
nand U26909 (N_26909,N_26096,N_26314);
or U26910 (N_26910,N_25924,N_25941);
nor U26911 (N_26911,N_26076,N_26333);
nor U26912 (N_26912,N_25805,N_25918);
or U26913 (N_26913,N_26349,N_25905);
and U26914 (N_26914,N_26353,N_26393);
and U26915 (N_26915,N_26243,N_26257);
nand U26916 (N_26916,N_26124,N_26363);
nand U26917 (N_26917,N_26101,N_26013);
xnor U26918 (N_26918,N_26074,N_25931);
or U26919 (N_26919,N_25854,N_25951);
or U26920 (N_26920,N_26348,N_25854);
nor U26921 (N_26921,N_26128,N_25894);
or U26922 (N_26922,N_26357,N_26056);
nand U26923 (N_26923,N_26060,N_25991);
xor U26924 (N_26924,N_26343,N_26321);
nor U26925 (N_26925,N_26385,N_26107);
xor U26926 (N_26926,N_25820,N_25994);
or U26927 (N_26927,N_26359,N_26372);
or U26928 (N_26928,N_25966,N_26223);
nand U26929 (N_26929,N_26020,N_26372);
xor U26930 (N_26930,N_26152,N_25853);
and U26931 (N_26931,N_26295,N_26139);
and U26932 (N_26932,N_25977,N_25803);
or U26933 (N_26933,N_26293,N_26182);
or U26934 (N_26934,N_26152,N_26319);
or U26935 (N_26935,N_26308,N_26120);
and U26936 (N_26936,N_26137,N_25896);
nand U26937 (N_26937,N_26353,N_26077);
nor U26938 (N_26938,N_25949,N_25837);
xnor U26939 (N_26939,N_25853,N_25892);
and U26940 (N_26940,N_25968,N_25806);
nor U26941 (N_26941,N_26089,N_26164);
xnor U26942 (N_26942,N_26178,N_25841);
nand U26943 (N_26943,N_25913,N_25980);
nor U26944 (N_26944,N_25801,N_25948);
nor U26945 (N_26945,N_26201,N_26390);
xor U26946 (N_26946,N_26308,N_25844);
and U26947 (N_26947,N_25852,N_26304);
nand U26948 (N_26948,N_26291,N_26343);
or U26949 (N_26949,N_25880,N_26077);
nand U26950 (N_26950,N_26051,N_25870);
xor U26951 (N_26951,N_26294,N_26341);
nor U26952 (N_26952,N_25958,N_25952);
nand U26953 (N_26953,N_26059,N_26032);
nand U26954 (N_26954,N_26276,N_26095);
and U26955 (N_26955,N_25961,N_26177);
nor U26956 (N_26956,N_25976,N_26089);
or U26957 (N_26957,N_25815,N_26024);
or U26958 (N_26958,N_26109,N_26041);
or U26959 (N_26959,N_25889,N_26346);
nor U26960 (N_26960,N_25812,N_26031);
nor U26961 (N_26961,N_26141,N_26368);
and U26962 (N_26962,N_26051,N_26200);
or U26963 (N_26963,N_26211,N_26209);
and U26964 (N_26964,N_26171,N_26194);
xnor U26965 (N_26965,N_26207,N_26376);
xor U26966 (N_26966,N_26246,N_26141);
nor U26967 (N_26967,N_26276,N_26279);
or U26968 (N_26968,N_26017,N_25933);
and U26969 (N_26969,N_26334,N_26281);
xor U26970 (N_26970,N_26023,N_25982);
and U26971 (N_26971,N_26191,N_25982);
and U26972 (N_26972,N_25800,N_26290);
or U26973 (N_26973,N_26025,N_25817);
and U26974 (N_26974,N_25850,N_26248);
nand U26975 (N_26975,N_25917,N_26221);
and U26976 (N_26976,N_26190,N_26032);
or U26977 (N_26977,N_26145,N_25874);
xnor U26978 (N_26978,N_25819,N_26017);
xor U26979 (N_26979,N_26281,N_25873);
nor U26980 (N_26980,N_26125,N_26170);
or U26981 (N_26981,N_26303,N_26176);
xor U26982 (N_26982,N_25901,N_26070);
nand U26983 (N_26983,N_25856,N_26223);
and U26984 (N_26984,N_25934,N_26296);
or U26985 (N_26985,N_25879,N_26295);
nor U26986 (N_26986,N_26305,N_26206);
nor U26987 (N_26987,N_26289,N_26291);
xor U26988 (N_26988,N_26127,N_26095);
and U26989 (N_26989,N_25929,N_26011);
xor U26990 (N_26990,N_26071,N_26260);
nor U26991 (N_26991,N_25961,N_26166);
nor U26992 (N_26992,N_26047,N_26247);
nand U26993 (N_26993,N_26180,N_26119);
nand U26994 (N_26994,N_26129,N_25935);
xnor U26995 (N_26995,N_26208,N_26081);
nor U26996 (N_26996,N_26389,N_26380);
xor U26997 (N_26997,N_26309,N_26003);
or U26998 (N_26998,N_26273,N_26134);
xor U26999 (N_26999,N_26340,N_26304);
or U27000 (N_27000,N_26477,N_26440);
nand U27001 (N_27001,N_26445,N_26682);
and U27002 (N_27002,N_26688,N_26967);
nand U27003 (N_27003,N_26531,N_26559);
nor U27004 (N_27004,N_26500,N_26599);
xor U27005 (N_27005,N_26777,N_26730);
nor U27006 (N_27006,N_26697,N_26853);
nand U27007 (N_27007,N_26683,N_26762);
nand U27008 (N_27008,N_26653,N_26416);
nor U27009 (N_27009,N_26737,N_26489);
nor U27010 (N_27010,N_26917,N_26887);
nand U27011 (N_27011,N_26888,N_26522);
nor U27012 (N_27012,N_26744,N_26767);
and U27013 (N_27013,N_26785,N_26422);
xor U27014 (N_27014,N_26441,N_26756);
nor U27015 (N_27015,N_26454,N_26444);
xor U27016 (N_27016,N_26886,N_26977);
nand U27017 (N_27017,N_26891,N_26474);
nand U27018 (N_27018,N_26790,N_26947);
and U27019 (N_27019,N_26950,N_26834);
xor U27020 (N_27020,N_26548,N_26698);
nor U27021 (N_27021,N_26585,N_26666);
or U27022 (N_27022,N_26504,N_26401);
xor U27023 (N_27023,N_26722,N_26406);
or U27024 (N_27024,N_26897,N_26782);
nor U27025 (N_27025,N_26753,N_26575);
and U27026 (N_27026,N_26818,N_26966);
xor U27027 (N_27027,N_26494,N_26924);
or U27028 (N_27028,N_26600,N_26909);
nor U27029 (N_27029,N_26515,N_26764);
nand U27030 (N_27030,N_26750,N_26501);
nand U27031 (N_27031,N_26847,N_26578);
and U27032 (N_27032,N_26411,N_26775);
nand U27033 (N_27033,N_26569,N_26594);
and U27034 (N_27034,N_26631,N_26632);
and U27035 (N_27035,N_26984,N_26420);
nand U27036 (N_27036,N_26889,N_26997);
and U27037 (N_27037,N_26668,N_26447);
xnor U27038 (N_27038,N_26582,N_26634);
nand U27039 (N_27039,N_26752,N_26604);
xor U27040 (N_27040,N_26603,N_26649);
and U27041 (N_27041,N_26946,N_26996);
or U27042 (N_27042,N_26890,N_26719);
or U27043 (N_27043,N_26506,N_26598);
nand U27044 (N_27044,N_26759,N_26707);
nor U27045 (N_27045,N_26677,N_26667);
xnor U27046 (N_27046,N_26922,N_26532);
or U27047 (N_27047,N_26488,N_26469);
xnor U27048 (N_27048,N_26971,N_26449);
nand U27049 (N_27049,N_26805,N_26681);
nand U27050 (N_27050,N_26560,N_26542);
nand U27051 (N_27051,N_26874,N_26959);
xnor U27052 (N_27052,N_26758,N_26591);
xnor U27053 (N_27053,N_26620,N_26651);
and U27054 (N_27054,N_26590,N_26473);
nor U27055 (N_27055,N_26654,N_26754);
nand U27056 (N_27056,N_26686,N_26828);
nand U27057 (N_27057,N_26524,N_26640);
nand U27058 (N_27058,N_26413,N_26679);
nor U27059 (N_27059,N_26982,N_26806);
nor U27060 (N_27060,N_26956,N_26544);
nand U27061 (N_27061,N_26659,N_26846);
nor U27062 (N_27062,N_26804,N_26492);
nor U27063 (N_27063,N_26672,N_26910);
nand U27064 (N_27064,N_26812,N_26741);
nor U27065 (N_27065,N_26687,N_26658);
and U27066 (N_27066,N_26882,N_26881);
or U27067 (N_27067,N_26944,N_26797);
or U27068 (N_27068,N_26734,N_26926);
and U27069 (N_27069,N_26995,N_26872);
or U27070 (N_27070,N_26432,N_26557);
nor U27071 (N_27071,N_26616,N_26404);
xor U27072 (N_27072,N_26918,N_26450);
nand U27073 (N_27073,N_26919,N_26403);
nor U27074 (N_27074,N_26438,N_26803);
and U27075 (N_27075,N_26972,N_26930);
nor U27076 (N_27076,N_26661,N_26990);
nor U27077 (N_27077,N_26729,N_26993);
nand U27078 (N_27078,N_26624,N_26907);
xor U27079 (N_27079,N_26895,N_26771);
or U27080 (N_27080,N_26665,N_26580);
nand U27081 (N_27081,N_26482,N_26773);
xor U27082 (N_27082,N_26629,N_26826);
and U27083 (N_27083,N_26466,N_26637);
or U27084 (N_27084,N_26699,N_26541);
xor U27085 (N_27085,N_26772,N_26615);
or U27086 (N_27086,N_26840,N_26951);
nand U27087 (N_27087,N_26457,N_26927);
and U27088 (N_27088,N_26923,N_26938);
xor U27089 (N_27089,N_26788,N_26538);
xor U27090 (N_27090,N_26418,N_26836);
or U27091 (N_27091,N_26948,N_26776);
nand U27092 (N_27092,N_26829,N_26791);
nor U27093 (N_27093,N_26675,N_26407);
nand U27094 (N_27094,N_26832,N_26628);
nor U27095 (N_27095,N_26702,N_26412);
nand U27096 (N_27096,N_26543,N_26724);
nand U27097 (N_27097,N_26817,N_26610);
or U27098 (N_27098,N_26400,N_26931);
nor U27099 (N_27099,N_26921,N_26572);
or U27100 (N_27100,N_26770,N_26861);
xnor U27101 (N_27101,N_26455,N_26475);
and U27102 (N_27102,N_26901,N_26958);
nand U27103 (N_27103,N_26973,N_26857);
nand U27104 (N_27104,N_26448,N_26978);
nor U27105 (N_27105,N_26553,N_26991);
xor U27106 (N_27106,N_26650,N_26587);
nand U27107 (N_27107,N_26467,N_26745);
xor U27108 (N_27108,N_26845,N_26565);
or U27109 (N_27109,N_26472,N_26505);
or U27110 (N_27110,N_26674,N_26979);
and U27111 (N_27111,N_26660,N_26528);
nand U27112 (N_27112,N_26914,N_26822);
xnor U27113 (N_27113,N_26983,N_26521);
nor U27114 (N_27114,N_26540,N_26796);
xnor U27115 (N_27115,N_26647,N_26798);
or U27116 (N_27116,N_26906,N_26811);
or U27117 (N_27117,N_26405,N_26549);
nand U27118 (N_27118,N_26755,N_26483);
or U27119 (N_27119,N_26639,N_26986);
or U27120 (N_27120,N_26815,N_26761);
and U27121 (N_27121,N_26415,N_26430);
and U27122 (N_27122,N_26608,N_26487);
or U27123 (N_27123,N_26760,N_26558);
nand U27124 (N_27124,N_26689,N_26463);
and U27125 (N_27125,N_26904,N_26607);
xnor U27126 (N_27126,N_26436,N_26497);
and U27127 (N_27127,N_26456,N_26622);
and U27128 (N_27128,N_26529,N_26446);
or U27129 (N_27129,N_26915,N_26725);
nand U27130 (N_27130,N_26708,N_26439);
nor U27131 (N_27131,N_26664,N_26425);
nor U27132 (N_27132,N_26518,N_26525);
or U27133 (N_27133,N_26480,N_26852);
and U27134 (N_27134,N_26410,N_26943);
and U27135 (N_27135,N_26417,N_26908);
and U27136 (N_27136,N_26484,N_26636);
nand U27137 (N_27137,N_26539,N_26617);
nand U27138 (N_27138,N_26913,N_26676);
and U27139 (N_27139,N_26747,N_26526);
nand U27140 (N_27140,N_26739,N_26824);
nand U27141 (N_27141,N_26563,N_26715);
or U27142 (N_27142,N_26733,N_26584);
nand U27143 (N_27143,N_26987,N_26641);
nor U27144 (N_27144,N_26460,N_26774);
xnor U27145 (N_27145,N_26427,N_26855);
nor U27146 (N_27146,N_26612,N_26648);
and U27147 (N_27147,N_26793,N_26769);
nand U27148 (N_27148,N_26989,N_26833);
or U27149 (N_27149,N_26988,N_26534);
and U27150 (N_27150,N_26547,N_26428);
or U27151 (N_27151,N_26691,N_26821);
or U27152 (N_27152,N_26856,N_26499);
nor U27153 (N_27153,N_26700,N_26655);
nor U27154 (N_27154,N_26935,N_26451);
and U27155 (N_27155,N_26513,N_26876);
and U27156 (N_27156,N_26794,N_26479);
nor U27157 (N_27157,N_26727,N_26414);
and U27158 (N_27158,N_26596,N_26925);
nand U27159 (N_27159,N_26704,N_26985);
nor U27160 (N_27160,N_26858,N_26928);
nand U27161 (N_27161,N_26564,N_26865);
nor U27162 (N_27162,N_26723,N_26609);
nor U27163 (N_27163,N_26952,N_26514);
and U27164 (N_27164,N_26442,N_26728);
nand U27165 (N_27165,N_26490,N_26570);
xnor U27166 (N_27166,N_26537,N_26644);
and U27167 (N_27167,N_26517,N_26884);
or U27168 (N_27168,N_26671,N_26940);
and U27169 (N_27169,N_26789,N_26933);
nor U27170 (N_27170,N_26885,N_26476);
and U27171 (N_27171,N_26718,N_26566);
nor U27172 (N_27172,N_26530,N_26732);
nand U27173 (N_27173,N_26562,N_26523);
nand U27174 (N_27174,N_26813,N_26437);
xor U27175 (N_27175,N_26696,N_26621);
nor U27176 (N_27176,N_26503,N_26519);
xor U27177 (N_27177,N_26942,N_26408);
nand U27178 (N_27178,N_26520,N_26916);
and U27179 (N_27179,N_26426,N_26962);
xor U27180 (N_27180,N_26831,N_26809);
and U27181 (N_27181,N_26611,N_26626);
nand U27182 (N_27182,N_26742,N_26920);
and U27183 (N_27183,N_26567,N_26712);
nor U27184 (N_27184,N_26875,N_26841);
nor U27185 (N_27185,N_26738,N_26898);
xnor U27186 (N_27186,N_26894,N_26512);
nand U27187 (N_27187,N_26502,N_26588);
nand U27188 (N_27188,N_26980,N_26957);
and U27189 (N_27189,N_26975,N_26453);
xnor U27190 (N_27190,N_26743,N_26556);
nand U27191 (N_27191,N_26606,N_26835);
and U27192 (N_27192,N_26863,N_26625);
or U27193 (N_27193,N_26545,N_26561);
nand U27194 (N_27194,N_26932,N_26792);
or U27195 (N_27195,N_26896,N_26554);
xnor U27196 (N_27196,N_26879,N_26779);
nor U27197 (N_27197,N_26527,N_26934);
xnor U27198 (N_27198,N_26871,N_26652);
nor U27199 (N_27199,N_26716,N_26878);
nor U27200 (N_27200,N_26864,N_26941);
or U27201 (N_27201,N_26516,N_26905);
nor U27202 (N_27202,N_26464,N_26577);
nor U27203 (N_27203,N_26657,N_26510);
nor U27204 (N_27204,N_26830,N_26713);
and U27205 (N_27205,N_26709,N_26486);
and U27206 (N_27206,N_26646,N_26736);
nand U27207 (N_27207,N_26471,N_26850);
and U27208 (N_27208,N_26869,N_26452);
nand U27209 (N_27209,N_26731,N_26862);
nor U27210 (N_27210,N_26690,N_26508);
or U27211 (N_27211,N_26695,N_26902);
and U27212 (N_27212,N_26586,N_26746);
and U27213 (N_27213,N_26900,N_26535);
and U27214 (N_27214,N_26802,N_26692);
nand U27215 (N_27215,N_26867,N_26842);
xor U27216 (N_27216,N_26478,N_26583);
xnor U27217 (N_27217,N_26574,N_26435);
xor U27218 (N_27218,N_26602,N_26468);
and U27219 (N_27219,N_26953,N_26751);
nand U27220 (N_27220,N_26550,N_26678);
xor U27221 (N_27221,N_26877,N_26633);
nor U27222 (N_27222,N_26423,N_26680);
and U27223 (N_27223,N_26735,N_26714);
xnor U27224 (N_27224,N_26964,N_26507);
or U27225 (N_27225,N_26801,N_26883);
nand U27226 (N_27226,N_26409,N_26994);
and U27227 (N_27227,N_26495,N_26568);
nor U27228 (N_27228,N_26892,N_26536);
nor U27229 (N_27229,N_26693,N_26592);
and U27230 (N_27230,N_26605,N_26684);
and U27231 (N_27231,N_26673,N_26837);
nor U27232 (N_27232,N_26462,N_26999);
nand U27233 (N_27233,N_26757,N_26571);
or U27234 (N_27234,N_26546,N_26825);
xnor U27235 (N_27235,N_26778,N_26685);
or U27236 (N_27236,N_26787,N_26981);
and U27237 (N_27237,N_26965,N_26763);
nand U27238 (N_27238,N_26929,N_26939);
xnor U27239 (N_27239,N_26424,N_26663);
nand U27240 (N_27240,N_26481,N_26711);
or U27241 (N_27241,N_26721,N_26814);
and U27242 (N_27242,N_26643,N_26860);
or U27243 (N_27243,N_26843,N_26810);
or U27244 (N_27244,N_26795,N_26496);
nand U27245 (N_27245,N_26461,N_26573);
nand U27246 (N_27246,N_26768,N_26694);
or U27247 (N_27247,N_26595,N_26669);
nor U27248 (N_27248,N_26786,N_26579);
nor U27249 (N_27249,N_26765,N_26630);
nor U27250 (N_27250,N_26859,N_26470);
and U27251 (N_27251,N_26866,N_26870);
nor U27252 (N_27252,N_26740,N_26970);
nand U27253 (N_27253,N_26880,N_26799);
or U27254 (N_27254,N_26465,N_26498);
xor U27255 (N_27255,N_26493,N_26838);
or U27256 (N_27256,N_26848,N_26954);
and U27257 (N_27257,N_26717,N_26839);
nor U27258 (N_27258,N_26618,N_26868);
or U27259 (N_27259,N_26851,N_26533);
nand U27260 (N_27260,N_26485,N_26597);
xnor U27261 (N_27261,N_26429,N_26911);
xor U27262 (N_27262,N_26955,N_26783);
or U27263 (N_27263,N_26960,N_26662);
nor U27264 (N_27264,N_26748,N_26720);
nor U27265 (N_27265,N_26903,N_26749);
and U27266 (N_27266,N_26781,N_26576);
nor U27267 (N_27267,N_26601,N_26827);
and U27268 (N_27268,N_26816,N_26703);
xor U27269 (N_27269,N_26614,N_26433);
nor U27270 (N_27270,N_26968,N_26402);
xor U27271 (N_27271,N_26849,N_26992);
or U27272 (N_27272,N_26726,N_26873);
and U27273 (N_27273,N_26589,N_26808);
and U27274 (N_27274,N_26936,N_26670);
or U27275 (N_27275,N_26766,N_26645);
nor U27276 (N_27276,N_26613,N_26784);
nand U27277 (N_27277,N_26627,N_26963);
nor U27278 (N_27278,N_26710,N_26431);
nand U27279 (N_27279,N_26780,N_26434);
nand U27280 (N_27280,N_26623,N_26705);
xor U27281 (N_27281,N_26619,N_26807);
nand U27282 (N_27282,N_26819,N_26912);
nor U27283 (N_27283,N_26551,N_26949);
xnor U27284 (N_27284,N_26656,N_26974);
nand U27285 (N_27285,N_26459,N_26491);
and U27286 (N_27286,N_26509,N_26701);
nor U27287 (N_27287,N_26635,N_26893);
or U27288 (N_27288,N_26593,N_26945);
xor U27289 (N_27289,N_26581,N_26706);
and U27290 (N_27290,N_26820,N_26511);
xor U27291 (N_27291,N_26421,N_26458);
xnor U27292 (N_27292,N_26844,N_26552);
nand U27293 (N_27293,N_26899,N_26937);
xnor U27294 (N_27294,N_26969,N_26800);
nand U27295 (N_27295,N_26823,N_26961);
xnor U27296 (N_27296,N_26419,N_26642);
or U27297 (N_27297,N_26443,N_26555);
nand U27298 (N_27298,N_26638,N_26976);
and U27299 (N_27299,N_26998,N_26854);
nor U27300 (N_27300,N_26765,N_26962);
nor U27301 (N_27301,N_26562,N_26486);
nor U27302 (N_27302,N_26975,N_26506);
nor U27303 (N_27303,N_26899,N_26670);
or U27304 (N_27304,N_26985,N_26562);
and U27305 (N_27305,N_26414,N_26595);
nand U27306 (N_27306,N_26686,N_26739);
or U27307 (N_27307,N_26797,N_26632);
or U27308 (N_27308,N_26909,N_26525);
or U27309 (N_27309,N_26829,N_26732);
xnor U27310 (N_27310,N_26424,N_26930);
and U27311 (N_27311,N_26566,N_26602);
and U27312 (N_27312,N_26875,N_26939);
xor U27313 (N_27313,N_26921,N_26613);
xor U27314 (N_27314,N_26971,N_26441);
and U27315 (N_27315,N_26790,N_26553);
nand U27316 (N_27316,N_26807,N_26409);
and U27317 (N_27317,N_26992,N_26560);
nor U27318 (N_27318,N_26829,N_26535);
and U27319 (N_27319,N_26713,N_26926);
or U27320 (N_27320,N_26997,N_26595);
nand U27321 (N_27321,N_26607,N_26418);
and U27322 (N_27322,N_26674,N_26848);
nor U27323 (N_27323,N_26531,N_26937);
or U27324 (N_27324,N_26903,N_26984);
and U27325 (N_27325,N_26808,N_26742);
nor U27326 (N_27326,N_26518,N_26991);
and U27327 (N_27327,N_26875,N_26586);
xnor U27328 (N_27328,N_26983,N_26924);
and U27329 (N_27329,N_26941,N_26448);
xnor U27330 (N_27330,N_26562,N_26745);
and U27331 (N_27331,N_26654,N_26844);
and U27332 (N_27332,N_26573,N_26718);
xor U27333 (N_27333,N_26724,N_26912);
and U27334 (N_27334,N_26707,N_26794);
xor U27335 (N_27335,N_26448,N_26813);
xor U27336 (N_27336,N_26693,N_26560);
or U27337 (N_27337,N_26433,N_26988);
and U27338 (N_27338,N_26872,N_26628);
nor U27339 (N_27339,N_26814,N_26529);
xnor U27340 (N_27340,N_26870,N_26458);
and U27341 (N_27341,N_26838,N_26871);
and U27342 (N_27342,N_26553,N_26662);
or U27343 (N_27343,N_26784,N_26856);
nor U27344 (N_27344,N_26897,N_26855);
xnor U27345 (N_27345,N_26531,N_26572);
xnor U27346 (N_27346,N_26828,N_26792);
nand U27347 (N_27347,N_26511,N_26936);
or U27348 (N_27348,N_26943,N_26657);
nor U27349 (N_27349,N_26769,N_26777);
and U27350 (N_27350,N_26413,N_26864);
xnor U27351 (N_27351,N_26976,N_26678);
and U27352 (N_27352,N_26976,N_26574);
nor U27353 (N_27353,N_26812,N_26994);
nor U27354 (N_27354,N_26897,N_26484);
and U27355 (N_27355,N_26814,N_26666);
xor U27356 (N_27356,N_26548,N_26429);
xor U27357 (N_27357,N_26714,N_26584);
nand U27358 (N_27358,N_26546,N_26648);
and U27359 (N_27359,N_26732,N_26686);
and U27360 (N_27360,N_26905,N_26642);
nor U27361 (N_27361,N_26743,N_26994);
xnor U27362 (N_27362,N_26482,N_26860);
nor U27363 (N_27363,N_26845,N_26744);
and U27364 (N_27364,N_26894,N_26750);
nand U27365 (N_27365,N_26603,N_26514);
xnor U27366 (N_27366,N_26800,N_26504);
nor U27367 (N_27367,N_26874,N_26544);
and U27368 (N_27368,N_26870,N_26693);
nor U27369 (N_27369,N_26914,N_26685);
or U27370 (N_27370,N_26897,N_26518);
nor U27371 (N_27371,N_26620,N_26409);
xor U27372 (N_27372,N_26757,N_26581);
or U27373 (N_27373,N_26841,N_26449);
xor U27374 (N_27374,N_26482,N_26790);
nor U27375 (N_27375,N_26438,N_26605);
and U27376 (N_27376,N_26507,N_26641);
xnor U27377 (N_27377,N_26829,N_26751);
or U27378 (N_27378,N_26912,N_26755);
nor U27379 (N_27379,N_26805,N_26706);
and U27380 (N_27380,N_26979,N_26621);
nand U27381 (N_27381,N_26949,N_26704);
and U27382 (N_27382,N_26551,N_26720);
xor U27383 (N_27383,N_26463,N_26904);
nor U27384 (N_27384,N_26548,N_26574);
or U27385 (N_27385,N_26434,N_26952);
xnor U27386 (N_27386,N_26818,N_26693);
nand U27387 (N_27387,N_26828,N_26763);
nand U27388 (N_27388,N_26694,N_26644);
or U27389 (N_27389,N_26547,N_26551);
nand U27390 (N_27390,N_26480,N_26954);
nor U27391 (N_27391,N_26419,N_26635);
nor U27392 (N_27392,N_26791,N_26709);
xor U27393 (N_27393,N_26896,N_26464);
and U27394 (N_27394,N_26447,N_26738);
nor U27395 (N_27395,N_26651,N_26712);
or U27396 (N_27396,N_26678,N_26559);
xor U27397 (N_27397,N_26772,N_26614);
xor U27398 (N_27398,N_26938,N_26446);
nand U27399 (N_27399,N_26518,N_26846);
xor U27400 (N_27400,N_26472,N_26817);
nand U27401 (N_27401,N_26734,N_26996);
nor U27402 (N_27402,N_26410,N_26492);
nor U27403 (N_27403,N_26910,N_26706);
nor U27404 (N_27404,N_26581,N_26872);
nand U27405 (N_27405,N_26977,N_26446);
nand U27406 (N_27406,N_26957,N_26842);
or U27407 (N_27407,N_26814,N_26973);
or U27408 (N_27408,N_26722,N_26826);
nand U27409 (N_27409,N_26927,N_26525);
nand U27410 (N_27410,N_26425,N_26886);
nand U27411 (N_27411,N_26576,N_26673);
or U27412 (N_27412,N_26537,N_26760);
nand U27413 (N_27413,N_26596,N_26684);
or U27414 (N_27414,N_26593,N_26655);
nand U27415 (N_27415,N_26543,N_26640);
and U27416 (N_27416,N_26977,N_26675);
and U27417 (N_27417,N_26539,N_26521);
nand U27418 (N_27418,N_26703,N_26760);
or U27419 (N_27419,N_26796,N_26621);
or U27420 (N_27420,N_26493,N_26565);
and U27421 (N_27421,N_26831,N_26524);
or U27422 (N_27422,N_26977,N_26753);
or U27423 (N_27423,N_26723,N_26447);
nand U27424 (N_27424,N_26838,N_26790);
xnor U27425 (N_27425,N_26421,N_26947);
nand U27426 (N_27426,N_26925,N_26595);
nor U27427 (N_27427,N_26928,N_26671);
or U27428 (N_27428,N_26534,N_26927);
and U27429 (N_27429,N_26996,N_26586);
and U27430 (N_27430,N_26840,N_26844);
xnor U27431 (N_27431,N_26614,N_26599);
xnor U27432 (N_27432,N_26950,N_26512);
and U27433 (N_27433,N_26964,N_26626);
or U27434 (N_27434,N_26851,N_26527);
xor U27435 (N_27435,N_26444,N_26721);
nand U27436 (N_27436,N_26993,N_26544);
nand U27437 (N_27437,N_26427,N_26453);
nand U27438 (N_27438,N_26805,N_26836);
nor U27439 (N_27439,N_26997,N_26789);
and U27440 (N_27440,N_26491,N_26541);
xor U27441 (N_27441,N_26773,N_26919);
nand U27442 (N_27442,N_26754,N_26672);
nor U27443 (N_27443,N_26795,N_26919);
nand U27444 (N_27444,N_26777,N_26929);
xor U27445 (N_27445,N_26985,N_26846);
or U27446 (N_27446,N_26648,N_26913);
nor U27447 (N_27447,N_26877,N_26430);
nand U27448 (N_27448,N_26742,N_26890);
and U27449 (N_27449,N_26720,N_26654);
nor U27450 (N_27450,N_26519,N_26886);
or U27451 (N_27451,N_26402,N_26625);
xor U27452 (N_27452,N_26447,N_26863);
xor U27453 (N_27453,N_26581,N_26430);
xor U27454 (N_27454,N_26901,N_26513);
or U27455 (N_27455,N_26965,N_26796);
nand U27456 (N_27456,N_26463,N_26808);
or U27457 (N_27457,N_26788,N_26729);
nand U27458 (N_27458,N_26486,N_26403);
xor U27459 (N_27459,N_26982,N_26793);
nand U27460 (N_27460,N_26650,N_26631);
and U27461 (N_27461,N_26518,N_26406);
nor U27462 (N_27462,N_26632,N_26986);
and U27463 (N_27463,N_26881,N_26775);
or U27464 (N_27464,N_26746,N_26447);
nor U27465 (N_27465,N_26994,N_26656);
nor U27466 (N_27466,N_26604,N_26522);
xnor U27467 (N_27467,N_26834,N_26548);
nand U27468 (N_27468,N_26577,N_26812);
nand U27469 (N_27469,N_26899,N_26526);
nand U27470 (N_27470,N_26945,N_26676);
and U27471 (N_27471,N_26685,N_26835);
or U27472 (N_27472,N_26889,N_26566);
and U27473 (N_27473,N_26608,N_26821);
and U27474 (N_27474,N_26919,N_26575);
xor U27475 (N_27475,N_26895,N_26476);
or U27476 (N_27476,N_26903,N_26797);
nor U27477 (N_27477,N_26411,N_26929);
or U27478 (N_27478,N_26589,N_26815);
nand U27479 (N_27479,N_26917,N_26855);
or U27480 (N_27480,N_26950,N_26428);
nor U27481 (N_27481,N_26962,N_26508);
and U27482 (N_27482,N_26894,N_26640);
nand U27483 (N_27483,N_26863,N_26785);
nand U27484 (N_27484,N_26679,N_26631);
xnor U27485 (N_27485,N_26659,N_26622);
or U27486 (N_27486,N_26815,N_26881);
or U27487 (N_27487,N_26752,N_26425);
xnor U27488 (N_27488,N_26476,N_26922);
nor U27489 (N_27489,N_26571,N_26864);
or U27490 (N_27490,N_26413,N_26700);
and U27491 (N_27491,N_26649,N_26784);
or U27492 (N_27492,N_26942,N_26765);
xnor U27493 (N_27493,N_26630,N_26404);
nor U27494 (N_27494,N_26950,N_26602);
or U27495 (N_27495,N_26855,N_26509);
xor U27496 (N_27496,N_26550,N_26735);
or U27497 (N_27497,N_26485,N_26818);
and U27498 (N_27498,N_26901,N_26663);
nand U27499 (N_27499,N_26666,N_26993);
and U27500 (N_27500,N_26528,N_26562);
xor U27501 (N_27501,N_26448,N_26663);
or U27502 (N_27502,N_26588,N_26613);
and U27503 (N_27503,N_26606,N_26434);
xor U27504 (N_27504,N_26943,N_26951);
nand U27505 (N_27505,N_26756,N_26527);
xor U27506 (N_27506,N_26558,N_26953);
xnor U27507 (N_27507,N_26855,N_26850);
nand U27508 (N_27508,N_26519,N_26884);
or U27509 (N_27509,N_26692,N_26499);
and U27510 (N_27510,N_26933,N_26976);
xor U27511 (N_27511,N_26431,N_26542);
nand U27512 (N_27512,N_26434,N_26890);
or U27513 (N_27513,N_26725,N_26769);
or U27514 (N_27514,N_26863,N_26546);
nand U27515 (N_27515,N_26939,N_26958);
nand U27516 (N_27516,N_26706,N_26640);
nor U27517 (N_27517,N_26691,N_26938);
xnor U27518 (N_27518,N_26584,N_26968);
nor U27519 (N_27519,N_26428,N_26587);
or U27520 (N_27520,N_26781,N_26495);
nor U27521 (N_27521,N_26818,N_26681);
and U27522 (N_27522,N_26823,N_26506);
xor U27523 (N_27523,N_26863,N_26869);
nand U27524 (N_27524,N_26561,N_26759);
xnor U27525 (N_27525,N_26520,N_26565);
xor U27526 (N_27526,N_26854,N_26618);
nor U27527 (N_27527,N_26866,N_26821);
xnor U27528 (N_27528,N_26958,N_26676);
nand U27529 (N_27529,N_26549,N_26924);
nor U27530 (N_27530,N_26596,N_26469);
and U27531 (N_27531,N_26596,N_26863);
and U27532 (N_27532,N_26989,N_26760);
and U27533 (N_27533,N_26737,N_26671);
nor U27534 (N_27534,N_26617,N_26411);
nand U27535 (N_27535,N_26414,N_26580);
nor U27536 (N_27536,N_26562,N_26636);
or U27537 (N_27537,N_26936,N_26541);
xnor U27538 (N_27538,N_26604,N_26942);
xnor U27539 (N_27539,N_26597,N_26621);
and U27540 (N_27540,N_26797,N_26544);
xnor U27541 (N_27541,N_26423,N_26961);
or U27542 (N_27542,N_26526,N_26898);
xor U27543 (N_27543,N_26838,N_26476);
xnor U27544 (N_27544,N_26852,N_26701);
or U27545 (N_27545,N_26447,N_26939);
or U27546 (N_27546,N_26498,N_26404);
or U27547 (N_27547,N_26921,N_26644);
or U27548 (N_27548,N_26916,N_26567);
or U27549 (N_27549,N_26621,N_26912);
and U27550 (N_27550,N_26448,N_26550);
nand U27551 (N_27551,N_26606,N_26774);
or U27552 (N_27552,N_26828,N_26557);
and U27553 (N_27553,N_26528,N_26828);
or U27554 (N_27554,N_26589,N_26782);
and U27555 (N_27555,N_26489,N_26640);
or U27556 (N_27556,N_26996,N_26454);
nand U27557 (N_27557,N_26734,N_26506);
nor U27558 (N_27558,N_26627,N_26891);
nand U27559 (N_27559,N_26712,N_26996);
nor U27560 (N_27560,N_26507,N_26847);
nand U27561 (N_27561,N_26784,N_26474);
nand U27562 (N_27562,N_26609,N_26993);
nor U27563 (N_27563,N_26483,N_26716);
or U27564 (N_27564,N_26849,N_26703);
and U27565 (N_27565,N_26683,N_26837);
or U27566 (N_27566,N_26541,N_26564);
nor U27567 (N_27567,N_26458,N_26737);
nor U27568 (N_27568,N_26999,N_26532);
nor U27569 (N_27569,N_26791,N_26703);
nor U27570 (N_27570,N_26408,N_26548);
nor U27571 (N_27571,N_26929,N_26713);
nand U27572 (N_27572,N_26841,N_26952);
nand U27573 (N_27573,N_26991,N_26985);
nor U27574 (N_27574,N_26636,N_26916);
nor U27575 (N_27575,N_26805,N_26727);
nand U27576 (N_27576,N_26930,N_26625);
or U27577 (N_27577,N_26541,N_26456);
or U27578 (N_27578,N_26920,N_26443);
or U27579 (N_27579,N_26708,N_26456);
xnor U27580 (N_27580,N_26740,N_26442);
nor U27581 (N_27581,N_26438,N_26475);
nor U27582 (N_27582,N_26647,N_26778);
or U27583 (N_27583,N_26739,N_26841);
or U27584 (N_27584,N_26790,N_26919);
and U27585 (N_27585,N_26897,N_26913);
nor U27586 (N_27586,N_26550,N_26429);
nand U27587 (N_27587,N_26920,N_26881);
xnor U27588 (N_27588,N_26991,N_26629);
xor U27589 (N_27589,N_26962,N_26621);
nor U27590 (N_27590,N_26622,N_26821);
xor U27591 (N_27591,N_26570,N_26776);
and U27592 (N_27592,N_26431,N_26925);
xor U27593 (N_27593,N_26555,N_26934);
or U27594 (N_27594,N_26697,N_26799);
or U27595 (N_27595,N_26421,N_26648);
and U27596 (N_27596,N_26939,N_26863);
nor U27597 (N_27597,N_26599,N_26752);
or U27598 (N_27598,N_26815,N_26440);
or U27599 (N_27599,N_26892,N_26474);
nand U27600 (N_27600,N_27309,N_27046);
nor U27601 (N_27601,N_27334,N_27428);
nand U27602 (N_27602,N_27330,N_27347);
xnor U27603 (N_27603,N_27335,N_27114);
and U27604 (N_27604,N_27265,N_27413);
xnor U27605 (N_27605,N_27587,N_27386);
and U27606 (N_27606,N_27368,N_27180);
xor U27607 (N_27607,N_27344,N_27465);
and U27608 (N_27608,N_27138,N_27302);
nand U27609 (N_27609,N_27203,N_27132);
or U27610 (N_27610,N_27201,N_27189);
xor U27611 (N_27611,N_27224,N_27153);
and U27612 (N_27612,N_27495,N_27359);
nor U27613 (N_27613,N_27425,N_27556);
xor U27614 (N_27614,N_27086,N_27356);
or U27615 (N_27615,N_27107,N_27374);
xnor U27616 (N_27616,N_27006,N_27575);
and U27617 (N_27617,N_27526,N_27393);
and U27618 (N_27618,N_27295,N_27226);
or U27619 (N_27619,N_27118,N_27555);
or U27620 (N_27620,N_27594,N_27277);
nor U27621 (N_27621,N_27026,N_27510);
nand U27622 (N_27622,N_27025,N_27324);
and U27623 (N_27623,N_27409,N_27089);
and U27624 (N_27624,N_27035,N_27476);
or U27625 (N_27625,N_27582,N_27112);
nand U27626 (N_27626,N_27363,N_27452);
xnor U27627 (N_27627,N_27167,N_27438);
or U27628 (N_27628,N_27401,N_27172);
nor U27629 (N_27629,N_27162,N_27319);
or U27630 (N_27630,N_27375,N_27539);
or U27631 (N_27631,N_27494,N_27047);
and U27632 (N_27632,N_27420,N_27216);
xnor U27633 (N_27633,N_27151,N_27155);
nand U27634 (N_27634,N_27503,N_27337);
xnor U27635 (N_27635,N_27514,N_27084);
xnor U27636 (N_27636,N_27061,N_27546);
nand U27637 (N_27637,N_27161,N_27573);
xnor U27638 (N_27638,N_27507,N_27541);
and U27639 (N_27639,N_27257,N_27268);
or U27640 (N_27640,N_27345,N_27398);
and U27641 (N_27641,N_27190,N_27444);
and U27642 (N_27642,N_27000,N_27517);
and U27643 (N_27643,N_27327,N_27414);
and U27644 (N_27644,N_27412,N_27518);
nand U27645 (N_27645,N_27157,N_27031);
nor U27646 (N_27646,N_27014,N_27017);
nand U27647 (N_27647,N_27247,N_27264);
and U27648 (N_27648,N_27463,N_27097);
xnor U27649 (N_27649,N_27562,N_27131);
nand U27650 (N_27650,N_27559,N_27547);
nor U27651 (N_27651,N_27099,N_27271);
nand U27652 (N_27652,N_27236,N_27055);
nor U27653 (N_27653,N_27064,N_27049);
or U27654 (N_27654,N_27288,N_27280);
or U27655 (N_27655,N_27571,N_27037);
nand U27656 (N_27656,N_27360,N_27551);
nor U27657 (N_27657,N_27235,N_27001);
or U27658 (N_27658,N_27152,N_27544);
nand U27659 (N_27659,N_27584,N_27377);
nand U27660 (N_27660,N_27147,N_27029);
xor U27661 (N_27661,N_27455,N_27230);
and U27662 (N_27662,N_27273,N_27536);
xor U27663 (N_27663,N_27053,N_27593);
and U27664 (N_27664,N_27490,N_27456);
nand U27665 (N_27665,N_27419,N_27183);
or U27666 (N_27666,N_27116,N_27169);
nor U27667 (N_27667,N_27072,N_27125);
xnor U27668 (N_27668,N_27239,N_27210);
or U27669 (N_27669,N_27383,N_27486);
nor U27670 (N_27670,N_27437,N_27340);
xnor U27671 (N_27671,N_27290,N_27382);
nand U27672 (N_27672,N_27417,N_27069);
and U27673 (N_27673,N_27148,N_27208);
nor U27674 (N_27674,N_27166,N_27480);
nand U27675 (N_27675,N_27580,N_27322);
nand U27676 (N_27676,N_27243,N_27133);
xnor U27677 (N_27677,N_27044,N_27156);
or U27678 (N_27678,N_27149,N_27198);
nand U27679 (N_27679,N_27042,N_27548);
or U27680 (N_27680,N_27205,N_27472);
and U27681 (N_27681,N_27531,N_27564);
or U27682 (N_27682,N_27193,N_27371);
nand U27683 (N_27683,N_27135,N_27079);
or U27684 (N_27684,N_27105,N_27569);
or U27685 (N_27685,N_27498,N_27574);
nand U27686 (N_27686,N_27202,N_27396);
or U27687 (N_27687,N_27350,N_27355);
and U27688 (N_27688,N_27276,N_27123);
and U27689 (N_27689,N_27188,N_27098);
nor U27690 (N_27690,N_27073,N_27174);
and U27691 (N_27691,N_27050,N_27275);
nor U27692 (N_27692,N_27246,N_27397);
nor U27693 (N_27693,N_27181,N_27540);
nand U27694 (N_27694,N_27286,N_27285);
nand U27695 (N_27695,N_27364,N_27365);
and U27696 (N_27696,N_27033,N_27457);
nor U27697 (N_27697,N_27379,N_27165);
xnor U27698 (N_27698,N_27178,N_27328);
xor U27699 (N_27699,N_27010,N_27292);
xor U27700 (N_27700,N_27576,N_27008);
or U27701 (N_27701,N_27291,N_27483);
xor U27702 (N_27702,N_27361,N_27093);
nand U27703 (N_27703,N_27372,N_27145);
and U27704 (N_27704,N_27535,N_27598);
xnor U27705 (N_27705,N_27595,N_27012);
xor U27706 (N_27706,N_27134,N_27523);
nand U27707 (N_27707,N_27308,N_27212);
and U27708 (N_27708,N_27176,N_27300);
xor U27709 (N_27709,N_27170,N_27113);
nor U27710 (N_27710,N_27206,N_27222);
xnor U27711 (N_27711,N_27101,N_27357);
nand U27712 (N_27712,N_27082,N_27023);
nand U27713 (N_27713,N_27248,N_27043);
and U27714 (N_27714,N_27532,N_27108);
nand U27715 (N_27715,N_27599,N_27088);
nor U27716 (N_27716,N_27519,N_27392);
or U27717 (N_27717,N_27109,N_27331);
and U27718 (N_27718,N_27056,N_27515);
or U27719 (N_27719,N_27126,N_27561);
or U27720 (N_27720,N_27045,N_27467);
xnor U27721 (N_27721,N_27525,N_27445);
and U27722 (N_27722,N_27410,N_27094);
xor U27723 (N_27723,N_27404,N_27423);
or U27724 (N_27724,N_27120,N_27032);
xnor U27725 (N_27725,N_27034,N_27085);
and U27726 (N_27726,N_27278,N_27381);
xnor U27727 (N_27727,N_27092,N_27543);
nor U27728 (N_27728,N_27020,N_27421);
nor U27729 (N_27729,N_27550,N_27127);
nor U27730 (N_27730,N_27237,N_27245);
and U27731 (N_27731,N_27004,N_27339);
or U27732 (N_27732,N_27013,N_27373);
nor U27733 (N_27733,N_27468,N_27348);
nor U27734 (N_27734,N_27279,N_27513);
and U27735 (N_27735,N_27447,N_27542);
or U27736 (N_27736,N_27469,N_27333);
or U27737 (N_27737,N_27301,N_27549);
and U27738 (N_27738,N_27454,N_27362);
or U27739 (N_27739,N_27287,N_27493);
xor U27740 (N_27740,N_27553,N_27171);
xor U27741 (N_27741,N_27378,N_27427);
and U27742 (N_27742,N_27065,N_27080);
and U27743 (N_27743,N_27225,N_27563);
nand U27744 (N_27744,N_27238,N_27242);
nor U27745 (N_27745,N_27411,N_27433);
nor U27746 (N_27746,N_27117,N_27284);
and U27747 (N_27747,N_27102,N_27527);
nand U27748 (N_27748,N_27255,N_27592);
nor U27749 (N_27749,N_27234,N_27137);
nor U27750 (N_27750,N_27538,N_27529);
xnor U27751 (N_27751,N_27311,N_27260);
nand U27752 (N_27752,N_27177,N_27095);
and U27753 (N_27753,N_27314,N_27263);
xor U27754 (N_27754,N_27520,N_27002);
xor U27755 (N_27755,N_27070,N_27482);
and U27756 (N_27756,N_27103,N_27293);
xnor U27757 (N_27757,N_27464,N_27254);
nor U27758 (N_27758,N_27076,N_27441);
nor U27759 (N_27759,N_27213,N_27481);
or U27760 (N_27760,N_27121,N_27349);
and U27761 (N_27761,N_27192,N_27390);
nand U27762 (N_27762,N_27321,N_27475);
and U27763 (N_27763,N_27566,N_27142);
nor U27764 (N_27764,N_27430,N_27304);
nand U27765 (N_27765,N_27141,N_27380);
xnor U27766 (N_27766,N_27228,N_27122);
or U27767 (N_27767,N_27415,N_27274);
nor U27768 (N_27768,N_27015,N_27077);
and U27769 (N_27769,N_27496,N_27596);
nor U27770 (N_27770,N_27497,N_27241);
and U27771 (N_27771,N_27506,N_27219);
or U27772 (N_27772,N_27450,N_27351);
and U27773 (N_27773,N_27261,N_27154);
xor U27774 (N_27774,N_27159,N_27303);
nor U27775 (N_27775,N_27585,N_27590);
and U27776 (N_27776,N_27283,N_27106);
nor U27777 (N_27777,N_27338,N_27066);
nand U27778 (N_27778,N_27466,N_27139);
nand U27779 (N_27779,N_27136,N_27318);
nor U27780 (N_27780,N_27353,N_27028);
xor U27781 (N_27781,N_27146,N_27583);
xor U27782 (N_27782,N_27018,N_27578);
nand U27783 (N_27783,N_27389,N_27063);
xnor U27784 (N_27784,N_27403,N_27346);
xor U27785 (N_27785,N_27299,N_27453);
and U27786 (N_27786,N_27185,N_27220);
or U27787 (N_27787,N_27129,N_27431);
and U27788 (N_27788,N_27267,N_27075);
and U27789 (N_27789,N_27168,N_27232);
nor U27790 (N_27790,N_27173,N_27565);
or U27791 (N_27791,N_27024,N_27163);
nand U27792 (N_27792,N_27272,N_27187);
nand U27793 (N_27793,N_27416,N_27019);
nor U27794 (N_27794,N_27579,N_27376);
xnor U27795 (N_27795,N_27270,N_27227);
nor U27796 (N_27796,N_27387,N_27048);
nor U27797 (N_27797,N_27458,N_27307);
and U27798 (N_27798,N_27317,N_27196);
xnor U27799 (N_27799,N_27577,N_27312);
or U27800 (N_27800,N_27492,N_27477);
nor U27801 (N_27801,N_27186,N_27289);
nand U27802 (N_27802,N_27552,N_27516);
or U27803 (N_27803,N_27557,N_27060);
or U27804 (N_27804,N_27104,N_27195);
xor U27805 (N_27805,N_27144,N_27325);
xnor U27806 (N_27806,N_27435,N_27266);
and U27807 (N_27807,N_27009,N_27408);
and U27808 (N_27808,N_27229,N_27570);
nor U27809 (N_27809,N_27459,N_27487);
and U27810 (N_27810,N_27588,N_27367);
nand U27811 (N_27811,N_27568,N_27119);
xnor U27812 (N_27812,N_27252,N_27011);
nor U27813 (N_27813,N_27460,N_27394);
xor U27814 (N_27814,N_27537,N_27038);
nand U27815 (N_27815,N_27491,N_27111);
and U27816 (N_27816,N_27258,N_27343);
and U27817 (N_27817,N_27407,N_27062);
or U27818 (N_27818,N_27215,N_27310);
nor U27819 (N_27819,N_27511,N_27436);
or U27820 (N_27820,N_27479,N_27130);
or U27821 (N_27821,N_27326,N_27016);
nand U27822 (N_27822,N_27096,N_27067);
xnor U27823 (N_27823,N_27354,N_27499);
nor U27824 (N_27824,N_27432,N_27399);
nor U27825 (N_27825,N_27140,N_27058);
and U27826 (N_27826,N_27451,N_27110);
and U27827 (N_27827,N_27059,N_27589);
nor U27828 (N_27828,N_27439,N_27211);
nor U27829 (N_27829,N_27504,N_27298);
or U27830 (N_27830,N_27164,N_27244);
and U27831 (N_27831,N_27449,N_27484);
nand U27832 (N_27832,N_27395,N_27448);
nand U27833 (N_27833,N_27091,N_27488);
nor U27834 (N_27834,N_27221,N_27259);
nand U27835 (N_27835,N_27081,N_27087);
and U27836 (N_27836,N_27027,N_27030);
nand U27837 (N_27837,N_27384,N_27336);
and U27838 (N_27838,N_27533,N_27184);
or U27839 (N_27839,N_27315,N_27528);
nand U27840 (N_27840,N_27402,N_27200);
nand U27841 (N_27841,N_27316,N_27100);
nor U27842 (N_27842,N_27470,N_27332);
and U27843 (N_27843,N_27068,N_27158);
nor U27844 (N_27844,N_27545,N_27231);
or U27845 (N_27845,N_27406,N_27143);
nor U27846 (N_27846,N_27461,N_27296);
nor U27847 (N_27847,N_27352,N_27071);
xnor U27848 (N_27848,N_27567,N_27007);
and U27849 (N_27849,N_27240,N_27204);
xor U27850 (N_27850,N_27305,N_27366);
xnor U27851 (N_27851,N_27249,N_27442);
nor U27852 (N_27852,N_27251,N_27209);
nand U27853 (N_27853,N_27485,N_27446);
xor U27854 (N_27854,N_27558,N_27306);
nor U27855 (N_27855,N_27489,N_27036);
nor U27856 (N_27856,N_27021,N_27074);
or U27857 (N_27857,N_27294,N_27179);
nand U27858 (N_27858,N_27385,N_27253);
nand U27859 (N_27859,N_27509,N_27057);
xor U27860 (N_27860,N_27040,N_27313);
nand U27861 (N_27861,N_27051,N_27281);
and U27862 (N_27862,N_27426,N_27003);
nor U27863 (N_27863,N_27591,N_27521);
nand U27864 (N_27864,N_27572,N_27052);
nor U27865 (N_27865,N_27124,N_27522);
xor U27866 (N_27866,N_27250,N_27524);
or U27867 (N_27867,N_27217,N_27090);
nor U27868 (N_27868,N_27505,N_27083);
and U27869 (N_27869,N_27478,N_27197);
nand U27870 (N_27870,N_27500,N_27440);
nand U27871 (N_27871,N_27370,N_27434);
and U27872 (N_27872,N_27422,N_27022);
and U27873 (N_27873,N_27369,N_27429);
nor U27874 (N_27874,N_27388,N_27473);
xnor U27875 (N_27875,N_27508,N_27041);
and U27876 (N_27876,N_27218,N_27391);
and U27877 (N_27877,N_27424,N_27256);
nand U27878 (N_27878,N_27501,N_27586);
and U27879 (N_27879,N_27358,N_27554);
nor U27880 (N_27880,N_27214,N_27512);
or U27881 (N_27881,N_27262,N_27182);
nor U27882 (N_27882,N_27005,N_27342);
xor U27883 (N_27883,N_27534,N_27128);
or U27884 (N_27884,N_27329,N_27530);
nor U27885 (N_27885,N_27269,N_27323);
xnor U27886 (N_27886,N_27405,N_27474);
xnor U27887 (N_27887,N_27297,N_27560);
nor U27888 (N_27888,N_27115,N_27400);
xor U27889 (N_27889,N_27223,N_27320);
nor U27890 (N_27890,N_27462,N_27443);
nand U27891 (N_27891,N_27282,N_27502);
nand U27892 (N_27892,N_27194,N_27039);
nand U27893 (N_27893,N_27471,N_27581);
nand U27894 (N_27894,N_27418,N_27199);
and U27895 (N_27895,N_27078,N_27207);
nand U27896 (N_27896,N_27233,N_27150);
or U27897 (N_27897,N_27160,N_27597);
and U27898 (N_27898,N_27054,N_27341);
or U27899 (N_27899,N_27191,N_27175);
or U27900 (N_27900,N_27012,N_27374);
nand U27901 (N_27901,N_27233,N_27228);
nand U27902 (N_27902,N_27558,N_27590);
nand U27903 (N_27903,N_27129,N_27522);
nor U27904 (N_27904,N_27230,N_27071);
or U27905 (N_27905,N_27551,N_27155);
or U27906 (N_27906,N_27069,N_27434);
nor U27907 (N_27907,N_27340,N_27496);
xor U27908 (N_27908,N_27352,N_27022);
or U27909 (N_27909,N_27294,N_27395);
and U27910 (N_27910,N_27109,N_27530);
or U27911 (N_27911,N_27570,N_27290);
nor U27912 (N_27912,N_27356,N_27476);
or U27913 (N_27913,N_27324,N_27118);
nand U27914 (N_27914,N_27160,N_27522);
and U27915 (N_27915,N_27451,N_27408);
nand U27916 (N_27916,N_27126,N_27518);
or U27917 (N_27917,N_27186,N_27434);
or U27918 (N_27918,N_27265,N_27291);
and U27919 (N_27919,N_27556,N_27084);
or U27920 (N_27920,N_27250,N_27473);
or U27921 (N_27921,N_27277,N_27218);
nand U27922 (N_27922,N_27386,N_27385);
xnor U27923 (N_27923,N_27216,N_27091);
nor U27924 (N_27924,N_27299,N_27009);
and U27925 (N_27925,N_27009,N_27104);
or U27926 (N_27926,N_27356,N_27538);
or U27927 (N_27927,N_27546,N_27501);
and U27928 (N_27928,N_27468,N_27448);
or U27929 (N_27929,N_27035,N_27306);
and U27930 (N_27930,N_27235,N_27180);
nor U27931 (N_27931,N_27070,N_27061);
and U27932 (N_27932,N_27283,N_27339);
xor U27933 (N_27933,N_27176,N_27588);
and U27934 (N_27934,N_27086,N_27423);
nor U27935 (N_27935,N_27059,N_27584);
nor U27936 (N_27936,N_27169,N_27446);
nand U27937 (N_27937,N_27495,N_27351);
nor U27938 (N_27938,N_27152,N_27521);
and U27939 (N_27939,N_27494,N_27395);
nor U27940 (N_27940,N_27250,N_27027);
and U27941 (N_27941,N_27028,N_27115);
or U27942 (N_27942,N_27183,N_27239);
and U27943 (N_27943,N_27568,N_27315);
and U27944 (N_27944,N_27465,N_27115);
nand U27945 (N_27945,N_27052,N_27000);
and U27946 (N_27946,N_27178,N_27446);
nor U27947 (N_27947,N_27148,N_27593);
or U27948 (N_27948,N_27098,N_27320);
nand U27949 (N_27949,N_27404,N_27579);
nor U27950 (N_27950,N_27096,N_27573);
and U27951 (N_27951,N_27263,N_27106);
or U27952 (N_27952,N_27219,N_27301);
and U27953 (N_27953,N_27362,N_27160);
nand U27954 (N_27954,N_27530,N_27262);
or U27955 (N_27955,N_27547,N_27322);
xnor U27956 (N_27956,N_27412,N_27192);
and U27957 (N_27957,N_27492,N_27338);
nand U27958 (N_27958,N_27521,N_27216);
and U27959 (N_27959,N_27238,N_27174);
and U27960 (N_27960,N_27308,N_27325);
nor U27961 (N_27961,N_27526,N_27298);
nor U27962 (N_27962,N_27378,N_27391);
and U27963 (N_27963,N_27546,N_27135);
nand U27964 (N_27964,N_27105,N_27006);
nor U27965 (N_27965,N_27307,N_27472);
nand U27966 (N_27966,N_27153,N_27066);
nor U27967 (N_27967,N_27594,N_27588);
or U27968 (N_27968,N_27320,N_27444);
nand U27969 (N_27969,N_27394,N_27323);
nor U27970 (N_27970,N_27090,N_27227);
and U27971 (N_27971,N_27468,N_27404);
nor U27972 (N_27972,N_27596,N_27142);
and U27973 (N_27973,N_27246,N_27194);
and U27974 (N_27974,N_27268,N_27510);
and U27975 (N_27975,N_27100,N_27175);
xnor U27976 (N_27976,N_27449,N_27257);
xor U27977 (N_27977,N_27394,N_27375);
xor U27978 (N_27978,N_27475,N_27018);
xnor U27979 (N_27979,N_27033,N_27176);
nand U27980 (N_27980,N_27593,N_27353);
or U27981 (N_27981,N_27350,N_27118);
and U27982 (N_27982,N_27217,N_27488);
xnor U27983 (N_27983,N_27056,N_27133);
and U27984 (N_27984,N_27164,N_27161);
or U27985 (N_27985,N_27280,N_27269);
and U27986 (N_27986,N_27069,N_27079);
and U27987 (N_27987,N_27267,N_27257);
and U27988 (N_27988,N_27549,N_27452);
and U27989 (N_27989,N_27364,N_27340);
nand U27990 (N_27990,N_27588,N_27290);
nor U27991 (N_27991,N_27012,N_27140);
nor U27992 (N_27992,N_27240,N_27100);
nor U27993 (N_27993,N_27231,N_27243);
nand U27994 (N_27994,N_27092,N_27007);
nand U27995 (N_27995,N_27226,N_27132);
nor U27996 (N_27996,N_27038,N_27042);
xor U27997 (N_27997,N_27063,N_27045);
nor U27998 (N_27998,N_27150,N_27132);
or U27999 (N_27999,N_27472,N_27537);
nand U28000 (N_28000,N_27216,N_27348);
xor U28001 (N_28001,N_27442,N_27540);
xnor U28002 (N_28002,N_27229,N_27147);
xnor U28003 (N_28003,N_27534,N_27253);
and U28004 (N_28004,N_27266,N_27094);
xor U28005 (N_28005,N_27597,N_27157);
or U28006 (N_28006,N_27019,N_27378);
nor U28007 (N_28007,N_27145,N_27532);
nand U28008 (N_28008,N_27502,N_27414);
or U28009 (N_28009,N_27051,N_27301);
xor U28010 (N_28010,N_27454,N_27146);
and U28011 (N_28011,N_27365,N_27368);
or U28012 (N_28012,N_27105,N_27190);
or U28013 (N_28013,N_27500,N_27337);
nor U28014 (N_28014,N_27475,N_27588);
nand U28015 (N_28015,N_27077,N_27300);
nand U28016 (N_28016,N_27434,N_27210);
nand U28017 (N_28017,N_27099,N_27563);
nand U28018 (N_28018,N_27057,N_27464);
and U28019 (N_28019,N_27062,N_27237);
or U28020 (N_28020,N_27394,N_27164);
xor U28021 (N_28021,N_27185,N_27397);
nor U28022 (N_28022,N_27566,N_27150);
or U28023 (N_28023,N_27446,N_27137);
nor U28024 (N_28024,N_27176,N_27410);
nand U28025 (N_28025,N_27435,N_27366);
or U28026 (N_28026,N_27085,N_27141);
and U28027 (N_28027,N_27069,N_27041);
nor U28028 (N_28028,N_27317,N_27164);
and U28029 (N_28029,N_27227,N_27086);
and U28030 (N_28030,N_27400,N_27081);
nand U28031 (N_28031,N_27062,N_27368);
nand U28032 (N_28032,N_27239,N_27353);
and U28033 (N_28033,N_27266,N_27032);
or U28034 (N_28034,N_27080,N_27472);
or U28035 (N_28035,N_27152,N_27328);
nor U28036 (N_28036,N_27155,N_27565);
nor U28037 (N_28037,N_27249,N_27499);
or U28038 (N_28038,N_27134,N_27068);
xnor U28039 (N_28039,N_27116,N_27504);
nor U28040 (N_28040,N_27138,N_27570);
nor U28041 (N_28041,N_27022,N_27589);
xor U28042 (N_28042,N_27243,N_27125);
nand U28043 (N_28043,N_27557,N_27055);
and U28044 (N_28044,N_27338,N_27269);
nor U28045 (N_28045,N_27517,N_27069);
xnor U28046 (N_28046,N_27462,N_27069);
and U28047 (N_28047,N_27475,N_27243);
nor U28048 (N_28048,N_27367,N_27136);
and U28049 (N_28049,N_27213,N_27590);
nor U28050 (N_28050,N_27448,N_27211);
nor U28051 (N_28051,N_27592,N_27273);
and U28052 (N_28052,N_27466,N_27081);
or U28053 (N_28053,N_27515,N_27368);
or U28054 (N_28054,N_27061,N_27302);
and U28055 (N_28055,N_27493,N_27437);
nand U28056 (N_28056,N_27058,N_27462);
and U28057 (N_28057,N_27183,N_27226);
xor U28058 (N_28058,N_27555,N_27311);
nand U28059 (N_28059,N_27457,N_27363);
or U28060 (N_28060,N_27106,N_27400);
xnor U28061 (N_28061,N_27550,N_27219);
or U28062 (N_28062,N_27296,N_27102);
nand U28063 (N_28063,N_27210,N_27564);
xor U28064 (N_28064,N_27561,N_27070);
nand U28065 (N_28065,N_27275,N_27593);
and U28066 (N_28066,N_27545,N_27063);
nor U28067 (N_28067,N_27466,N_27463);
nand U28068 (N_28068,N_27094,N_27162);
xor U28069 (N_28069,N_27189,N_27250);
or U28070 (N_28070,N_27105,N_27175);
xnor U28071 (N_28071,N_27389,N_27545);
nand U28072 (N_28072,N_27500,N_27063);
and U28073 (N_28073,N_27321,N_27268);
xnor U28074 (N_28074,N_27446,N_27510);
and U28075 (N_28075,N_27205,N_27193);
xor U28076 (N_28076,N_27421,N_27459);
or U28077 (N_28077,N_27099,N_27296);
xor U28078 (N_28078,N_27563,N_27452);
and U28079 (N_28079,N_27448,N_27514);
xnor U28080 (N_28080,N_27422,N_27528);
or U28081 (N_28081,N_27599,N_27409);
xnor U28082 (N_28082,N_27113,N_27014);
nand U28083 (N_28083,N_27488,N_27215);
or U28084 (N_28084,N_27417,N_27453);
and U28085 (N_28085,N_27229,N_27176);
nand U28086 (N_28086,N_27187,N_27106);
xor U28087 (N_28087,N_27247,N_27540);
nand U28088 (N_28088,N_27398,N_27031);
xnor U28089 (N_28089,N_27339,N_27539);
and U28090 (N_28090,N_27505,N_27482);
nand U28091 (N_28091,N_27428,N_27144);
or U28092 (N_28092,N_27490,N_27540);
nor U28093 (N_28093,N_27384,N_27314);
nor U28094 (N_28094,N_27572,N_27424);
nand U28095 (N_28095,N_27001,N_27545);
nand U28096 (N_28096,N_27139,N_27340);
xnor U28097 (N_28097,N_27059,N_27448);
xnor U28098 (N_28098,N_27153,N_27340);
and U28099 (N_28099,N_27068,N_27272);
xnor U28100 (N_28100,N_27423,N_27140);
or U28101 (N_28101,N_27118,N_27371);
and U28102 (N_28102,N_27249,N_27044);
nand U28103 (N_28103,N_27164,N_27110);
xnor U28104 (N_28104,N_27377,N_27521);
or U28105 (N_28105,N_27562,N_27289);
xor U28106 (N_28106,N_27106,N_27273);
nand U28107 (N_28107,N_27225,N_27525);
nand U28108 (N_28108,N_27199,N_27226);
nor U28109 (N_28109,N_27347,N_27413);
nand U28110 (N_28110,N_27031,N_27309);
nand U28111 (N_28111,N_27050,N_27288);
xor U28112 (N_28112,N_27179,N_27197);
nor U28113 (N_28113,N_27301,N_27472);
nand U28114 (N_28114,N_27198,N_27014);
nand U28115 (N_28115,N_27192,N_27014);
or U28116 (N_28116,N_27110,N_27373);
or U28117 (N_28117,N_27419,N_27308);
or U28118 (N_28118,N_27301,N_27415);
and U28119 (N_28119,N_27513,N_27594);
and U28120 (N_28120,N_27289,N_27523);
or U28121 (N_28121,N_27306,N_27130);
nand U28122 (N_28122,N_27151,N_27388);
xnor U28123 (N_28123,N_27267,N_27353);
nand U28124 (N_28124,N_27386,N_27561);
and U28125 (N_28125,N_27051,N_27422);
nand U28126 (N_28126,N_27443,N_27590);
or U28127 (N_28127,N_27202,N_27306);
nand U28128 (N_28128,N_27272,N_27165);
xor U28129 (N_28129,N_27177,N_27193);
or U28130 (N_28130,N_27367,N_27448);
nand U28131 (N_28131,N_27304,N_27185);
or U28132 (N_28132,N_27388,N_27439);
nor U28133 (N_28133,N_27472,N_27303);
xnor U28134 (N_28134,N_27194,N_27138);
or U28135 (N_28135,N_27088,N_27472);
and U28136 (N_28136,N_27546,N_27484);
or U28137 (N_28137,N_27150,N_27036);
nor U28138 (N_28138,N_27540,N_27549);
nand U28139 (N_28139,N_27173,N_27242);
nor U28140 (N_28140,N_27570,N_27425);
nor U28141 (N_28141,N_27054,N_27541);
and U28142 (N_28142,N_27497,N_27186);
and U28143 (N_28143,N_27340,N_27329);
or U28144 (N_28144,N_27254,N_27538);
and U28145 (N_28145,N_27164,N_27357);
nor U28146 (N_28146,N_27188,N_27368);
nor U28147 (N_28147,N_27238,N_27478);
xnor U28148 (N_28148,N_27255,N_27127);
nor U28149 (N_28149,N_27132,N_27138);
or U28150 (N_28150,N_27352,N_27097);
or U28151 (N_28151,N_27516,N_27511);
nor U28152 (N_28152,N_27408,N_27595);
xnor U28153 (N_28153,N_27327,N_27125);
nand U28154 (N_28154,N_27153,N_27370);
xnor U28155 (N_28155,N_27151,N_27200);
and U28156 (N_28156,N_27574,N_27594);
or U28157 (N_28157,N_27421,N_27561);
and U28158 (N_28158,N_27228,N_27358);
or U28159 (N_28159,N_27344,N_27426);
nor U28160 (N_28160,N_27280,N_27250);
or U28161 (N_28161,N_27298,N_27043);
or U28162 (N_28162,N_27041,N_27550);
xor U28163 (N_28163,N_27217,N_27001);
or U28164 (N_28164,N_27480,N_27359);
or U28165 (N_28165,N_27040,N_27330);
and U28166 (N_28166,N_27403,N_27041);
xor U28167 (N_28167,N_27526,N_27574);
or U28168 (N_28168,N_27165,N_27398);
nor U28169 (N_28169,N_27040,N_27392);
nand U28170 (N_28170,N_27269,N_27555);
or U28171 (N_28171,N_27137,N_27370);
and U28172 (N_28172,N_27004,N_27059);
xnor U28173 (N_28173,N_27166,N_27185);
or U28174 (N_28174,N_27133,N_27067);
and U28175 (N_28175,N_27489,N_27349);
nand U28176 (N_28176,N_27227,N_27536);
xor U28177 (N_28177,N_27487,N_27509);
and U28178 (N_28178,N_27527,N_27597);
or U28179 (N_28179,N_27330,N_27365);
and U28180 (N_28180,N_27421,N_27211);
or U28181 (N_28181,N_27347,N_27097);
or U28182 (N_28182,N_27559,N_27538);
xor U28183 (N_28183,N_27584,N_27099);
and U28184 (N_28184,N_27455,N_27403);
nor U28185 (N_28185,N_27442,N_27166);
or U28186 (N_28186,N_27241,N_27089);
nor U28187 (N_28187,N_27151,N_27445);
xor U28188 (N_28188,N_27163,N_27104);
or U28189 (N_28189,N_27153,N_27576);
xor U28190 (N_28190,N_27597,N_27594);
and U28191 (N_28191,N_27172,N_27002);
and U28192 (N_28192,N_27213,N_27294);
xnor U28193 (N_28193,N_27505,N_27363);
and U28194 (N_28194,N_27551,N_27511);
or U28195 (N_28195,N_27505,N_27435);
nor U28196 (N_28196,N_27119,N_27500);
and U28197 (N_28197,N_27379,N_27376);
xor U28198 (N_28198,N_27596,N_27566);
and U28199 (N_28199,N_27285,N_27235);
or U28200 (N_28200,N_27902,N_28046);
or U28201 (N_28201,N_28108,N_28080);
nor U28202 (N_28202,N_27978,N_28186);
nand U28203 (N_28203,N_28105,N_27922);
and U28204 (N_28204,N_28119,N_27688);
nand U28205 (N_28205,N_27920,N_27947);
xor U28206 (N_28206,N_27952,N_27830);
xnor U28207 (N_28207,N_28093,N_27740);
nand U28208 (N_28208,N_28136,N_28182);
xnor U28209 (N_28209,N_27829,N_28142);
nor U28210 (N_28210,N_27743,N_27854);
nor U28211 (N_28211,N_28154,N_28082);
nand U28212 (N_28212,N_27974,N_27933);
and U28213 (N_28213,N_27926,N_27600);
and U28214 (N_28214,N_27898,N_27791);
nor U28215 (N_28215,N_28191,N_27623);
nor U28216 (N_28216,N_28079,N_27754);
or U28217 (N_28217,N_27836,N_27847);
xnor U28218 (N_28218,N_27726,N_27723);
nand U28219 (N_28219,N_28148,N_27907);
and U28220 (N_28220,N_27993,N_27940);
and U28221 (N_28221,N_27962,N_28107);
or U28222 (N_28222,N_27963,N_28134);
xor U28223 (N_28223,N_28097,N_28054);
xor U28224 (N_28224,N_28006,N_27931);
or U28225 (N_28225,N_27739,N_27633);
and U28226 (N_28226,N_27887,N_27879);
xnor U28227 (N_28227,N_27606,N_27760);
and U28228 (N_28228,N_27775,N_27742);
xor U28229 (N_28229,N_27778,N_27801);
nor U28230 (N_28230,N_27826,N_28092);
or U28231 (N_28231,N_27849,N_27965);
nand U28232 (N_28232,N_27783,N_28139);
or U28233 (N_28233,N_27724,N_28020);
xor U28234 (N_28234,N_28030,N_28069);
and U28235 (N_28235,N_27883,N_28034);
nor U28236 (N_28236,N_27881,N_27753);
or U28237 (N_28237,N_27820,N_27911);
nand U28238 (N_28238,N_27927,N_28122);
nand U28239 (N_28239,N_27719,N_27840);
and U28240 (N_28240,N_28192,N_28089);
nand U28241 (N_28241,N_27700,N_28028);
nand U28242 (N_28242,N_28130,N_27690);
nand U28243 (N_28243,N_27950,N_28026);
nand U28244 (N_28244,N_28145,N_27875);
xnor U28245 (N_28245,N_28061,N_27752);
or U28246 (N_28246,N_28086,N_27825);
xor U28247 (N_28247,N_28125,N_27811);
nor U28248 (N_28248,N_27808,N_27725);
and U28249 (N_28249,N_27785,N_27661);
nor U28250 (N_28250,N_27814,N_28194);
xnor U28251 (N_28251,N_28042,N_27917);
xnor U28252 (N_28252,N_27607,N_27873);
and U28253 (N_28253,N_27809,N_27908);
nand U28254 (N_28254,N_27738,N_28041);
and U28255 (N_28255,N_27648,N_27624);
nor U28256 (N_28256,N_27781,N_28022);
or U28257 (N_28257,N_27968,N_27627);
and U28258 (N_28258,N_27604,N_27741);
nand U28259 (N_28259,N_27789,N_27953);
nor U28260 (N_28260,N_28038,N_28178);
nand U28261 (N_28261,N_28123,N_28101);
and U28262 (N_28262,N_27712,N_27960);
nand U28263 (N_28263,N_27749,N_27680);
and U28264 (N_28264,N_27780,N_28155);
and U28265 (N_28265,N_27964,N_27602);
or U28266 (N_28266,N_27924,N_27870);
and U28267 (N_28267,N_28100,N_27876);
nor U28268 (N_28268,N_28156,N_27971);
nor U28269 (N_28269,N_27689,N_27949);
xor U28270 (N_28270,N_27997,N_28132);
or U28271 (N_28271,N_27795,N_28121);
xnor U28272 (N_28272,N_27656,N_28173);
and U28273 (N_28273,N_28117,N_28065);
nand U28274 (N_28274,N_27831,N_27747);
and U28275 (N_28275,N_27804,N_28106);
xor U28276 (N_28276,N_27822,N_28181);
and U28277 (N_28277,N_28070,N_27930);
xor U28278 (N_28278,N_27695,N_28021);
xor U28279 (N_28279,N_27787,N_27672);
xnor U28280 (N_28280,N_27982,N_27685);
nor U28281 (N_28281,N_27649,N_27709);
and U28282 (N_28282,N_28138,N_27698);
xnor U28283 (N_28283,N_27620,N_28165);
nand U28284 (N_28284,N_27605,N_28064);
and U28285 (N_28285,N_27641,N_27764);
nor U28286 (N_28286,N_27652,N_27736);
or U28287 (N_28287,N_27970,N_27660);
xnor U28288 (N_28288,N_28032,N_27731);
xnor U28289 (N_28289,N_27866,N_27897);
nand U28290 (N_28290,N_27852,N_27972);
or U28291 (N_28291,N_28098,N_27617);
nor U28292 (N_28292,N_27891,N_27824);
xnor U28293 (N_28293,N_27722,N_27991);
nand U28294 (N_28294,N_28072,N_27976);
or U28295 (N_28295,N_27892,N_27793);
nand U28296 (N_28296,N_27986,N_27704);
nor U28297 (N_28297,N_28025,N_28179);
nor U28298 (N_28298,N_27610,N_28018);
nand U28299 (N_28299,N_27957,N_28014);
nor U28300 (N_28300,N_27810,N_27834);
xnor U28301 (N_28301,N_27630,N_27612);
and U28302 (N_28302,N_27608,N_27702);
nor U28303 (N_28303,N_27805,N_27796);
and U28304 (N_28304,N_27903,N_27694);
nor U28305 (N_28305,N_27999,N_27967);
nor U28306 (N_28306,N_27877,N_27915);
and U28307 (N_28307,N_28039,N_28043);
or U28308 (N_28308,N_27951,N_27954);
nand U28309 (N_28309,N_27794,N_27647);
xor U28310 (N_28310,N_28051,N_27663);
nor U28311 (N_28311,N_27973,N_27913);
xnor U28312 (N_28312,N_28033,N_27899);
xnor U28313 (N_28313,N_27727,N_27782);
nor U28314 (N_28314,N_27683,N_27961);
nand U28315 (N_28315,N_27842,N_27681);
nand U28316 (N_28316,N_28141,N_27861);
xor U28317 (N_28317,N_27730,N_28040);
or U28318 (N_28318,N_27646,N_27639);
and U28319 (N_28319,N_27856,N_27886);
xnor U28320 (N_28320,N_28005,N_27687);
nor U28321 (N_28321,N_27654,N_28147);
nand U28322 (N_28322,N_28077,N_27958);
nand U28323 (N_28323,N_27645,N_28174);
nor U28324 (N_28324,N_27827,N_27880);
nor U28325 (N_28325,N_27621,N_28187);
xnor U28326 (N_28326,N_28185,N_28045);
nor U28327 (N_28327,N_28002,N_28103);
xnor U28328 (N_28328,N_27844,N_28044);
nand U28329 (N_28329,N_28113,N_27716);
nor U28330 (N_28330,N_28094,N_28160);
nand U28331 (N_28331,N_28078,N_27677);
or U28332 (N_28332,N_27912,N_27692);
or U28333 (N_28333,N_28009,N_28198);
and U28334 (N_28334,N_27664,N_27955);
or U28335 (N_28335,N_27987,N_27691);
or U28336 (N_28336,N_27860,N_27786);
xor U28337 (N_28337,N_27928,N_27817);
and U28338 (N_28338,N_27850,N_27618);
and U28339 (N_28339,N_27944,N_27790);
and U28340 (N_28340,N_27855,N_28062);
or U28341 (N_28341,N_28166,N_27632);
nand U28342 (N_28342,N_27750,N_28090);
nor U28343 (N_28343,N_27721,N_28088);
nor U28344 (N_28344,N_27909,N_27864);
or U28345 (N_28345,N_28193,N_28152);
or U28346 (N_28346,N_27684,N_27802);
or U28347 (N_28347,N_28015,N_27846);
xnor U28348 (N_28348,N_28199,N_28067);
xor U28349 (N_28349,N_28167,N_27772);
and U28350 (N_28350,N_27653,N_28172);
and U28351 (N_28351,N_27673,N_27788);
xor U28352 (N_28352,N_27765,N_27626);
and U28353 (N_28353,N_27706,N_27751);
or U28354 (N_28354,N_27705,N_27872);
xor U28355 (N_28355,N_28140,N_27714);
nor U28356 (N_28356,N_27888,N_27773);
or U28357 (N_28357,N_27910,N_28190);
xnor U28358 (N_28358,N_27867,N_28029);
or U28359 (N_28359,N_27635,N_27779);
nand U28360 (N_28360,N_28161,N_28011);
and U28361 (N_28361,N_28164,N_27884);
or U28362 (N_28362,N_27882,N_27946);
or U28363 (N_28363,N_27900,N_27853);
nand U28364 (N_28364,N_28149,N_27732);
nor U28365 (N_28365,N_27757,N_27662);
and U28366 (N_28366,N_28104,N_28170);
and U28367 (N_28367,N_27718,N_27869);
xor U28368 (N_28368,N_27699,N_28177);
or U28369 (N_28369,N_28031,N_27771);
or U28370 (N_28370,N_28013,N_27665);
xor U28371 (N_28371,N_28184,N_27998);
and U28372 (N_28372,N_27735,N_27756);
or U28373 (N_28373,N_28169,N_28036);
or U28374 (N_28374,N_27988,N_27923);
xnor U28375 (N_28375,N_27679,N_27770);
and U28376 (N_28376,N_28099,N_27625);
and U28377 (N_28377,N_28055,N_28159);
nor U28378 (N_28378,N_28057,N_27675);
nand U28379 (N_28379,N_27818,N_27995);
xnor U28380 (N_28380,N_27938,N_27769);
or U28381 (N_28381,N_27701,N_28197);
xor U28382 (N_28382,N_27893,N_27966);
nor U28383 (N_28383,N_28171,N_28076);
nor U28384 (N_28384,N_27835,N_27729);
or U28385 (N_28385,N_28053,N_27674);
nand U28386 (N_28386,N_28095,N_27977);
nand U28387 (N_28387,N_28068,N_27631);
nor U28388 (N_28388,N_27774,N_27768);
or U28389 (N_28389,N_28114,N_27916);
xnor U28390 (N_28390,N_27807,N_27761);
nand U28391 (N_28391,N_28111,N_28047);
nor U28392 (N_28392,N_27936,N_27763);
or U28393 (N_28393,N_27619,N_28049);
or U28394 (N_28394,N_27696,N_27655);
or U28395 (N_28395,N_28073,N_28183);
nor U28396 (N_28396,N_27734,N_28091);
nor U28397 (N_28397,N_28083,N_28081);
xnor U28398 (N_28398,N_28109,N_28003);
xnor U28399 (N_28399,N_28195,N_28163);
nor U28400 (N_28400,N_28124,N_28075);
xor U28401 (N_28401,N_27843,N_27823);
or U28402 (N_28402,N_27762,N_27848);
and U28403 (N_28403,N_27906,N_27925);
and U28404 (N_28404,N_28096,N_27905);
nor U28405 (N_28405,N_27746,N_27989);
xor U28406 (N_28406,N_27603,N_27932);
nand U28407 (N_28407,N_27668,N_27862);
nor U28408 (N_28408,N_28137,N_27642);
or U28409 (N_28409,N_27707,N_27609);
xnor U28410 (N_28410,N_28087,N_27667);
nor U28411 (N_28411,N_27914,N_27670);
nand U28412 (N_28412,N_27929,N_27613);
or U28413 (N_28413,N_28024,N_28066);
and U28414 (N_28414,N_28052,N_27616);
nand U28415 (N_28415,N_28158,N_28157);
nor U28416 (N_28416,N_27838,N_27728);
nor U28417 (N_28417,N_28176,N_27666);
nand U28418 (N_28418,N_27939,N_28180);
nor U28419 (N_28419,N_28071,N_28128);
xnor U28420 (N_28420,N_27839,N_27601);
nand U28421 (N_28421,N_27792,N_27798);
or U28422 (N_28422,N_27934,N_27697);
xnor U28423 (N_28423,N_27833,N_27767);
xor U28424 (N_28424,N_27969,N_28084);
or U28425 (N_28425,N_27733,N_27737);
nor U28426 (N_28426,N_27943,N_27918);
or U28427 (N_28427,N_28016,N_28143);
nand U28428 (N_28428,N_28127,N_27806);
nand U28429 (N_28429,N_27682,N_27711);
xor U28430 (N_28430,N_27766,N_27703);
and U28431 (N_28431,N_27799,N_27650);
or U28432 (N_28432,N_28008,N_27636);
nand U28433 (N_28433,N_27874,N_27992);
or U28434 (N_28434,N_27921,N_27980);
nand U28435 (N_28435,N_28012,N_27979);
and U28436 (N_28436,N_27815,N_27686);
nand U28437 (N_28437,N_27956,N_28035);
nand U28438 (N_28438,N_27858,N_28037);
nor U28439 (N_28439,N_27671,N_27851);
and U28440 (N_28440,N_28102,N_27676);
and U28441 (N_28441,N_28023,N_27996);
nor U28442 (N_28442,N_27813,N_27659);
or U28443 (N_28443,N_28050,N_28000);
xor U28444 (N_28444,N_28188,N_27800);
nor U28445 (N_28445,N_28115,N_28135);
and U28446 (N_28446,N_27857,N_27945);
xnor U28447 (N_28447,N_27859,N_28196);
xnor U28448 (N_28448,N_27622,N_27935);
or U28449 (N_28449,N_27816,N_28131);
and U28450 (N_28450,N_27643,N_27828);
or U28451 (N_28451,N_28133,N_28116);
or U28452 (N_28452,N_27744,N_27896);
nor U28453 (N_28453,N_28063,N_27748);
nor U28454 (N_28454,N_28129,N_27871);
or U28455 (N_28455,N_27959,N_27715);
nor U28456 (N_28456,N_27878,N_27901);
and U28457 (N_28457,N_28019,N_28027);
xor U28458 (N_28458,N_27994,N_27637);
nor U28459 (N_28459,N_27638,N_28017);
and U28460 (N_28460,N_28060,N_27797);
nand U28461 (N_28461,N_27868,N_27904);
xnor U28462 (N_28462,N_27984,N_28110);
or U28463 (N_28463,N_27615,N_28126);
xnor U28464 (N_28464,N_27678,N_28153);
or U28465 (N_28465,N_28120,N_28007);
xor U28466 (N_28466,N_28085,N_27759);
nand U28467 (N_28467,N_27717,N_28146);
or U28468 (N_28468,N_27658,N_27819);
xnor U28469 (N_28469,N_27894,N_27669);
and U28470 (N_28470,N_28175,N_27634);
nand U28471 (N_28471,N_27821,N_27890);
nand U28472 (N_28472,N_27657,N_27941);
and U28473 (N_28473,N_28004,N_27713);
nand U28474 (N_28474,N_27611,N_28118);
and U28475 (N_28475,N_27895,N_27776);
nand U28476 (N_28476,N_27837,N_27863);
or U28477 (N_28477,N_27812,N_27937);
xor U28478 (N_28478,N_27985,N_27777);
and U28479 (N_28479,N_28001,N_27832);
and U28480 (N_28480,N_27758,N_28144);
nand U28481 (N_28481,N_27803,N_27720);
nor U28482 (N_28482,N_27983,N_27865);
nor U28483 (N_28483,N_28162,N_27889);
nand U28484 (N_28484,N_28150,N_27640);
xor U28485 (N_28485,N_28059,N_27942);
or U28486 (N_28486,N_27845,N_27629);
xnor U28487 (N_28487,N_27784,N_27990);
nor U28488 (N_28488,N_28074,N_27948);
xnor U28489 (N_28489,N_27919,N_27981);
nor U28490 (N_28490,N_27628,N_28058);
and U28491 (N_28491,N_27651,N_28151);
or U28492 (N_28492,N_27708,N_27614);
nor U28493 (N_28493,N_27841,N_28010);
nand U28494 (N_28494,N_27693,N_28048);
nor U28495 (N_28495,N_27755,N_28189);
or U28496 (N_28496,N_28112,N_27644);
and U28497 (N_28497,N_27975,N_28168);
xor U28498 (N_28498,N_28056,N_27710);
or U28499 (N_28499,N_27745,N_27885);
and U28500 (N_28500,N_27923,N_27789);
nor U28501 (N_28501,N_27991,N_28047);
xor U28502 (N_28502,N_27665,N_28020);
or U28503 (N_28503,N_27851,N_27690);
and U28504 (N_28504,N_27691,N_27724);
nand U28505 (N_28505,N_28073,N_28001);
nor U28506 (N_28506,N_28171,N_27989);
nor U28507 (N_28507,N_27873,N_27942);
and U28508 (N_28508,N_28034,N_27803);
xor U28509 (N_28509,N_28057,N_27922);
xnor U28510 (N_28510,N_28001,N_27785);
nor U28511 (N_28511,N_27986,N_28122);
and U28512 (N_28512,N_27905,N_28098);
nand U28513 (N_28513,N_27940,N_27825);
xor U28514 (N_28514,N_27909,N_27891);
nand U28515 (N_28515,N_28129,N_28126);
or U28516 (N_28516,N_28048,N_27801);
nor U28517 (N_28517,N_27881,N_27855);
nor U28518 (N_28518,N_28017,N_27741);
nand U28519 (N_28519,N_27839,N_27906);
or U28520 (N_28520,N_27971,N_27699);
nor U28521 (N_28521,N_27735,N_27847);
or U28522 (N_28522,N_27620,N_27911);
and U28523 (N_28523,N_28112,N_27831);
or U28524 (N_28524,N_28075,N_27736);
nand U28525 (N_28525,N_27921,N_27863);
and U28526 (N_28526,N_27773,N_27899);
nand U28527 (N_28527,N_28077,N_27908);
nand U28528 (N_28528,N_27601,N_27613);
or U28529 (N_28529,N_27653,N_27704);
xnor U28530 (N_28530,N_28060,N_28026);
xnor U28531 (N_28531,N_27773,N_28038);
or U28532 (N_28532,N_28159,N_27975);
nor U28533 (N_28533,N_27683,N_28065);
nor U28534 (N_28534,N_27793,N_28033);
nand U28535 (N_28535,N_27984,N_27996);
xor U28536 (N_28536,N_27927,N_27676);
xor U28537 (N_28537,N_27771,N_28025);
nor U28538 (N_28538,N_27771,N_27823);
and U28539 (N_28539,N_27766,N_27900);
nand U28540 (N_28540,N_27604,N_27952);
or U28541 (N_28541,N_27769,N_27944);
and U28542 (N_28542,N_28027,N_27894);
nand U28543 (N_28543,N_27915,N_28082);
nand U28544 (N_28544,N_27643,N_27625);
and U28545 (N_28545,N_27843,N_28071);
or U28546 (N_28546,N_27942,N_27795);
nand U28547 (N_28547,N_27756,N_27962);
or U28548 (N_28548,N_28119,N_27990);
nand U28549 (N_28549,N_28080,N_27617);
and U28550 (N_28550,N_27976,N_27777);
nor U28551 (N_28551,N_27883,N_28153);
or U28552 (N_28552,N_28018,N_28045);
xor U28553 (N_28553,N_27928,N_27867);
nor U28554 (N_28554,N_27949,N_27969);
nor U28555 (N_28555,N_27973,N_27925);
nor U28556 (N_28556,N_27740,N_27979);
or U28557 (N_28557,N_28185,N_27606);
or U28558 (N_28558,N_28143,N_28057);
and U28559 (N_28559,N_27953,N_27989);
and U28560 (N_28560,N_28002,N_27812);
nor U28561 (N_28561,N_27713,N_28150);
or U28562 (N_28562,N_27887,N_27712);
and U28563 (N_28563,N_27960,N_28043);
nand U28564 (N_28564,N_27889,N_27801);
nand U28565 (N_28565,N_27773,N_27911);
nand U28566 (N_28566,N_27719,N_28135);
xor U28567 (N_28567,N_27919,N_27785);
nand U28568 (N_28568,N_28128,N_27905);
or U28569 (N_28569,N_28120,N_27786);
xor U28570 (N_28570,N_28065,N_28054);
nor U28571 (N_28571,N_27653,N_28003);
and U28572 (N_28572,N_28181,N_27806);
nand U28573 (N_28573,N_27842,N_28186);
nand U28574 (N_28574,N_28032,N_28138);
or U28575 (N_28575,N_28181,N_27705);
or U28576 (N_28576,N_28022,N_27621);
or U28577 (N_28577,N_27637,N_27671);
xnor U28578 (N_28578,N_28095,N_28055);
xor U28579 (N_28579,N_27883,N_27916);
nor U28580 (N_28580,N_27886,N_28172);
nor U28581 (N_28581,N_27786,N_27673);
nand U28582 (N_28582,N_27667,N_27995);
nand U28583 (N_28583,N_27807,N_28026);
nor U28584 (N_28584,N_27821,N_27960);
xor U28585 (N_28585,N_27902,N_28066);
xor U28586 (N_28586,N_27937,N_28163);
and U28587 (N_28587,N_27859,N_28071);
nor U28588 (N_28588,N_27963,N_27786);
and U28589 (N_28589,N_28110,N_27827);
and U28590 (N_28590,N_27974,N_28151);
and U28591 (N_28591,N_27921,N_28040);
and U28592 (N_28592,N_28074,N_27832);
and U28593 (N_28593,N_28186,N_28184);
xor U28594 (N_28594,N_27809,N_28145);
nor U28595 (N_28595,N_27684,N_27707);
or U28596 (N_28596,N_27971,N_28049);
nor U28597 (N_28597,N_27910,N_27831);
nor U28598 (N_28598,N_27798,N_27649);
and U28599 (N_28599,N_28080,N_27661);
or U28600 (N_28600,N_28085,N_28029);
xnor U28601 (N_28601,N_28028,N_27896);
and U28602 (N_28602,N_27716,N_28146);
or U28603 (N_28603,N_27984,N_27775);
xnor U28604 (N_28604,N_27847,N_28196);
nor U28605 (N_28605,N_27739,N_27909);
nand U28606 (N_28606,N_27817,N_27657);
and U28607 (N_28607,N_28026,N_28000);
nor U28608 (N_28608,N_28111,N_27983);
nor U28609 (N_28609,N_28049,N_27843);
and U28610 (N_28610,N_28018,N_28156);
or U28611 (N_28611,N_27898,N_27754);
xor U28612 (N_28612,N_27679,N_27833);
xor U28613 (N_28613,N_27768,N_28034);
or U28614 (N_28614,N_27840,N_28177);
nor U28615 (N_28615,N_27647,N_27691);
nor U28616 (N_28616,N_28186,N_27846);
nor U28617 (N_28617,N_27799,N_27862);
or U28618 (N_28618,N_27680,N_28016);
nand U28619 (N_28619,N_27802,N_27668);
xnor U28620 (N_28620,N_28179,N_27713);
nand U28621 (N_28621,N_27720,N_27892);
or U28622 (N_28622,N_27822,N_27730);
xor U28623 (N_28623,N_27930,N_27758);
nand U28624 (N_28624,N_28151,N_27980);
nor U28625 (N_28625,N_28063,N_27698);
and U28626 (N_28626,N_28098,N_28078);
nor U28627 (N_28627,N_27694,N_27855);
xnor U28628 (N_28628,N_28051,N_27776);
nor U28629 (N_28629,N_27720,N_27781);
or U28630 (N_28630,N_27989,N_28196);
nand U28631 (N_28631,N_27930,N_27899);
nor U28632 (N_28632,N_27924,N_28172);
or U28633 (N_28633,N_27987,N_28191);
nand U28634 (N_28634,N_27832,N_27785);
nand U28635 (N_28635,N_28153,N_27867);
or U28636 (N_28636,N_28110,N_28105);
xnor U28637 (N_28637,N_27656,N_28172);
nand U28638 (N_28638,N_27862,N_28150);
and U28639 (N_28639,N_27657,N_28028);
xor U28640 (N_28640,N_28088,N_27606);
xnor U28641 (N_28641,N_27615,N_27956);
nor U28642 (N_28642,N_28126,N_27973);
xor U28643 (N_28643,N_27814,N_28175);
nor U28644 (N_28644,N_27674,N_28131);
or U28645 (N_28645,N_27661,N_27744);
nor U28646 (N_28646,N_28175,N_27675);
or U28647 (N_28647,N_27794,N_28072);
or U28648 (N_28648,N_27657,N_28119);
and U28649 (N_28649,N_27877,N_27826);
xor U28650 (N_28650,N_27790,N_27967);
and U28651 (N_28651,N_27762,N_28109);
nand U28652 (N_28652,N_27974,N_27899);
or U28653 (N_28653,N_28010,N_27695);
or U28654 (N_28654,N_27748,N_28064);
xnor U28655 (N_28655,N_28018,N_27862);
xnor U28656 (N_28656,N_28103,N_27637);
xor U28657 (N_28657,N_28046,N_28132);
and U28658 (N_28658,N_27891,N_27877);
or U28659 (N_28659,N_27730,N_27753);
or U28660 (N_28660,N_28156,N_28089);
nand U28661 (N_28661,N_27610,N_27747);
nand U28662 (N_28662,N_27843,N_27721);
and U28663 (N_28663,N_27844,N_28153);
nand U28664 (N_28664,N_28060,N_28165);
xor U28665 (N_28665,N_28001,N_28163);
nand U28666 (N_28666,N_27712,N_28045);
xor U28667 (N_28667,N_27730,N_27909);
nor U28668 (N_28668,N_27957,N_27876);
and U28669 (N_28669,N_27823,N_27976);
and U28670 (N_28670,N_27802,N_27940);
nor U28671 (N_28671,N_27650,N_27928);
or U28672 (N_28672,N_27760,N_27824);
nor U28673 (N_28673,N_27888,N_27882);
and U28674 (N_28674,N_28133,N_27968);
nor U28675 (N_28675,N_27683,N_28123);
or U28676 (N_28676,N_28135,N_27641);
or U28677 (N_28677,N_27957,N_27709);
nor U28678 (N_28678,N_27864,N_27915);
nor U28679 (N_28679,N_27986,N_27602);
xnor U28680 (N_28680,N_27850,N_27877);
nor U28681 (N_28681,N_28172,N_28140);
and U28682 (N_28682,N_27954,N_27779);
nor U28683 (N_28683,N_27827,N_28056);
xnor U28684 (N_28684,N_27899,N_27878);
nand U28685 (N_28685,N_27904,N_27669);
and U28686 (N_28686,N_28110,N_27988);
or U28687 (N_28687,N_27638,N_27862);
and U28688 (N_28688,N_27700,N_27952);
and U28689 (N_28689,N_27975,N_27909);
and U28690 (N_28690,N_27935,N_27930);
or U28691 (N_28691,N_28166,N_28082);
nor U28692 (N_28692,N_27788,N_28073);
and U28693 (N_28693,N_28095,N_28075);
and U28694 (N_28694,N_28032,N_27620);
or U28695 (N_28695,N_27678,N_27807);
nand U28696 (N_28696,N_27993,N_28017);
nor U28697 (N_28697,N_27641,N_28116);
and U28698 (N_28698,N_27904,N_28027);
nand U28699 (N_28699,N_28159,N_27672);
xor U28700 (N_28700,N_28095,N_27993);
xnor U28701 (N_28701,N_27886,N_27607);
xor U28702 (N_28702,N_28096,N_28005);
or U28703 (N_28703,N_28107,N_28067);
and U28704 (N_28704,N_28037,N_27671);
xnor U28705 (N_28705,N_27834,N_27673);
nor U28706 (N_28706,N_27751,N_27715);
xor U28707 (N_28707,N_27971,N_27685);
and U28708 (N_28708,N_28145,N_27972);
nand U28709 (N_28709,N_28179,N_27670);
nor U28710 (N_28710,N_28105,N_28170);
nand U28711 (N_28711,N_27842,N_27686);
nor U28712 (N_28712,N_27681,N_27804);
nor U28713 (N_28713,N_27815,N_28121);
xor U28714 (N_28714,N_28166,N_27633);
xor U28715 (N_28715,N_27813,N_27916);
xnor U28716 (N_28716,N_27930,N_27620);
nor U28717 (N_28717,N_27939,N_27813);
nor U28718 (N_28718,N_28131,N_27773);
xnor U28719 (N_28719,N_27870,N_28024);
nor U28720 (N_28720,N_27779,N_27892);
nor U28721 (N_28721,N_27828,N_27781);
or U28722 (N_28722,N_28167,N_27733);
and U28723 (N_28723,N_27756,N_27722);
or U28724 (N_28724,N_27746,N_27695);
nand U28725 (N_28725,N_28011,N_28103);
xnor U28726 (N_28726,N_27788,N_27954);
xor U28727 (N_28727,N_28185,N_28067);
xnor U28728 (N_28728,N_27759,N_28074);
and U28729 (N_28729,N_27798,N_27732);
and U28730 (N_28730,N_27753,N_27740);
nand U28731 (N_28731,N_27776,N_27751);
nand U28732 (N_28732,N_27673,N_27881);
nor U28733 (N_28733,N_28052,N_27750);
nand U28734 (N_28734,N_27985,N_28118);
nor U28735 (N_28735,N_27691,N_28039);
xnor U28736 (N_28736,N_28051,N_27680);
or U28737 (N_28737,N_27623,N_28104);
xnor U28738 (N_28738,N_27669,N_27761);
or U28739 (N_28739,N_27892,N_28013);
nand U28740 (N_28740,N_27793,N_28030);
and U28741 (N_28741,N_27682,N_27842);
and U28742 (N_28742,N_27765,N_27900);
and U28743 (N_28743,N_28100,N_27824);
or U28744 (N_28744,N_27688,N_27981);
or U28745 (N_28745,N_28166,N_28006);
xnor U28746 (N_28746,N_27980,N_28024);
or U28747 (N_28747,N_27746,N_27725);
and U28748 (N_28748,N_27705,N_27866);
nor U28749 (N_28749,N_27782,N_27930);
xnor U28750 (N_28750,N_27612,N_27931);
and U28751 (N_28751,N_27607,N_27876);
and U28752 (N_28752,N_28049,N_27941);
nand U28753 (N_28753,N_27886,N_27947);
nand U28754 (N_28754,N_27957,N_27609);
xnor U28755 (N_28755,N_28077,N_28128);
nand U28756 (N_28756,N_28059,N_27865);
nor U28757 (N_28757,N_28019,N_27776);
xnor U28758 (N_28758,N_27837,N_27942);
xor U28759 (N_28759,N_27929,N_27868);
xnor U28760 (N_28760,N_28159,N_28169);
xor U28761 (N_28761,N_28085,N_28192);
nand U28762 (N_28762,N_28131,N_27691);
nor U28763 (N_28763,N_28122,N_27775);
xnor U28764 (N_28764,N_27807,N_28100);
nand U28765 (N_28765,N_27792,N_27806);
nor U28766 (N_28766,N_27775,N_27735);
nand U28767 (N_28767,N_27716,N_28097);
or U28768 (N_28768,N_27809,N_27778);
nand U28769 (N_28769,N_27617,N_28180);
or U28770 (N_28770,N_28119,N_27982);
nor U28771 (N_28771,N_28067,N_28092);
or U28772 (N_28772,N_28024,N_27873);
or U28773 (N_28773,N_27620,N_27953);
xnor U28774 (N_28774,N_28078,N_27960);
and U28775 (N_28775,N_27825,N_28194);
nor U28776 (N_28776,N_27689,N_27960);
xor U28777 (N_28777,N_28109,N_28062);
nor U28778 (N_28778,N_27971,N_27941);
nand U28779 (N_28779,N_27604,N_27688);
nor U28780 (N_28780,N_27658,N_27975);
and U28781 (N_28781,N_28099,N_27875);
and U28782 (N_28782,N_27649,N_27866);
nand U28783 (N_28783,N_28057,N_27733);
or U28784 (N_28784,N_28020,N_28153);
or U28785 (N_28785,N_27725,N_27650);
xnor U28786 (N_28786,N_27604,N_28194);
and U28787 (N_28787,N_27711,N_27814);
nor U28788 (N_28788,N_28054,N_27742);
and U28789 (N_28789,N_27801,N_27639);
nand U28790 (N_28790,N_28187,N_28069);
and U28791 (N_28791,N_28168,N_28148);
nand U28792 (N_28792,N_27795,N_27898);
nand U28793 (N_28793,N_27785,N_27609);
nand U28794 (N_28794,N_27742,N_28056);
nand U28795 (N_28795,N_28165,N_27936);
or U28796 (N_28796,N_28028,N_27832);
nand U28797 (N_28797,N_27935,N_28196);
or U28798 (N_28798,N_27925,N_28079);
nor U28799 (N_28799,N_27834,N_27748);
nor U28800 (N_28800,N_28708,N_28574);
nand U28801 (N_28801,N_28352,N_28288);
nand U28802 (N_28802,N_28509,N_28525);
nor U28803 (N_28803,N_28203,N_28629);
nand U28804 (N_28804,N_28799,N_28404);
xnor U28805 (N_28805,N_28244,N_28587);
nor U28806 (N_28806,N_28546,N_28528);
or U28807 (N_28807,N_28502,N_28726);
nand U28808 (N_28808,N_28275,N_28327);
xnor U28809 (N_28809,N_28453,N_28610);
nand U28810 (N_28810,N_28754,N_28594);
nand U28811 (N_28811,N_28556,N_28326);
and U28812 (N_28812,N_28294,N_28265);
nand U28813 (N_28813,N_28691,N_28224);
nor U28814 (N_28814,N_28335,N_28599);
or U28815 (N_28815,N_28664,N_28670);
xor U28816 (N_28816,N_28282,N_28758);
nand U28817 (N_28817,N_28416,N_28504);
nand U28818 (N_28818,N_28591,N_28257);
xnor U28819 (N_28819,N_28560,N_28766);
or U28820 (N_28820,N_28314,N_28709);
xor U28821 (N_28821,N_28261,N_28748);
or U28822 (N_28822,N_28618,N_28447);
xor U28823 (N_28823,N_28503,N_28713);
and U28824 (N_28824,N_28479,N_28354);
nand U28825 (N_28825,N_28566,N_28559);
or U28826 (N_28826,N_28222,N_28297);
nand U28827 (N_28827,N_28508,N_28434);
xnor U28828 (N_28828,N_28572,N_28392);
nor U28829 (N_28829,N_28728,N_28607);
and U28830 (N_28830,N_28789,N_28755);
nand U28831 (N_28831,N_28237,N_28285);
and U28832 (N_28832,N_28299,N_28692);
and U28833 (N_28833,N_28321,N_28476);
xor U28834 (N_28834,N_28620,N_28338);
nor U28835 (N_28835,N_28281,N_28756);
nand U28836 (N_28836,N_28346,N_28760);
and U28837 (N_28837,N_28358,N_28557);
xor U28838 (N_28838,N_28783,N_28584);
and U28839 (N_28839,N_28201,N_28682);
or U28840 (N_28840,N_28400,N_28384);
xor U28841 (N_28841,N_28795,N_28483);
nor U28842 (N_28842,N_28268,N_28649);
nor U28843 (N_28843,N_28459,N_28598);
or U28844 (N_28844,N_28383,N_28370);
and U28845 (N_28845,N_28633,N_28570);
nor U28846 (N_28846,N_28717,N_28262);
and U28847 (N_28847,N_28341,N_28291);
nor U28848 (N_28848,N_28636,N_28589);
nor U28849 (N_28849,N_28251,N_28298);
and U28850 (N_28850,N_28538,N_28233);
nand U28851 (N_28851,N_28277,N_28641);
nor U28852 (N_28852,N_28628,N_28736);
nand U28853 (N_28853,N_28438,N_28531);
xor U28854 (N_28854,N_28676,N_28622);
nand U28855 (N_28855,N_28389,N_28548);
xor U28856 (N_28856,N_28724,N_28240);
nor U28857 (N_28857,N_28227,N_28207);
nor U28858 (N_28858,N_28465,N_28242);
or U28859 (N_28859,N_28444,N_28302);
and U28860 (N_28860,N_28308,N_28774);
nor U28861 (N_28861,N_28600,N_28428);
and U28862 (N_28862,N_28450,N_28613);
xor U28863 (N_28863,N_28549,N_28284);
or U28864 (N_28864,N_28510,N_28456);
or U28865 (N_28865,N_28655,N_28597);
or U28866 (N_28866,N_28707,N_28675);
or U28867 (N_28867,N_28543,N_28443);
nor U28868 (N_28868,N_28605,N_28455);
nor U28869 (N_28869,N_28727,N_28394);
nor U28870 (N_28870,N_28669,N_28309);
and U28871 (N_28871,N_28506,N_28787);
or U28872 (N_28872,N_28374,N_28289);
or U28873 (N_28873,N_28753,N_28554);
nand U28874 (N_28874,N_28577,N_28419);
and U28875 (N_28875,N_28396,N_28377);
nand U28876 (N_28876,N_28463,N_28778);
nand U28877 (N_28877,N_28360,N_28494);
xor U28878 (N_28878,N_28482,N_28292);
nand U28879 (N_28879,N_28445,N_28208);
nand U28880 (N_28880,N_28501,N_28779);
or U28881 (N_28881,N_28684,N_28290);
and U28882 (N_28882,N_28446,N_28334);
nor U28883 (N_28883,N_28611,N_28763);
or U28884 (N_28884,N_28712,N_28263);
and U28885 (N_28885,N_28656,N_28359);
nor U28886 (N_28886,N_28612,N_28530);
and U28887 (N_28887,N_28274,N_28380);
xnor U28888 (N_28888,N_28686,N_28313);
and U28889 (N_28889,N_28330,N_28775);
nor U28890 (N_28890,N_28466,N_28704);
nor U28891 (N_28891,N_28700,N_28634);
nand U28892 (N_28892,N_28345,N_28423);
or U28893 (N_28893,N_28410,N_28220);
or U28894 (N_28894,N_28513,N_28792);
or U28895 (N_28895,N_28322,N_28544);
and U28896 (N_28896,N_28542,N_28286);
or U28897 (N_28897,N_28451,N_28588);
nor U28898 (N_28898,N_28209,N_28514);
nor U28899 (N_28899,N_28376,N_28395);
nand U28900 (N_28900,N_28499,N_28433);
and U28901 (N_28901,N_28351,N_28498);
or U28902 (N_28902,N_28462,N_28470);
nand U28903 (N_28903,N_28536,N_28517);
nand U28904 (N_28904,N_28661,N_28399);
xor U28905 (N_28905,N_28752,N_28361);
xnor U28906 (N_28906,N_28743,N_28604);
nor U28907 (N_28907,N_28586,N_28683);
or U28908 (N_28908,N_28718,N_28417);
nand U28909 (N_28909,N_28414,N_28468);
nand U28910 (N_28910,N_28312,N_28333);
and U28911 (N_28911,N_28595,N_28614);
nor U28912 (N_28912,N_28214,N_28762);
and U28913 (N_28913,N_28307,N_28635);
xnor U28914 (N_28914,N_28735,N_28402);
or U28915 (N_28915,N_28545,N_28720);
nor U28916 (N_28916,N_28658,N_28674);
xor U28917 (N_28917,N_28678,N_28798);
or U28918 (N_28918,N_28253,N_28537);
nand U28919 (N_28919,N_28436,N_28272);
nand U28920 (N_28920,N_28715,N_28256);
nor U28921 (N_28921,N_28271,N_28353);
nor U28922 (N_28922,N_28780,N_28315);
nand U28923 (N_28923,N_28391,N_28551);
or U28924 (N_28924,N_28300,N_28212);
nand U28925 (N_28925,N_28637,N_28473);
or U28926 (N_28926,N_28681,N_28491);
and U28927 (N_28927,N_28356,N_28532);
and U28928 (N_28928,N_28238,N_28344);
nor U28929 (N_28929,N_28642,N_28461);
xnor U28930 (N_28930,N_28460,N_28487);
and U28931 (N_28931,N_28425,N_28699);
nor U28932 (N_28932,N_28511,N_28663);
nor U28933 (N_28933,N_28247,N_28608);
xor U28934 (N_28934,N_28547,N_28449);
and U28935 (N_28935,N_28342,N_28492);
xor U28936 (N_28936,N_28403,N_28388);
or U28937 (N_28937,N_28606,N_28363);
nand U28938 (N_28938,N_28200,N_28258);
nor U28939 (N_28939,N_28386,N_28585);
xnor U28940 (N_28940,N_28793,N_28236);
or U28941 (N_28941,N_28582,N_28615);
xor U28942 (N_28942,N_28710,N_28381);
nor U28943 (N_28943,N_28702,N_28471);
and U28944 (N_28944,N_28405,N_28540);
nor U28945 (N_28945,N_28287,N_28228);
or U28946 (N_28946,N_28719,N_28219);
or U28947 (N_28947,N_28519,N_28293);
nor U28948 (N_28948,N_28750,N_28500);
xor U28949 (N_28949,N_28393,N_28329);
xor U28950 (N_28950,N_28533,N_28490);
nor U28951 (N_28951,N_28467,N_28527);
nor U28952 (N_28952,N_28362,N_28680);
nand U28953 (N_28953,N_28378,N_28472);
xor U28954 (N_28954,N_28442,N_28507);
or U28955 (N_28955,N_28521,N_28331);
nand U28956 (N_28956,N_28458,N_28348);
or U28957 (N_28957,N_28685,N_28552);
or U28958 (N_28958,N_28617,N_28497);
or U28959 (N_28959,N_28254,N_28406);
xnor U28960 (N_28960,N_28318,N_28368);
or U28961 (N_28961,N_28316,N_28535);
xnor U28962 (N_28962,N_28235,N_28662);
and U28963 (N_28963,N_28706,N_28243);
nand U28964 (N_28964,N_28731,N_28665);
nand U28965 (N_28965,N_28379,N_28448);
or U28966 (N_28966,N_28304,N_28323);
and U28967 (N_28967,N_28569,N_28474);
nand U28968 (N_28968,N_28301,N_28751);
xnor U28969 (N_28969,N_28246,N_28215);
xnor U28970 (N_28970,N_28695,N_28529);
nand U28971 (N_28971,N_28580,N_28796);
xor U28972 (N_28972,N_28276,N_28267);
nand U28973 (N_28973,N_28689,N_28457);
nor U28974 (N_28974,N_28581,N_28625);
nor U28975 (N_28975,N_28364,N_28260);
or U28976 (N_28976,N_28431,N_28679);
and U28977 (N_28977,N_28365,N_28630);
or U28978 (N_28978,N_28744,N_28657);
nand U28979 (N_28979,N_28213,N_28310);
xnor U28980 (N_28980,N_28204,N_28740);
nand U28981 (N_28981,N_28624,N_28369);
nand U28982 (N_28982,N_28454,N_28452);
or U28983 (N_28983,N_28772,N_28279);
and U28984 (N_28984,N_28324,N_28218);
nand U28985 (N_28985,N_28325,N_28248);
xor U28986 (N_28986,N_28469,N_28421);
nor U28987 (N_28987,N_28375,N_28645);
and U28988 (N_28988,N_28512,N_28269);
or U28989 (N_28989,N_28648,N_28283);
nand U28990 (N_28990,N_28477,N_28734);
nor U28991 (N_28991,N_28765,N_28266);
nor U28992 (N_28992,N_28385,N_28343);
or U28993 (N_28993,N_28553,N_28576);
nand U28994 (N_28994,N_28439,N_28534);
and U28995 (N_28995,N_28273,N_28688);
nor U28996 (N_28996,N_28722,N_28305);
nand U28997 (N_28997,N_28252,N_28231);
nor U28998 (N_28998,N_28741,N_28716);
and U28999 (N_28999,N_28210,N_28573);
and U29000 (N_29000,N_28328,N_28568);
and U29001 (N_29001,N_28484,N_28366);
xor U29002 (N_29002,N_28794,N_28601);
or U29003 (N_29003,N_28563,N_28621);
nor U29004 (N_29004,N_28673,N_28690);
nor U29005 (N_29005,N_28562,N_28697);
and U29006 (N_29006,N_28522,N_28784);
or U29007 (N_29007,N_28632,N_28475);
xnor U29008 (N_29008,N_28739,N_28422);
or U29009 (N_29009,N_28644,N_28721);
nand U29010 (N_29010,N_28303,N_28347);
nand U29011 (N_29011,N_28781,N_28420);
xor U29012 (N_29012,N_28249,N_28647);
nor U29013 (N_29013,N_28541,N_28478);
nor U29014 (N_29014,N_28603,N_28349);
and U29015 (N_29015,N_28782,N_28495);
xor U29016 (N_29016,N_28785,N_28245);
nor U29017 (N_29017,N_28761,N_28232);
nand U29018 (N_29018,N_28486,N_28437);
nor U29019 (N_29019,N_28745,N_28653);
or U29020 (N_29020,N_28205,N_28759);
nor U29021 (N_29021,N_28424,N_28367);
nand U29022 (N_29022,N_28723,N_28229);
nand U29023 (N_29023,N_28650,N_28769);
nor U29024 (N_29024,N_28429,N_28311);
xnor U29025 (N_29025,N_28730,N_28590);
or U29026 (N_29026,N_28555,N_28703);
xnor U29027 (N_29027,N_28320,N_28742);
nand U29028 (N_29028,N_28771,N_28578);
nor U29029 (N_29029,N_28667,N_28426);
and U29030 (N_29030,N_28440,N_28481);
and U29031 (N_29031,N_28790,N_28415);
and U29032 (N_29032,N_28666,N_28216);
nor U29033 (N_29033,N_28797,N_28732);
nor U29034 (N_29034,N_28640,N_28738);
xor U29035 (N_29035,N_28239,N_28340);
or U29036 (N_29036,N_28561,N_28764);
and U29037 (N_29037,N_28631,N_28217);
or U29038 (N_29038,N_28652,N_28671);
or U29039 (N_29039,N_28623,N_28639);
and U29040 (N_29040,N_28770,N_28776);
nor U29041 (N_29041,N_28295,N_28278);
and U29042 (N_29042,N_28523,N_28518);
or U29043 (N_29043,N_28432,N_28317);
nand U29044 (N_29044,N_28435,N_28259);
or U29045 (N_29045,N_28592,N_28332);
xnor U29046 (N_29046,N_28693,N_28651);
nand U29047 (N_29047,N_28694,N_28526);
nand U29048 (N_29048,N_28306,N_28791);
and U29049 (N_29049,N_28409,N_28619);
or U29050 (N_29050,N_28387,N_28638);
and U29051 (N_29051,N_28737,N_28505);
xnor U29052 (N_29052,N_28733,N_28264);
nand U29053 (N_29053,N_28677,N_28539);
and U29054 (N_29054,N_28583,N_28609);
nor U29055 (N_29055,N_28729,N_28280);
nor U29056 (N_29056,N_28646,N_28225);
nand U29057 (N_29057,N_28296,N_28211);
nand U29058 (N_29058,N_28788,N_28660);
and U29059 (N_29059,N_28408,N_28616);
nor U29060 (N_29060,N_28223,N_28565);
or U29061 (N_29061,N_28319,N_28337);
or U29062 (N_29062,N_28520,N_28747);
nor U29063 (N_29063,N_28596,N_28786);
or U29064 (N_29064,N_28749,N_28496);
and U29065 (N_29065,N_28390,N_28241);
or U29066 (N_29066,N_28698,N_28626);
nor U29067 (N_29067,N_28373,N_28357);
nor U29068 (N_29068,N_28602,N_28643);
or U29069 (N_29069,N_28480,N_28593);
or U29070 (N_29070,N_28221,N_28768);
and U29071 (N_29071,N_28711,N_28372);
nor U29072 (N_29072,N_28575,N_28206);
nand U29073 (N_29073,N_28564,N_28202);
or U29074 (N_29074,N_28397,N_28411);
or U29075 (N_29075,N_28401,N_28714);
nor U29076 (N_29076,N_28336,N_28427);
nand U29077 (N_29077,N_28382,N_28430);
or U29078 (N_29078,N_28413,N_28339);
or U29079 (N_29079,N_28627,N_28571);
nand U29080 (N_29080,N_28668,N_28407);
and U29081 (N_29081,N_28255,N_28757);
and U29082 (N_29082,N_28516,N_28489);
or U29083 (N_29083,N_28696,N_28398);
nor U29084 (N_29084,N_28488,N_28558);
and U29085 (N_29085,N_28659,N_28515);
nor U29086 (N_29086,N_28464,N_28654);
nand U29087 (N_29087,N_28687,N_28579);
and U29088 (N_29088,N_28746,N_28493);
or U29089 (N_29089,N_28441,N_28250);
xor U29090 (N_29090,N_28567,N_28767);
nor U29091 (N_29091,N_28777,N_28672);
nor U29092 (N_29092,N_28270,N_28725);
xnor U29093 (N_29093,N_28524,N_28412);
xnor U29094 (N_29094,N_28371,N_28550);
xnor U29095 (N_29095,N_28705,N_28350);
nand U29096 (N_29096,N_28773,N_28485);
nand U29097 (N_29097,N_28226,N_28701);
nand U29098 (N_29098,N_28230,N_28355);
or U29099 (N_29099,N_28418,N_28234);
or U29100 (N_29100,N_28589,N_28225);
nor U29101 (N_29101,N_28688,N_28361);
xnor U29102 (N_29102,N_28424,N_28299);
and U29103 (N_29103,N_28234,N_28731);
nor U29104 (N_29104,N_28307,N_28727);
xor U29105 (N_29105,N_28700,N_28286);
or U29106 (N_29106,N_28516,N_28284);
nor U29107 (N_29107,N_28477,N_28490);
nor U29108 (N_29108,N_28202,N_28605);
xor U29109 (N_29109,N_28232,N_28641);
or U29110 (N_29110,N_28364,N_28722);
nand U29111 (N_29111,N_28621,N_28200);
or U29112 (N_29112,N_28224,N_28527);
or U29113 (N_29113,N_28520,N_28614);
and U29114 (N_29114,N_28539,N_28626);
or U29115 (N_29115,N_28591,N_28712);
nand U29116 (N_29116,N_28648,N_28232);
and U29117 (N_29117,N_28769,N_28764);
nand U29118 (N_29118,N_28621,N_28693);
xor U29119 (N_29119,N_28318,N_28683);
and U29120 (N_29120,N_28223,N_28528);
xnor U29121 (N_29121,N_28454,N_28242);
xnor U29122 (N_29122,N_28557,N_28449);
and U29123 (N_29123,N_28437,N_28756);
and U29124 (N_29124,N_28796,N_28239);
and U29125 (N_29125,N_28432,N_28771);
nand U29126 (N_29126,N_28229,N_28378);
and U29127 (N_29127,N_28433,N_28612);
and U29128 (N_29128,N_28754,N_28753);
nor U29129 (N_29129,N_28517,N_28767);
nand U29130 (N_29130,N_28493,N_28468);
nor U29131 (N_29131,N_28357,N_28493);
xnor U29132 (N_29132,N_28756,N_28421);
nand U29133 (N_29133,N_28235,N_28207);
or U29134 (N_29134,N_28419,N_28381);
or U29135 (N_29135,N_28654,N_28670);
nor U29136 (N_29136,N_28627,N_28684);
nand U29137 (N_29137,N_28484,N_28549);
and U29138 (N_29138,N_28791,N_28408);
nand U29139 (N_29139,N_28241,N_28598);
nand U29140 (N_29140,N_28725,N_28312);
nor U29141 (N_29141,N_28329,N_28651);
nand U29142 (N_29142,N_28677,N_28299);
nand U29143 (N_29143,N_28542,N_28425);
nor U29144 (N_29144,N_28699,N_28390);
nor U29145 (N_29145,N_28512,N_28264);
nand U29146 (N_29146,N_28289,N_28538);
or U29147 (N_29147,N_28769,N_28561);
nand U29148 (N_29148,N_28409,N_28430);
nor U29149 (N_29149,N_28736,N_28616);
and U29150 (N_29150,N_28404,N_28311);
or U29151 (N_29151,N_28243,N_28672);
xor U29152 (N_29152,N_28798,N_28704);
or U29153 (N_29153,N_28305,N_28333);
and U29154 (N_29154,N_28272,N_28688);
xor U29155 (N_29155,N_28499,N_28223);
and U29156 (N_29156,N_28622,N_28481);
and U29157 (N_29157,N_28719,N_28380);
nand U29158 (N_29158,N_28530,N_28587);
nand U29159 (N_29159,N_28696,N_28377);
nand U29160 (N_29160,N_28593,N_28471);
or U29161 (N_29161,N_28432,N_28423);
and U29162 (N_29162,N_28409,N_28237);
and U29163 (N_29163,N_28555,N_28243);
xor U29164 (N_29164,N_28388,N_28590);
xor U29165 (N_29165,N_28426,N_28203);
nor U29166 (N_29166,N_28433,N_28720);
xnor U29167 (N_29167,N_28570,N_28553);
or U29168 (N_29168,N_28252,N_28364);
nor U29169 (N_29169,N_28460,N_28302);
nor U29170 (N_29170,N_28221,N_28263);
or U29171 (N_29171,N_28478,N_28598);
nand U29172 (N_29172,N_28685,N_28369);
nor U29173 (N_29173,N_28694,N_28277);
or U29174 (N_29174,N_28573,N_28489);
and U29175 (N_29175,N_28722,N_28597);
nand U29176 (N_29176,N_28307,N_28257);
or U29177 (N_29177,N_28474,N_28791);
or U29178 (N_29178,N_28523,N_28339);
nor U29179 (N_29179,N_28400,N_28540);
or U29180 (N_29180,N_28637,N_28499);
or U29181 (N_29181,N_28657,N_28502);
nand U29182 (N_29182,N_28710,N_28480);
or U29183 (N_29183,N_28416,N_28574);
and U29184 (N_29184,N_28224,N_28799);
xnor U29185 (N_29185,N_28628,N_28312);
or U29186 (N_29186,N_28533,N_28590);
or U29187 (N_29187,N_28285,N_28398);
nor U29188 (N_29188,N_28769,N_28452);
xor U29189 (N_29189,N_28770,N_28591);
nand U29190 (N_29190,N_28580,N_28600);
and U29191 (N_29191,N_28270,N_28532);
xor U29192 (N_29192,N_28288,N_28541);
nand U29193 (N_29193,N_28691,N_28515);
nor U29194 (N_29194,N_28736,N_28310);
nor U29195 (N_29195,N_28324,N_28458);
xor U29196 (N_29196,N_28504,N_28590);
or U29197 (N_29197,N_28311,N_28474);
or U29198 (N_29198,N_28356,N_28349);
or U29199 (N_29199,N_28727,N_28554);
xor U29200 (N_29200,N_28330,N_28755);
and U29201 (N_29201,N_28626,N_28357);
xor U29202 (N_29202,N_28520,N_28444);
xnor U29203 (N_29203,N_28702,N_28366);
xor U29204 (N_29204,N_28417,N_28575);
and U29205 (N_29205,N_28573,N_28296);
xnor U29206 (N_29206,N_28381,N_28596);
nand U29207 (N_29207,N_28678,N_28737);
xnor U29208 (N_29208,N_28404,N_28682);
nor U29209 (N_29209,N_28536,N_28348);
and U29210 (N_29210,N_28273,N_28571);
xor U29211 (N_29211,N_28254,N_28280);
xnor U29212 (N_29212,N_28338,N_28368);
and U29213 (N_29213,N_28339,N_28375);
nor U29214 (N_29214,N_28734,N_28406);
or U29215 (N_29215,N_28647,N_28247);
nor U29216 (N_29216,N_28503,N_28324);
or U29217 (N_29217,N_28537,N_28515);
or U29218 (N_29218,N_28716,N_28779);
xnor U29219 (N_29219,N_28599,N_28292);
or U29220 (N_29220,N_28698,N_28642);
or U29221 (N_29221,N_28792,N_28411);
nand U29222 (N_29222,N_28737,N_28771);
and U29223 (N_29223,N_28677,N_28384);
or U29224 (N_29224,N_28392,N_28427);
xor U29225 (N_29225,N_28296,N_28464);
nor U29226 (N_29226,N_28721,N_28638);
and U29227 (N_29227,N_28752,N_28314);
and U29228 (N_29228,N_28554,N_28785);
nand U29229 (N_29229,N_28643,N_28719);
nand U29230 (N_29230,N_28646,N_28200);
xnor U29231 (N_29231,N_28447,N_28454);
nand U29232 (N_29232,N_28620,N_28293);
or U29233 (N_29233,N_28281,N_28464);
and U29234 (N_29234,N_28615,N_28416);
or U29235 (N_29235,N_28786,N_28335);
or U29236 (N_29236,N_28797,N_28768);
nand U29237 (N_29237,N_28784,N_28685);
nor U29238 (N_29238,N_28730,N_28753);
or U29239 (N_29239,N_28398,N_28294);
nand U29240 (N_29240,N_28260,N_28671);
xor U29241 (N_29241,N_28205,N_28518);
nor U29242 (N_29242,N_28461,N_28596);
nor U29243 (N_29243,N_28204,N_28480);
or U29244 (N_29244,N_28520,N_28423);
nor U29245 (N_29245,N_28781,N_28557);
nand U29246 (N_29246,N_28487,N_28603);
nor U29247 (N_29247,N_28745,N_28631);
nor U29248 (N_29248,N_28426,N_28687);
and U29249 (N_29249,N_28552,N_28712);
nand U29250 (N_29250,N_28339,N_28344);
nand U29251 (N_29251,N_28242,N_28277);
or U29252 (N_29252,N_28618,N_28237);
nor U29253 (N_29253,N_28263,N_28497);
nand U29254 (N_29254,N_28236,N_28530);
and U29255 (N_29255,N_28596,N_28726);
nand U29256 (N_29256,N_28594,N_28557);
nand U29257 (N_29257,N_28626,N_28795);
nand U29258 (N_29258,N_28268,N_28482);
nor U29259 (N_29259,N_28796,N_28338);
xnor U29260 (N_29260,N_28311,N_28296);
nor U29261 (N_29261,N_28353,N_28303);
or U29262 (N_29262,N_28461,N_28400);
or U29263 (N_29263,N_28572,N_28469);
nand U29264 (N_29264,N_28239,N_28740);
nand U29265 (N_29265,N_28224,N_28760);
xnor U29266 (N_29266,N_28752,N_28708);
xor U29267 (N_29267,N_28297,N_28541);
nor U29268 (N_29268,N_28313,N_28286);
nand U29269 (N_29269,N_28757,N_28414);
and U29270 (N_29270,N_28629,N_28410);
xnor U29271 (N_29271,N_28335,N_28414);
or U29272 (N_29272,N_28592,N_28287);
or U29273 (N_29273,N_28575,N_28460);
xnor U29274 (N_29274,N_28730,N_28576);
or U29275 (N_29275,N_28486,N_28742);
xnor U29276 (N_29276,N_28213,N_28369);
nand U29277 (N_29277,N_28648,N_28563);
nand U29278 (N_29278,N_28271,N_28740);
nor U29279 (N_29279,N_28349,N_28572);
nor U29280 (N_29280,N_28689,N_28509);
nand U29281 (N_29281,N_28770,N_28434);
nand U29282 (N_29282,N_28294,N_28455);
and U29283 (N_29283,N_28513,N_28355);
or U29284 (N_29284,N_28580,N_28435);
nand U29285 (N_29285,N_28571,N_28221);
nand U29286 (N_29286,N_28691,N_28728);
nor U29287 (N_29287,N_28397,N_28774);
and U29288 (N_29288,N_28317,N_28789);
and U29289 (N_29289,N_28409,N_28687);
and U29290 (N_29290,N_28504,N_28652);
xor U29291 (N_29291,N_28425,N_28735);
nand U29292 (N_29292,N_28751,N_28642);
and U29293 (N_29293,N_28432,N_28414);
or U29294 (N_29294,N_28735,N_28415);
or U29295 (N_29295,N_28475,N_28298);
or U29296 (N_29296,N_28444,N_28717);
nand U29297 (N_29297,N_28585,N_28798);
nand U29298 (N_29298,N_28723,N_28458);
and U29299 (N_29299,N_28454,N_28519);
and U29300 (N_29300,N_28484,N_28608);
nor U29301 (N_29301,N_28424,N_28626);
xnor U29302 (N_29302,N_28479,N_28688);
xor U29303 (N_29303,N_28415,N_28456);
or U29304 (N_29304,N_28290,N_28744);
or U29305 (N_29305,N_28700,N_28402);
nand U29306 (N_29306,N_28719,N_28680);
nand U29307 (N_29307,N_28372,N_28453);
xnor U29308 (N_29308,N_28257,N_28236);
nor U29309 (N_29309,N_28733,N_28271);
xor U29310 (N_29310,N_28262,N_28477);
and U29311 (N_29311,N_28340,N_28274);
nor U29312 (N_29312,N_28571,N_28325);
nor U29313 (N_29313,N_28225,N_28617);
nand U29314 (N_29314,N_28673,N_28598);
xnor U29315 (N_29315,N_28406,N_28259);
nand U29316 (N_29316,N_28250,N_28505);
xnor U29317 (N_29317,N_28507,N_28571);
xor U29318 (N_29318,N_28342,N_28576);
nand U29319 (N_29319,N_28719,N_28663);
and U29320 (N_29320,N_28722,N_28443);
nor U29321 (N_29321,N_28311,N_28343);
nand U29322 (N_29322,N_28320,N_28210);
nor U29323 (N_29323,N_28271,N_28227);
xor U29324 (N_29324,N_28336,N_28776);
and U29325 (N_29325,N_28638,N_28438);
nor U29326 (N_29326,N_28213,N_28203);
nand U29327 (N_29327,N_28378,N_28559);
and U29328 (N_29328,N_28501,N_28689);
nor U29329 (N_29329,N_28435,N_28745);
xnor U29330 (N_29330,N_28470,N_28503);
nand U29331 (N_29331,N_28780,N_28700);
xnor U29332 (N_29332,N_28525,N_28215);
xnor U29333 (N_29333,N_28736,N_28446);
or U29334 (N_29334,N_28497,N_28741);
and U29335 (N_29335,N_28467,N_28423);
nand U29336 (N_29336,N_28286,N_28556);
nor U29337 (N_29337,N_28469,N_28567);
nand U29338 (N_29338,N_28516,N_28764);
and U29339 (N_29339,N_28428,N_28755);
or U29340 (N_29340,N_28377,N_28302);
nor U29341 (N_29341,N_28529,N_28711);
or U29342 (N_29342,N_28370,N_28796);
xor U29343 (N_29343,N_28239,N_28237);
xor U29344 (N_29344,N_28546,N_28269);
or U29345 (N_29345,N_28389,N_28243);
nor U29346 (N_29346,N_28286,N_28754);
xor U29347 (N_29347,N_28207,N_28545);
xor U29348 (N_29348,N_28422,N_28700);
nor U29349 (N_29349,N_28292,N_28208);
or U29350 (N_29350,N_28667,N_28293);
nor U29351 (N_29351,N_28780,N_28708);
xor U29352 (N_29352,N_28390,N_28456);
nand U29353 (N_29353,N_28406,N_28599);
or U29354 (N_29354,N_28735,N_28310);
or U29355 (N_29355,N_28210,N_28652);
and U29356 (N_29356,N_28304,N_28628);
nor U29357 (N_29357,N_28665,N_28408);
and U29358 (N_29358,N_28304,N_28624);
nand U29359 (N_29359,N_28510,N_28753);
or U29360 (N_29360,N_28613,N_28768);
and U29361 (N_29361,N_28264,N_28583);
nand U29362 (N_29362,N_28368,N_28580);
nor U29363 (N_29363,N_28333,N_28415);
or U29364 (N_29364,N_28368,N_28414);
or U29365 (N_29365,N_28676,N_28585);
nor U29366 (N_29366,N_28731,N_28611);
or U29367 (N_29367,N_28339,N_28759);
nand U29368 (N_29368,N_28731,N_28322);
and U29369 (N_29369,N_28537,N_28442);
or U29370 (N_29370,N_28599,N_28207);
and U29371 (N_29371,N_28282,N_28772);
or U29372 (N_29372,N_28607,N_28269);
nand U29373 (N_29373,N_28380,N_28318);
xnor U29374 (N_29374,N_28668,N_28365);
and U29375 (N_29375,N_28207,N_28518);
nor U29376 (N_29376,N_28472,N_28627);
xnor U29377 (N_29377,N_28799,N_28546);
and U29378 (N_29378,N_28275,N_28570);
and U29379 (N_29379,N_28777,N_28710);
nand U29380 (N_29380,N_28437,N_28294);
nor U29381 (N_29381,N_28511,N_28543);
xor U29382 (N_29382,N_28311,N_28553);
nand U29383 (N_29383,N_28486,N_28285);
and U29384 (N_29384,N_28543,N_28513);
or U29385 (N_29385,N_28261,N_28404);
nor U29386 (N_29386,N_28646,N_28472);
or U29387 (N_29387,N_28399,N_28634);
xor U29388 (N_29388,N_28262,N_28476);
nor U29389 (N_29389,N_28618,N_28348);
xor U29390 (N_29390,N_28606,N_28640);
and U29391 (N_29391,N_28702,N_28688);
or U29392 (N_29392,N_28719,N_28245);
or U29393 (N_29393,N_28342,N_28499);
and U29394 (N_29394,N_28727,N_28530);
nor U29395 (N_29395,N_28310,N_28464);
nor U29396 (N_29396,N_28443,N_28223);
nor U29397 (N_29397,N_28302,N_28684);
or U29398 (N_29398,N_28590,N_28636);
and U29399 (N_29399,N_28322,N_28318);
nand U29400 (N_29400,N_29386,N_29117);
or U29401 (N_29401,N_28860,N_29321);
nand U29402 (N_29402,N_29052,N_29089);
nor U29403 (N_29403,N_29061,N_29300);
nor U29404 (N_29404,N_29056,N_28868);
or U29405 (N_29405,N_29265,N_29335);
and U29406 (N_29406,N_29088,N_29077);
nand U29407 (N_29407,N_29139,N_29241);
or U29408 (N_29408,N_29200,N_28960);
nor U29409 (N_29409,N_29282,N_29342);
nor U29410 (N_29410,N_28904,N_28878);
nand U29411 (N_29411,N_29155,N_28979);
or U29412 (N_29412,N_29186,N_29110);
and U29413 (N_29413,N_29344,N_28942);
nor U29414 (N_29414,N_28905,N_28973);
or U29415 (N_29415,N_28806,N_28836);
nor U29416 (N_29416,N_28914,N_29010);
nor U29417 (N_29417,N_28989,N_29387);
or U29418 (N_29418,N_29033,N_28978);
xor U29419 (N_29419,N_29041,N_29148);
nand U29420 (N_29420,N_29381,N_29390);
nor U29421 (N_29421,N_29246,N_28883);
nor U29422 (N_29422,N_28864,N_29190);
or U29423 (N_29423,N_29023,N_28801);
xor U29424 (N_29424,N_28893,N_29192);
and U29425 (N_29425,N_28928,N_29207);
xor U29426 (N_29426,N_29206,N_29328);
nor U29427 (N_29427,N_29244,N_29198);
nor U29428 (N_29428,N_28941,N_29007);
nand U29429 (N_29429,N_28911,N_29288);
nand U29430 (N_29430,N_28877,N_28940);
or U29431 (N_29431,N_28974,N_28968);
xor U29432 (N_29432,N_28885,N_28855);
nor U29433 (N_29433,N_28993,N_29039);
nor U29434 (N_29434,N_29219,N_29114);
nor U29435 (N_29435,N_28804,N_29369);
nor U29436 (N_29436,N_29374,N_29152);
nand U29437 (N_29437,N_29055,N_29256);
nor U29438 (N_29438,N_28998,N_29174);
xnor U29439 (N_29439,N_29296,N_29370);
or U29440 (N_29440,N_29120,N_28896);
nor U29441 (N_29441,N_29216,N_29281);
nand U29442 (N_29442,N_28972,N_28848);
and U29443 (N_29443,N_28943,N_29118);
nor U29444 (N_29444,N_29020,N_29225);
xor U29445 (N_29445,N_29022,N_29213);
nor U29446 (N_29446,N_29261,N_29323);
nor U29447 (N_29447,N_29326,N_29314);
nor U29448 (N_29448,N_28997,N_29310);
and U29449 (N_29449,N_29283,N_29157);
and U29450 (N_29450,N_29373,N_29294);
xor U29451 (N_29451,N_29030,N_29350);
nor U29452 (N_29452,N_28859,N_29129);
or U29453 (N_29453,N_29392,N_29170);
or U29454 (N_29454,N_29325,N_29000);
xnor U29455 (N_29455,N_29015,N_29204);
or U29456 (N_29456,N_29124,N_29247);
and U29457 (N_29457,N_29008,N_28976);
nor U29458 (N_29458,N_28892,N_28886);
or U29459 (N_29459,N_29107,N_29202);
nand U29460 (N_29460,N_29315,N_29329);
nor U29461 (N_29461,N_29222,N_28924);
xnor U29462 (N_29462,N_28839,N_28995);
nor U29463 (N_29463,N_28807,N_29371);
or U29464 (N_29464,N_29252,N_29357);
nor U29465 (N_29465,N_28994,N_29025);
nand U29466 (N_29466,N_29362,N_29218);
or U29467 (N_29467,N_28837,N_29229);
nand U29468 (N_29468,N_28831,N_29279);
and U29469 (N_29469,N_28948,N_28817);
or U29470 (N_29470,N_29049,N_29162);
nand U29471 (N_29471,N_29076,N_28984);
nand U29472 (N_29472,N_29084,N_29276);
xnor U29473 (N_29473,N_29193,N_29156);
nor U29474 (N_29474,N_28835,N_29340);
nor U29475 (N_29475,N_28996,N_28988);
or U29476 (N_29476,N_28956,N_28909);
and U29477 (N_29477,N_29073,N_29116);
or U29478 (N_29478,N_29201,N_29187);
or U29479 (N_29479,N_28854,N_29349);
and U29480 (N_29480,N_28844,N_29179);
and U29481 (N_29481,N_28800,N_29103);
xnor U29482 (N_29482,N_28918,N_28999);
or U29483 (N_29483,N_29345,N_29309);
nand U29484 (N_29484,N_29239,N_28919);
nor U29485 (N_29485,N_29299,N_29263);
and U29486 (N_29486,N_29368,N_29259);
or U29487 (N_29487,N_28805,N_29021);
nor U29488 (N_29488,N_29292,N_29062);
and U29489 (N_29489,N_29286,N_29348);
or U29490 (N_29490,N_28992,N_29150);
or U29491 (N_29491,N_29134,N_29237);
or U29492 (N_29492,N_29173,N_29178);
and U29493 (N_29493,N_29172,N_29255);
or U29494 (N_29494,N_28927,N_28857);
nor U29495 (N_29495,N_29228,N_28832);
xnor U29496 (N_29496,N_29014,N_29011);
xnor U29497 (N_29497,N_29379,N_28949);
nor U29498 (N_29498,N_29053,N_28810);
nand U29499 (N_29499,N_29135,N_29195);
nand U29500 (N_29500,N_29184,N_29017);
or U29501 (N_29501,N_29377,N_29306);
or U29502 (N_29502,N_29024,N_29127);
and U29503 (N_29503,N_28816,N_29060);
nor U29504 (N_29504,N_29128,N_29230);
and U29505 (N_29505,N_29217,N_29395);
or U29506 (N_29506,N_28964,N_29046);
and U29507 (N_29507,N_29075,N_29043);
nand U29508 (N_29508,N_28834,N_29199);
xnor U29509 (N_29509,N_29058,N_28841);
xnor U29510 (N_29510,N_29164,N_29316);
nand U29511 (N_29511,N_28921,N_28980);
xnor U29512 (N_29512,N_29019,N_28891);
xnor U29513 (N_29513,N_28966,N_28959);
nand U29514 (N_29514,N_29289,N_28845);
and U29515 (N_29515,N_29298,N_28953);
nor U29516 (N_29516,N_29269,N_28840);
nand U29517 (N_29517,N_29231,N_29066);
nand U29518 (N_29518,N_29018,N_29301);
nor U29519 (N_29519,N_28920,N_28982);
nor U29520 (N_29520,N_29074,N_29347);
nand U29521 (N_29521,N_29317,N_28900);
and U29522 (N_29522,N_29303,N_29208);
and U29523 (N_29523,N_29236,N_28873);
and U29524 (N_29524,N_28969,N_29376);
xnor U29525 (N_29525,N_29273,N_28818);
or U29526 (N_29526,N_29113,N_29092);
nor U29527 (N_29527,N_29346,N_28843);
xor U29528 (N_29528,N_29136,N_29224);
or U29529 (N_29529,N_29009,N_29048);
nor U29530 (N_29530,N_29050,N_28866);
or U29531 (N_29531,N_29338,N_29068);
nand U29532 (N_29532,N_29277,N_28881);
xor U29533 (N_29533,N_28879,N_28926);
xnor U29534 (N_29534,N_29057,N_29153);
xnor U29535 (N_29535,N_29069,N_28925);
nand U29536 (N_29536,N_29356,N_28929);
xor U29537 (N_29537,N_28954,N_29330);
nor U29538 (N_29538,N_29122,N_29151);
or U29539 (N_29539,N_28932,N_29284);
or U29540 (N_29540,N_29235,N_29214);
and U29541 (N_29541,N_29163,N_29095);
xnor U29542 (N_29542,N_29320,N_28910);
and U29543 (N_29543,N_29038,N_29394);
and U29544 (N_29544,N_28811,N_28906);
or U29545 (N_29545,N_29180,N_29313);
and U29546 (N_29546,N_29391,N_29005);
or U29547 (N_29547,N_28937,N_28901);
or U29548 (N_29548,N_29233,N_29154);
nor U29549 (N_29549,N_29091,N_28970);
nor U29550 (N_29550,N_28951,N_28902);
or U29551 (N_29551,N_29125,N_29258);
or U29552 (N_29552,N_29324,N_28829);
nand U29553 (N_29553,N_28962,N_29364);
and U29554 (N_29554,N_29027,N_29166);
nand U29555 (N_29555,N_29399,N_29396);
nor U29556 (N_29556,N_28852,N_29042);
or U29557 (N_29557,N_28803,N_29112);
xor U29558 (N_29558,N_29119,N_29319);
or U29559 (N_29559,N_29383,N_29177);
xnor U29560 (N_29560,N_29274,N_29086);
nand U29561 (N_29561,N_29140,N_28861);
or U29562 (N_29562,N_28944,N_29165);
xor U29563 (N_29563,N_28894,N_29251);
nor U29564 (N_29564,N_28912,N_29365);
nor U29565 (N_29565,N_29271,N_28820);
or U29566 (N_29566,N_29176,N_29266);
nor U29567 (N_29567,N_29045,N_28977);
nor U29568 (N_29568,N_29211,N_29013);
and U29569 (N_29569,N_29322,N_29267);
nor U29570 (N_29570,N_29249,N_28863);
nand U29571 (N_29571,N_28888,N_29026);
nand U29572 (N_29572,N_29070,N_28952);
nor U29573 (N_29573,N_28865,N_29106);
or U29574 (N_29574,N_29359,N_28819);
and U29575 (N_29575,N_29227,N_29308);
xnor U29576 (N_29576,N_29360,N_28853);
or U29577 (N_29577,N_29339,N_29367);
or U29578 (N_29578,N_29185,N_29147);
or U29579 (N_29579,N_29385,N_29078);
nand U29580 (N_29580,N_29232,N_28833);
xnor U29581 (N_29581,N_28822,N_28851);
xor U29582 (N_29582,N_29126,N_29366);
or U29583 (N_29583,N_29293,N_28975);
nand U29584 (N_29584,N_28828,N_29181);
nor U29585 (N_29585,N_29318,N_29253);
or U29586 (N_29586,N_29389,N_29380);
nor U29587 (N_29587,N_29245,N_28825);
or U29588 (N_29588,N_29397,N_29003);
or U29589 (N_29589,N_29002,N_29311);
or U29590 (N_29590,N_29096,N_29090);
or U29591 (N_29591,N_29260,N_29004);
nand U29592 (N_29592,N_28826,N_29130);
or U29593 (N_29593,N_28812,N_29372);
nand U29594 (N_29594,N_28827,N_28985);
nor U29595 (N_29595,N_28931,N_29093);
xor U29596 (N_29596,N_28933,N_28875);
and U29597 (N_29597,N_29209,N_28938);
xnor U29598 (N_29598,N_29132,N_29102);
nand U29599 (N_29599,N_29032,N_29071);
or U29600 (N_29600,N_29034,N_28809);
and U29601 (N_29601,N_28870,N_29109);
nor U29602 (N_29602,N_28903,N_29393);
nand U29603 (N_29603,N_28967,N_28813);
or U29604 (N_29604,N_29285,N_29333);
or U29605 (N_29605,N_29243,N_29115);
or U29606 (N_29606,N_29210,N_29072);
and U29607 (N_29607,N_29302,N_29234);
nand U29608 (N_29608,N_28830,N_29188);
nand U29609 (N_29609,N_29044,N_29137);
or U29610 (N_29610,N_28874,N_28815);
xnor U29611 (N_29611,N_29197,N_29221);
xnor U29612 (N_29612,N_29028,N_28930);
xnor U29613 (N_29613,N_29361,N_29238);
and U29614 (N_29614,N_28922,N_29029);
or U29615 (N_29615,N_29159,N_29341);
or U29616 (N_29616,N_29087,N_28939);
and U29617 (N_29617,N_29080,N_29171);
nand U29618 (N_29618,N_29035,N_29169);
nor U29619 (N_29619,N_29182,N_29270);
or U29620 (N_29620,N_29191,N_29220);
and U29621 (N_29621,N_29194,N_29079);
or U29622 (N_29622,N_28957,N_29099);
and U29623 (N_29623,N_29105,N_29353);
nand U29624 (N_29624,N_29250,N_28955);
nor U29625 (N_29625,N_28850,N_29336);
nor U29626 (N_29626,N_29226,N_29104);
or U29627 (N_29627,N_28983,N_29203);
nand U29628 (N_29628,N_28872,N_29031);
or U29629 (N_29629,N_29196,N_29142);
and U29630 (N_29630,N_29257,N_29354);
xnor U29631 (N_29631,N_28991,N_28838);
or U29632 (N_29632,N_28935,N_29145);
nor U29633 (N_29633,N_28907,N_28946);
xor U29634 (N_29634,N_28917,N_29059);
xnor U29635 (N_29635,N_28899,N_28971);
nand U29636 (N_29636,N_29146,N_29212);
nand U29637 (N_29637,N_28965,N_29141);
nand U29638 (N_29638,N_29175,N_28871);
nand U29639 (N_29639,N_28842,N_29268);
nand U29640 (N_29640,N_29355,N_29183);
and U29641 (N_29641,N_29307,N_29001);
xnor U29642 (N_29642,N_29272,N_29158);
and U29643 (N_29643,N_29312,N_29161);
xor U29644 (N_29644,N_28990,N_29398);
nand U29645 (N_29645,N_29168,N_28950);
or U29646 (N_29646,N_29264,N_29343);
xor U29647 (N_29647,N_29297,N_29280);
and U29648 (N_29648,N_28963,N_29144);
nand U29649 (N_29649,N_29351,N_29248);
or U29650 (N_29650,N_28802,N_29334);
or U29651 (N_29651,N_28889,N_28916);
or U29652 (N_29652,N_29240,N_28908);
or U29653 (N_29653,N_29123,N_29133);
nor U29654 (N_29654,N_29063,N_29082);
and U29655 (N_29655,N_29167,N_28814);
nor U29656 (N_29656,N_29384,N_29054);
nor U29657 (N_29657,N_28981,N_28867);
nand U29658 (N_29658,N_29006,N_29304);
xor U29659 (N_29659,N_29037,N_28876);
nand U29660 (N_29660,N_29331,N_29100);
xor U29661 (N_29661,N_29160,N_29388);
or U29662 (N_29662,N_29275,N_28823);
nand U29663 (N_29663,N_29083,N_29012);
and U29664 (N_29664,N_29205,N_28987);
xor U29665 (N_29665,N_28898,N_28934);
nand U29666 (N_29666,N_28895,N_28897);
xnor U29667 (N_29667,N_29149,N_28915);
nand U29668 (N_29668,N_28986,N_29067);
nand U29669 (N_29669,N_29295,N_29378);
or U29670 (N_29670,N_29036,N_29131);
or U29671 (N_29671,N_28869,N_28947);
nor U29672 (N_29672,N_29382,N_29094);
or U29673 (N_29673,N_28890,N_28884);
nand U29674 (N_29674,N_29101,N_28824);
and U29675 (N_29675,N_28923,N_29215);
and U29676 (N_29676,N_28847,N_29305);
xor U29677 (N_29677,N_28913,N_29064);
or U29678 (N_29678,N_29108,N_29121);
nand U29679 (N_29679,N_29352,N_29051);
nor U29680 (N_29680,N_28858,N_29040);
or U29681 (N_29681,N_28882,N_29111);
or U29682 (N_29682,N_29047,N_29337);
xor U29683 (N_29683,N_28846,N_29287);
and U29684 (N_29684,N_29097,N_29143);
and U29685 (N_29685,N_28856,N_28887);
nor U29686 (N_29686,N_29327,N_29085);
xnor U29687 (N_29687,N_28849,N_28821);
nand U29688 (N_29688,N_29290,N_29363);
nand U29689 (N_29689,N_28862,N_29223);
and U29690 (N_29690,N_29375,N_28936);
xnor U29691 (N_29691,N_29332,N_28880);
xnor U29692 (N_29692,N_29098,N_29065);
and U29693 (N_29693,N_29278,N_28808);
nor U29694 (N_29694,N_29358,N_29081);
or U29695 (N_29695,N_29291,N_28961);
nor U29696 (N_29696,N_28958,N_29189);
nor U29697 (N_29697,N_28945,N_29016);
xnor U29698 (N_29698,N_29242,N_29262);
nor U29699 (N_29699,N_29138,N_29254);
and U29700 (N_29700,N_28975,N_29319);
or U29701 (N_29701,N_28813,N_29022);
or U29702 (N_29702,N_28841,N_28867);
or U29703 (N_29703,N_29206,N_29253);
nor U29704 (N_29704,N_29351,N_29260);
or U29705 (N_29705,N_29056,N_28897);
xor U29706 (N_29706,N_29278,N_29328);
nand U29707 (N_29707,N_29008,N_29309);
nor U29708 (N_29708,N_28965,N_29338);
or U29709 (N_29709,N_29297,N_28855);
nor U29710 (N_29710,N_29084,N_29136);
xnor U29711 (N_29711,N_28844,N_29037);
nand U29712 (N_29712,N_28961,N_29265);
xnor U29713 (N_29713,N_29239,N_28960);
nor U29714 (N_29714,N_29367,N_29301);
and U29715 (N_29715,N_29027,N_29383);
and U29716 (N_29716,N_29089,N_28990);
nand U29717 (N_29717,N_28970,N_29147);
xnor U29718 (N_29718,N_29237,N_29066);
xor U29719 (N_29719,N_29210,N_29340);
nand U29720 (N_29720,N_28848,N_29180);
or U29721 (N_29721,N_28866,N_29192);
nor U29722 (N_29722,N_28977,N_28823);
xnor U29723 (N_29723,N_29049,N_28964);
nand U29724 (N_29724,N_28925,N_28947);
nand U29725 (N_29725,N_28854,N_28863);
and U29726 (N_29726,N_29223,N_29019);
nand U29727 (N_29727,N_29094,N_29305);
nor U29728 (N_29728,N_28980,N_28957);
and U29729 (N_29729,N_29163,N_28892);
nand U29730 (N_29730,N_29324,N_28845);
nor U29731 (N_29731,N_28979,N_29078);
and U29732 (N_29732,N_29005,N_28889);
and U29733 (N_29733,N_29165,N_29358);
or U29734 (N_29734,N_28975,N_29222);
and U29735 (N_29735,N_28946,N_29235);
and U29736 (N_29736,N_29009,N_28963);
and U29737 (N_29737,N_29169,N_29123);
xnor U29738 (N_29738,N_29136,N_28919);
nor U29739 (N_29739,N_29307,N_29025);
xnor U29740 (N_29740,N_29328,N_29234);
nand U29741 (N_29741,N_29247,N_29086);
xnor U29742 (N_29742,N_29320,N_28848);
or U29743 (N_29743,N_29107,N_29069);
nand U29744 (N_29744,N_29116,N_29279);
xnor U29745 (N_29745,N_29316,N_29240);
nand U29746 (N_29746,N_29343,N_28929);
nor U29747 (N_29747,N_29382,N_28885);
nand U29748 (N_29748,N_29134,N_28810);
xor U29749 (N_29749,N_28950,N_29336);
xnor U29750 (N_29750,N_29020,N_29346);
xnor U29751 (N_29751,N_29075,N_29134);
or U29752 (N_29752,N_29180,N_29315);
nand U29753 (N_29753,N_29102,N_29315);
nor U29754 (N_29754,N_29380,N_29214);
nand U29755 (N_29755,N_29241,N_29018);
xor U29756 (N_29756,N_29322,N_29245);
xor U29757 (N_29757,N_28889,N_29268);
nor U29758 (N_29758,N_29219,N_28904);
nand U29759 (N_29759,N_29277,N_28811);
nand U29760 (N_29760,N_28925,N_29334);
nor U29761 (N_29761,N_29221,N_29371);
xor U29762 (N_29762,N_29169,N_28815);
or U29763 (N_29763,N_28910,N_29048);
nor U29764 (N_29764,N_29012,N_29087);
or U29765 (N_29765,N_29293,N_28878);
and U29766 (N_29766,N_29182,N_29109);
or U29767 (N_29767,N_29331,N_28865);
or U29768 (N_29768,N_29267,N_29284);
xor U29769 (N_29769,N_29076,N_29011);
and U29770 (N_29770,N_28946,N_29390);
and U29771 (N_29771,N_29162,N_29094);
or U29772 (N_29772,N_28857,N_29236);
nand U29773 (N_29773,N_28932,N_28888);
and U29774 (N_29774,N_29357,N_29271);
xor U29775 (N_29775,N_29279,N_29122);
and U29776 (N_29776,N_29187,N_29350);
nand U29777 (N_29777,N_29125,N_29347);
xor U29778 (N_29778,N_29124,N_29346);
and U29779 (N_29779,N_29093,N_29376);
nand U29780 (N_29780,N_28873,N_28956);
and U29781 (N_29781,N_29293,N_29132);
or U29782 (N_29782,N_29004,N_28867);
nand U29783 (N_29783,N_29108,N_29390);
and U29784 (N_29784,N_29098,N_28981);
nand U29785 (N_29785,N_29373,N_29291);
xor U29786 (N_29786,N_29053,N_29370);
or U29787 (N_29787,N_28950,N_28944);
nor U29788 (N_29788,N_28996,N_29212);
nor U29789 (N_29789,N_29205,N_29304);
and U29790 (N_29790,N_28995,N_29397);
or U29791 (N_29791,N_28977,N_28946);
nor U29792 (N_29792,N_29091,N_29386);
nor U29793 (N_29793,N_29115,N_28902);
nand U29794 (N_29794,N_28959,N_28996);
nor U29795 (N_29795,N_29052,N_29302);
xor U29796 (N_29796,N_29088,N_29118);
nand U29797 (N_29797,N_28865,N_29268);
nand U29798 (N_29798,N_29115,N_29004);
xnor U29799 (N_29799,N_29243,N_29241);
xor U29800 (N_29800,N_28961,N_29394);
nand U29801 (N_29801,N_29319,N_29322);
nand U29802 (N_29802,N_29031,N_29265);
or U29803 (N_29803,N_29308,N_28976);
or U29804 (N_29804,N_29116,N_29077);
nor U29805 (N_29805,N_28992,N_28925);
nor U29806 (N_29806,N_29268,N_29198);
xor U29807 (N_29807,N_29048,N_29013);
nand U29808 (N_29808,N_29197,N_29347);
nand U29809 (N_29809,N_29078,N_29274);
or U29810 (N_29810,N_28817,N_29112);
nand U29811 (N_29811,N_29185,N_28897);
and U29812 (N_29812,N_28863,N_29022);
nand U29813 (N_29813,N_29090,N_29000);
xnor U29814 (N_29814,N_29360,N_29313);
and U29815 (N_29815,N_29262,N_29343);
nor U29816 (N_29816,N_29364,N_28909);
nand U29817 (N_29817,N_29299,N_29131);
or U29818 (N_29818,N_29073,N_28847);
nand U29819 (N_29819,N_29280,N_29108);
nor U29820 (N_29820,N_29349,N_28860);
or U29821 (N_29821,N_28811,N_29251);
nor U29822 (N_29822,N_29036,N_28906);
nor U29823 (N_29823,N_29398,N_29167);
and U29824 (N_29824,N_29319,N_29144);
or U29825 (N_29825,N_28803,N_29123);
and U29826 (N_29826,N_28947,N_29261);
xor U29827 (N_29827,N_29399,N_29019);
xnor U29828 (N_29828,N_28841,N_29162);
nand U29829 (N_29829,N_29373,N_29146);
nand U29830 (N_29830,N_29162,N_29096);
and U29831 (N_29831,N_28947,N_29123);
and U29832 (N_29832,N_28912,N_29298);
or U29833 (N_29833,N_29267,N_29353);
nor U29834 (N_29834,N_29150,N_29304);
nor U29835 (N_29835,N_29382,N_29032);
nand U29836 (N_29836,N_29391,N_29137);
xor U29837 (N_29837,N_29168,N_28826);
xor U29838 (N_29838,N_29024,N_29101);
xor U29839 (N_29839,N_28960,N_29082);
xor U29840 (N_29840,N_29136,N_29369);
or U29841 (N_29841,N_29288,N_29068);
nor U29842 (N_29842,N_29128,N_28928);
nor U29843 (N_29843,N_29398,N_28863);
and U29844 (N_29844,N_29349,N_29231);
nand U29845 (N_29845,N_29166,N_29367);
nand U29846 (N_29846,N_28864,N_29084);
or U29847 (N_29847,N_29277,N_29194);
nor U29848 (N_29848,N_29290,N_29015);
and U29849 (N_29849,N_29230,N_29218);
or U29850 (N_29850,N_29043,N_29138);
xnor U29851 (N_29851,N_29322,N_29077);
nand U29852 (N_29852,N_29216,N_28828);
nor U29853 (N_29853,N_29051,N_28898);
nor U29854 (N_29854,N_29048,N_29298);
nor U29855 (N_29855,N_28953,N_29066);
and U29856 (N_29856,N_29038,N_28850);
nand U29857 (N_29857,N_29272,N_29315);
nand U29858 (N_29858,N_29279,N_29241);
and U29859 (N_29859,N_29227,N_29128);
nand U29860 (N_29860,N_29159,N_28907);
and U29861 (N_29861,N_29278,N_28982);
xnor U29862 (N_29862,N_29320,N_29103);
and U29863 (N_29863,N_29042,N_29376);
nand U29864 (N_29864,N_28970,N_28956);
or U29865 (N_29865,N_29213,N_29141);
xnor U29866 (N_29866,N_29018,N_29201);
and U29867 (N_29867,N_28878,N_29141);
or U29868 (N_29868,N_29169,N_28963);
xor U29869 (N_29869,N_29063,N_29227);
nor U29870 (N_29870,N_29015,N_29392);
nor U29871 (N_29871,N_28848,N_29162);
xor U29872 (N_29872,N_29368,N_29059);
and U29873 (N_29873,N_29121,N_29097);
or U29874 (N_29874,N_29076,N_28881);
nand U29875 (N_29875,N_29299,N_28899);
and U29876 (N_29876,N_28941,N_29238);
and U29877 (N_29877,N_28976,N_29072);
xnor U29878 (N_29878,N_28894,N_29257);
nor U29879 (N_29879,N_28816,N_29137);
or U29880 (N_29880,N_28817,N_28972);
xor U29881 (N_29881,N_29047,N_29218);
or U29882 (N_29882,N_28965,N_28875);
nand U29883 (N_29883,N_29161,N_29172);
nor U29884 (N_29884,N_29080,N_29308);
and U29885 (N_29885,N_29345,N_28996);
or U29886 (N_29886,N_29347,N_29089);
nor U29887 (N_29887,N_29345,N_29370);
nor U29888 (N_29888,N_29362,N_29035);
nor U29889 (N_29889,N_29371,N_29010);
xnor U29890 (N_29890,N_29132,N_29015);
xnor U29891 (N_29891,N_28842,N_29088);
and U29892 (N_29892,N_29329,N_29320);
nor U29893 (N_29893,N_29027,N_29121);
or U29894 (N_29894,N_29170,N_29299);
xnor U29895 (N_29895,N_28916,N_28870);
and U29896 (N_29896,N_29088,N_28912);
nor U29897 (N_29897,N_28893,N_28878);
nand U29898 (N_29898,N_28876,N_29219);
nand U29899 (N_29899,N_29376,N_29291);
or U29900 (N_29900,N_29131,N_29276);
nand U29901 (N_29901,N_29015,N_29371);
or U29902 (N_29902,N_29234,N_28952);
xnor U29903 (N_29903,N_29316,N_29278);
xnor U29904 (N_29904,N_29030,N_29178);
or U29905 (N_29905,N_28904,N_29238);
xnor U29906 (N_29906,N_29039,N_29358);
or U29907 (N_29907,N_29175,N_29348);
nand U29908 (N_29908,N_29049,N_28917);
or U29909 (N_29909,N_29264,N_29300);
nand U29910 (N_29910,N_29210,N_29260);
and U29911 (N_29911,N_29237,N_28866);
or U29912 (N_29912,N_29282,N_29061);
and U29913 (N_29913,N_28955,N_29079);
or U29914 (N_29914,N_29097,N_29149);
xnor U29915 (N_29915,N_29063,N_29307);
and U29916 (N_29916,N_29303,N_28976);
xor U29917 (N_29917,N_28931,N_29067);
nor U29918 (N_29918,N_29130,N_28801);
nand U29919 (N_29919,N_28823,N_29167);
nand U29920 (N_29920,N_29287,N_29142);
nand U29921 (N_29921,N_29267,N_28834);
nor U29922 (N_29922,N_28936,N_29051);
xnor U29923 (N_29923,N_29141,N_28993);
nand U29924 (N_29924,N_29065,N_28950);
xnor U29925 (N_29925,N_29030,N_29089);
nor U29926 (N_29926,N_28972,N_29128);
or U29927 (N_29927,N_29391,N_29105);
nor U29928 (N_29928,N_29248,N_28957);
and U29929 (N_29929,N_28973,N_29219);
or U29930 (N_29930,N_29045,N_28860);
and U29931 (N_29931,N_28879,N_29283);
and U29932 (N_29932,N_28993,N_29349);
nor U29933 (N_29933,N_29010,N_29194);
or U29934 (N_29934,N_29317,N_29118);
or U29935 (N_29935,N_28953,N_29350);
xnor U29936 (N_29936,N_29062,N_29367);
nand U29937 (N_29937,N_28834,N_29080);
and U29938 (N_29938,N_29231,N_28875);
nor U29939 (N_29939,N_29398,N_29178);
nor U29940 (N_29940,N_28889,N_29253);
xnor U29941 (N_29941,N_29317,N_28952);
nor U29942 (N_29942,N_28879,N_28890);
or U29943 (N_29943,N_29124,N_29273);
xnor U29944 (N_29944,N_29386,N_28861);
and U29945 (N_29945,N_28842,N_29060);
and U29946 (N_29946,N_28894,N_29334);
xor U29947 (N_29947,N_28919,N_29058);
xnor U29948 (N_29948,N_28808,N_29063);
and U29949 (N_29949,N_29158,N_28814);
or U29950 (N_29950,N_29126,N_29224);
and U29951 (N_29951,N_28861,N_28952);
and U29952 (N_29952,N_29382,N_29368);
nor U29953 (N_29953,N_29042,N_29267);
and U29954 (N_29954,N_28874,N_29201);
and U29955 (N_29955,N_28849,N_29271);
and U29956 (N_29956,N_29386,N_29112);
or U29957 (N_29957,N_29022,N_28998);
nor U29958 (N_29958,N_29179,N_29152);
nor U29959 (N_29959,N_28816,N_29206);
xnor U29960 (N_29960,N_29067,N_29362);
and U29961 (N_29961,N_29052,N_29247);
nand U29962 (N_29962,N_28801,N_29085);
xor U29963 (N_29963,N_29008,N_29086);
or U29964 (N_29964,N_29202,N_29050);
or U29965 (N_29965,N_28844,N_29060);
nor U29966 (N_29966,N_29208,N_29337);
or U29967 (N_29967,N_28903,N_29229);
or U29968 (N_29968,N_29237,N_29081);
nand U29969 (N_29969,N_29168,N_29041);
or U29970 (N_29970,N_29104,N_28946);
xor U29971 (N_29971,N_28995,N_28810);
xnor U29972 (N_29972,N_29291,N_29221);
nor U29973 (N_29973,N_29266,N_28846);
and U29974 (N_29974,N_28998,N_29027);
xnor U29975 (N_29975,N_29025,N_29262);
nand U29976 (N_29976,N_29143,N_29162);
nor U29977 (N_29977,N_29222,N_28903);
nor U29978 (N_29978,N_29277,N_29328);
nand U29979 (N_29979,N_29303,N_29384);
xor U29980 (N_29980,N_29028,N_29029);
xor U29981 (N_29981,N_28979,N_29186);
nor U29982 (N_29982,N_29271,N_28941);
or U29983 (N_29983,N_28968,N_28872);
xnor U29984 (N_29984,N_29153,N_29078);
or U29985 (N_29985,N_29092,N_28820);
xnor U29986 (N_29986,N_29373,N_28943);
or U29987 (N_29987,N_29270,N_29107);
and U29988 (N_29988,N_28896,N_29342);
nand U29989 (N_29989,N_28837,N_28862);
and U29990 (N_29990,N_29237,N_29356);
or U29991 (N_29991,N_29163,N_28916);
nand U29992 (N_29992,N_28999,N_29356);
xnor U29993 (N_29993,N_29354,N_29305);
or U29994 (N_29994,N_28855,N_29128);
nand U29995 (N_29995,N_29190,N_29069);
nor U29996 (N_29996,N_28805,N_29372);
xnor U29997 (N_29997,N_28878,N_29320);
nor U29998 (N_29998,N_29028,N_29303);
nor U29999 (N_29999,N_28859,N_28803);
nand UO_0 (O_0,N_29555,N_29715);
nand UO_1 (O_1,N_29630,N_29881);
or UO_2 (O_2,N_29955,N_29776);
or UO_3 (O_3,N_29459,N_29569);
and UO_4 (O_4,N_29949,N_29452);
or UO_5 (O_5,N_29573,N_29581);
or UO_6 (O_6,N_29787,N_29904);
or UO_7 (O_7,N_29481,N_29863);
and UO_8 (O_8,N_29731,N_29844);
and UO_9 (O_9,N_29862,N_29605);
or UO_10 (O_10,N_29436,N_29603);
and UO_11 (O_11,N_29465,N_29400);
xnor UO_12 (O_12,N_29695,N_29855);
nor UO_13 (O_13,N_29655,N_29757);
or UO_14 (O_14,N_29914,N_29667);
or UO_15 (O_15,N_29568,N_29824);
nand UO_16 (O_16,N_29642,N_29554);
xor UO_17 (O_17,N_29438,N_29446);
or UO_18 (O_18,N_29689,N_29781);
nor UO_19 (O_19,N_29976,N_29876);
nor UO_20 (O_20,N_29526,N_29745);
nand UO_21 (O_21,N_29448,N_29780);
nor UO_22 (O_22,N_29579,N_29531);
nor UO_23 (O_23,N_29494,N_29430);
xnor UO_24 (O_24,N_29996,N_29724);
or UO_25 (O_25,N_29434,N_29616);
nand UO_26 (O_26,N_29671,N_29702);
or UO_27 (O_27,N_29815,N_29545);
or UO_28 (O_28,N_29500,N_29962);
xor UO_29 (O_29,N_29482,N_29468);
nand UO_30 (O_30,N_29750,N_29574);
nand UO_31 (O_31,N_29547,N_29674);
nor UO_32 (O_32,N_29889,N_29618);
or UO_33 (O_33,N_29931,N_29773);
nor UO_34 (O_34,N_29930,N_29402);
nor UO_35 (O_35,N_29980,N_29946);
and UO_36 (O_36,N_29758,N_29622);
nand UO_37 (O_37,N_29754,N_29585);
and UO_38 (O_38,N_29917,N_29772);
or UO_39 (O_39,N_29846,N_29840);
nand UO_40 (O_40,N_29453,N_29471);
xor UO_41 (O_41,N_29788,N_29417);
and UO_42 (O_42,N_29782,N_29937);
nand UO_43 (O_43,N_29463,N_29498);
and UO_44 (O_44,N_29928,N_29886);
and UO_45 (O_45,N_29948,N_29943);
xnor UO_46 (O_46,N_29519,N_29462);
or UO_47 (O_47,N_29791,N_29419);
nand UO_48 (O_48,N_29550,N_29884);
or UO_49 (O_49,N_29813,N_29838);
or UO_50 (O_50,N_29627,N_29795);
nor UO_51 (O_51,N_29546,N_29756);
xor UO_52 (O_52,N_29637,N_29493);
and UO_53 (O_53,N_29720,N_29940);
nand UO_54 (O_54,N_29877,N_29563);
and UO_55 (O_55,N_29523,N_29464);
nor UO_56 (O_56,N_29577,N_29693);
nor UO_57 (O_57,N_29615,N_29990);
xnor UO_58 (O_58,N_29918,N_29764);
xnor UO_59 (O_59,N_29413,N_29852);
xor UO_60 (O_60,N_29658,N_29892);
nor UO_61 (O_61,N_29847,N_29851);
and UO_62 (O_62,N_29979,N_29822);
nand UO_63 (O_63,N_29460,N_29437);
or UO_64 (O_64,N_29698,N_29708);
nor UO_65 (O_65,N_29933,N_29817);
and UO_66 (O_66,N_29684,N_29888);
nand UO_67 (O_67,N_29625,N_29935);
xor UO_68 (O_68,N_29898,N_29520);
or UO_69 (O_69,N_29488,N_29834);
xor UO_70 (O_70,N_29461,N_29534);
nor UO_71 (O_71,N_29726,N_29811);
or UO_72 (O_72,N_29763,N_29429);
nand UO_73 (O_73,N_29447,N_29511);
nand UO_74 (O_74,N_29502,N_29723);
xor UO_75 (O_75,N_29418,N_29475);
nor UO_76 (O_76,N_29826,N_29639);
or UO_77 (O_77,N_29845,N_29633);
or UO_78 (O_78,N_29727,N_29414);
nand UO_79 (O_79,N_29919,N_29623);
nand UO_80 (O_80,N_29730,N_29985);
xor UO_81 (O_81,N_29506,N_29472);
xnor UO_82 (O_82,N_29858,N_29964);
or UO_83 (O_83,N_29604,N_29653);
or UO_84 (O_84,N_29939,N_29590);
or UO_85 (O_85,N_29729,N_29528);
or UO_86 (O_86,N_29944,N_29607);
or UO_87 (O_87,N_29992,N_29882);
or UO_88 (O_88,N_29551,N_29536);
xnor UO_89 (O_89,N_29663,N_29451);
or UO_90 (O_90,N_29868,N_29995);
xnor UO_91 (O_91,N_29433,N_29539);
and UO_92 (O_92,N_29404,N_29982);
and UO_93 (O_93,N_29687,N_29476);
nand UO_94 (O_94,N_29784,N_29830);
and UO_95 (O_95,N_29945,N_29697);
or UO_96 (O_96,N_29856,N_29799);
xnor UO_97 (O_97,N_29905,N_29835);
nor UO_98 (O_98,N_29759,N_29983);
nand UO_99 (O_99,N_29975,N_29432);
and UO_100 (O_100,N_29941,N_29444);
xnor UO_101 (O_101,N_29443,N_29592);
nand UO_102 (O_102,N_29548,N_29412);
nand UO_103 (O_103,N_29602,N_29768);
xnor UO_104 (O_104,N_29848,N_29644);
or UO_105 (O_105,N_29825,N_29869);
xnor UO_106 (O_106,N_29790,N_29606);
nand UO_107 (O_107,N_29542,N_29609);
nand UO_108 (O_108,N_29612,N_29672);
or UO_109 (O_109,N_29679,N_29712);
or UO_110 (O_110,N_29969,N_29853);
or UO_111 (O_111,N_29911,N_29636);
and UO_112 (O_112,N_29860,N_29938);
nand UO_113 (O_113,N_29556,N_29427);
xor UO_114 (O_114,N_29805,N_29875);
nand UO_115 (O_115,N_29880,N_29613);
nor UO_116 (O_116,N_29755,N_29837);
nand UO_117 (O_117,N_29864,N_29713);
or UO_118 (O_118,N_29685,N_29797);
nand UO_119 (O_119,N_29973,N_29567);
or UO_120 (O_120,N_29497,N_29743);
and UO_121 (O_121,N_29582,N_29450);
nand UO_122 (O_122,N_29913,N_29651);
xor UO_123 (O_123,N_29711,N_29833);
xnor UO_124 (O_124,N_29587,N_29692);
or UO_125 (O_125,N_29491,N_29648);
nand UO_126 (O_126,N_29570,N_29871);
xnor UO_127 (O_127,N_29660,N_29704);
and UO_128 (O_128,N_29424,N_29705);
nor UO_129 (O_129,N_29934,N_29922);
nand UO_130 (O_130,N_29737,N_29649);
nand UO_131 (O_131,N_29971,N_29496);
and UO_132 (O_132,N_29495,N_29647);
and UO_133 (O_133,N_29564,N_29611);
nor UO_134 (O_134,N_29406,N_29421);
or UO_135 (O_135,N_29735,N_29678);
xor UO_136 (O_136,N_29707,N_29749);
nand UO_137 (O_137,N_29821,N_29593);
and UO_138 (O_138,N_29789,N_29690);
or UO_139 (O_139,N_29455,N_29652);
and UO_140 (O_140,N_29596,N_29956);
nand UO_141 (O_141,N_29832,N_29553);
nor UO_142 (O_142,N_29558,N_29703);
and UO_143 (O_143,N_29706,N_29986);
xor UO_144 (O_144,N_29410,N_29599);
or UO_145 (O_145,N_29540,N_29819);
nand UO_146 (O_146,N_29879,N_29909);
and UO_147 (O_147,N_29458,N_29796);
and UO_148 (O_148,N_29970,N_29640);
nor UO_149 (O_149,N_29747,N_29614);
nor UO_150 (O_150,N_29449,N_29890);
or UO_151 (O_151,N_29719,N_29489);
nor UO_152 (O_152,N_29870,N_29562);
nor UO_153 (O_153,N_29894,N_29510);
or UO_154 (O_154,N_29677,N_29798);
or UO_155 (O_155,N_29961,N_29978);
and UO_156 (O_156,N_29901,N_29699);
nand UO_157 (O_157,N_29896,N_29580);
nand UO_158 (O_158,N_29467,N_29859);
and UO_159 (O_159,N_29718,N_29897);
or UO_160 (O_160,N_29578,N_29765);
and UO_161 (O_161,N_29786,N_29575);
and UO_162 (O_162,N_29409,N_29408);
xnor UO_163 (O_163,N_29774,N_29802);
or UO_164 (O_164,N_29907,N_29664);
xnor UO_165 (O_165,N_29816,N_29895);
nor UO_166 (O_166,N_29586,N_29810);
and UO_167 (O_167,N_29900,N_29525);
nand UO_168 (O_168,N_29766,N_29537);
or UO_169 (O_169,N_29857,N_29974);
nor UO_170 (O_170,N_29942,N_29994);
or UO_171 (O_171,N_29801,N_29646);
or UO_172 (O_172,N_29591,N_29775);
xor UO_173 (O_173,N_29874,N_29908);
or UO_174 (O_174,N_29680,N_29626);
nor UO_175 (O_175,N_29479,N_29527);
or UO_176 (O_176,N_29501,N_29929);
xor UO_177 (O_177,N_29915,N_29522);
xnor UO_178 (O_178,N_29722,N_29507);
nor UO_179 (O_179,N_29829,N_29872);
nand UO_180 (O_180,N_29549,N_29921);
xnor UO_181 (O_181,N_29778,N_29617);
and UO_182 (O_182,N_29513,N_29405);
nand UO_183 (O_183,N_29624,N_29634);
or UO_184 (O_184,N_29899,N_29977);
or UO_185 (O_185,N_29841,N_29426);
nand UO_186 (O_186,N_29533,N_29411);
nand UO_187 (O_187,N_29748,N_29407);
nand UO_188 (O_188,N_29657,N_29682);
nor UO_189 (O_189,N_29661,N_29742);
nand UO_190 (O_190,N_29425,N_29621);
nor UO_191 (O_191,N_29836,N_29827);
xnor UO_192 (O_192,N_29650,N_29560);
or UO_193 (O_193,N_29435,N_29806);
nor UO_194 (O_194,N_29710,N_29668);
or UO_195 (O_195,N_29401,N_29454);
nor UO_196 (O_196,N_29998,N_29968);
nand UO_197 (O_197,N_29867,N_29769);
and UO_198 (O_198,N_29891,N_29800);
xor UO_199 (O_199,N_29508,N_29620);
or UO_200 (O_200,N_29878,N_29809);
and UO_201 (O_201,N_29484,N_29883);
nand UO_202 (O_202,N_29566,N_29594);
nor UO_203 (O_203,N_29512,N_29681);
and UO_204 (O_204,N_29839,N_29993);
nor UO_205 (O_205,N_29641,N_29807);
and UO_206 (O_206,N_29916,N_29486);
xor UO_207 (O_207,N_29721,N_29638);
or UO_208 (O_208,N_29598,N_29517);
nor UO_209 (O_209,N_29541,N_29457);
and UO_210 (O_210,N_29589,N_29632);
nor UO_211 (O_211,N_29873,N_29610);
and UO_212 (O_212,N_29984,N_29415);
and UO_213 (O_213,N_29988,N_29628);
or UO_214 (O_214,N_29499,N_29804);
or UO_215 (O_215,N_29544,N_29752);
xnor UO_216 (O_216,N_29910,N_29694);
or UO_217 (O_217,N_29893,N_29991);
xor UO_218 (O_218,N_29559,N_29673);
xnor UO_219 (O_219,N_29420,N_29843);
nor UO_220 (O_220,N_29584,N_29714);
or UO_221 (O_221,N_29902,N_29999);
nand UO_222 (O_222,N_29485,N_29503);
and UO_223 (O_223,N_29767,N_29732);
and UO_224 (O_224,N_29492,N_29963);
nor UO_225 (O_225,N_29989,N_29740);
or UO_226 (O_226,N_29473,N_29515);
or UO_227 (O_227,N_29588,N_29478);
nor UO_228 (O_228,N_29850,N_29717);
or UO_229 (O_229,N_29887,N_29656);
nor UO_230 (O_230,N_29514,N_29565);
or UO_231 (O_231,N_29770,N_29709);
or UO_232 (O_232,N_29854,N_29601);
and UO_233 (O_233,N_29659,N_29666);
and UO_234 (O_234,N_29700,N_29619);
and UO_235 (O_235,N_29771,N_29957);
xnor UO_236 (O_236,N_29716,N_29926);
xor UO_237 (O_237,N_29792,N_29529);
nand UO_238 (O_238,N_29952,N_29524);
nor UO_239 (O_239,N_29803,N_29812);
nand UO_240 (O_240,N_29865,N_29967);
xor UO_241 (O_241,N_29474,N_29981);
and UO_242 (O_242,N_29762,N_29814);
nand UO_243 (O_243,N_29932,N_29927);
and UO_244 (O_244,N_29431,N_29521);
nor UO_245 (O_245,N_29572,N_29728);
xor UO_246 (O_246,N_29849,N_29785);
and UO_247 (O_247,N_29987,N_29490);
and UO_248 (O_248,N_29631,N_29760);
xnor UO_249 (O_249,N_29483,N_29480);
nand UO_250 (O_250,N_29818,N_29997);
and UO_251 (O_251,N_29953,N_29783);
nor UO_252 (O_252,N_29794,N_29552);
xnor UO_253 (O_253,N_29543,N_29428);
nor UO_254 (O_254,N_29477,N_29885);
and UO_255 (O_255,N_29736,N_29532);
nor UO_256 (O_256,N_29793,N_29779);
and UO_257 (O_257,N_29403,N_29505);
and UO_258 (O_258,N_29777,N_29751);
and UO_259 (O_259,N_29441,N_29936);
nor UO_260 (O_260,N_29571,N_29823);
and UO_261 (O_261,N_29972,N_29906);
nand UO_262 (O_262,N_29456,N_29422);
nor UO_263 (O_263,N_29924,N_29958);
xor UO_264 (O_264,N_29920,N_29635);
xor UO_265 (O_265,N_29530,N_29960);
xor UO_266 (O_266,N_29516,N_29954);
nor UO_267 (O_267,N_29966,N_29959);
nor UO_268 (O_268,N_29746,N_29439);
nand UO_269 (O_269,N_29866,N_29608);
xnor UO_270 (O_270,N_29675,N_29669);
nor UO_271 (O_271,N_29665,N_29820);
nand UO_272 (O_272,N_29831,N_29595);
or UO_273 (O_273,N_29701,N_29691);
nand UO_274 (O_274,N_29738,N_29965);
or UO_275 (O_275,N_29753,N_29654);
and UO_276 (O_276,N_29416,N_29583);
or UO_277 (O_277,N_29629,N_29557);
xor UO_278 (O_278,N_29739,N_29442);
xnor UO_279 (O_279,N_29828,N_29733);
xnor UO_280 (O_280,N_29741,N_29861);
nor UO_281 (O_281,N_29662,N_29744);
nor UO_282 (O_282,N_29670,N_29469);
and UO_283 (O_283,N_29504,N_29561);
and UO_284 (O_284,N_29686,N_29734);
nand UO_285 (O_285,N_29538,N_29470);
and UO_286 (O_286,N_29912,N_29683);
nor UO_287 (O_287,N_29950,N_29597);
or UO_288 (O_288,N_29535,N_29440);
nor UO_289 (O_289,N_29761,N_29676);
nand UO_290 (O_290,N_29645,N_29925);
and UO_291 (O_291,N_29903,N_29518);
and UO_292 (O_292,N_29808,N_29923);
nand UO_293 (O_293,N_29951,N_29423);
nor UO_294 (O_294,N_29487,N_29643);
and UO_295 (O_295,N_29445,N_29842);
nand UO_296 (O_296,N_29600,N_29509);
or UO_297 (O_297,N_29725,N_29947);
or UO_298 (O_298,N_29466,N_29576);
xnor UO_299 (O_299,N_29688,N_29696);
nor UO_300 (O_300,N_29964,N_29600);
and UO_301 (O_301,N_29948,N_29601);
nor UO_302 (O_302,N_29575,N_29533);
nand UO_303 (O_303,N_29857,N_29477);
or UO_304 (O_304,N_29993,N_29894);
nor UO_305 (O_305,N_29615,N_29516);
nor UO_306 (O_306,N_29706,N_29776);
and UO_307 (O_307,N_29420,N_29985);
nor UO_308 (O_308,N_29671,N_29579);
nand UO_309 (O_309,N_29739,N_29853);
nor UO_310 (O_310,N_29490,N_29700);
nand UO_311 (O_311,N_29792,N_29603);
and UO_312 (O_312,N_29770,N_29455);
or UO_313 (O_313,N_29549,N_29617);
nor UO_314 (O_314,N_29790,N_29666);
xor UO_315 (O_315,N_29855,N_29506);
nor UO_316 (O_316,N_29425,N_29527);
xnor UO_317 (O_317,N_29677,N_29681);
xor UO_318 (O_318,N_29863,N_29860);
or UO_319 (O_319,N_29501,N_29590);
nand UO_320 (O_320,N_29688,N_29477);
or UO_321 (O_321,N_29703,N_29756);
nor UO_322 (O_322,N_29781,N_29941);
nand UO_323 (O_323,N_29494,N_29671);
nand UO_324 (O_324,N_29479,N_29483);
or UO_325 (O_325,N_29539,N_29445);
xnor UO_326 (O_326,N_29669,N_29702);
and UO_327 (O_327,N_29606,N_29858);
and UO_328 (O_328,N_29472,N_29603);
nand UO_329 (O_329,N_29911,N_29940);
nand UO_330 (O_330,N_29877,N_29473);
or UO_331 (O_331,N_29943,N_29496);
nand UO_332 (O_332,N_29953,N_29795);
nor UO_333 (O_333,N_29708,N_29679);
nor UO_334 (O_334,N_29780,N_29540);
nand UO_335 (O_335,N_29587,N_29922);
or UO_336 (O_336,N_29782,N_29635);
or UO_337 (O_337,N_29601,N_29730);
or UO_338 (O_338,N_29714,N_29999);
and UO_339 (O_339,N_29557,N_29408);
and UO_340 (O_340,N_29842,N_29835);
and UO_341 (O_341,N_29613,N_29743);
xor UO_342 (O_342,N_29626,N_29519);
or UO_343 (O_343,N_29783,N_29753);
and UO_344 (O_344,N_29879,N_29535);
xor UO_345 (O_345,N_29742,N_29598);
nand UO_346 (O_346,N_29839,N_29442);
nor UO_347 (O_347,N_29425,N_29614);
and UO_348 (O_348,N_29861,N_29817);
or UO_349 (O_349,N_29885,N_29421);
nand UO_350 (O_350,N_29926,N_29554);
xor UO_351 (O_351,N_29585,N_29869);
or UO_352 (O_352,N_29988,N_29620);
nand UO_353 (O_353,N_29865,N_29958);
xnor UO_354 (O_354,N_29887,N_29544);
and UO_355 (O_355,N_29563,N_29986);
or UO_356 (O_356,N_29777,N_29423);
xor UO_357 (O_357,N_29489,N_29658);
nor UO_358 (O_358,N_29798,N_29933);
nor UO_359 (O_359,N_29907,N_29696);
xor UO_360 (O_360,N_29439,N_29680);
or UO_361 (O_361,N_29450,N_29475);
nand UO_362 (O_362,N_29903,N_29817);
or UO_363 (O_363,N_29524,N_29633);
nor UO_364 (O_364,N_29523,N_29979);
and UO_365 (O_365,N_29801,N_29851);
and UO_366 (O_366,N_29894,N_29416);
and UO_367 (O_367,N_29684,N_29894);
xnor UO_368 (O_368,N_29649,N_29513);
xnor UO_369 (O_369,N_29967,N_29403);
xnor UO_370 (O_370,N_29551,N_29910);
xnor UO_371 (O_371,N_29420,N_29490);
or UO_372 (O_372,N_29814,N_29839);
nand UO_373 (O_373,N_29880,N_29745);
nand UO_374 (O_374,N_29425,N_29435);
nor UO_375 (O_375,N_29589,N_29855);
nand UO_376 (O_376,N_29917,N_29622);
or UO_377 (O_377,N_29409,N_29889);
or UO_378 (O_378,N_29515,N_29903);
xor UO_379 (O_379,N_29422,N_29541);
nor UO_380 (O_380,N_29434,N_29976);
and UO_381 (O_381,N_29663,N_29634);
xor UO_382 (O_382,N_29798,N_29793);
xnor UO_383 (O_383,N_29574,N_29547);
xnor UO_384 (O_384,N_29656,N_29491);
or UO_385 (O_385,N_29918,N_29961);
xor UO_386 (O_386,N_29666,N_29949);
nor UO_387 (O_387,N_29722,N_29978);
or UO_388 (O_388,N_29623,N_29578);
and UO_389 (O_389,N_29637,N_29783);
xor UO_390 (O_390,N_29856,N_29508);
and UO_391 (O_391,N_29488,N_29934);
xor UO_392 (O_392,N_29534,N_29838);
and UO_393 (O_393,N_29503,N_29584);
nand UO_394 (O_394,N_29698,N_29450);
or UO_395 (O_395,N_29837,N_29700);
nand UO_396 (O_396,N_29410,N_29595);
and UO_397 (O_397,N_29902,N_29933);
or UO_398 (O_398,N_29704,N_29762);
nor UO_399 (O_399,N_29804,N_29451);
or UO_400 (O_400,N_29989,N_29515);
xnor UO_401 (O_401,N_29839,N_29792);
and UO_402 (O_402,N_29618,N_29935);
nand UO_403 (O_403,N_29778,N_29861);
nand UO_404 (O_404,N_29755,N_29779);
nand UO_405 (O_405,N_29913,N_29725);
xnor UO_406 (O_406,N_29502,N_29514);
or UO_407 (O_407,N_29612,N_29708);
nor UO_408 (O_408,N_29542,N_29843);
xor UO_409 (O_409,N_29702,N_29726);
or UO_410 (O_410,N_29640,N_29451);
or UO_411 (O_411,N_29731,N_29876);
nand UO_412 (O_412,N_29718,N_29769);
and UO_413 (O_413,N_29418,N_29763);
nand UO_414 (O_414,N_29760,N_29480);
xor UO_415 (O_415,N_29696,N_29534);
or UO_416 (O_416,N_29536,N_29736);
or UO_417 (O_417,N_29620,N_29565);
nor UO_418 (O_418,N_29637,N_29787);
nor UO_419 (O_419,N_29464,N_29964);
or UO_420 (O_420,N_29467,N_29770);
or UO_421 (O_421,N_29538,N_29439);
nor UO_422 (O_422,N_29789,N_29637);
or UO_423 (O_423,N_29953,N_29683);
and UO_424 (O_424,N_29437,N_29519);
or UO_425 (O_425,N_29754,N_29487);
or UO_426 (O_426,N_29766,N_29727);
nand UO_427 (O_427,N_29874,N_29792);
nand UO_428 (O_428,N_29575,N_29971);
xnor UO_429 (O_429,N_29783,N_29459);
and UO_430 (O_430,N_29466,N_29438);
nor UO_431 (O_431,N_29616,N_29449);
and UO_432 (O_432,N_29804,N_29864);
xnor UO_433 (O_433,N_29961,N_29667);
and UO_434 (O_434,N_29509,N_29681);
or UO_435 (O_435,N_29475,N_29777);
nand UO_436 (O_436,N_29927,N_29805);
or UO_437 (O_437,N_29630,N_29499);
nor UO_438 (O_438,N_29420,N_29960);
nand UO_439 (O_439,N_29662,N_29413);
or UO_440 (O_440,N_29857,N_29782);
xor UO_441 (O_441,N_29442,N_29452);
xor UO_442 (O_442,N_29489,N_29609);
nand UO_443 (O_443,N_29992,N_29430);
nand UO_444 (O_444,N_29485,N_29418);
nand UO_445 (O_445,N_29618,N_29531);
xor UO_446 (O_446,N_29762,N_29421);
and UO_447 (O_447,N_29665,N_29689);
nor UO_448 (O_448,N_29983,N_29633);
nor UO_449 (O_449,N_29783,N_29941);
xor UO_450 (O_450,N_29763,N_29624);
and UO_451 (O_451,N_29564,N_29954);
nand UO_452 (O_452,N_29887,N_29669);
xnor UO_453 (O_453,N_29524,N_29963);
or UO_454 (O_454,N_29623,N_29883);
xnor UO_455 (O_455,N_29429,N_29501);
nor UO_456 (O_456,N_29439,N_29739);
nand UO_457 (O_457,N_29449,N_29898);
and UO_458 (O_458,N_29468,N_29960);
or UO_459 (O_459,N_29621,N_29823);
xnor UO_460 (O_460,N_29439,N_29411);
or UO_461 (O_461,N_29769,N_29597);
and UO_462 (O_462,N_29659,N_29966);
and UO_463 (O_463,N_29592,N_29570);
xnor UO_464 (O_464,N_29412,N_29849);
or UO_465 (O_465,N_29739,N_29454);
and UO_466 (O_466,N_29713,N_29941);
or UO_467 (O_467,N_29856,N_29614);
or UO_468 (O_468,N_29458,N_29845);
xor UO_469 (O_469,N_29592,N_29873);
nand UO_470 (O_470,N_29465,N_29593);
and UO_471 (O_471,N_29860,N_29937);
nand UO_472 (O_472,N_29687,N_29723);
and UO_473 (O_473,N_29768,N_29440);
and UO_474 (O_474,N_29616,N_29730);
and UO_475 (O_475,N_29813,N_29716);
and UO_476 (O_476,N_29594,N_29543);
xnor UO_477 (O_477,N_29487,N_29933);
or UO_478 (O_478,N_29979,N_29504);
or UO_479 (O_479,N_29696,N_29637);
nor UO_480 (O_480,N_29711,N_29466);
nand UO_481 (O_481,N_29938,N_29479);
xor UO_482 (O_482,N_29687,N_29951);
nor UO_483 (O_483,N_29528,N_29591);
nand UO_484 (O_484,N_29688,N_29533);
nor UO_485 (O_485,N_29568,N_29845);
or UO_486 (O_486,N_29580,N_29455);
nor UO_487 (O_487,N_29777,N_29716);
or UO_488 (O_488,N_29917,N_29539);
xnor UO_489 (O_489,N_29826,N_29945);
or UO_490 (O_490,N_29762,N_29807);
nor UO_491 (O_491,N_29497,N_29411);
xor UO_492 (O_492,N_29470,N_29832);
xor UO_493 (O_493,N_29420,N_29941);
xor UO_494 (O_494,N_29724,N_29660);
xnor UO_495 (O_495,N_29682,N_29897);
xnor UO_496 (O_496,N_29422,N_29402);
and UO_497 (O_497,N_29637,N_29680);
and UO_498 (O_498,N_29996,N_29965);
nand UO_499 (O_499,N_29547,N_29680);
and UO_500 (O_500,N_29963,N_29478);
and UO_501 (O_501,N_29467,N_29567);
xnor UO_502 (O_502,N_29984,N_29997);
nor UO_503 (O_503,N_29616,N_29750);
nand UO_504 (O_504,N_29975,N_29509);
xor UO_505 (O_505,N_29810,N_29685);
nor UO_506 (O_506,N_29783,N_29448);
and UO_507 (O_507,N_29763,N_29985);
xnor UO_508 (O_508,N_29826,N_29500);
nor UO_509 (O_509,N_29517,N_29918);
nor UO_510 (O_510,N_29956,N_29748);
or UO_511 (O_511,N_29906,N_29745);
nand UO_512 (O_512,N_29869,N_29512);
nand UO_513 (O_513,N_29426,N_29549);
xor UO_514 (O_514,N_29747,N_29599);
and UO_515 (O_515,N_29770,N_29673);
and UO_516 (O_516,N_29669,N_29451);
or UO_517 (O_517,N_29553,N_29556);
nor UO_518 (O_518,N_29895,N_29496);
nand UO_519 (O_519,N_29610,N_29662);
xor UO_520 (O_520,N_29905,N_29424);
and UO_521 (O_521,N_29471,N_29895);
or UO_522 (O_522,N_29870,N_29478);
nand UO_523 (O_523,N_29568,N_29605);
nand UO_524 (O_524,N_29432,N_29594);
nor UO_525 (O_525,N_29614,N_29812);
nand UO_526 (O_526,N_29706,N_29453);
nand UO_527 (O_527,N_29632,N_29615);
nand UO_528 (O_528,N_29728,N_29403);
xor UO_529 (O_529,N_29758,N_29636);
xnor UO_530 (O_530,N_29656,N_29450);
nor UO_531 (O_531,N_29978,N_29492);
nand UO_532 (O_532,N_29888,N_29869);
nor UO_533 (O_533,N_29839,N_29419);
and UO_534 (O_534,N_29973,N_29895);
or UO_535 (O_535,N_29882,N_29704);
or UO_536 (O_536,N_29831,N_29436);
xor UO_537 (O_537,N_29671,N_29706);
nand UO_538 (O_538,N_29611,N_29517);
xor UO_539 (O_539,N_29915,N_29706);
nand UO_540 (O_540,N_29853,N_29849);
nor UO_541 (O_541,N_29645,N_29648);
xnor UO_542 (O_542,N_29827,N_29502);
and UO_543 (O_543,N_29665,N_29466);
nor UO_544 (O_544,N_29513,N_29583);
nor UO_545 (O_545,N_29675,N_29679);
nand UO_546 (O_546,N_29575,N_29682);
and UO_547 (O_547,N_29706,N_29581);
nand UO_548 (O_548,N_29547,N_29461);
nor UO_549 (O_549,N_29906,N_29840);
nand UO_550 (O_550,N_29861,N_29953);
or UO_551 (O_551,N_29752,N_29860);
and UO_552 (O_552,N_29688,N_29982);
nor UO_553 (O_553,N_29450,N_29513);
nand UO_554 (O_554,N_29781,N_29907);
and UO_555 (O_555,N_29721,N_29635);
or UO_556 (O_556,N_29850,N_29770);
xor UO_557 (O_557,N_29484,N_29509);
nor UO_558 (O_558,N_29813,N_29937);
nand UO_559 (O_559,N_29614,N_29951);
or UO_560 (O_560,N_29568,N_29545);
or UO_561 (O_561,N_29745,N_29972);
nand UO_562 (O_562,N_29851,N_29857);
and UO_563 (O_563,N_29403,N_29566);
xor UO_564 (O_564,N_29834,N_29929);
nor UO_565 (O_565,N_29794,N_29943);
and UO_566 (O_566,N_29525,N_29983);
and UO_567 (O_567,N_29588,N_29975);
nand UO_568 (O_568,N_29722,N_29950);
or UO_569 (O_569,N_29582,N_29550);
nand UO_570 (O_570,N_29473,N_29886);
and UO_571 (O_571,N_29778,N_29577);
nor UO_572 (O_572,N_29725,N_29778);
nand UO_573 (O_573,N_29623,N_29781);
xnor UO_574 (O_574,N_29411,N_29485);
nand UO_575 (O_575,N_29660,N_29435);
nor UO_576 (O_576,N_29500,N_29897);
xnor UO_577 (O_577,N_29450,N_29740);
nand UO_578 (O_578,N_29854,N_29450);
and UO_579 (O_579,N_29926,N_29572);
nor UO_580 (O_580,N_29725,N_29474);
and UO_581 (O_581,N_29417,N_29623);
nand UO_582 (O_582,N_29552,N_29890);
nor UO_583 (O_583,N_29859,N_29445);
or UO_584 (O_584,N_29857,N_29827);
xor UO_585 (O_585,N_29452,N_29819);
xnor UO_586 (O_586,N_29507,N_29674);
and UO_587 (O_587,N_29536,N_29994);
nor UO_588 (O_588,N_29700,N_29499);
and UO_589 (O_589,N_29407,N_29605);
or UO_590 (O_590,N_29614,N_29611);
and UO_591 (O_591,N_29531,N_29868);
xnor UO_592 (O_592,N_29990,N_29512);
or UO_593 (O_593,N_29659,N_29738);
xor UO_594 (O_594,N_29759,N_29769);
or UO_595 (O_595,N_29960,N_29546);
and UO_596 (O_596,N_29442,N_29830);
or UO_597 (O_597,N_29810,N_29406);
or UO_598 (O_598,N_29820,N_29712);
or UO_599 (O_599,N_29597,N_29990);
nand UO_600 (O_600,N_29632,N_29813);
or UO_601 (O_601,N_29625,N_29692);
nand UO_602 (O_602,N_29732,N_29979);
nand UO_603 (O_603,N_29572,N_29576);
nor UO_604 (O_604,N_29532,N_29496);
xnor UO_605 (O_605,N_29655,N_29512);
and UO_606 (O_606,N_29489,N_29815);
xor UO_607 (O_607,N_29697,N_29665);
and UO_608 (O_608,N_29802,N_29799);
nand UO_609 (O_609,N_29603,N_29406);
or UO_610 (O_610,N_29864,N_29808);
nor UO_611 (O_611,N_29873,N_29641);
and UO_612 (O_612,N_29562,N_29924);
and UO_613 (O_613,N_29892,N_29638);
nor UO_614 (O_614,N_29898,N_29425);
nand UO_615 (O_615,N_29711,N_29710);
xnor UO_616 (O_616,N_29613,N_29630);
and UO_617 (O_617,N_29856,N_29808);
nand UO_618 (O_618,N_29727,N_29730);
or UO_619 (O_619,N_29524,N_29888);
and UO_620 (O_620,N_29981,N_29432);
and UO_621 (O_621,N_29546,N_29971);
xor UO_622 (O_622,N_29815,N_29931);
and UO_623 (O_623,N_29512,N_29550);
xor UO_624 (O_624,N_29584,N_29810);
nor UO_625 (O_625,N_29424,N_29810);
or UO_626 (O_626,N_29535,N_29485);
xor UO_627 (O_627,N_29950,N_29443);
and UO_628 (O_628,N_29412,N_29727);
nor UO_629 (O_629,N_29786,N_29692);
nand UO_630 (O_630,N_29514,N_29473);
nand UO_631 (O_631,N_29520,N_29613);
nor UO_632 (O_632,N_29945,N_29536);
and UO_633 (O_633,N_29631,N_29480);
and UO_634 (O_634,N_29628,N_29984);
nand UO_635 (O_635,N_29728,N_29820);
and UO_636 (O_636,N_29717,N_29826);
and UO_637 (O_637,N_29974,N_29983);
nor UO_638 (O_638,N_29710,N_29957);
nand UO_639 (O_639,N_29795,N_29440);
or UO_640 (O_640,N_29447,N_29733);
nand UO_641 (O_641,N_29501,N_29534);
nand UO_642 (O_642,N_29914,N_29517);
nor UO_643 (O_643,N_29934,N_29884);
and UO_644 (O_644,N_29481,N_29820);
nor UO_645 (O_645,N_29837,N_29610);
xnor UO_646 (O_646,N_29633,N_29577);
and UO_647 (O_647,N_29971,N_29914);
xnor UO_648 (O_648,N_29632,N_29629);
and UO_649 (O_649,N_29643,N_29813);
xnor UO_650 (O_650,N_29512,N_29820);
xnor UO_651 (O_651,N_29735,N_29494);
nand UO_652 (O_652,N_29715,N_29730);
xor UO_653 (O_653,N_29806,N_29752);
xnor UO_654 (O_654,N_29952,N_29749);
xor UO_655 (O_655,N_29878,N_29986);
xor UO_656 (O_656,N_29677,N_29568);
and UO_657 (O_657,N_29423,N_29490);
nand UO_658 (O_658,N_29461,N_29912);
or UO_659 (O_659,N_29939,N_29578);
nand UO_660 (O_660,N_29652,N_29989);
and UO_661 (O_661,N_29882,N_29469);
and UO_662 (O_662,N_29922,N_29663);
nand UO_663 (O_663,N_29458,N_29908);
nor UO_664 (O_664,N_29981,N_29405);
and UO_665 (O_665,N_29739,N_29538);
nor UO_666 (O_666,N_29818,N_29966);
nor UO_667 (O_667,N_29804,N_29437);
and UO_668 (O_668,N_29633,N_29821);
nand UO_669 (O_669,N_29403,N_29955);
or UO_670 (O_670,N_29817,N_29694);
xor UO_671 (O_671,N_29709,N_29828);
or UO_672 (O_672,N_29827,N_29978);
nand UO_673 (O_673,N_29835,N_29627);
nor UO_674 (O_674,N_29460,N_29967);
or UO_675 (O_675,N_29804,N_29537);
xnor UO_676 (O_676,N_29430,N_29860);
nor UO_677 (O_677,N_29819,N_29433);
nand UO_678 (O_678,N_29978,N_29521);
and UO_679 (O_679,N_29410,N_29809);
xor UO_680 (O_680,N_29967,N_29542);
or UO_681 (O_681,N_29996,N_29719);
or UO_682 (O_682,N_29992,N_29702);
and UO_683 (O_683,N_29504,N_29872);
nor UO_684 (O_684,N_29780,N_29665);
nand UO_685 (O_685,N_29877,N_29924);
or UO_686 (O_686,N_29858,N_29827);
or UO_687 (O_687,N_29713,N_29711);
and UO_688 (O_688,N_29651,N_29930);
nor UO_689 (O_689,N_29855,N_29566);
or UO_690 (O_690,N_29841,N_29443);
and UO_691 (O_691,N_29526,N_29702);
and UO_692 (O_692,N_29721,N_29440);
nor UO_693 (O_693,N_29772,N_29415);
xor UO_694 (O_694,N_29421,N_29977);
or UO_695 (O_695,N_29458,N_29686);
xor UO_696 (O_696,N_29688,N_29689);
nor UO_697 (O_697,N_29758,N_29544);
nand UO_698 (O_698,N_29675,N_29520);
xnor UO_699 (O_699,N_29477,N_29797);
nor UO_700 (O_700,N_29450,N_29744);
nand UO_701 (O_701,N_29818,N_29495);
xor UO_702 (O_702,N_29778,N_29818);
and UO_703 (O_703,N_29972,N_29943);
or UO_704 (O_704,N_29943,N_29873);
xnor UO_705 (O_705,N_29566,N_29741);
nor UO_706 (O_706,N_29589,N_29660);
xor UO_707 (O_707,N_29637,N_29874);
xnor UO_708 (O_708,N_29529,N_29508);
and UO_709 (O_709,N_29666,N_29821);
and UO_710 (O_710,N_29909,N_29408);
xnor UO_711 (O_711,N_29646,N_29498);
nand UO_712 (O_712,N_29852,N_29565);
xor UO_713 (O_713,N_29892,N_29767);
and UO_714 (O_714,N_29526,N_29831);
nor UO_715 (O_715,N_29945,N_29481);
and UO_716 (O_716,N_29543,N_29492);
nor UO_717 (O_717,N_29988,N_29916);
nor UO_718 (O_718,N_29990,N_29409);
nand UO_719 (O_719,N_29925,N_29455);
xnor UO_720 (O_720,N_29739,N_29587);
nor UO_721 (O_721,N_29616,N_29825);
nand UO_722 (O_722,N_29428,N_29752);
or UO_723 (O_723,N_29990,N_29900);
xnor UO_724 (O_724,N_29607,N_29709);
nand UO_725 (O_725,N_29437,N_29444);
and UO_726 (O_726,N_29505,N_29829);
xor UO_727 (O_727,N_29842,N_29895);
and UO_728 (O_728,N_29913,N_29836);
and UO_729 (O_729,N_29703,N_29522);
or UO_730 (O_730,N_29480,N_29511);
nor UO_731 (O_731,N_29608,N_29913);
xor UO_732 (O_732,N_29920,N_29690);
nand UO_733 (O_733,N_29444,N_29591);
or UO_734 (O_734,N_29755,N_29862);
xnor UO_735 (O_735,N_29885,N_29588);
or UO_736 (O_736,N_29928,N_29755);
and UO_737 (O_737,N_29589,N_29938);
or UO_738 (O_738,N_29481,N_29735);
nor UO_739 (O_739,N_29468,N_29437);
xnor UO_740 (O_740,N_29543,N_29653);
or UO_741 (O_741,N_29980,N_29869);
or UO_742 (O_742,N_29583,N_29829);
nor UO_743 (O_743,N_29611,N_29573);
nand UO_744 (O_744,N_29574,N_29524);
nor UO_745 (O_745,N_29787,N_29842);
nand UO_746 (O_746,N_29493,N_29404);
nor UO_747 (O_747,N_29844,N_29833);
and UO_748 (O_748,N_29459,N_29557);
nand UO_749 (O_749,N_29620,N_29615);
and UO_750 (O_750,N_29618,N_29573);
nand UO_751 (O_751,N_29807,N_29715);
or UO_752 (O_752,N_29732,N_29677);
xnor UO_753 (O_753,N_29479,N_29400);
nand UO_754 (O_754,N_29462,N_29483);
nand UO_755 (O_755,N_29906,N_29923);
nand UO_756 (O_756,N_29829,N_29581);
and UO_757 (O_757,N_29693,N_29962);
nor UO_758 (O_758,N_29536,N_29716);
and UO_759 (O_759,N_29628,N_29598);
or UO_760 (O_760,N_29989,N_29481);
xnor UO_761 (O_761,N_29700,N_29933);
and UO_762 (O_762,N_29995,N_29767);
nand UO_763 (O_763,N_29646,N_29792);
nand UO_764 (O_764,N_29475,N_29454);
nand UO_765 (O_765,N_29572,N_29796);
nor UO_766 (O_766,N_29581,N_29935);
nand UO_767 (O_767,N_29865,N_29669);
and UO_768 (O_768,N_29890,N_29617);
nand UO_769 (O_769,N_29785,N_29689);
xnor UO_770 (O_770,N_29863,N_29683);
or UO_771 (O_771,N_29566,N_29770);
nor UO_772 (O_772,N_29408,N_29956);
or UO_773 (O_773,N_29572,N_29758);
nor UO_774 (O_774,N_29581,N_29995);
nor UO_775 (O_775,N_29739,N_29475);
and UO_776 (O_776,N_29832,N_29778);
or UO_777 (O_777,N_29724,N_29863);
or UO_778 (O_778,N_29795,N_29993);
or UO_779 (O_779,N_29459,N_29733);
and UO_780 (O_780,N_29678,N_29443);
xor UO_781 (O_781,N_29444,N_29415);
or UO_782 (O_782,N_29432,N_29915);
xor UO_783 (O_783,N_29695,N_29740);
or UO_784 (O_784,N_29685,N_29727);
nand UO_785 (O_785,N_29910,N_29843);
nor UO_786 (O_786,N_29714,N_29420);
and UO_787 (O_787,N_29730,N_29612);
and UO_788 (O_788,N_29665,N_29761);
nor UO_789 (O_789,N_29688,N_29930);
xor UO_790 (O_790,N_29857,N_29907);
nand UO_791 (O_791,N_29726,N_29882);
and UO_792 (O_792,N_29905,N_29608);
nand UO_793 (O_793,N_29796,N_29982);
xor UO_794 (O_794,N_29815,N_29424);
or UO_795 (O_795,N_29913,N_29638);
or UO_796 (O_796,N_29844,N_29715);
nand UO_797 (O_797,N_29723,N_29447);
xnor UO_798 (O_798,N_29960,N_29455);
and UO_799 (O_799,N_29668,N_29815);
nor UO_800 (O_800,N_29481,N_29886);
xor UO_801 (O_801,N_29731,N_29661);
or UO_802 (O_802,N_29651,N_29457);
nor UO_803 (O_803,N_29978,N_29657);
nand UO_804 (O_804,N_29911,N_29451);
nand UO_805 (O_805,N_29427,N_29856);
nor UO_806 (O_806,N_29451,N_29887);
and UO_807 (O_807,N_29436,N_29583);
nand UO_808 (O_808,N_29928,N_29724);
and UO_809 (O_809,N_29683,N_29733);
nor UO_810 (O_810,N_29624,N_29815);
nand UO_811 (O_811,N_29880,N_29776);
or UO_812 (O_812,N_29978,N_29465);
nand UO_813 (O_813,N_29700,N_29838);
or UO_814 (O_814,N_29766,N_29527);
nand UO_815 (O_815,N_29927,N_29746);
and UO_816 (O_816,N_29762,N_29767);
nor UO_817 (O_817,N_29859,N_29410);
and UO_818 (O_818,N_29991,N_29848);
and UO_819 (O_819,N_29474,N_29759);
or UO_820 (O_820,N_29936,N_29433);
or UO_821 (O_821,N_29971,N_29488);
nor UO_822 (O_822,N_29893,N_29809);
or UO_823 (O_823,N_29482,N_29856);
nor UO_824 (O_824,N_29989,N_29696);
or UO_825 (O_825,N_29463,N_29627);
nand UO_826 (O_826,N_29741,N_29773);
or UO_827 (O_827,N_29436,N_29969);
nand UO_828 (O_828,N_29830,N_29884);
nor UO_829 (O_829,N_29793,N_29509);
nor UO_830 (O_830,N_29800,N_29420);
nand UO_831 (O_831,N_29683,N_29588);
nor UO_832 (O_832,N_29962,N_29967);
or UO_833 (O_833,N_29681,N_29752);
xor UO_834 (O_834,N_29882,N_29841);
and UO_835 (O_835,N_29980,N_29696);
and UO_836 (O_836,N_29516,N_29691);
nor UO_837 (O_837,N_29760,N_29947);
and UO_838 (O_838,N_29476,N_29668);
and UO_839 (O_839,N_29679,N_29465);
xnor UO_840 (O_840,N_29911,N_29879);
xor UO_841 (O_841,N_29899,N_29878);
nor UO_842 (O_842,N_29451,N_29664);
xnor UO_843 (O_843,N_29971,N_29789);
xnor UO_844 (O_844,N_29768,N_29686);
and UO_845 (O_845,N_29457,N_29755);
nor UO_846 (O_846,N_29932,N_29749);
and UO_847 (O_847,N_29448,N_29577);
xnor UO_848 (O_848,N_29547,N_29666);
or UO_849 (O_849,N_29823,N_29609);
nand UO_850 (O_850,N_29941,N_29558);
or UO_851 (O_851,N_29916,N_29526);
nor UO_852 (O_852,N_29948,N_29801);
xnor UO_853 (O_853,N_29989,N_29764);
nand UO_854 (O_854,N_29675,N_29871);
and UO_855 (O_855,N_29768,N_29789);
and UO_856 (O_856,N_29623,N_29407);
xnor UO_857 (O_857,N_29673,N_29413);
nor UO_858 (O_858,N_29495,N_29556);
or UO_859 (O_859,N_29556,N_29419);
nand UO_860 (O_860,N_29722,N_29456);
nor UO_861 (O_861,N_29714,N_29973);
xnor UO_862 (O_862,N_29581,N_29824);
or UO_863 (O_863,N_29961,N_29627);
and UO_864 (O_864,N_29625,N_29906);
nand UO_865 (O_865,N_29503,N_29952);
or UO_866 (O_866,N_29754,N_29943);
or UO_867 (O_867,N_29787,N_29453);
and UO_868 (O_868,N_29511,N_29535);
or UO_869 (O_869,N_29963,N_29730);
nor UO_870 (O_870,N_29871,N_29818);
nand UO_871 (O_871,N_29956,N_29526);
nand UO_872 (O_872,N_29940,N_29569);
and UO_873 (O_873,N_29640,N_29595);
xnor UO_874 (O_874,N_29499,N_29447);
nand UO_875 (O_875,N_29493,N_29762);
nand UO_876 (O_876,N_29710,N_29426);
nor UO_877 (O_877,N_29874,N_29400);
xnor UO_878 (O_878,N_29643,N_29846);
nand UO_879 (O_879,N_29695,N_29960);
xnor UO_880 (O_880,N_29938,N_29524);
and UO_881 (O_881,N_29736,N_29963);
and UO_882 (O_882,N_29942,N_29419);
xor UO_883 (O_883,N_29979,N_29759);
xor UO_884 (O_884,N_29443,N_29493);
or UO_885 (O_885,N_29526,N_29586);
or UO_886 (O_886,N_29626,N_29537);
xor UO_887 (O_887,N_29708,N_29945);
nand UO_888 (O_888,N_29492,N_29461);
xor UO_889 (O_889,N_29972,N_29653);
and UO_890 (O_890,N_29629,N_29771);
nand UO_891 (O_891,N_29565,N_29893);
nand UO_892 (O_892,N_29782,N_29574);
or UO_893 (O_893,N_29546,N_29769);
nor UO_894 (O_894,N_29684,N_29725);
or UO_895 (O_895,N_29741,N_29461);
nor UO_896 (O_896,N_29462,N_29746);
or UO_897 (O_897,N_29744,N_29801);
nor UO_898 (O_898,N_29498,N_29452);
or UO_899 (O_899,N_29905,N_29670);
nor UO_900 (O_900,N_29703,N_29659);
nor UO_901 (O_901,N_29962,N_29753);
and UO_902 (O_902,N_29437,N_29916);
and UO_903 (O_903,N_29540,N_29921);
xor UO_904 (O_904,N_29759,N_29414);
nand UO_905 (O_905,N_29718,N_29961);
xor UO_906 (O_906,N_29632,N_29691);
nand UO_907 (O_907,N_29583,N_29924);
nand UO_908 (O_908,N_29864,N_29718);
and UO_909 (O_909,N_29810,N_29963);
nand UO_910 (O_910,N_29562,N_29644);
and UO_911 (O_911,N_29829,N_29677);
xnor UO_912 (O_912,N_29614,N_29786);
nand UO_913 (O_913,N_29897,N_29908);
and UO_914 (O_914,N_29835,N_29514);
nand UO_915 (O_915,N_29724,N_29794);
and UO_916 (O_916,N_29416,N_29749);
nand UO_917 (O_917,N_29826,N_29834);
nor UO_918 (O_918,N_29655,N_29971);
nor UO_919 (O_919,N_29554,N_29863);
nand UO_920 (O_920,N_29539,N_29756);
nand UO_921 (O_921,N_29701,N_29650);
nor UO_922 (O_922,N_29727,N_29425);
and UO_923 (O_923,N_29645,N_29939);
and UO_924 (O_924,N_29928,N_29925);
nand UO_925 (O_925,N_29427,N_29921);
nor UO_926 (O_926,N_29755,N_29692);
nor UO_927 (O_927,N_29684,N_29939);
nor UO_928 (O_928,N_29528,N_29456);
and UO_929 (O_929,N_29880,N_29661);
nor UO_930 (O_930,N_29531,N_29505);
nand UO_931 (O_931,N_29914,N_29524);
xnor UO_932 (O_932,N_29812,N_29811);
nor UO_933 (O_933,N_29495,N_29856);
nand UO_934 (O_934,N_29475,N_29714);
or UO_935 (O_935,N_29780,N_29890);
or UO_936 (O_936,N_29509,N_29508);
nand UO_937 (O_937,N_29444,N_29723);
and UO_938 (O_938,N_29659,N_29569);
and UO_939 (O_939,N_29841,N_29713);
xnor UO_940 (O_940,N_29784,N_29826);
nor UO_941 (O_941,N_29439,N_29531);
xor UO_942 (O_942,N_29678,N_29840);
or UO_943 (O_943,N_29793,N_29791);
and UO_944 (O_944,N_29715,N_29734);
or UO_945 (O_945,N_29571,N_29485);
nand UO_946 (O_946,N_29642,N_29610);
or UO_947 (O_947,N_29466,N_29849);
or UO_948 (O_948,N_29824,N_29734);
nor UO_949 (O_949,N_29989,N_29889);
xor UO_950 (O_950,N_29941,N_29416);
and UO_951 (O_951,N_29879,N_29729);
nor UO_952 (O_952,N_29997,N_29623);
or UO_953 (O_953,N_29735,N_29662);
nor UO_954 (O_954,N_29687,N_29969);
or UO_955 (O_955,N_29931,N_29537);
and UO_956 (O_956,N_29823,N_29822);
and UO_957 (O_957,N_29932,N_29526);
xor UO_958 (O_958,N_29768,N_29542);
nor UO_959 (O_959,N_29883,N_29411);
and UO_960 (O_960,N_29943,N_29426);
or UO_961 (O_961,N_29972,N_29555);
and UO_962 (O_962,N_29787,N_29960);
nor UO_963 (O_963,N_29656,N_29617);
nand UO_964 (O_964,N_29931,N_29875);
and UO_965 (O_965,N_29878,N_29668);
xor UO_966 (O_966,N_29745,N_29840);
nand UO_967 (O_967,N_29674,N_29710);
or UO_968 (O_968,N_29540,N_29459);
nor UO_969 (O_969,N_29988,N_29502);
and UO_970 (O_970,N_29779,N_29528);
nor UO_971 (O_971,N_29415,N_29587);
nand UO_972 (O_972,N_29417,N_29627);
or UO_973 (O_973,N_29638,N_29663);
xor UO_974 (O_974,N_29899,N_29770);
xor UO_975 (O_975,N_29656,N_29565);
nor UO_976 (O_976,N_29850,N_29861);
or UO_977 (O_977,N_29864,N_29881);
or UO_978 (O_978,N_29596,N_29825);
nand UO_979 (O_979,N_29716,N_29670);
xnor UO_980 (O_980,N_29829,N_29885);
nand UO_981 (O_981,N_29863,N_29416);
nor UO_982 (O_982,N_29571,N_29808);
xor UO_983 (O_983,N_29406,N_29510);
nor UO_984 (O_984,N_29756,N_29531);
and UO_985 (O_985,N_29651,N_29437);
xnor UO_986 (O_986,N_29493,N_29693);
nor UO_987 (O_987,N_29845,N_29906);
xor UO_988 (O_988,N_29926,N_29809);
or UO_989 (O_989,N_29415,N_29837);
xor UO_990 (O_990,N_29829,N_29465);
and UO_991 (O_991,N_29592,N_29576);
nor UO_992 (O_992,N_29697,N_29746);
or UO_993 (O_993,N_29435,N_29875);
nor UO_994 (O_994,N_29408,N_29897);
and UO_995 (O_995,N_29654,N_29748);
or UO_996 (O_996,N_29568,N_29729);
xor UO_997 (O_997,N_29657,N_29412);
xor UO_998 (O_998,N_29446,N_29685);
nor UO_999 (O_999,N_29862,N_29635);
xnor UO_1000 (O_1000,N_29851,N_29831);
nand UO_1001 (O_1001,N_29727,N_29879);
and UO_1002 (O_1002,N_29766,N_29535);
nor UO_1003 (O_1003,N_29481,N_29969);
or UO_1004 (O_1004,N_29856,N_29577);
nand UO_1005 (O_1005,N_29524,N_29498);
nand UO_1006 (O_1006,N_29732,N_29999);
nor UO_1007 (O_1007,N_29658,N_29559);
or UO_1008 (O_1008,N_29411,N_29647);
xnor UO_1009 (O_1009,N_29924,N_29437);
xnor UO_1010 (O_1010,N_29959,N_29796);
and UO_1011 (O_1011,N_29428,N_29941);
or UO_1012 (O_1012,N_29576,N_29907);
xnor UO_1013 (O_1013,N_29644,N_29629);
and UO_1014 (O_1014,N_29584,N_29695);
xnor UO_1015 (O_1015,N_29415,N_29416);
xor UO_1016 (O_1016,N_29595,N_29409);
or UO_1017 (O_1017,N_29511,N_29411);
and UO_1018 (O_1018,N_29495,N_29489);
and UO_1019 (O_1019,N_29698,N_29895);
and UO_1020 (O_1020,N_29753,N_29569);
and UO_1021 (O_1021,N_29991,N_29675);
nand UO_1022 (O_1022,N_29623,N_29918);
or UO_1023 (O_1023,N_29845,N_29841);
and UO_1024 (O_1024,N_29991,N_29896);
nand UO_1025 (O_1025,N_29609,N_29416);
or UO_1026 (O_1026,N_29976,N_29523);
or UO_1027 (O_1027,N_29661,N_29780);
xor UO_1028 (O_1028,N_29995,N_29673);
xor UO_1029 (O_1029,N_29795,N_29705);
or UO_1030 (O_1030,N_29542,N_29518);
nor UO_1031 (O_1031,N_29457,N_29976);
and UO_1032 (O_1032,N_29641,N_29911);
xor UO_1033 (O_1033,N_29570,N_29772);
xor UO_1034 (O_1034,N_29591,N_29923);
xnor UO_1035 (O_1035,N_29767,N_29666);
xor UO_1036 (O_1036,N_29897,N_29430);
and UO_1037 (O_1037,N_29973,N_29874);
nor UO_1038 (O_1038,N_29656,N_29483);
xnor UO_1039 (O_1039,N_29632,N_29756);
nor UO_1040 (O_1040,N_29607,N_29706);
and UO_1041 (O_1041,N_29953,N_29919);
or UO_1042 (O_1042,N_29574,N_29495);
xnor UO_1043 (O_1043,N_29489,N_29756);
xor UO_1044 (O_1044,N_29819,N_29794);
nand UO_1045 (O_1045,N_29734,N_29678);
or UO_1046 (O_1046,N_29793,N_29865);
nor UO_1047 (O_1047,N_29873,N_29655);
nand UO_1048 (O_1048,N_29659,N_29692);
and UO_1049 (O_1049,N_29529,N_29604);
nor UO_1050 (O_1050,N_29943,N_29771);
nand UO_1051 (O_1051,N_29971,N_29818);
nand UO_1052 (O_1052,N_29595,N_29861);
and UO_1053 (O_1053,N_29733,N_29693);
xor UO_1054 (O_1054,N_29707,N_29625);
nor UO_1055 (O_1055,N_29879,N_29623);
and UO_1056 (O_1056,N_29894,N_29676);
or UO_1057 (O_1057,N_29888,N_29473);
or UO_1058 (O_1058,N_29484,N_29469);
nor UO_1059 (O_1059,N_29501,N_29747);
nor UO_1060 (O_1060,N_29796,N_29437);
nor UO_1061 (O_1061,N_29973,N_29949);
nor UO_1062 (O_1062,N_29827,N_29657);
or UO_1063 (O_1063,N_29572,N_29763);
or UO_1064 (O_1064,N_29438,N_29591);
and UO_1065 (O_1065,N_29785,N_29495);
nand UO_1066 (O_1066,N_29753,N_29592);
or UO_1067 (O_1067,N_29879,N_29964);
nand UO_1068 (O_1068,N_29761,N_29856);
xor UO_1069 (O_1069,N_29942,N_29534);
nor UO_1070 (O_1070,N_29873,N_29811);
nand UO_1071 (O_1071,N_29534,N_29768);
and UO_1072 (O_1072,N_29776,N_29600);
and UO_1073 (O_1073,N_29795,N_29966);
or UO_1074 (O_1074,N_29446,N_29552);
xor UO_1075 (O_1075,N_29992,N_29497);
nand UO_1076 (O_1076,N_29957,N_29410);
or UO_1077 (O_1077,N_29601,N_29650);
nor UO_1078 (O_1078,N_29403,N_29795);
or UO_1079 (O_1079,N_29898,N_29418);
and UO_1080 (O_1080,N_29481,N_29526);
and UO_1081 (O_1081,N_29576,N_29904);
nor UO_1082 (O_1082,N_29987,N_29756);
nand UO_1083 (O_1083,N_29700,N_29936);
xor UO_1084 (O_1084,N_29905,N_29654);
and UO_1085 (O_1085,N_29483,N_29748);
xor UO_1086 (O_1086,N_29922,N_29606);
nor UO_1087 (O_1087,N_29927,N_29481);
nor UO_1088 (O_1088,N_29876,N_29920);
and UO_1089 (O_1089,N_29954,N_29840);
and UO_1090 (O_1090,N_29401,N_29561);
or UO_1091 (O_1091,N_29484,N_29504);
or UO_1092 (O_1092,N_29538,N_29661);
nor UO_1093 (O_1093,N_29926,N_29844);
xor UO_1094 (O_1094,N_29995,N_29572);
or UO_1095 (O_1095,N_29743,N_29778);
xnor UO_1096 (O_1096,N_29996,N_29915);
or UO_1097 (O_1097,N_29781,N_29590);
nand UO_1098 (O_1098,N_29401,N_29498);
and UO_1099 (O_1099,N_29406,N_29633);
nor UO_1100 (O_1100,N_29547,N_29811);
nor UO_1101 (O_1101,N_29950,N_29840);
and UO_1102 (O_1102,N_29603,N_29851);
nand UO_1103 (O_1103,N_29865,N_29508);
and UO_1104 (O_1104,N_29479,N_29893);
nand UO_1105 (O_1105,N_29956,N_29862);
and UO_1106 (O_1106,N_29790,N_29567);
xnor UO_1107 (O_1107,N_29891,N_29634);
xor UO_1108 (O_1108,N_29874,N_29678);
nor UO_1109 (O_1109,N_29431,N_29501);
nand UO_1110 (O_1110,N_29913,N_29578);
nand UO_1111 (O_1111,N_29577,N_29800);
xor UO_1112 (O_1112,N_29453,N_29464);
nor UO_1113 (O_1113,N_29426,N_29997);
and UO_1114 (O_1114,N_29744,N_29722);
xor UO_1115 (O_1115,N_29897,N_29855);
xor UO_1116 (O_1116,N_29760,N_29624);
nand UO_1117 (O_1117,N_29888,N_29486);
xor UO_1118 (O_1118,N_29412,N_29589);
xnor UO_1119 (O_1119,N_29894,N_29801);
xnor UO_1120 (O_1120,N_29667,N_29935);
or UO_1121 (O_1121,N_29473,N_29457);
nand UO_1122 (O_1122,N_29957,N_29842);
nor UO_1123 (O_1123,N_29982,N_29761);
nor UO_1124 (O_1124,N_29415,N_29540);
nand UO_1125 (O_1125,N_29684,N_29417);
xor UO_1126 (O_1126,N_29428,N_29632);
and UO_1127 (O_1127,N_29583,N_29490);
and UO_1128 (O_1128,N_29509,N_29925);
and UO_1129 (O_1129,N_29626,N_29937);
nand UO_1130 (O_1130,N_29585,N_29767);
and UO_1131 (O_1131,N_29406,N_29681);
nand UO_1132 (O_1132,N_29414,N_29904);
xor UO_1133 (O_1133,N_29558,N_29501);
xnor UO_1134 (O_1134,N_29642,N_29720);
and UO_1135 (O_1135,N_29687,N_29662);
nand UO_1136 (O_1136,N_29772,N_29649);
nand UO_1137 (O_1137,N_29985,N_29498);
nor UO_1138 (O_1138,N_29458,N_29421);
or UO_1139 (O_1139,N_29664,N_29892);
xnor UO_1140 (O_1140,N_29810,N_29949);
nand UO_1141 (O_1141,N_29914,N_29584);
nor UO_1142 (O_1142,N_29941,N_29846);
or UO_1143 (O_1143,N_29618,N_29919);
or UO_1144 (O_1144,N_29465,N_29442);
nor UO_1145 (O_1145,N_29889,N_29947);
nor UO_1146 (O_1146,N_29776,N_29720);
and UO_1147 (O_1147,N_29755,N_29541);
nor UO_1148 (O_1148,N_29587,N_29900);
or UO_1149 (O_1149,N_29789,N_29691);
xnor UO_1150 (O_1150,N_29727,N_29837);
nand UO_1151 (O_1151,N_29834,N_29883);
xnor UO_1152 (O_1152,N_29754,N_29517);
xnor UO_1153 (O_1153,N_29702,N_29935);
xor UO_1154 (O_1154,N_29403,N_29976);
xnor UO_1155 (O_1155,N_29556,N_29987);
nor UO_1156 (O_1156,N_29958,N_29472);
nor UO_1157 (O_1157,N_29993,N_29955);
nand UO_1158 (O_1158,N_29579,N_29680);
or UO_1159 (O_1159,N_29518,N_29475);
xor UO_1160 (O_1160,N_29463,N_29684);
and UO_1161 (O_1161,N_29619,N_29735);
xor UO_1162 (O_1162,N_29484,N_29689);
or UO_1163 (O_1163,N_29525,N_29450);
or UO_1164 (O_1164,N_29666,N_29447);
xor UO_1165 (O_1165,N_29682,N_29612);
nand UO_1166 (O_1166,N_29494,N_29499);
nand UO_1167 (O_1167,N_29533,N_29924);
and UO_1168 (O_1168,N_29866,N_29953);
nand UO_1169 (O_1169,N_29665,N_29601);
nand UO_1170 (O_1170,N_29563,N_29833);
nor UO_1171 (O_1171,N_29828,N_29651);
or UO_1172 (O_1172,N_29517,N_29547);
nor UO_1173 (O_1173,N_29407,N_29488);
nor UO_1174 (O_1174,N_29634,N_29866);
and UO_1175 (O_1175,N_29611,N_29955);
or UO_1176 (O_1176,N_29634,N_29623);
or UO_1177 (O_1177,N_29880,N_29738);
nor UO_1178 (O_1178,N_29731,N_29943);
nand UO_1179 (O_1179,N_29579,N_29911);
xor UO_1180 (O_1180,N_29824,N_29798);
or UO_1181 (O_1181,N_29547,N_29495);
or UO_1182 (O_1182,N_29968,N_29531);
or UO_1183 (O_1183,N_29957,N_29474);
xor UO_1184 (O_1184,N_29957,N_29559);
or UO_1185 (O_1185,N_29414,N_29446);
and UO_1186 (O_1186,N_29977,N_29550);
nand UO_1187 (O_1187,N_29886,N_29457);
and UO_1188 (O_1188,N_29970,N_29943);
or UO_1189 (O_1189,N_29492,N_29418);
and UO_1190 (O_1190,N_29696,N_29853);
nor UO_1191 (O_1191,N_29788,N_29470);
nor UO_1192 (O_1192,N_29452,N_29449);
and UO_1193 (O_1193,N_29906,N_29973);
nand UO_1194 (O_1194,N_29737,N_29765);
xnor UO_1195 (O_1195,N_29787,N_29725);
xor UO_1196 (O_1196,N_29836,N_29984);
nor UO_1197 (O_1197,N_29421,N_29523);
or UO_1198 (O_1198,N_29590,N_29567);
nand UO_1199 (O_1199,N_29904,N_29430);
and UO_1200 (O_1200,N_29764,N_29571);
or UO_1201 (O_1201,N_29793,N_29970);
nor UO_1202 (O_1202,N_29875,N_29984);
or UO_1203 (O_1203,N_29438,N_29624);
nand UO_1204 (O_1204,N_29479,N_29931);
nor UO_1205 (O_1205,N_29697,N_29568);
xnor UO_1206 (O_1206,N_29671,N_29941);
nor UO_1207 (O_1207,N_29474,N_29662);
xor UO_1208 (O_1208,N_29874,N_29859);
xor UO_1209 (O_1209,N_29604,N_29924);
and UO_1210 (O_1210,N_29500,N_29699);
nand UO_1211 (O_1211,N_29622,N_29722);
nor UO_1212 (O_1212,N_29768,N_29443);
and UO_1213 (O_1213,N_29666,N_29872);
nor UO_1214 (O_1214,N_29767,N_29769);
or UO_1215 (O_1215,N_29566,N_29881);
nor UO_1216 (O_1216,N_29740,N_29867);
and UO_1217 (O_1217,N_29431,N_29920);
and UO_1218 (O_1218,N_29913,N_29639);
and UO_1219 (O_1219,N_29614,N_29893);
or UO_1220 (O_1220,N_29997,N_29440);
nor UO_1221 (O_1221,N_29591,N_29650);
and UO_1222 (O_1222,N_29425,N_29441);
or UO_1223 (O_1223,N_29406,N_29621);
and UO_1224 (O_1224,N_29414,N_29611);
nand UO_1225 (O_1225,N_29459,N_29695);
nand UO_1226 (O_1226,N_29973,N_29823);
and UO_1227 (O_1227,N_29645,N_29938);
nor UO_1228 (O_1228,N_29428,N_29931);
and UO_1229 (O_1229,N_29955,N_29688);
nand UO_1230 (O_1230,N_29491,N_29689);
and UO_1231 (O_1231,N_29995,N_29672);
nand UO_1232 (O_1232,N_29800,N_29794);
and UO_1233 (O_1233,N_29850,N_29634);
nor UO_1234 (O_1234,N_29846,N_29981);
and UO_1235 (O_1235,N_29623,N_29715);
and UO_1236 (O_1236,N_29945,N_29745);
xnor UO_1237 (O_1237,N_29607,N_29759);
nor UO_1238 (O_1238,N_29547,N_29499);
or UO_1239 (O_1239,N_29618,N_29647);
and UO_1240 (O_1240,N_29537,N_29798);
nor UO_1241 (O_1241,N_29662,N_29454);
nand UO_1242 (O_1242,N_29953,N_29559);
nor UO_1243 (O_1243,N_29551,N_29548);
and UO_1244 (O_1244,N_29623,N_29905);
nor UO_1245 (O_1245,N_29719,N_29473);
nor UO_1246 (O_1246,N_29864,N_29542);
nand UO_1247 (O_1247,N_29435,N_29800);
nor UO_1248 (O_1248,N_29829,N_29835);
and UO_1249 (O_1249,N_29655,N_29659);
or UO_1250 (O_1250,N_29687,N_29633);
nand UO_1251 (O_1251,N_29889,N_29707);
or UO_1252 (O_1252,N_29490,N_29520);
and UO_1253 (O_1253,N_29895,N_29759);
nand UO_1254 (O_1254,N_29513,N_29880);
nand UO_1255 (O_1255,N_29447,N_29434);
nor UO_1256 (O_1256,N_29833,N_29716);
xnor UO_1257 (O_1257,N_29463,N_29732);
nand UO_1258 (O_1258,N_29574,N_29991);
and UO_1259 (O_1259,N_29904,N_29949);
and UO_1260 (O_1260,N_29930,N_29724);
nor UO_1261 (O_1261,N_29432,N_29551);
nor UO_1262 (O_1262,N_29596,N_29747);
or UO_1263 (O_1263,N_29444,N_29760);
nand UO_1264 (O_1264,N_29493,N_29900);
nand UO_1265 (O_1265,N_29428,N_29997);
and UO_1266 (O_1266,N_29420,N_29712);
nand UO_1267 (O_1267,N_29822,N_29980);
nand UO_1268 (O_1268,N_29817,N_29603);
and UO_1269 (O_1269,N_29463,N_29768);
and UO_1270 (O_1270,N_29407,N_29821);
nor UO_1271 (O_1271,N_29563,N_29521);
nand UO_1272 (O_1272,N_29676,N_29948);
xnor UO_1273 (O_1273,N_29558,N_29807);
nand UO_1274 (O_1274,N_29735,N_29487);
and UO_1275 (O_1275,N_29824,N_29875);
xor UO_1276 (O_1276,N_29813,N_29967);
or UO_1277 (O_1277,N_29939,N_29481);
or UO_1278 (O_1278,N_29874,N_29625);
and UO_1279 (O_1279,N_29796,N_29465);
nor UO_1280 (O_1280,N_29495,N_29847);
nand UO_1281 (O_1281,N_29483,N_29476);
nand UO_1282 (O_1282,N_29712,N_29499);
xor UO_1283 (O_1283,N_29462,N_29401);
nor UO_1284 (O_1284,N_29855,N_29697);
nor UO_1285 (O_1285,N_29869,N_29509);
xnor UO_1286 (O_1286,N_29761,N_29492);
or UO_1287 (O_1287,N_29834,N_29635);
nand UO_1288 (O_1288,N_29408,N_29989);
xnor UO_1289 (O_1289,N_29658,N_29866);
and UO_1290 (O_1290,N_29723,N_29586);
xnor UO_1291 (O_1291,N_29568,N_29510);
nand UO_1292 (O_1292,N_29493,N_29872);
and UO_1293 (O_1293,N_29667,N_29590);
xnor UO_1294 (O_1294,N_29649,N_29748);
or UO_1295 (O_1295,N_29458,N_29974);
or UO_1296 (O_1296,N_29506,N_29613);
or UO_1297 (O_1297,N_29520,N_29791);
xnor UO_1298 (O_1298,N_29479,N_29750);
or UO_1299 (O_1299,N_29925,N_29678);
or UO_1300 (O_1300,N_29583,N_29534);
nand UO_1301 (O_1301,N_29900,N_29812);
nor UO_1302 (O_1302,N_29759,N_29965);
nor UO_1303 (O_1303,N_29996,N_29902);
xnor UO_1304 (O_1304,N_29639,N_29532);
nor UO_1305 (O_1305,N_29938,N_29773);
xor UO_1306 (O_1306,N_29946,N_29901);
xnor UO_1307 (O_1307,N_29659,N_29505);
nor UO_1308 (O_1308,N_29522,N_29524);
nand UO_1309 (O_1309,N_29656,N_29880);
or UO_1310 (O_1310,N_29993,N_29455);
nor UO_1311 (O_1311,N_29815,N_29766);
nor UO_1312 (O_1312,N_29763,N_29785);
xor UO_1313 (O_1313,N_29599,N_29889);
and UO_1314 (O_1314,N_29503,N_29430);
nand UO_1315 (O_1315,N_29980,N_29801);
xnor UO_1316 (O_1316,N_29877,N_29945);
xnor UO_1317 (O_1317,N_29949,N_29755);
and UO_1318 (O_1318,N_29488,N_29678);
nor UO_1319 (O_1319,N_29915,N_29981);
xnor UO_1320 (O_1320,N_29854,N_29700);
xor UO_1321 (O_1321,N_29644,N_29836);
xor UO_1322 (O_1322,N_29456,N_29621);
nor UO_1323 (O_1323,N_29869,N_29526);
xor UO_1324 (O_1324,N_29506,N_29458);
or UO_1325 (O_1325,N_29493,N_29804);
or UO_1326 (O_1326,N_29964,N_29587);
or UO_1327 (O_1327,N_29658,N_29541);
nand UO_1328 (O_1328,N_29703,N_29734);
nand UO_1329 (O_1329,N_29804,N_29969);
nor UO_1330 (O_1330,N_29734,N_29553);
or UO_1331 (O_1331,N_29890,N_29422);
and UO_1332 (O_1332,N_29529,N_29971);
or UO_1333 (O_1333,N_29799,N_29561);
and UO_1334 (O_1334,N_29998,N_29723);
or UO_1335 (O_1335,N_29635,N_29513);
nor UO_1336 (O_1336,N_29921,N_29464);
xnor UO_1337 (O_1337,N_29727,N_29420);
or UO_1338 (O_1338,N_29710,N_29523);
and UO_1339 (O_1339,N_29459,N_29587);
nor UO_1340 (O_1340,N_29629,N_29848);
nand UO_1341 (O_1341,N_29553,N_29808);
xnor UO_1342 (O_1342,N_29806,N_29572);
and UO_1343 (O_1343,N_29784,N_29461);
and UO_1344 (O_1344,N_29868,N_29794);
or UO_1345 (O_1345,N_29842,N_29746);
nor UO_1346 (O_1346,N_29566,N_29608);
or UO_1347 (O_1347,N_29505,N_29962);
and UO_1348 (O_1348,N_29426,N_29823);
nor UO_1349 (O_1349,N_29619,N_29511);
or UO_1350 (O_1350,N_29839,N_29787);
and UO_1351 (O_1351,N_29844,N_29784);
nand UO_1352 (O_1352,N_29798,N_29484);
xnor UO_1353 (O_1353,N_29750,N_29572);
and UO_1354 (O_1354,N_29921,N_29911);
and UO_1355 (O_1355,N_29938,N_29650);
nor UO_1356 (O_1356,N_29995,N_29922);
nand UO_1357 (O_1357,N_29657,N_29819);
xnor UO_1358 (O_1358,N_29873,N_29910);
nand UO_1359 (O_1359,N_29986,N_29884);
and UO_1360 (O_1360,N_29592,N_29870);
or UO_1361 (O_1361,N_29951,N_29586);
xor UO_1362 (O_1362,N_29639,N_29438);
xnor UO_1363 (O_1363,N_29841,N_29460);
and UO_1364 (O_1364,N_29667,N_29671);
and UO_1365 (O_1365,N_29577,N_29661);
xor UO_1366 (O_1366,N_29924,N_29938);
nor UO_1367 (O_1367,N_29536,N_29816);
nor UO_1368 (O_1368,N_29888,N_29716);
nand UO_1369 (O_1369,N_29731,N_29604);
and UO_1370 (O_1370,N_29643,N_29844);
nor UO_1371 (O_1371,N_29797,N_29763);
or UO_1372 (O_1372,N_29517,N_29594);
nand UO_1373 (O_1373,N_29926,N_29996);
nor UO_1374 (O_1374,N_29843,N_29461);
xnor UO_1375 (O_1375,N_29762,N_29992);
nor UO_1376 (O_1376,N_29403,N_29789);
xor UO_1377 (O_1377,N_29899,N_29568);
nand UO_1378 (O_1378,N_29486,N_29925);
nand UO_1379 (O_1379,N_29890,N_29415);
nor UO_1380 (O_1380,N_29705,N_29690);
nor UO_1381 (O_1381,N_29713,N_29424);
or UO_1382 (O_1382,N_29912,N_29512);
xor UO_1383 (O_1383,N_29799,N_29785);
and UO_1384 (O_1384,N_29652,N_29754);
and UO_1385 (O_1385,N_29818,N_29790);
or UO_1386 (O_1386,N_29887,N_29440);
and UO_1387 (O_1387,N_29653,N_29498);
nor UO_1388 (O_1388,N_29686,N_29428);
or UO_1389 (O_1389,N_29752,N_29679);
and UO_1390 (O_1390,N_29475,N_29651);
nand UO_1391 (O_1391,N_29519,N_29544);
nor UO_1392 (O_1392,N_29571,N_29555);
nand UO_1393 (O_1393,N_29768,N_29800);
or UO_1394 (O_1394,N_29951,N_29874);
nand UO_1395 (O_1395,N_29700,N_29642);
and UO_1396 (O_1396,N_29837,N_29710);
xnor UO_1397 (O_1397,N_29821,N_29816);
or UO_1398 (O_1398,N_29489,N_29697);
or UO_1399 (O_1399,N_29449,N_29764);
nor UO_1400 (O_1400,N_29796,N_29647);
nand UO_1401 (O_1401,N_29954,N_29627);
xnor UO_1402 (O_1402,N_29633,N_29835);
nor UO_1403 (O_1403,N_29420,N_29561);
and UO_1404 (O_1404,N_29843,N_29447);
nor UO_1405 (O_1405,N_29803,N_29697);
and UO_1406 (O_1406,N_29475,N_29896);
nand UO_1407 (O_1407,N_29798,N_29560);
xnor UO_1408 (O_1408,N_29650,N_29566);
nand UO_1409 (O_1409,N_29986,N_29598);
or UO_1410 (O_1410,N_29516,N_29444);
and UO_1411 (O_1411,N_29866,N_29577);
xnor UO_1412 (O_1412,N_29526,N_29491);
and UO_1413 (O_1413,N_29666,N_29722);
and UO_1414 (O_1414,N_29804,N_29834);
or UO_1415 (O_1415,N_29719,N_29980);
or UO_1416 (O_1416,N_29891,N_29638);
and UO_1417 (O_1417,N_29433,N_29630);
and UO_1418 (O_1418,N_29469,N_29730);
and UO_1419 (O_1419,N_29756,N_29731);
or UO_1420 (O_1420,N_29474,N_29419);
xor UO_1421 (O_1421,N_29528,N_29669);
nand UO_1422 (O_1422,N_29745,N_29570);
nor UO_1423 (O_1423,N_29523,N_29553);
and UO_1424 (O_1424,N_29907,N_29587);
xor UO_1425 (O_1425,N_29686,N_29617);
and UO_1426 (O_1426,N_29477,N_29800);
nor UO_1427 (O_1427,N_29857,N_29868);
xor UO_1428 (O_1428,N_29961,N_29506);
nand UO_1429 (O_1429,N_29512,N_29866);
xnor UO_1430 (O_1430,N_29464,N_29828);
nand UO_1431 (O_1431,N_29846,N_29935);
nor UO_1432 (O_1432,N_29808,N_29801);
xor UO_1433 (O_1433,N_29897,N_29830);
and UO_1434 (O_1434,N_29955,N_29836);
or UO_1435 (O_1435,N_29715,N_29523);
and UO_1436 (O_1436,N_29613,N_29775);
xnor UO_1437 (O_1437,N_29578,N_29738);
xor UO_1438 (O_1438,N_29436,N_29631);
xnor UO_1439 (O_1439,N_29621,N_29798);
or UO_1440 (O_1440,N_29571,N_29791);
nand UO_1441 (O_1441,N_29813,N_29872);
nand UO_1442 (O_1442,N_29813,N_29860);
xor UO_1443 (O_1443,N_29623,N_29624);
nor UO_1444 (O_1444,N_29442,N_29696);
xor UO_1445 (O_1445,N_29913,N_29408);
nor UO_1446 (O_1446,N_29922,N_29459);
nor UO_1447 (O_1447,N_29592,N_29658);
or UO_1448 (O_1448,N_29646,N_29468);
nand UO_1449 (O_1449,N_29833,N_29698);
nand UO_1450 (O_1450,N_29854,N_29816);
nand UO_1451 (O_1451,N_29702,N_29537);
and UO_1452 (O_1452,N_29724,N_29669);
or UO_1453 (O_1453,N_29868,N_29440);
nor UO_1454 (O_1454,N_29964,N_29785);
xnor UO_1455 (O_1455,N_29823,N_29833);
nor UO_1456 (O_1456,N_29905,N_29936);
or UO_1457 (O_1457,N_29771,N_29510);
nand UO_1458 (O_1458,N_29426,N_29731);
and UO_1459 (O_1459,N_29445,N_29545);
and UO_1460 (O_1460,N_29537,N_29951);
or UO_1461 (O_1461,N_29963,N_29981);
and UO_1462 (O_1462,N_29927,N_29873);
nor UO_1463 (O_1463,N_29636,N_29417);
or UO_1464 (O_1464,N_29552,N_29835);
xnor UO_1465 (O_1465,N_29610,N_29539);
nand UO_1466 (O_1466,N_29480,N_29935);
and UO_1467 (O_1467,N_29774,N_29421);
and UO_1468 (O_1468,N_29814,N_29454);
or UO_1469 (O_1469,N_29692,N_29799);
xor UO_1470 (O_1470,N_29852,N_29639);
nor UO_1471 (O_1471,N_29842,N_29961);
or UO_1472 (O_1472,N_29551,N_29561);
nand UO_1473 (O_1473,N_29837,N_29585);
and UO_1474 (O_1474,N_29696,N_29589);
nor UO_1475 (O_1475,N_29737,N_29715);
and UO_1476 (O_1476,N_29759,N_29748);
nor UO_1477 (O_1477,N_29688,N_29561);
nand UO_1478 (O_1478,N_29686,N_29534);
nand UO_1479 (O_1479,N_29518,N_29925);
or UO_1480 (O_1480,N_29634,N_29619);
or UO_1481 (O_1481,N_29428,N_29976);
nand UO_1482 (O_1482,N_29681,N_29665);
nand UO_1483 (O_1483,N_29950,N_29601);
xnor UO_1484 (O_1484,N_29479,N_29449);
nand UO_1485 (O_1485,N_29891,N_29424);
and UO_1486 (O_1486,N_29849,N_29731);
nand UO_1487 (O_1487,N_29908,N_29729);
xnor UO_1488 (O_1488,N_29996,N_29685);
and UO_1489 (O_1489,N_29952,N_29890);
or UO_1490 (O_1490,N_29571,N_29735);
and UO_1491 (O_1491,N_29486,N_29584);
or UO_1492 (O_1492,N_29779,N_29949);
nand UO_1493 (O_1493,N_29795,N_29886);
or UO_1494 (O_1494,N_29936,N_29965);
or UO_1495 (O_1495,N_29889,N_29675);
nand UO_1496 (O_1496,N_29502,N_29950);
and UO_1497 (O_1497,N_29696,N_29561);
or UO_1498 (O_1498,N_29997,N_29988);
and UO_1499 (O_1499,N_29800,N_29806);
nor UO_1500 (O_1500,N_29774,N_29498);
and UO_1501 (O_1501,N_29805,N_29583);
xor UO_1502 (O_1502,N_29532,N_29945);
nor UO_1503 (O_1503,N_29607,N_29532);
nor UO_1504 (O_1504,N_29940,N_29913);
nand UO_1505 (O_1505,N_29407,N_29898);
nor UO_1506 (O_1506,N_29516,N_29426);
nand UO_1507 (O_1507,N_29469,N_29770);
and UO_1508 (O_1508,N_29910,N_29541);
and UO_1509 (O_1509,N_29810,N_29733);
or UO_1510 (O_1510,N_29703,N_29804);
nand UO_1511 (O_1511,N_29478,N_29863);
xor UO_1512 (O_1512,N_29576,N_29951);
nor UO_1513 (O_1513,N_29420,N_29456);
and UO_1514 (O_1514,N_29920,N_29512);
xor UO_1515 (O_1515,N_29903,N_29547);
or UO_1516 (O_1516,N_29498,N_29578);
nor UO_1517 (O_1517,N_29619,N_29760);
xnor UO_1518 (O_1518,N_29483,N_29446);
nand UO_1519 (O_1519,N_29440,N_29412);
xor UO_1520 (O_1520,N_29599,N_29765);
nand UO_1521 (O_1521,N_29407,N_29703);
and UO_1522 (O_1522,N_29865,N_29881);
nor UO_1523 (O_1523,N_29562,N_29755);
or UO_1524 (O_1524,N_29966,N_29525);
nor UO_1525 (O_1525,N_29588,N_29959);
or UO_1526 (O_1526,N_29495,N_29759);
and UO_1527 (O_1527,N_29893,N_29534);
xor UO_1528 (O_1528,N_29876,N_29959);
nand UO_1529 (O_1529,N_29904,N_29450);
xnor UO_1530 (O_1530,N_29789,N_29672);
nor UO_1531 (O_1531,N_29699,N_29497);
or UO_1532 (O_1532,N_29550,N_29694);
and UO_1533 (O_1533,N_29676,N_29896);
and UO_1534 (O_1534,N_29475,N_29748);
nor UO_1535 (O_1535,N_29444,N_29628);
xnor UO_1536 (O_1536,N_29764,N_29932);
nand UO_1537 (O_1537,N_29646,N_29954);
and UO_1538 (O_1538,N_29964,N_29844);
or UO_1539 (O_1539,N_29840,N_29838);
xor UO_1540 (O_1540,N_29998,N_29947);
or UO_1541 (O_1541,N_29576,N_29972);
xor UO_1542 (O_1542,N_29954,N_29843);
nand UO_1543 (O_1543,N_29644,N_29470);
nand UO_1544 (O_1544,N_29829,N_29637);
nand UO_1545 (O_1545,N_29706,N_29503);
nand UO_1546 (O_1546,N_29829,N_29432);
or UO_1547 (O_1547,N_29556,N_29905);
nand UO_1548 (O_1548,N_29993,N_29920);
and UO_1549 (O_1549,N_29494,N_29837);
nand UO_1550 (O_1550,N_29676,N_29764);
and UO_1551 (O_1551,N_29556,N_29931);
nor UO_1552 (O_1552,N_29493,N_29584);
or UO_1553 (O_1553,N_29913,N_29887);
or UO_1554 (O_1554,N_29872,N_29833);
or UO_1555 (O_1555,N_29821,N_29409);
and UO_1556 (O_1556,N_29902,N_29450);
or UO_1557 (O_1557,N_29994,N_29983);
nor UO_1558 (O_1558,N_29923,N_29436);
or UO_1559 (O_1559,N_29669,N_29881);
and UO_1560 (O_1560,N_29456,N_29430);
nor UO_1561 (O_1561,N_29610,N_29816);
or UO_1562 (O_1562,N_29918,N_29590);
or UO_1563 (O_1563,N_29699,N_29763);
or UO_1564 (O_1564,N_29418,N_29852);
or UO_1565 (O_1565,N_29940,N_29690);
nand UO_1566 (O_1566,N_29627,N_29656);
xor UO_1567 (O_1567,N_29786,N_29404);
nand UO_1568 (O_1568,N_29568,N_29876);
nand UO_1569 (O_1569,N_29965,N_29770);
nor UO_1570 (O_1570,N_29938,N_29621);
and UO_1571 (O_1571,N_29552,N_29785);
nand UO_1572 (O_1572,N_29644,N_29415);
xnor UO_1573 (O_1573,N_29796,N_29759);
nor UO_1574 (O_1574,N_29438,N_29750);
and UO_1575 (O_1575,N_29460,N_29709);
nor UO_1576 (O_1576,N_29976,N_29855);
or UO_1577 (O_1577,N_29566,N_29485);
nand UO_1578 (O_1578,N_29856,N_29841);
or UO_1579 (O_1579,N_29524,N_29990);
nand UO_1580 (O_1580,N_29458,N_29577);
or UO_1581 (O_1581,N_29716,N_29627);
xnor UO_1582 (O_1582,N_29482,N_29855);
nor UO_1583 (O_1583,N_29515,N_29761);
nor UO_1584 (O_1584,N_29921,N_29719);
and UO_1585 (O_1585,N_29882,N_29817);
xor UO_1586 (O_1586,N_29720,N_29762);
xnor UO_1587 (O_1587,N_29477,N_29779);
and UO_1588 (O_1588,N_29763,N_29958);
and UO_1589 (O_1589,N_29770,N_29430);
and UO_1590 (O_1590,N_29404,N_29901);
nand UO_1591 (O_1591,N_29732,N_29866);
or UO_1592 (O_1592,N_29758,N_29756);
and UO_1593 (O_1593,N_29787,N_29880);
nor UO_1594 (O_1594,N_29983,N_29774);
xor UO_1595 (O_1595,N_29896,N_29635);
nand UO_1596 (O_1596,N_29842,N_29851);
or UO_1597 (O_1597,N_29513,N_29577);
xnor UO_1598 (O_1598,N_29678,N_29758);
nor UO_1599 (O_1599,N_29528,N_29650);
nand UO_1600 (O_1600,N_29941,N_29722);
or UO_1601 (O_1601,N_29685,N_29535);
and UO_1602 (O_1602,N_29831,N_29973);
and UO_1603 (O_1603,N_29433,N_29606);
nor UO_1604 (O_1604,N_29468,N_29665);
nand UO_1605 (O_1605,N_29854,N_29976);
nand UO_1606 (O_1606,N_29875,N_29585);
and UO_1607 (O_1607,N_29918,N_29450);
nand UO_1608 (O_1608,N_29951,N_29536);
or UO_1609 (O_1609,N_29864,N_29739);
and UO_1610 (O_1610,N_29598,N_29422);
xor UO_1611 (O_1611,N_29494,N_29762);
xor UO_1612 (O_1612,N_29538,N_29572);
nand UO_1613 (O_1613,N_29454,N_29744);
and UO_1614 (O_1614,N_29474,N_29882);
nand UO_1615 (O_1615,N_29505,N_29888);
nor UO_1616 (O_1616,N_29969,N_29712);
nor UO_1617 (O_1617,N_29901,N_29750);
nor UO_1618 (O_1618,N_29969,N_29775);
xnor UO_1619 (O_1619,N_29992,N_29898);
nand UO_1620 (O_1620,N_29906,N_29837);
nand UO_1621 (O_1621,N_29454,N_29819);
xor UO_1622 (O_1622,N_29892,N_29613);
nand UO_1623 (O_1623,N_29984,N_29633);
xnor UO_1624 (O_1624,N_29487,N_29720);
or UO_1625 (O_1625,N_29930,N_29942);
and UO_1626 (O_1626,N_29862,N_29675);
or UO_1627 (O_1627,N_29594,N_29529);
nor UO_1628 (O_1628,N_29461,N_29961);
xor UO_1629 (O_1629,N_29777,N_29455);
or UO_1630 (O_1630,N_29623,N_29796);
or UO_1631 (O_1631,N_29591,N_29875);
and UO_1632 (O_1632,N_29741,N_29865);
or UO_1633 (O_1633,N_29438,N_29846);
and UO_1634 (O_1634,N_29655,N_29811);
and UO_1635 (O_1635,N_29760,N_29433);
and UO_1636 (O_1636,N_29643,N_29728);
or UO_1637 (O_1637,N_29451,N_29916);
and UO_1638 (O_1638,N_29450,N_29465);
nand UO_1639 (O_1639,N_29858,N_29452);
or UO_1640 (O_1640,N_29435,N_29762);
and UO_1641 (O_1641,N_29824,N_29849);
nand UO_1642 (O_1642,N_29726,N_29457);
or UO_1643 (O_1643,N_29713,N_29677);
nor UO_1644 (O_1644,N_29478,N_29821);
nor UO_1645 (O_1645,N_29577,N_29990);
nor UO_1646 (O_1646,N_29709,N_29554);
nor UO_1647 (O_1647,N_29669,N_29433);
nand UO_1648 (O_1648,N_29483,N_29420);
nor UO_1649 (O_1649,N_29552,N_29727);
nand UO_1650 (O_1650,N_29768,N_29934);
nor UO_1651 (O_1651,N_29883,N_29923);
nor UO_1652 (O_1652,N_29864,N_29515);
nand UO_1653 (O_1653,N_29620,N_29921);
nor UO_1654 (O_1654,N_29512,N_29507);
nor UO_1655 (O_1655,N_29498,N_29698);
xor UO_1656 (O_1656,N_29707,N_29503);
and UO_1657 (O_1657,N_29768,N_29446);
or UO_1658 (O_1658,N_29991,N_29579);
nand UO_1659 (O_1659,N_29871,N_29641);
and UO_1660 (O_1660,N_29456,N_29979);
and UO_1661 (O_1661,N_29892,N_29485);
nor UO_1662 (O_1662,N_29567,N_29924);
xor UO_1663 (O_1663,N_29542,N_29915);
xor UO_1664 (O_1664,N_29591,N_29909);
and UO_1665 (O_1665,N_29750,N_29619);
or UO_1666 (O_1666,N_29531,N_29477);
xnor UO_1667 (O_1667,N_29463,N_29766);
and UO_1668 (O_1668,N_29647,N_29725);
or UO_1669 (O_1669,N_29857,N_29663);
xnor UO_1670 (O_1670,N_29590,N_29864);
or UO_1671 (O_1671,N_29501,N_29655);
and UO_1672 (O_1672,N_29489,N_29594);
or UO_1673 (O_1673,N_29797,N_29770);
or UO_1674 (O_1674,N_29520,N_29491);
xor UO_1675 (O_1675,N_29740,N_29458);
and UO_1676 (O_1676,N_29751,N_29485);
nor UO_1677 (O_1677,N_29724,N_29636);
xnor UO_1678 (O_1678,N_29967,N_29859);
nor UO_1679 (O_1679,N_29946,N_29679);
xnor UO_1680 (O_1680,N_29474,N_29712);
nor UO_1681 (O_1681,N_29768,N_29799);
and UO_1682 (O_1682,N_29896,N_29707);
xor UO_1683 (O_1683,N_29888,N_29910);
xor UO_1684 (O_1684,N_29940,N_29995);
xnor UO_1685 (O_1685,N_29562,N_29621);
xor UO_1686 (O_1686,N_29939,N_29529);
nor UO_1687 (O_1687,N_29684,N_29439);
xnor UO_1688 (O_1688,N_29703,N_29917);
xnor UO_1689 (O_1689,N_29917,N_29559);
xor UO_1690 (O_1690,N_29635,N_29601);
nand UO_1691 (O_1691,N_29496,N_29859);
nor UO_1692 (O_1692,N_29932,N_29566);
nand UO_1693 (O_1693,N_29775,N_29487);
nor UO_1694 (O_1694,N_29584,N_29981);
or UO_1695 (O_1695,N_29529,N_29757);
nand UO_1696 (O_1696,N_29953,N_29936);
nor UO_1697 (O_1697,N_29577,N_29453);
nand UO_1698 (O_1698,N_29477,N_29512);
or UO_1699 (O_1699,N_29945,N_29989);
or UO_1700 (O_1700,N_29401,N_29530);
xor UO_1701 (O_1701,N_29555,N_29755);
or UO_1702 (O_1702,N_29528,N_29412);
and UO_1703 (O_1703,N_29504,N_29638);
xnor UO_1704 (O_1704,N_29711,N_29454);
xor UO_1705 (O_1705,N_29788,N_29805);
nor UO_1706 (O_1706,N_29752,N_29567);
xnor UO_1707 (O_1707,N_29684,N_29512);
xor UO_1708 (O_1708,N_29808,N_29524);
xnor UO_1709 (O_1709,N_29923,N_29780);
or UO_1710 (O_1710,N_29800,N_29583);
nand UO_1711 (O_1711,N_29837,N_29979);
and UO_1712 (O_1712,N_29742,N_29731);
nor UO_1713 (O_1713,N_29488,N_29973);
nor UO_1714 (O_1714,N_29461,N_29445);
or UO_1715 (O_1715,N_29480,N_29436);
nand UO_1716 (O_1716,N_29980,N_29796);
nor UO_1717 (O_1717,N_29853,N_29962);
nor UO_1718 (O_1718,N_29968,N_29549);
nand UO_1719 (O_1719,N_29787,N_29952);
nand UO_1720 (O_1720,N_29409,N_29875);
xor UO_1721 (O_1721,N_29429,N_29419);
and UO_1722 (O_1722,N_29668,N_29745);
and UO_1723 (O_1723,N_29647,N_29759);
or UO_1724 (O_1724,N_29795,N_29679);
nand UO_1725 (O_1725,N_29949,N_29880);
nor UO_1726 (O_1726,N_29557,N_29548);
and UO_1727 (O_1727,N_29674,N_29942);
or UO_1728 (O_1728,N_29956,N_29983);
xor UO_1729 (O_1729,N_29929,N_29585);
xnor UO_1730 (O_1730,N_29886,N_29744);
nor UO_1731 (O_1731,N_29788,N_29777);
nor UO_1732 (O_1732,N_29593,N_29495);
nand UO_1733 (O_1733,N_29648,N_29973);
xnor UO_1734 (O_1734,N_29435,N_29814);
xnor UO_1735 (O_1735,N_29892,N_29775);
and UO_1736 (O_1736,N_29522,N_29561);
and UO_1737 (O_1737,N_29428,N_29681);
nor UO_1738 (O_1738,N_29807,N_29728);
and UO_1739 (O_1739,N_29583,N_29628);
or UO_1740 (O_1740,N_29823,N_29736);
nand UO_1741 (O_1741,N_29962,N_29637);
nor UO_1742 (O_1742,N_29911,N_29959);
or UO_1743 (O_1743,N_29892,N_29801);
nand UO_1744 (O_1744,N_29770,N_29520);
or UO_1745 (O_1745,N_29773,N_29611);
xnor UO_1746 (O_1746,N_29558,N_29450);
or UO_1747 (O_1747,N_29839,N_29510);
xor UO_1748 (O_1748,N_29878,N_29573);
and UO_1749 (O_1749,N_29621,N_29639);
xor UO_1750 (O_1750,N_29926,N_29419);
nand UO_1751 (O_1751,N_29472,N_29554);
nor UO_1752 (O_1752,N_29481,N_29734);
nand UO_1753 (O_1753,N_29468,N_29863);
nor UO_1754 (O_1754,N_29427,N_29728);
or UO_1755 (O_1755,N_29835,N_29818);
nand UO_1756 (O_1756,N_29576,N_29514);
and UO_1757 (O_1757,N_29957,N_29908);
nand UO_1758 (O_1758,N_29743,N_29557);
nor UO_1759 (O_1759,N_29412,N_29875);
or UO_1760 (O_1760,N_29493,N_29446);
nor UO_1761 (O_1761,N_29657,N_29872);
nand UO_1762 (O_1762,N_29537,N_29666);
or UO_1763 (O_1763,N_29857,N_29749);
xnor UO_1764 (O_1764,N_29592,N_29971);
xnor UO_1765 (O_1765,N_29819,N_29551);
nand UO_1766 (O_1766,N_29970,N_29888);
and UO_1767 (O_1767,N_29765,N_29635);
or UO_1768 (O_1768,N_29820,N_29980);
or UO_1769 (O_1769,N_29619,N_29699);
nor UO_1770 (O_1770,N_29702,N_29657);
or UO_1771 (O_1771,N_29616,N_29491);
or UO_1772 (O_1772,N_29658,N_29630);
or UO_1773 (O_1773,N_29997,N_29887);
and UO_1774 (O_1774,N_29855,N_29520);
nor UO_1775 (O_1775,N_29538,N_29839);
nor UO_1776 (O_1776,N_29779,N_29933);
nor UO_1777 (O_1777,N_29598,N_29833);
xor UO_1778 (O_1778,N_29652,N_29447);
nor UO_1779 (O_1779,N_29590,N_29892);
nor UO_1780 (O_1780,N_29967,N_29504);
xnor UO_1781 (O_1781,N_29826,N_29875);
and UO_1782 (O_1782,N_29956,N_29668);
xnor UO_1783 (O_1783,N_29464,N_29570);
and UO_1784 (O_1784,N_29803,N_29714);
and UO_1785 (O_1785,N_29738,N_29605);
and UO_1786 (O_1786,N_29593,N_29528);
nand UO_1787 (O_1787,N_29640,N_29469);
xor UO_1788 (O_1788,N_29985,N_29509);
xor UO_1789 (O_1789,N_29778,N_29486);
or UO_1790 (O_1790,N_29666,N_29530);
xnor UO_1791 (O_1791,N_29589,N_29716);
nor UO_1792 (O_1792,N_29887,N_29709);
and UO_1793 (O_1793,N_29685,N_29771);
nor UO_1794 (O_1794,N_29535,N_29664);
and UO_1795 (O_1795,N_29504,N_29550);
nand UO_1796 (O_1796,N_29625,N_29633);
and UO_1797 (O_1797,N_29971,N_29560);
xor UO_1798 (O_1798,N_29762,N_29624);
and UO_1799 (O_1799,N_29780,N_29755);
xor UO_1800 (O_1800,N_29945,N_29450);
xor UO_1801 (O_1801,N_29511,N_29705);
nand UO_1802 (O_1802,N_29518,N_29988);
and UO_1803 (O_1803,N_29772,N_29948);
nor UO_1804 (O_1804,N_29935,N_29985);
nor UO_1805 (O_1805,N_29475,N_29558);
nand UO_1806 (O_1806,N_29820,N_29543);
and UO_1807 (O_1807,N_29926,N_29987);
xnor UO_1808 (O_1808,N_29513,N_29631);
or UO_1809 (O_1809,N_29733,N_29972);
nor UO_1810 (O_1810,N_29766,N_29807);
and UO_1811 (O_1811,N_29836,N_29530);
xnor UO_1812 (O_1812,N_29437,N_29907);
and UO_1813 (O_1813,N_29547,N_29410);
nor UO_1814 (O_1814,N_29428,N_29420);
or UO_1815 (O_1815,N_29779,N_29947);
or UO_1816 (O_1816,N_29940,N_29798);
nand UO_1817 (O_1817,N_29428,N_29899);
or UO_1818 (O_1818,N_29891,N_29952);
and UO_1819 (O_1819,N_29913,N_29529);
xor UO_1820 (O_1820,N_29514,N_29953);
nor UO_1821 (O_1821,N_29911,N_29969);
nand UO_1822 (O_1822,N_29892,N_29885);
xor UO_1823 (O_1823,N_29590,N_29634);
or UO_1824 (O_1824,N_29834,N_29828);
nand UO_1825 (O_1825,N_29444,N_29848);
or UO_1826 (O_1826,N_29424,N_29529);
nor UO_1827 (O_1827,N_29945,N_29484);
xor UO_1828 (O_1828,N_29570,N_29991);
or UO_1829 (O_1829,N_29825,N_29705);
xor UO_1830 (O_1830,N_29562,N_29514);
nand UO_1831 (O_1831,N_29582,N_29408);
xnor UO_1832 (O_1832,N_29890,N_29679);
xor UO_1833 (O_1833,N_29493,N_29687);
nand UO_1834 (O_1834,N_29785,N_29810);
nor UO_1835 (O_1835,N_29510,N_29466);
nand UO_1836 (O_1836,N_29829,N_29422);
or UO_1837 (O_1837,N_29875,N_29573);
or UO_1838 (O_1838,N_29570,N_29856);
or UO_1839 (O_1839,N_29540,N_29655);
or UO_1840 (O_1840,N_29436,N_29953);
nor UO_1841 (O_1841,N_29809,N_29534);
xor UO_1842 (O_1842,N_29576,N_29817);
or UO_1843 (O_1843,N_29816,N_29661);
nor UO_1844 (O_1844,N_29444,N_29736);
nor UO_1845 (O_1845,N_29498,N_29759);
or UO_1846 (O_1846,N_29493,N_29577);
and UO_1847 (O_1847,N_29532,N_29591);
nor UO_1848 (O_1848,N_29889,N_29710);
or UO_1849 (O_1849,N_29630,N_29973);
and UO_1850 (O_1850,N_29738,N_29413);
nand UO_1851 (O_1851,N_29997,N_29949);
nand UO_1852 (O_1852,N_29440,N_29406);
or UO_1853 (O_1853,N_29849,N_29699);
or UO_1854 (O_1854,N_29841,N_29760);
xnor UO_1855 (O_1855,N_29729,N_29945);
and UO_1856 (O_1856,N_29809,N_29462);
and UO_1857 (O_1857,N_29950,N_29709);
xnor UO_1858 (O_1858,N_29558,N_29777);
nor UO_1859 (O_1859,N_29958,N_29789);
and UO_1860 (O_1860,N_29868,N_29487);
nor UO_1861 (O_1861,N_29431,N_29485);
or UO_1862 (O_1862,N_29693,N_29833);
nand UO_1863 (O_1863,N_29460,N_29426);
xnor UO_1864 (O_1864,N_29698,N_29458);
xor UO_1865 (O_1865,N_29975,N_29416);
or UO_1866 (O_1866,N_29732,N_29433);
xnor UO_1867 (O_1867,N_29691,N_29400);
or UO_1868 (O_1868,N_29520,N_29850);
nand UO_1869 (O_1869,N_29975,N_29811);
or UO_1870 (O_1870,N_29425,N_29968);
or UO_1871 (O_1871,N_29409,N_29705);
nor UO_1872 (O_1872,N_29894,N_29734);
nor UO_1873 (O_1873,N_29564,N_29769);
or UO_1874 (O_1874,N_29605,N_29667);
or UO_1875 (O_1875,N_29658,N_29862);
or UO_1876 (O_1876,N_29706,N_29829);
and UO_1877 (O_1877,N_29795,N_29404);
and UO_1878 (O_1878,N_29601,N_29606);
xor UO_1879 (O_1879,N_29782,N_29558);
xor UO_1880 (O_1880,N_29642,N_29644);
xor UO_1881 (O_1881,N_29736,N_29437);
nor UO_1882 (O_1882,N_29943,N_29852);
nor UO_1883 (O_1883,N_29583,N_29646);
nor UO_1884 (O_1884,N_29956,N_29901);
xnor UO_1885 (O_1885,N_29720,N_29836);
nor UO_1886 (O_1886,N_29451,N_29704);
or UO_1887 (O_1887,N_29444,N_29506);
or UO_1888 (O_1888,N_29583,N_29623);
and UO_1889 (O_1889,N_29460,N_29997);
or UO_1890 (O_1890,N_29749,N_29446);
nand UO_1891 (O_1891,N_29893,N_29849);
or UO_1892 (O_1892,N_29822,N_29952);
nor UO_1893 (O_1893,N_29985,N_29652);
nor UO_1894 (O_1894,N_29774,N_29676);
or UO_1895 (O_1895,N_29594,N_29665);
xor UO_1896 (O_1896,N_29896,N_29867);
nor UO_1897 (O_1897,N_29700,N_29957);
and UO_1898 (O_1898,N_29724,N_29428);
xnor UO_1899 (O_1899,N_29592,N_29848);
nand UO_1900 (O_1900,N_29807,N_29466);
and UO_1901 (O_1901,N_29497,N_29550);
nor UO_1902 (O_1902,N_29610,N_29621);
and UO_1903 (O_1903,N_29955,N_29772);
and UO_1904 (O_1904,N_29418,N_29799);
and UO_1905 (O_1905,N_29898,N_29772);
xor UO_1906 (O_1906,N_29470,N_29980);
nand UO_1907 (O_1907,N_29425,N_29551);
or UO_1908 (O_1908,N_29798,N_29556);
and UO_1909 (O_1909,N_29963,N_29749);
xor UO_1910 (O_1910,N_29697,N_29732);
nor UO_1911 (O_1911,N_29939,N_29962);
nand UO_1912 (O_1912,N_29789,N_29962);
nor UO_1913 (O_1913,N_29966,N_29521);
and UO_1914 (O_1914,N_29791,N_29727);
nand UO_1915 (O_1915,N_29405,N_29765);
nand UO_1916 (O_1916,N_29691,N_29903);
or UO_1917 (O_1917,N_29845,N_29963);
nor UO_1918 (O_1918,N_29657,N_29796);
and UO_1919 (O_1919,N_29639,N_29740);
or UO_1920 (O_1920,N_29797,N_29869);
xor UO_1921 (O_1921,N_29563,N_29894);
xnor UO_1922 (O_1922,N_29646,N_29551);
xor UO_1923 (O_1923,N_29767,N_29838);
and UO_1924 (O_1924,N_29875,N_29611);
or UO_1925 (O_1925,N_29895,N_29991);
nor UO_1926 (O_1926,N_29836,N_29757);
xor UO_1927 (O_1927,N_29643,N_29639);
or UO_1928 (O_1928,N_29489,N_29571);
nor UO_1929 (O_1929,N_29874,N_29762);
xnor UO_1930 (O_1930,N_29938,N_29754);
xor UO_1931 (O_1931,N_29888,N_29541);
or UO_1932 (O_1932,N_29959,N_29710);
and UO_1933 (O_1933,N_29738,N_29671);
or UO_1934 (O_1934,N_29530,N_29715);
or UO_1935 (O_1935,N_29501,N_29869);
or UO_1936 (O_1936,N_29856,N_29674);
or UO_1937 (O_1937,N_29557,N_29633);
nand UO_1938 (O_1938,N_29853,N_29815);
nor UO_1939 (O_1939,N_29962,N_29950);
nor UO_1940 (O_1940,N_29908,N_29910);
and UO_1941 (O_1941,N_29544,N_29843);
and UO_1942 (O_1942,N_29641,N_29744);
nand UO_1943 (O_1943,N_29607,N_29783);
nand UO_1944 (O_1944,N_29935,N_29496);
xnor UO_1945 (O_1945,N_29710,N_29744);
xnor UO_1946 (O_1946,N_29942,N_29720);
and UO_1947 (O_1947,N_29732,N_29409);
xor UO_1948 (O_1948,N_29699,N_29510);
xnor UO_1949 (O_1949,N_29462,N_29928);
nor UO_1950 (O_1950,N_29499,N_29719);
and UO_1951 (O_1951,N_29838,N_29923);
and UO_1952 (O_1952,N_29683,N_29897);
or UO_1953 (O_1953,N_29560,N_29504);
xnor UO_1954 (O_1954,N_29405,N_29882);
and UO_1955 (O_1955,N_29920,N_29807);
or UO_1956 (O_1956,N_29900,N_29988);
xnor UO_1957 (O_1957,N_29785,N_29990);
and UO_1958 (O_1958,N_29956,N_29590);
or UO_1959 (O_1959,N_29908,N_29943);
nor UO_1960 (O_1960,N_29701,N_29639);
or UO_1961 (O_1961,N_29983,N_29843);
nor UO_1962 (O_1962,N_29442,N_29756);
or UO_1963 (O_1963,N_29837,N_29935);
or UO_1964 (O_1964,N_29534,N_29417);
and UO_1965 (O_1965,N_29557,N_29691);
nand UO_1966 (O_1966,N_29513,N_29761);
nor UO_1967 (O_1967,N_29952,N_29988);
and UO_1968 (O_1968,N_29718,N_29848);
and UO_1969 (O_1969,N_29510,N_29796);
nand UO_1970 (O_1970,N_29480,N_29999);
or UO_1971 (O_1971,N_29816,N_29931);
nor UO_1972 (O_1972,N_29451,N_29712);
and UO_1973 (O_1973,N_29713,N_29474);
xor UO_1974 (O_1974,N_29590,N_29422);
xor UO_1975 (O_1975,N_29706,N_29995);
nand UO_1976 (O_1976,N_29461,N_29601);
and UO_1977 (O_1977,N_29415,N_29607);
xnor UO_1978 (O_1978,N_29583,N_29966);
nor UO_1979 (O_1979,N_29984,N_29932);
or UO_1980 (O_1980,N_29707,N_29834);
nor UO_1981 (O_1981,N_29853,N_29963);
nand UO_1982 (O_1982,N_29407,N_29887);
or UO_1983 (O_1983,N_29687,N_29934);
and UO_1984 (O_1984,N_29519,N_29669);
and UO_1985 (O_1985,N_29805,N_29920);
nand UO_1986 (O_1986,N_29826,N_29792);
or UO_1987 (O_1987,N_29493,N_29597);
and UO_1988 (O_1988,N_29978,N_29425);
or UO_1989 (O_1989,N_29892,N_29879);
and UO_1990 (O_1990,N_29979,N_29475);
and UO_1991 (O_1991,N_29709,N_29439);
xor UO_1992 (O_1992,N_29638,N_29682);
nand UO_1993 (O_1993,N_29696,N_29668);
xnor UO_1994 (O_1994,N_29755,N_29632);
and UO_1995 (O_1995,N_29502,N_29618);
nor UO_1996 (O_1996,N_29917,N_29467);
xnor UO_1997 (O_1997,N_29804,N_29665);
nor UO_1998 (O_1998,N_29858,N_29449);
nand UO_1999 (O_1999,N_29667,N_29889);
or UO_2000 (O_2000,N_29574,N_29633);
xor UO_2001 (O_2001,N_29999,N_29773);
and UO_2002 (O_2002,N_29527,N_29858);
nand UO_2003 (O_2003,N_29897,N_29576);
and UO_2004 (O_2004,N_29820,N_29518);
or UO_2005 (O_2005,N_29820,N_29754);
xnor UO_2006 (O_2006,N_29625,N_29828);
and UO_2007 (O_2007,N_29765,N_29697);
and UO_2008 (O_2008,N_29403,N_29807);
nor UO_2009 (O_2009,N_29682,N_29405);
nor UO_2010 (O_2010,N_29961,N_29614);
xnor UO_2011 (O_2011,N_29647,N_29883);
xor UO_2012 (O_2012,N_29890,N_29656);
and UO_2013 (O_2013,N_29829,N_29971);
nand UO_2014 (O_2014,N_29440,N_29746);
or UO_2015 (O_2015,N_29502,N_29558);
nor UO_2016 (O_2016,N_29440,N_29606);
nand UO_2017 (O_2017,N_29531,N_29631);
nand UO_2018 (O_2018,N_29914,N_29859);
xnor UO_2019 (O_2019,N_29993,N_29764);
or UO_2020 (O_2020,N_29904,N_29811);
nor UO_2021 (O_2021,N_29420,N_29691);
nor UO_2022 (O_2022,N_29617,N_29931);
nor UO_2023 (O_2023,N_29669,N_29986);
nor UO_2024 (O_2024,N_29430,N_29502);
and UO_2025 (O_2025,N_29802,N_29655);
xnor UO_2026 (O_2026,N_29632,N_29843);
nor UO_2027 (O_2027,N_29797,N_29982);
nand UO_2028 (O_2028,N_29812,N_29595);
xor UO_2029 (O_2029,N_29575,N_29836);
nor UO_2030 (O_2030,N_29821,N_29426);
nand UO_2031 (O_2031,N_29790,N_29901);
nor UO_2032 (O_2032,N_29978,N_29500);
and UO_2033 (O_2033,N_29530,N_29897);
and UO_2034 (O_2034,N_29866,N_29982);
xor UO_2035 (O_2035,N_29470,N_29527);
nor UO_2036 (O_2036,N_29519,N_29419);
xor UO_2037 (O_2037,N_29716,N_29895);
or UO_2038 (O_2038,N_29454,N_29693);
xnor UO_2039 (O_2039,N_29931,N_29738);
xnor UO_2040 (O_2040,N_29460,N_29896);
xnor UO_2041 (O_2041,N_29674,N_29432);
nor UO_2042 (O_2042,N_29819,N_29411);
nor UO_2043 (O_2043,N_29649,N_29950);
nand UO_2044 (O_2044,N_29818,N_29540);
or UO_2045 (O_2045,N_29488,N_29733);
and UO_2046 (O_2046,N_29639,N_29620);
and UO_2047 (O_2047,N_29662,N_29756);
or UO_2048 (O_2048,N_29908,N_29923);
nor UO_2049 (O_2049,N_29968,N_29498);
nand UO_2050 (O_2050,N_29742,N_29861);
xnor UO_2051 (O_2051,N_29590,N_29960);
and UO_2052 (O_2052,N_29759,N_29584);
and UO_2053 (O_2053,N_29948,N_29808);
xor UO_2054 (O_2054,N_29943,N_29563);
and UO_2055 (O_2055,N_29671,N_29839);
xnor UO_2056 (O_2056,N_29993,N_29797);
or UO_2057 (O_2057,N_29785,N_29857);
nand UO_2058 (O_2058,N_29818,N_29478);
or UO_2059 (O_2059,N_29892,N_29909);
nand UO_2060 (O_2060,N_29610,N_29650);
nand UO_2061 (O_2061,N_29876,N_29418);
nand UO_2062 (O_2062,N_29632,N_29983);
nor UO_2063 (O_2063,N_29802,N_29444);
nor UO_2064 (O_2064,N_29923,N_29705);
nor UO_2065 (O_2065,N_29858,N_29746);
nand UO_2066 (O_2066,N_29946,N_29749);
nor UO_2067 (O_2067,N_29995,N_29944);
xor UO_2068 (O_2068,N_29613,N_29897);
nand UO_2069 (O_2069,N_29868,N_29755);
nand UO_2070 (O_2070,N_29415,N_29755);
and UO_2071 (O_2071,N_29715,N_29691);
and UO_2072 (O_2072,N_29977,N_29670);
nor UO_2073 (O_2073,N_29502,N_29457);
nand UO_2074 (O_2074,N_29848,N_29628);
nor UO_2075 (O_2075,N_29506,N_29688);
xor UO_2076 (O_2076,N_29747,N_29840);
nor UO_2077 (O_2077,N_29415,N_29650);
xnor UO_2078 (O_2078,N_29965,N_29447);
xnor UO_2079 (O_2079,N_29754,N_29826);
nor UO_2080 (O_2080,N_29747,N_29485);
nand UO_2081 (O_2081,N_29615,N_29617);
or UO_2082 (O_2082,N_29445,N_29892);
nor UO_2083 (O_2083,N_29744,N_29605);
xnor UO_2084 (O_2084,N_29930,N_29515);
or UO_2085 (O_2085,N_29515,N_29471);
xor UO_2086 (O_2086,N_29714,N_29740);
nor UO_2087 (O_2087,N_29960,N_29418);
or UO_2088 (O_2088,N_29812,N_29828);
or UO_2089 (O_2089,N_29945,N_29501);
nor UO_2090 (O_2090,N_29486,N_29836);
xnor UO_2091 (O_2091,N_29457,N_29966);
nand UO_2092 (O_2092,N_29500,N_29404);
and UO_2093 (O_2093,N_29994,N_29940);
nand UO_2094 (O_2094,N_29451,N_29496);
xnor UO_2095 (O_2095,N_29924,N_29872);
xnor UO_2096 (O_2096,N_29743,N_29865);
nor UO_2097 (O_2097,N_29463,N_29453);
or UO_2098 (O_2098,N_29845,N_29613);
nand UO_2099 (O_2099,N_29410,N_29828);
nand UO_2100 (O_2100,N_29509,N_29965);
or UO_2101 (O_2101,N_29483,N_29457);
and UO_2102 (O_2102,N_29454,N_29494);
or UO_2103 (O_2103,N_29570,N_29579);
nand UO_2104 (O_2104,N_29498,N_29781);
nor UO_2105 (O_2105,N_29889,N_29737);
or UO_2106 (O_2106,N_29952,N_29976);
and UO_2107 (O_2107,N_29484,N_29603);
nand UO_2108 (O_2108,N_29601,N_29757);
and UO_2109 (O_2109,N_29494,N_29742);
xnor UO_2110 (O_2110,N_29497,N_29946);
xnor UO_2111 (O_2111,N_29516,N_29581);
xnor UO_2112 (O_2112,N_29941,N_29984);
nand UO_2113 (O_2113,N_29590,N_29862);
xor UO_2114 (O_2114,N_29772,N_29874);
xnor UO_2115 (O_2115,N_29963,N_29977);
xor UO_2116 (O_2116,N_29658,N_29536);
or UO_2117 (O_2117,N_29664,N_29968);
nand UO_2118 (O_2118,N_29619,N_29548);
xor UO_2119 (O_2119,N_29723,N_29617);
xor UO_2120 (O_2120,N_29853,N_29660);
nor UO_2121 (O_2121,N_29657,N_29668);
xnor UO_2122 (O_2122,N_29603,N_29758);
or UO_2123 (O_2123,N_29839,N_29416);
xnor UO_2124 (O_2124,N_29539,N_29692);
and UO_2125 (O_2125,N_29662,N_29447);
or UO_2126 (O_2126,N_29802,N_29979);
nand UO_2127 (O_2127,N_29987,N_29916);
or UO_2128 (O_2128,N_29924,N_29889);
or UO_2129 (O_2129,N_29646,N_29483);
nand UO_2130 (O_2130,N_29823,N_29888);
and UO_2131 (O_2131,N_29845,N_29615);
and UO_2132 (O_2132,N_29974,N_29521);
nand UO_2133 (O_2133,N_29507,N_29854);
and UO_2134 (O_2134,N_29416,N_29536);
nand UO_2135 (O_2135,N_29461,N_29990);
nor UO_2136 (O_2136,N_29929,N_29619);
nand UO_2137 (O_2137,N_29855,N_29985);
and UO_2138 (O_2138,N_29858,N_29498);
and UO_2139 (O_2139,N_29906,N_29693);
or UO_2140 (O_2140,N_29794,N_29723);
nand UO_2141 (O_2141,N_29908,N_29830);
or UO_2142 (O_2142,N_29897,N_29674);
nor UO_2143 (O_2143,N_29854,N_29983);
xor UO_2144 (O_2144,N_29612,N_29506);
or UO_2145 (O_2145,N_29474,N_29672);
xor UO_2146 (O_2146,N_29544,N_29597);
and UO_2147 (O_2147,N_29563,N_29501);
nor UO_2148 (O_2148,N_29948,N_29814);
nor UO_2149 (O_2149,N_29932,N_29442);
xnor UO_2150 (O_2150,N_29658,N_29602);
nand UO_2151 (O_2151,N_29924,N_29784);
nand UO_2152 (O_2152,N_29432,N_29978);
and UO_2153 (O_2153,N_29590,N_29478);
xnor UO_2154 (O_2154,N_29679,N_29516);
and UO_2155 (O_2155,N_29666,N_29619);
xnor UO_2156 (O_2156,N_29972,N_29942);
or UO_2157 (O_2157,N_29633,N_29732);
nor UO_2158 (O_2158,N_29791,N_29581);
or UO_2159 (O_2159,N_29889,N_29617);
nor UO_2160 (O_2160,N_29536,N_29999);
nand UO_2161 (O_2161,N_29521,N_29512);
xnor UO_2162 (O_2162,N_29724,N_29844);
nor UO_2163 (O_2163,N_29736,N_29992);
nor UO_2164 (O_2164,N_29722,N_29851);
and UO_2165 (O_2165,N_29863,N_29885);
and UO_2166 (O_2166,N_29576,N_29560);
or UO_2167 (O_2167,N_29621,N_29667);
or UO_2168 (O_2168,N_29713,N_29924);
and UO_2169 (O_2169,N_29870,N_29790);
nor UO_2170 (O_2170,N_29888,N_29962);
xnor UO_2171 (O_2171,N_29932,N_29850);
xor UO_2172 (O_2172,N_29492,N_29992);
and UO_2173 (O_2173,N_29604,N_29558);
and UO_2174 (O_2174,N_29411,N_29793);
nor UO_2175 (O_2175,N_29948,N_29694);
and UO_2176 (O_2176,N_29857,N_29913);
and UO_2177 (O_2177,N_29717,N_29705);
nand UO_2178 (O_2178,N_29934,N_29569);
and UO_2179 (O_2179,N_29882,N_29751);
or UO_2180 (O_2180,N_29876,N_29835);
or UO_2181 (O_2181,N_29741,N_29618);
xor UO_2182 (O_2182,N_29729,N_29832);
nand UO_2183 (O_2183,N_29695,N_29703);
and UO_2184 (O_2184,N_29770,N_29706);
xor UO_2185 (O_2185,N_29801,N_29524);
or UO_2186 (O_2186,N_29478,N_29643);
or UO_2187 (O_2187,N_29467,N_29772);
xnor UO_2188 (O_2188,N_29757,N_29584);
or UO_2189 (O_2189,N_29476,N_29791);
or UO_2190 (O_2190,N_29817,N_29412);
nand UO_2191 (O_2191,N_29786,N_29978);
and UO_2192 (O_2192,N_29435,N_29963);
and UO_2193 (O_2193,N_29486,N_29927);
nor UO_2194 (O_2194,N_29571,N_29728);
xnor UO_2195 (O_2195,N_29846,N_29863);
xnor UO_2196 (O_2196,N_29501,N_29537);
xor UO_2197 (O_2197,N_29428,N_29585);
or UO_2198 (O_2198,N_29639,N_29608);
xnor UO_2199 (O_2199,N_29751,N_29506);
xor UO_2200 (O_2200,N_29678,N_29842);
nand UO_2201 (O_2201,N_29505,N_29489);
nor UO_2202 (O_2202,N_29620,N_29874);
xnor UO_2203 (O_2203,N_29788,N_29812);
and UO_2204 (O_2204,N_29725,N_29612);
nand UO_2205 (O_2205,N_29636,N_29827);
nand UO_2206 (O_2206,N_29957,N_29588);
xnor UO_2207 (O_2207,N_29429,N_29438);
xor UO_2208 (O_2208,N_29643,N_29444);
nor UO_2209 (O_2209,N_29796,N_29692);
nor UO_2210 (O_2210,N_29654,N_29971);
xnor UO_2211 (O_2211,N_29832,N_29587);
or UO_2212 (O_2212,N_29850,N_29714);
xnor UO_2213 (O_2213,N_29908,N_29410);
nand UO_2214 (O_2214,N_29719,N_29468);
or UO_2215 (O_2215,N_29885,N_29663);
xor UO_2216 (O_2216,N_29910,N_29932);
nor UO_2217 (O_2217,N_29937,N_29906);
xnor UO_2218 (O_2218,N_29721,N_29701);
nor UO_2219 (O_2219,N_29976,N_29419);
or UO_2220 (O_2220,N_29705,N_29741);
and UO_2221 (O_2221,N_29694,N_29637);
xor UO_2222 (O_2222,N_29916,N_29858);
nor UO_2223 (O_2223,N_29800,N_29900);
xor UO_2224 (O_2224,N_29865,N_29509);
and UO_2225 (O_2225,N_29861,N_29999);
and UO_2226 (O_2226,N_29871,N_29429);
xnor UO_2227 (O_2227,N_29708,N_29933);
xor UO_2228 (O_2228,N_29974,N_29513);
xnor UO_2229 (O_2229,N_29445,N_29432);
nor UO_2230 (O_2230,N_29422,N_29586);
nor UO_2231 (O_2231,N_29784,N_29400);
nor UO_2232 (O_2232,N_29575,N_29861);
nor UO_2233 (O_2233,N_29730,N_29922);
and UO_2234 (O_2234,N_29652,N_29516);
xor UO_2235 (O_2235,N_29962,N_29649);
or UO_2236 (O_2236,N_29428,N_29579);
or UO_2237 (O_2237,N_29413,N_29853);
nor UO_2238 (O_2238,N_29800,N_29991);
xnor UO_2239 (O_2239,N_29414,N_29586);
and UO_2240 (O_2240,N_29798,N_29978);
and UO_2241 (O_2241,N_29624,N_29599);
nor UO_2242 (O_2242,N_29662,N_29840);
xnor UO_2243 (O_2243,N_29780,N_29928);
and UO_2244 (O_2244,N_29516,N_29797);
nor UO_2245 (O_2245,N_29914,N_29868);
xnor UO_2246 (O_2246,N_29488,N_29495);
nor UO_2247 (O_2247,N_29919,N_29822);
nor UO_2248 (O_2248,N_29609,N_29959);
nand UO_2249 (O_2249,N_29839,N_29783);
or UO_2250 (O_2250,N_29960,N_29506);
xnor UO_2251 (O_2251,N_29400,N_29856);
or UO_2252 (O_2252,N_29561,N_29556);
or UO_2253 (O_2253,N_29438,N_29519);
xor UO_2254 (O_2254,N_29829,N_29699);
nand UO_2255 (O_2255,N_29537,N_29929);
and UO_2256 (O_2256,N_29939,N_29853);
or UO_2257 (O_2257,N_29594,N_29812);
nor UO_2258 (O_2258,N_29438,N_29770);
and UO_2259 (O_2259,N_29648,N_29418);
and UO_2260 (O_2260,N_29507,N_29614);
xor UO_2261 (O_2261,N_29505,N_29763);
xor UO_2262 (O_2262,N_29666,N_29759);
or UO_2263 (O_2263,N_29530,N_29653);
nand UO_2264 (O_2264,N_29665,N_29691);
and UO_2265 (O_2265,N_29569,N_29778);
xor UO_2266 (O_2266,N_29577,N_29941);
nand UO_2267 (O_2267,N_29596,N_29707);
or UO_2268 (O_2268,N_29637,N_29747);
nor UO_2269 (O_2269,N_29533,N_29669);
and UO_2270 (O_2270,N_29489,N_29682);
or UO_2271 (O_2271,N_29877,N_29644);
and UO_2272 (O_2272,N_29996,N_29740);
nand UO_2273 (O_2273,N_29757,N_29528);
xor UO_2274 (O_2274,N_29584,N_29953);
nor UO_2275 (O_2275,N_29639,N_29416);
nor UO_2276 (O_2276,N_29629,N_29516);
and UO_2277 (O_2277,N_29917,N_29466);
nand UO_2278 (O_2278,N_29535,N_29949);
or UO_2279 (O_2279,N_29712,N_29471);
xnor UO_2280 (O_2280,N_29551,N_29837);
nor UO_2281 (O_2281,N_29430,N_29871);
nand UO_2282 (O_2282,N_29817,N_29618);
or UO_2283 (O_2283,N_29674,N_29867);
xnor UO_2284 (O_2284,N_29772,N_29956);
or UO_2285 (O_2285,N_29580,N_29841);
nand UO_2286 (O_2286,N_29962,N_29421);
or UO_2287 (O_2287,N_29407,N_29592);
nor UO_2288 (O_2288,N_29429,N_29729);
nor UO_2289 (O_2289,N_29855,N_29668);
xor UO_2290 (O_2290,N_29627,N_29608);
nand UO_2291 (O_2291,N_29647,N_29584);
nand UO_2292 (O_2292,N_29654,N_29979);
nor UO_2293 (O_2293,N_29556,N_29918);
or UO_2294 (O_2294,N_29560,N_29875);
xnor UO_2295 (O_2295,N_29763,N_29619);
and UO_2296 (O_2296,N_29898,N_29921);
xor UO_2297 (O_2297,N_29715,N_29600);
nand UO_2298 (O_2298,N_29680,N_29468);
xnor UO_2299 (O_2299,N_29560,N_29915);
xnor UO_2300 (O_2300,N_29632,N_29794);
nand UO_2301 (O_2301,N_29444,N_29462);
nand UO_2302 (O_2302,N_29605,N_29743);
and UO_2303 (O_2303,N_29414,N_29624);
nand UO_2304 (O_2304,N_29807,N_29733);
nor UO_2305 (O_2305,N_29638,N_29774);
xor UO_2306 (O_2306,N_29442,N_29546);
xor UO_2307 (O_2307,N_29836,N_29745);
and UO_2308 (O_2308,N_29568,N_29770);
nor UO_2309 (O_2309,N_29552,N_29532);
nor UO_2310 (O_2310,N_29654,N_29512);
xor UO_2311 (O_2311,N_29484,N_29846);
or UO_2312 (O_2312,N_29509,N_29884);
or UO_2313 (O_2313,N_29411,N_29800);
xor UO_2314 (O_2314,N_29546,N_29404);
or UO_2315 (O_2315,N_29950,N_29823);
nand UO_2316 (O_2316,N_29815,N_29728);
nand UO_2317 (O_2317,N_29452,N_29591);
or UO_2318 (O_2318,N_29672,N_29415);
xnor UO_2319 (O_2319,N_29870,N_29971);
xnor UO_2320 (O_2320,N_29878,N_29995);
and UO_2321 (O_2321,N_29977,N_29960);
xnor UO_2322 (O_2322,N_29587,N_29970);
nor UO_2323 (O_2323,N_29850,N_29749);
and UO_2324 (O_2324,N_29946,N_29743);
nor UO_2325 (O_2325,N_29943,N_29876);
nor UO_2326 (O_2326,N_29977,N_29480);
and UO_2327 (O_2327,N_29629,N_29713);
xnor UO_2328 (O_2328,N_29450,N_29733);
xnor UO_2329 (O_2329,N_29538,N_29720);
or UO_2330 (O_2330,N_29901,N_29948);
xor UO_2331 (O_2331,N_29833,N_29945);
nor UO_2332 (O_2332,N_29539,N_29436);
xor UO_2333 (O_2333,N_29944,N_29613);
xor UO_2334 (O_2334,N_29862,N_29438);
or UO_2335 (O_2335,N_29455,N_29905);
and UO_2336 (O_2336,N_29835,N_29682);
and UO_2337 (O_2337,N_29884,N_29683);
and UO_2338 (O_2338,N_29467,N_29476);
nor UO_2339 (O_2339,N_29862,N_29677);
nor UO_2340 (O_2340,N_29897,N_29789);
and UO_2341 (O_2341,N_29934,N_29867);
nand UO_2342 (O_2342,N_29472,N_29476);
or UO_2343 (O_2343,N_29503,N_29723);
or UO_2344 (O_2344,N_29916,N_29466);
nor UO_2345 (O_2345,N_29671,N_29501);
or UO_2346 (O_2346,N_29640,N_29419);
nand UO_2347 (O_2347,N_29704,N_29817);
and UO_2348 (O_2348,N_29744,N_29936);
nand UO_2349 (O_2349,N_29465,N_29470);
and UO_2350 (O_2350,N_29711,N_29422);
or UO_2351 (O_2351,N_29517,N_29556);
or UO_2352 (O_2352,N_29483,N_29485);
xor UO_2353 (O_2353,N_29462,N_29578);
xor UO_2354 (O_2354,N_29559,N_29820);
xnor UO_2355 (O_2355,N_29409,N_29542);
or UO_2356 (O_2356,N_29538,N_29702);
nand UO_2357 (O_2357,N_29604,N_29997);
xor UO_2358 (O_2358,N_29511,N_29949);
xnor UO_2359 (O_2359,N_29411,N_29592);
nand UO_2360 (O_2360,N_29897,N_29490);
xnor UO_2361 (O_2361,N_29993,N_29668);
xor UO_2362 (O_2362,N_29546,N_29941);
nand UO_2363 (O_2363,N_29560,N_29508);
and UO_2364 (O_2364,N_29922,N_29926);
nand UO_2365 (O_2365,N_29909,N_29972);
nand UO_2366 (O_2366,N_29629,N_29692);
and UO_2367 (O_2367,N_29790,N_29966);
nand UO_2368 (O_2368,N_29821,N_29499);
nand UO_2369 (O_2369,N_29898,N_29897);
nor UO_2370 (O_2370,N_29696,N_29579);
xor UO_2371 (O_2371,N_29855,N_29893);
xor UO_2372 (O_2372,N_29446,N_29915);
nor UO_2373 (O_2373,N_29900,N_29736);
xnor UO_2374 (O_2374,N_29838,N_29886);
nand UO_2375 (O_2375,N_29554,N_29639);
nor UO_2376 (O_2376,N_29921,N_29698);
and UO_2377 (O_2377,N_29916,N_29853);
xor UO_2378 (O_2378,N_29755,N_29573);
and UO_2379 (O_2379,N_29878,N_29891);
nand UO_2380 (O_2380,N_29541,N_29886);
nand UO_2381 (O_2381,N_29991,N_29866);
nor UO_2382 (O_2382,N_29595,N_29539);
and UO_2383 (O_2383,N_29629,N_29805);
nand UO_2384 (O_2384,N_29813,N_29759);
nand UO_2385 (O_2385,N_29789,N_29934);
xnor UO_2386 (O_2386,N_29955,N_29658);
or UO_2387 (O_2387,N_29839,N_29642);
nand UO_2388 (O_2388,N_29941,N_29791);
xor UO_2389 (O_2389,N_29937,N_29783);
nor UO_2390 (O_2390,N_29855,N_29769);
nor UO_2391 (O_2391,N_29631,N_29569);
and UO_2392 (O_2392,N_29711,N_29792);
or UO_2393 (O_2393,N_29823,N_29403);
nand UO_2394 (O_2394,N_29891,N_29944);
and UO_2395 (O_2395,N_29472,N_29678);
xor UO_2396 (O_2396,N_29699,N_29646);
or UO_2397 (O_2397,N_29771,N_29422);
or UO_2398 (O_2398,N_29862,N_29642);
or UO_2399 (O_2399,N_29666,N_29768);
nand UO_2400 (O_2400,N_29766,N_29854);
nor UO_2401 (O_2401,N_29415,N_29630);
nand UO_2402 (O_2402,N_29786,N_29856);
or UO_2403 (O_2403,N_29628,N_29430);
or UO_2404 (O_2404,N_29928,N_29817);
or UO_2405 (O_2405,N_29975,N_29960);
or UO_2406 (O_2406,N_29812,N_29979);
and UO_2407 (O_2407,N_29886,N_29490);
or UO_2408 (O_2408,N_29780,N_29789);
xor UO_2409 (O_2409,N_29545,N_29514);
xor UO_2410 (O_2410,N_29853,N_29434);
nor UO_2411 (O_2411,N_29419,N_29767);
xor UO_2412 (O_2412,N_29849,N_29966);
or UO_2413 (O_2413,N_29432,N_29784);
xnor UO_2414 (O_2414,N_29979,N_29400);
nor UO_2415 (O_2415,N_29515,N_29542);
nor UO_2416 (O_2416,N_29586,N_29934);
xor UO_2417 (O_2417,N_29641,N_29437);
or UO_2418 (O_2418,N_29514,N_29629);
or UO_2419 (O_2419,N_29520,N_29829);
nand UO_2420 (O_2420,N_29476,N_29490);
and UO_2421 (O_2421,N_29737,N_29942);
nor UO_2422 (O_2422,N_29712,N_29830);
nand UO_2423 (O_2423,N_29754,N_29770);
nand UO_2424 (O_2424,N_29925,N_29712);
nor UO_2425 (O_2425,N_29866,N_29675);
nor UO_2426 (O_2426,N_29733,N_29817);
or UO_2427 (O_2427,N_29782,N_29997);
and UO_2428 (O_2428,N_29730,N_29546);
and UO_2429 (O_2429,N_29851,N_29989);
and UO_2430 (O_2430,N_29570,N_29580);
or UO_2431 (O_2431,N_29767,N_29554);
or UO_2432 (O_2432,N_29786,N_29634);
xnor UO_2433 (O_2433,N_29915,N_29463);
or UO_2434 (O_2434,N_29680,N_29711);
nor UO_2435 (O_2435,N_29754,N_29762);
xnor UO_2436 (O_2436,N_29952,N_29480);
or UO_2437 (O_2437,N_29940,N_29590);
or UO_2438 (O_2438,N_29869,N_29910);
nor UO_2439 (O_2439,N_29605,N_29510);
xor UO_2440 (O_2440,N_29655,N_29764);
or UO_2441 (O_2441,N_29953,N_29540);
or UO_2442 (O_2442,N_29520,N_29999);
or UO_2443 (O_2443,N_29685,N_29435);
nand UO_2444 (O_2444,N_29654,N_29915);
nand UO_2445 (O_2445,N_29643,N_29545);
nor UO_2446 (O_2446,N_29402,N_29448);
nand UO_2447 (O_2447,N_29724,N_29696);
or UO_2448 (O_2448,N_29588,N_29603);
nor UO_2449 (O_2449,N_29510,N_29689);
nand UO_2450 (O_2450,N_29848,N_29402);
xor UO_2451 (O_2451,N_29555,N_29925);
or UO_2452 (O_2452,N_29951,N_29669);
nor UO_2453 (O_2453,N_29569,N_29611);
and UO_2454 (O_2454,N_29618,N_29996);
or UO_2455 (O_2455,N_29757,N_29712);
or UO_2456 (O_2456,N_29687,N_29449);
nor UO_2457 (O_2457,N_29651,N_29448);
nor UO_2458 (O_2458,N_29835,N_29897);
and UO_2459 (O_2459,N_29777,N_29682);
or UO_2460 (O_2460,N_29751,N_29551);
or UO_2461 (O_2461,N_29554,N_29788);
nand UO_2462 (O_2462,N_29754,N_29949);
and UO_2463 (O_2463,N_29441,N_29989);
nor UO_2464 (O_2464,N_29854,N_29784);
nand UO_2465 (O_2465,N_29971,N_29904);
nor UO_2466 (O_2466,N_29780,N_29802);
or UO_2467 (O_2467,N_29489,N_29634);
nor UO_2468 (O_2468,N_29819,N_29866);
xnor UO_2469 (O_2469,N_29811,N_29450);
xor UO_2470 (O_2470,N_29825,N_29839);
nand UO_2471 (O_2471,N_29413,N_29998);
xor UO_2472 (O_2472,N_29492,N_29966);
nor UO_2473 (O_2473,N_29511,N_29856);
or UO_2474 (O_2474,N_29607,N_29467);
and UO_2475 (O_2475,N_29965,N_29909);
xnor UO_2476 (O_2476,N_29480,N_29692);
nor UO_2477 (O_2477,N_29408,N_29996);
nor UO_2478 (O_2478,N_29760,N_29474);
nand UO_2479 (O_2479,N_29562,N_29863);
nor UO_2480 (O_2480,N_29586,N_29846);
xor UO_2481 (O_2481,N_29518,N_29763);
xor UO_2482 (O_2482,N_29468,N_29456);
xnor UO_2483 (O_2483,N_29717,N_29583);
nand UO_2484 (O_2484,N_29671,N_29927);
or UO_2485 (O_2485,N_29833,N_29423);
and UO_2486 (O_2486,N_29428,N_29922);
nand UO_2487 (O_2487,N_29900,N_29441);
xor UO_2488 (O_2488,N_29765,N_29831);
xor UO_2489 (O_2489,N_29476,N_29861);
or UO_2490 (O_2490,N_29435,N_29786);
and UO_2491 (O_2491,N_29923,N_29889);
xnor UO_2492 (O_2492,N_29499,N_29860);
or UO_2493 (O_2493,N_29404,N_29575);
nand UO_2494 (O_2494,N_29419,N_29551);
nand UO_2495 (O_2495,N_29928,N_29516);
nand UO_2496 (O_2496,N_29903,N_29902);
and UO_2497 (O_2497,N_29533,N_29839);
nor UO_2498 (O_2498,N_29664,N_29442);
xnor UO_2499 (O_2499,N_29897,N_29681);
nand UO_2500 (O_2500,N_29958,N_29661);
xor UO_2501 (O_2501,N_29543,N_29984);
xnor UO_2502 (O_2502,N_29662,N_29887);
nand UO_2503 (O_2503,N_29835,N_29631);
and UO_2504 (O_2504,N_29525,N_29446);
xnor UO_2505 (O_2505,N_29485,N_29688);
nor UO_2506 (O_2506,N_29909,N_29881);
and UO_2507 (O_2507,N_29447,N_29432);
nor UO_2508 (O_2508,N_29642,N_29465);
and UO_2509 (O_2509,N_29517,N_29835);
and UO_2510 (O_2510,N_29440,N_29756);
xnor UO_2511 (O_2511,N_29534,N_29868);
and UO_2512 (O_2512,N_29441,N_29492);
or UO_2513 (O_2513,N_29747,N_29740);
and UO_2514 (O_2514,N_29986,N_29928);
nand UO_2515 (O_2515,N_29809,N_29623);
and UO_2516 (O_2516,N_29783,N_29402);
or UO_2517 (O_2517,N_29435,N_29658);
nor UO_2518 (O_2518,N_29762,N_29947);
nand UO_2519 (O_2519,N_29710,N_29790);
and UO_2520 (O_2520,N_29551,N_29989);
nor UO_2521 (O_2521,N_29713,N_29826);
xnor UO_2522 (O_2522,N_29428,N_29425);
and UO_2523 (O_2523,N_29544,N_29937);
and UO_2524 (O_2524,N_29473,N_29938);
nand UO_2525 (O_2525,N_29935,N_29743);
and UO_2526 (O_2526,N_29950,N_29870);
nor UO_2527 (O_2527,N_29545,N_29448);
xor UO_2528 (O_2528,N_29738,N_29635);
xnor UO_2529 (O_2529,N_29492,N_29986);
and UO_2530 (O_2530,N_29401,N_29757);
xnor UO_2531 (O_2531,N_29824,N_29953);
and UO_2532 (O_2532,N_29845,N_29410);
and UO_2533 (O_2533,N_29587,N_29761);
or UO_2534 (O_2534,N_29982,N_29943);
and UO_2535 (O_2535,N_29560,N_29440);
nor UO_2536 (O_2536,N_29844,N_29875);
xor UO_2537 (O_2537,N_29424,N_29509);
nor UO_2538 (O_2538,N_29812,N_29573);
nand UO_2539 (O_2539,N_29960,N_29600);
and UO_2540 (O_2540,N_29703,N_29501);
or UO_2541 (O_2541,N_29798,N_29982);
nand UO_2542 (O_2542,N_29953,N_29589);
or UO_2543 (O_2543,N_29688,N_29589);
and UO_2544 (O_2544,N_29570,N_29593);
nand UO_2545 (O_2545,N_29727,N_29966);
xor UO_2546 (O_2546,N_29898,N_29572);
nand UO_2547 (O_2547,N_29454,N_29677);
or UO_2548 (O_2548,N_29489,N_29776);
nand UO_2549 (O_2549,N_29698,N_29466);
nor UO_2550 (O_2550,N_29857,N_29566);
xor UO_2551 (O_2551,N_29805,N_29551);
nor UO_2552 (O_2552,N_29725,N_29592);
and UO_2553 (O_2553,N_29798,N_29459);
and UO_2554 (O_2554,N_29533,N_29962);
nand UO_2555 (O_2555,N_29663,N_29506);
nand UO_2556 (O_2556,N_29777,N_29414);
xor UO_2557 (O_2557,N_29429,N_29471);
and UO_2558 (O_2558,N_29942,N_29705);
nand UO_2559 (O_2559,N_29729,N_29697);
xnor UO_2560 (O_2560,N_29433,N_29925);
and UO_2561 (O_2561,N_29531,N_29804);
nand UO_2562 (O_2562,N_29556,N_29528);
and UO_2563 (O_2563,N_29513,N_29675);
nor UO_2564 (O_2564,N_29650,N_29705);
nor UO_2565 (O_2565,N_29714,N_29906);
or UO_2566 (O_2566,N_29458,N_29926);
xor UO_2567 (O_2567,N_29849,N_29998);
nand UO_2568 (O_2568,N_29470,N_29724);
nand UO_2569 (O_2569,N_29417,N_29590);
nor UO_2570 (O_2570,N_29818,N_29855);
nor UO_2571 (O_2571,N_29856,N_29418);
xor UO_2572 (O_2572,N_29665,N_29611);
and UO_2573 (O_2573,N_29673,N_29541);
or UO_2574 (O_2574,N_29457,N_29896);
or UO_2575 (O_2575,N_29731,N_29576);
or UO_2576 (O_2576,N_29864,N_29581);
and UO_2577 (O_2577,N_29789,N_29802);
or UO_2578 (O_2578,N_29672,N_29923);
nand UO_2579 (O_2579,N_29973,N_29893);
and UO_2580 (O_2580,N_29569,N_29758);
and UO_2581 (O_2581,N_29808,N_29667);
or UO_2582 (O_2582,N_29603,N_29429);
nor UO_2583 (O_2583,N_29936,N_29735);
nor UO_2584 (O_2584,N_29600,N_29764);
nand UO_2585 (O_2585,N_29436,N_29410);
or UO_2586 (O_2586,N_29498,N_29574);
nor UO_2587 (O_2587,N_29736,N_29486);
xor UO_2588 (O_2588,N_29428,N_29875);
or UO_2589 (O_2589,N_29605,N_29485);
nand UO_2590 (O_2590,N_29470,N_29759);
and UO_2591 (O_2591,N_29638,N_29972);
xor UO_2592 (O_2592,N_29906,N_29658);
or UO_2593 (O_2593,N_29531,N_29708);
or UO_2594 (O_2594,N_29780,N_29952);
nor UO_2595 (O_2595,N_29747,N_29510);
nor UO_2596 (O_2596,N_29532,N_29942);
nand UO_2597 (O_2597,N_29797,N_29426);
nor UO_2598 (O_2598,N_29485,N_29719);
xnor UO_2599 (O_2599,N_29574,N_29948);
nand UO_2600 (O_2600,N_29650,N_29708);
nor UO_2601 (O_2601,N_29725,N_29544);
nor UO_2602 (O_2602,N_29939,N_29400);
and UO_2603 (O_2603,N_29885,N_29893);
or UO_2604 (O_2604,N_29905,N_29795);
nand UO_2605 (O_2605,N_29931,N_29581);
nand UO_2606 (O_2606,N_29587,N_29701);
xnor UO_2607 (O_2607,N_29424,N_29983);
or UO_2608 (O_2608,N_29719,N_29427);
nor UO_2609 (O_2609,N_29515,N_29834);
xor UO_2610 (O_2610,N_29669,N_29773);
or UO_2611 (O_2611,N_29660,N_29840);
and UO_2612 (O_2612,N_29609,N_29817);
and UO_2613 (O_2613,N_29873,N_29824);
nor UO_2614 (O_2614,N_29775,N_29824);
xnor UO_2615 (O_2615,N_29925,N_29931);
or UO_2616 (O_2616,N_29419,N_29511);
or UO_2617 (O_2617,N_29825,N_29853);
and UO_2618 (O_2618,N_29870,N_29630);
or UO_2619 (O_2619,N_29859,N_29476);
xnor UO_2620 (O_2620,N_29797,N_29661);
and UO_2621 (O_2621,N_29624,N_29934);
nor UO_2622 (O_2622,N_29655,N_29434);
and UO_2623 (O_2623,N_29506,N_29515);
and UO_2624 (O_2624,N_29540,N_29699);
nor UO_2625 (O_2625,N_29932,N_29720);
nor UO_2626 (O_2626,N_29932,N_29664);
nand UO_2627 (O_2627,N_29607,N_29638);
nor UO_2628 (O_2628,N_29852,N_29456);
nor UO_2629 (O_2629,N_29722,N_29889);
and UO_2630 (O_2630,N_29645,N_29849);
and UO_2631 (O_2631,N_29767,N_29739);
xor UO_2632 (O_2632,N_29537,N_29672);
nand UO_2633 (O_2633,N_29824,N_29452);
or UO_2634 (O_2634,N_29682,N_29664);
nand UO_2635 (O_2635,N_29567,N_29581);
or UO_2636 (O_2636,N_29799,N_29833);
and UO_2637 (O_2637,N_29500,N_29579);
nand UO_2638 (O_2638,N_29737,N_29911);
nor UO_2639 (O_2639,N_29558,N_29514);
or UO_2640 (O_2640,N_29749,N_29746);
and UO_2641 (O_2641,N_29490,N_29844);
nand UO_2642 (O_2642,N_29418,N_29759);
and UO_2643 (O_2643,N_29764,N_29770);
nand UO_2644 (O_2644,N_29466,N_29815);
xor UO_2645 (O_2645,N_29480,N_29567);
and UO_2646 (O_2646,N_29632,N_29732);
xor UO_2647 (O_2647,N_29910,N_29809);
nor UO_2648 (O_2648,N_29558,N_29987);
or UO_2649 (O_2649,N_29937,N_29901);
nor UO_2650 (O_2650,N_29450,N_29873);
nor UO_2651 (O_2651,N_29813,N_29710);
or UO_2652 (O_2652,N_29781,N_29452);
nand UO_2653 (O_2653,N_29742,N_29716);
and UO_2654 (O_2654,N_29924,N_29519);
and UO_2655 (O_2655,N_29913,N_29588);
nor UO_2656 (O_2656,N_29442,N_29721);
and UO_2657 (O_2657,N_29859,N_29431);
or UO_2658 (O_2658,N_29476,N_29595);
nor UO_2659 (O_2659,N_29853,N_29986);
nor UO_2660 (O_2660,N_29770,N_29898);
nor UO_2661 (O_2661,N_29496,N_29780);
and UO_2662 (O_2662,N_29941,N_29564);
and UO_2663 (O_2663,N_29874,N_29916);
nor UO_2664 (O_2664,N_29957,N_29675);
xnor UO_2665 (O_2665,N_29781,N_29871);
and UO_2666 (O_2666,N_29700,N_29990);
nor UO_2667 (O_2667,N_29412,N_29415);
nand UO_2668 (O_2668,N_29640,N_29422);
or UO_2669 (O_2669,N_29532,N_29662);
and UO_2670 (O_2670,N_29679,N_29774);
and UO_2671 (O_2671,N_29741,N_29409);
and UO_2672 (O_2672,N_29434,N_29916);
nand UO_2673 (O_2673,N_29687,N_29730);
xor UO_2674 (O_2674,N_29872,N_29718);
xnor UO_2675 (O_2675,N_29731,N_29727);
nand UO_2676 (O_2676,N_29988,N_29417);
nor UO_2677 (O_2677,N_29645,N_29905);
or UO_2678 (O_2678,N_29434,N_29639);
nor UO_2679 (O_2679,N_29629,N_29717);
or UO_2680 (O_2680,N_29686,N_29843);
xnor UO_2681 (O_2681,N_29560,N_29750);
xor UO_2682 (O_2682,N_29596,N_29506);
or UO_2683 (O_2683,N_29914,N_29424);
or UO_2684 (O_2684,N_29651,N_29973);
xor UO_2685 (O_2685,N_29970,N_29457);
nand UO_2686 (O_2686,N_29549,N_29452);
xor UO_2687 (O_2687,N_29594,N_29929);
and UO_2688 (O_2688,N_29502,N_29443);
nor UO_2689 (O_2689,N_29404,N_29482);
nand UO_2690 (O_2690,N_29933,N_29980);
or UO_2691 (O_2691,N_29413,N_29493);
or UO_2692 (O_2692,N_29832,N_29588);
or UO_2693 (O_2693,N_29669,N_29527);
or UO_2694 (O_2694,N_29602,N_29847);
xnor UO_2695 (O_2695,N_29774,N_29445);
nand UO_2696 (O_2696,N_29699,N_29553);
nand UO_2697 (O_2697,N_29463,N_29764);
nor UO_2698 (O_2698,N_29697,N_29882);
or UO_2699 (O_2699,N_29938,N_29568);
and UO_2700 (O_2700,N_29890,N_29705);
and UO_2701 (O_2701,N_29780,N_29769);
xnor UO_2702 (O_2702,N_29403,N_29583);
nor UO_2703 (O_2703,N_29642,N_29867);
and UO_2704 (O_2704,N_29638,N_29407);
or UO_2705 (O_2705,N_29933,N_29493);
and UO_2706 (O_2706,N_29713,N_29510);
and UO_2707 (O_2707,N_29866,N_29896);
nand UO_2708 (O_2708,N_29475,N_29864);
xnor UO_2709 (O_2709,N_29868,N_29527);
nor UO_2710 (O_2710,N_29954,N_29410);
or UO_2711 (O_2711,N_29524,N_29951);
nand UO_2712 (O_2712,N_29994,N_29867);
or UO_2713 (O_2713,N_29567,N_29446);
and UO_2714 (O_2714,N_29845,N_29560);
or UO_2715 (O_2715,N_29461,N_29526);
or UO_2716 (O_2716,N_29457,N_29658);
and UO_2717 (O_2717,N_29819,N_29544);
nand UO_2718 (O_2718,N_29819,N_29561);
or UO_2719 (O_2719,N_29728,N_29542);
or UO_2720 (O_2720,N_29931,N_29833);
and UO_2721 (O_2721,N_29921,N_29843);
nor UO_2722 (O_2722,N_29775,N_29925);
nor UO_2723 (O_2723,N_29876,N_29490);
or UO_2724 (O_2724,N_29876,N_29641);
nor UO_2725 (O_2725,N_29400,N_29438);
nor UO_2726 (O_2726,N_29458,N_29905);
nor UO_2727 (O_2727,N_29820,N_29959);
nand UO_2728 (O_2728,N_29834,N_29962);
xor UO_2729 (O_2729,N_29481,N_29759);
nand UO_2730 (O_2730,N_29520,N_29609);
and UO_2731 (O_2731,N_29878,N_29960);
xor UO_2732 (O_2732,N_29568,N_29995);
and UO_2733 (O_2733,N_29441,N_29819);
nand UO_2734 (O_2734,N_29728,N_29478);
nand UO_2735 (O_2735,N_29469,N_29736);
nand UO_2736 (O_2736,N_29907,N_29686);
nand UO_2737 (O_2737,N_29739,N_29533);
and UO_2738 (O_2738,N_29915,N_29810);
xnor UO_2739 (O_2739,N_29416,N_29574);
and UO_2740 (O_2740,N_29409,N_29417);
nor UO_2741 (O_2741,N_29862,N_29958);
nor UO_2742 (O_2742,N_29419,N_29544);
xor UO_2743 (O_2743,N_29917,N_29933);
nor UO_2744 (O_2744,N_29645,N_29462);
and UO_2745 (O_2745,N_29428,N_29658);
and UO_2746 (O_2746,N_29493,N_29899);
and UO_2747 (O_2747,N_29912,N_29927);
nor UO_2748 (O_2748,N_29433,N_29430);
xnor UO_2749 (O_2749,N_29826,N_29859);
or UO_2750 (O_2750,N_29612,N_29910);
xor UO_2751 (O_2751,N_29559,N_29679);
nand UO_2752 (O_2752,N_29591,N_29845);
or UO_2753 (O_2753,N_29534,N_29812);
nor UO_2754 (O_2754,N_29482,N_29782);
nor UO_2755 (O_2755,N_29525,N_29607);
and UO_2756 (O_2756,N_29593,N_29560);
or UO_2757 (O_2757,N_29876,N_29637);
or UO_2758 (O_2758,N_29707,N_29770);
nand UO_2759 (O_2759,N_29402,N_29480);
xor UO_2760 (O_2760,N_29490,N_29417);
or UO_2761 (O_2761,N_29519,N_29695);
and UO_2762 (O_2762,N_29860,N_29463);
and UO_2763 (O_2763,N_29881,N_29611);
or UO_2764 (O_2764,N_29931,N_29497);
and UO_2765 (O_2765,N_29769,N_29760);
or UO_2766 (O_2766,N_29996,N_29506);
xnor UO_2767 (O_2767,N_29513,N_29665);
nand UO_2768 (O_2768,N_29660,N_29722);
or UO_2769 (O_2769,N_29970,N_29575);
nor UO_2770 (O_2770,N_29649,N_29944);
nand UO_2771 (O_2771,N_29749,N_29808);
or UO_2772 (O_2772,N_29464,N_29745);
nand UO_2773 (O_2773,N_29794,N_29525);
nor UO_2774 (O_2774,N_29899,N_29764);
nand UO_2775 (O_2775,N_29918,N_29843);
xor UO_2776 (O_2776,N_29412,N_29854);
or UO_2777 (O_2777,N_29914,N_29993);
xor UO_2778 (O_2778,N_29448,N_29583);
nand UO_2779 (O_2779,N_29577,N_29942);
and UO_2780 (O_2780,N_29893,N_29934);
nor UO_2781 (O_2781,N_29485,N_29977);
nand UO_2782 (O_2782,N_29791,N_29437);
or UO_2783 (O_2783,N_29425,N_29740);
xor UO_2784 (O_2784,N_29933,N_29822);
or UO_2785 (O_2785,N_29937,N_29748);
or UO_2786 (O_2786,N_29809,N_29737);
xnor UO_2787 (O_2787,N_29402,N_29735);
and UO_2788 (O_2788,N_29472,N_29856);
or UO_2789 (O_2789,N_29662,N_29968);
xnor UO_2790 (O_2790,N_29946,N_29636);
or UO_2791 (O_2791,N_29661,N_29665);
xnor UO_2792 (O_2792,N_29953,N_29483);
xnor UO_2793 (O_2793,N_29479,N_29539);
xor UO_2794 (O_2794,N_29680,N_29848);
nand UO_2795 (O_2795,N_29482,N_29830);
and UO_2796 (O_2796,N_29520,N_29871);
or UO_2797 (O_2797,N_29778,N_29741);
xor UO_2798 (O_2798,N_29906,N_29465);
nand UO_2799 (O_2799,N_29887,N_29700);
and UO_2800 (O_2800,N_29729,N_29857);
and UO_2801 (O_2801,N_29998,N_29583);
nor UO_2802 (O_2802,N_29471,N_29875);
or UO_2803 (O_2803,N_29629,N_29475);
nor UO_2804 (O_2804,N_29859,N_29474);
xnor UO_2805 (O_2805,N_29813,N_29524);
and UO_2806 (O_2806,N_29660,N_29954);
and UO_2807 (O_2807,N_29987,N_29959);
or UO_2808 (O_2808,N_29772,N_29906);
xor UO_2809 (O_2809,N_29697,N_29671);
nor UO_2810 (O_2810,N_29990,N_29833);
and UO_2811 (O_2811,N_29685,N_29950);
nor UO_2812 (O_2812,N_29475,N_29697);
and UO_2813 (O_2813,N_29791,N_29736);
nor UO_2814 (O_2814,N_29688,N_29491);
nand UO_2815 (O_2815,N_29703,N_29677);
nand UO_2816 (O_2816,N_29577,N_29684);
or UO_2817 (O_2817,N_29680,N_29972);
or UO_2818 (O_2818,N_29820,N_29484);
and UO_2819 (O_2819,N_29782,N_29833);
or UO_2820 (O_2820,N_29468,N_29797);
and UO_2821 (O_2821,N_29577,N_29731);
xor UO_2822 (O_2822,N_29543,N_29501);
and UO_2823 (O_2823,N_29623,N_29733);
nand UO_2824 (O_2824,N_29873,N_29916);
nor UO_2825 (O_2825,N_29686,N_29665);
or UO_2826 (O_2826,N_29528,N_29510);
xor UO_2827 (O_2827,N_29831,N_29664);
xnor UO_2828 (O_2828,N_29469,N_29435);
or UO_2829 (O_2829,N_29893,N_29907);
nand UO_2830 (O_2830,N_29772,N_29527);
nor UO_2831 (O_2831,N_29802,N_29409);
xnor UO_2832 (O_2832,N_29445,N_29659);
xor UO_2833 (O_2833,N_29566,N_29476);
nand UO_2834 (O_2834,N_29569,N_29568);
or UO_2835 (O_2835,N_29864,N_29737);
nor UO_2836 (O_2836,N_29631,N_29662);
xor UO_2837 (O_2837,N_29880,N_29915);
xor UO_2838 (O_2838,N_29470,N_29651);
nor UO_2839 (O_2839,N_29744,N_29592);
and UO_2840 (O_2840,N_29707,N_29515);
nand UO_2841 (O_2841,N_29781,N_29805);
nor UO_2842 (O_2842,N_29479,N_29821);
nand UO_2843 (O_2843,N_29888,N_29732);
and UO_2844 (O_2844,N_29583,N_29419);
nand UO_2845 (O_2845,N_29890,N_29640);
or UO_2846 (O_2846,N_29921,N_29860);
or UO_2847 (O_2847,N_29620,N_29443);
nor UO_2848 (O_2848,N_29593,N_29591);
xnor UO_2849 (O_2849,N_29549,N_29812);
or UO_2850 (O_2850,N_29675,N_29817);
nor UO_2851 (O_2851,N_29927,N_29813);
nor UO_2852 (O_2852,N_29430,N_29883);
xor UO_2853 (O_2853,N_29585,N_29856);
nor UO_2854 (O_2854,N_29667,N_29929);
nor UO_2855 (O_2855,N_29440,N_29951);
or UO_2856 (O_2856,N_29889,N_29899);
nor UO_2857 (O_2857,N_29856,N_29733);
xor UO_2858 (O_2858,N_29564,N_29902);
or UO_2859 (O_2859,N_29813,N_29817);
or UO_2860 (O_2860,N_29510,N_29711);
nor UO_2861 (O_2861,N_29739,N_29501);
or UO_2862 (O_2862,N_29966,N_29898);
nor UO_2863 (O_2863,N_29946,N_29808);
nor UO_2864 (O_2864,N_29731,N_29965);
nor UO_2865 (O_2865,N_29725,N_29445);
nor UO_2866 (O_2866,N_29838,N_29749);
or UO_2867 (O_2867,N_29522,N_29483);
xnor UO_2868 (O_2868,N_29541,N_29832);
nand UO_2869 (O_2869,N_29701,N_29490);
nor UO_2870 (O_2870,N_29978,N_29488);
and UO_2871 (O_2871,N_29586,N_29609);
nand UO_2872 (O_2872,N_29778,N_29883);
xor UO_2873 (O_2873,N_29766,N_29973);
xnor UO_2874 (O_2874,N_29762,N_29923);
or UO_2875 (O_2875,N_29452,N_29870);
or UO_2876 (O_2876,N_29567,N_29460);
or UO_2877 (O_2877,N_29639,N_29835);
or UO_2878 (O_2878,N_29758,N_29975);
or UO_2879 (O_2879,N_29427,N_29482);
nand UO_2880 (O_2880,N_29964,N_29625);
nor UO_2881 (O_2881,N_29897,N_29453);
nor UO_2882 (O_2882,N_29713,N_29460);
nand UO_2883 (O_2883,N_29540,N_29633);
nor UO_2884 (O_2884,N_29545,N_29923);
and UO_2885 (O_2885,N_29991,N_29517);
nand UO_2886 (O_2886,N_29586,N_29732);
or UO_2887 (O_2887,N_29411,N_29826);
and UO_2888 (O_2888,N_29922,N_29991);
xor UO_2889 (O_2889,N_29877,N_29951);
or UO_2890 (O_2890,N_29824,N_29569);
or UO_2891 (O_2891,N_29641,N_29988);
xnor UO_2892 (O_2892,N_29946,N_29528);
xnor UO_2893 (O_2893,N_29661,N_29705);
nand UO_2894 (O_2894,N_29892,N_29539);
nor UO_2895 (O_2895,N_29529,N_29815);
and UO_2896 (O_2896,N_29865,N_29536);
xnor UO_2897 (O_2897,N_29670,N_29908);
nor UO_2898 (O_2898,N_29801,N_29845);
and UO_2899 (O_2899,N_29858,N_29677);
or UO_2900 (O_2900,N_29944,N_29698);
xnor UO_2901 (O_2901,N_29633,N_29781);
and UO_2902 (O_2902,N_29504,N_29575);
nand UO_2903 (O_2903,N_29418,N_29870);
nor UO_2904 (O_2904,N_29707,N_29645);
and UO_2905 (O_2905,N_29696,N_29773);
nand UO_2906 (O_2906,N_29990,N_29909);
xnor UO_2907 (O_2907,N_29406,N_29625);
nor UO_2908 (O_2908,N_29431,N_29514);
xor UO_2909 (O_2909,N_29876,N_29891);
and UO_2910 (O_2910,N_29688,N_29656);
nand UO_2911 (O_2911,N_29681,N_29580);
or UO_2912 (O_2912,N_29439,N_29421);
nor UO_2913 (O_2913,N_29598,N_29672);
nand UO_2914 (O_2914,N_29761,N_29696);
nor UO_2915 (O_2915,N_29676,N_29409);
xnor UO_2916 (O_2916,N_29640,N_29529);
and UO_2917 (O_2917,N_29947,N_29927);
nand UO_2918 (O_2918,N_29830,N_29696);
nor UO_2919 (O_2919,N_29839,N_29851);
nand UO_2920 (O_2920,N_29547,N_29750);
and UO_2921 (O_2921,N_29939,N_29896);
xor UO_2922 (O_2922,N_29659,N_29684);
nand UO_2923 (O_2923,N_29579,N_29720);
or UO_2924 (O_2924,N_29515,N_29535);
or UO_2925 (O_2925,N_29559,N_29685);
xnor UO_2926 (O_2926,N_29753,N_29793);
nand UO_2927 (O_2927,N_29944,N_29509);
nor UO_2928 (O_2928,N_29410,N_29434);
nor UO_2929 (O_2929,N_29424,N_29405);
or UO_2930 (O_2930,N_29731,N_29423);
or UO_2931 (O_2931,N_29725,N_29628);
or UO_2932 (O_2932,N_29879,N_29912);
and UO_2933 (O_2933,N_29981,N_29763);
nand UO_2934 (O_2934,N_29840,N_29515);
xor UO_2935 (O_2935,N_29891,N_29736);
or UO_2936 (O_2936,N_29979,N_29926);
nor UO_2937 (O_2937,N_29586,N_29709);
nor UO_2938 (O_2938,N_29985,N_29418);
or UO_2939 (O_2939,N_29955,N_29722);
nor UO_2940 (O_2940,N_29941,N_29814);
or UO_2941 (O_2941,N_29498,N_29456);
or UO_2942 (O_2942,N_29988,N_29428);
and UO_2943 (O_2943,N_29712,N_29993);
xor UO_2944 (O_2944,N_29813,N_29789);
and UO_2945 (O_2945,N_29460,N_29644);
and UO_2946 (O_2946,N_29408,N_29762);
and UO_2947 (O_2947,N_29464,N_29738);
nand UO_2948 (O_2948,N_29717,N_29970);
nand UO_2949 (O_2949,N_29736,N_29867);
and UO_2950 (O_2950,N_29452,N_29943);
or UO_2951 (O_2951,N_29897,N_29820);
and UO_2952 (O_2952,N_29698,N_29684);
and UO_2953 (O_2953,N_29610,N_29549);
xor UO_2954 (O_2954,N_29979,N_29553);
xor UO_2955 (O_2955,N_29956,N_29878);
nor UO_2956 (O_2956,N_29582,N_29706);
xor UO_2957 (O_2957,N_29571,N_29903);
xor UO_2958 (O_2958,N_29698,N_29799);
xnor UO_2959 (O_2959,N_29559,N_29706);
xor UO_2960 (O_2960,N_29878,N_29881);
nand UO_2961 (O_2961,N_29567,N_29912);
or UO_2962 (O_2962,N_29736,N_29524);
or UO_2963 (O_2963,N_29764,N_29838);
xnor UO_2964 (O_2964,N_29701,N_29716);
xnor UO_2965 (O_2965,N_29521,N_29968);
and UO_2966 (O_2966,N_29786,N_29581);
or UO_2967 (O_2967,N_29681,N_29718);
or UO_2968 (O_2968,N_29566,N_29647);
nor UO_2969 (O_2969,N_29960,N_29595);
nand UO_2970 (O_2970,N_29679,N_29779);
nor UO_2971 (O_2971,N_29527,N_29927);
nand UO_2972 (O_2972,N_29606,N_29712);
or UO_2973 (O_2973,N_29442,N_29750);
or UO_2974 (O_2974,N_29552,N_29492);
nor UO_2975 (O_2975,N_29608,N_29442);
and UO_2976 (O_2976,N_29834,N_29859);
or UO_2977 (O_2977,N_29616,N_29896);
nand UO_2978 (O_2978,N_29751,N_29728);
or UO_2979 (O_2979,N_29573,N_29904);
nor UO_2980 (O_2980,N_29865,N_29475);
xor UO_2981 (O_2981,N_29900,N_29740);
nor UO_2982 (O_2982,N_29800,N_29492);
xnor UO_2983 (O_2983,N_29499,N_29522);
or UO_2984 (O_2984,N_29866,N_29444);
nor UO_2985 (O_2985,N_29903,N_29735);
nand UO_2986 (O_2986,N_29827,N_29871);
nor UO_2987 (O_2987,N_29430,N_29500);
and UO_2988 (O_2988,N_29755,N_29654);
nor UO_2989 (O_2989,N_29910,N_29408);
or UO_2990 (O_2990,N_29983,N_29829);
and UO_2991 (O_2991,N_29546,N_29974);
nand UO_2992 (O_2992,N_29426,N_29784);
xnor UO_2993 (O_2993,N_29853,N_29823);
nand UO_2994 (O_2994,N_29508,N_29877);
nor UO_2995 (O_2995,N_29498,N_29497);
xnor UO_2996 (O_2996,N_29400,N_29953);
or UO_2997 (O_2997,N_29913,N_29736);
or UO_2998 (O_2998,N_29466,N_29423);
and UO_2999 (O_2999,N_29782,N_29459);
xnor UO_3000 (O_3000,N_29987,N_29611);
or UO_3001 (O_3001,N_29963,N_29400);
nor UO_3002 (O_3002,N_29725,N_29863);
and UO_3003 (O_3003,N_29489,N_29427);
or UO_3004 (O_3004,N_29425,N_29641);
and UO_3005 (O_3005,N_29785,N_29743);
and UO_3006 (O_3006,N_29674,N_29457);
nand UO_3007 (O_3007,N_29874,N_29596);
nand UO_3008 (O_3008,N_29827,N_29862);
nor UO_3009 (O_3009,N_29863,N_29654);
and UO_3010 (O_3010,N_29876,N_29611);
and UO_3011 (O_3011,N_29973,N_29681);
nand UO_3012 (O_3012,N_29416,N_29880);
nor UO_3013 (O_3013,N_29788,N_29592);
and UO_3014 (O_3014,N_29689,N_29920);
xnor UO_3015 (O_3015,N_29762,N_29889);
xor UO_3016 (O_3016,N_29659,N_29914);
and UO_3017 (O_3017,N_29767,N_29636);
and UO_3018 (O_3018,N_29928,N_29981);
nand UO_3019 (O_3019,N_29611,N_29519);
or UO_3020 (O_3020,N_29757,N_29775);
or UO_3021 (O_3021,N_29558,N_29612);
and UO_3022 (O_3022,N_29860,N_29420);
nor UO_3023 (O_3023,N_29446,N_29776);
nor UO_3024 (O_3024,N_29839,N_29926);
nor UO_3025 (O_3025,N_29839,N_29900);
nor UO_3026 (O_3026,N_29481,N_29860);
or UO_3027 (O_3027,N_29777,N_29797);
nand UO_3028 (O_3028,N_29918,N_29872);
or UO_3029 (O_3029,N_29709,N_29772);
xor UO_3030 (O_3030,N_29774,N_29835);
xnor UO_3031 (O_3031,N_29755,N_29420);
and UO_3032 (O_3032,N_29852,N_29589);
or UO_3033 (O_3033,N_29401,N_29873);
xnor UO_3034 (O_3034,N_29831,N_29638);
xnor UO_3035 (O_3035,N_29490,N_29514);
and UO_3036 (O_3036,N_29555,N_29845);
nor UO_3037 (O_3037,N_29939,N_29480);
or UO_3038 (O_3038,N_29522,N_29834);
nand UO_3039 (O_3039,N_29427,N_29847);
or UO_3040 (O_3040,N_29631,N_29418);
xnor UO_3041 (O_3041,N_29797,N_29944);
nor UO_3042 (O_3042,N_29568,N_29615);
xor UO_3043 (O_3043,N_29475,N_29402);
and UO_3044 (O_3044,N_29895,N_29613);
xor UO_3045 (O_3045,N_29814,N_29742);
and UO_3046 (O_3046,N_29897,N_29946);
nand UO_3047 (O_3047,N_29879,N_29986);
nor UO_3048 (O_3048,N_29708,N_29785);
xor UO_3049 (O_3049,N_29791,N_29622);
xor UO_3050 (O_3050,N_29655,N_29959);
or UO_3051 (O_3051,N_29547,N_29787);
or UO_3052 (O_3052,N_29872,N_29835);
or UO_3053 (O_3053,N_29492,N_29838);
nand UO_3054 (O_3054,N_29926,N_29898);
nor UO_3055 (O_3055,N_29848,N_29824);
and UO_3056 (O_3056,N_29927,N_29797);
and UO_3057 (O_3057,N_29934,N_29682);
xor UO_3058 (O_3058,N_29755,N_29865);
and UO_3059 (O_3059,N_29684,N_29650);
and UO_3060 (O_3060,N_29893,N_29842);
nor UO_3061 (O_3061,N_29690,N_29657);
nor UO_3062 (O_3062,N_29530,N_29595);
xor UO_3063 (O_3063,N_29944,N_29935);
nor UO_3064 (O_3064,N_29416,N_29768);
or UO_3065 (O_3065,N_29871,N_29459);
nor UO_3066 (O_3066,N_29996,N_29764);
nor UO_3067 (O_3067,N_29774,N_29909);
and UO_3068 (O_3068,N_29780,N_29570);
nand UO_3069 (O_3069,N_29479,N_29711);
and UO_3070 (O_3070,N_29465,N_29581);
xor UO_3071 (O_3071,N_29617,N_29920);
xor UO_3072 (O_3072,N_29962,N_29912);
or UO_3073 (O_3073,N_29862,N_29797);
xor UO_3074 (O_3074,N_29509,N_29626);
xor UO_3075 (O_3075,N_29739,N_29459);
nor UO_3076 (O_3076,N_29978,N_29941);
nor UO_3077 (O_3077,N_29842,N_29711);
or UO_3078 (O_3078,N_29665,N_29493);
xnor UO_3079 (O_3079,N_29623,N_29843);
xor UO_3080 (O_3080,N_29867,N_29877);
and UO_3081 (O_3081,N_29865,N_29915);
and UO_3082 (O_3082,N_29632,N_29959);
nor UO_3083 (O_3083,N_29840,N_29569);
nor UO_3084 (O_3084,N_29968,N_29527);
or UO_3085 (O_3085,N_29463,N_29509);
nand UO_3086 (O_3086,N_29779,N_29553);
and UO_3087 (O_3087,N_29627,N_29406);
and UO_3088 (O_3088,N_29830,N_29448);
and UO_3089 (O_3089,N_29883,N_29869);
or UO_3090 (O_3090,N_29434,N_29494);
nand UO_3091 (O_3091,N_29637,N_29419);
nor UO_3092 (O_3092,N_29602,N_29692);
nand UO_3093 (O_3093,N_29512,N_29706);
nand UO_3094 (O_3094,N_29980,N_29420);
xnor UO_3095 (O_3095,N_29624,N_29655);
nor UO_3096 (O_3096,N_29852,N_29962);
and UO_3097 (O_3097,N_29608,N_29449);
and UO_3098 (O_3098,N_29646,N_29616);
xnor UO_3099 (O_3099,N_29900,N_29641);
xnor UO_3100 (O_3100,N_29585,N_29531);
nand UO_3101 (O_3101,N_29848,N_29745);
xnor UO_3102 (O_3102,N_29591,N_29538);
or UO_3103 (O_3103,N_29964,N_29617);
nor UO_3104 (O_3104,N_29936,N_29434);
xor UO_3105 (O_3105,N_29718,N_29777);
or UO_3106 (O_3106,N_29980,N_29938);
nand UO_3107 (O_3107,N_29909,N_29431);
and UO_3108 (O_3108,N_29852,N_29791);
and UO_3109 (O_3109,N_29514,N_29517);
xnor UO_3110 (O_3110,N_29914,N_29936);
or UO_3111 (O_3111,N_29710,N_29586);
xnor UO_3112 (O_3112,N_29827,N_29849);
nor UO_3113 (O_3113,N_29417,N_29792);
nor UO_3114 (O_3114,N_29825,N_29400);
xor UO_3115 (O_3115,N_29401,N_29571);
nor UO_3116 (O_3116,N_29415,N_29693);
nand UO_3117 (O_3117,N_29720,N_29552);
nand UO_3118 (O_3118,N_29474,N_29506);
or UO_3119 (O_3119,N_29815,N_29596);
or UO_3120 (O_3120,N_29415,N_29482);
or UO_3121 (O_3121,N_29450,N_29909);
nor UO_3122 (O_3122,N_29641,N_29489);
or UO_3123 (O_3123,N_29857,N_29669);
and UO_3124 (O_3124,N_29908,N_29727);
xnor UO_3125 (O_3125,N_29519,N_29415);
or UO_3126 (O_3126,N_29585,N_29473);
or UO_3127 (O_3127,N_29575,N_29497);
and UO_3128 (O_3128,N_29700,N_29823);
and UO_3129 (O_3129,N_29706,N_29709);
xnor UO_3130 (O_3130,N_29670,N_29765);
nand UO_3131 (O_3131,N_29441,N_29967);
and UO_3132 (O_3132,N_29685,N_29747);
nand UO_3133 (O_3133,N_29456,N_29521);
nand UO_3134 (O_3134,N_29547,N_29701);
and UO_3135 (O_3135,N_29554,N_29779);
or UO_3136 (O_3136,N_29706,N_29472);
nor UO_3137 (O_3137,N_29997,N_29845);
nand UO_3138 (O_3138,N_29547,N_29544);
xor UO_3139 (O_3139,N_29941,N_29976);
or UO_3140 (O_3140,N_29566,N_29889);
or UO_3141 (O_3141,N_29515,N_29751);
and UO_3142 (O_3142,N_29516,N_29405);
and UO_3143 (O_3143,N_29663,N_29871);
and UO_3144 (O_3144,N_29419,N_29723);
and UO_3145 (O_3145,N_29521,N_29962);
nand UO_3146 (O_3146,N_29810,N_29827);
nor UO_3147 (O_3147,N_29922,N_29930);
nand UO_3148 (O_3148,N_29456,N_29518);
or UO_3149 (O_3149,N_29540,N_29409);
or UO_3150 (O_3150,N_29604,N_29931);
xnor UO_3151 (O_3151,N_29904,N_29833);
nor UO_3152 (O_3152,N_29984,N_29679);
nand UO_3153 (O_3153,N_29730,N_29710);
and UO_3154 (O_3154,N_29468,N_29407);
nor UO_3155 (O_3155,N_29690,N_29930);
xnor UO_3156 (O_3156,N_29835,N_29699);
xor UO_3157 (O_3157,N_29583,N_29798);
xnor UO_3158 (O_3158,N_29527,N_29600);
and UO_3159 (O_3159,N_29651,N_29752);
nor UO_3160 (O_3160,N_29436,N_29863);
nor UO_3161 (O_3161,N_29810,N_29842);
and UO_3162 (O_3162,N_29913,N_29984);
nor UO_3163 (O_3163,N_29437,N_29863);
nand UO_3164 (O_3164,N_29873,N_29966);
nor UO_3165 (O_3165,N_29598,N_29820);
nand UO_3166 (O_3166,N_29724,N_29484);
xnor UO_3167 (O_3167,N_29440,N_29778);
xor UO_3168 (O_3168,N_29689,N_29790);
nand UO_3169 (O_3169,N_29502,N_29534);
nor UO_3170 (O_3170,N_29905,N_29693);
nand UO_3171 (O_3171,N_29847,N_29573);
xor UO_3172 (O_3172,N_29604,N_29400);
nand UO_3173 (O_3173,N_29722,N_29411);
nor UO_3174 (O_3174,N_29552,N_29596);
nand UO_3175 (O_3175,N_29703,N_29939);
nor UO_3176 (O_3176,N_29735,N_29451);
nor UO_3177 (O_3177,N_29424,N_29444);
nand UO_3178 (O_3178,N_29854,N_29725);
or UO_3179 (O_3179,N_29597,N_29545);
xnor UO_3180 (O_3180,N_29630,N_29441);
nand UO_3181 (O_3181,N_29872,N_29801);
nand UO_3182 (O_3182,N_29781,N_29429);
and UO_3183 (O_3183,N_29808,N_29961);
xor UO_3184 (O_3184,N_29964,N_29424);
or UO_3185 (O_3185,N_29594,N_29984);
xnor UO_3186 (O_3186,N_29788,N_29657);
nand UO_3187 (O_3187,N_29835,N_29461);
nor UO_3188 (O_3188,N_29567,N_29477);
xnor UO_3189 (O_3189,N_29799,N_29505);
and UO_3190 (O_3190,N_29671,N_29843);
or UO_3191 (O_3191,N_29840,N_29680);
nand UO_3192 (O_3192,N_29491,N_29456);
nand UO_3193 (O_3193,N_29970,N_29840);
and UO_3194 (O_3194,N_29460,N_29718);
and UO_3195 (O_3195,N_29728,N_29552);
nor UO_3196 (O_3196,N_29703,N_29812);
xnor UO_3197 (O_3197,N_29988,N_29725);
and UO_3198 (O_3198,N_29762,N_29993);
and UO_3199 (O_3199,N_29758,N_29909);
nor UO_3200 (O_3200,N_29890,N_29728);
xnor UO_3201 (O_3201,N_29499,N_29729);
or UO_3202 (O_3202,N_29550,N_29946);
and UO_3203 (O_3203,N_29812,N_29750);
or UO_3204 (O_3204,N_29494,N_29686);
nand UO_3205 (O_3205,N_29638,N_29912);
nor UO_3206 (O_3206,N_29842,N_29631);
nand UO_3207 (O_3207,N_29612,N_29471);
xor UO_3208 (O_3208,N_29721,N_29497);
or UO_3209 (O_3209,N_29482,N_29551);
xor UO_3210 (O_3210,N_29669,N_29449);
xor UO_3211 (O_3211,N_29493,N_29992);
and UO_3212 (O_3212,N_29873,N_29862);
or UO_3213 (O_3213,N_29838,N_29661);
xnor UO_3214 (O_3214,N_29760,N_29520);
nand UO_3215 (O_3215,N_29708,N_29700);
and UO_3216 (O_3216,N_29790,N_29552);
nand UO_3217 (O_3217,N_29969,N_29987);
nand UO_3218 (O_3218,N_29752,N_29510);
xnor UO_3219 (O_3219,N_29869,N_29892);
nor UO_3220 (O_3220,N_29593,N_29741);
nor UO_3221 (O_3221,N_29586,N_29448);
and UO_3222 (O_3222,N_29877,N_29857);
or UO_3223 (O_3223,N_29748,N_29709);
nor UO_3224 (O_3224,N_29451,N_29701);
nand UO_3225 (O_3225,N_29745,N_29917);
or UO_3226 (O_3226,N_29811,N_29798);
or UO_3227 (O_3227,N_29910,N_29974);
or UO_3228 (O_3228,N_29852,N_29474);
xnor UO_3229 (O_3229,N_29474,N_29692);
xor UO_3230 (O_3230,N_29683,N_29491);
nand UO_3231 (O_3231,N_29476,N_29626);
nor UO_3232 (O_3232,N_29894,N_29846);
xnor UO_3233 (O_3233,N_29406,N_29581);
or UO_3234 (O_3234,N_29823,N_29876);
nand UO_3235 (O_3235,N_29472,N_29893);
or UO_3236 (O_3236,N_29810,N_29515);
and UO_3237 (O_3237,N_29991,N_29676);
nor UO_3238 (O_3238,N_29629,N_29452);
nand UO_3239 (O_3239,N_29916,N_29891);
nor UO_3240 (O_3240,N_29845,N_29540);
nor UO_3241 (O_3241,N_29610,N_29709);
and UO_3242 (O_3242,N_29486,N_29545);
nand UO_3243 (O_3243,N_29650,N_29754);
nand UO_3244 (O_3244,N_29741,N_29839);
nor UO_3245 (O_3245,N_29580,N_29712);
nand UO_3246 (O_3246,N_29576,N_29482);
xor UO_3247 (O_3247,N_29977,N_29475);
or UO_3248 (O_3248,N_29452,N_29972);
and UO_3249 (O_3249,N_29865,N_29664);
and UO_3250 (O_3250,N_29613,N_29634);
nand UO_3251 (O_3251,N_29419,N_29444);
xor UO_3252 (O_3252,N_29556,N_29649);
and UO_3253 (O_3253,N_29422,N_29905);
nor UO_3254 (O_3254,N_29571,N_29577);
and UO_3255 (O_3255,N_29687,N_29765);
nor UO_3256 (O_3256,N_29929,N_29976);
xor UO_3257 (O_3257,N_29617,N_29777);
nor UO_3258 (O_3258,N_29884,N_29632);
nand UO_3259 (O_3259,N_29769,N_29561);
or UO_3260 (O_3260,N_29964,N_29554);
xor UO_3261 (O_3261,N_29970,N_29428);
nand UO_3262 (O_3262,N_29861,N_29597);
xnor UO_3263 (O_3263,N_29451,N_29808);
xnor UO_3264 (O_3264,N_29403,N_29938);
or UO_3265 (O_3265,N_29580,N_29772);
and UO_3266 (O_3266,N_29486,N_29665);
xor UO_3267 (O_3267,N_29508,N_29617);
or UO_3268 (O_3268,N_29764,N_29518);
xor UO_3269 (O_3269,N_29869,N_29648);
or UO_3270 (O_3270,N_29867,N_29914);
nor UO_3271 (O_3271,N_29407,N_29477);
or UO_3272 (O_3272,N_29627,N_29508);
nor UO_3273 (O_3273,N_29988,N_29671);
nor UO_3274 (O_3274,N_29644,N_29812);
or UO_3275 (O_3275,N_29949,N_29662);
and UO_3276 (O_3276,N_29763,N_29662);
nor UO_3277 (O_3277,N_29510,N_29989);
nor UO_3278 (O_3278,N_29541,N_29612);
and UO_3279 (O_3279,N_29552,N_29545);
xnor UO_3280 (O_3280,N_29994,N_29570);
or UO_3281 (O_3281,N_29856,N_29883);
nor UO_3282 (O_3282,N_29933,N_29814);
nand UO_3283 (O_3283,N_29997,N_29812);
xnor UO_3284 (O_3284,N_29727,N_29706);
and UO_3285 (O_3285,N_29809,N_29849);
and UO_3286 (O_3286,N_29603,N_29984);
or UO_3287 (O_3287,N_29721,N_29963);
xor UO_3288 (O_3288,N_29475,N_29830);
xor UO_3289 (O_3289,N_29683,N_29534);
nand UO_3290 (O_3290,N_29441,N_29488);
nor UO_3291 (O_3291,N_29995,N_29912);
nor UO_3292 (O_3292,N_29881,N_29919);
xnor UO_3293 (O_3293,N_29955,N_29812);
nor UO_3294 (O_3294,N_29700,N_29713);
xor UO_3295 (O_3295,N_29890,N_29606);
and UO_3296 (O_3296,N_29943,N_29421);
and UO_3297 (O_3297,N_29490,N_29923);
and UO_3298 (O_3298,N_29727,N_29662);
or UO_3299 (O_3299,N_29772,N_29794);
and UO_3300 (O_3300,N_29724,N_29708);
and UO_3301 (O_3301,N_29955,N_29765);
or UO_3302 (O_3302,N_29679,N_29540);
xnor UO_3303 (O_3303,N_29556,N_29557);
nand UO_3304 (O_3304,N_29814,N_29997);
nand UO_3305 (O_3305,N_29468,N_29861);
nand UO_3306 (O_3306,N_29672,N_29631);
xor UO_3307 (O_3307,N_29586,N_29643);
and UO_3308 (O_3308,N_29623,N_29982);
nand UO_3309 (O_3309,N_29737,N_29723);
nor UO_3310 (O_3310,N_29877,N_29995);
or UO_3311 (O_3311,N_29977,N_29791);
xor UO_3312 (O_3312,N_29415,N_29733);
nand UO_3313 (O_3313,N_29643,N_29466);
and UO_3314 (O_3314,N_29656,N_29444);
or UO_3315 (O_3315,N_29704,N_29452);
and UO_3316 (O_3316,N_29979,N_29805);
nor UO_3317 (O_3317,N_29831,N_29857);
xor UO_3318 (O_3318,N_29904,N_29952);
xor UO_3319 (O_3319,N_29572,N_29531);
xor UO_3320 (O_3320,N_29412,N_29550);
xnor UO_3321 (O_3321,N_29470,N_29799);
nand UO_3322 (O_3322,N_29417,N_29577);
nand UO_3323 (O_3323,N_29541,N_29568);
or UO_3324 (O_3324,N_29657,N_29759);
and UO_3325 (O_3325,N_29856,N_29770);
xor UO_3326 (O_3326,N_29815,N_29430);
nand UO_3327 (O_3327,N_29681,N_29836);
nand UO_3328 (O_3328,N_29986,N_29992);
or UO_3329 (O_3329,N_29479,N_29860);
or UO_3330 (O_3330,N_29946,N_29446);
xor UO_3331 (O_3331,N_29916,N_29497);
nand UO_3332 (O_3332,N_29652,N_29898);
or UO_3333 (O_3333,N_29580,N_29957);
nand UO_3334 (O_3334,N_29683,N_29945);
or UO_3335 (O_3335,N_29586,N_29900);
xnor UO_3336 (O_3336,N_29953,N_29464);
or UO_3337 (O_3337,N_29825,N_29660);
nor UO_3338 (O_3338,N_29693,N_29448);
nand UO_3339 (O_3339,N_29790,N_29794);
or UO_3340 (O_3340,N_29524,N_29612);
nand UO_3341 (O_3341,N_29669,N_29695);
xor UO_3342 (O_3342,N_29721,N_29429);
xnor UO_3343 (O_3343,N_29491,N_29552);
nand UO_3344 (O_3344,N_29549,N_29765);
nor UO_3345 (O_3345,N_29609,N_29746);
or UO_3346 (O_3346,N_29671,N_29633);
nor UO_3347 (O_3347,N_29706,N_29800);
or UO_3348 (O_3348,N_29722,N_29719);
and UO_3349 (O_3349,N_29849,N_29856);
xnor UO_3350 (O_3350,N_29744,N_29868);
or UO_3351 (O_3351,N_29523,N_29884);
xor UO_3352 (O_3352,N_29424,N_29751);
nor UO_3353 (O_3353,N_29568,N_29656);
nand UO_3354 (O_3354,N_29511,N_29539);
or UO_3355 (O_3355,N_29633,N_29951);
nor UO_3356 (O_3356,N_29422,N_29766);
and UO_3357 (O_3357,N_29559,N_29529);
xnor UO_3358 (O_3358,N_29518,N_29908);
nand UO_3359 (O_3359,N_29939,N_29785);
nor UO_3360 (O_3360,N_29682,N_29941);
nand UO_3361 (O_3361,N_29680,N_29934);
nand UO_3362 (O_3362,N_29956,N_29863);
and UO_3363 (O_3363,N_29560,N_29728);
xor UO_3364 (O_3364,N_29541,N_29649);
or UO_3365 (O_3365,N_29739,N_29688);
nand UO_3366 (O_3366,N_29429,N_29567);
xnor UO_3367 (O_3367,N_29578,N_29951);
and UO_3368 (O_3368,N_29838,N_29880);
and UO_3369 (O_3369,N_29532,N_29895);
nand UO_3370 (O_3370,N_29983,N_29428);
or UO_3371 (O_3371,N_29601,N_29634);
nand UO_3372 (O_3372,N_29400,N_29544);
nand UO_3373 (O_3373,N_29481,N_29796);
xnor UO_3374 (O_3374,N_29916,N_29540);
and UO_3375 (O_3375,N_29470,N_29732);
nor UO_3376 (O_3376,N_29688,N_29869);
nor UO_3377 (O_3377,N_29836,N_29552);
nor UO_3378 (O_3378,N_29759,N_29893);
nor UO_3379 (O_3379,N_29683,N_29456);
or UO_3380 (O_3380,N_29655,N_29853);
or UO_3381 (O_3381,N_29461,N_29560);
nand UO_3382 (O_3382,N_29892,N_29697);
and UO_3383 (O_3383,N_29488,N_29601);
or UO_3384 (O_3384,N_29409,N_29437);
xor UO_3385 (O_3385,N_29550,N_29449);
or UO_3386 (O_3386,N_29412,N_29434);
nor UO_3387 (O_3387,N_29627,N_29703);
nor UO_3388 (O_3388,N_29503,N_29580);
or UO_3389 (O_3389,N_29905,N_29988);
and UO_3390 (O_3390,N_29661,N_29979);
and UO_3391 (O_3391,N_29983,N_29776);
xor UO_3392 (O_3392,N_29464,N_29848);
xnor UO_3393 (O_3393,N_29622,N_29424);
xnor UO_3394 (O_3394,N_29587,N_29466);
nand UO_3395 (O_3395,N_29953,N_29661);
or UO_3396 (O_3396,N_29518,N_29675);
nor UO_3397 (O_3397,N_29512,N_29454);
or UO_3398 (O_3398,N_29741,N_29659);
nor UO_3399 (O_3399,N_29775,N_29736);
nand UO_3400 (O_3400,N_29997,N_29558);
nor UO_3401 (O_3401,N_29440,N_29971);
nor UO_3402 (O_3402,N_29484,N_29605);
and UO_3403 (O_3403,N_29656,N_29927);
xnor UO_3404 (O_3404,N_29904,N_29832);
or UO_3405 (O_3405,N_29887,N_29918);
and UO_3406 (O_3406,N_29939,N_29488);
nand UO_3407 (O_3407,N_29712,N_29713);
and UO_3408 (O_3408,N_29641,N_29847);
and UO_3409 (O_3409,N_29431,N_29978);
nand UO_3410 (O_3410,N_29720,N_29944);
or UO_3411 (O_3411,N_29682,N_29532);
nand UO_3412 (O_3412,N_29638,N_29684);
or UO_3413 (O_3413,N_29872,N_29584);
xnor UO_3414 (O_3414,N_29848,N_29481);
xnor UO_3415 (O_3415,N_29490,N_29614);
nor UO_3416 (O_3416,N_29423,N_29419);
xor UO_3417 (O_3417,N_29884,N_29861);
or UO_3418 (O_3418,N_29420,N_29443);
and UO_3419 (O_3419,N_29853,N_29408);
nor UO_3420 (O_3420,N_29608,N_29514);
and UO_3421 (O_3421,N_29640,N_29407);
and UO_3422 (O_3422,N_29897,N_29587);
and UO_3423 (O_3423,N_29415,N_29670);
xor UO_3424 (O_3424,N_29664,N_29617);
nand UO_3425 (O_3425,N_29702,N_29764);
and UO_3426 (O_3426,N_29774,N_29646);
xor UO_3427 (O_3427,N_29631,N_29857);
or UO_3428 (O_3428,N_29858,N_29576);
or UO_3429 (O_3429,N_29954,N_29465);
nand UO_3430 (O_3430,N_29662,N_29746);
nand UO_3431 (O_3431,N_29938,N_29717);
and UO_3432 (O_3432,N_29651,N_29456);
and UO_3433 (O_3433,N_29486,N_29632);
xor UO_3434 (O_3434,N_29576,N_29982);
or UO_3435 (O_3435,N_29790,N_29898);
and UO_3436 (O_3436,N_29463,N_29558);
nand UO_3437 (O_3437,N_29633,N_29569);
or UO_3438 (O_3438,N_29520,N_29862);
nand UO_3439 (O_3439,N_29628,N_29765);
or UO_3440 (O_3440,N_29528,N_29756);
xor UO_3441 (O_3441,N_29993,N_29526);
and UO_3442 (O_3442,N_29611,N_29598);
and UO_3443 (O_3443,N_29823,N_29497);
xnor UO_3444 (O_3444,N_29881,N_29980);
nand UO_3445 (O_3445,N_29757,N_29678);
nor UO_3446 (O_3446,N_29533,N_29981);
nand UO_3447 (O_3447,N_29707,N_29652);
xor UO_3448 (O_3448,N_29940,N_29707);
xnor UO_3449 (O_3449,N_29608,N_29654);
and UO_3450 (O_3450,N_29591,N_29434);
nand UO_3451 (O_3451,N_29562,N_29626);
xnor UO_3452 (O_3452,N_29784,N_29836);
nor UO_3453 (O_3453,N_29733,N_29978);
or UO_3454 (O_3454,N_29856,N_29985);
nor UO_3455 (O_3455,N_29868,N_29552);
nand UO_3456 (O_3456,N_29885,N_29693);
xor UO_3457 (O_3457,N_29613,N_29788);
or UO_3458 (O_3458,N_29438,N_29442);
nor UO_3459 (O_3459,N_29827,N_29747);
and UO_3460 (O_3460,N_29970,N_29581);
and UO_3461 (O_3461,N_29685,N_29527);
and UO_3462 (O_3462,N_29946,N_29935);
or UO_3463 (O_3463,N_29990,N_29751);
and UO_3464 (O_3464,N_29413,N_29940);
xnor UO_3465 (O_3465,N_29970,N_29868);
nand UO_3466 (O_3466,N_29655,N_29991);
or UO_3467 (O_3467,N_29884,N_29724);
nand UO_3468 (O_3468,N_29533,N_29948);
xnor UO_3469 (O_3469,N_29628,N_29502);
and UO_3470 (O_3470,N_29913,N_29959);
and UO_3471 (O_3471,N_29754,N_29807);
nor UO_3472 (O_3472,N_29881,N_29479);
nand UO_3473 (O_3473,N_29915,N_29578);
nand UO_3474 (O_3474,N_29601,N_29695);
and UO_3475 (O_3475,N_29704,N_29620);
or UO_3476 (O_3476,N_29536,N_29456);
xnor UO_3477 (O_3477,N_29417,N_29618);
nor UO_3478 (O_3478,N_29908,N_29706);
or UO_3479 (O_3479,N_29598,N_29898);
or UO_3480 (O_3480,N_29460,N_29465);
nand UO_3481 (O_3481,N_29479,N_29894);
or UO_3482 (O_3482,N_29891,N_29910);
or UO_3483 (O_3483,N_29567,N_29967);
nand UO_3484 (O_3484,N_29919,N_29541);
xor UO_3485 (O_3485,N_29644,N_29958);
nor UO_3486 (O_3486,N_29407,N_29782);
nand UO_3487 (O_3487,N_29604,N_29508);
or UO_3488 (O_3488,N_29624,N_29402);
nor UO_3489 (O_3489,N_29477,N_29959);
or UO_3490 (O_3490,N_29823,N_29407);
or UO_3491 (O_3491,N_29573,N_29684);
and UO_3492 (O_3492,N_29978,N_29980);
xor UO_3493 (O_3493,N_29672,N_29983);
nor UO_3494 (O_3494,N_29974,N_29997);
nor UO_3495 (O_3495,N_29627,N_29585);
xnor UO_3496 (O_3496,N_29468,N_29644);
nor UO_3497 (O_3497,N_29851,N_29493);
and UO_3498 (O_3498,N_29808,N_29677);
or UO_3499 (O_3499,N_29636,N_29989);
endmodule