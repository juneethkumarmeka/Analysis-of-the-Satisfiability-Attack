module basic_750_5000_1000_2_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2501,N_2502,N_2503,N_2504,N_2505,N_2508,N_2513,N_2514,N_2515,N_2516,N_2518,N_2519,N_2520,N_2521,N_2522,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2533,N_2534,N_2535,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2545,N_2547,N_2548,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2573,N_2575,N_2576,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2586,N_2587,N_2588,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2598,N_2600,N_2601,N_2602,N_2603,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2616,N_2619,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2663,N_2664,N_2665,N_2666,N_2668,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2726,N_2727,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2748,N_2749,N_2750,N_2751,N_2752,N_2754,N_2756,N_2759,N_2760,N_2761,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2775,N_2779,N_2780,N_2782,N_2783,N_2784,N_2788,N_2789,N_2790,N_2791,N_2792,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2802,N_2803,N_2806,N_2807,N_2809,N_2810,N_2811,N_2812,N_2813,N_2815,N_2817,N_2819,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2832,N_2833,N_2834,N_2837,N_2838,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2848,N_2849,N_2850,N_2852,N_2855,N_2856,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2867,N_2868,N_2870,N_2871,N_2872,N_2873,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2883,N_2884,N_2885,N_2886,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2915,N_2916,N_2917,N_2919,N_2920,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2943,N_2944,N_2945,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2980,N_2983,N_2984,N_2987,N_2988,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3008,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3054,N_3057,N_3058,N_3061,N_3062,N_3064,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3075,N_3076,N_3077,N_3079,N_3081,N_3082,N_3083,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3092,N_3094,N_3096,N_3097,N_3100,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3109,N_3111,N_3113,N_3114,N_3115,N_3116,N_3118,N_3119,N_3121,N_3122,N_3123,N_3124,N_3126,N_3128,N_3129,N_3130,N_3131,N_3132,N_3134,N_3136,N_3138,N_3139,N_3141,N_3142,N_3143,N_3148,N_3151,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3163,N_3164,N_3165,N_3167,N_3169,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3197,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3250,N_3251,N_3252,N_3254,N_3255,N_3256,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3274,N_3275,N_3276,N_3277,N_3278,N_3280,N_3281,N_3282,N_3283,N_3285,N_3286,N_3289,N_3290,N_3291,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3302,N_3303,N_3304,N_3308,N_3309,N_3310,N_3311,N_3312,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3323,N_3325,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3339,N_3341,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3351,N_3352,N_3353,N_3354,N_3356,N_3357,N_3358,N_3360,N_3361,N_3362,N_3364,N_3366,N_3368,N_3369,N_3370,N_3371,N_3372,N_3374,N_3376,N_3377,N_3378,N_3380,N_3381,N_3382,N_3383,N_3384,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3393,N_3394,N_3395,N_3396,N_3397,N_3399,N_3400,N_3401,N_3402,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3411,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3421,N_3422,N_3424,N_3426,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3448,N_3450,N_3451,N_3454,N_3455,N_3456,N_3457,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3485,N_3486,N_3487,N_3488,N_3489,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3506,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3542,N_3543,N_3547,N_3550,N_3552,N_3553,N_3554,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3568,N_3569,N_3571,N_3572,N_3573,N_3575,N_3576,N_3577,N_3578,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3589,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3613,N_3614,N_3615,N_3616,N_3618,N_3621,N_3622,N_3624,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3634,N_3635,N_3636,N_3639,N_3640,N_3642,N_3643,N_3644,N_3645,N_3647,N_3648,N_3649,N_3650,N_3651,N_3653,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3665,N_3666,N_3668,N_3669,N_3671,N_3672,N_3674,N_3675,N_3676,N_3677,N_3678,N_3680,N_3681,N_3682,N_3685,N_3687,N_3689,N_3691,N_3692,N_3693,N_3694,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3718,N_3719,N_3720,N_3721,N_3722,N_3724,N_3725,N_3726,N_3729,N_3730,N_3731,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3758,N_3759,N_3760,N_3761,N_3762,N_3764,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3785,N_3787,N_3788,N_3789,N_3790,N_3791,N_3793,N_3794,N_3795,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3804,N_3806,N_3807,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3818,N_3819,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3830,N_3831,N_3832,N_3834,N_3835,N_3837,N_3838,N_3839,N_3840,N_3843,N_3844,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3856,N_3857,N_3860,N_3861,N_3862,N_3864,N_3865,N_3866,N_3868,N_3869,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3878,N_3879,N_3880,N_3881,N_3883,N_3886,N_3887,N_3888,N_3891,N_3892,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3952,N_3954,N_3955,N_3956,N_3958,N_3959,N_3960,N_3961,N_3962,N_3964,N_3965,N_3966,N_3967,N_3968,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_4000,N_4001,N_4002,N_4003,N_4004,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4016,N_4017,N_4018,N_4019,N_4020,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4030,N_4031,N_4032,N_4033,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4056,N_4057,N_4059,N_4062,N_4063,N_4064,N_4065,N_4067,N_4069,N_4071,N_4072,N_4073,N_4074,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4091,N_4093,N_4095,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4137,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4154,N_4155,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4167,N_4168,N_4169,N_4171,N_4172,N_4173,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4200,N_4201,N_4202,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4216,N_4218,N_4219,N_4220,N_4222,N_4223,N_4224,N_4225,N_4227,N_4228,N_4230,N_4231,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4240,N_4241,N_4242,N_4243,N_4245,N_4246,N_4247,N_4248,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4258,N_4259,N_4260,N_4262,N_4263,N_4264,N_4265,N_4266,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4289,N_4291,N_4293,N_4294,N_4295,N_4297,N_4298,N_4300,N_4302,N_4303,N_4304,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4328,N_4330,N_4332,N_4336,N_4337,N_4338,N_4339,N_4340,N_4342,N_4343,N_4344,N_4346,N_4347,N_4348,N_4349,N_4351,N_4352,N_4353,N_4354,N_4355,N_4357,N_4358,N_4359,N_4361,N_4362,N_4364,N_4365,N_4366,N_4368,N_4369,N_4371,N_4372,N_4373,N_4374,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4383,N_4384,N_4385,N_4386,N_4389,N_4390,N_4391,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4464,N_4465,N_4466,N_4467,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4488,N_4489,N_4491,N_4493,N_4494,N_4495,N_4496,N_4497,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4507,N_4509,N_4511,N_4512,N_4513,N_4514,N_4516,N_4517,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4549,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4557,N_4558,N_4559,N_4561,N_4562,N_4563,N_4565,N_4566,N_4568,N_4569,N_4570,N_4572,N_4574,N_4575,N_4578,N_4579,N_4580,N_4581,N_4582,N_4584,N_4585,N_4586,N_4588,N_4590,N_4592,N_4593,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4603,N_4604,N_4605,N_4606,N_4607,N_4609,N_4610,N_4611,N_4613,N_4614,N_4615,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4659,N_4660,N_4661,N_4662,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4675,N_4676,N_4677,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4697,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4709,N_4710,N_4711,N_4712,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4724,N_4725,N_4726,N_4727,N_4729,N_4730,N_4731,N_4733,N_4734,N_4735,N_4736,N_4737,N_4739,N_4740,N_4741,N_4743,N_4744,N_4745,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4761,N_4762,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4777,N_4778,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4789,N_4790,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4801,N_4803,N_4804,N_4806,N_4807,N_4808,N_4809,N_4811,N_4814,N_4815,N_4816,N_4818,N_4819,N_4820,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4845,N_4846,N_4847,N_4849,N_4851,N_4853,N_4854,N_4855,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4892,N_4893,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4902,N_4903,N_4904,N_4905,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4922,N_4924,N_4925,N_4927,N_4928,N_4930,N_4931,N_4932,N_4933,N_4935,N_4936,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4946,N_4947,N_4948,N_4949,N_4951,N_4953,N_4954,N_4956,N_4957,N_4958,N_4959,N_4960,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4970,N_4971,N_4973,N_4974,N_4975,N_4976,N_4978,N_4980,N_4981,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_345,In_504);
nor U1 (N_1,In_638,In_224);
nor U2 (N_2,In_512,In_325);
nor U3 (N_3,In_651,In_195);
nor U4 (N_4,In_683,In_405);
or U5 (N_5,In_602,In_98);
or U6 (N_6,In_358,In_362);
nand U7 (N_7,In_181,In_377);
and U8 (N_8,In_334,In_408);
nand U9 (N_9,In_655,In_124);
nor U10 (N_10,In_149,In_446);
nor U11 (N_11,In_747,In_180);
nand U12 (N_12,In_511,In_129);
and U13 (N_13,In_383,In_508);
or U14 (N_14,In_617,In_62);
nor U15 (N_15,In_144,In_453);
nand U16 (N_16,In_242,In_163);
and U17 (N_17,In_419,In_733);
or U18 (N_18,In_344,In_313);
nand U19 (N_19,In_705,In_629);
nor U20 (N_20,In_35,In_145);
nor U21 (N_21,In_555,In_55);
nor U22 (N_22,In_454,In_713);
or U23 (N_23,In_670,In_645);
nor U24 (N_24,In_436,In_160);
nand U25 (N_25,In_142,In_317);
and U26 (N_26,In_697,In_351);
or U27 (N_27,In_54,In_710);
or U28 (N_28,In_201,In_521);
nor U29 (N_29,In_380,In_462);
or U30 (N_30,In_281,In_105);
nor U31 (N_31,In_3,In_140);
or U32 (N_32,In_122,In_654);
xnor U33 (N_33,In_126,In_104);
nand U34 (N_34,In_298,In_715);
and U35 (N_35,In_192,In_514);
nor U36 (N_36,In_13,In_736);
nand U37 (N_37,In_112,In_245);
nand U38 (N_38,In_559,In_694);
and U39 (N_39,In_726,In_593);
or U40 (N_40,In_553,In_650);
nand U41 (N_41,In_532,In_45);
nand U42 (N_42,In_47,In_416);
nor U43 (N_43,In_554,In_341);
or U44 (N_44,In_369,In_601);
and U45 (N_45,In_337,In_422);
nand U46 (N_46,In_718,In_328);
or U47 (N_47,In_674,In_169);
and U48 (N_48,In_734,In_262);
nand U49 (N_49,In_722,In_412);
or U50 (N_50,In_246,In_564);
nand U51 (N_51,In_95,In_33);
or U52 (N_52,In_266,In_20);
and U53 (N_53,In_202,In_572);
nand U54 (N_54,In_339,In_319);
nor U55 (N_55,In_65,In_477);
nor U56 (N_56,In_528,In_493);
nor U57 (N_57,In_85,In_481);
nor U58 (N_58,In_361,In_570);
xor U59 (N_59,In_647,In_23);
nand U60 (N_60,In_204,In_6);
xor U61 (N_61,In_631,In_165);
or U62 (N_62,In_205,In_237);
nor U63 (N_63,In_724,In_576);
nor U64 (N_64,In_367,In_107);
xor U65 (N_65,In_608,In_111);
nand U66 (N_66,In_61,In_322);
or U67 (N_67,In_355,In_60);
nor U68 (N_68,In_677,In_208);
or U69 (N_69,In_605,In_686);
xor U70 (N_70,In_250,In_233);
and U71 (N_71,In_652,In_745);
or U72 (N_72,In_379,In_5);
nand U73 (N_73,In_267,In_286);
xnor U74 (N_74,In_640,In_290);
nor U75 (N_75,In_539,In_110);
xor U76 (N_76,In_384,In_583);
and U77 (N_77,In_77,In_81);
nor U78 (N_78,In_143,In_644);
xnor U79 (N_79,In_627,In_82);
nand U80 (N_80,In_269,In_225);
or U81 (N_81,In_499,In_738);
nand U82 (N_82,In_546,In_372);
nor U83 (N_83,In_561,In_103);
nor U84 (N_84,In_100,In_155);
nor U85 (N_85,In_11,In_1);
and U86 (N_86,In_461,In_458);
and U87 (N_87,In_681,In_594);
or U88 (N_88,In_548,In_421);
nand U89 (N_89,In_15,In_146);
nand U90 (N_90,In_474,In_698);
nand U91 (N_91,In_311,In_413);
nor U92 (N_92,In_130,In_376);
and U93 (N_93,In_302,In_92);
nor U94 (N_94,In_136,In_513);
or U95 (N_95,In_125,In_99);
nor U96 (N_96,In_44,In_611);
nand U97 (N_97,In_531,In_116);
nand U98 (N_98,In_721,In_52);
nor U99 (N_99,In_121,In_428);
nor U100 (N_100,In_342,In_600);
nand U101 (N_101,In_26,In_392);
or U102 (N_102,In_218,In_324);
nand U103 (N_103,In_723,In_479);
nor U104 (N_104,In_491,In_212);
nand U105 (N_105,In_106,In_349);
nor U106 (N_106,In_42,In_354);
nand U107 (N_107,In_497,In_133);
nor U108 (N_108,In_673,In_614);
and U109 (N_109,In_312,In_487);
or U110 (N_110,In_565,In_279);
or U111 (N_111,In_375,In_308);
nand U112 (N_112,In_171,In_476);
or U113 (N_113,In_174,In_101);
nand U114 (N_114,In_265,In_53);
nor U115 (N_115,In_148,In_393);
nor U116 (N_116,In_524,In_310);
or U117 (N_117,In_475,In_727);
and U118 (N_118,In_333,In_340);
and U119 (N_119,In_50,In_271);
nor U120 (N_120,In_215,In_9);
and U121 (N_121,In_441,In_717);
nand U122 (N_122,In_543,In_223);
or U123 (N_123,In_578,In_626);
or U124 (N_124,In_582,In_556);
nand U125 (N_125,In_520,In_604);
or U126 (N_126,In_630,In_643);
nor U127 (N_127,In_691,In_127);
nor U128 (N_128,In_471,In_326);
nor U129 (N_129,In_57,In_459);
nor U130 (N_130,In_418,In_228);
nor U131 (N_131,In_283,In_294);
nand U132 (N_132,In_581,In_251);
or U133 (N_133,In_282,In_221);
nor U134 (N_134,In_327,In_131);
nand U135 (N_135,In_357,In_307);
nor U136 (N_136,In_526,In_501);
nor U137 (N_137,In_74,In_219);
nor U138 (N_138,In_449,In_712);
nand U139 (N_139,In_19,In_389);
or U140 (N_140,In_612,In_48);
and U141 (N_141,In_37,In_186);
or U142 (N_142,In_537,In_235);
xor U143 (N_143,In_658,In_735);
nor U144 (N_144,In_8,In_547);
nor U145 (N_145,In_278,In_275);
nand U146 (N_146,In_443,In_414);
nand U147 (N_147,In_634,In_482);
nor U148 (N_148,In_183,In_230);
or U149 (N_149,In_260,In_115);
nor U150 (N_150,In_447,In_177);
nand U151 (N_151,In_56,In_580);
nor U152 (N_152,In_226,In_741);
nor U153 (N_153,In_210,In_86);
and U154 (N_154,In_196,In_247);
nor U155 (N_155,In_530,In_444);
or U156 (N_156,In_467,In_305);
nor U157 (N_157,In_529,In_430);
nand U158 (N_158,In_607,In_296);
nor U159 (N_159,In_12,In_590);
or U160 (N_160,In_687,In_71);
nand U161 (N_161,In_536,In_280);
or U162 (N_162,In_17,In_696);
nand U163 (N_163,In_457,In_434);
nand U164 (N_164,In_360,In_69);
nor U165 (N_165,In_470,In_321);
or U166 (N_166,In_429,In_588);
or U167 (N_167,In_469,In_366);
or U168 (N_168,In_615,In_29);
nor U169 (N_169,In_185,In_199);
and U170 (N_170,In_541,In_109);
nor U171 (N_171,In_66,In_273);
nor U172 (N_172,In_18,In_663);
nand U173 (N_173,In_193,In_154);
and U174 (N_174,In_743,In_549);
and U175 (N_175,In_34,In_303);
nor U176 (N_176,In_287,In_374);
nand U177 (N_177,In_648,In_639);
or U178 (N_178,In_244,In_32);
nand U179 (N_179,In_503,In_272);
nor U180 (N_180,In_692,In_460);
nor U181 (N_181,In_359,In_138);
and U182 (N_182,In_299,In_455);
nor U183 (N_183,In_137,In_173);
nor U184 (N_184,In_49,In_252);
or U185 (N_185,In_402,In_188);
nand U186 (N_186,In_117,In_494);
and U187 (N_187,In_403,In_270);
or U188 (N_188,In_178,In_438);
and U189 (N_189,In_64,In_574);
nand U190 (N_190,In_706,In_519);
or U191 (N_191,In_30,In_141);
or U192 (N_192,In_320,In_399);
and U193 (N_193,In_584,In_288);
nor U194 (N_194,In_496,In_284);
nand U195 (N_195,In_240,In_113);
nand U196 (N_196,In_365,In_708);
and U197 (N_197,In_184,In_709);
nor U198 (N_198,In_197,In_159);
and U199 (N_199,In_350,In_685);
or U200 (N_200,In_68,In_216);
nor U201 (N_201,In_472,In_432);
nor U202 (N_202,In_675,In_41);
or U203 (N_203,In_268,In_119);
nor U204 (N_204,In_238,In_669);
and U205 (N_205,In_36,In_737);
nor U206 (N_206,In_387,In_78);
and U207 (N_207,In_410,In_297);
nor U208 (N_208,In_390,In_128);
nand U209 (N_209,In_488,In_448);
nand U210 (N_210,In_108,In_435);
nor U211 (N_211,In_231,In_417);
and U212 (N_212,In_39,In_175);
nand U213 (N_213,In_373,In_707);
nand U214 (N_214,In_211,In_442);
or U215 (N_215,In_450,In_209);
and U216 (N_216,In_484,In_649);
nand U217 (N_217,In_254,In_550);
nor U218 (N_218,In_610,In_385);
or U219 (N_219,In_426,In_76);
and U220 (N_220,In_22,In_415);
nor U221 (N_221,In_306,In_510);
nand U222 (N_222,In_263,In_59);
nor U223 (N_223,In_558,In_364);
xor U224 (N_224,In_404,In_207);
nand U225 (N_225,In_353,In_619);
and U226 (N_226,In_318,In_277);
or U227 (N_227,In_84,In_500);
and U228 (N_228,In_304,In_517);
nand U229 (N_229,In_335,In_606);
and U230 (N_230,In_382,In_540);
nor U231 (N_231,In_217,In_190);
nor U232 (N_232,In_167,In_182);
and U233 (N_233,In_628,In_682);
or U234 (N_234,In_292,In_609);
nor U235 (N_235,In_700,In_259);
nand U236 (N_236,In_70,In_660);
and U237 (N_237,In_731,In_506);
nand U238 (N_238,In_595,In_336);
nand U239 (N_239,In_485,In_329);
nor U240 (N_240,In_567,In_176);
or U241 (N_241,In_168,In_621);
and U242 (N_242,In_249,In_563);
or U243 (N_243,In_749,In_676);
and U244 (N_244,In_498,In_664);
nand U245 (N_245,In_4,In_388);
and U246 (N_246,In_147,In_28);
or U247 (N_247,In_439,In_229);
nor U248 (N_248,In_603,In_566);
and U249 (N_249,In_507,In_332);
nor U250 (N_250,In_613,In_2);
or U251 (N_251,In_732,In_352);
or U252 (N_252,In_347,In_586);
or U253 (N_253,In_693,In_25);
and U254 (N_254,In_623,In_94);
nor U255 (N_255,In_348,In_492);
nor U256 (N_256,In_592,In_88);
nor U257 (N_257,In_622,In_153);
nand U258 (N_258,In_678,In_552);
xor U259 (N_259,In_203,In_123);
nand U260 (N_260,In_515,In_338);
and U261 (N_261,In_24,In_679);
or U262 (N_262,In_585,In_478);
or U263 (N_263,In_14,In_680);
or U264 (N_264,In_719,In_10);
and U265 (N_265,In_409,In_659);
nand U266 (N_266,In_396,In_91);
or U267 (N_267,In_624,In_27);
nor U268 (N_268,In_527,In_97);
nand U269 (N_269,In_346,In_330);
nand U270 (N_270,In_716,In_538);
and U271 (N_271,In_533,In_579);
nand U272 (N_272,In_489,In_31);
or U273 (N_273,In_742,In_43);
nand U274 (N_274,In_411,In_495);
nor U275 (N_275,In_616,In_702);
or U276 (N_276,In_463,In_668);
nand U277 (N_277,In_689,In_542);
nor U278 (N_278,In_40,In_206);
or U279 (N_279,In_368,In_688);
and U280 (N_280,In_120,In_598);
or U281 (N_281,In_381,In_544);
xnor U282 (N_282,In_551,In_222);
or U283 (N_283,In_577,In_518);
nand U284 (N_284,In_391,In_96);
nand U285 (N_285,In_440,In_525);
nor U286 (N_286,In_378,In_398);
nor U287 (N_287,In_420,In_67);
nand U288 (N_288,In_452,In_672);
and U289 (N_289,In_89,In_83);
or U290 (N_290,In_739,In_456);
or U291 (N_291,In_740,In_425);
nand U292 (N_292,In_748,In_371);
and U293 (N_293,In_730,In_703);
nand U294 (N_294,In_363,In_468);
nor U295 (N_295,In_316,In_227);
or U296 (N_296,In_662,In_534);
nand U297 (N_297,In_483,In_72);
and U298 (N_298,In_172,In_473);
or U299 (N_299,In_690,In_191);
nand U300 (N_300,In_407,In_401);
nor U301 (N_301,In_241,In_632);
nand U302 (N_302,In_255,In_437);
and U303 (N_303,In_243,In_0);
nand U304 (N_304,In_486,In_400);
nor U305 (N_305,In_170,In_523);
nor U306 (N_306,In_464,In_502);
nand U307 (N_307,In_21,In_516);
or U308 (N_308,In_620,In_509);
nand U309 (N_309,In_433,In_46);
xnor U310 (N_310,In_665,In_699);
nand U311 (N_311,In_725,In_314);
or U312 (N_312,In_701,In_562);
nand U313 (N_313,In_597,In_568);
and U314 (N_314,In_16,In_466);
and U315 (N_315,In_38,In_51);
nor U316 (N_316,In_156,In_261);
or U317 (N_317,In_132,In_150);
nand U318 (N_318,In_200,In_744);
nand U319 (N_319,In_505,In_657);
nor U320 (N_320,In_587,In_625);
or U321 (N_321,In_194,In_162);
nand U322 (N_322,In_343,In_397);
or U323 (N_323,In_465,In_695);
or U324 (N_324,In_220,In_139);
or U325 (N_325,In_535,In_596);
nand U326 (N_326,In_164,In_656);
and U327 (N_327,In_118,In_285);
or U328 (N_328,In_490,In_560);
nor U329 (N_329,In_158,In_423);
nor U330 (N_330,In_161,In_522);
nor U331 (N_331,In_102,In_248);
nand U332 (N_332,In_395,In_79);
and U333 (N_333,In_309,In_264);
nor U334 (N_334,In_661,In_315);
nand U335 (N_335,In_90,In_642);
or U336 (N_336,In_720,In_545);
or U337 (N_337,In_666,In_667);
nor U338 (N_338,In_575,In_653);
nor U339 (N_339,In_569,In_214);
nor U340 (N_340,In_636,In_618);
nor U341 (N_341,In_276,In_274);
and U342 (N_342,In_684,In_134);
and U343 (N_343,In_711,In_571);
or U344 (N_344,In_671,In_189);
or U345 (N_345,In_394,In_187);
nor U346 (N_346,In_232,In_295);
or U347 (N_347,In_331,In_151);
or U348 (N_348,In_239,In_236);
nor U349 (N_349,In_406,In_63);
nor U350 (N_350,In_73,In_704);
nor U351 (N_351,In_256,In_135);
or U352 (N_352,In_641,In_152);
or U353 (N_353,In_480,In_637);
nor U354 (N_354,In_633,In_293);
or U355 (N_355,In_356,In_646);
or U356 (N_356,In_75,In_728);
or U357 (N_357,In_213,In_93);
or U358 (N_358,In_300,In_589);
nand U359 (N_359,In_370,In_635);
xor U360 (N_360,In_114,In_591);
xor U361 (N_361,In_253,In_427);
nor U362 (N_362,In_386,In_424);
and U363 (N_363,In_166,In_289);
nand U364 (N_364,In_714,In_573);
or U365 (N_365,In_7,In_234);
and U366 (N_366,In_729,In_599);
and U367 (N_367,In_291,In_445);
nand U368 (N_368,In_58,In_179);
and U369 (N_369,In_323,In_258);
or U370 (N_370,In_87,In_257);
or U371 (N_371,In_746,In_451);
nand U372 (N_372,In_198,In_80);
nor U373 (N_373,In_157,In_557);
nand U374 (N_374,In_301,In_431);
and U375 (N_375,In_728,In_545);
nand U376 (N_376,In_114,In_444);
nand U377 (N_377,In_669,In_109);
and U378 (N_378,In_218,In_727);
nand U379 (N_379,In_584,In_270);
nand U380 (N_380,In_655,In_28);
nor U381 (N_381,In_547,In_415);
nor U382 (N_382,In_235,In_33);
or U383 (N_383,In_639,In_295);
or U384 (N_384,In_738,In_149);
and U385 (N_385,In_310,In_422);
nor U386 (N_386,In_434,In_618);
or U387 (N_387,In_257,In_602);
or U388 (N_388,In_91,In_727);
or U389 (N_389,In_598,In_710);
or U390 (N_390,In_344,In_467);
nand U391 (N_391,In_0,In_443);
nand U392 (N_392,In_273,In_223);
nor U393 (N_393,In_326,In_277);
nor U394 (N_394,In_33,In_149);
nor U395 (N_395,In_539,In_311);
and U396 (N_396,In_558,In_174);
or U397 (N_397,In_485,In_652);
nor U398 (N_398,In_647,In_581);
nand U399 (N_399,In_730,In_186);
nor U400 (N_400,In_477,In_692);
and U401 (N_401,In_366,In_175);
nand U402 (N_402,In_517,In_521);
and U403 (N_403,In_396,In_200);
and U404 (N_404,In_637,In_309);
or U405 (N_405,In_739,In_45);
nand U406 (N_406,In_681,In_133);
and U407 (N_407,In_332,In_574);
or U408 (N_408,In_642,In_379);
nor U409 (N_409,In_356,In_145);
and U410 (N_410,In_654,In_663);
or U411 (N_411,In_6,In_283);
nand U412 (N_412,In_476,In_423);
nor U413 (N_413,In_283,In_49);
nand U414 (N_414,In_646,In_383);
and U415 (N_415,In_183,In_362);
or U416 (N_416,In_517,In_245);
nor U417 (N_417,In_734,In_610);
or U418 (N_418,In_399,In_124);
nor U419 (N_419,In_366,In_130);
and U420 (N_420,In_442,In_681);
nand U421 (N_421,In_367,In_266);
or U422 (N_422,In_539,In_86);
and U423 (N_423,In_296,In_201);
or U424 (N_424,In_344,In_86);
nor U425 (N_425,In_391,In_381);
nor U426 (N_426,In_665,In_714);
and U427 (N_427,In_713,In_64);
xnor U428 (N_428,In_381,In_261);
nor U429 (N_429,In_384,In_85);
or U430 (N_430,In_589,In_638);
or U431 (N_431,In_45,In_280);
nor U432 (N_432,In_266,In_13);
nor U433 (N_433,In_267,In_724);
or U434 (N_434,In_551,In_660);
and U435 (N_435,In_556,In_421);
or U436 (N_436,In_485,In_268);
or U437 (N_437,In_520,In_466);
or U438 (N_438,In_598,In_536);
or U439 (N_439,In_232,In_377);
or U440 (N_440,In_462,In_676);
nand U441 (N_441,In_732,In_580);
or U442 (N_442,In_100,In_93);
and U443 (N_443,In_187,In_735);
and U444 (N_444,In_553,In_245);
nor U445 (N_445,In_605,In_391);
nor U446 (N_446,In_566,In_346);
nor U447 (N_447,In_377,In_352);
and U448 (N_448,In_286,In_12);
and U449 (N_449,In_633,In_615);
and U450 (N_450,In_742,In_326);
xnor U451 (N_451,In_273,In_339);
and U452 (N_452,In_435,In_219);
nor U453 (N_453,In_528,In_175);
and U454 (N_454,In_205,In_484);
nor U455 (N_455,In_102,In_16);
nand U456 (N_456,In_567,In_650);
nor U457 (N_457,In_687,In_737);
or U458 (N_458,In_629,In_504);
nand U459 (N_459,In_550,In_556);
and U460 (N_460,In_603,In_453);
nor U461 (N_461,In_382,In_541);
nor U462 (N_462,In_381,In_451);
or U463 (N_463,In_339,In_347);
and U464 (N_464,In_316,In_48);
nand U465 (N_465,In_116,In_441);
nor U466 (N_466,In_552,In_257);
or U467 (N_467,In_579,In_288);
nor U468 (N_468,In_345,In_193);
nand U469 (N_469,In_440,In_447);
and U470 (N_470,In_128,In_11);
and U471 (N_471,In_653,In_278);
xnor U472 (N_472,In_101,In_49);
nor U473 (N_473,In_313,In_594);
nand U474 (N_474,In_390,In_711);
xor U475 (N_475,In_504,In_95);
nand U476 (N_476,In_702,In_547);
nand U477 (N_477,In_714,In_652);
and U478 (N_478,In_533,In_468);
and U479 (N_479,In_738,In_408);
nor U480 (N_480,In_262,In_467);
nor U481 (N_481,In_705,In_454);
or U482 (N_482,In_683,In_341);
nor U483 (N_483,In_645,In_305);
nor U484 (N_484,In_295,In_160);
nor U485 (N_485,In_194,In_219);
nor U486 (N_486,In_706,In_33);
and U487 (N_487,In_214,In_111);
and U488 (N_488,In_595,In_72);
nand U489 (N_489,In_225,In_464);
or U490 (N_490,In_272,In_416);
or U491 (N_491,In_541,In_244);
and U492 (N_492,In_310,In_518);
and U493 (N_493,In_407,In_498);
and U494 (N_494,In_589,In_243);
and U495 (N_495,In_698,In_719);
and U496 (N_496,In_144,In_708);
and U497 (N_497,In_263,In_60);
and U498 (N_498,In_319,In_23);
and U499 (N_499,In_89,In_575);
or U500 (N_500,In_224,In_367);
nand U501 (N_501,In_52,In_335);
and U502 (N_502,In_551,In_309);
and U503 (N_503,In_430,In_237);
xnor U504 (N_504,In_119,In_304);
nand U505 (N_505,In_196,In_311);
nor U506 (N_506,In_531,In_161);
nor U507 (N_507,In_550,In_85);
nand U508 (N_508,In_227,In_129);
xnor U509 (N_509,In_85,In_467);
or U510 (N_510,In_428,In_328);
or U511 (N_511,In_289,In_717);
nand U512 (N_512,In_337,In_297);
nand U513 (N_513,In_520,In_571);
nand U514 (N_514,In_191,In_540);
nand U515 (N_515,In_739,In_495);
nand U516 (N_516,In_231,In_704);
nor U517 (N_517,In_59,In_483);
and U518 (N_518,In_645,In_192);
xor U519 (N_519,In_518,In_618);
or U520 (N_520,In_178,In_673);
and U521 (N_521,In_407,In_25);
nand U522 (N_522,In_229,In_419);
nand U523 (N_523,In_338,In_694);
or U524 (N_524,In_326,In_360);
and U525 (N_525,In_70,In_645);
or U526 (N_526,In_242,In_314);
nand U527 (N_527,In_118,In_159);
or U528 (N_528,In_452,In_382);
and U529 (N_529,In_60,In_258);
and U530 (N_530,In_11,In_73);
and U531 (N_531,In_446,In_413);
nor U532 (N_532,In_308,In_107);
and U533 (N_533,In_695,In_554);
nor U534 (N_534,In_23,In_589);
nor U535 (N_535,In_291,In_201);
or U536 (N_536,In_173,In_387);
nor U537 (N_537,In_31,In_479);
xnor U538 (N_538,In_241,In_389);
or U539 (N_539,In_402,In_489);
nand U540 (N_540,In_16,In_475);
xnor U541 (N_541,In_739,In_121);
nand U542 (N_542,In_552,In_77);
nor U543 (N_543,In_556,In_621);
nor U544 (N_544,In_510,In_78);
or U545 (N_545,In_361,In_592);
or U546 (N_546,In_646,In_499);
and U547 (N_547,In_490,In_480);
nor U548 (N_548,In_88,In_319);
and U549 (N_549,In_45,In_451);
and U550 (N_550,In_315,In_361);
nor U551 (N_551,In_483,In_119);
nand U552 (N_552,In_144,In_749);
and U553 (N_553,In_737,In_70);
or U554 (N_554,In_707,In_364);
or U555 (N_555,In_608,In_469);
nand U556 (N_556,In_673,In_537);
xnor U557 (N_557,In_638,In_349);
or U558 (N_558,In_133,In_466);
nand U559 (N_559,In_645,In_178);
nor U560 (N_560,In_5,In_655);
nand U561 (N_561,In_238,In_746);
or U562 (N_562,In_497,In_42);
nor U563 (N_563,In_534,In_451);
nor U564 (N_564,In_589,In_39);
or U565 (N_565,In_245,In_344);
or U566 (N_566,In_344,In_310);
nor U567 (N_567,In_34,In_85);
nor U568 (N_568,In_600,In_413);
and U569 (N_569,In_137,In_497);
and U570 (N_570,In_208,In_119);
and U571 (N_571,In_170,In_606);
nor U572 (N_572,In_323,In_52);
nand U573 (N_573,In_358,In_460);
and U574 (N_574,In_328,In_680);
nand U575 (N_575,In_466,In_726);
nor U576 (N_576,In_333,In_273);
and U577 (N_577,In_610,In_576);
or U578 (N_578,In_420,In_579);
nor U579 (N_579,In_342,In_696);
or U580 (N_580,In_325,In_312);
nor U581 (N_581,In_648,In_584);
nand U582 (N_582,In_447,In_605);
nor U583 (N_583,In_116,In_80);
or U584 (N_584,In_594,In_566);
xor U585 (N_585,In_569,In_251);
and U586 (N_586,In_423,In_671);
nand U587 (N_587,In_443,In_677);
and U588 (N_588,In_79,In_357);
nand U589 (N_589,In_744,In_180);
or U590 (N_590,In_138,In_344);
xnor U591 (N_591,In_53,In_95);
nand U592 (N_592,In_299,In_256);
and U593 (N_593,In_494,In_297);
nor U594 (N_594,In_394,In_339);
nor U595 (N_595,In_738,In_57);
and U596 (N_596,In_745,In_551);
or U597 (N_597,In_339,In_202);
nor U598 (N_598,In_576,In_659);
nand U599 (N_599,In_19,In_676);
or U600 (N_600,In_270,In_406);
nor U601 (N_601,In_405,In_569);
nand U602 (N_602,In_444,In_223);
nand U603 (N_603,In_742,In_235);
and U604 (N_604,In_547,In_462);
nor U605 (N_605,In_87,In_644);
and U606 (N_606,In_464,In_176);
or U607 (N_607,In_720,In_320);
and U608 (N_608,In_617,In_597);
nand U609 (N_609,In_481,In_190);
nand U610 (N_610,In_260,In_197);
and U611 (N_611,In_345,In_617);
nand U612 (N_612,In_739,In_469);
nand U613 (N_613,In_80,In_418);
nand U614 (N_614,In_55,In_87);
or U615 (N_615,In_400,In_254);
and U616 (N_616,In_236,In_611);
nor U617 (N_617,In_222,In_478);
nand U618 (N_618,In_482,In_584);
or U619 (N_619,In_464,In_40);
or U620 (N_620,In_318,In_246);
or U621 (N_621,In_219,In_617);
and U622 (N_622,In_540,In_480);
nor U623 (N_623,In_650,In_41);
nor U624 (N_624,In_690,In_705);
or U625 (N_625,In_248,In_124);
nand U626 (N_626,In_260,In_67);
nand U627 (N_627,In_243,In_175);
nor U628 (N_628,In_597,In_55);
nor U629 (N_629,In_624,In_595);
or U630 (N_630,In_472,In_686);
or U631 (N_631,In_587,In_410);
nand U632 (N_632,In_657,In_171);
nor U633 (N_633,In_225,In_278);
or U634 (N_634,In_382,In_28);
and U635 (N_635,In_655,In_60);
nand U636 (N_636,In_589,In_291);
nand U637 (N_637,In_52,In_242);
xnor U638 (N_638,In_723,In_497);
nand U639 (N_639,In_634,In_393);
and U640 (N_640,In_330,In_532);
and U641 (N_641,In_573,In_408);
nor U642 (N_642,In_617,In_549);
nor U643 (N_643,In_477,In_338);
or U644 (N_644,In_396,In_557);
and U645 (N_645,In_411,In_358);
nand U646 (N_646,In_546,In_322);
nor U647 (N_647,In_683,In_195);
nand U648 (N_648,In_245,In_557);
nand U649 (N_649,In_16,In_286);
nand U650 (N_650,In_503,In_95);
and U651 (N_651,In_541,In_624);
or U652 (N_652,In_408,In_146);
nor U653 (N_653,In_709,In_390);
nor U654 (N_654,In_40,In_398);
nor U655 (N_655,In_632,In_116);
nand U656 (N_656,In_20,In_357);
and U657 (N_657,In_452,In_537);
nand U658 (N_658,In_369,In_312);
nor U659 (N_659,In_318,In_745);
and U660 (N_660,In_523,In_49);
nand U661 (N_661,In_264,In_135);
nor U662 (N_662,In_567,In_325);
and U663 (N_663,In_557,In_49);
and U664 (N_664,In_339,In_313);
or U665 (N_665,In_162,In_247);
and U666 (N_666,In_53,In_661);
and U667 (N_667,In_392,In_137);
or U668 (N_668,In_379,In_459);
nor U669 (N_669,In_511,In_81);
or U670 (N_670,In_352,In_150);
xor U671 (N_671,In_607,In_439);
and U672 (N_672,In_621,In_0);
nand U673 (N_673,In_224,In_38);
or U674 (N_674,In_374,In_545);
and U675 (N_675,In_529,In_712);
nor U676 (N_676,In_511,In_377);
nand U677 (N_677,In_227,In_409);
nand U678 (N_678,In_337,In_689);
nor U679 (N_679,In_590,In_669);
nor U680 (N_680,In_713,In_420);
nand U681 (N_681,In_532,In_313);
nand U682 (N_682,In_258,In_201);
nor U683 (N_683,In_430,In_448);
nor U684 (N_684,In_406,In_646);
and U685 (N_685,In_328,In_115);
nand U686 (N_686,In_549,In_730);
and U687 (N_687,In_296,In_118);
and U688 (N_688,In_178,In_732);
or U689 (N_689,In_204,In_390);
nor U690 (N_690,In_572,In_361);
or U691 (N_691,In_420,In_668);
and U692 (N_692,In_617,In_150);
or U693 (N_693,In_548,In_381);
nor U694 (N_694,In_362,In_589);
nand U695 (N_695,In_608,In_23);
and U696 (N_696,In_399,In_311);
nor U697 (N_697,In_87,In_729);
or U698 (N_698,In_6,In_156);
nand U699 (N_699,In_552,In_305);
nand U700 (N_700,In_378,In_579);
or U701 (N_701,In_578,In_424);
nand U702 (N_702,In_179,In_464);
nand U703 (N_703,In_471,In_261);
nand U704 (N_704,In_391,In_159);
and U705 (N_705,In_641,In_302);
nand U706 (N_706,In_379,In_390);
or U707 (N_707,In_740,In_578);
nand U708 (N_708,In_280,In_668);
nand U709 (N_709,In_90,In_508);
and U710 (N_710,In_483,In_624);
or U711 (N_711,In_215,In_232);
nor U712 (N_712,In_237,In_103);
and U713 (N_713,In_139,In_222);
and U714 (N_714,In_429,In_72);
or U715 (N_715,In_506,In_325);
nor U716 (N_716,In_512,In_602);
nor U717 (N_717,In_354,In_462);
xnor U718 (N_718,In_316,In_739);
and U719 (N_719,In_732,In_11);
nor U720 (N_720,In_41,In_51);
nand U721 (N_721,In_439,In_57);
or U722 (N_722,In_568,In_677);
nor U723 (N_723,In_506,In_721);
nand U724 (N_724,In_229,In_131);
nand U725 (N_725,In_670,In_734);
nand U726 (N_726,In_341,In_66);
or U727 (N_727,In_178,In_71);
nand U728 (N_728,In_669,In_427);
and U729 (N_729,In_92,In_709);
and U730 (N_730,In_141,In_252);
or U731 (N_731,In_586,In_63);
nand U732 (N_732,In_87,In_287);
or U733 (N_733,In_516,In_189);
and U734 (N_734,In_513,In_151);
nor U735 (N_735,In_646,In_98);
and U736 (N_736,In_302,In_322);
nor U737 (N_737,In_336,In_687);
nor U738 (N_738,In_620,In_336);
or U739 (N_739,In_519,In_477);
or U740 (N_740,In_516,In_611);
and U741 (N_741,In_589,In_683);
and U742 (N_742,In_47,In_481);
nor U743 (N_743,In_647,In_501);
xor U744 (N_744,In_316,In_138);
and U745 (N_745,In_378,In_449);
nand U746 (N_746,In_348,In_711);
nor U747 (N_747,In_82,In_286);
and U748 (N_748,In_315,In_489);
nand U749 (N_749,In_498,In_728);
nor U750 (N_750,In_534,In_278);
and U751 (N_751,In_330,In_156);
nor U752 (N_752,In_431,In_453);
and U753 (N_753,In_714,In_185);
nor U754 (N_754,In_535,In_200);
nand U755 (N_755,In_494,In_128);
xor U756 (N_756,In_16,In_189);
nand U757 (N_757,In_445,In_90);
and U758 (N_758,In_306,In_154);
and U759 (N_759,In_63,In_28);
nor U760 (N_760,In_651,In_516);
or U761 (N_761,In_566,In_70);
or U762 (N_762,In_726,In_221);
nor U763 (N_763,In_246,In_732);
or U764 (N_764,In_147,In_379);
nor U765 (N_765,In_517,In_728);
or U766 (N_766,In_384,In_628);
nand U767 (N_767,In_298,In_186);
or U768 (N_768,In_102,In_83);
nor U769 (N_769,In_479,In_151);
nor U770 (N_770,In_56,In_6);
or U771 (N_771,In_113,In_620);
xnor U772 (N_772,In_36,In_337);
nor U773 (N_773,In_172,In_321);
nand U774 (N_774,In_617,In_162);
xor U775 (N_775,In_0,In_700);
or U776 (N_776,In_581,In_436);
and U777 (N_777,In_700,In_627);
or U778 (N_778,In_678,In_577);
or U779 (N_779,In_627,In_648);
or U780 (N_780,In_441,In_177);
or U781 (N_781,In_549,In_487);
nor U782 (N_782,In_37,In_441);
and U783 (N_783,In_301,In_147);
nand U784 (N_784,In_731,In_296);
or U785 (N_785,In_299,In_261);
nand U786 (N_786,In_148,In_327);
and U787 (N_787,In_470,In_251);
and U788 (N_788,In_159,In_304);
nand U789 (N_789,In_56,In_548);
nor U790 (N_790,In_564,In_493);
and U791 (N_791,In_94,In_554);
nand U792 (N_792,In_248,In_682);
nor U793 (N_793,In_412,In_278);
nand U794 (N_794,In_663,In_179);
and U795 (N_795,In_98,In_126);
nor U796 (N_796,In_717,In_424);
or U797 (N_797,In_609,In_306);
nor U798 (N_798,In_390,In_502);
nor U799 (N_799,In_432,In_312);
or U800 (N_800,In_565,In_721);
nor U801 (N_801,In_181,In_361);
nand U802 (N_802,In_581,In_330);
or U803 (N_803,In_461,In_343);
and U804 (N_804,In_683,In_689);
nor U805 (N_805,In_288,In_85);
or U806 (N_806,In_373,In_110);
and U807 (N_807,In_457,In_157);
nand U808 (N_808,In_185,In_549);
nand U809 (N_809,In_236,In_553);
and U810 (N_810,In_588,In_490);
or U811 (N_811,In_690,In_568);
nor U812 (N_812,In_250,In_530);
nor U813 (N_813,In_521,In_334);
nor U814 (N_814,In_119,In_325);
nand U815 (N_815,In_195,In_249);
and U816 (N_816,In_367,In_518);
or U817 (N_817,In_703,In_200);
or U818 (N_818,In_660,In_557);
nand U819 (N_819,In_202,In_36);
or U820 (N_820,In_480,In_137);
or U821 (N_821,In_12,In_210);
and U822 (N_822,In_482,In_291);
and U823 (N_823,In_56,In_732);
nand U824 (N_824,In_21,In_485);
and U825 (N_825,In_320,In_333);
nand U826 (N_826,In_512,In_463);
and U827 (N_827,In_714,In_227);
and U828 (N_828,In_662,In_506);
nor U829 (N_829,In_499,In_251);
nor U830 (N_830,In_664,In_747);
nand U831 (N_831,In_197,In_701);
and U832 (N_832,In_652,In_46);
and U833 (N_833,In_333,In_219);
nor U834 (N_834,In_737,In_114);
nor U835 (N_835,In_29,In_501);
nand U836 (N_836,In_81,In_138);
xor U837 (N_837,In_28,In_336);
or U838 (N_838,In_319,In_289);
and U839 (N_839,In_108,In_370);
and U840 (N_840,In_223,In_83);
or U841 (N_841,In_429,In_687);
nor U842 (N_842,In_640,In_504);
nand U843 (N_843,In_635,In_63);
nand U844 (N_844,In_110,In_72);
nand U845 (N_845,In_691,In_601);
nor U846 (N_846,In_104,In_595);
and U847 (N_847,In_487,In_168);
nand U848 (N_848,In_514,In_20);
nand U849 (N_849,In_449,In_42);
nor U850 (N_850,In_143,In_377);
nand U851 (N_851,In_216,In_574);
nand U852 (N_852,In_496,In_63);
and U853 (N_853,In_327,In_235);
or U854 (N_854,In_355,In_298);
nand U855 (N_855,In_201,In_607);
nand U856 (N_856,In_292,In_194);
xnor U857 (N_857,In_505,In_270);
or U858 (N_858,In_473,In_134);
nor U859 (N_859,In_312,In_156);
and U860 (N_860,In_154,In_459);
nand U861 (N_861,In_547,In_642);
or U862 (N_862,In_432,In_338);
nand U863 (N_863,In_336,In_329);
nand U864 (N_864,In_319,In_28);
and U865 (N_865,In_7,In_389);
or U866 (N_866,In_631,In_326);
and U867 (N_867,In_81,In_123);
nor U868 (N_868,In_427,In_339);
nand U869 (N_869,In_339,In_71);
nor U870 (N_870,In_115,In_272);
nand U871 (N_871,In_404,In_547);
nand U872 (N_872,In_373,In_288);
nor U873 (N_873,In_451,In_392);
and U874 (N_874,In_142,In_230);
xor U875 (N_875,In_228,In_700);
nor U876 (N_876,In_327,In_97);
nand U877 (N_877,In_104,In_109);
nand U878 (N_878,In_222,In_174);
or U879 (N_879,In_566,In_369);
nand U880 (N_880,In_57,In_396);
nand U881 (N_881,In_17,In_484);
and U882 (N_882,In_661,In_111);
nor U883 (N_883,In_465,In_437);
nand U884 (N_884,In_174,In_434);
nand U885 (N_885,In_748,In_575);
nand U886 (N_886,In_641,In_49);
and U887 (N_887,In_279,In_388);
or U888 (N_888,In_574,In_168);
or U889 (N_889,In_374,In_145);
nor U890 (N_890,In_321,In_402);
and U891 (N_891,In_568,In_570);
nand U892 (N_892,In_479,In_156);
nand U893 (N_893,In_639,In_348);
or U894 (N_894,In_338,In_399);
nand U895 (N_895,In_491,In_607);
and U896 (N_896,In_712,In_671);
and U897 (N_897,In_230,In_686);
or U898 (N_898,In_499,In_447);
or U899 (N_899,In_657,In_464);
and U900 (N_900,In_122,In_271);
and U901 (N_901,In_747,In_672);
and U902 (N_902,In_275,In_89);
or U903 (N_903,In_29,In_633);
and U904 (N_904,In_648,In_96);
or U905 (N_905,In_29,In_747);
or U906 (N_906,In_436,In_171);
nand U907 (N_907,In_152,In_435);
or U908 (N_908,In_242,In_560);
or U909 (N_909,In_503,In_604);
nor U910 (N_910,In_286,In_500);
or U911 (N_911,In_7,In_324);
nor U912 (N_912,In_731,In_176);
or U913 (N_913,In_566,In_446);
and U914 (N_914,In_98,In_690);
and U915 (N_915,In_483,In_493);
nor U916 (N_916,In_51,In_182);
nand U917 (N_917,In_535,In_176);
nor U918 (N_918,In_365,In_1);
nor U919 (N_919,In_633,In_309);
nor U920 (N_920,In_18,In_598);
or U921 (N_921,In_418,In_12);
xor U922 (N_922,In_337,In_298);
nand U923 (N_923,In_504,In_91);
nor U924 (N_924,In_473,In_61);
nor U925 (N_925,In_129,In_143);
nor U926 (N_926,In_457,In_251);
or U927 (N_927,In_659,In_112);
nor U928 (N_928,In_403,In_508);
nand U929 (N_929,In_52,In_405);
xnor U930 (N_930,In_330,In_485);
nor U931 (N_931,In_545,In_439);
xor U932 (N_932,In_325,In_709);
nor U933 (N_933,In_698,In_693);
nand U934 (N_934,In_411,In_310);
nand U935 (N_935,In_60,In_120);
nor U936 (N_936,In_504,In_727);
or U937 (N_937,In_343,In_151);
or U938 (N_938,In_343,In_49);
or U939 (N_939,In_517,In_623);
and U940 (N_940,In_85,In_254);
and U941 (N_941,In_151,In_587);
nor U942 (N_942,In_440,In_486);
and U943 (N_943,In_367,In_191);
and U944 (N_944,In_715,In_552);
and U945 (N_945,In_64,In_669);
or U946 (N_946,In_536,In_62);
nand U947 (N_947,In_305,In_167);
nor U948 (N_948,In_353,In_719);
or U949 (N_949,In_19,In_478);
or U950 (N_950,In_745,In_520);
nor U951 (N_951,In_578,In_489);
or U952 (N_952,In_306,In_742);
nor U953 (N_953,In_588,In_374);
and U954 (N_954,In_181,In_383);
nand U955 (N_955,In_272,In_181);
and U956 (N_956,In_467,In_322);
nor U957 (N_957,In_705,In_4);
nand U958 (N_958,In_214,In_397);
nand U959 (N_959,In_659,In_86);
and U960 (N_960,In_68,In_25);
nand U961 (N_961,In_115,In_285);
nand U962 (N_962,In_377,In_30);
or U963 (N_963,In_376,In_623);
or U964 (N_964,In_356,In_365);
nor U965 (N_965,In_24,In_45);
or U966 (N_966,In_73,In_301);
and U967 (N_967,In_196,In_519);
nand U968 (N_968,In_129,In_149);
and U969 (N_969,In_497,In_227);
or U970 (N_970,In_534,In_410);
nand U971 (N_971,In_262,In_639);
nand U972 (N_972,In_155,In_165);
and U973 (N_973,In_294,In_13);
or U974 (N_974,In_632,In_208);
and U975 (N_975,In_720,In_157);
nor U976 (N_976,In_195,In_427);
nand U977 (N_977,In_604,In_237);
or U978 (N_978,In_633,In_742);
and U979 (N_979,In_257,In_290);
nand U980 (N_980,In_627,In_255);
nor U981 (N_981,In_192,In_75);
or U982 (N_982,In_568,In_258);
or U983 (N_983,In_246,In_427);
and U984 (N_984,In_552,In_517);
and U985 (N_985,In_352,In_365);
nand U986 (N_986,In_420,In_431);
and U987 (N_987,In_196,In_326);
nor U988 (N_988,In_367,In_153);
or U989 (N_989,In_669,In_479);
or U990 (N_990,In_694,In_730);
nand U991 (N_991,In_572,In_426);
nand U992 (N_992,In_509,In_687);
nor U993 (N_993,In_565,In_336);
nand U994 (N_994,In_141,In_309);
nand U995 (N_995,In_705,In_435);
nor U996 (N_996,In_263,In_306);
and U997 (N_997,In_341,In_318);
nand U998 (N_998,In_579,In_664);
nand U999 (N_999,In_88,In_160);
or U1000 (N_1000,In_137,In_552);
nand U1001 (N_1001,In_101,In_8);
nor U1002 (N_1002,In_240,In_175);
or U1003 (N_1003,In_428,In_187);
or U1004 (N_1004,In_644,In_178);
nand U1005 (N_1005,In_338,In_688);
nor U1006 (N_1006,In_115,In_492);
or U1007 (N_1007,In_284,In_357);
or U1008 (N_1008,In_591,In_738);
nor U1009 (N_1009,In_79,In_201);
nor U1010 (N_1010,In_74,In_180);
nand U1011 (N_1011,In_731,In_367);
nand U1012 (N_1012,In_409,In_610);
nand U1013 (N_1013,In_286,In_698);
or U1014 (N_1014,In_454,In_23);
nand U1015 (N_1015,In_171,In_41);
and U1016 (N_1016,In_134,In_612);
nand U1017 (N_1017,In_281,In_670);
nor U1018 (N_1018,In_741,In_472);
nor U1019 (N_1019,In_504,In_538);
nand U1020 (N_1020,In_272,In_745);
and U1021 (N_1021,In_116,In_542);
or U1022 (N_1022,In_289,In_521);
nor U1023 (N_1023,In_623,In_167);
nor U1024 (N_1024,In_539,In_504);
nor U1025 (N_1025,In_261,In_17);
or U1026 (N_1026,In_197,In_725);
and U1027 (N_1027,In_31,In_378);
nand U1028 (N_1028,In_226,In_625);
nor U1029 (N_1029,In_101,In_562);
or U1030 (N_1030,In_457,In_595);
nor U1031 (N_1031,In_673,In_712);
or U1032 (N_1032,In_479,In_419);
and U1033 (N_1033,In_330,In_488);
nand U1034 (N_1034,In_93,In_414);
or U1035 (N_1035,In_75,In_685);
nand U1036 (N_1036,In_180,In_169);
or U1037 (N_1037,In_35,In_164);
or U1038 (N_1038,In_525,In_240);
and U1039 (N_1039,In_394,In_582);
or U1040 (N_1040,In_434,In_564);
nor U1041 (N_1041,In_288,In_19);
and U1042 (N_1042,In_42,In_664);
nand U1043 (N_1043,In_694,In_54);
or U1044 (N_1044,In_398,In_112);
nand U1045 (N_1045,In_75,In_109);
and U1046 (N_1046,In_492,In_633);
nor U1047 (N_1047,In_368,In_17);
or U1048 (N_1048,In_370,In_339);
and U1049 (N_1049,In_649,In_719);
and U1050 (N_1050,In_482,In_286);
nand U1051 (N_1051,In_662,In_474);
and U1052 (N_1052,In_723,In_623);
and U1053 (N_1053,In_587,In_249);
and U1054 (N_1054,In_30,In_608);
or U1055 (N_1055,In_328,In_59);
and U1056 (N_1056,In_379,In_440);
or U1057 (N_1057,In_365,In_531);
nor U1058 (N_1058,In_41,In_531);
or U1059 (N_1059,In_690,In_236);
nor U1060 (N_1060,In_327,In_4);
nand U1061 (N_1061,In_295,In_417);
nand U1062 (N_1062,In_192,In_456);
and U1063 (N_1063,In_234,In_180);
and U1064 (N_1064,In_456,In_448);
nand U1065 (N_1065,In_398,In_304);
and U1066 (N_1066,In_468,In_716);
nand U1067 (N_1067,In_489,In_132);
nand U1068 (N_1068,In_3,In_703);
nand U1069 (N_1069,In_670,In_501);
nor U1070 (N_1070,In_377,In_342);
or U1071 (N_1071,In_433,In_633);
and U1072 (N_1072,In_598,In_422);
nand U1073 (N_1073,In_453,In_639);
nor U1074 (N_1074,In_109,In_315);
and U1075 (N_1075,In_450,In_385);
nor U1076 (N_1076,In_47,In_497);
nand U1077 (N_1077,In_130,In_49);
nand U1078 (N_1078,In_600,In_152);
xnor U1079 (N_1079,In_172,In_340);
or U1080 (N_1080,In_630,In_687);
and U1081 (N_1081,In_474,In_306);
nand U1082 (N_1082,In_61,In_44);
and U1083 (N_1083,In_625,In_90);
and U1084 (N_1084,In_713,In_654);
nand U1085 (N_1085,In_309,In_545);
nor U1086 (N_1086,In_97,In_277);
nand U1087 (N_1087,In_525,In_230);
or U1088 (N_1088,In_214,In_331);
or U1089 (N_1089,In_630,In_579);
and U1090 (N_1090,In_105,In_20);
nand U1091 (N_1091,In_624,In_581);
and U1092 (N_1092,In_30,In_635);
or U1093 (N_1093,In_88,In_178);
or U1094 (N_1094,In_176,In_565);
or U1095 (N_1095,In_190,In_311);
and U1096 (N_1096,In_96,In_643);
and U1097 (N_1097,In_342,In_188);
and U1098 (N_1098,In_645,In_404);
nand U1099 (N_1099,In_738,In_712);
nand U1100 (N_1100,In_279,In_328);
or U1101 (N_1101,In_341,In_648);
nor U1102 (N_1102,In_338,In_741);
and U1103 (N_1103,In_745,In_218);
or U1104 (N_1104,In_599,In_244);
nand U1105 (N_1105,In_104,In_707);
nor U1106 (N_1106,In_491,In_626);
nand U1107 (N_1107,In_32,In_191);
nor U1108 (N_1108,In_416,In_249);
nand U1109 (N_1109,In_513,In_28);
nand U1110 (N_1110,In_105,In_632);
nor U1111 (N_1111,In_501,In_253);
nand U1112 (N_1112,In_671,In_151);
or U1113 (N_1113,In_589,In_722);
nand U1114 (N_1114,In_496,In_725);
or U1115 (N_1115,In_716,In_350);
or U1116 (N_1116,In_542,In_213);
nor U1117 (N_1117,In_93,In_125);
xnor U1118 (N_1118,In_177,In_523);
nor U1119 (N_1119,In_231,In_271);
nor U1120 (N_1120,In_69,In_394);
nor U1121 (N_1121,In_89,In_191);
nand U1122 (N_1122,In_78,In_12);
nand U1123 (N_1123,In_65,In_359);
and U1124 (N_1124,In_588,In_319);
xor U1125 (N_1125,In_154,In_216);
and U1126 (N_1126,In_522,In_615);
xnor U1127 (N_1127,In_387,In_329);
and U1128 (N_1128,In_32,In_439);
and U1129 (N_1129,In_205,In_100);
and U1130 (N_1130,In_308,In_205);
or U1131 (N_1131,In_429,In_239);
and U1132 (N_1132,In_461,In_137);
nand U1133 (N_1133,In_149,In_152);
nor U1134 (N_1134,In_131,In_424);
and U1135 (N_1135,In_341,In_10);
and U1136 (N_1136,In_748,In_319);
or U1137 (N_1137,In_544,In_528);
nor U1138 (N_1138,In_236,In_172);
nand U1139 (N_1139,In_689,In_651);
nand U1140 (N_1140,In_451,In_709);
and U1141 (N_1141,In_345,In_333);
nand U1142 (N_1142,In_83,In_344);
or U1143 (N_1143,In_381,In_241);
or U1144 (N_1144,In_303,In_650);
nand U1145 (N_1145,In_705,In_56);
or U1146 (N_1146,In_282,In_357);
and U1147 (N_1147,In_5,In_21);
and U1148 (N_1148,In_208,In_400);
or U1149 (N_1149,In_110,In_114);
nor U1150 (N_1150,In_341,In_71);
nor U1151 (N_1151,In_390,In_650);
and U1152 (N_1152,In_740,In_508);
nor U1153 (N_1153,In_688,In_446);
nor U1154 (N_1154,In_293,In_420);
or U1155 (N_1155,In_161,In_421);
and U1156 (N_1156,In_527,In_271);
and U1157 (N_1157,In_490,In_634);
and U1158 (N_1158,In_335,In_438);
nor U1159 (N_1159,In_112,In_654);
or U1160 (N_1160,In_170,In_26);
nor U1161 (N_1161,In_191,In_124);
or U1162 (N_1162,In_312,In_350);
nor U1163 (N_1163,In_618,In_617);
nand U1164 (N_1164,In_680,In_251);
or U1165 (N_1165,In_325,In_275);
nand U1166 (N_1166,In_13,In_69);
nand U1167 (N_1167,In_740,In_435);
or U1168 (N_1168,In_106,In_415);
or U1169 (N_1169,In_222,In_469);
or U1170 (N_1170,In_89,In_706);
or U1171 (N_1171,In_410,In_156);
or U1172 (N_1172,In_385,In_477);
and U1173 (N_1173,In_240,In_392);
or U1174 (N_1174,In_53,In_106);
and U1175 (N_1175,In_502,In_506);
nor U1176 (N_1176,In_710,In_402);
or U1177 (N_1177,In_565,In_275);
and U1178 (N_1178,In_635,In_394);
or U1179 (N_1179,In_350,In_255);
nor U1180 (N_1180,In_137,In_476);
or U1181 (N_1181,In_704,In_285);
nor U1182 (N_1182,In_570,In_611);
and U1183 (N_1183,In_147,In_713);
or U1184 (N_1184,In_10,In_120);
nor U1185 (N_1185,In_34,In_30);
or U1186 (N_1186,In_128,In_350);
nand U1187 (N_1187,In_692,In_274);
nor U1188 (N_1188,In_612,In_529);
and U1189 (N_1189,In_263,In_726);
or U1190 (N_1190,In_744,In_361);
or U1191 (N_1191,In_334,In_547);
nor U1192 (N_1192,In_543,In_120);
or U1193 (N_1193,In_470,In_377);
nor U1194 (N_1194,In_424,In_431);
or U1195 (N_1195,In_524,In_594);
or U1196 (N_1196,In_735,In_61);
nand U1197 (N_1197,In_230,In_568);
nor U1198 (N_1198,In_605,In_204);
or U1199 (N_1199,In_507,In_513);
nand U1200 (N_1200,In_20,In_383);
nand U1201 (N_1201,In_496,In_109);
nor U1202 (N_1202,In_679,In_247);
nand U1203 (N_1203,In_571,In_700);
nor U1204 (N_1204,In_719,In_508);
xnor U1205 (N_1205,In_649,In_443);
nand U1206 (N_1206,In_185,In_684);
nor U1207 (N_1207,In_14,In_238);
or U1208 (N_1208,In_396,In_704);
or U1209 (N_1209,In_158,In_152);
or U1210 (N_1210,In_85,In_563);
xor U1211 (N_1211,In_722,In_596);
nor U1212 (N_1212,In_100,In_456);
xnor U1213 (N_1213,In_450,In_252);
nand U1214 (N_1214,In_207,In_729);
nor U1215 (N_1215,In_607,In_580);
nor U1216 (N_1216,In_443,In_652);
or U1217 (N_1217,In_497,In_267);
nor U1218 (N_1218,In_450,In_521);
nor U1219 (N_1219,In_295,In_141);
nor U1220 (N_1220,In_10,In_565);
nor U1221 (N_1221,In_447,In_114);
and U1222 (N_1222,In_352,In_422);
nand U1223 (N_1223,In_639,In_304);
nand U1224 (N_1224,In_196,In_615);
nor U1225 (N_1225,In_264,In_17);
and U1226 (N_1226,In_35,In_218);
and U1227 (N_1227,In_537,In_169);
nor U1228 (N_1228,In_312,In_297);
and U1229 (N_1229,In_41,In_163);
nor U1230 (N_1230,In_149,In_32);
or U1231 (N_1231,In_115,In_688);
or U1232 (N_1232,In_694,In_94);
and U1233 (N_1233,In_601,In_325);
nor U1234 (N_1234,In_725,In_301);
and U1235 (N_1235,In_729,In_601);
nor U1236 (N_1236,In_175,In_415);
nand U1237 (N_1237,In_536,In_479);
nor U1238 (N_1238,In_196,In_286);
nand U1239 (N_1239,In_589,In_6);
nand U1240 (N_1240,In_113,In_132);
nor U1241 (N_1241,In_364,In_426);
nand U1242 (N_1242,In_665,In_231);
or U1243 (N_1243,In_76,In_407);
and U1244 (N_1244,In_79,In_585);
or U1245 (N_1245,In_318,In_457);
and U1246 (N_1246,In_243,In_321);
or U1247 (N_1247,In_379,In_343);
and U1248 (N_1248,In_85,In_238);
nand U1249 (N_1249,In_295,In_354);
nand U1250 (N_1250,In_82,In_436);
nand U1251 (N_1251,In_517,In_462);
or U1252 (N_1252,In_629,In_654);
and U1253 (N_1253,In_712,In_469);
xnor U1254 (N_1254,In_80,In_325);
nand U1255 (N_1255,In_511,In_484);
or U1256 (N_1256,In_686,In_39);
or U1257 (N_1257,In_399,In_71);
nor U1258 (N_1258,In_639,In_226);
nand U1259 (N_1259,In_121,In_705);
and U1260 (N_1260,In_21,In_313);
nor U1261 (N_1261,In_295,In_610);
xnor U1262 (N_1262,In_250,In_157);
or U1263 (N_1263,In_90,In_701);
nand U1264 (N_1264,In_667,In_313);
nand U1265 (N_1265,In_135,In_486);
and U1266 (N_1266,In_207,In_522);
and U1267 (N_1267,In_133,In_398);
or U1268 (N_1268,In_199,In_217);
nor U1269 (N_1269,In_562,In_732);
nand U1270 (N_1270,In_714,In_724);
nor U1271 (N_1271,In_693,In_539);
or U1272 (N_1272,In_458,In_174);
nor U1273 (N_1273,In_601,In_427);
and U1274 (N_1274,In_188,In_508);
nand U1275 (N_1275,In_446,In_388);
or U1276 (N_1276,In_50,In_577);
nor U1277 (N_1277,In_209,In_377);
or U1278 (N_1278,In_277,In_575);
nor U1279 (N_1279,In_671,In_266);
nor U1280 (N_1280,In_682,In_449);
or U1281 (N_1281,In_344,In_80);
or U1282 (N_1282,In_684,In_462);
nand U1283 (N_1283,In_135,In_352);
nand U1284 (N_1284,In_347,In_443);
and U1285 (N_1285,In_201,In_593);
nor U1286 (N_1286,In_23,In_649);
or U1287 (N_1287,In_257,In_375);
and U1288 (N_1288,In_280,In_598);
and U1289 (N_1289,In_560,In_459);
nor U1290 (N_1290,In_736,In_621);
nand U1291 (N_1291,In_435,In_482);
or U1292 (N_1292,In_214,In_676);
and U1293 (N_1293,In_208,In_25);
or U1294 (N_1294,In_200,In_408);
and U1295 (N_1295,In_252,In_388);
nand U1296 (N_1296,In_300,In_100);
nor U1297 (N_1297,In_642,In_111);
or U1298 (N_1298,In_164,In_230);
nor U1299 (N_1299,In_624,In_132);
and U1300 (N_1300,In_611,In_453);
and U1301 (N_1301,In_70,In_45);
or U1302 (N_1302,In_219,In_536);
and U1303 (N_1303,In_353,In_583);
and U1304 (N_1304,In_468,In_222);
nor U1305 (N_1305,In_319,In_273);
and U1306 (N_1306,In_187,In_167);
and U1307 (N_1307,In_241,In_723);
nor U1308 (N_1308,In_677,In_216);
nor U1309 (N_1309,In_464,In_334);
and U1310 (N_1310,In_339,In_448);
or U1311 (N_1311,In_511,In_355);
nand U1312 (N_1312,In_43,In_475);
and U1313 (N_1313,In_118,In_179);
and U1314 (N_1314,In_207,In_555);
and U1315 (N_1315,In_142,In_268);
and U1316 (N_1316,In_627,In_28);
or U1317 (N_1317,In_156,In_578);
and U1318 (N_1318,In_476,In_199);
nor U1319 (N_1319,In_237,In_299);
or U1320 (N_1320,In_134,In_504);
and U1321 (N_1321,In_571,In_585);
nor U1322 (N_1322,In_624,In_255);
nand U1323 (N_1323,In_205,In_126);
or U1324 (N_1324,In_566,In_14);
and U1325 (N_1325,In_136,In_206);
nand U1326 (N_1326,In_622,In_552);
or U1327 (N_1327,In_283,In_237);
xor U1328 (N_1328,In_527,In_209);
and U1329 (N_1329,In_325,In_607);
or U1330 (N_1330,In_568,In_215);
nand U1331 (N_1331,In_51,In_436);
nand U1332 (N_1332,In_741,In_210);
and U1333 (N_1333,In_342,In_184);
or U1334 (N_1334,In_226,In_247);
nor U1335 (N_1335,In_649,In_44);
nor U1336 (N_1336,In_613,In_740);
nor U1337 (N_1337,In_98,In_246);
nor U1338 (N_1338,In_495,In_448);
nor U1339 (N_1339,In_38,In_15);
nor U1340 (N_1340,In_104,In_330);
nand U1341 (N_1341,In_270,In_675);
nor U1342 (N_1342,In_383,In_700);
and U1343 (N_1343,In_229,In_581);
nor U1344 (N_1344,In_565,In_558);
or U1345 (N_1345,In_149,In_77);
nor U1346 (N_1346,In_604,In_236);
nand U1347 (N_1347,In_711,In_746);
and U1348 (N_1348,In_10,In_518);
and U1349 (N_1349,In_293,In_749);
or U1350 (N_1350,In_240,In_484);
nor U1351 (N_1351,In_590,In_696);
or U1352 (N_1352,In_452,In_455);
nand U1353 (N_1353,In_313,In_388);
nand U1354 (N_1354,In_648,In_58);
nand U1355 (N_1355,In_545,In_650);
nor U1356 (N_1356,In_468,In_458);
nand U1357 (N_1357,In_169,In_452);
nand U1358 (N_1358,In_674,In_390);
nor U1359 (N_1359,In_726,In_195);
nand U1360 (N_1360,In_29,In_527);
nand U1361 (N_1361,In_532,In_612);
and U1362 (N_1362,In_364,In_348);
nand U1363 (N_1363,In_649,In_688);
or U1364 (N_1364,In_76,In_430);
nand U1365 (N_1365,In_212,In_560);
or U1366 (N_1366,In_219,In_731);
nor U1367 (N_1367,In_163,In_467);
or U1368 (N_1368,In_91,In_693);
or U1369 (N_1369,In_434,In_690);
nor U1370 (N_1370,In_466,In_19);
nor U1371 (N_1371,In_647,In_251);
nand U1372 (N_1372,In_42,In_139);
nand U1373 (N_1373,In_168,In_714);
or U1374 (N_1374,In_54,In_447);
nor U1375 (N_1375,In_728,In_662);
and U1376 (N_1376,In_480,In_164);
nor U1377 (N_1377,In_379,In_498);
and U1378 (N_1378,In_125,In_559);
nand U1379 (N_1379,In_121,In_107);
nor U1380 (N_1380,In_491,In_320);
or U1381 (N_1381,In_730,In_369);
and U1382 (N_1382,In_615,In_679);
or U1383 (N_1383,In_524,In_521);
nor U1384 (N_1384,In_639,In_359);
and U1385 (N_1385,In_47,In_339);
nor U1386 (N_1386,In_233,In_131);
and U1387 (N_1387,In_707,In_556);
or U1388 (N_1388,In_548,In_664);
or U1389 (N_1389,In_163,In_722);
and U1390 (N_1390,In_71,In_714);
or U1391 (N_1391,In_534,In_19);
nor U1392 (N_1392,In_356,In_547);
nand U1393 (N_1393,In_305,In_76);
nor U1394 (N_1394,In_313,In_442);
and U1395 (N_1395,In_107,In_543);
and U1396 (N_1396,In_71,In_694);
or U1397 (N_1397,In_319,In_447);
or U1398 (N_1398,In_355,In_371);
nand U1399 (N_1399,In_491,In_451);
nand U1400 (N_1400,In_235,In_593);
nor U1401 (N_1401,In_5,In_693);
nor U1402 (N_1402,In_406,In_7);
nand U1403 (N_1403,In_177,In_40);
nand U1404 (N_1404,In_723,In_163);
or U1405 (N_1405,In_563,In_493);
nand U1406 (N_1406,In_349,In_612);
nand U1407 (N_1407,In_234,In_425);
and U1408 (N_1408,In_531,In_154);
or U1409 (N_1409,In_488,In_128);
nand U1410 (N_1410,In_109,In_300);
and U1411 (N_1411,In_88,In_364);
and U1412 (N_1412,In_700,In_147);
nand U1413 (N_1413,In_29,In_123);
nor U1414 (N_1414,In_10,In_152);
or U1415 (N_1415,In_108,In_737);
and U1416 (N_1416,In_573,In_10);
and U1417 (N_1417,In_426,In_613);
nor U1418 (N_1418,In_428,In_707);
nand U1419 (N_1419,In_635,In_501);
nor U1420 (N_1420,In_683,In_128);
or U1421 (N_1421,In_238,In_640);
and U1422 (N_1422,In_394,In_161);
or U1423 (N_1423,In_363,In_54);
and U1424 (N_1424,In_402,In_427);
and U1425 (N_1425,In_54,In_412);
nand U1426 (N_1426,In_325,In_363);
or U1427 (N_1427,In_560,In_587);
xnor U1428 (N_1428,In_217,In_663);
nor U1429 (N_1429,In_537,In_692);
or U1430 (N_1430,In_153,In_724);
and U1431 (N_1431,In_483,In_16);
or U1432 (N_1432,In_208,In_192);
or U1433 (N_1433,In_675,In_150);
nor U1434 (N_1434,In_419,In_497);
xnor U1435 (N_1435,In_600,In_50);
nand U1436 (N_1436,In_596,In_196);
nand U1437 (N_1437,In_675,In_439);
nand U1438 (N_1438,In_237,In_162);
or U1439 (N_1439,In_20,In_289);
and U1440 (N_1440,In_674,In_658);
nand U1441 (N_1441,In_740,In_602);
nand U1442 (N_1442,In_297,In_235);
and U1443 (N_1443,In_628,In_167);
nand U1444 (N_1444,In_672,In_682);
or U1445 (N_1445,In_675,In_578);
or U1446 (N_1446,In_200,In_64);
xnor U1447 (N_1447,In_652,In_738);
and U1448 (N_1448,In_281,In_667);
and U1449 (N_1449,In_130,In_468);
and U1450 (N_1450,In_154,In_705);
or U1451 (N_1451,In_684,In_537);
nand U1452 (N_1452,In_1,In_100);
nor U1453 (N_1453,In_389,In_662);
or U1454 (N_1454,In_246,In_705);
nand U1455 (N_1455,In_41,In_570);
and U1456 (N_1456,In_737,In_703);
xor U1457 (N_1457,In_556,In_696);
nand U1458 (N_1458,In_606,In_554);
and U1459 (N_1459,In_644,In_524);
or U1460 (N_1460,In_23,In_284);
nand U1461 (N_1461,In_153,In_15);
nand U1462 (N_1462,In_392,In_132);
nor U1463 (N_1463,In_63,In_325);
nand U1464 (N_1464,In_220,In_204);
and U1465 (N_1465,In_748,In_737);
nand U1466 (N_1466,In_405,In_459);
nor U1467 (N_1467,In_96,In_249);
xor U1468 (N_1468,In_23,In_480);
or U1469 (N_1469,In_81,In_522);
nor U1470 (N_1470,In_714,In_69);
and U1471 (N_1471,In_583,In_726);
or U1472 (N_1472,In_340,In_291);
nor U1473 (N_1473,In_280,In_87);
nor U1474 (N_1474,In_60,In_641);
and U1475 (N_1475,In_246,In_271);
nor U1476 (N_1476,In_610,In_45);
nand U1477 (N_1477,In_528,In_574);
or U1478 (N_1478,In_342,In_241);
and U1479 (N_1479,In_653,In_698);
nor U1480 (N_1480,In_583,In_484);
and U1481 (N_1481,In_235,In_45);
or U1482 (N_1482,In_41,In_250);
nand U1483 (N_1483,In_679,In_2);
or U1484 (N_1484,In_34,In_43);
and U1485 (N_1485,In_394,In_317);
or U1486 (N_1486,In_157,In_468);
nor U1487 (N_1487,In_423,In_537);
and U1488 (N_1488,In_36,In_97);
or U1489 (N_1489,In_648,In_143);
nor U1490 (N_1490,In_631,In_628);
and U1491 (N_1491,In_223,In_89);
nand U1492 (N_1492,In_517,In_402);
and U1493 (N_1493,In_454,In_372);
or U1494 (N_1494,In_248,In_450);
or U1495 (N_1495,In_199,In_414);
and U1496 (N_1496,In_567,In_366);
and U1497 (N_1497,In_668,In_505);
or U1498 (N_1498,In_219,In_188);
or U1499 (N_1499,In_506,In_351);
or U1500 (N_1500,In_695,In_384);
nor U1501 (N_1501,In_743,In_111);
nor U1502 (N_1502,In_101,In_119);
nand U1503 (N_1503,In_643,In_680);
and U1504 (N_1504,In_582,In_364);
nor U1505 (N_1505,In_512,In_198);
or U1506 (N_1506,In_434,In_185);
nand U1507 (N_1507,In_321,In_34);
nand U1508 (N_1508,In_672,In_34);
or U1509 (N_1509,In_138,In_367);
or U1510 (N_1510,In_99,In_37);
or U1511 (N_1511,In_577,In_198);
nor U1512 (N_1512,In_225,In_709);
nand U1513 (N_1513,In_604,In_617);
nor U1514 (N_1514,In_741,In_343);
nor U1515 (N_1515,In_417,In_489);
nand U1516 (N_1516,In_547,In_616);
nand U1517 (N_1517,In_588,In_180);
nor U1518 (N_1518,In_516,In_548);
and U1519 (N_1519,In_357,In_546);
nor U1520 (N_1520,In_489,In_531);
nand U1521 (N_1521,In_228,In_348);
nand U1522 (N_1522,In_600,In_614);
or U1523 (N_1523,In_646,In_689);
xnor U1524 (N_1524,In_287,In_383);
or U1525 (N_1525,In_385,In_358);
nand U1526 (N_1526,In_220,In_463);
nor U1527 (N_1527,In_716,In_356);
nor U1528 (N_1528,In_139,In_170);
and U1529 (N_1529,In_252,In_329);
nor U1530 (N_1530,In_464,In_80);
or U1531 (N_1531,In_545,In_294);
or U1532 (N_1532,In_146,In_553);
or U1533 (N_1533,In_575,In_665);
nand U1534 (N_1534,In_110,In_245);
and U1535 (N_1535,In_12,In_84);
nand U1536 (N_1536,In_375,In_404);
and U1537 (N_1537,In_4,In_396);
or U1538 (N_1538,In_523,In_120);
nand U1539 (N_1539,In_353,In_577);
and U1540 (N_1540,In_651,In_620);
nand U1541 (N_1541,In_290,In_74);
nand U1542 (N_1542,In_487,In_139);
nor U1543 (N_1543,In_47,In_390);
or U1544 (N_1544,In_610,In_531);
nand U1545 (N_1545,In_330,In_426);
or U1546 (N_1546,In_632,In_694);
nand U1547 (N_1547,In_713,In_631);
nand U1548 (N_1548,In_232,In_163);
nand U1549 (N_1549,In_381,In_462);
or U1550 (N_1550,In_124,In_32);
nor U1551 (N_1551,In_34,In_653);
nand U1552 (N_1552,In_60,In_342);
and U1553 (N_1553,In_670,In_157);
nand U1554 (N_1554,In_687,In_624);
nor U1555 (N_1555,In_151,In_318);
and U1556 (N_1556,In_20,In_144);
nand U1557 (N_1557,In_468,In_419);
nor U1558 (N_1558,In_545,In_138);
nor U1559 (N_1559,In_27,In_619);
xnor U1560 (N_1560,In_344,In_34);
nor U1561 (N_1561,In_694,In_2);
and U1562 (N_1562,In_102,In_233);
nand U1563 (N_1563,In_18,In_613);
nor U1564 (N_1564,In_261,In_449);
nor U1565 (N_1565,In_550,In_645);
and U1566 (N_1566,In_560,In_620);
nor U1567 (N_1567,In_236,In_333);
nand U1568 (N_1568,In_543,In_318);
and U1569 (N_1569,In_276,In_53);
or U1570 (N_1570,In_688,In_295);
nor U1571 (N_1571,In_109,In_319);
or U1572 (N_1572,In_723,In_642);
and U1573 (N_1573,In_298,In_676);
and U1574 (N_1574,In_159,In_439);
and U1575 (N_1575,In_143,In_265);
nor U1576 (N_1576,In_541,In_4);
nand U1577 (N_1577,In_118,In_184);
nor U1578 (N_1578,In_313,In_548);
nor U1579 (N_1579,In_132,In_276);
or U1580 (N_1580,In_545,In_402);
nand U1581 (N_1581,In_87,In_246);
and U1582 (N_1582,In_527,In_715);
nor U1583 (N_1583,In_633,In_650);
or U1584 (N_1584,In_379,In_493);
and U1585 (N_1585,In_294,In_219);
and U1586 (N_1586,In_386,In_30);
and U1587 (N_1587,In_518,In_521);
nor U1588 (N_1588,In_636,In_562);
or U1589 (N_1589,In_527,In_658);
nor U1590 (N_1590,In_391,In_698);
and U1591 (N_1591,In_158,In_169);
nor U1592 (N_1592,In_120,In_297);
and U1593 (N_1593,In_133,In_675);
and U1594 (N_1594,In_26,In_662);
and U1595 (N_1595,In_613,In_108);
nand U1596 (N_1596,In_391,In_87);
nand U1597 (N_1597,In_459,In_544);
nand U1598 (N_1598,In_204,In_346);
and U1599 (N_1599,In_126,In_691);
or U1600 (N_1600,In_188,In_301);
and U1601 (N_1601,In_30,In_291);
nand U1602 (N_1602,In_493,In_41);
nor U1603 (N_1603,In_746,In_134);
nor U1604 (N_1604,In_284,In_471);
and U1605 (N_1605,In_204,In_46);
or U1606 (N_1606,In_672,In_171);
or U1607 (N_1607,In_545,In_312);
nor U1608 (N_1608,In_608,In_738);
nand U1609 (N_1609,In_436,In_135);
and U1610 (N_1610,In_610,In_130);
nand U1611 (N_1611,In_143,In_303);
or U1612 (N_1612,In_376,In_207);
nand U1613 (N_1613,In_399,In_357);
nand U1614 (N_1614,In_648,In_489);
nand U1615 (N_1615,In_409,In_378);
or U1616 (N_1616,In_477,In_666);
xnor U1617 (N_1617,In_105,In_193);
nor U1618 (N_1618,In_122,In_692);
or U1619 (N_1619,In_710,In_122);
nor U1620 (N_1620,In_315,In_5);
xnor U1621 (N_1621,In_58,In_403);
and U1622 (N_1622,In_366,In_592);
nand U1623 (N_1623,In_113,In_682);
or U1624 (N_1624,In_57,In_380);
or U1625 (N_1625,In_627,In_270);
nor U1626 (N_1626,In_690,In_187);
nand U1627 (N_1627,In_686,In_268);
nand U1628 (N_1628,In_72,In_2);
and U1629 (N_1629,In_618,In_425);
nor U1630 (N_1630,In_235,In_575);
and U1631 (N_1631,In_332,In_469);
nor U1632 (N_1632,In_178,In_272);
nor U1633 (N_1633,In_268,In_711);
nor U1634 (N_1634,In_391,In_108);
nand U1635 (N_1635,In_123,In_98);
nor U1636 (N_1636,In_651,In_102);
nor U1637 (N_1637,In_670,In_565);
nor U1638 (N_1638,In_707,In_187);
nor U1639 (N_1639,In_374,In_293);
or U1640 (N_1640,In_91,In_457);
or U1641 (N_1641,In_419,In_730);
nor U1642 (N_1642,In_447,In_650);
and U1643 (N_1643,In_533,In_526);
nand U1644 (N_1644,In_194,In_518);
nand U1645 (N_1645,In_722,In_10);
nor U1646 (N_1646,In_661,In_458);
and U1647 (N_1647,In_403,In_24);
or U1648 (N_1648,In_578,In_610);
and U1649 (N_1649,In_543,In_367);
nor U1650 (N_1650,In_709,In_445);
nand U1651 (N_1651,In_581,In_594);
nand U1652 (N_1652,In_55,In_224);
and U1653 (N_1653,In_284,In_520);
or U1654 (N_1654,In_687,In_441);
nand U1655 (N_1655,In_142,In_572);
nor U1656 (N_1656,In_685,In_347);
or U1657 (N_1657,In_128,In_365);
and U1658 (N_1658,In_164,In_616);
and U1659 (N_1659,In_210,In_270);
or U1660 (N_1660,In_275,In_634);
and U1661 (N_1661,In_340,In_109);
xor U1662 (N_1662,In_440,In_734);
and U1663 (N_1663,In_340,In_170);
and U1664 (N_1664,In_590,In_39);
nand U1665 (N_1665,In_236,In_235);
or U1666 (N_1666,In_354,In_15);
nor U1667 (N_1667,In_288,In_306);
nand U1668 (N_1668,In_15,In_555);
or U1669 (N_1669,In_6,In_723);
and U1670 (N_1670,In_420,In_105);
nand U1671 (N_1671,In_38,In_45);
nand U1672 (N_1672,In_161,In_638);
and U1673 (N_1673,In_729,In_460);
nor U1674 (N_1674,In_30,In_590);
nand U1675 (N_1675,In_295,In_143);
or U1676 (N_1676,In_738,In_103);
nand U1677 (N_1677,In_64,In_139);
nor U1678 (N_1678,In_119,In_463);
nand U1679 (N_1679,In_196,In_10);
xor U1680 (N_1680,In_722,In_398);
and U1681 (N_1681,In_174,In_652);
nand U1682 (N_1682,In_695,In_700);
nand U1683 (N_1683,In_410,In_644);
nor U1684 (N_1684,In_707,In_484);
or U1685 (N_1685,In_421,In_150);
or U1686 (N_1686,In_670,In_474);
nor U1687 (N_1687,In_400,In_86);
nand U1688 (N_1688,In_99,In_534);
xor U1689 (N_1689,In_153,In_619);
and U1690 (N_1690,In_407,In_440);
nor U1691 (N_1691,In_711,In_233);
and U1692 (N_1692,In_222,In_442);
nand U1693 (N_1693,In_164,In_351);
and U1694 (N_1694,In_158,In_206);
nand U1695 (N_1695,In_159,In_233);
or U1696 (N_1696,In_659,In_140);
xor U1697 (N_1697,In_45,In_730);
or U1698 (N_1698,In_619,In_683);
or U1699 (N_1699,In_611,In_191);
nor U1700 (N_1700,In_500,In_18);
or U1701 (N_1701,In_68,In_607);
nand U1702 (N_1702,In_487,In_10);
nand U1703 (N_1703,In_532,In_555);
xnor U1704 (N_1704,In_557,In_17);
nor U1705 (N_1705,In_512,In_290);
nand U1706 (N_1706,In_313,In_511);
and U1707 (N_1707,In_373,In_712);
nand U1708 (N_1708,In_35,In_105);
and U1709 (N_1709,In_78,In_428);
nand U1710 (N_1710,In_198,In_329);
nand U1711 (N_1711,In_482,In_718);
or U1712 (N_1712,In_35,In_334);
nor U1713 (N_1713,In_308,In_440);
nor U1714 (N_1714,In_86,In_530);
or U1715 (N_1715,In_381,In_580);
or U1716 (N_1716,In_547,In_60);
nand U1717 (N_1717,In_357,In_302);
nor U1718 (N_1718,In_48,In_177);
or U1719 (N_1719,In_491,In_663);
nand U1720 (N_1720,In_709,In_254);
or U1721 (N_1721,In_258,In_702);
nand U1722 (N_1722,In_718,In_68);
nand U1723 (N_1723,In_38,In_210);
nor U1724 (N_1724,In_481,In_43);
nand U1725 (N_1725,In_85,In_92);
and U1726 (N_1726,In_636,In_631);
nor U1727 (N_1727,In_492,In_707);
and U1728 (N_1728,In_46,In_483);
nand U1729 (N_1729,In_291,In_27);
or U1730 (N_1730,In_679,In_731);
and U1731 (N_1731,In_603,In_214);
nor U1732 (N_1732,In_686,In_681);
or U1733 (N_1733,In_576,In_215);
nor U1734 (N_1734,In_438,In_140);
and U1735 (N_1735,In_350,In_550);
or U1736 (N_1736,In_225,In_206);
or U1737 (N_1737,In_543,In_140);
nor U1738 (N_1738,In_530,In_664);
xnor U1739 (N_1739,In_380,In_495);
or U1740 (N_1740,In_575,In_404);
and U1741 (N_1741,In_505,In_723);
and U1742 (N_1742,In_42,In_691);
nor U1743 (N_1743,In_531,In_465);
nand U1744 (N_1744,In_621,In_563);
or U1745 (N_1745,In_358,In_399);
nor U1746 (N_1746,In_90,In_601);
or U1747 (N_1747,In_368,In_304);
and U1748 (N_1748,In_325,In_220);
or U1749 (N_1749,In_64,In_427);
or U1750 (N_1750,In_317,In_628);
and U1751 (N_1751,In_414,In_446);
or U1752 (N_1752,In_338,In_543);
nand U1753 (N_1753,In_333,In_573);
nand U1754 (N_1754,In_574,In_741);
nand U1755 (N_1755,In_4,In_368);
and U1756 (N_1756,In_120,In_746);
nor U1757 (N_1757,In_632,In_600);
and U1758 (N_1758,In_686,In_199);
and U1759 (N_1759,In_140,In_521);
nor U1760 (N_1760,In_543,In_40);
or U1761 (N_1761,In_40,In_238);
nor U1762 (N_1762,In_711,In_743);
or U1763 (N_1763,In_444,In_745);
and U1764 (N_1764,In_307,In_46);
nor U1765 (N_1765,In_420,In_367);
nor U1766 (N_1766,In_120,In_725);
nand U1767 (N_1767,In_679,In_397);
nand U1768 (N_1768,In_442,In_676);
nand U1769 (N_1769,In_476,In_58);
nor U1770 (N_1770,In_608,In_436);
nor U1771 (N_1771,In_41,In_0);
nand U1772 (N_1772,In_532,In_643);
or U1773 (N_1773,In_48,In_456);
or U1774 (N_1774,In_539,In_471);
nor U1775 (N_1775,In_373,In_113);
and U1776 (N_1776,In_423,In_58);
and U1777 (N_1777,In_564,In_632);
xnor U1778 (N_1778,In_601,In_230);
and U1779 (N_1779,In_165,In_97);
nand U1780 (N_1780,In_206,In_733);
or U1781 (N_1781,In_375,In_547);
nand U1782 (N_1782,In_99,In_23);
nor U1783 (N_1783,In_699,In_106);
nor U1784 (N_1784,In_154,In_46);
nor U1785 (N_1785,In_329,In_545);
or U1786 (N_1786,In_312,In_116);
nor U1787 (N_1787,In_56,In_725);
nand U1788 (N_1788,In_709,In_79);
or U1789 (N_1789,In_622,In_312);
nor U1790 (N_1790,In_613,In_152);
and U1791 (N_1791,In_597,In_20);
or U1792 (N_1792,In_555,In_417);
nand U1793 (N_1793,In_275,In_93);
nor U1794 (N_1794,In_233,In_30);
nand U1795 (N_1795,In_410,In_81);
or U1796 (N_1796,In_689,In_567);
nand U1797 (N_1797,In_176,In_227);
nand U1798 (N_1798,In_607,In_239);
nand U1799 (N_1799,In_398,In_195);
nand U1800 (N_1800,In_360,In_78);
or U1801 (N_1801,In_713,In_610);
nand U1802 (N_1802,In_431,In_662);
and U1803 (N_1803,In_20,In_395);
or U1804 (N_1804,In_468,In_97);
or U1805 (N_1805,In_635,In_443);
or U1806 (N_1806,In_359,In_264);
nand U1807 (N_1807,In_442,In_598);
nand U1808 (N_1808,In_119,In_398);
and U1809 (N_1809,In_172,In_309);
or U1810 (N_1810,In_476,In_528);
nand U1811 (N_1811,In_695,In_58);
or U1812 (N_1812,In_601,In_292);
nand U1813 (N_1813,In_468,In_465);
nor U1814 (N_1814,In_304,In_593);
or U1815 (N_1815,In_74,In_31);
and U1816 (N_1816,In_670,In_427);
and U1817 (N_1817,In_243,In_453);
and U1818 (N_1818,In_566,In_365);
nor U1819 (N_1819,In_687,In_356);
or U1820 (N_1820,In_641,In_633);
and U1821 (N_1821,In_373,In_65);
nand U1822 (N_1822,In_15,In_35);
or U1823 (N_1823,In_386,In_459);
nor U1824 (N_1824,In_246,In_259);
nor U1825 (N_1825,In_307,In_656);
or U1826 (N_1826,In_315,In_253);
or U1827 (N_1827,In_578,In_183);
nand U1828 (N_1828,In_692,In_132);
nand U1829 (N_1829,In_243,In_296);
nand U1830 (N_1830,In_54,In_314);
and U1831 (N_1831,In_292,In_719);
nand U1832 (N_1832,In_409,In_125);
or U1833 (N_1833,In_101,In_666);
or U1834 (N_1834,In_19,In_266);
and U1835 (N_1835,In_221,In_479);
and U1836 (N_1836,In_464,In_167);
nor U1837 (N_1837,In_549,In_148);
nand U1838 (N_1838,In_61,In_446);
nor U1839 (N_1839,In_312,In_290);
or U1840 (N_1840,In_440,In_618);
or U1841 (N_1841,In_599,In_330);
nor U1842 (N_1842,In_511,In_410);
nand U1843 (N_1843,In_400,In_99);
or U1844 (N_1844,In_502,In_692);
and U1845 (N_1845,In_609,In_196);
or U1846 (N_1846,In_475,In_449);
and U1847 (N_1847,In_327,In_250);
nand U1848 (N_1848,In_596,In_5);
nand U1849 (N_1849,In_632,In_155);
nor U1850 (N_1850,In_200,In_725);
and U1851 (N_1851,In_45,In_540);
nand U1852 (N_1852,In_605,In_440);
or U1853 (N_1853,In_566,In_215);
and U1854 (N_1854,In_228,In_103);
nor U1855 (N_1855,In_424,In_356);
or U1856 (N_1856,In_318,In_286);
or U1857 (N_1857,In_609,In_738);
nand U1858 (N_1858,In_231,In_107);
nand U1859 (N_1859,In_127,In_365);
nand U1860 (N_1860,In_21,In_111);
and U1861 (N_1861,In_638,In_346);
nor U1862 (N_1862,In_93,In_19);
and U1863 (N_1863,In_167,In_408);
xor U1864 (N_1864,In_648,In_741);
or U1865 (N_1865,In_155,In_413);
nor U1866 (N_1866,In_5,In_574);
or U1867 (N_1867,In_56,In_649);
nand U1868 (N_1868,In_164,In_40);
nand U1869 (N_1869,In_261,In_648);
or U1870 (N_1870,In_350,In_252);
xor U1871 (N_1871,In_328,In_37);
or U1872 (N_1872,In_663,In_669);
and U1873 (N_1873,In_235,In_409);
nand U1874 (N_1874,In_118,In_129);
nor U1875 (N_1875,In_70,In_422);
nand U1876 (N_1876,In_528,In_72);
nand U1877 (N_1877,In_246,In_176);
and U1878 (N_1878,In_430,In_579);
nor U1879 (N_1879,In_68,In_342);
nor U1880 (N_1880,In_98,In_188);
nand U1881 (N_1881,In_552,In_217);
nand U1882 (N_1882,In_184,In_482);
or U1883 (N_1883,In_263,In_369);
nand U1884 (N_1884,In_682,In_539);
and U1885 (N_1885,In_189,In_649);
or U1886 (N_1886,In_698,In_686);
nand U1887 (N_1887,In_658,In_728);
and U1888 (N_1888,In_286,In_348);
or U1889 (N_1889,In_399,In_653);
or U1890 (N_1890,In_335,In_388);
and U1891 (N_1891,In_341,In_437);
and U1892 (N_1892,In_408,In_455);
or U1893 (N_1893,In_385,In_433);
or U1894 (N_1894,In_200,In_483);
or U1895 (N_1895,In_405,In_45);
and U1896 (N_1896,In_421,In_145);
nand U1897 (N_1897,In_249,In_684);
and U1898 (N_1898,In_333,In_458);
and U1899 (N_1899,In_370,In_202);
or U1900 (N_1900,In_571,In_51);
nand U1901 (N_1901,In_617,In_709);
nor U1902 (N_1902,In_714,In_557);
xnor U1903 (N_1903,In_236,In_692);
or U1904 (N_1904,In_719,In_290);
and U1905 (N_1905,In_281,In_384);
xnor U1906 (N_1906,In_622,In_19);
nor U1907 (N_1907,In_429,In_209);
or U1908 (N_1908,In_406,In_285);
and U1909 (N_1909,In_285,In_390);
nand U1910 (N_1910,In_324,In_243);
nor U1911 (N_1911,In_649,In_441);
and U1912 (N_1912,In_558,In_394);
nand U1913 (N_1913,In_534,In_1);
nor U1914 (N_1914,In_606,In_0);
nand U1915 (N_1915,In_17,In_133);
and U1916 (N_1916,In_168,In_559);
xor U1917 (N_1917,In_353,In_595);
and U1918 (N_1918,In_293,In_305);
nand U1919 (N_1919,In_63,In_450);
nor U1920 (N_1920,In_426,In_658);
nor U1921 (N_1921,In_539,In_269);
nor U1922 (N_1922,In_398,In_459);
nor U1923 (N_1923,In_562,In_535);
nor U1924 (N_1924,In_59,In_394);
nand U1925 (N_1925,In_253,In_608);
or U1926 (N_1926,In_655,In_475);
and U1927 (N_1927,In_747,In_508);
nor U1928 (N_1928,In_5,In_26);
and U1929 (N_1929,In_521,In_445);
nand U1930 (N_1930,In_445,In_704);
nor U1931 (N_1931,In_499,In_27);
nand U1932 (N_1932,In_326,In_624);
or U1933 (N_1933,In_274,In_435);
or U1934 (N_1934,In_709,In_507);
and U1935 (N_1935,In_339,In_622);
nand U1936 (N_1936,In_492,In_363);
nand U1937 (N_1937,In_625,In_633);
or U1938 (N_1938,In_664,In_650);
nor U1939 (N_1939,In_555,In_369);
or U1940 (N_1940,In_706,In_147);
nand U1941 (N_1941,In_640,In_538);
nor U1942 (N_1942,In_58,In_266);
or U1943 (N_1943,In_47,In_20);
nand U1944 (N_1944,In_605,In_228);
or U1945 (N_1945,In_121,In_89);
nand U1946 (N_1946,In_86,In_357);
nor U1947 (N_1947,In_230,In_133);
or U1948 (N_1948,In_368,In_600);
xnor U1949 (N_1949,In_90,In_418);
and U1950 (N_1950,In_17,In_190);
nor U1951 (N_1951,In_698,In_740);
nor U1952 (N_1952,In_39,In_239);
nor U1953 (N_1953,In_594,In_160);
and U1954 (N_1954,In_611,In_166);
nand U1955 (N_1955,In_178,In_198);
nor U1956 (N_1956,In_655,In_350);
and U1957 (N_1957,In_462,In_189);
and U1958 (N_1958,In_207,In_649);
nand U1959 (N_1959,In_732,In_494);
nand U1960 (N_1960,In_666,In_551);
nor U1961 (N_1961,In_187,In_439);
and U1962 (N_1962,In_490,In_631);
nand U1963 (N_1963,In_547,In_698);
nor U1964 (N_1964,In_361,In_112);
nor U1965 (N_1965,In_103,In_270);
or U1966 (N_1966,In_2,In_142);
and U1967 (N_1967,In_467,In_142);
nor U1968 (N_1968,In_22,In_194);
nor U1969 (N_1969,In_641,In_288);
nor U1970 (N_1970,In_204,In_407);
or U1971 (N_1971,In_321,In_203);
or U1972 (N_1972,In_551,In_292);
nor U1973 (N_1973,In_484,In_254);
and U1974 (N_1974,In_589,In_215);
or U1975 (N_1975,In_326,In_704);
nand U1976 (N_1976,In_269,In_664);
xor U1977 (N_1977,In_501,In_395);
nor U1978 (N_1978,In_486,In_661);
nor U1979 (N_1979,In_79,In_621);
and U1980 (N_1980,In_171,In_594);
or U1981 (N_1981,In_571,In_503);
nor U1982 (N_1982,In_108,In_616);
nand U1983 (N_1983,In_508,In_50);
or U1984 (N_1984,In_208,In_413);
nand U1985 (N_1985,In_289,In_314);
and U1986 (N_1986,In_548,In_532);
nor U1987 (N_1987,In_113,In_462);
and U1988 (N_1988,In_466,In_60);
and U1989 (N_1989,In_440,In_85);
nor U1990 (N_1990,In_63,In_230);
or U1991 (N_1991,In_481,In_630);
nand U1992 (N_1992,In_44,In_734);
and U1993 (N_1993,In_115,In_477);
and U1994 (N_1994,In_384,In_322);
nand U1995 (N_1995,In_434,In_43);
and U1996 (N_1996,In_693,In_215);
and U1997 (N_1997,In_706,In_630);
or U1998 (N_1998,In_348,In_483);
and U1999 (N_1999,In_618,In_591);
nor U2000 (N_2000,In_565,In_258);
nor U2001 (N_2001,In_467,In_342);
nor U2002 (N_2002,In_438,In_353);
and U2003 (N_2003,In_310,In_189);
nand U2004 (N_2004,In_235,In_61);
xor U2005 (N_2005,In_108,In_182);
or U2006 (N_2006,In_740,In_644);
nor U2007 (N_2007,In_565,In_505);
nand U2008 (N_2008,In_600,In_585);
nor U2009 (N_2009,In_422,In_417);
nor U2010 (N_2010,In_427,In_81);
and U2011 (N_2011,In_732,In_550);
nand U2012 (N_2012,In_448,In_88);
nand U2013 (N_2013,In_198,In_336);
nand U2014 (N_2014,In_202,In_680);
nand U2015 (N_2015,In_321,In_636);
or U2016 (N_2016,In_172,In_133);
or U2017 (N_2017,In_2,In_686);
nand U2018 (N_2018,In_521,In_420);
nand U2019 (N_2019,In_77,In_278);
nor U2020 (N_2020,In_385,In_376);
or U2021 (N_2021,In_677,In_482);
and U2022 (N_2022,In_401,In_726);
nand U2023 (N_2023,In_170,In_499);
nor U2024 (N_2024,In_444,In_391);
and U2025 (N_2025,In_4,In_745);
nor U2026 (N_2026,In_525,In_242);
and U2027 (N_2027,In_587,In_69);
and U2028 (N_2028,In_266,In_10);
nand U2029 (N_2029,In_229,In_181);
and U2030 (N_2030,In_222,In_432);
nand U2031 (N_2031,In_360,In_466);
nand U2032 (N_2032,In_465,In_278);
and U2033 (N_2033,In_492,In_655);
nand U2034 (N_2034,In_224,In_357);
nor U2035 (N_2035,In_721,In_530);
nor U2036 (N_2036,In_420,In_166);
and U2037 (N_2037,In_609,In_373);
nor U2038 (N_2038,In_431,In_287);
and U2039 (N_2039,In_431,In_276);
nand U2040 (N_2040,In_244,In_435);
nor U2041 (N_2041,In_743,In_748);
nand U2042 (N_2042,In_296,In_729);
nor U2043 (N_2043,In_34,In_438);
or U2044 (N_2044,In_33,In_160);
or U2045 (N_2045,In_687,In_391);
xnor U2046 (N_2046,In_227,In_403);
or U2047 (N_2047,In_540,In_241);
or U2048 (N_2048,In_14,In_163);
and U2049 (N_2049,In_169,In_123);
and U2050 (N_2050,In_26,In_739);
xor U2051 (N_2051,In_154,In_454);
and U2052 (N_2052,In_318,In_193);
nor U2053 (N_2053,In_373,In_180);
nand U2054 (N_2054,In_696,In_68);
nor U2055 (N_2055,In_708,In_570);
and U2056 (N_2056,In_690,In_737);
and U2057 (N_2057,In_373,In_397);
and U2058 (N_2058,In_251,In_703);
or U2059 (N_2059,In_482,In_615);
and U2060 (N_2060,In_363,In_260);
nor U2061 (N_2061,In_681,In_69);
or U2062 (N_2062,In_199,In_240);
or U2063 (N_2063,In_221,In_500);
nand U2064 (N_2064,In_272,In_723);
and U2065 (N_2065,In_190,In_185);
nand U2066 (N_2066,In_256,In_411);
nand U2067 (N_2067,In_347,In_722);
xnor U2068 (N_2068,In_91,In_218);
and U2069 (N_2069,In_404,In_664);
or U2070 (N_2070,In_218,In_81);
nor U2071 (N_2071,In_585,In_655);
nand U2072 (N_2072,In_233,In_444);
nor U2073 (N_2073,In_624,In_173);
nand U2074 (N_2074,In_578,In_728);
and U2075 (N_2075,In_53,In_235);
xnor U2076 (N_2076,In_273,In_90);
nor U2077 (N_2077,In_515,In_304);
nor U2078 (N_2078,In_59,In_232);
nor U2079 (N_2079,In_529,In_387);
nor U2080 (N_2080,In_41,In_24);
and U2081 (N_2081,In_68,In_694);
or U2082 (N_2082,In_183,In_695);
and U2083 (N_2083,In_411,In_515);
nor U2084 (N_2084,In_195,In_449);
nor U2085 (N_2085,In_482,In_519);
or U2086 (N_2086,In_237,In_213);
or U2087 (N_2087,In_362,In_688);
nand U2088 (N_2088,In_618,In_403);
nand U2089 (N_2089,In_323,In_239);
and U2090 (N_2090,In_740,In_266);
or U2091 (N_2091,In_680,In_538);
or U2092 (N_2092,In_664,In_511);
nand U2093 (N_2093,In_199,In_133);
nor U2094 (N_2094,In_686,In_410);
or U2095 (N_2095,In_216,In_35);
nand U2096 (N_2096,In_579,In_36);
nand U2097 (N_2097,In_380,In_497);
or U2098 (N_2098,In_399,In_734);
nand U2099 (N_2099,In_742,In_412);
or U2100 (N_2100,In_614,In_370);
and U2101 (N_2101,In_210,In_428);
or U2102 (N_2102,In_175,In_66);
nand U2103 (N_2103,In_357,In_524);
and U2104 (N_2104,In_576,In_66);
and U2105 (N_2105,In_249,In_188);
or U2106 (N_2106,In_604,In_338);
nor U2107 (N_2107,In_450,In_392);
or U2108 (N_2108,In_350,In_115);
nand U2109 (N_2109,In_657,In_25);
or U2110 (N_2110,In_382,In_513);
nor U2111 (N_2111,In_147,In_748);
and U2112 (N_2112,In_578,In_624);
nand U2113 (N_2113,In_450,In_722);
or U2114 (N_2114,In_614,In_150);
nor U2115 (N_2115,In_0,In_515);
nand U2116 (N_2116,In_185,In_554);
or U2117 (N_2117,In_546,In_155);
or U2118 (N_2118,In_560,In_360);
and U2119 (N_2119,In_382,In_234);
nor U2120 (N_2120,In_34,In_747);
nor U2121 (N_2121,In_27,In_93);
nand U2122 (N_2122,In_93,In_64);
and U2123 (N_2123,In_276,In_536);
nor U2124 (N_2124,In_261,In_424);
nor U2125 (N_2125,In_386,In_254);
xor U2126 (N_2126,In_361,In_11);
and U2127 (N_2127,In_450,In_231);
or U2128 (N_2128,In_170,In_111);
nor U2129 (N_2129,In_76,In_639);
or U2130 (N_2130,In_702,In_478);
or U2131 (N_2131,In_660,In_118);
or U2132 (N_2132,In_340,In_337);
and U2133 (N_2133,In_387,In_448);
nand U2134 (N_2134,In_82,In_155);
or U2135 (N_2135,In_375,In_154);
or U2136 (N_2136,In_243,In_672);
and U2137 (N_2137,In_254,In_687);
nand U2138 (N_2138,In_287,In_89);
nor U2139 (N_2139,In_733,In_682);
nand U2140 (N_2140,In_618,In_723);
and U2141 (N_2141,In_488,In_11);
xnor U2142 (N_2142,In_25,In_723);
nor U2143 (N_2143,In_207,In_541);
or U2144 (N_2144,In_628,In_252);
nand U2145 (N_2145,In_578,In_240);
nand U2146 (N_2146,In_344,In_222);
nor U2147 (N_2147,In_264,In_610);
and U2148 (N_2148,In_570,In_11);
nor U2149 (N_2149,In_547,In_542);
nand U2150 (N_2150,In_722,In_247);
or U2151 (N_2151,In_272,In_513);
xor U2152 (N_2152,In_119,In_140);
nor U2153 (N_2153,In_428,In_342);
and U2154 (N_2154,In_409,In_661);
or U2155 (N_2155,In_464,In_99);
nor U2156 (N_2156,In_360,In_526);
nand U2157 (N_2157,In_431,In_278);
and U2158 (N_2158,In_473,In_214);
or U2159 (N_2159,In_502,In_352);
or U2160 (N_2160,In_625,In_321);
or U2161 (N_2161,In_563,In_553);
nand U2162 (N_2162,In_1,In_406);
nand U2163 (N_2163,In_666,In_28);
and U2164 (N_2164,In_682,In_83);
nand U2165 (N_2165,In_489,In_223);
or U2166 (N_2166,In_427,In_631);
or U2167 (N_2167,In_100,In_749);
nand U2168 (N_2168,In_388,In_47);
and U2169 (N_2169,In_743,In_313);
nand U2170 (N_2170,In_23,In_610);
nor U2171 (N_2171,In_87,In_221);
nand U2172 (N_2172,In_57,In_289);
nor U2173 (N_2173,In_446,In_621);
nand U2174 (N_2174,In_485,In_187);
or U2175 (N_2175,In_268,In_406);
nor U2176 (N_2176,In_324,In_99);
nor U2177 (N_2177,In_536,In_368);
or U2178 (N_2178,In_120,In_649);
and U2179 (N_2179,In_513,In_404);
nand U2180 (N_2180,In_273,In_377);
or U2181 (N_2181,In_409,In_315);
and U2182 (N_2182,In_481,In_543);
nor U2183 (N_2183,In_397,In_213);
or U2184 (N_2184,In_437,In_504);
nand U2185 (N_2185,In_698,In_232);
nor U2186 (N_2186,In_83,In_596);
and U2187 (N_2187,In_91,In_472);
nand U2188 (N_2188,In_426,In_747);
and U2189 (N_2189,In_527,In_741);
and U2190 (N_2190,In_736,In_88);
or U2191 (N_2191,In_152,In_369);
nand U2192 (N_2192,In_33,In_284);
nand U2193 (N_2193,In_51,In_71);
nand U2194 (N_2194,In_285,In_645);
nor U2195 (N_2195,In_605,In_485);
and U2196 (N_2196,In_221,In_549);
nor U2197 (N_2197,In_320,In_303);
and U2198 (N_2198,In_417,In_322);
or U2199 (N_2199,In_698,In_692);
or U2200 (N_2200,In_476,In_10);
or U2201 (N_2201,In_636,In_741);
and U2202 (N_2202,In_63,In_332);
xnor U2203 (N_2203,In_661,In_342);
or U2204 (N_2204,In_132,In_458);
nor U2205 (N_2205,In_476,In_226);
or U2206 (N_2206,In_26,In_162);
or U2207 (N_2207,In_665,In_69);
nor U2208 (N_2208,In_287,In_320);
nor U2209 (N_2209,In_406,In_48);
nand U2210 (N_2210,In_54,In_544);
or U2211 (N_2211,In_184,In_575);
nand U2212 (N_2212,In_669,In_237);
nor U2213 (N_2213,In_240,In_680);
nand U2214 (N_2214,In_681,In_187);
xor U2215 (N_2215,In_468,In_338);
nand U2216 (N_2216,In_692,In_548);
or U2217 (N_2217,In_254,In_417);
or U2218 (N_2218,In_88,In_111);
and U2219 (N_2219,In_214,In_77);
nand U2220 (N_2220,In_286,In_86);
nor U2221 (N_2221,In_89,In_2);
nand U2222 (N_2222,In_47,In_345);
nor U2223 (N_2223,In_237,In_650);
and U2224 (N_2224,In_56,In_276);
xnor U2225 (N_2225,In_8,In_38);
nand U2226 (N_2226,In_417,In_35);
nand U2227 (N_2227,In_263,In_5);
and U2228 (N_2228,In_346,In_240);
nor U2229 (N_2229,In_545,In_246);
nand U2230 (N_2230,In_149,In_331);
nor U2231 (N_2231,In_49,In_678);
xnor U2232 (N_2232,In_59,In_23);
and U2233 (N_2233,In_437,In_665);
nand U2234 (N_2234,In_694,In_426);
nand U2235 (N_2235,In_748,In_425);
and U2236 (N_2236,In_485,In_677);
or U2237 (N_2237,In_539,In_742);
or U2238 (N_2238,In_554,In_150);
nand U2239 (N_2239,In_157,In_473);
nand U2240 (N_2240,In_90,In_647);
nand U2241 (N_2241,In_4,In_146);
or U2242 (N_2242,In_271,In_108);
or U2243 (N_2243,In_277,In_233);
and U2244 (N_2244,In_598,In_544);
or U2245 (N_2245,In_466,In_322);
nand U2246 (N_2246,In_732,In_446);
nand U2247 (N_2247,In_66,In_691);
and U2248 (N_2248,In_631,In_274);
or U2249 (N_2249,In_420,In_87);
nand U2250 (N_2250,In_311,In_289);
or U2251 (N_2251,In_413,In_444);
or U2252 (N_2252,In_21,In_72);
or U2253 (N_2253,In_5,In_69);
or U2254 (N_2254,In_145,In_147);
and U2255 (N_2255,In_339,In_691);
nor U2256 (N_2256,In_663,In_156);
nand U2257 (N_2257,In_196,In_472);
or U2258 (N_2258,In_597,In_262);
nand U2259 (N_2259,In_557,In_525);
and U2260 (N_2260,In_506,In_37);
nand U2261 (N_2261,In_300,In_195);
nor U2262 (N_2262,In_292,In_128);
nand U2263 (N_2263,In_15,In_258);
nand U2264 (N_2264,In_141,In_538);
nor U2265 (N_2265,In_377,In_223);
or U2266 (N_2266,In_17,In_223);
and U2267 (N_2267,In_181,In_635);
nand U2268 (N_2268,In_296,In_484);
nor U2269 (N_2269,In_237,In_33);
and U2270 (N_2270,In_558,In_278);
nand U2271 (N_2271,In_443,In_359);
nand U2272 (N_2272,In_569,In_161);
nor U2273 (N_2273,In_95,In_371);
or U2274 (N_2274,In_398,In_449);
and U2275 (N_2275,In_619,In_666);
nor U2276 (N_2276,In_481,In_677);
and U2277 (N_2277,In_143,In_266);
and U2278 (N_2278,In_739,In_734);
nand U2279 (N_2279,In_245,In_749);
or U2280 (N_2280,In_616,In_344);
nor U2281 (N_2281,In_106,In_693);
nand U2282 (N_2282,In_670,In_396);
or U2283 (N_2283,In_475,In_611);
nor U2284 (N_2284,In_723,In_621);
nand U2285 (N_2285,In_331,In_85);
and U2286 (N_2286,In_31,In_281);
and U2287 (N_2287,In_203,In_706);
and U2288 (N_2288,In_207,In_112);
and U2289 (N_2289,In_689,In_286);
or U2290 (N_2290,In_233,In_433);
or U2291 (N_2291,In_244,In_156);
or U2292 (N_2292,In_63,In_428);
and U2293 (N_2293,In_41,In_10);
nand U2294 (N_2294,In_39,In_338);
nand U2295 (N_2295,In_446,In_337);
and U2296 (N_2296,In_656,In_624);
nor U2297 (N_2297,In_497,In_557);
nand U2298 (N_2298,In_425,In_484);
or U2299 (N_2299,In_228,In_93);
and U2300 (N_2300,In_124,In_272);
and U2301 (N_2301,In_692,In_744);
nor U2302 (N_2302,In_681,In_2);
nor U2303 (N_2303,In_677,In_138);
nand U2304 (N_2304,In_15,In_483);
and U2305 (N_2305,In_502,In_272);
nor U2306 (N_2306,In_73,In_486);
nor U2307 (N_2307,In_482,In_28);
and U2308 (N_2308,In_162,In_166);
or U2309 (N_2309,In_208,In_89);
nand U2310 (N_2310,In_415,In_30);
nand U2311 (N_2311,In_232,In_661);
and U2312 (N_2312,In_337,In_388);
and U2313 (N_2313,In_232,In_662);
and U2314 (N_2314,In_23,In_108);
or U2315 (N_2315,In_635,In_676);
and U2316 (N_2316,In_325,In_42);
and U2317 (N_2317,In_58,In_214);
nor U2318 (N_2318,In_181,In_297);
or U2319 (N_2319,In_82,In_103);
nor U2320 (N_2320,In_237,In_638);
nand U2321 (N_2321,In_107,In_284);
nand U2322 (N_2322,In_139,In_736);
or U2323 (N_2323,In_127,In_285);
nor U2324 (N_2324,In_42,In_531);
nand U2325 (N_2325,In_376,In_77);
and U2326 (N_2326,In_547,In_603);
nand U2327 (N_2327,In_78,In_72);
nand U2328 (N_2328,In_444,In_188);
nand U2329 (N_2329,In_426,In_199);
nand U2330 (N_2330,In_424,In_68);
and U2331 (N_2331,In_561,In_658);
nand U2332 (N_2332,In_371,In_174);
and U2333 (N_2333,In_335,In_163);
nor U2334 (N_2334,In_261,In_733);
nor U2335 (N_2335,In_25,In_510);
nand U2336 (N_2336,In_378,In_387);
or U2337 (N_2337,In_672,In_228);
nor U2338 (N_2338,In_337,In_620);
xor U2339 (N_2339,In_38,In_211);
nand U2340 (N_2340,In_241,In_463);
or U2341 (N_2341,In_348,In_458);
or U2342 (N_2342,In_492,In_17);
nor U2343 (N_2343,In_482,In_466);
or U2344 (N_2344,In_749,In_118);
and U2345 (N_2345,In_715,In_684);
nor U2346 (N_2346,In_516,In_196);
nor U2347 (N_2347,In_525,In_2);
or U2348 (N_2348,In_699,In_362);
or U2349 (N_2349,In_562,In_283);
and U2350 (N_2350,In_60,In_571);
nand U2351 (N_2351,In_345,In_240);
or U2352 (N_2352,In_422,In_239);
nand U2353 (N_2353,In_91,In_688);
nand U2354 (N_2354,In_58,In_33);
nor U2355 (N_2355,In_267,In_317);
nor U2356 (N_2356,In_227,In_206);
or U2357 (N_2357,In_384,In_302);
nand U2358 (N_2358,In_436,In_557);
or U2359 (N_2359,In_701,In_380);
or U2360 (N_2360,In_372,In_517);
nand U2361 (N_2361,In_67,In_514);
nand U2362 (N_2362,In_347,In_232);
nand U2363 (N_2363,In_681,In_260);
and U2364 (N_2364,In_700,In_742);
or U2365 (N_2365,In_285,In_617);
nand U2366 (N_2366,In_251,In_617);
nor U2367 (N_2367,In_390,In_32);
or U2368 (N_2368,In_634,In_460);
nand U2369 (N_2369,In_486,In_454);
or U2370 (N_2370,In_502,In_106);
or U2371 (N_2371,In_353,In_69);
and U2372 (N_2372,In_130,In_154);
and U2373 (N_2373,In_327,In_234);
and U2374 (N_2374,In_507,In_573);
nand U2375 (N_2375,In_80,In_497);
and U2376 (N_2376,In_475,In_409);
nor U2377 (N_2377,In_715,In_613);
nand U2378 (N_2378,In_420,In_718);
or U2379 (N_2379,In_466,In_160);
and U2380 (N_2380,In_369,In_356);
nand U2381 (N_2381,In_115,In_226);
nand U2382 (N_2382,In_404,In_161);
nand U2383 (N_2383,In_196,In_648);
nand U2384 (N_2384,In_532,In_381);
or U2385 (N_2385,In_639,In_454);
or U2386 (N_2386,In_225,In_350);
nand U2387 (N_2387,In_690,In_604);
and U2388 (N_2388,In_375,In_692);
and U2389 (N_2389,In_286,In_27);
or U2390 (N_2390,In_142,In_3);
and U2391 (N_2391,In_456,In_475);
nor U2392 (N_2392,In_71,In_207);
or U2393 (N_2393,In_597,In_9);
xor U2394 (N_2394,In_131,In_732);
nand U2395 (N_2395,In_564,In_445);
and U2396 (N_2396,In_716,In_257);
and U2397 (N_2397,In_428,In_452);
or U2398 (N_2398,In_138,In_152);
nor U2399 (N_2399,In_536,In_621);
or U2400 (N_2400,In_189,In_712);
or U2401 (N_2401,In_243,In_245);
nand U2402 (N_2402,In_183,In_99);
or U2403 (N_2403,In_29,In_568);
nand U2404 (N_2404,In_287,In_0);
nand U2405 (N_2405,In_113,In_588);
or U2406 (N_2406,In_741,In_584);
and U2407 (N_2407,In_632,In_447);
nand U2408 (N_2408,In_176,In_548);
and U2409 (N_2409,In_694,In_582);
or U2410 (N_2410,In_438,In_638);
nand U2411 (N_2411,In_156,In_729);
nor U2412 (N_2412,In_625,In_80);
nor U2413 (N_2413,In_360,In_401);
and U2414 (N_2414,In_670,In_181);
and U2415 (N_2415,In_322,In_676);
or U2416 (N_2416,In_721,In_538);
and U2417 (N_2417,In_358,In_238);
nand U2418 (N_2418,In_202,In_171);
or U2419 (N_2419,In_604,In_243);
nor U2420 (N_2420,In_597,In_477);
and U2421 (N_2421,In_713,In_129);
or U2422 (N_2422,In_721,In_294);
nor U2423 (N_2423,In_269,In_339);
and U2424 (N_2424,In_725,In_639);
and U2425 (N_2425,In_582,In_384);
nand U2426 (N_2426,In_383,In_480);
or U2427 (N_2427,In_122,In_637);
nor U2428 (N_2428,In_483,In_438);
and U2429 (N_2429,In_702,In_324);
or U2430 (N_2430,In_455,In_436);
and U2431 (N_2431,In_726,In_374);
nor U2432 (N_2432,In_28,In_328);
nor U2433 (N_2433,In_412,In_220);
and U2434 (N_2434,In_510,In_281);
and U2435 (N_2435,In_646,In_278);
or U2436 (N_2436,In_158,In_643);
or U2437 (N_2437,In_635,In_470);
nand U2438 (N_2438,In_557,In_279);
nor U2439 (N_2439,In_734,In_173);
xor U2440 (N_2440,In_555,In_669);
or U2441 (N_2441,In_509,In_707);
xor U2442 (N_2442,In_639,In_254);
or U2443 (N_2443,In_265,In_701);
or U2444 (N_2444,In_696,In_339);
or U2445 (N_2445,In_625,In_437);
or U2446 (N_2446,In_32,In_387);
or U2447 (N_2447,In_152,In_460);
and U2448 (N_2448,In_308,In_408);
nand U2449 (N_2449,In_513,In_643);
nand U2450 (N_2450,In_77,In_44);
and U2451 (N_2451,In_43,In_417);
or U2452 (N_2452,In_54,In_22);
nand U2453 (N_2453,In_676,In_186);
or U2454 (N_2454,In_289,In_366);
nor U2455 (N_2455,In_445,In_194);
nand U2456 (N_2456,In_258,In_129);
xnor U2457 (N_2457,In_250,In_234);
and U2458 (N_2458,In_58,In_153);
and U2459 (N_2459,In_33,In_315);
nand U2460 (N_2460,In_139,In_534);
nand U2461 (N_2461,In_632,In_126);
nor U2462 (N_2462,In_586,In_689);
nand U2463 (N_2463,In_137,In_177);
or U2464 (N_2464,In_326,In_622);
or U2465 (N_2465,In_129,In_680);
nand U2466 (N_2466,In_252,In_580);
nor U2467 (N_2467,In_77,In_567);
and U2468 (N_2468,In_442,In_456);
nand U2469 (N_2469,In_425,In_376);
nor U2470 (N_2470,In_306,In_745);
or U2471 (N_2471,In_134,In_490);
or U2472 (N_2472,In_536,In_661);
nand U2473 (N_2473,In_464,In_660);
and U2474 (N_2474,In_648,In_515);
or U2475 (N_2475,In_244,In_505);
nand U2476 (N_2476,In_471,In_41);
nand U2477 (N_2477,In_246,In_350);
nor U2478 (N_2478,In_555,In_326);
nand U2479 (N_2479,In_442,In_489);
and U2480 (N_2480,In_533,In_113);
or U2481 (N_2481,In_414,In_459);
nand U2482 (N_2482,In_421,In_138);
xor U2483 (N_2483,In_221,In_678);
nand U2484 (N_2484,In_747,In_484);
nor U2485 (N_2485,In_7,In_655);
nand U2486 (N_2486,In_617,In_75);
nand U2487 (N_2487,In_618,In_122);
or U2488 (N_2488,In_28,In_632);
or U2489 (N_2489,In_371,In_299);
nand U2490 (N_2490,In_480,In_226);
nand U2491 (N_2491,In_496,In_667);
and U2492 (N_2492,In_414,In_27);
nor U2493 (N_2493,In_679,In_29);
and U2494 (N_2494,In_209,In_692);
nor U2495 (N_2495,In_388,In_505);
nor U2496 (N_2496,In_686,In_433);
nor U2497 (N_2497,In_387,In_498);
nor U2498 (N_2498,In_92,In_143);
or U2499 (N_2499,In_670,In_50);
nand U2500 (N_2500,N_404,N_2487);
and U2501 (N_2501,N_57,N_1259);
or U2502 (N_2502,N_1725,N_1606);
nand U2503 (N_2503,N_1336,N_1840);
and U2504 (N_2504,N_860,N_1838);
and U2505 (N_2505,N_2410,N_2196);
or U2506 (N_2506,N_966,N_2046);
or U2507 (N_2507,N_1181,N_2469);
nor U2508 (N_2508,N_241,N_1534);
nand U2509 (N_2509,N_1392,N_1962);
and U2510 (N_2510,N_1236,N_1868);
nor U2511 (N_2511,N_379,N_1282);
nand U2512 (N_2512,N_1496,N_1679);
nor U2513 (N_2513,N_1803,N_1950);
nor U2514 (N_2514,N_1576,N_1035);
and U2515 (N_2515,N_1034,N_2147);
or U2516 (N_2516,N_957,N_919);
or U2517 (N_2517,N_485,N_1712);
nand U2518 (N_2518,N_285,N_1190);
or U2519 (N_2519,N_614,N_1493);
nor U2520 (N_2520,N_1425,N_475);
nor U2521 (N_2521,N_1951,N_774);
nand U2522 (N_2522,N_984,N_708);
nand U2523 (N_2523,N_374,N_1882);
or U2524 (N_2524,N_1001,N_1571);
or U2525 (N_2525,N_2260,N_415);
nand U2526 (N_2526,N_837,N_625);
or U2527 (N_2527,N_93,N_1203);
nand U2528 (N_2528,N_1912,N_1981);
and U2529 (N_2529,N_1033,N_1498);
nor U2530 (N_2530,N_1697,N_272);
nor U2531 (N_2531,N_1941,N_1457);
nand U2532 (N_2532,N_200,N_540);
nor U2533 (N_2533,N_1660,N_1583);
nand U2534 (N_2534,N_399,N_1573);
and U2535 (N_2535,N_868,N_740);
or U2536 (N_2536,N_491,N_390);
or U2537 (N_2537,N_353,N_1161);
or U2538 (N_2538,N_883,N_6);
nor U2539 (N_2539,N_1351,N_1813);
and U2540 (N_2540,N_195,N_891);
nor U2541 (N_2541,N_842,N_401);
nor U2542 (N_2542,N_1329,N_1330);
nor U2543 (N_2543,N_2128,N_977);
or U2544 (N_2544,N_1672,N_2398);
or U2545 (N_2545,N_1323,N_1316);
or U2546 (N_2546,N_403,N_1286);
nand U2547 (N_2547,N_1475,N_739);
nand U2548 (N_2548,N_287,N_2471);
and U2549 (N_2549,N_554,N_1921);
nor U2550 (N_2550,N_313,N_1260);
and U2551 (N_2551,N_203,N_259);
nand U2552 (N_2552,N_566,N_2268);
or U2553 (N_2553,N_2276,N_278);
and U2554 (N_2554,N_1225,N_1165);
and U2555 (N_2555,N_1986,N_1271);
or U2556 (N_2556,N_1757,N_1961);
or U2557 (N_2557,N_25,N_1807);
and U2558 (N_2558,N_201,N_667);
or U2559 (N_2559,N_2430,N_603);
nand U2560 (N_2560,N_1238,N_653);
nor U2561 (N_2561,N_2053,N_516);
and U2562 (N_2562,N_1875,N_744);
nand U2563 (N_2563,N_443,N_2238);
or U2564 (N_2564,N_691,N_1845);
or U2565 (N_2565,N_388,N_1949);
or U2566 (N_2566,N_1309,N_198);
or U2567 (N_2567,N_1758,N_196);
and U2568 (N_2568,N_2373,N_2176);
xnor U2569 (N_2569,N_1189,N_1107);
nor U2570 (N_2570,N_2458,N_1406);
nand U2571 (N_2571,N_649,N_1526);
or U2572 (N_2572,N_1704,N_146);
or U2573 (N_2573,N_288,N_2381);
or U2574 (N_2574,N_787,N_383);
or U2575 (N_2575,N_1497,N_2250);
and U2576 (N_2576,N_32,N_1814);
and U2577 (N_2577,N_127,N_1995);
or U2578 (N_2578,N_116,N_2033);
or U2579 (N_2579,N_141,N_1081);
or U2580 (N_2580,N_326,N_757);
nand U2581 (N_2581,N_188,N_309);
xor U2582 (N_2582,N_1549,N_2026);
nand U2583 (N_2583,N_750,N_997);
nor U2584 (N_2584,N_2467,N_901);
nand U2585 (N_2585,N_1842,N_1415);
nand U2586 (N_2586,N_1111,N_1993);
xnor U2587 (N_2587,N_257,N_1088);
or U2588 (N_2588,N_477,N_946);
or U2589 (N_2589,N_1927,N_1918);
nor U2590 (N_2590,N_1249,N_1796);
nor U2591 (N_2591,N_441,N_1452);
xor U2592 (N_2592,N_1263,N_1825);
or U2593 (N_2593,N_1974,N_1418);
and U2594 (N_2594,N_2474,N_2479);
xor U2595 (N_2595,N_1861,N_445);
and U2596 (N_2596,N_2424,N_145);
or U2597 (N_2597,N_2329,N_50);
nand U2598 (N_2598,N_1117,N_980);
nor U2599 (N_2599,N_931,N_865);
nand U2600 (N_2600,N_847,N_599);
and U2601 (N_2601,N_2334,N_1503);
nor U2602 (N_2602,N_478,N_1850);
and U2603 (N_2603,N_1182,N_1970);
nand U2604 (N_2604,N_1664,N_1387);
nor U2605 (N_2605,N_297,N_437);
nand U2606 (N_2606,N_1087,N_1090);
nor U2607 (N_2607,N_674,N_216);
or U2608 (N_2608,N_1944,N_2378);
and U2609 (N_2609,N_1829,N_1805);
and U2610 (N_2610,N_1036,N_2435);
and U2611 (N_2611,N_1155,N_1565);
or U2612 (N_2612,N_92,N_1653);
nor U2613 (N_2613,N_2438,N_2486);
nand U2614 (N_2614,N_514,N_579);
nor U2615 (N_2615,N_1501,N_2376);
nand U2616 (N_2616,N_2210,N_395);
and U2617 (N_2617,N_1240,N_1340);
nor U2618 (N_2618,N_1625,N_2083);
and U2619 (N_2619,N_459,N_2194);
nor U2620 (N_2620,N_2375,N_2072);
nand U2621 (N_2621,N_2024,N_1032);
nand U2622 (N_2622,N_206,N_1585);
or U2623 (N_2623,N_397,N_1208);
nand U2624 (N_2624,N_2167,N_41);
nor U2625 (N_2625,N_113,N_1328);
nand U2626 (N_2626,N_1700,N_1063);
and U2627 (N_2627,N_1278,N_726);
and U2628 (N_2628,N_2264,N_684);
or U2629 (N_2629,N_1643,N_2068);
nand U2630 (N_2630,N_2237,N_882);
xor U2631 (N_2631,N_245,N_2456);
nand U2632 (N_2632,N_1654,N_271);
or U2633 (N_2633,N_381,N_451);
and U2634 (N_2634,N_2013,N_557);
and U2635 (N_2635,N_2137,N_1742);
nand U2636 (N_2636,N_1135,N_607);
nor U2637 (N_2637,N_1280,N_157);
nand U2638 (N_2638,N_1547,N_930);
or U2639 (N_2639,N_1202,N_1051);
nand U2640 (N_2640,N_1505,N_2001);
nor U2641 (N_2641,N_2234,N_2213);
or U2642 (N_2642,N_1123,N_2222);
nand U2643 (N_2643,N_1557,N_192);
and U2644 (N_2644,N_1586,N_2230);
nand U2645 (N_2645,N_150,N_519);
nand U2646 (N_2646,N_1297,N_1258);
and U2647 (N_2647,N_227,N_1535);
and U2648 (N_2648,N_43,N_732);
or U2649 (N_2649,N_626,N_2014);
and U2650 (N_2650,N_235,N_633);
or U2651 (N_2651,N_2223,N_1228);
or U2652 (N_2652,N_1568,N_851);
and U2653 (N_2653,N_831,N_844);
and U2654 (N_2654,N_764,N_1183);
and U2655 (N_2655,N_29,N_511);
nand U2656 (N_2656,N_1989,N_143);
or U2657 (N_2657,N_1396,N_2322);
and U2658 (N_2658,N_2172,N_52);
or U2659 (N_2659,N_595,N_1478);
nor U2660 (N_2660,N_564,N_698);
and U2661 (N_2661,N_887,N_2047);
and U2662 (N_2662,N_1613,N_593);
and U2663 (N_2663,N_623,N_2121);
or U2664 (N_2664,N_1611,N_904);
nor U2665 (N_2665,N_710,N_843);
and U2666 (N_2666,N_2008,N_1969);
and U2667 (N_2667,N_1551,N_87);
nand U2668 (N_2668,N_1633,N_2226);
and U2669 (N_2669,N_1647,N_527);
nor U2670 (N_2670,N_2212,N_719);
and U2671 (N_2671,N_746,N_2272);
nand U2672 (N_2672,N_1693,N_107);
nor U2673 (N_2673,N_1640,N_2459);
nand U2674 (N_2674,N_23,N_1164);
and U2675 (N_2675,N_1844,N_2231);
or U2676 (N_2676,N_853,N_17);
or U2677 (N_2677,N_1579,N_2245);
xor U2678 (N_2678,N_1076,N_2233);
and U2679 (N_2679,N_2342,N_2299);
nand U2680 (N_2680,N_2021,N_2484);
and U2681 (N_2681,N_2155,N_306);
and U2682 (N_2682,N_1283,N_812);
nor U2683 (N_2683,N_2045,N_2058);
and U2684 (N_2684,N_522,N_1809);
nand U2685 (N_2685,N_102,N_1116);
and U2686 (N_2686,N_2490,N_1686);
nor U2687 (N_2687,N_469,N_250);
or U2688 (N_2688,N_590,N_1652);
or U2689 (N_2689,N_2399,N_622);
or U2690 (N_2690,N_1602,N_1744);
or U2691 (N_2691,N_2071,N_442);
nand U2692 (N_2692,N_1147,N_1403);
nand U2693 (N_2693,N_1121,N_422);
nand U2694 (N_2694,N_1455,N_1086);
nor U2695 (N_2695,N_126,N_1901);
or U2696 (N_2696,N_1100,N_1341);
nor U2697 (N_2697,N_261,N_1619);
nor U2698 (N_2698,N_551,N_1473);
nor U2699 (N_2699,N_1562,N_103);
or U2700 (N_2700,N_1192,N_1674);
nor U2701 (N_2701,N_2078,N_1818);
nand U2702 (N_2702,N_2380,N_211);
nor U2703 (N_2703,N_2044,N_480);
and U2704 (N_2704,N_301,N_1622);
or U2705 (N_2705,N_717,N_2158);
nand U2706 (N_2706,N_1847,N_2029);
nand U2707 (N_2707,N_1936,N_528);
or U2708 (N_2708,N_168,N_2428);
nor U2709 (N_2709,N_1866,N_97);
or U2710 (N_2710,N_1062,N_1026);
or U2711 (N_2711,N_2187,N_800);
and U2712 (N_2712,N_269,N_926);
nand U2713 (N_2713,N_149,N_42);
and U2714 (N_2714,N_391,N_542);
and U2715 (N_2715,N_118,N_219);
nand U2716 (N_2716,N_55,N_239);
nor U2717 (N_2717,N_888,N_923);
and U2718 (N_2718,N_2280,N_2449);
and U2719 (N_2719,N_2270,N_819);
or U2720 (N_2720,N_2414,N_2081);
and U2721 (N_2721,N_61,N_902);
nand U2722 (N_2722,N_1637,N_440);
nand U2723 (N_2723,N_507,N_1281);
or U2724 (N_2724,N_840,N_988);
and U2725 (N_2725,N_181,N_735);
and U2726 (N_2726,N_1400,N_2447);
nor U2727 (N_2727,N_1293,N_2023);
and U2728 (N_2728,N_1287,N_1359);
and U2729 (N_2729,N_348,N_2207);
nand U2730 (N_2730,N_86,N_1792);
nand U2731 (N_2731,N_2110,N_2478);
nor U2732 (N_2732,N_1605,N_1886);
nor U2733 (N_2733,N_2279,N_1559);
nand U2734 (N_2734,N_1734,N_2472);
nand U2735 (N_2735,N_518,N_1003);
or U2736 (N_2736,N_985,N_1030);
and U2737 (N_2737,N_1662,N_334);
nand U2738 (N_2738,N_1333,N_1234);
xor U2739 (N_2739,N_363,N_417);
nor U2740 (N_2740,N_2154,N_1934);
nor U2741 (N_2741,N_1657,N_2096);
or U2742 (N_2742,N_2437,N_798);
nor U2743 (N_2743,N_1315,N_2303);
or U2744 (N_2744,N_472,N_1851);
nor U2745 (N_2745,N_2117,N_26);
and U2746 (N_2746,N_311,N_171);
nor U2747 (N_2747,N_138,N_315);
and U2748 (N_2748,N_1148,N_1617);
or U2749 (N_2749,N_749,N_700);
nand U2750 (N_2750,N_394,N_1491);
and U2751 (N_2751,N_2057,N_747);
nor U2752 (N_2752,N_925,N_1587);
xor U2753 (N_2753,N_2174,N_736);
nand U2754 (N_2754,N_1958,N_742);
and U2755 (N_2755,N_1867,N_2114);
and U2756 (N_2756,N_2049,N_1869);
nor U2757 (N_2757,N_166,N_1506);
and U2758 (N_2758,N_263,N_2099);
nand U2759 (N_2759,N_598,N_120);
nand U2760 (N_2760,N_2291,N_2002);
and U2761 (N_2761,N_811,N_1320);
nor U2762 (N_2762,N_2042,N_1764);
and U2763 (N_2763,N_2217,N_1154);
nor U2764 (N_2764,N_21,N_457);
nor U2765 (N_2765,N_1171,N_1675);
nor U2766 (N_2766,N_416,N_45);
nand U2767 (N_2767,N_1275,N_1344);
and U2768 (N_2768,N_1537,N_252);
or U2769 (N_2769,N_1865,N_1130);
nand U2770 (N_2770,N_1273,N_1760);
or U2771 (N_2771,N_961,N_367);
nor U2772 (N_2772,N_897,N_1381);
nor U2773 (N_2773,N_836,N_729);
nand U2774 (N_2774,N_2211,N_1159);
or U2775 (N_2775,N_796,N_657);
or U2776 (N_2776,N_382,N_771);
and U2777 (N_2777,N_461,N_734);
or U2778 (N_2778,N_1857,N_2448);
or U2779 (N_2779,N_58,N_577);
nand U2780 (N_2780,N_1823,N_1940);
or U2781 (N_2781,N_642,N_1288);
and U2782 (N_2782,N_123,N_2336);
or U2783 (N_2783,N_380,N_1773);
nand U2784 (N_2784,N_669,N_830);
and U2785 (N_2785,N_702,N_1984);
and U2786 (N_2786,N_918,N_944);
and U2787 (N_2787,N_2499,N_1820);
or U2788 (N_2788,N_1476,N_2221);
nor U2789 (N_2789,N_1431,N_2360);
nor U2790 (N_2790,N_1569,N_1916);
or U2791 (N_2791,N_106,N_779);
and U2792 (N_2792,N_1919,N_652);
nor U2793 (N_2793,N_2161,N_484);
nand U2794 (N_2794,N_7,N_164);
and U2795 (N_2795,N_2050,N_778);
nand U2796 (N_2796,N_1952,N_371);
or U2797 (N_2797,N_654,N_1310);
nand U2798 (N_2798,N_454,N_1474);
nor U2799 (N_2799,N_1331,N_619);
nor U2800 (N_2800,N_1701,N_857);
nand U2801 (N_2801,N_1061,N_142);
nand U2802 (N_2802,N_2417,N_1544);
xor U2803 (N_2803,N_576,N_1489);
nand U2804 (N_2804,N_1759,N_1313);
nand U2805 (N_2805,N_597,N_1614);
or U2806 (N_2806,N_979,N_378);
nand U2807 (N_2807,N_1930,N_1736);
and U2808 (N_2808,N_2027,N_180);
nor U2809 (N_2809,N_723,N_1705);
nand U2810 (N_2810,N_1976,N_2007);
nor U2811 (N_2811,N_572,N_2111);
or U2812 (N_2812,N_1364,N_2298);
or U2813 (N_2813,N_13,N_2020);
nand U2814 (N_2814,N_741,N_1118);
nor U2815 (N_2815,N_591,N_1824);
and U2816 (N_2816,N_638,N_72);
xor U2817 (N_2817,N_2089,N_68);
and U2818 (N_2818,N_238,N_1389);
nand U2819 (N_2819,N_162,N_1279);
and U2820 (N_2820,N_1651,N_2040);
and U2821 (N_2821,N_2331,N_234);
nor U2822 (N_2822,N_648,N_724);
and U2823 (N_2823,N_1427,N_1133);
and U2824 (N_2824,N_1956,N_360);
nor U2825 (N_2825,N_872,N_2318);
nand U2826 (N_2826,N_718,N_2429);
or U2827 (N_2827,N_254,N_1768);
nand U2828 (N_2828,N_680,N_587);
and U2829 (N_2829,N_1327,N_498);
nand U2830 (N_2830,N_1482,N_2374);
xor U2831 (N_2831,N_2177,N_1639);
nand U2832 (N_2832,N_1401,N_2135);
and U2833 (N_2833,N_545,N_1567);
or U2834 (N_2834,N_2080,N_538);
nand U2835 (N_2835,N_810,N_1750);
nor U2836 (N_2836,N_2030,N_1306);
or U2837 (N_2837,N_1852,N_1987);
or U2838 (N_2838,N_1447,N_2289);
nand U2839 (N_2839,N_1516,N_3);
and U2840 (N_2840,N_1991,N_350);
nand U2841 (N_2841,N_460,N_1488);
and U2842 (N_2842,N_1881,N_1718);
nand U2843 (N_2843,N_2444,N_1906);
nand U2844 (N_2844,N_2084,N_999);
and U2845 (N_2845,N_547,N_1676);
nand U2846 (N_2846,N_682,N_1015);
nand U2847 (N_2847,N_1379,N_410);
and U2848 (N_2848,N_679,N_232);
and U2849 (N_2849,N_1307,N_333);
or U2850 (N_2850,N_549,N_273);
and U2851 (N_2851,N_773,N_1685);
nand U2852 (N_2852,N_920,N_64);
or U2853 (N_2853,N_1141,N_167);
nand U2854 (N_2854,N_1769,N_2141);
nor U2855 (N_2855,N_2018,N_1683);
nor U2856 (N_2856,N_71,N_1859);
nor U2857 (N_2857,N_993,N_1348);
or U2858 (N_2858,N_949,N_956);
nor U2859 (N_2859,N_1413,N_81);
and U2860 (N_2860,N_16,N_1284);
nor U2861 (N_2861,N_1767,N_2288);
and U2862 (N_2862,N_1276,N_2338);
nor U2863 (N_2863,N_660,N_10);
xor U2864 (N_2864,N_807,N_1385);
or U2865 (N_2865,N_1603,N_1853);
or U2866 (N_2866,N_2395,N_2178);
nor U2867 (N_2867,N_637,N_242);
xor U2868 (N_2868,N_2139,N_1053);
nor U2869 (N_2869,N_1515,N_1082);
or U2870 (N_2870,N_1655,N_148);
or U2871 (N_2871,N_606,N_1717);
xnor U2872 (N_2872,N_74,N_848);
and U2873 (N_2873,N_121,N_1907);
or U2874 (N_2874,N_222,N_1084);
nand U2875 (N_2875,N_659,N_389);
nor U2876 (N_2876,N_124,N_1968);
nor U2877 (N_2877,N_1541,N_229);
nand U2878 (N_2878,N_1908,N_2418);
nor U2879 (N_2879,N_277,N_2060);
nor U2880 (N_2880,N_2372,N_1746);
nand U2881 (N_2881,N_1898,N_1593);
or U2882 (N_2882,N_228,N_2235);
and U2883 (N_2883,N_613,N_435);
or U2884 (N_2884,N_789,N_361);
nor U2885 (N_2885,N_1270,N_2498);
and U2886 (N_2886,N_1826,N_1714);
nand U2887 (N_2887,N_2074,N_2097);
xnor U2888 (N_2888,N_2152,N_1325);
nand U2889 (N_2889,N_1884,N_2411);
and U2890 (N_2890,N_291,N_1375);
nand U2891 (N_2891,N_1103,N_1180);
nor U2892 (N_2892,N_553,N_400);
nand U2893 (N_2893,N_687,N_51);
nand U2894 (N_2894,N_2457,N_1608);
nand U2895 (N_2895,N_2256,N_1913);
or U2896 (N_2896,N_1358,N_1132);
and U2897 (N_2897,N_1903,N_1391);
or U2898 (N_2898,N_621,N_1377);
nand U2899 (N_2899,N_2202,N_447);
and U2900 (N_2900,N_2287,N_2426);
and U2901 (N_2901,N_446,N_544);
xnor U2902 (N_2902,N_1440,N_989);
nor U2903 (N_2903,N_253,N_1518);
or U2904 (N_2904,N_713,N_1687);
nand U2905 (N_2905,N_1374,N_2006);
nand U2906 (N_2906,N_280,N_2366);
and U2907 (N_2907,N_1058,N_2214);
nor U2908 (N_2908,N_1176,N_0);
nor U2909 (N_2909,N_44,N_571);
nand U2910 (N_2910,N_300,N_1417);
nor U2911 (N_2911,N_2422,N_1253);
and U2912 (N_2912,N_678,N_405);
nand U2913 (N_2913,N_1011,N_1879);
and U2914 (N_2914,N_573,N_466);
xor U2915 (N_2915,N_2497,N_1963);
nand U2916 (N_2916,N_996,N_1665);
nor U2917 (N_2917,N_1638,N_335);
or U2918 (N_2918,N_790,N_983);
nand U2919 (N_2919,N_22,N_1612);
nor U2920 (N_2920,N_536,N_2286);
and U2921 (N_2921,N_938,N_1979);
or U2922 (N_2922,N_1029,N_801);
or U2923 (N_2923,N_2355,N_1193);
and U2924 (N_2924,N_817,N_650);
nor U2925 (N_2925,N_411,N_1716);
nor U2926 (N_2926,N_1289,N_1386);
or U2927 (N_2927,N_312,N_1771);
nand U2928 (N_2928,N_1129,N_1016);
nor U2929 (N_2929,N_1151,N_1302);
and U2930 (N_2930,N_432,N_1730);
or U2931 (N_2931,N_2156,N_1955);
and U2932 (N_2932,N_2065,N_47);
nor U2933 (N_2933,N_450,N_2170);
nor U2934 (N_2934,N_645,N_2452);
and U2935 (N_2935,N_1545,N_2239);
xor U2936 (N_2936,N_578,N_282);
or U2937 (N_2937,N_893,N_2339);
nand U2938 (N_2938,N_896,N_1412);
nand U2939 (N_2939,N_1739,N_497);
nor U2940 (N_2940,N_1831,N_1802);
or U2941 (N_2941,N_240,N_217);
or U2942 (N_2942,N_421,N_2382);
and U2943 (N_2943,N_1312,N_36);
and U2944 (N_2944,N_1223,N_2370);
nor U2945 (N_2945,N_1257,N_2048);
nor U2946 (N_2946,N_1982,N_592);
or U2947 (N_2947,N_2200,N_1460);
or U2948 (N_2948,N_1210,N_358);
or U2949 (N_2949,N_670,N_5);
and U2950 (N_2950,N_1115,N_1531);
nor U2951 (N_2951,N_1472,N_2341);
nor U2952 (N_2952,N_543,N_2052);
nand U2953 (N_2953,N_1343,N_1096);
and U2954 (N_2954,N_2224,N_1169);
nand U2955 (N_2955,N_1322,N_2009);
and U2956 (N_2956,N_210,N_1751);
nand U2957 (N_2957,N_1163,N_1504);
or U2958 (N_2958,N_1000,N_1841);
nand U2959 (N_2959,N_194,N_582);
nand U2960 (N_2960,N_1024,N_641);
and U2961 (N_2961,N_769,N_2189);
nand U2962 (N_2962,N_1661,N_1212);
or U2963 (N_2963,N_1980,N_531);
nand U2964 (N_2964,N_1409,N_2091);
nor U2965 (N_2965,N_1747,N_1079);
and U2966 (N_2966,N_636,N_586);
nand U2967 (N_2967,N_663,N_563);
nand U2968 (N_2968,N_186,N_2323);
nor U2969 (N_2969,N_398,N_38);
nor U2970 (N_2970,N_2282,N_1928);
nand U2971 (N_2971,N_683,N_274);
nand U2972 (N_2972,N_953,N_1360);
or U2973 (N_2973,N_513,N_125);
or U2974 (N_2974,N_347,N_418);
nor U2975 (N_2975,N_1226,N_2454);
nor U2976 (N_2976,N_1871,N_1698);
nor U2977 (N_2977,N_1815,N_1074);
or U2978 (N_2978,N_2462,N_244);
nor U2979 (N_2979,N_294,N_950);
nor U2980 (N_2980,N_1947,N_917);
or U2981 (N_2981,N_423,N_2340);
nor U2982 (N_2982,N_964,N_1337);
or U2983 (N_2983,N_721,N_731);
or U2984 (N_2984,N_1971,N_1205);
and U2985 (N_2985,N_1067,N_431);
or U2986 (N_2986,N_2168,N_829);
xor U2987 (N_2987,N_1513,N_1626);
or U2988 (N_2988,N_1218,N_799);
nand U2989 (N_2989,N_560,N_1383);
and U2990 (N_2990,N_927,N_1300);
nand U2991 (N_2991,N_2025,N_1996);
or U2992 (N_2992,N_960,N_304);
or U2993 (N_2993,N_2421,N_1862);
and U2994 (N_2994,N_2337,N_385);
and U2995 (N_2995,N_1581,N_1791);
and U2996 (N_2996,N_1694,N_1519);
nor U2997 (N_2997,N_295,N_1102);
or U2998 (N_2998,N_2227,N_1376);
nand U2999 (N_2999,N_618,N_1254);
nand U3000 (N_3000,N_644,N_1536);
nand U3001 (N_3001,N_791,N_962);
nand U3002 (N_3002,N_1156,N_369);
and U3003 (N_3003,N_412,N_1797);
and U3004 (N_3004,N_1338,N_805);
or U3005 (N_3005,N_2258,N_1992);
nor U3006 (N_3006,N_2283,N_1630);
nand U3007 (N_3007,N_783,N_444);
nor U3008 (N_3008,N_1816,N_711);
nor U3009 (N_3009,N_788,N_1217);
nor U3010 (N_3010,N_2451,N_170);
nand U3011 (N_3011,N_2144,N_804);
nor U3012 (N_3012,N_2393,N_2311);
nor U3013 (N_3013,N_2066,N_743);
nand U3014 (N_3014,N_2122,N_797);
nand U3015 (N_3015,N_1204,N_1774);
or U3016 (N_3016,N_900,N_1352);
nor U3017 (N_3017,N_1469,N_90);
and U3018 (N_3018,N_286,N_689);
and U3019 (N_3019,N_1932,N_2324);
and U3020 (N_3020,N_1729,N_2427);
and U3021 (N_3021,N_9,N_2357);
nand U3022 (N_3022,N_1889,N_187);
or U3023 (N_3023,N_2266,N_2293);
or U3024 (N_3024,N_2105,N_2326);
and U3025 (N_3025,N_2365,N_2138);
and U3026 (N_3026,N_2295,N_65);
nor U3027 (N_3027,N_1247,N_1524);
nor U3028 (N_3028,N_368,N_1658);
or U3029 (N_3029,N_890,N_174);
and U3030 (N_3030,N_1314,N_1911);
nand U3031 (N_3031,N_906,N_640);
or U3032 (N_3032,N_878,N_1104);
nand U3033 (N_3033,N_321,N_2095);
nor U3034 (N_3034,N_204,N_1858);
and U3035 (N_3035,N_226,N_354);
or U3036 (N_3036,N_534,N_79);
or U3037 (N_3037,N_488,N_2463);
nor U3038 (N_3038,N_1248,N_1542);
or U3039 (N_3039,N_2201,N_1398);
and U3040 (N_3040,N_990,N_777);
nor U3041 (N_3041,N_69,N_1883);
or U3042 (N_3042,N_1938,N_1663);
and U3043 (N_3043,N_193,N_1776);
or U3044 (N_3044,N_2252,N_96);
nor U3045 (N_3045,N_1727,N_948);
nand U3046 (N_3046,N_854,N_856);
or U3047 (N_3047,N_574,N_1502);
nor U3048 (N_3048,N_786,N_2229);
nand U3049 (N_3049,N_34,N_2208);
nor U3050 (N_3050,N_1239,N_190);
and U3051 (N_3051,N_2063,N_2285);
nand U3052 (N_3052,N_346,N_1766);
nor U3053 (N_3053,N_866,N_2085);
nor U3054 (N_3054,N_2003,N_561);
or U3055 (N_3055,N_503,N_1197);
or U3056 (N_3056,N_1167,N_1429);
nor U3057 (N_3057,N_822,N_2396);
or U3058 (N_3058,N_2255,N_1960);
nand U3059 (N_3059,N_2278,N_1269);
or U3060 (N_3060,N_2134,N_1010);
or U3061 (N_3061,N_359,N_78);
nor U3062 (N_3062,N_2402,N_1357);
or U3063 (N_3063,N_852,N_1828);
and U3064 (N_3064,N_1018,N_1623);
and U3065 (N_3065,N_1874,N_2169);
nor U3066 (N_3066,N_1353,N_982);
nand U3067 (N_3067,N_1810,N_1175);
nand U3068 (N_3068,N_2401,N_1483);
and U3069 (N_3069,N_1801,N_1463);
nor U3070 (N_3070,N_420,N_407);
nand U3071 (N_3071,N_1785,N_2394);
or U3072 (N_3072,N_762,N_594);
nor U3073 (N_3073,N_1356,N_1038);
nor U3074 (N_3074,N_2246,N_54);
nor U3075 (N_3075,N_482,N_1682);
and U3076 (N_3076,N_2219,N_676);
nand U3077 (N_3077,N_651,N_139);
nand U3078 (N_3078,N_1787,N_2436);
nor U3079 (N_3079,N_159,N_1339);
nor U3080 (N_3080,N_213,N_1411);
nand U3081 (N_3081,N_978,N_1789);
and U3082 (N_3082,N_14,N_1244);
nand U3083 (N_3083,N_1368,N_2460);
or U3084 (N_3084,N_2319,N_392);
xor U3085 (N_3085,N_994,N_1895);
nand U3086 (N_3086,N_688,N_1667);
or U3087 (N_3087,N_970,N_515);
or U3088 (N_3088,N_2113,N_508);
and U3089 (N_3089,N_655,N_1410);
nand U3090 (N_3090,N_728,N_429);
nor U3091 (N_3091,N_2317,N_1837);
nor U3092 (N_3092,N_1720,N_2408);
xor U3093 (N_3093,N_2489,N_104);
nor U3094 (N_3094,N_279,N_158);
and U3095 (N_3095,N_1948,N_1220);
or U3096 (N_3096,N_1237,N_2349);
and U3097 (N_3097,N_986,N_1347);
or U3098 (N_3098,N_2441,N_1106);
or U3099 (N_3099,N_991,N_1528);
nand U3100 (N_3100,N_317,N_1120);
or U3101 (N_3101,N_1540,N_1077);
xor U3102 (N_3102,N_2243,N_2308);
nand U3103 (N_3103,N_1763,N_951);
and U3104 (N_3104,N_1231,N_869);
or U3105 (N_3105,N_567,N_589);
or U3106 (N_3106,N_505,N_802);
or U3107 (N_3107,N_885,N_247);
nand U3108 (N_3108,N_1566,N_2351);
nand U3109 (N_3109,N_548,N_1670);
nor U3110 (N_3110,N_2102,N_751);
and U3111 (N_3111,N_1977,N_2082);
or U3112 (N_3112,N_176,N_1945);
and U3113 (N_3113,N_1125,N_2482);
and U3114 (N_3114,N_1438,N_1245);
nand U3115 (N_3115,N_828,N_387);
nor U3116 (N_3116,N_1201,N_1721);
or U3117 (N_3117,N_2358,N_877);
nand U3118 (N_3118,N_685,N_1935);
xor U3119 (N_3119,N_2362,N_892);
and U3120 (N_3120,N_2384,N_2124);
nand U3121 (N_3121,N_119,N_281);
nor U3122 (N_3122,N_153,N_1795);
nor U3123 (N_3123,N_2019,N_1066);
and U3124 (N_3124,N_1023,N_504);
nor U3125 (N_3125,N_1914,N_2445);
and U3126 (N_3126,N_1043,N_781);
nand U3127 (N_3127,N_2363,N_1572);
nand U3128 (N_3128,N_2251,N_2450);
nor U3129 (N_3129,N_889,N_316);
or U3130 (N_3130,N_1456,N_175);
and U3131 (N_3131,N_2242,N_647);
nor U3132 (N_3132,N_873,N_1085);
nor U3133 (N_3133,N_331,N_165);
xor U3134 (N_3134,N_1953,N_1091);
nand U3135 (N_3135,N_2185,N_1600);
xnor U3136 (N_3136,N_898,N_178);
nor U3137 (N_3137,N_2310,N_2269);
nor U3138 (N_3138,N_1681,N_2190);
or U3139 (N_3139,N_1964,N_870);
nand U3140 (N_3140,N_173,N_1168);
or U3141 (N_3141,N_2038,N_1246);
and U3142 (N_3142,N_2004,N_223);
nand U3143 (N_3143,N_681,N_1436);
xor U3144 (N_3144,N_2000,N_114);
nor U3145 (N_3145,N_1832,N_481);
and U3146 (N_3146,N_1500,N_2112);
nand U3147 (N_3147,N_70,N_1126);
nor U3148 (N_3148,N_464,N_1142);
and U3149 (N_3149,N_850,N_832);
nor U3150 (N_3150,N_324,N_1507);
xnor U3151 (N_3151,N_570,N_487);
and U3152 (N_3152,N_341,N_1349);
nor U3153 (N_3153,N_2193,N_2316);
and U3154 (N_3154,N_2132,N_1490);
nor U3155 (N_3155,N_1873,N_1527);
or U3156 (N_3156,N_813,N_763);
and U3157 (N_3157,N_998,N_2405);
and U3158 (N_3158,N_2348,N_486);
or U3159 (N_3159,N_129,N_1749);
or U3160 (N_3160,N_1185,N_1839);
nor U3161 (N_3161,N_2386,N_2016);
or U3162 (N_3162,N_2294,N_2145);
nor U3163 (N_3163,N_1607,N_1355);
nor U3164 (N_3164,N_2496,N_1435);
nand U3165 (N_3165,N_2088,N_2206);
and U3166 (N_3166,N_1049,N_191);
and U3167 (N_3167,N_2468,N_1394);
nand U3168 (N_3168,N_182,N_972);
nor U3169 (N_3169,N_895,N_1471);
nand U3170 (N_3170,N_1707,N_179);
and U3171 (N_3171,N_2069,N_1441);
nor U3172 (N_3172,N_1812,N_305);
and U3173 (N_3173,N_258,N_1574);
nor U3174 (N_3174,N_2171,N_974);
nor U3175 (N_3175,N_1532,N_1420);
nor U3176 (N_3176,N_2059,N_863);
or U3177 (N_3177,N_1743,N_2387);
nor U3178 (N_3178,N_1450,N_225);
nor U3179 (N_3179,N_1892,N_1421);
nand U3180 (N_3180,N_2476,N_929);
nor U3181 (N_3181,N_1775,N_1272);
nand U3182 (N_3182,N_100,N_1709);
and U3183 (N_3183,N_1596,N_1708);
nand U3184 (N_3184,N_163,N_376);
nand U3185 (N_3185,N_1779,N_1893);
nor U3186 (N_3186,N_1671,N_841);
nor U3187 (N_3187,N_2480,N_2146);
or U3188 (N_3188,N_677,N_134);
nor U3189 (N_3189,N_455,N_1629);
nand U3190 (N_3190,N_809,N_1041);
nor U3191 (N_3191,N_1924,N_565);
nor U3192 (N_3192,N_1134,N_634);
nand U3193 (N_3193,N_284,N_1520);
nand U3194 (N_3194,N_2182,N_2162);
nor U3195 (N_3195,N_220,N_1372);
and U3196 (N_3196,N_2086,N_343);
nand U3197 (N_3197,N_1031,N_532);
nand U3198 (N_3198,N_56,N_2130);
nor U3199 (N_3199,N_2404,N_1480);
nand U3200 (N_3200,N_2495,N_2120);
nor U3201 (N_3201,N_1618,N_342);
nand U3202 (N_3202,N_584,N_2271);
and U3203 (N_3203,N_754,N_707);
or U3204 (N_3204,N_1972,N_2254);
or U3205 (N_3205,N_1321,N_2216);
nand U3206 (N_3206,N_2263,N_199);
and U3207 (N_3207,N_2273,N_1399);
or U3208 (N_3208,N_1426,N_818);
nand U3209 (N_3209,N_617,N_1998);
and U3210 (N_3210,N_725,N_329);
or U3211 (N_3211,N_1556,N_1335);
nand U3212 (N_3212,N_1466,N_704);
or U3213 (N_3213,N_714,N_1213);
nor U3214 (N_3214,N_1380,N_696);
and U3215 (N_3215,N_2175,N_83);
nor U3216 (N_3216,N_1601,N_814);
and U3217 (N_3217,N_1199,N_473);
nand U3218 (N_3218,N_117,N_1703);
or U3219 (N_3219,N_517,N_1487);
nand U3220 (N_3220,N_1732,N_1174);
or U3221 (N_3221,N_35,N_2232);
xnor U3222 (N_3222,N_1099,N_600);
nor U3223 (N_3223,N_1691,N_1595);
or U3224 (N_3224,N_1136,N_2034);
nand U3225 (N_3225,N_609,N_2367);
nand U3226 (N_3226,N_1243,N_1885);
or U3227 (N_3227,N_2215,N_2332);
nand U3228 (N_3228,N_765,N_730);
and U3229 (N_3229,N_40,N_1966);
or U3230 (N_3230,N_356,N_1388);
nand U3231 (N_3231,N_209,N_2125);
and U3232 (N_3232,N_492,N_631);
and U3233 (N_3233,N_915,N_1728);
nor U3234 (N_3234,N_1646,N_434);
nand U3235 (N_3235,N_2415,N_89);
nand U3236 (N_3236,N_2356,N_656);
and U3237 (N_3237,N_1214,N_205);
and U3238 (N_3238,N_2064,N_1756);
and U3239 (N_3239,N_672,N_393);
nand U3240 (N_3240,N_427,N_884);
nor U3241 (N_3241,N_1509,N_115);
nor U3242 (N_3242,N_611,N_2153);
nand U3243 (N_3243,N_1207,N_2409);
xnor U3244 (N_3244,N_2151,N_1529);
nand U3245 (N_3245,N_583,N_496);
xnor U3246 (N_3246,N_1114,N_1177);
xor U3247 (N_3247,N_720,N_2181);
nand U3248 (N_3248,N_1187,N_275);
and U3249 (N_3249,N_1702,N_1461);
nand U3250 (N_3250,N_1929,N_775);
xnor U3251 (N_3251,N_493,N_963);
nand U3252 (N_3252,N_1632,N_1071);
and U3253 (N_3253,N_1110,N_30);
nor U3254 (N_3254,N_608,N_355);
nor U3255 (N_3255,N_952,N_1723);
or U3256 (N_3256,N_959,N_2247);
or U3257 (N_3257,N_2305,N_1468);
or U3258 (N_3258,N_233,N_2307);
or U3259 (N_3259,N_449,N_2123);
nand U3260 (N_3260,N_483,N_2192);
and U3261 (N_3261,N_2037,N_2012);
nor U3262 (N_3262,N_2118,N_99);
nand U3263 (N_3263,N_1097,N_1423);
nor U3264 (N_3264,N_1722,N_260);
or U3265 (N_3265,N_2180,N_1139);
or U3266 (N_3266,N_2166,N_1954);
nor U3267 (N_3267,N_1860,N_969);
nor U3268 (N_3268,N_1362,N_2440);
and U3269 (N_3269,N_1678,N_1609);
or U3270 (N_3270,N_2195,N_344);
and U3271 (N_3271,N_2056,N_351);
or U3272 (N_3272,N_2389,N_1404);
or U3273 (N_3273,N_1072,N_849);
nor U3274 (N_3274,N_803,N_2407);
and U3275 (N_3275,N_237,N_230);
or U3276 (N_3276,N_1817,N_699);
or U3277 (N_3277,N_2119,N_462);
nand U3278 (N_3278,N_701,N_112);
nand U3279 (N_3279,N_1990,N_825);
nand U3280 (N_3280,N_2108,N_1268);
or U3281 (N_3281,N_320,N_1459);
nand U3282 (N_3282,N_965,N_2425);
or U3283 (N_3283,N_1848,N_1370);
nand U3284 (N_3284,N_345,N_1827);
or U3285 (N_3285,N_2327,N_49);
or U3286 (N_3286,N_2364,N_471);
nor U3287 (N_3287,N_169,N_1052);
nor U3288 (N_3288,N_414,N_1706);
and U3289 (N_3289,N_635,N_1094);
nor U3290 (N_3290,N_2062,N_559);
and U3291 (N_3291,N_768,N_601);
and U3292 (N_3292,N_541,N_2354);
nand U3293 (N_3293,N_894,N_1946);
nand U3294 (N_3294,N_1872,N_1230);
nor U3295 (N_3295,N_1008,N_207);
xnor U3296 (N_3296,N_924,N_265);
and U3297 (N_3297,N_1146,N_1999);
and U3298 (N_3298,N_864,N_243);
nand U3299 (N_3299,N_1897,N_879);
nor U3300 (N_3300,N_1430,N_1888);
or U3301 (N_3301,N_761,N_755);
or U3302 (N_3302,N_1453,N_1870);
nand U3303 (N_3303,N_861,N_936);
nor U3304 (N_3304,N_512,N_874);
nor U3305 (N_3305,N_1311,N_73);
nor U3306 (N_3306,N_1724,N_795);
nand U3307 (N_3307,N_933,N_1449);
or U3308 (N_3308,N_1397,N_604);
or U3309 (N_3309,N_63,N_1037);
nand U3310 (N_3310,N_2203,N_1153);
nor U3311 (N_3311,N_2115,N_1692);
nand U3312 (N_3312,N_310,N_1224);
and U3313 (N_3313,N_1428,N_248);
nand U3314 (N_3314,N_1434,N_1393);
or U3315 (N_3315,N_1317,N_1846);
or U3316 (N_3316,N_1262,N_907);
xnor U3317 (N_3317,N_1162,N_823);
nor U3318 (N_3318,N_2361,N_1973);
nor U3319 (N_3319,N_643,N_876);
and U3320 (N_3320,N_2106,N_1318);
nor U3321 (N_3321,N_266,N_2079);
nor U3322 (N_3322,N_2149,N_2032);
and U3323 (N_3323,N_2352,N_1740);
or U3324 (N_3324,N_1462,N_2453);
or U3325 (N_3325,N_1836,N_1092);
and U3326 (N_3326,N_303,N_937);
nand U3327 (N_3327,N_2075,N_712);
nand U3328 (N_3328,N_1521,N_1046);
and U3329 (N_3329,N_88,N_1696);
nor U3330 (N_3330,N_846,N_1324);
nor U3331 (N_3331,N_256,N_2328);
and U3332 (N_3332,N_1628,N_37);
and U3333 (N_3333,N_386,N_1864);
nor U3334 (N_3334,N_533,N_59);
and U3335 (N_3335,N_1635,N_160);
nor U3336 (N_3336,N_575,N_867);
nand U3337 (N_3337,N_108,N_270);
or U3338 (N_3338,N_1508,N_1196);
and U3339 (N_3339,N_1184,N_675);
xor U3340 (N_3340,N_1552,N_585);
nand U3341 (N_3341,N_705,N_1382);
and U3342 (N_3342,N_2051,N_101);
and U3343 (N_3343,N_2236,N_154);
nor U3344 (N_3344,N_2244,N_1849);
nor U3345 (N_3345,N_502,N_1905);
or U3346 (N_3346,N_662,N_24);
nor U3347 (N_3347,N_1621,N_28);
xnor U3348 (N_3348,N_1334,N_2446);
and U3349 (N_3349,N_967,N_2126);
and U3350 (N_3350,N_424,N_1216);
nand U3351 (N_3351,N_1048,N_1553);
nor U3352 (N_3352,N_558,N_1754);
nor U3353 (N_3353,N_373,N_1959);
and U3354 (N_3354,N_2284,N_629);
or U3355 (N_3355,N_826,N_1499);
or U3356 (N_3356,N_419,N_1433);
nand U3357 (N_3357,N_298,N_1910);
and U3358 (N_3358,N_470,N_2315);
nor U3359 (N_3359,N_1822,N_602);
nand U3360 (N_3360,N_658,N_2225);
or U3361 (N_3361,N_1668,N_1975);
or U3362 (N_3362,N_1584,N_1451);
nor U3363 (N_3363,N_467,N_2481);
or U3364 (N_3364,N_2335,N_1363);
and U3365 (N_3365,N_1128,N_221);
nand U3366 (N_3366,N_871,N_1830);
and U3367 (N_3367,N_1752,N_911);
and U3368 (N_3368,N_98,N_2432);
nand U3369 (N_3369,N_2173,N_1285);
nand U3370 (N_3370,N_1523,N_1748);
xnor U3371 (N_3371,N_941,N_1405);
nand U3372 (N_3372,N_903,N_1582);
and U3373 (N_3373,N_1688,N_2179);
and U3374 (N_3374,N_1083,N_1345);
and U3375 (N_3375,N_943,N_2198);
or U3376 (N_3376,N_135,N_628);
and U3377 (N_3377,N_197,N_1615);
nor U3378 (N_3378,N_1105,N_1064);
nand U3379 (N_3379,N_1191,N_2035);
or U3380 (N_3380,N_185,N_453);
or U3381 (N_3381,N_1144,N_1648);
nand U3382 (N_3382,N_2070,N_122);
or U3383 (N_3383,N_463,N_1863);
and U3384 (N_3384,N_2371,N_2302);
or U3385 (N_3385,N_2439,N_995);
or U3386 (N_3386,N_1854,N_1012);
and U3387 (N_3387,N_2485,N_1575);
nand U3388 (N_3388,N_33,N_384);
nor U3389 (N_3389,N_1599,N_733);
nor U3390 (N_3390,N_1424,N_1781);
nor U3391 (N_3391,N_1416,N_2442);
nor U3392 (N_3392,N_2359,N_2031);
nor U3393 (N_3393,N_2267,N_2094);
or U3394 (N_3394,N_555,N_2419);
and U3395 (N_3395,N_2165,N_1194);
and U3396 (N_3396,N_2275,N_1887);
or U3397 (N_3397,N_2077,N_2475);
and U3398 (N_3398,N_1878,N_612);
or U3399 (N_3399,N_1265,N_1059);
and U3400 (N_3400,N_202,N_231);
or U3401 (N_3401,N_912,N_1558);
nand U3402 (N_3402,N_307,N_976);
nor U3403 (N_3403,N_973,N_1578);
nand U3404 (N_3404,N_2377,N_136);
nand U3405 (N_3405,N_588,N_364);
nand U3406 (N_3406,N_1778,N_792);
nand U3407 (N_3407,N_703,N_328);
xor U3408 (N_3408,N_2061,N_212);
nand U3409 (N_3409,N_2312,N_1022);
nand U3410 (N_3410,N_1641,N_2093);
and U3411 (N_3411,N_815,N_4);
nor U3412 (N_3412,N_2369,N_520);
nor U3413 (N_3413,N_1978,N_913);
nand U3414 (N_3414,N_1131,N_1227);
nand U3415 (N_3415,N_1467,N_958);
nor U3416 (N_3416,N_916,N_766);
and U3417 (N_3417,N_793,N_550);
nor U3418 (N_3418,N_1634,N_67);
or U3419 (N_3419,N_2388,N_880);
and U3420 (N_3420,N_2015,N_1298);
and U3421 (N_3421,N_130,N_2423);
xor U3422 (N_3422,N_2274,N_1124);
nand U3423 (N_3423,N_365,N_752);
and U3424 (N_3424,N_2133,N_2041);
and U3425 (N_3425,N_319,N_1098);
or U3426 (N_3426,N_337,N_1834);
nand U3427 (N_3427,N_1926,N_1710);
nor U3428 (N_3428,N_1080,N_1782);
nand U3429 (N_3429,N_1025,N_1988);
or U3430 (N_3430,N_408,N_905);
and U3431 (N_3431,N_436,N_1013);
or U3432 (N_3432,N_340,N_448);
nand U3433 (N_3433,N_758,N_1408);
nor U3434 (N_3434,N_1777,N_155);
or U3435 (N_3435,N_1179,N_1101);
and U3436 (N_3436,N_1689,N_1160);
nand U3437 (N_3437,N_1819,N_218);
nand U3438 (N_3438,N_1985,N_693);
nor U3439 (N_3439,N_1464,N_1437);
and U3440 (N_3440,N_1465,N_1492);
nor U3441 (N_3441,N_1095,N_465);
nand U3442 (N_3442,N_1909,N_1793);
or U3443 (N_3443,N_327,N_510);
nand U3444 (N_3444,N_370,N_1877);
nor U3445 (N_3445,N_914,N_1019);
nor U3446 (N_3446,N_1232,N_296);
nand U3447 (N_3447,N_1856,N_276);
nand U3448 (N_3448,N_53,N_1650);
or U3449 (N_3449,N_336,N_1477);
and U3450 (N_3450,N_694,N_1735);
or U3451 (N_3451,N_1811,N_268);
nand U3452 (N_3452,N_1580,N_1378);
and U3453 (N_3453,N_322,N_987);
nor U3454 (N_3454,N_2043,N_60);
or U3455 (N_3455,N_2443,N_406);
xnor U3456 (N_3456,N_945,N_94);
and U3457 (N_3457,N_147,N_413);
nand U3458 (N_3458,N_2333,N_323);
nor U3459 (N_3459,N_1994,N_1439);
nand U3460 (N_3460,N_2259,N_2466);
or U3461 (N_3461,N_1904,N_1186);
or U3462 (N_3462,N_1548,N_338);
nor U3463 (N_3463,N_1915,N_2368);
nand U3464 (N_3464,N_494,N_1127);
nor U3465 (N_3465,N_2277,N_1448);
nand U3466 (N_3466,N_1555,N_2488);
and U3467 (N_3467,N_2473,N_1261);
nor U3468 (N_3468,N_27,N_1020);
nand U3469 (N_3469,N_1666,N_2306);
nor U3470 (N_3470,N_133,N_928);
or U3471 (N_3471,N_2470,N_172);
nor U3472 (N_3472,N_753,N_1479);
nor U3473 (N_3473,N_939,N_1178);
nand U3474 (N_3474,N_426,N_1255);
and U3475 (N_3475,N_521,N_246);
and U3476 (N_3476,N_2205,N_1684);
nor U3477 (N_3477,N_1800,N_1755);
nor U3478 (N_3478,N_425,N_539);
nand U3479 (N_3479,N_1550,N_921);
and U3480 (N_3480,N_580,N_1808);
and U3481 (N_3481,N_1624,N_2054);
or U3482 (N_3482,N_1054,N_1899);
nor U3483 (N_3483,N_1699,N_1089);
nand U3484 (N_3484,N_1902,N_2343);
and U3485 (N_3485,N_2477,N_1780);
or U3486 (N_3486,N_935,N_1211);
nor U3487 (N_3487,N_1900,N_886);
nand U3488 (N_3488,N_283,N_2320);
nand U3489 (N_3489,N_1266,N_1149);
nor U3490 (N_3490,N_1122,N_1419);
nand U3491 (N_3491,N_1308,N_2262);
nand U3492 (N_3492,N_2240,N_183);
or U3493 (N_3493,N_2184,N_1219);
or U3494 (N_3494,N_632,N_1784);
and U3495 (N_3495,N_1005,N_1510);
and U3496 (N_3496,N_727,N_1644);
or U3497 (N_3497,N_1009,N_289);
xor U3498 (N_3498,N_782,N_1060);
nand U3499 (N_3499,N_1604,N_1589);
nor U3500 (N_3500,N_748,N_695);
nor U3501 (N_3501,N_910,N_402);
nor U3502 (N_3502,N_838,N_1446);
or U3503 (N_3503,N_1,N_2036);
nand U3504 (N_3504,N_1680,N_2412);
nor U3505 (N_3505,N_981,N_1138);
or U3506 (N_3506,N_110,N_690);
or U3507 (N_3507,N_1108,N_1274);
and U3508 (N_3508,N_1395,N_1292);
nor U3509 (N_3509,N_1304,N_537);
or U3510 (N_3510,N_530,N_111);
and U3511 (N_3511,N_2455,N_2281);
and U3512 (N_3512,N_1631,N_1923);
nor U3513 (N_3513,N_968,N_1342);
nand U3514 (N_3514,N_1166,N_11);
nor U3515 (N_3515,N_2107,N_1113);
or U3516 (N_3516,N_2420,N_546);
nand U3517 (N_3517,N_140,N_2067);
or U3518 (N_3518,N_947,N_1119);
or U3519 (N_3519,N_1922,N_20);
nand U3520 (N_3520,N_1677,N_1481);
nand U3521 (N_3521,N_1786,N_673);
and U3522 (N_3522,N_2143,N_1152);
nor U3523 (N_3523,N_1039,N_91);
nand U3524 (N_3524,N_2220,N_314);
nor U3525 (N_3525,N_501,N_845);
or U3526 (N_3526,N_686,N_1068);
nor U3527 (N_3527,N_616,N_820);
nand U3528 (N_3528,N_827,N_881);
or U3529 (N_3529,N_2292,N_2253);
nor U3530 (N_3530,N_1093,N_2347);
nand U3531 (N_3531,N_1109,N_2087);
and U3532 (N_3532,N_1407,N_251);
or U3533 (N_3533,N_1616,N_2321);
nor U3534 (N_3534,N_605,N_1050);
and U3535 (N_3535,N_2022,N_1511);
nor U3536 (N_3536,N_610,N_1821);
nor U3537 (N_3537,N_1690,N_526);
nand U3538 (N_3538,N_2116,N_264);
or U3539 (N_3539,N_1222,N_1933);
and U3540 (N_3540,N_1442,N_2392);
and U3541 (N_3541,N_1264,N_1806);
and U3542 (N_3542,N_1713,N_1788);
or U3543 (N_3543,N_615,N_1299);
and U3544 (N_3544,N_858,N_1044);
or U3545 (N_3545,N_934,N_1235);
and U3546 (N_3546,N_109,N_1173);
and U3547 (N_3547,N_1673,N_1538);
nor U3548 (N_3548,N_430,N_2104);
nand U3549 (N_3549,N_302,N_2494);
and U3550 (N_3550,N_1597,N_1458);
nand U3551 (N_3551,N_1943,N_46);
or U3552 (N_3552,N_2313,N_1711);
or U3553 (N_3553,N_1570,N_1636);
and U3554 (N_3554,N_2191,N_95);
nor U3555 (N_3555,N_255,N_1296);
and U3556 (N_3556,N_2197,N_1075);
nand U3557 (N_3557,N_908,N_500);
or U3558 (N_3558,N_1332,N_1659);
nor U3559 (N_3559,N_152,N_738);
xnor U3560 (N_3560,N_1303,N_581);
or U3561 (N_3561,N_2296,N_1251);
nand U3562 (N_3562,N_2150,N_1145);
and U3563 (N_3563,N_922,N_476);
nand U3564 (N_3564,N_1170,N_760);
nor U3565 (N_3565,N_1669,N_784);
or U3566 (N_3566,N_332,N_1002);
and U3567 (N_3567,N_377,N_1027);
and U3568 (N_3568,N_39,N_438);
and U3569 (N_3569,N_2157,N_2140);
or U3570 (N_3570,N_1056,N_668);
or U3571 (N_3571,N_1305,N_1588);
nor U3572 (N_3572,N_1140,N_2142);
nor U3573 (N_3573,N_1112,N_2076);
and U3574 (N_3574,N_1291,N_665);
nand U3575 (N_3575,N_2148,N_569);
nor U3576 (N_3576,N_2164,N_1195);
nand U3577 (N_3577,N_1522,N_2136);
nand U3578 (N_3578,N_1917,N_2028);
nand U3579 (N_3579,N_630,N_151);
nor U3580 (N_3580,N_639,N_940);
or U3581 (N_3581,N_932,N_1772);
or U3582 (N_3582,N_824,N_1794);
or U3583 (N_3583,N_1215,N_875);
and U3584 (N_3584,N_2218,N_1517);
nand U3585 (N_3585,N_293,N_855);
nor U3586 (N_3586,N_2092,N_1731);
nand U3587 (N_3587,N_1890,N_2385);
nand U3588 (N_3588,N_671,N_2353);
nand U3589 (N_3589,N_716,N_128);
or U3590 (N_3590,N_1494,N_1157);
nor U3591 (N_3591,N_1290,N_1137);
nand U3592 (N_3592,N_1454,N_1592);
or U3593 (N_3593,N_722,N_2434);
or U3594 (N_3594,N_1200,N_770);
or U3595 (N_3595,N_975,N_1564);
nor U3596 (N_3596,N_1242,N_1957);
or U3597 (N_3597,N_568,N_1591);
nand U3598 (N_3598,N_1514,N_692);
and U3599 (N_3599,N_780,N_1188);
nand U3600 (N_3600,N_1833,N_2483);
and U3601 (N_3601,N_1028,N_2406);
and U3602 (N_3602,N_2383,N_1733);
and U3603 (N_3603,N_1367,N_661);
or U3604 (N_3604,N_2160,N_2345);
nand U3605 (N_3605,N_1561,N_1554);
nor U3606 (N_3606,N_18,N_1695);
nor U3607 (N_3607,N_2005,N_1719);
and U3608 (N_3608,N_75,N_1371);
nor U3609 (N_3609,N_1486,N_1365);
and U3610 (N_3610,N_15,N_82);
nor U3611 (N_3611,N_697,N_954);
nand U3612 (N_3612,N_2073,N_2465);
nor U3613 (N_3613,N_1876,N_366);
and U3614 (N_3614,N_1301,N_2309);
or U3615 (N_3615,N_1627,N_1925);
or U3616 (N_3616,N_955,N_2461);
and U3617 (N_3617,N_1256,N_1444);
and U3618 (N_3618,N_2241,N_2261);
and U3619 (N_3619,N_66,N_433);
nand U3620 (N_3620,N_2433,N_85);
and U3621 (N_3621,N_2204,N_1610);
or U3622 (N_3622,N_1880,N_706);
and U3623 (N_3623,N_1070,N_1563);
nor U3624 (N_3624,N_808,N_1939);
or U3625 (N_3625,N_1384,N_177);
nor U3626 (N_3626,N_249,N_2304);
or U3627 (N_3627,N_2011,N_1443);
nor U3628 (N_3628,N_1590,N_299);
nand U3629 (N_3629,N_490,N_1891);
nor U3630 (N_3630,N_318,N_2257);
nand U3631 (N_3631,N_535,N_452);
nand U3632 (N_3632,N_62,N_1277);
nor U3633 (N_3633,N_834,N_1055);
and U3634 (N_3634,N_1997,N_1445);
or U3635 (N_3635,N_715,N_1233);
nor U3636 (N_3636,N_1040,N_2391);
or U3637 (N_3637,N_161,N_1530);
and U3638 (N_3638,N_1649,N_2297);
nand U3639 (N_3639,N_839,N_2413);
and U3640 (N_3640,N_12,N_1642);
nor U3641 (N_3641,N_772,N_330);
nor U3642 (N_3642,N_1350,N_349);
nor U3643 (N_3643,N_523,N_428);
or U3644 (N_3644,N_1762,N_666);
or U3645 (N_3645,N_1294,N_1143);
and U3646 (N_3646,N_2314,N_509);
and U3647 (N_3647,N_48,N_1252);
nor U3648 (N_3648,N_1598,N_1745);
or U3649 (N_3649,N_2493,N_137);
nand U3650 (N_3650,N_1206,N_2491);
and U3651 (N_3651,N_794,N_756);
nand U3652 (N_3652,N_624,N_357);
and U3653 (N_3653,N_2228,N_236);
and U3654 (N_3654,N_1006,N_627);
or U3655 (N_3655,N_1346,N_474);
nand U3656 (N_3656,N_2492,N_1656);
nand U3657 (N_3657,N_1065,N_1007);
and U3658 (N_3658,N_745,N_1014);
and U3659 (N_3659,N_2330,N_1229);
and U3660 (N_3660,N_339,N_2400);
nor U3661 (N_3661,N_1512,N_156);
xor U3662 (N_3662,N_1221,N_2159);
and U3663 (N_3663,N_495,N_1770);
nand U3664 (N_3664,N_2183,N_835);
or U3665 (N_3665,N_899,N_909);
and U3666 (N_3666,N_821,N_1422);
or U3667 (N_3667,N_2416,N_409);
or U3668 (N_3668,N_76,N_1319);
nor U3669 (N_3669,N_1073,N_1738);
nor U3670 (N_3670,N_1942,N_1069);
and U3671 (N_3671,N_1543,N_1250);
or U3672 (N_3672,N_1835,N_2290);
nor U3673 (N_3673,N_2431,N_1741);
nand U3674 (N_3674,N_816,N_1402);
and U3675 (N_3675,N_1965,N_8);
nor U3676 (N_3676,N_1414,N_1369);
or U3677 (N_3677,N_2039,N_1539);
nor U3678 (N_3678,N_556,N_2379);
nand U3679 (N_3679,N_2010,N_1158);
nor U3680 (N_3680,N_208,N_2209);
and U3681 (N_3681,N_375,N_2397);
nand U3682 (N_3682,N_1172,N_1390);
and U3683 (N_3683,N_737,N_1021);
nor U3684 (N_3684,N_2188,N_1737);
or U3685 (N_3685,N_664,N_1047);
and U3686 (N_3686,N_1354,N_2464);
nand U3687 (N_3687,N_352,N_1432);
or U3688 (N_3688,N_2248,N_1495);
and U3689 (N_3689,N_2,N_2249);
and U3690 (N_3690,N_525,N_1783);
nand U3691 (N_3691,N_1843,N_1484);
nor U3692 (N_3692,N_224,N_1366);
and U3693 (N_3693,N_1017,N_439);
or U3694 (N_3694,N_80,N_1645);
xor U3695 (N_3695,N_506,N_1485);
or U3696 (N_3696,N_31,N_529);
nand U3697 (N_3697,N_144,N_759);
nand U3698 (N_3698,N_646,N_1150);
and U3699 (N_3699,N_1198,N_489);
and U3700 (N_3700,N_184,N_2301);
or U3701 (N_3701,N_862,N_105);
nand U3702 (N_3702,N_2300,N_1577);
nor U3703 (N_3703,N_1799,N_709);
xor U3704 (N_3704,N_2325,N_971);
nor U3705 (N_3705,N_2129,N_524);
nor U3706 (N_3706,N_132,N_1078);
and U3707 (N_3707,N_2127,N_776);
nand U3708 (N_3708,N_1326,N_552);
or U3709 (N_3709,N_2055,N_308);
nand U3710 (N_3710,N_1045,N_1931);
and U3711 (N_3711,N_1855,N_806);
or U3712 (N_3712,N_2131,N_1295);
and U3713 (N_3713,N_1620,N_1525);
nor U3714 (N_3714,N_372,N_262);
or U3715 (N_3715,N_131,N_325);
and U3716 (N_3716,N_1042,N_214);
nor U3717 (N_3717,N_396,N_189);
or U3718 (N_3718,N_2199,N_1753);
or U3719 (N_3719,N_19,N_1560);
or U3720 (N_3720,N_1790,N_1546);
and U3721 (N_3721,N_2101,N_1361);
and U3722 (N_3722,N_942,N_77);
nand U3723 (N_3723,N_2403,N_2344);
nor U3724 (N_3724,N_2350,N_1004);
and U3725 (N_3725,N_1241,N_2017);
nand U3726 (N_3726,N_2265,N_1967);
nor U3727 (N_3727,N_2098,N_1804);
nor U3728 (N_3728,N_620,N_2103);
nor U3729 (N_3729,N_267,N_215);
nand U3730 (N_3730,N_833,N_1896);
nand U3731 (N_3731,N_2100,N_1765);
and U3732 (N_3732,N_1533,N_859);
and U3733 (N_3733,N_456,N_2090);
or U3734 (N_3734,N_479,N_1057);
and U3735 (N_3735,N_1470,N_1209);
and U3736 (N_3736,N_1920,N_562);
nor U3737 (N_3737,N_1726,N_992);
nand U3738 (N_3738,N_362,N_1715);
nand U3739 (N_3739,N_292,N_2163);
or U3740 (N_3740,N_1937,N_499);
or U3741 (N_3741,N_1983,N_596);
nand U3742 (N_3742,N_1761,N_468);
nor U3743 (N_3743,N_2186,N_458);
nand U3744 (N_3744,N_1594,N_84);
and U3745 (N_3745,N_1894,N_1798);
and U3746 (N_3746,N_767,N_785);
nor U3747 (N_3747,N_1373,N_1267);
and U3748 (N_3748,N_2109,N_2390);
nand U3749 (N_3749,N_2346,N_290);
or U3750 (N_3750,N_1341,N_1414);
or U3751 (N_3751,N_2244,N_1314);
and U3752 (N_3752,N_1795,N_581);
xnor U3753 (N_3753,N_1677,N_2493);
nand U3754 (N_3754,N_1103,N_467);
nor U3755 (N_3755,N_1444,N_235);
and U3756 (N_3756,N_1930,N_1346);
and U3757 (N_3757,N_84,N_658);
nor U3758 (N_3758,N_156,N_399);
or U3759 (N_3759,N_1260,N_480);
or U3760 (N_3760,N_2243,N_974);
or U3761 (N_3761,N_2164,N_1057);
or U3762 (N_3762,N_1835,N_629);
or U3763 (N_3763,N_1147,N_1530);
or U3764 (N_3764,N_2105,N_1310);
nand U3765 (N_3765,N_750,N_221);
nor U3766 (N_3766,N_4,N_718);
nor U3767 (N_3767,N_2280,N_2361);
or U3768 (N_3768,N_939,N_2130);
and U3769 (N_3769,N_1103,N_748);
nand U3770 (N_3770,N_561,N_1070);
nor U3771 (N_3771,N_394,N_1394);
nand U3772 (N_3772,N_2340,N_1838);
nand U3773 (N_3773,N_1281,N_364);
nand U3774 (N_3774,N_1657,N_759);
and U3775 (N_3775,N_983,N_1496);
nor U3776 (N_3776,N_1509,N_638);
nor U3777 (N_3777,N_2378,N_104);
and U3778 (N_3778,N_2117,N_439);
or U3779 (N_3779,N_193,N_839);
and U3780 (N_3780,N_1753,N_441);
nand U3781 (N_3781,N_2107,N_1485);
and U3782 (N_3782,N_1184,N_1984);
nor U3783 (N_3783,N_1025,N_2082);
nor U3784 (N_3784,N_2493,N_1944);
or U3785 (N_3785,N_414,N_242);
nand U3786 (N_3786,N_1005,N_2103);
or U3787 (N_3787,N_1797,N_2436);
and U3788 (N_3788,N_1411,N_835);
nor U3789 (N_3789,N_15,N_2431);
nand U3790 (N_3790,N_474,N_1124);
xnor U3791 (N_3791,N_1761,N_383);
nand U3792 (N_3792,N_427,N_1002);
xor U3793 (N_3793,N_902,N_1804);
nor U3794 (N_3794,N_1016,N_1303);
nor U3795 (N_3795,N_674,N_1322);
nor U3796 (N_3796,N_1481,N_679);
nand U3797 (N_3797,N_1303,N_1149);
xor U3798 (N_3798,N_963,N_127);
or U3799 (N_3799,N_1430,N_1225);
nand U3800 (N_3800,N_1548,N_1426);
or U3801 (N_3801,N_2143,N_496);
or U3802 (N_3802,N_890,N_1023);
nor U3803 (N_3803,N_1629,N_2318);
and U3804 (N_3804,N_1908,N_814);
nor U3805 (N_3805,N_1034,N_1252);
and U3806 (N_3806,N_325,N_1658);
xor U3807 (N_3807,N_336,N_2246);
nand U3808 (N_3808,N_473,N_2400);
nor U3809 (N_3809,N_2284,N_708);
nor U3810 (N_3810,N_798,N_2137);
and U3811 (N_3811,N_125,N_2051);
or U3812 (N_3812,N_1281,N_537);
nor U3813 (N_3813,N_1336,N_756);
and U3814 (N_3814,N_712,N_1153);
or U3815 (N_3815,N_1981,N_1644);
nor U3816 (N_3816,N_1877,N_633);
nor U3817 (N_3817,N_2478,N_1749);
or U3818 (N_3818,N_52,N_1929);
nor U3819 (N_3819,N_222,N_1284);
and U3820 (N_3820,N_248,N_1990);
nor U3821 (N_3821,N_734,N_541);
nor U3822 (N_3822,N_996,N_832);
nand U3823 (N_3823,N_907,N_891);
nand U3824 (N_3824,N_1506,N_1028);
nor U3825 (N_3825,N_1587,N_706);
and U3826 (N_3826,N_1016,N_1352);
nor U3827 (N_3827,N_1239,N_1608);
or U3828 (N_3828,N_1025,N_847);
nor U3829 (N_3829,N_468,N_1973);
nor U3830 (N_3830,N_365,N_1138);
nand U3831 (N_3831,N_1021,N_848);
and U3832 (N_3832,N_1021,N_2023);
nand U3833 (N_3833,N_198,N_418);
and U3834 (N_3834,N_1634,N_1740);
nand U3835 (N_3835,N_1747,N_1243);
or U3836 (N_3836,N_1229,N_1428);
or U3837 (N_3837,N_627,N_1672);
nor U3838 (N_3838,N_2261,N_1180);
and U3839 (N_3839,N_103,N_2020);
nor U3840 (N_3840,N_1505,N_1971);
nand U3841 (N_3841,N_193,N_1879);
nor U3842 (N_3842,N_974,N_143);
and U3843 (N_3843,N_1302,N_1531);
and U3844 (N_3844,N_1105,N_1292);
or U3845 (N_3845,N_74,N_2486);
and U3846 (N_3846,N_1561,N_2403);
or U3847 (N_3847,N_597,N_1072);
nand U3848 (N_3848,N_1523,N_225);
and U3849 (N_3849,N_582,N_1852);
and U3850 (N_3850,N_1501,N_259);
or U3851 (N_3851,N_112,N_891);
nor U3852 (N_3852,N_641,N_1120);
and U3853 (N_3853,N_1397,N_1134);
nor U3854 (N_3854,N_1882,N_940);
nand U3855 (N_3855,N_534,N_394);
nand U3856 (N_3856,N_544,N_1727);
and U3857 (N_3857,N_1029,N_2226);
nand U3858 (N_3858,N_436,N_72);
nand U3859 (N_3859,N_2400,N_2256);
or U3860 (N_3860,N_1867,N_123);
nor U3861 (N_3861,N_884,N_1017);
and U3862 (N_3862,N_558,N_84);
nor U3863 (N_3863,N_32,N_882);
nor U3864 (N_3864,N_2323,N_1774);
nand U3865 (N_3865,N_2498,N_756);
or U3866 (N_3866,N_2189,N_1862);
and U3867 (N_3867,N_1546,N_939);
or U3868 (N_3868,N_587,N_2260);
nor U3869 (N_3869,N_800,N_854);
or U3870 (N_3870,N_1916,N_140);
and U3871 (N_3871,N_1193,N_224);
or U3872 (N_3872,N_261,N_650);
and U3873 (N_3873,N_941,N_1685);
xor U3874 (N_3874,N_1856,N_964);
nor U3875 (N_3875,N_982,N_2423);
nand U3876 (N_3876,N_639,N_793);
and U3877 (N_3877,N_2458,N_1203);
and U3878 (N_3878,N_825,N_888);
and U3879 (N_3879,N_29,N_1927);
and U3880 (N_3880,N_1511,N_1683);
nor U3881 (N_3881,N_19,N_473);
and U3882 (N_3882,N_1329,N_523);
and U3883 (N_3883,N_1759,N_1371);
and U3884 (N_3884,N_429,N_256);
nor U3885 (N_3885,N_982,N_481);
or U3886 (N_3886,N_1149,N_71);
or U3887 (N_3887,N_22,N_1889);
or U3888 (N_3888,N_678,N_815);
nand U3889 (N_3889,N_1407,N_2291);
or U3890 (N_3890,N_1442,N_931);
nor U3891 (N_3891,N_2135,N_1994);
nand U3892 (N_3892,N_230,N_242);
and U3893 (N_3893,N_1206,N_191);
nand U3894 (N_3894,N_1725,N_681);
and U3895 (N_3895,N_2029,N_1322);
nand U3896 (N_3896,N_773,N_2002);
nand U3897 (N_3897,N_2365,N_1659);
or U3898 (N_3898,N_2395,N_1662);
nand U3899 (N_3899,N_1717,N_1639);
or U3900 (N_3900,N_2260,N_1882);
nor U3901 (N_3901,N_717,N_1592);
nand U3902 (N_3902,N_417,N_2070);
nor U3903 (N_3903,N_1948,N_1609);
or U3904 (N_3904,N_388,N_2170);
and U3905 (N_3905,N_1595,N_1695);
and U3906 (N_3906,N_1022,N_2350);
and U3907 (N_3907,N_2264,N_1865);
nand U3908 (N_3908,N_334,N_2308);
or U3909 (N_3909,N_946,N_2478);
nand U3910 (N_3910,N_768,N_582);
xor U3911 (N_3911,N_2077,N_1885);
nand U3912 (N_3912,N_232,N_1670);
nor U3913 (N_3913,N_420,N_270);
and U3914 (N_3914,N_1569,N_1276);
or U3915 (N_3915,N_1686,N_548);
or U3916 (N_3916,N_1553,N_1177);
nand U3917 (N_3917,N_1806,N_309);
nor U3918 (N_3918,N_2297,N_1281);
and U3919 (N_3919,N_310,N_81);
or U3920 (N_3920,N_2330,N_2367);
or U3921 (N_3921,N_1488,N_2345);
and U3922 (N_3922,N_1866,N_840);
nand U3923 (N_3923,N_1962,N_1447);
nand U3924 (N_3924,N_2488,N_790);
and U3925 (N_3925,N_978,N_895);
nand U3926 (N_3926,N_2159,N_1847);
nor U3927 (N_3927,N_1081,N_996);
nand U3928 (N_3928,N_133,N_468);
nand U3929 (N_3929,N_801,N_139);
nand U3930 (N_3930,N_2461,N_2356);
and U3931 (N_3931,N_237,N_1285);
or U3932 (N_3932,N_1464,N_1958);
or U3933 (N_3933,N_1651,N_1689);
nand U3934 (N_3934,N_866,N_1646);
and U3935 (N_3935,N_1189,N_2467);
nor U3936 (N_3936,N_2429,N_944);
nor U3937 (N_3937,N_163,N_873);
nor U3938 (N_3938,N_1454,N_388);
and U3939 (N_3939,N_1692,N_2387);
or U3940 (N_3940,N_1715,N_587);
nor U3941 (N_3941,N_470,N_2063);
and U3942 (N_3942,N_1585,N_1533);
or U3943 (N_3943,N_1219,N_470);
xnor U3944 (N_3944,N_1398,N_454);
nand U3945 (N_3945,N_315,N_1927);
nor U3946 (N_3946,N_1292,N_1494);
or U3947 (N_3947,N_731,N_1699);
nor U3948 (N_3948,N_1637,N_1202);
nand U3949 (N_3949,N_1500,N_1427);
nor U3950 (N_3950,N_2227,N_1729);
or U3951 (N_3951,N_1946,N_695);
nand U3952 (N_3952,N_1385,N_1135);
and U3953 (N_3953,N_1904,N_2181);
and U3954 (N_3954,N_129,N_2113);
and U3955 (N_3955,N_74,N_424);
nand U3956 (N_3956,N_1960,N_2);
or U3957 (N_3957,N_1401,N_1841);
nor U3958 (N_3958,N_246,N_101);
nand U3959 (N_3959,N_1228,N_819);
nor U3960 (N_3960,N_453,N_1527);
and U3961 (N_3961,N_1460,N_787);
and U3962 (N_3962,N_480,N_1279);
or U3963 (N_3963,N_495,N_2127);
or U3964 (N_3964,N_1801,N_1007);
or U3965 (N_3965,N_421,N_2426);
nand U3966 (N_3966,N_2139,N_1581);
and U3967 (N_3967,N_946,N_1857);
or U3968 (N_3968,N_1252,N_465);
or U3969 (N_3969,N_1226,N_2157);
nand U3970 (N_3970,N_319,N_2473);
nor U3971 (N_3971,N_837,N_1950);
nor U3972 (N_3972,N_2039,N_1887);
or U3973 (N_3973,N_2251,N_1510);
nor U3974 (N_3974,N_2028,N_935);
nand U3975 (N_3975,N_933,N_1467);
nor U3976 (N_3976,N_487,N_996);
or U3977 (N_3977,N_2168,N_1143);
nor U3978 (N_3978,N_1702,N_1678);
nor U3979 (N_3979,N_925,N_1722);
and U3980 (N_3980,N_1236,N_828);
or U3981 (N_3981,N_348,N_855);
and U3982 (N_3982,N_2081,N_1752);
and U3983 (N_3983,N_158,N_1982);
or U3984 (N_3984,N_925,N_2380);
or U3985 (N_3985,N_712,N_561);
nor U3986 (N_3986,N_1261,N_1236);
or U3987 (N_3987,N_320,N_419);
nor U3988 (N_3988,N_1207,N_2280);
and U3989 (N_3989,N_584,N_1086);
nand U3990 (N_3990,N_902,N_992);
nor U3991 (N_3991,N_414,N_947);
or U3992 (N_3992,N_664,N_25);
or U3993 (N_3993,N_836,N_666);
nor U3994 (N_3994,N_378,N_2352);
or U3995 (N_3995,N_84,N_1674);
and U3996 (N_3996,N_11,N_1427);
nor U3997 (N_3997,N_241,N_2431);
nor U3998 (N_3998,N_1354,N_1780);
or U3999 (N_3999,N_2,N_847);
and U4000 (N_4000,N_286,N_672);
and U4001 (N_4001,N_2213,N_910);
or U4002 (N_4002,N_1105,N_1010);
and U4003 (N_4003,N_1361,N_2162);
nand U4004 (N_4004,N_1807,N_1722);
and U4005 (N_4005,N_886,N_1127);
and U4006 (N_4006,N_1254,N_979);
and U4007 (N_4007,N_459,N_973);
or U4008 (N_4008,N_1294,N_2061);
nor U4009 (N_4009,N_988,N_1452);
or U4010 (N_4010,N_25,N_1218);
and U4011 (N_4011,N_2144,N_995);
and U4012 (N_4012,N_1202,N_7);
and U4013 (N_4013,N_1653,N_1829);
nand U4014 (N_4014,N_2465,N_1077);
or U4015 (N_4015,N_2151,N_1193);
nor U4016 (N_4016,N_478,N_761);
nor U4017 (N_4017,N_1467,N_1941);
and U4018 (N_4018,N_580,N_418);
xnor U4019 (N_4019,N_1078,N_925);
nor U4020 (N_4020,N_1873,N_1733);
nor U4021 (N_4021,N_6,N_373);
or U4022 (N_4022,N_1305,N_843);
nand U4023 (N_4023,N_1287,N_1810);
nor U4024 (N_4024,N_1812,N_89);
nand U4025 (N_4025,N_740,N_1429);
nor U4026 (N_4026,N_1300,N_541);
nand U4027 (N_4027,N_1409,N_1812);
and U4028 (N_4028,N_1548,N_671);
nand U4029 (N_4029,N_59,N_638);
or U4030 (N_4030,N_2060,N_548);
nor U4031 (N_4031,N_308,N_140);
nand U4032 (N_4032,N_913,N_517);
or U4033 (N_4033,N_1708,N_1579);
xnor U4034 (N_4034,N_1112,N_2256);
and U4035 (N_4035,N_1948,N_1892);
xnor U4036 (N_4036,N_105,N_1452);
or U4037 (N_4037,N_1938,N_2444);
and U4038 (N_4038,N_1316,N_2252);
nand U4039 (N_4039,N_502,N_214);
or U4040 (N_4040,N_711,N_2325);
or U4041 (N_4041,N_1469,N_2221);
xor U4042 (N_4042,N_1918,N_778);
nand U4043 (N_4043,N_501,N_858);
and U4044 (N_4044,N_2438,N_2026);
nand U4045 (N_4045,N_239,N_1689);
and U4046 (N_4046,N_12,N_1171);
and U4047 (N_4047,N_1973,N_566);
and U4048 (N_4048,N_1052,N_321);
nor U4049 (N_4049,N_106,N_386);
and U4050 (N_4050,N_2164,N_2095);
or U4051 (N_4051,N_1601,N_2110);
nand U4052 (N_4052,N_1786,N_628);
nor U4053 (N_4053,N_2455,N_371);
and U4054 (N_4054,N_1521,N_2000);
nand U4055 (N_4055,N_1421,N_15);
and U4056 (N_4056,N_1912,N_1407);
nor U4057 (N_4057,N_652,N_61);
nor U4058 (N_4058,N_1139,N_185);
or U4059 (N_4059,N_572,N_1856);
nor U4060 (N_4060,N_2063,N_30);
and U4061 (N_4061,N_137,N_1998);
nand U4062 (N_4062,N_627,N_805);
and U4063 (N_4063,N_2288,N_260);
nand U4064 (N_4064,N_662,N_340);
nor U4065 (N_4065,N_2283,N_2388);
nand U4066 (N_4066,N_715,N_886);
and U4067 (N_4067,N_2473,N_632);
nand U4068 (N_4068,N_2396,N_2323);
or U4069 (N_4069,N_957,N_124);
nand U4070 (N_4070,N_663,N_1741);
nand U4071 (N_4071,N_1275,N_359);
and U4072 (N_4072,N_745,N_2496);
and U4073 (N_4073,N_1716,N_583);
xnor U4074 (N_4074,N_1684,N_575);
and U4075 (N_4075,N_258,N_1332);
and U4076 (N_4076,N_823,N_1664);
or U4077 (N_4077,N_74,N_489);
nand U4078 (N_4078,N_330,N_321);
or U4079 (N_4079,N_1607,N_1490);
or U4080 (N_4080,N_2227,N_881);
or U4081 (N_4081,N_246,N_609);
nor U4082 (N_4082,N_1047,N_590);
nor U4083 (N_4083,N_2247,N_1424);
and U4084 (N_4084,N_1841,N_180);
xor U4085 (N_4085,N_664,N_550);
xor U4086 (N_4086,N_581,N_271);
nand U4087 (N_4087,N_819,N_1468);
and U4088 (N_4088,N_1416,N_2204);
nand U4089 (N_4089,N_1633,N_437);
or U4090 (N_4090,N_1239,N_670);
nand U4091 (N_4091,N_2085,N_1807);
or U4092 (N_4092,N_911,N_741);
and U4093 (N_4093,N_2184,N_26);
nand U4094 (N_4094,N_1461,N_2221);
nand U4095 (N_4095,N_694,N_919);
nand U4096 (N_4096,N_750,N_1383);
or U4097 (N_4097,N_1270,N_733);
or U4098 (N_4098,N_1624,N_1983);
or U4099 (N_4099,N_2333,N_1144);
nor U4100 (N_4100,N_930,N_398);
and U4101 (N_4101,N_2486,N_1831);
and U4102 (N_4102,N_298,N_2485);
nor U4103 (N_4103,N_1555,N_442);
and U4104 (N_4104,N_116,N_642);
nor U4105 (N_4105,N_1698,N_692);
nand U4106 (N_4106,N_1817,N_2002);
nor U4107 (N_4107,N_1586,N_846);
and U4108 (N_4108,N_2123,N_257);
or U4109 (N_4109,N_2421,N_514);
or U4110 (N_4110,N_2252,N_1884);
nor U4111 (N_4111,N_591,N_2225);
xor U4112 (N_4112,N_2261,N_380);
xnor U4113 (N_4113,N_1454,N_1834);
nand U4114 (N_4114,N_74,N_2499);
nor U4115 (N_4115,N_1275,N_34);
or U4116 (N_4116,N_1302,N_322);
nor U4117 (N_4117,N_1753,N_1361);
nor U4118 (N_4118,N_831,N_860);
nor U4119 (N_4119,N_242,N_900);
and U4120 (N_4120,N_365,N_2154);
and U4121 (N_4121,N_952,N_1162);
nand U4122 (N_4122,N_560,N_951);
and U4123 (N_4123,N_1511,N_1660);
nor U4124 (N_4124,N_644,N_866);
nor U4125 (N_4125,N_1124,N_1701);
nor U4126 (N_4126,N_715,N_1324);
nor U4127 (N_4127,N_2396,N_2333);
nand U4128 (N_4128,N_787,N_1422);
nor U4129 (N_4129,N_1698,N_1344);
nand U4130 (N_4130,N_597,N_1886);
nor U4131 (N_4131,N_1182,N_2408);
and U4132 (N_4132,N_1193,N_612);
nand U4133 (N_4133,N_279,N_539);
nor U4134 (N_4134,N_734,N_1863);
and U4135 (N_4135,N_874,N_1759);
nor U4136 (N_4136,N_995,N_1025);
or U4137 (N_4137,N_616,N_1829);
nor U4138 (N_4138,N_317,N_291);
or U4139 (N_4139,N_749,N_1587);
nor U4140 (N_4140,N_38,N_1721);
and U4141 (N_4141,N_379,N_55);
or U4142 (N_4142,N_1669,N_1576);
nand U4143 (N_4143,N_1592,N_340);
nand U4144 (N_4144,N_1869,N_1752);
or U4145 (N_4145,N_1975,N_616);
and U4146 (N_4146,N_2045,N_1407);
or U4147 (N_4147,N_1434,N_1367);
nand U4148 (N_4148,N_96,N_988);
or U4149 (N_4149,N_920,N_2108);
and U4150 (N_4150,N_493,N_1215);
and U4151 (N_4151,N_1592,N_243);
nand U4152 (N_4152,N_2486,N_678);
and U4153 (N_4153,N_741,N_399);
and U4154 (N_4154,N_392,N_2403);
xnor U4155 (N_4155,N_1353,N_1541);
nand U4156 (N_4156,N_2168,N_1760);
nand U4157 (N_4157,N_1567,N_1776);
nor U4158 (N_4158,N_1559,N_346);
nand U4159 (N_4159,N_1937,N_632);
nor U4160 (N_4160,N_1716,N_2309);
xor U4161 (N_4161,N_1986,N_1316);
or U4162 (N_4162,N_191,N_1389);
or U4163 (N_4163,N_1183,N_1729);
nor U4164 (N_4164,N_586,N_1182);
and U4165 (N_4165,N_1558,N_1135);
and U4166 (N_4166,N_2016,N_850);
nor U4167 (N_4167,N_833,N_1222);
nor U4168 (N_4168,N_1514,N_131);
and U4169 (N_4169,N_5,N_1644);
nor U4170 (N_4170,N_2369,N_2479);
or U4171 (N_4171,N_1642,N_1266);
and U4172 (N_4172,N_350,N_136);
nand U4173 (N_4173,N_1054,N_1173);
nor U4174 (N_4174,N_2151,N_1448);
nor U4175 (N_4175,N_2262,N_820);
nand U4176 (N_4176,N_954,N_770);
nand U4177 (N_4177,N_396,N_547);
and U4178 (N_4178,N_1156,N_620);
or U4179 (N_4179,N_1527,N_1019);
nand U4180 (N_4180,N_56,N_117);
nand U4181 (N_4181,N_2183,N_1217);
or U4182 (N_4182,N_519,N_1879);
and U4183 (N_4183,N_184,N_448);
and U4184 (N_4184,N_75,N_899);
nand U4185 (N_4185,N_790,N_2477);
and U4186 (N_4186,N_2323,N_190);
nor U4187 (N_4187,N_1383,N_2017);
nand U4188 (N_4188,N_882,N_1544);
or U4189 (N_4189,N_1015,N_1529);
or U4190 (N_4190,N_1945,N_1819);
nand U4191 (N_4191,N_585,N_275);
nor U4192 (N_4192,N_634,N_1558);
nor U4193 (N_4193,N_1453,N_1867);
and U4194 (N_4194,N_1772,N_1570);
xor U4195 (N_4195,N_50,N_25);
nand U4196 (N_4196,N_1523,N_191);
and U4197 (N_4197,N_1951,N_1551);
nor U4198 (N_4198,N_1931,N_2439);
nand U4199 (N_4199,N_1980,N_144);
and U4200 (N_4200,N_523,N_849);
nand U4201 (N_4201,N_758,N_894);
or U4202 (N_4202,N_1980,N_19);
nand U4203 (N_4203,N_1201,N_1685);
nor U4204 (N_4204,N_110,N_1475);
nor U4205 (N_4205,N_925,N_778);
nand U4206 (N_4206,N_538,N_216);
and U4207 (N_4207,N_295,N_173);
or U4208 (N_4208,N_1234,N_2260);
or U4209 (N_4209,N_402,N_2400);
nor U4210 (N_4210,N_1051,N_1210);
nand U4211 (N_4211,N_1198,N_1907);
or U4212 (N_4212,N_1461,N_1235);
and U4213 (N_4213,N_1117,N_1101);
nor U4214 (N_4214,N_1988,N_2206);
or U4215 (N_4215,N_2385,N_1983);
and U4216 (N_4216,N_2359,N_1783);
nand U4217 (N_4217,N_2381,N_2442);
nor U4218 (N_4218,N_988,N_1250);
nor U4219 (N_4219,N_592,N_209);
nand U4220 (N_4220,N_2063,N_1967);
nor U4221 (N_4221,N_812,N_1431);
and U4222 (N_4222,N_1522,N_2028);
nand U4223 (N_4223,N_36,N_1254);
and U4224 (N_4224,N_914,N_1332);
and U4225 (N_4225,N_107,N_1048);
nor U4226 (N_4226,N_138,N_825);
nor U4227 (N_4227,N_489,N_1717);
nor U4228 (N_4228,N_1017,N_1043);
nor U4229 (N_4229,N_801,N_1985);
or U4230 (N_4230,N_415,N_1088);
nand U4231 (N_4231,N_2022,N_2402);
nand U4232 (N_4232,N_766,N_256);
and U4233 (N_4233,N_1670,N_2139);
nor U4234 (N_4234,N_2357,N_2051);
nand U4235 (N_4235,N_192,N_515);
nor U4236 (N_4236,N_614,N_2129);
nand U4237 (N_4237,N_288,N_1469);
and U4238 (N_4238,N_1574,N_1207);
nand U4239 (N_4239,N_2255,N_465);
nor U4240 (N_4240,N_900,N_1385);
nand U4241 (N_4241,N_1487,N_422);
nand U4242 (N_4242,N_2035,N_485);
and U4243 (N_4243,N_292,N_221);
nand U4244 (N_4244,N_1026,N_1118);
or U4245 (N_4245,N_1788,N_1549);
and U4246 (N_4246,N_907,N_827);
and U4247 (N_4247,N_1396,N_1627);
and U4248 (N_4248,N_1345,N_1786);
and U4249 (N_4249,N_1419,N_1310);
and U4250 (N_4250,N_1231,N_325);
and U4251 (N_4251,N_1193,N_319);
or U4252 (N_4252,N_1494,N_1927);
and U4253 (N_4253,N_2006,N_1499);
and U4254 (N_4254,N_677,N_2087);
and U4255 (N_4255,N_1505,N_872);
and U4256 (N_4256,N_2231,N_377);
nand U4257 (N_4257,N_148,N_716);
or U4258 (N_4258,N_1131,N_1021);
nor U4259 (N_4259,N_59,N_2140);
and U4260 (N_4260,N_100,N_1205);
or U4261 (N_4261,N_39,N_226);
or U4262 (N_4262,N_797,N_1751);
and U4263 (N_4263,N_1746,N_2307);
or U4264 (N_4264,N_934,N_1439);
nand U4265 (N_4265,N_2233,N_2103);
nand U4266 (N_4266,N_1962,N_183);
nand U4267 (N_4267,N_695,N_1428);
and U4268 (N_4268,N_1511,N_2249);
or U4269 (N_4269,N_12,N_1513);
and U4270 (N_4270,N_2430,N_62);
nor U4271 (N_4271,N_1096,N_1250);
nor U4272 (N_4272,N_2330,N_1774);
and U4273 (N_4273,N_1509,N_2303);
and U4274 (N_4274,N_1143,N_1168);
and U4275 (N_4275,N_1378,N_1757);
nand U4276 (N_4276,N_1313,N_1967);
and U4277 (N_4277,N_2375,N_1207);
nand U4278 (N_4278,N_2392,N_281);
and U4279 (N_4279,N_773,N_1010);
nand U4280 (N_4280,N_2375,N_743);
nor U4281 (N_4281,N_2148,N_731);
nor U4282 (N_4282,N_102,N_321);
and U4283 (N_4283,N_1457,N_2441);
nor U4284 (N_4284,N_393,N_50);
nand U4285 (N_4285,N_184,N_1771);
nand U4286 (N_4286,N_1856,N_2336);
and U4287 (N_4287,N_1862,N_502);
nor U4288 (N_4288,N_2228,N_189);
or U4289 (N_4289,N_1976,N_478);
nand U4290 (N_4290,N_1553,N_1208);
nand U4291 (N_4291,N_1203,N_575);
or U4292 (N_4292,N_437,N_975);
nor U4293 (N_4293,N_606,N_189);
nor U4294 (N_4294,N_947,N_2485);
or U4295 (N_4295,N_133,N_998);
nand U4296 (N_4296,N_1899,N_1885);
or U4297 (N_4297,N_827,N_621);
nor U4298 (N_4298,N_2486,N_2219);
nor U4299 (N_4299,N_1,N_665);
and U4300 (N_4300,N_264,N_435);
nor U4301 (N_4301,N_1302,N_198);
nand U4302 (N_4302,N_1935,N_926);
and U4303 (N_4303,N_552,N_2070);
nor U4304 (N_4304,N_245,N_588);
or U4305 (N_4305,N_1683,N_608);
nor U4306 (N_4306,N_1541,N_263);
nor U4307 (N_4307,N_2047,N_351);
or U4308 (N_4308,N_1394,N_540);
and U4309 (N_4309,N_962,N_1448);
and U4310 (N_4310,N_1923,N_1929);
and U4311 (N_4311,N_1909,N_286);
nor U4312 (N_4312,N_926,N_639);
or U4313 (N_4313,N_454,N_771);
nand U4314 (N_4314,N_730,N_534);
or U4315 (N_4315,N_432,N_458);
nand U4316 (N_4316,N_2077,N_1562);
nor U4317 (N_4317,N_1116,N_117);
nand U4318 (N_4318,N_2315,N_1384);
nor U4319 (N_4319,N_99,N_869);
nor U4320 (N_4320,N_157,N_1304);
nand U4321 (N_4321,N_1081,N_904);
and U4322 (N_4322,N_1971,N_1811);
or U4323 (N_4323,N_219,N_1039);
or U4324 (N_4324,N_182,N_2206);
and U4325 (N_4325,N_1202,N_624);
and U4326 (N_4326,N_1467,N_1263);
nor U4327 (N_4327,N_1636,N_1109);
and U4328 (N_4328,N_2258,N_1207);
and U4329 (N_4329,N_1266,N_1467);
nor U4330 (N_4330,N_174,N_0);
nand U4331 (N_4331,N_1083,N_1524);
or U4332 (N_4332,N_1966,N_348);
nand U4333 (N_4333,N_789,N_876);
nand U4334 (N_4334,N_1829,N_1285);
or U4335 (N_4335,N_1985,N_40);
or U4336 (N_4336,N_975,N_863);
or U4337 (N_4337,N_1613,N_1529);
and U4338 (N_4338,N_423,N_959);
nand U4339 (N_4339,N_268,N_2398);
nand U4340 (N_4340,N_2389,N_1104);
nand U4341 (N_4341,N_2309,N_156);
nor U4342 (N_4342,N_1235,N_1847);
or U4343 (N_4343,N_2406,N_2006);
nor U4344 (N_4344,N_1327,N_1059);
and U4345 (N_4345,N_570,N_100);
and U4346 (N_4346,N_88,N_1739);
and U4347 (N_4347,N_1869,N_1071);
nor U4348 (N_4348,N_160,N_1818);
nor U4349 (N_4349,N_344,N_2258);
or U4350 (N_4350,N_1502,N_1731);
or U4351 (N_4351,N_660,N_1442);
and U4352 (N_4352,N_609,N_632);
nor U4353 (N_4353,N_2222,N_391);
and U4354 (N_4354,N_838,N_562);
or U4355 (N_4355,N_19,N_1382);
xor U4356 (N_4356,N_1813,N_1737);
and U4357 (N_4357,N_1836,N_1202);
nand U4358 (N_4358,N_18,N_2118);
nand U4359 (N_4359,N_1422,N_1307);
nand U4360 (N_4360,N_1885,N_84);
and U4361 (N_4361,N_1603,N_1056);
and U4362 (N_4362,N_977,N_609);
or U4363 (N_4363,N_717,N_2290);
and U4364 (N_4364,N_1950,N_831);
or U4365 (N_4365,N_1760,N_2170);
and U4366 (N_4366,N_469,N_605);
or U4367 (N_4367,N_769,N_153);
and U4368 (N_4368,N_302,N_228);
and U4369 (N_4369,N_1231,N_2111);
nand U4370 (N_4370,N_1285,N_215);
nand U4371 (N_4371,N_580,N_1118);
and U4372 (N_4372,N_473,N_761);
or U4373 (N_4373,N_330,N_812);
or U4374 (N_4374,N_517,N_1395);
or U4375 (N_4375,N_1873,N_2467);
nand U4376 (N_4376,N_1026,N_1651);
nor U4377 (N_4377,N_2429,N_1426);
nor U4378 (N_4378,N_181,N_799);
or U4379 (N_4379,N_1659,N_1695);
or U4380 (N_4380,N_343,N_1481);
nor U4381 (N_4381,N_1811,N_2118);
nor U4382 (N_4382,N_1828,N_1959);
nand U4383 (N_4383,N_748,N_769);
nor U4384 (N_4384,N_602,N_1470);
and U4385 (N_4385,N_834,N_2239);
or U4386 (N_4386,N_1573,N_1038);
xnor U4387 (N_4387,N_584,N_352);
nand U4388 (N_4388,N_944,N_1153);
nand U4389 (N_4389,N_357,N_927);
nand U4390 (N_4390,N_1190,N_1427);
nor U4391 (N_4391,N_364,N_2308);
or U4392 (N_4392,N_18,N_36);
or U4393 (N_4393,N_1070,N_867);
or U4394 (N_4394,N_1000,N_1100);
or U4395 (N_4395,N_1724,N_1720);
nor U4396 (N_4396,N_1093,N_1695);
and U4397 (N_4397,N_1900,N_2384);
nor U4398 (N_4398,N_292,N_71);
and U4399 (N_4399,N_1612,N_1871);
and U4400 (N_4400,N_237,N_1265);
nor U4401 (N_4401,N_789,N_199);
or U4402 (N_4402,N_1211,N_1313);
and U4403 (N_4403,N_745,N_1694);
nor U4404 (N_4404,N_473,N_1532);
or U4405 (N_4405,N_1684,N_853);
nor U4406 (N_4406,N_1576,N_1936);
nor U4407 (N_4407,N_1784,N_424);
nor U4408 (N_4408,N_838,N_1614);
and U4409 (N_4409,N_2465,N_2151);
nand U4410 (N_4410,N_210,N_2350);
and U4411 (N_4411,N_1849,N_1527);
nand U4412 (N_4412,N_520,N_1383);
xnor U4413 (N_4413,N_436,N_1476);
nor U4414 (N_4414,N_1912,N_2066);
and U4415 (N_4415,N_1088,N_2293);
nor U4416 (N_4416,N_717,N_743);
and U4417 (N_4417,N_1785,N_1610);
or U4418 (N_4418,N_2426,N_830);
nand U4419 (N_4419,N_1691,N_5);
nand U4420 (N_4420,N_1327,N_639);
or U4421 (N_4421,N_1825,N_987);
and U4422 (N_4422,N_934,N_621);
nand U4423 (N_4423,N_1590,N_830);
nand U4424 (N_4424,N_1683,N_204);
xnor U4425 (N_4425,N_807,N_728);
or U4426 (N_4426,N_523,N_1212);
nand U4427 (N_4427,N_2343,N_1621);
nand U4428 (N_4428,N_1635,N_1432);
nor U4429 (N_4429,N_534,N_2318);
and U4430 (N_4430,N_247,N_2339);
nand U4431 (N_4431,N_2185,N_509);
or U4432 (N_4432,N_1698,N_2017);
nand U4433 (N_4433,N_1929,N_1151);
or U4434 (N_4434,N_469,N_153);
nand U4435 (N_4435,N_927,N_729);
nor U4436 (N_4436,N_1316,N_0);
nor U4437 (N_4437,N_353,N_638);
xor U4438 (N_4438,N_100,N_562);
nand U4439 (N_4439,N_1748,N_456);
or U4440 (N_4440,N_448,N_1655);
xnor U4441 (N_4441,N_356,N_2451);
or U4442 (N_4442,N_218,N_2325);
or U4443 (N_4443,N_1966,N_1996);
nand U4444 (N_4444,N_1795,N_1085);
nand U4445 (N_4445,N_318,N_593);
nor U4446 (N_4446,N_386,N_2088);
and U4447 (N_4447,N_288,N_813);
xnor U4448 (N_4448,N_1567,N_893);
nand U4449 (N_4449,N_1070,N_2152);
or U4450 (N_4450,N_1946,N_291);
or U4451 (N_4451,N_483,N_933);
nor U4452 (N_4452,N_1691,N_217);
nor U4453 (N_4453,N_2320,N_1899);
or U4454 (N_4454,N_1272,N_2061);
nor U4455 (N_4455,N_1079,N_1496);
and U4456 (N_4456,N_1084,N_624);
nor U4457 (N_4457,N_926,N_1788);
nor U4458 (N_4458,N_270,N_607);
nor U4459 (N_4459,N_656,N_464);
nand U4460 (N_4460,N_1323,N_2271);
and U4461 (N_4461,N_1786,N_56);
and U4462 (N_4462,N_1909,N_2233);
nor U4463 (N_4463,N_2278,N_1534);
and U4464 (N_4464,N_314,N_1308);
or U4465 (N_4465,N_425,N_774);
nor U4466 (N_4466,N_1808,N_1188);
nand U4467 (N_4467,N_2191,N_1188);
and U4468 (N_4468,N_2249,N_1627);
and U4469 (N_4469,N_1964,N_407);
and U4470 (N_4470,N_1416,N_2440);
and U4471 (N_4471,N_1113,N_2029);
and U4472 (N_4472,N_2040,N_18);
or U4473 (N_4473,N_1368,N_632);
xnor U4474 (N_4474,N_691,N_2045);
nand U4475 (N_4475,N_471,N_1755);
and U4476 (N_4476,N_262,N_1498);
nand U4477 (N_4477,N_2385,N_1338);
and U4478 (N_4478,N_1311,N_235);
and U4479 (N_4479,N_2087,N_843);
or U4480 (N_4480,N_152,N_1002);
and U4481 (N_4481,N_1133,N_991);
nand U4482 (N_4482,N_1539,N_2356);
nand U4483 (N_4483,N_2044,N_1535);
nor U4484 (N_4484,N_862,N_2059);
nand U4485 (N_4485,N_425,N_437);
nand U4486 (N_4486,N_1458,N_834);
or U4487 (N_4487,N_128,N_1169);
nand U4488 (N_4488,N_665,N_2412);
nand U4489 (N_4489,N_482,N_1096);
nor U4490 (N_4490,N_2247,N_717);
or U4491 (N_4491,N_817,N_1479);
and U4492 (N_4492,N_668,N_187);
and U4493 (N_4493,N_421,N_487);
or U4494 (N_4494,N_640,N_209);
and U4495 (N_4495,N_2011,N_1780);
or U4496 (N_4496,N_1762,N_1655);
and U4497 (N_4497,N_766,N_1191);
nor U4498 (N_4498,N_2141,N_1421);
or U4499 (N_4499,N_288,N_430);
nor U4500 (N_4500,N_506,N_747);
nor U4501 (N_4501,N_119,N_395);
and U4502 (N_4502,N_2423,N_612);
nand U4503 (N_4503,N_2181,N_2342);
nor U4504 (N_4504,N_634,N_1050);
nor U4505 (N_4505,N_1993,N_1125);
nor U4506 (N_4506,N_1781,N_1369);
or U4507 (N_4507,N_1201,N_2084);
nand U4508 (N_4508,N_1997,N_1040);
nand U4509 (N_4509,N_842,N_1719);
and U4510 (N_4510,N_1798,N_457);
or U4511 (N_4511,N_2481,N_1538);
nor U4512 (N_4512,N_1489,N_2020);
nor U4513 (N_4513,N_379,N_1772);
nand U4514 (N_4514,N_667,N_1723);
nor U4515 (N_4515,N_89,N_1647);
and U4516 (N_4516,N_1652,N_1688);
and U4517 (N_4517,N_848,N_250);
nor U4518 (N_4518,N_1546,N_1756);
or U4519 (N_4519,N_1765,N_1966);
nand U4520 (N_4520,N_1749,N_215);
nand U4521 (N_4521,N_1675,N_614);
nor U4522 (N_4522,N_249,N_2196);
nor U4523 (N_4523,N_160,N_2396);
or U4524 (N_4524,N_1772,N_81);
nand U4525 (N_4525,N_368,N_457);
nor U4526 (N_4526,N_2321,N_1951);
or U4527 (N_4527,N_1903,N_2042);
nand U4528 (N_4528,N_386,N_136);
or U4529 (N_4529,N_894,N_243);
nor U4530 (N_4530,N_1243,N_1437);
nor U4531 (N_4531,N_71,N_441);
or U4532 (N_4532,N_992,N_2193);
nor U4533 (N_4533,N_335,N_956);
or U4534 (N_4534,N_389,N_2291);
or U4535 (N_4535,N_891,N_105);
or U4536 (N_4536,N_1909,N_1397);
or U4537 (N_4537,N_514,N_865);
and U4538 (N_4538,N_1353,N_1380);
or U4539 (N_4539,N_34,N_1615);
nor U4540 (N_4540,N_1171,N_1662);
or U4541 (N_4541,N_740,N_1617);
nand U4542 (N_4542,N_2427,N_2072);
nor U4543 (N_4543,N_371,N_607);
nor U4544 (N_4544,N_781,N_737);
and U4545 (N_4545,N_1714,N_2462);
and U4546 (N_4546,N_1600,N_1404);
or U4547 (N_4547,N_473,N_366);
and U4548 (N_4548,N_2347,N_2253);
nor U4549 (N_4549,N_95,N_1971);
and U4550 (N_4550,N_2297,N_1519);
or U4551 (N_4551,N_13,N_937);
nand U4552 (N_4552,N_60,N_214);
nand U4553 (N_4553,N_1984,N_1885);
nor U4554 (N_4554,N_1600,N_682);
or U4555 (N_4555,N_1161,N_1108);
nand U4556 (N_4556,N_686,N_1604);
nor U4557 (N_4557,N_2461,N_1469);
or U4558 (N_4558,N_883,N_1726);
or U4559 (N_4559,N_1573,N_1089);
or U4560 (N_4560,N_1390,N_370);
nor U4561 (N_4561,N_2402,N_515);
or U4562 (N_4562,N_1655,N_60);
and U4563 (N_4563,N_1517,N_2201);
nor U4564 (N_4564,N_405,N_926);
nor U4565 (N_4565,N_1634,N_219);
and U4566 (N_4566,N_788,N_1565);
xor U4567 (N_4567,N_192,N_1962);
or U4568 (N_4568,N_2009,N_1706);
or U4569 (N_4569,N_2464,N_1838);
or U4570 (N_4570,N_479,N_1302);
and U4571 (N_4571,N_648,N_1255);
and U4572 (N_4572,N_194,N_847);
or U4573 (N_4573,N_1894,N_1834);
and U4574 (N_4574,N_1610,N_905);
nor U4575 (N_4575,N_1380,N_1207);
and U4576 (N_4576,N_250,N_2187);
or U4577 (N_4577,N_2182,N_577);
or U4578 (N_4578,N_512,N_2268);
xor U4579 (N_4579,N_427,N_1732);
or U4580 (N_4580,N_459,N_1943);
or U4581 (N_4581,N_591,N_240);
nor U4582 (N_4582,N_683,N_623);
nor U4583 (N_4583,N_918,N_784);
or U4584 (N_4584,N_908,N_329);
and U4585 (N_4585,N_2322,N_1177);
nand U4586 (N_4586,N_1920,N_1175);
nand U4587 (N_4587,N_622,N_2200);
or U4588 (N_4588,N_1864,N_1772);
and U4589 (N_4589,N_254,N_1686);
or U4590 (N_4590,N_2091,N_1733);
nor U4591 (N_4591,N_375,N_417);
nor U4592 (N_4592,N_2040,N_1973);
nor U4593 (N_4593,N_836,N_2163);
nand U4594 (N_4594,N_986,N_1248);
and U4595 (N_4595,N_714,N_26);
or U4596 (N_4596,N_2231,N_272);
nand U4597 (N_4597,N_27,N_1622);
and U4598 (N_4598,N_705,N_1400);
nor U4599 (N_4599,N_1780,N_1674);
and U4600 (N_4600,N_228,N_1920);
and U4601 (N_4601,N_1439,N_64);
or U4602 (N_4602,N_2007,N_329);
and U4603 (N_4603,N_17,N_2341);
nor U4604 (N_4604,N_816,N_202);
nand U4605 (N_4605,N_1633,N_789);
and U4606 (N_4606,N_1585,N_1999);
nand U4607 (N_4607,N_576,N_1679);
nor U4608 (N_4608,N_488,N_2396);
xnor U4609 (N_4609,N_80,N_2285);
and U4610 (N_4610,N_7,N_1752);
and U4611 (N_4611,N_2414,N_1934);
nor U4612 (N_4612,N_554,N_984);
nor U4613 (N_4613,N_984,N_888);
or U4614 (N_4614,N_553,N_1204);
nor U4615 (N_4615,N_125,N_2218);
nand U4616 (N_4616,N_1632,N_1036);
or U4617 (N_4617,N_361,N_1384);
nor U4618 (N_4618,N_1584,N_209);
and U4619 (N_4619,N_1855,N_354);
nand U4620 (N_4620,N_1069,N_1544);
and U4621 (N_4621,N_1116,N_2050);
and U4622 (N_4622,N_194,N_529);
or U4623 (N_4623,N_2339,N_2310);
and U4624 (N_4624,N_109,N_1762);
or U4625 (N_4625,N_668,N_1993);
or U4626 (N_4626,N_2498,N_2151);
and U4627 (N_4627,N_1343,N_334);
nand U4628 (N_4628,N_2189,N_118);
or U4629 (N_4629,N_1632,N_1666);
nor U4630 (N_4630,N_2291,N_2340);
or U4631 (N_4631,N_1133,N_230);
and U4632 (N_4632,N_403,N_1804);
and U4633 (N_4633,N_2272,N_76);
and U4634 (N_4634,N_1494,N_2234);
nor U4635 (N_4635,N_427,N_2251);
nor U4636 (N_4636,N_1829,N_1676);
or U4637 (N_4637,N_1152,N_1958);
nor U4638 (N_4638,N_380,N_973);
and U4639 (N_4639,N_1857,N_196);
or U4640 (N_4640,N_1097,N_394);
or U4641 (N_4641,N_2290,N_243);
nor U4642 (N_4642,N_1866,N_1524);
or U4643 (N_4643,N_931,N_1409);
or U4644 (N_4644,N_2037,N_1117);
nor U4645 (N_4645,N_79,N_2330);
or U4646 (N_4646,N_1072,N_772);
and U4647 (N_4647,N_1074,N_275);
or U4648 (N_4648,N_798,N_957);
and U4649 (N_4649,N_1372,N_98);
nor U4650 (N_4650,N_1057,N_1617);
and U4651 (N_4651,N_320,N_792);
nand U4652 (N_4652,N_951,N_2027);
or U4653 (N_4653,N_605,N_472);
nand U4654 (N_4654,N_1189,N_985);
nand U4655 (N_4655,N_1860,N_2036);
nand U4656 (N_4656,N_1672,N_2271);
or U4657 (N_4657,N_981,N_1493);
or U4658 (N_4658,N_751,N_546);
nor U4659 (N_4659,N_1393,N_1675);
nand U4660 (N_4660,N_1222,N_1806);
or U4661 (N_4661,N_1065,N_2480);
and U4662 (N_4662,N_834,N_983);
or U4663 (N_4663,N_796,N_860);
nand U4664 (N_4664,N_1816,N_414);
nor U4665 (N_4665,N_2370,N_2003);
or U4666 (N_4666,N_1144,N_45);
nor U4667 (N_4667,N_2322,N_511);
nor U4668 (N_4668,N_2398,N_1767);
or U4669 (N_4669,N_637,N_1043);
and U4670 (N_4670,N_1627,N_925);
nor U4671 (N_4671,N_1109,N_197);
nand U4672 (N_4672,N_741,N_2460);
nor U4673 (N_4673,N_1545,N_458);
nand U4674 (N_4674,N_2460,N_327);
nand U4675 (N_4675,N_1694,N_1612);
xnor U4676 (N_4676,N_72,N_872);
or U4677 (N_4677,N_1725,N_2349);
xnor U4678 (N_4678,N_2134,N_1514);
nand U4679 (N_4679,N_2437,N_539);
and U4680 (N_4680,N_2089,N_2425);
and U4681 (N_4681,N_2017,N_255);
nor U4682 (N_4682,N_1012,N_799);
and U4683 (N_4683,N_2114,N_347);
or U4684 (N_4684,N_2245,N_685);
nor U4685 (N_4685,N_2428,N_1688);
and U4686 (N_4686,N_1352,N_1823);
nor U4687 (N_4687,N_1233,N_771);
xor U4688 (N_4688,N_1833,N_1738);
or U4689 (N_4689,N_1944,N_65);
and U4690 (N_4690,N_576,N_2400);
nand U4691 (N_4691,N_810,N_751);
nor U4692 (N_4692,N_2401,N_2176);
nor U4693 (N_4693,N_1752,N_2410);
or U4694 (N_4694,N_521,N_1443);
nor U4695 (N_4695,N_206,N_303);
and U4696 (N_4696,N_2387,N_1645);
nand U4697 (N_4697,N_1526,N_285);
or U4698 (N_4698,N_1281,N_1886);
or U4699 (N_4699,N_2124,N_1635);
nand U4700 (N_4700,N_28,N_1973);
and U4701 (N_4701,N_1057,N_67);
nor U4702 (N_4702,N_401,N_1821);
and U4703 (N_4703,N_1718,N_2372);
nand U4704 (N_4704,N_660,N_2154);
nand U4705 (N_4705,N_34,N_505);
nand U4706 (N_4706,N_2452,N_1203);
nor U4707 (N_4707,N_1781,N_783);
or U4708 (N_4708,N_2452,N_2082);
nor U4709 (N_4709,N_829,N_1012);
or U4710 (N_4710,N_1763,N_2395);
and U4711 (N_4711,N_1104,N_2063);
xnor U4712 (N_4712,N_934,N_1319);
and U4713 (N_4713,N_1532,N_2326);
or U4714 (N_4714,N_883,N_282);
or U4715 (N_4715,N_1085,N_1370);
nor U4716 (N_4716,N_2122,N_406);
xor U4717 (N_4717,N_1480,N_1461);
nor U4718 (N_4718,N_1544,N_1703);
and U4719 (N_4719,N_1935,N_1087);
nor U4720 (N_4720,N_431,N_1769);
and U4721 (N_4721,N_80,N_1313);
nand U4722 (N_4722,N_290,N_1075);
and U4723 (N_4723,N_1648,N_1440);
nor U4724 (N_4724,N_1293,N_451);
nor U4725 (N_4725,N_2409,N_1540);
or U4726 (N_4726,N_2286,N_1831);
xnor U4727 (N_4727,N_13,N_1095);
nor U4728 (N_4728,N_2474,N_1083);
nor U4729 (N_4729,N_1301,N_105);
and U4730 (N_4730,N_1776,N_2080);
nor U4731 (N_4731,N_1409,N_1145);
or U4732 (N_4732,N_194,N_2002);
and U4733 (N_4733,N_1816,N_1542);
or U4734 (N_4734,N_709,N_2195);
or U4735 (N_4735,N_1922,N_2132);
nand U4736 (N_4736,N_2057,N_1380);
or U4737 (N_4737,N_152,N_397);
nand U4738 (N_4738,N_214,N_1735);
or U4739 (N_4739,N_2113,N_505);
nand U4740 (N_4740,N_932,N_2030);
or U4741 (N_4741,N_2439,N_2288);
or U4742 (N_4742,N_637,N_112);
nor U4743 (N_4743,N_84,N_934);
and U4744 (N_4744,N_1795,N_1186);
nor U4745 (N_4745,N_1315,N_901);
nor U4746 (N_4746,N_1264,N_1998);
and U4747 (N_4747,N_1051,N_2048);
or U4748 (N_4748,N_1359,N_1713);
or U4749 (N_4749,N_512,N_2310);
or U4750 (N_4750,N_1845,N_2380);
and U4751 (N_4751,N_982,N_350);
nand U4752 (N_4752,N_2065,N_1980);
nor U4753 (N_4753,N_2076,N_539);
and U4754 (N_4754,N_107,N_1269);
nor U4755 (N_4755,N_904,N_2033);
and U4756 (N_4756,N_1413,N_131);
and U4757 (N_4757,N_657,N_1278);
nor U4758 (N_4758,N_1394,N_2499);
nor U4759 (N_4759,N_922,N_1265);
nand U4760 (N_4760,N_1800,N_323);
nand U4761 (N_4761,N_1775,N_1391);
nor U4762 (N_4762,N_1507,N_1014);
or U4763 (N_4763,N_1375,N_826);
nand U4764 (N_4764,N_2208,N_78);
or U4765 (N_4765,N_1829,N_2154);
nor U4766 (N_4766,N_2490,N_1497);
nor U4767 (N_4767,N_546,N_1321);
nor U4768 (N_4768,N_849,N_1945);
nand U4769 (N_4769,N_706,N_1242);
and U4770 (N_4770,N_1698,N_1835);
and U4771 (N_4771,N_2077,N_1593);
or U4772 (N_4772,N_1365,N_573);
nor U4773 (N_4773,N_2408,N_988);
and U4774 (N_4774,N_2342,N_926);
and U4775 (N_4775,N_218,N_339);
nor U4776 (N_4776,N_1545,N_1352);
and U4777 (N_4777,N_1559,N_596);
nor U4778 (N_4778,N_747,N_362);
or U4779 (N_4779,N_154,N_2346);
or U4780 (N_4780,N_1404,N_2327);
or U4781 (N_4781,N_846,N_351);
nand U4782 (N_4782,N_1965,N_662);
nand U4783 (N_4783,N_384,N_1084);
or U4784 (N_4784,N_2412,N_1564);
and U4785 (N_4785,N_77,N_496);
and U4786 (N_4786,N_918,N_933);
or U4787 (N_4787,N_2255,N_1254);
or U4788 (N_4788,N_771,N_257);
nand U4789 (N_4789,N_1824,N_604);
nand U4790 (N_4790,N_57,N_1408);
nor U4791 (N_4791,N_702,N_191);
nand U4792 (N_4792,N_17,N_743);
and U4793 (N_4793,N_2229,N_2183);
and U4794 (N_4794,N_2144,N_1111);
or U4795 (N_4795,N_1064,N_1346);
or U4796 (N_4796,N_2256,N_301);
nand U4797 (N_4797,N_158,N_1576);
or U4798 (N_4798,N_466,N_555);
nand U4799 (N_4799,N_1404,N_1002);
nand U4800 (N_4800,N_1875,N_1788);
nand U4801 (N_4801,N_2395,N_1263);
nand U4802 (N_4802,N_1722,N_1615);
or U4803 (N_4803,N_206,N_1264);
xor U4804 (N_4804,N_1822,N_2433);
nand U4805 (N_4805,N_407,N_1673);
nor U4806 (N_4806,N_481,N_1930);
or U4807 (N_4807,N_401,N_836);
or U4808 (N_4808,N_621,N_929);
nand U4809 (N_4809,N_1256,N_1528);
nand U4810 (N_4810,N_1133,N_2376);
nand U4811 (N_4811,N_1446,N_1881);
or U4812 (N_4812,N_1890,N_15);
and U4813 (N_4813,N_2493,N_902);
or U4814 (N_4814,N_838,N_1523);
nor U4815 (N_4815,N_209,N_1920);
and U4816 (N_4816,N_1978,N_885);
and U4817 (N_4817,N_46,N_273);
or U4818 (N_4818,N_1874,N_637);
nor U4819 (N_4819,N_2319,N_1064);
and U4820 (N_4820,N_638,N_1058);
and U4821 (N_4821,N_1866,N_151);
or U4822 (N_4822,N_362,N_1902);
nand U4823 (N_4823,N_2407,N_1166);
nor U4824 (N_4824,N_851,N_1537);
nand U4825 (N_4825,N_2428,N_1366);
nor U4826 (N_4826,N_1946,N_609);
nor U4827 (N_4827,N_1066,N_1711);
and U4828 (N_4828,N_2320,N_1533);
and U4829 (N_4829,N_861,N_2459);
or U4830 (N_4830,N_2325,N_348);
or U4831 (N_4831,N_328,N_2449);
and U4832 (N_4832,N_314,N_679);
nand U4833 (N_4833,N_1612,N_415);
nor U4834 (N_4834,N_2028,N_482);
nand U4835 (N_4835,N_1383,N_736);
or U4836 (N_4836,N_1831,N_2467);
nand U4837 (N_4837,N_2276,N_921);
nor U4838 (N_4838,N_1795,N_158);
nor U4839 (N_4839,N_2108,N_2397);
or U4840 (N_4840,N_1468,N_890);
nor U4841 (N_4841,N_1063,N_245);
nor U4842 (N_4842,N_1764,N_1329);
and U4843 (N_4843,N_1220,N_1598);
xor U4844 (N_4844,N_990,N_886);
nand U4845 (N_4845,N_2216,N_555);
nor U4846 (N_4846,N_1165,N_1352);
and U4847 (N_4847,N_1543,N_2136);
or U4848 (N_4848,N_1571,N_1013);
nor U4849 (N_4849,N_269,N_1930);
or U4850 (N_4850,N_1747,N_2007);
nor U4851 (N_4851,N_117,N_320);
nor U4852 (N_4852,N_2089,N_842);
nand U4853 (N_4853,N_9,N_1150);
nor U4854 (N_4854,N_817,N_1359);
nand U4855 (N_4855,N_1874,N_2421);
and U4856 (N_4856,N_649,N_2133);
nand U4857 (N_4857,N_765,N_359);
and U4858 (N_4858,N_1897,N_1038);
and U4859 (N_4859,N_923,N_1358);
nand U4860 (N_4860,N_2125,N_246);
nand U4861 (N_4861,N_1055,N_1756);
or U4862 (N_4862,N_1704,N_291);
and U4863 (N_4863,N_927,N_2468);
nor U4864 (N_4864,N_234,N_1903);
or U4865 (N_4865,N_1113,N_1919);
nor U4866 (N_4866,N_2134,N_1539);
nand U4867 (N_4867,N_603,N_434);
or U4868 (N_4868,N_1224,N_1119);
or U4869 (N_4869,N_2158,N_944);
nand U4870 (N_4870,N_577,N_744);
or U4871 (N_4871,N_249,N_961);
or U4872 (N_4872,N_39,N_697);
nor U4873 (N_4873,N_282,N_1702);
and U4874 (N_4874,N_1192,N_1223);
nand U4875 (N_4875,N_1608,N_273);
and U4876 (N_4876,N_1159,N_652);
or U4877 (N_4877,N_1424,N_453);
and U4878 (N_4878,N_677,N_919);
and U4879 (N_4879,N_2152,N_1363);
and U4880 (N_4880,N_1745,N_2357);
or U4881 (N_4881,N_2089,N_191);
nand U4882 (N_4882,N_2257,N_1685);
nor U4883 (N_4883,N_335,N_585);
and U4884 (N_4884,N_1469,N_201);
and U4885 (N_4885,N_809,N_373);
nand U4886 (N_4886,N_316,N_1225);
nand U4887 (N_4887,N_716,N_1792);
and U4888 (N_4888,N_534,N_1277);
nor U4889 (N_4889,N_1244,N_272);
and U4890 (N_4890,N_793,N_2381);
nand U4891 (N_4891,N_1415,N_1210);
nand U4892 (N_4892,N_741,N_199);
nor U4893 (N_4893,N_454,N_256);
nand U4894 (N_4894,N_2163,N_787);
or U4895 (N_4895,N_2444,N_1552);
nand U4896 (N_4896,N_2141,N_1817);
and U4897 (N_4897,N_1253,N_2358);
nor U4898 (N_4898,N_496,N_1316);
and U4899 (N_4899,N_58,N_1031);
nand U4900 (N_4900,N_843,N_1510);
nand U4901 (N_4901,N_1190,N_1625);
nand U4902 (N_4902,N_1134,N_1758);
nand U4903 (N_4903,N_1739,N_2196);
or U4904 (N_4904,N_1309,N_1822);
nand U4905 (N_4905,N_974,N_124);
nand U4906 (N_4906,N_641,N_1653);
nor U4907 (N_4907,N_986,N_2122);
and U4908 (N_4908,N_243,N_446);
nor U4909 (N_4909,N_1976,N_538);
nand U4910 (N_4910,N_1728,N_594);
or U4911 (N_4911,N_949,N_2467);
or U4912 (N_4912,N_2199,N_2240);
nand U4913 (N_4913,N_975,N_546);
nand U4914 (N_4914,N_546,N_619);
xor U4915 (N_4915,N_801,N_1386);
nor U4916 (N_4916,N_1116,N_2229);
or U4917 (N_4917,N_1360,N_229);
or U4918 (N_4918,N_2349,N_2062);
or U4919 (N_4919,N_1389,N_779);
nand U4920 (N_4920,N_1789,N_612);
and U4921 (N_4921,N_2201,N_1660);
and U4922 (N_4922,N_1248,N_1986);
and U4923 (N_4923,N_1775,N_753);
nand U4924 (N_4924,N_184,N_135);
or U4925 (N_4925,N_1033,N_1310);
and U4926 (N_4926,N_1450,N_472);
nor U4927 (N_4927,N_1017,N_1896);
or U4928 (N_4928,N_1012,N_853);
nor U4929 (N_4929,N_1266,N_984);
xor U4930 (N_4930,N_182,N_1932);
xor U4931 (N_4931,N_2499,N_2123);
or U4932 (N_4932,N_306,N_1296);
or U4933 (N_4933,N_1612,N_2242);
or U4934 (N_4934,N_102,N_912);
nand U4935 (N_4935,N_1449,N_552);
and U4936 (N_4936,N_2412,N_691);
and U4937 (N_4937,N_74,N_1651);
nor U4938 (N_4938,N_106,N_2273);
nand U4939 (N_4939,N_333,N_180);
xnor U4940 (N_4940,N_960,N_2221);
nor U4941 (N_4941,N_832,N_40);
nand U4942 (N_4942,N_2119,N_1391);
or U4943 (N_4943,N_2003,N_205);
nor U4944 (N_4944,N_1217,N_1846);
and U4945 (N_4945,N_75,N_1870);
or U4946 (N_4946,N_2161,N_2136);
and U4947 (N_4947,N_753,N_20);
and U4948 (N_4948,N_1944,N_41);
or U4949 (N_4949,N_1351,N_1634);
and U4950 (N_4950,N_659,N_1635);
and U4951 (N_4951,N_1967,N_246);
nor U4952 (N_4952,N_1102,N_1000);
and U4953 (N_4953,N_1810,N_739);
and U4954 (N_4954,N_24,N_486);
or U4955 (N_4955,N_235,N_461);
and U4956 (N_4956,N_1431,N_728);
nor U4957 (N_4957,N_98,N_774);
and U4958 (N_4958,N_224,N_100);
and U4959 (N_4959,N_1124,N_2358);
nor U4960 (N_4960,N_2011,N_1767);
and U4961 (N_4961,N_886,N_368);
and U4962 (N_4962,N_232,N_929);
nor U4963 (N_4963,N_2305,N_1918);
and U4964 (N_4964,N_562,N_2024);
and U4965 (N_4965,N_966,N_1878);
nand U4966 (N_4966,N_2232,N_142);
nor U4967 (N_4967,N_36,N_536);
nor U4968 (N_4968,N_1495,N_2367);
nor U4969 (N_4969,N_1905,N_394);
and U4970 (N_4970,N_951,N_4);
nor U4971 (N_4971,N_1128,N_394);
or U4972 (N_4972,N_1537,N_1813);
and U4973 (N_4973,N_1131,N_1586);
nor U4974 (N_4974,N_162,N_2440);
nor U4975 (N_4975,N_89,N_437);
nand U4976 (N_4976,N_301,N_1610);
nand U4977 (N_4977,N_89,N_2160);
and U4978 (N_4978,N_1291,N_1583);
and U4979 (N_4979,N_1276,N_740);
or U4980 (N_4980,N_994,N_2335);
or U4981 (N_4981,N_1487,N_2278);
nand U4982 (N_4982,N_1393,N_2036);
nor U4983 (N_4983,N_1808,N_1475);
or U4984 (N_4984,N_1029,N_324);
nor U4985 (N_4985,N_2357,N_1756);
nand U4986 (N_4986,N_1728,N_1931);
nor U4987 (N_4987,N_264,N_873);
and U4988 (N_4988,N_1143,N_1876);
nor U4989 (N_4989,N_1870,N_1230);
or U4990 (N_4990,N_1799,N_1756);
or U4991 (N_4991,N_1502,N_2223);
and U4992 (N_4992,N_843,N_1069);
nand U4993 (N_4993,N_1325,N_1261);
or U4994 (N_4994,N_441,N_532);
or U4995 (N_4995,N_2120,N_1484);
nor U4996 (N_4996,N_190,N_1345);
nand U4997 (N_4997,N_2166,N_2336);
nand U4998 (N_4998,N_1405,N_806);
or U4999 (N_4999,N_1594,N_373);
or UO_0 (O_0,N_3501,N_2829);
and UO_1 (O_1,N_4309,N_4022);
and UO_2 (O_2,N_4796,N_3875);
nand UO_3 (O_3,N_4983,N_3022);
xor UO_4 (O_4,N_4835,N_4499);
nor UO_5 (O_5,N_3744,N_4545);
nand UO_6 (O_6,N_3298,N_3086);
and UO_7 (O_7,N_2730,N_3861);
and UO_8 (O_8,N_4413,N_3798);
nor UO_9 (O_9,N_3180,N_3115);
and UO_10 (O_10,N_4651,N_2726);
nor UO_11 (O_11,N_4311,N_4159);
nor UO_12 (O_12,N_3012,N_4098);
nand UO_13 (O_13,N_4789,N_2660);
nor UO_14 (O_14,N_4711,N_3630);
or UO_15 (O_15,N_2702,N_4403);
and UO_16 (O_16,N_2508,N_4025);
or UO_17 (O_17,N_2852,N_3153);
and UO_18 (O_18,N_3128,N_4552);
nor UO_19 (O_19,N_2579,N_3358);
and UO_20 (O_20,N_4458,N_3285);
nand UO_21 (O_21,N_3050,N_4772);
or UO_22 (O_22,N_3531,N_4169);
and UO_23 (O_23,N_3402,N_4118);
nand UO_24 (O_24,N_3160,N_2911);
nor UO_25 (O_25,N_3430,N_3333);
or UO_26 (O_26,N_4503,N_2632);
nor UO_27 (O_27,N_3908,N_4057);
nor UO_28 (O_28,N_4380,N_2716);
nor UO_29 (O_29,N_2907,N_2830);
or UO_30 (O_30,N_3107,N_4834);
nand UO_31 (O_31,N_4748,N_2575);
or UO_32 (O_32,N_4707,N_4747);
and UO_33 (O_33,N_4168,N_3445);
nor UO_34 (O_34,N_2849,N_4832);
nand UO_35 (O_35,N_2780,N_3041);
and UO_36 (O_36,N_2609,N_3222);
and UO_37 (O_37,N_4086,N_4521);
nand UO_38 (O_38,N_3366,N_3242);
or UO_39 (O_39,N_4951,N_3843);
and UO_40 (O_40,N_4213,N_3959);
and UO_41 (O_41,N_3990,N_4028);
nand UO_42 (O_42,N_4580,N_4563);
nand UO_43 (O_43,N_2885,N_3530);
nor UO_44 (O_44,N_3880,N_3591);
nand UO_45 (O_45,N_3749,N_2936);
nand UO_46 (O_46,N_3628,N_2765);
nor UO_47 (O_47,N_4797,N_3037);
or UO_48 (O_48,N_4941,N_3790);
and UO_49 (O_49,N_2693,N_3347);
nor UO_50 (O_50,N_3925,N_3730);
nor UO_51 (O_51,N_4722,N_4248);
nand UO_52 (O_52,N_4668,N_4473);
and UO_53 (O_53,N_3699,N_4676);
nor UO_54 (O_54,N_3669,N_4558);
nand UO_55 (O_55,N_3439,N_4216);
or UO_56 (O_56,N_3123,N_3914);
nor UO_57 (O_57,N_2679,N_3952);
and UO_58 (O_58,N_3794,N_2782);
nor UO_59 (O_59,N_2950,N_3195);
nand UO_60 (O_60,N_3583,N_4725);
nand UO_61 (O_61,N_3559,N_2601);
and UO_62 (O_62,N_3849,N_2640);
nand UO_63 (O_63,N_4302,N_4140);
xor UO_64 (O_64,N_4001,N_4987);
or UO_65 (O_65,N_2619,N_4911);
or UO_66 (O_66,N_4497,N_4562);
nor UO_67 (O_67,N_4648,N_2896);
nor UO_68 (O_68,N_2736,N_4986);
nor UO_69 (O_69,N_4122,N_2733);
or UO_70 (O_70,N_4909,N_3399);
nor UO_71 (O_71,N_2560,N_4051);
and UO_72 (O_72,N_4131,N_3655);
and UO_73 (O_73,N_3263,N_3103);
or UO_74 (O_74,N_3337,N_4298);
nand UO_75 (O_75,N_3122,N_2654);
and UO_76 (O_76,N_4085,N_4915);
or UO_77 (O_77,N_3136,N_3045);
nand UO_78 (O_78,N_3205,N_4523);
nand UO_79 (O_79,N_4448,N_2720);
nand UO_80 (O_80,N_2751,N_4078);
and UO_81 (O_81,N_3926,N_2824);
nand UO_82 (O_82,N_2822,N_4259);
and UO_83 (O_83,N_4761,N_4039);
nand UO_84 (O_84,N_2588,N_2664);
nor UO_85 (O_85,N_4030,N_3408);
nor UO_86 (O_86,N_3443,N_4874);
xnor UO_87 (O_87,N_4441,N_3735);
nor UO_88 (O_88,N_3704,N_4970);
nand UO_89 (O_89,N_3563,N_4220);
nand UO_90 (O_90,N_2645,N_2668);
or UO_91 (O_91,N_4727,N_4378);
or UO_92 (O_92,N_3818,N_3994);
and UO_93 (O_93,N_4500,N_3345);
and UO_94 (O_94,N_2594,N_2954);
or UO_95 (O_95,N_2727,N_2813);
or UO_96 (O_96,N_3824,N_2945);
nor UO_97 (O_97,N_4262,N_2825);
xor UO_98 (O_98,N_4253,N_4179);
or UO_99 (O_99,N_2873,N_2859);
nor UO_100 (O_100,N_2530,N_4593);
nand UO_101 (O_101,N_4454,N_3762);
or UO_102 (O_102,N_4640,N_3778);
nand UO_103 (O_103,N_2924,N_4582);
xor UO_104 (O_104,N_4605,N_3163);
nand UO_105 (O_105,N_3424,N_3062);
and UO_106 (O_106,N_3309,N_3418);
nand UO_107 (O_107,N_2877,N_2784);
and UO_108 (O_108,N_4598,N_4757);
nor UO_109 (O_109,N_4330,N_4694);
nor UO_110 (O_110,N_3475,N_2909);
xnor UO_111 (O_111,N_2631,N_2744);
and UO_112 (O_112,N_3003,N_3685);
or UO_113 (O_113,N_2799,N_3519);
or UO_114 (O_114,N_4289,N_2977);
and UO_115 (O_115,N_3272,N_2797);
and UO_116 (O_116,N_3457,N_4774);
and UO_117 (O_117,N_3265,N_4898);
or UO_118 (O_118,N_4799,N_3986);
nand UO_119 (O_119,N_4342,N_3962);
or UO_120 (O_120,N_3944,N_3703);
and UO_121 (O_121,N_3391,N_4524);
nand UO_122 (O_122,N_3797,N_4247);
nand UO_123 (O_123,N_4764,N_3208);
or UO_124 (O_124,N_3077,N_3888);
nor UO_125 (O_125,N_4869,N_4218);
nor UO_126 (O_126,N_3776,N_4755);
nor UO_127 (O_127,N_4264,N_4902);
and UO_128 (O_128,N_4161,N_4867);
nor UO_129 (O_129,N_4080,N_4099);
nor UO_130 (O_130,N_3598,N_3293);
or UO_131 (O_131,N_3404,N_3052);
or UO_132 (O_132,N_3460,N_2515);
nor UO_133 (O_133,N_4409,N_3377);
xnor UO_134 (O_134,N_4044,N_3226);
nand UO_135 (O_135,N_2567,N_3188);
nor UO_136 (O_136,N_4730,N_3589);
or UO_137 (O_137,N_2691,N_4931);
or UO_138 (O_138,N_3711,N_3639);
nand UO_139 (O_139,N_4549,N_4621);
nand UO_140 (O_140,N_4632,N_4176);
and UO_141 (O_141,N_3436,N_2966);
and UO_142 (O_142,N_4815,N_3795);
nor UO_143 (O_143,N_4417,N_4925);
or UO_144 (O_144,N_3532,N_4816);
and UO_145 (O_145,N_3577,N_3520);
nand UO_146 (O_146,N_3977,N_3246);
nor UO_147 (O_147,N_4003,N_3650);
and UO_148 (O_148,N_3978,N_3374);
nand UO_149 (O_149,N_4871,N_3874);
nor UO_150 (O_150,N_4254,N_4575);
or UO_151 (O_151,N_4241,N_3419);
nand UO_152 (O_152,N_4634,N_3613);
nor UO_153 (O_153,N_2843,N_3736);
and UO_154 (O_154,N_3481,N_2621);
nand UO_155 (O_155,N_2923,N_3886);
and UO_156 (O_156,N_3466,N_4995);
or UO_157 (O_157,N_4146,N_3255);
nor UO_158 (O_158,N_3148,N_3585);
nor UO_159 (O_159,N_4617,N_4900);
xnor UO_160 (O_160,N_4297,N_3913);
nor UO_161 (O_161,N_3689,N_4397);
xnor UO_162 (O_162,N_4574,N_3276);
nor UO_163 (O_163,N_4056,N_3068);
or UO_164 (O_164,N_2522,N_3663);
nand UO_165 (O_165,N_2613,N_4372);
nor UO_166 (O_166,N_3756,N_3879);
nor UO_167 (O_167,N_2858,N_4536);
nand UO_168 (O_168,N_3158,N_3516);
nand UO_169 (O_169,N_4611,N_3070);
nand UO_170 (O_170,N_4184,N_2686);
nor UO_171 (O_171,N_4328,N_3599);
and UO_172 (O_172,N_3260,N_2552);
nor UO_173 (O_173,N_4669,N_4758);
or UO_174 (O_174,N_4148,N_2842);
nor UO_175 (O_175,N_4767,N_4106);
nor UO_176 (O_176,N_3437,N_3827);
or UO_177 (O_177,N_2935,N_3814);
or UO_178 (O_178,N_3019,N_4561);
and UO_179 (O_179,N_3779,N_2891);
or UO_180 (O_180,N_4720,N_4765);
and UO_181 (O_181,N_2925,N_2856);
nor UO_182 (O_182,N_4917,N_4944);
nand UO_183 (O_183,N_3116,N_4332);
nand UO_184 (O_184,N_4233,N_4000);
nor UO_185 (O_185,N_3336,N_3348);
xor UO_186 (O_186,N_2558,N_4888);
nand UO_187 (O_187,N_2731,N_4968);
and UO_188 (O_188,N_3393,N_4178);
and UO_189 (O_189,N_2772,N_4349);
nand UO_190 (O_190,N_2650,N_4471);
nand UO_191 (O_191,N_3970,N_3090);
and UO_192 (O_192,N_3975,N_4556);
or UO_193 (O_193,N_4809,N_4736);
nor UO_194 (O_194,N_2682,N_2685);
or UO_195 (O_195,N_3834,N_4418);
nand UO_196 (O_196,N_4113,N_4134);
and UO_197 (O_197,N_3984,N_4892);
xnor UO_198 (O_198,N_3282,N_4541);
nand UO_199 (O_199,N_3627,N_4513);
and UO_200 (O_200,N_4187,N_4101);
and UO_201 (O_201,N_3937,N_4196);
nor UO_202 (O_202,N_2637,N_4845);
nand UO_203 (O_203,N_3965,N_3609);
and UO_204 (O_204,N_4590,N_4235);
or UO_205 (O_205,N_4399,N_3513);
nand UO_206 (O_206,N_4896,N_3331);
and UO_207 (O_207,N_3968,N_3018);
xnor UO_208 (O_208,N_4875,N_3887);
and UO_209 (O_209,N_4637,N_3787);
nor UO_210 (O_210,N_4933,N_3344);
nand UO_211 (O_211,N_3229,N_2596);
nor UO_212 (O_212,N_4319,N_3054);
nor UO_213 (O_213,N_3771,N_4386);
nand UO_214 (O_214,N_3511,N_4444);
nor UO_215 (O_215,N_3810,N_2819);
nand UO_216 (O_216,N_3130,N_4528);
and UO_217 (O_217,N_4191,N_4189);
and UO_218 (O_218,N_3194,N_3184);
nor UO_219 (O_219,N_4864,N_4786);
and UO_220 (O_220,N_3141,N_4496);
nand UO_221 (O_221,N_4245,N_3026);
and UO_222 (O_222,N_3643,N_3261);
nand UO_223 (O_223,N_4876,N_2624);
and UO_224 (O_224,N_4826,N_4509);
nor UO_225 (O_225,N_4599,N_4618);
and UO_226 (O_226,N_4703,N_4004);
nand UO_227 (O_227,N_4701,N_4020);
nor UO_228 (O_228,N_3409,N_4132);
nor UO_229 (O_229,N_4569,N_3215);
nor UO_230 (O_230,N_4323,N_4103);
or UO_231 (O_231,N_2868,N_3676);
or UO_232 (O_232,N_4224,N_2889);
nor UO_233 (O_233,N_3239,N_4863);
and UO_234 (O_234,N_3243,N_2996);
and UO_235 (O_235,N_3151,N_4540);
nor UO_236 (O_236,N_3218,N_3316);
or UO_237 (O_237,N_4491,N_3584);
nor UO_238 (O_238,N_4303,N_4534);
nand UO_239 (O_239,N_4155,N_4287);
nor UO_240 (O_240,N_4808,N_2749);
and UO_241 (O_241,N_4973,N_2673);
or UO_242 (O_242,N_3918,N_3044);
or UO_243 (O_243,N_2671,N_3600);
nand UO_244 (O_244,N_3710,N_4936);
nor UO_245 (O_245,N_2748,N_3998);
nor UO_246 (O_246,N_2742,N_3606);
nor UO_247 (O_247,N_3433,N_4127);
nor UO_248 (O_248,N_4859,N_4962);
or UO_249 (O_249,N_2993,N_2745);
nor UO_250 (O_250,N_3109,N_3720);
nor UO_251 (O_251,N_3983,N_3210);
nor UO_252 (O_252,N_4460,N_4265);
nand UO_253 (O_253,N_3456,N_3523);
and UO_254 (O_254,N_4778,N_3748);
or UO_255 (O_255,N_3259,N_3200);
or UO_256 (O_256,N_4827,N_3621);
nor UO_257 (O_257,N_3682,N_3321);
nor UO_258 (O_258,N_3414,N_4204);
and UO_259 (O_259,N_3181,N_4948);
or UO_260 (O_260,N_4715,N_4501);
or UO_261 (O_261,N_4147,N_4836);
or UO_262 (O_262,N_3167,N_4719);
nor UO_263 (O_263,N_4785,N_2545);
nand UO_264 (O_264,N_3791,N_3576);
and UO_265 (O_265,N_4677,N_4449);
nand UO_266 (O_266,N_2994,N_2520);
nand UO_267 (O_267,N_3072,N_2944);
nand UO_268 (O_268,N_2837,N_4457);
or UO_269 (O_269,N_4337,N_3601);
or UO_270 (O_270,N_4985,N_4295);
or UO_271 (O_271,N_4801,N_4046);
nor UO_272 (O_272,N_3468,N_3853);
nand UO_273 (O_273,N_3830,N_3479);
nor UO_274 (O_274,N_3881,N_4263);
nand UO_275 (O_275,N_3939,N_3949);
and UO_276 (O_276,N_3948,N_4365);
nand UO_277 (O_277,N_4313,N_3346);
and UO_278 (O_278,N_3750,N_4692);
or UO_279 (O_279,N_3995,N_3334);
or UO_280 (O_280,N_2962,N_4307);
nand UO_281 (O_281,N_3774,N_4899);
nor UO_282 (O_282,N_4943,N_3035);
and UO_283 (O_283,N_4745,N_3610);
nand UO_284 (O_284,N_3595,N_3607);
nand UO_285 (O_285,N_3159,N_2697);
nor UO_286 (O_286,N_4726,N_3847);
nand UO_287 (O_287,N_2568,N_3596);
and UO_288 (O_288,N_3821,N_4354);
xnor UO_289 (O_289,N_2657,N_3075);
or UO_290 (O_290,N_3800,N_4505);
nand UO_291 (O_291,N_4773,N_3111);
nand UO_292 (O_292,N_4423,N_4947);
and UO_293 (O_293,N_2592,N_2722);
nand UO_294 (O_294,N_3693,N_2658);
and UO_295 (O_295,N_3283,N_2655);
and UO_296 (O_296,N_4824,N_4697);
nand UO_297 (O_297,N_4308,N_3547);
and UO_298 (O_298,N_3248,N_2959);
and UO_299 (O_299,N_2893,N_2602);
nor UO_300 (O_300,N_2732,N_3946);
nor UO_301 (O_301,N_2681,N_3190);
nand UO_302 (O_302,N_3864,N_4410);
and UO_303 (O_303,N_4841,N_4953);
and UO_304 (O_304,N_4777,N_3237);
nor UO_305 (O_305,N_3973,N_3296);
xor UO_306 (O_306,N_2978,N_4193);
and UO_307 (O_307,N_4811,N_4183);
nor UO_308 (O_308,N_2612,N_3241);
and UO_309 (O_309,N_4150,N_3397);
and UO_310 (O_310,N_3979,N_4489);
or UO_311 (O_311,N_3486,N_2649);
nand UO_312 (O_312,N_3139,N_2541);
and UO_313 (O_313,N_4729,N_3993);
nand UO_314 (O_314,N_2502,N_3114);
or UO_315 (O_315,N_2792,N_4861);
nor UO_316 (O_316,N_4718,N_4642);
xnor UO_317 (O_317,N_3240,N_4084);
or UO_318 (O_318,N_3329,N_3189);
nor UO_319 (O_319,N_3008,N_3212);
nor UO_320 (O_320,N_4604,N_3838);
or UO_321 (O_321,N_3300,N_4662);
nand UO_322 (O_322,N_3804,N_4770);
nand UO_323 (O_323,N_3562,N_4011);
nor UO_324 (O_324,N_3976,N_3608);
nand UO_325 (O_325,N_4108,N_3653);
nor UO_326 (O_326,N_3429,N_3777);
and UO_327 (O_327,N_2952,N_3383);
nand UO_328 (O_328,N_4325,N_2513);
nand UO_329 (O_329,N_2855,N_4435);
or UO_330 (O_330,N_4924,N_2884);
and UO_331 (O_331,N_3622,N_3634);
nor UO_332 (O_332,N_3936,N_3647);
nor UO_333 (O_333,N_4753,N_4504);
nor UO_334 (O_334,N_3903,N_3286);
nor UO_335 (O_335,N_3361,N_3264);
and UO_336 (O_336,N_4206,N_4320);
and UO_337 (O_337,N_2740,N_4405);
nor UO_338 (O_338,N_3058,N_4043);
and UO_339 (O_339,N_2587,N_3500);
nand UO_340 (O_340,N_2647,N_4272);
nor UO_341 (O_341,N_3105,N_3413);
or UO_342 (O_342,N_3724,N_4539);
nand UO_343 (O_343,N_4316,N_3097);
and UO_344 (O_344,N_2960,N_3758);
and UO_345 (O_345,N_4942,N_3769);
and UO_346 (O_346,N_2768,N_2965);
nor UO_347 (O_347,N_4596,N_2844);
and UO_348 (O_348,N_4483,N_4194);
nand UO_349 (O_349,N_3182,N_2938);
nor UO_350 (O_350,N_3575,N_3572);
and UO_351 (O_351,N_2922,N_2672);
nor UO_352 (O_352,N_3343,N_2881);
nor UO_353 (O_353,N_3071,N_3290);
and UO_354 (O_354,N_3892,N_4088);
nand UO_355 (O_355,N_2548,N_4484);
nand UO_356 (O_356,N_3665,N_4097);
nor UO_357 (O_357,N_3533,N_4436);
or UO_358 (O_358,N_4293,N_4362);
and UO_359 (O_359,N_3660,N_4520);
or UO_360 (O_360,N_3506,N_4731);
nand UO_361 (O_361,N_2759,N_4243);
nor UO_362 (O_362,N_3502,N_3691);
and UO_363 (O_363,N_3025,N_2539);
or UO_364 (O_364,N_3542,N_4100);
nand UO_365 (O_365,N_2648,N_2912);
or UO_366 (O_366,N_3024,N_2800);
or UO_367 (O_367,N_4890,N_3406);
or UO_368 (O_368,N_3680,N_2803);
nor UO_369 (O_369,N_3741,N_4989);
or UO_370 (O_370,N_3742,N_3203);
nor UO_371 (O_371,N_2516,N_3121);
and UO_372 (O_372,N_2526,N_3192);
or UO_373 (O_373,N_4273,N_4230);
nor UO_374 (O_374,N_2937,N_2951);
nor UO_375 (O_375,N_3177,N_2576);
nor UO_376 (O_376,N_3927,N_2721);
or UO_377 (O_377,N_3225,N_4597);
nand UO_378 (O_378,N_2779,N_3485);
or UO_379 (O_379,N_4568,N_2525);
and UO_380 (O_380,N_4477,N_2554);
nand UO_381 (O_381,N_2713,N_4762);
or UO_382 (O_382,N_3328,N_4978);
nand UO_383 (O_383,N_3303,N_3876);
xnor UO_384 (O_384,N_4291,N_4017);
and UO_385 (O_385,N_4833,N_3659);
nand UO_386 (O_386,N_2968,N_2943);
xnor UO_387 (O_387,N_3764,N_3270);
and UO_388 (O_388,N_3015,N_2862);
or UO_389 (O_389,N_3027,N_4201);
and UO_390 (O_390,N_2556,N_4688);
nor UO_391 (O_391,N_4304,N_4361);
nor UO_392 (O_392,N_2614,N_2642);
or UO_393 (O_393,N_4355,N_3185);
nor UO_394 (O_394,N_2633,N_3118);
nor UO_395 (O_395,N_4087,N_4649);
or UO_396 (O_396,N_3958,N_3698);
nand UO_397 (O_397,N_3694,N_4453);
nand UO_398 (O_398,N_4373,N_2967);
nor UO_399 (O_399,N_4737,N_2901);
nand UO_400 (O_400,N_2916,N_3057);
nand UO_401 (O_401,N_3157,N_3451);
or UO_402 (O_402,N_4884,N_2628);
nor UO_403 (O_403,N_2723,N_2564);
nor UO_404 (O_404,N_3852,N_4467);
nor UO_405 (O_405,N_4881,N_3354);
and UO_406 (O_406,N_3016,N_3236);
and UO_407 (O_407,N_4389,N_3088);
or UO_408 (O_408,N_4974,N_3480);
nor UO_409 (O_409,N_4734,N_2783);
nor UO_410 (O_410,N_3631,N_2984);
or UO_411 (O_411,N_3349,N_4228);
nor UO_412 (O_412,N_3076,N_3911);
nor UO_413 (O_413,N_3102,N_4069);
nor UO_414 (O_414,N_3510,N_2687);
nor UO_415 (O_415,N_3868,N_2809);
or UO_416 (O_416,N_2598,N_3472);
or UO_417 (O_417,N_3878,N_4519);
or UO_418 (O_418,N_4091,N_4434);
and UO_419 (O_419,N_4872,N_2930);
and UO_420 (O_420,N_4343,N_4588);
and UO_421 (O_421,N_4339,N_3793);
and UO_422 (O_422,N_3751,N_4065);
nor UO_423 (O_423,N_4286,N_3169);
and UO_424 (O_424,N_4465,N_4322);
nor UO_425 (O_425,N_2955,N_3183);
and UO_426 (O_426,N_4493,N_4935);
nor UO_427 (O_427,N_3330,N_4795);
nand UO_428 (O_428,N_2698,N_3517);
nand UO_429 (O_429,N_2910,N_4638);
or UO_430 (O_430,N_2734,N_3840);
nand UO_431 (O_431,N_4222,N_3933);
nand UO_432 (O_432,N_4932,N_2865);
nand UO_433 (O_433,N_3119,N_4082);
nor UO_434 (O_434,N_3005,N_3785);
nand UO_435 (O_435,N_2949,N_4526);
or UO_436 (O_436,N_3594,N_3524);
or UO_437 (O_437,N_4447,N_2543);
and UO_438 (O_438,N_4984,N_4712);
or UO_439 (O_439,N_3924,N_3431);
nand UO_440 (O_440,N_2934,N_2607);
nand UO_441 (O_441,N_3557,N_2553);
nand UO_442 (O_442,N_2521,N_4223);
nor UO_443 (O_443,N_3362,N_4026);
and UO_444 (O_444,N_3454,N_3981);
and UO_445 (O_445,N_2665,N_3483);
or UO_446 (O_446,N_4172,N_3644);
or UO_447 (O_447,N_4175,N_4988);
nor UO_448 (O_448,N_4188,N_3256);
nor UO_449 (O_449,N_3219,N_2848);
and UO_450 (O_450,N_4455,N_3206);
nand UO_451 (O_451,N_4480,N_3389);
or UO_452 (O_452,N_3854,N_3235);
nor UO_453 (O_453,N_4914,N_4527);
nand UO_454 (O_454,N_4716,N_3214);
or UO_455 (O_455,N_2920,N_3898);
nor UO_456 (O_456,N_3900,N_4553);
and UO_457 (O_457,N_4475,N_2636);
nor UO_458 (O_458,N_4687,N_3311);
or UO_459 (O_459,N_4255,N_4693);
nor UO_460 (O_460,N_3988,N_4421);
nand UO_461 (O_461,N_4584,N_2703);
and UO_462 (O_462,N_3964,N_2611);
nand UO_463 (O_463,N_4256,N_3491);
or UO_464 (O_464,N_3357,N_4671);
nand UO_465 (O_465,N_2763,N_4390);
and UO_466 (O_466,N_4269,N_4837);
nand UO_467 (O_467,N_2927,N_4416);
or UO_468 (O_468,N_4570,N_3266);
nor UO_469 (O_469,N_2917,N_4242);
nor UO_470 (O_470,N_3503,N_4829);
nand UO_471 (O_471,N_4476,N_2817);
xnor UO_472 (O_472,N_2595,N_4958);
or UO_473 (O_473,N_3476,N_4016);
or UO_474 (O_474,N_3733,N_4522);
nand UO_475 (O_475,N_3172,N_4428);
or UO_476 (O_476,N_3294,N_3780);
nand UO_477 (O_477,N_4672,N_4756);
and UO_478 (O_478,N_4840,N_2690);
nor UO_479 (O_479,N_3705,N_3895);
nand UO_480 (O_480,N_3143,N_2975);
nand UO_481 (O_481,N_4959,N_2915);
and UO_482 (O_482,N_3106,N_3681);
or UO_483 (O_483,N_3816,N_2528);
nor UO_484 (O_484,N_2610,N_2603);
nand UO_485 (O_485,N_4200,N_2961);
nand UO_486 (O_486,N_3390,N_4754);
nor UO_487 (O_487,N_4893,N_3497);
nor UO_488 (O_488,N_4076,N_4581);
and UO_489 (O_489,N_3267,N_3568);
xnor UO_490 (O_490,N_3561,N_4049);
or UO_491 (O_491,N_2919,N_4227);
and UO_492 (O_492,N_3550,N_4624);
and UO_493 (O_493,N_3801,N_3269);
xnor UO_494 (O_494,N_3438,N_4803);
nand UO_495 (O_495,N_2752,N_3310);
xor UO_496 (O_496,N_4572,N_4414);
nor UO_497 (O_497,N_3799,N_3380);
nor UO_498 (O_498,N_4197,N_2953);
and UO_499 (O_499,N_2990,N_3862);
nor UO_500 (O_500,N_3815,N_3142);
and UO_501 (O_501,N_4019,N_4154);
nor UO_502 (O_502,N_3325,N_3731);
or UO_503 (O_503,N_4771,N_4321);
or UO_504 (O_504,N_4283,N_4535);
and UO_505 (O_505,N_2563,N_4766);
nor UO_506 (O_506,N_4928,N_4680);
or UO_507 (O_507,N_4260,N_3618);
nand UO_508 (O_508,N_4398,N_2957);
or UO_509 (O_509,N_3001,N_4190);
nand UO_510 (O_510,N_3386,N_3061);
nor UO_511 (O_511,N_3991,N_4905);
nand UO_512 (O_512,N_3202,N_2666);
nand UO_513 (O_513,N_4622,N_4865);
nand UO_514 (O_514,N_4271,N_4895);
or UO_515 (O_515,N_3906,N_4683);
nor UO_516 (O_516,N_3508,N_4266);
and UO_517 (O_517,N_3478,N_2771);
nand UO_518 (O_518,N_2898,N_2503);
nor UO_519 (O_519,N_2766,N_2675);
or UO_520 (O_520,N_2683,N_2867);
or UO_521 (O_521,N_4125,N_4395);
and UO_522 (O_522,N_4429,N_3244);
and UO_523 (O_523,N_3696,N_3857);
and UO_524 (O_524,N_3448,N_3387);
and UO_525 (O_525,N_4252,N_3865);
and UO_526 (O_526,N_4877,N_4042);
nor UO_527 (O_527,N_3234,N_2656);
xor UO_528 (O_528,N_2827,N_2581);
nor UO_529 (O_529,N_4721,N_4631);
or UO_530 (O_530,N_2578,N_4063);
xnor UO_531 (O_531,N_4600,N_2832);
nor UO_532 (O_532,N_4284,N_2789);
nand UO_533 (O_533,N_2841,N_3543);
or UO_534 (O_534,N_4744,N_4609);
nor UO_535 (O_535,N_3224,N_2987);
nor UO_536 (O_536,N_4024,N_3187);
nand UO_537 (O_537,N_3275,N_3658);
nand UO_538 (O_538,N_4661,N_3851);
or UO_539 (O_539,N_3807,N_3232);
or UO_540 (O_540,N_3537,N_3211);
nand UO_541 (O_541,N_3193,N_2963);
or UO_542 (O_542,N_4461,N_3761);
and UO_543 (O_543,N_3972,N_4806);
nand UO_544 (O_544,N_4684,N_3421);
nor UO_545 (O_545,N_3825,N_3565);
nor UO_546 (O_546,N_4424,N_4285);
and UO_547 (O_547,N_4401,N_4883);
nor UO_548 (O_548,N_2995,N_4585);
nand UO_549 (O_549,N_4054,N_4798);
or UO_550 (O_550,N_2540,N_4889);
or UO_551 (O_551,N_4358,N_3934);
nor UO_552 (O_552,N_4904,N_3716);
or UO_553 (O_553,N_4650,N_3789);
nand UO_554 (O_554,N_2828,N_4079);
and UO_555 (O_555,N_4312,N_2729);
nor UO_556 (O_556,N_4887,N_4282);
nor UO_557 (O_557,N_4610,N_3578);
nand UO_558 (O_558,N_4445,N_3339);
or UO_559 (O_559,N_3529,N_4750);
nor UO_560 (O_560,N_3614,N_3640);
or UO_561 (O_561,N_4967,N_4037);
and UO_562 (O_562,N_2706,N_3245);
and UO_563 (O_563,N_3422,N_3945);
nand UO_564 (O_564,N_2524,N_2880);
nand UO_565 (O_565,N_3624,N_3079);
nand UO_566 (O_566,N_3000,N_2708);
nor UO_567 (O_567,N_3473,N_3426);
nor UO_568 (O_568,N_2791,N_4402);
and UO_569 (O_569,N_4538,N_3931);
and UO_570 (O_570,N_4768,N_2794);
or UO_571 (O_571,N_4916,N_3132);
nor UO_572 (O_572,N_3291,N_4511);
nand UO_573 (O_573,N_2788,N_4126);
nand UO_574 (O_574,N_4897,N_2997);
nand UO_575 (O_575,N_4565,N_3740);
or UO_576 (O_576,N_3046,N_4681);
and UO_577 (O_577,N_2505,N_3384);
nor UO_578 (O_578,N_2802,N_4740);
nor UO_579 (O_579,N_3737,N_4171);
nor UO_580 (O_580,N_2644,N_3405);
and UO_581 (O_581,N_4665,N_2833);
xnor UO_582 (O_582,N_3586,N_3048);
and UO_583 (O_583,N_2878,N_4481);
and UO_584 (O_584,N_4868,N_2969);
and UO_585 (O_585,N_2860,N_4660);
nor UO_586 (O_586,N_2719,N_3201);
nor UO_587 (O_587,N_2600,N_2622);
nor UO_588 (O_588,N_3191,N_4407);
and UO_589 (O_589,N_4927,N_3254);
nand UO_590 (O_590,N_4783,N_2764);
or UO_591 (O_591,N_4633,N_2964);
nor UO_592 (O_592,N_3721,N_3277);
nor UO_593 (O_593,N_3131,N_3871);
and UO_594 (O_594,N_4371,N_2840);
or UO_595 (O_595,N_2542,N_3602);
and UO_596 (O_596,N_3087,N_4459);
or UO_597 (O_597,N_3922,N_4120);
or UO_598 (O_598,N_4769,N_4014);
nand UO_599 (O_599,N_3042,N_4814);
or UO_600 (O_600,N_3352,N_4452);
nand UO_601 (O_601,N_4074,N_2970);
nor UO_602 (O_602,N_2811,N_3773);
or UO_603 (O_603,N_4913,N_4225);
and UO_604 (O_604,N_3415,N_4516);
nor UO_605 (O_605,N_4426,N_4031);
or UO_606 (O_606,N_4050,N_3955);
nand UO_607 (O_607,N_4586,N_4347);
or UO_608 (O_608,N_4438,N_4400);
nand UO_609 (O_609,N_3216,N_2890);
nand UO_610 (O_610,N_2823,N_3943);
and UO_611 (O_611,N_3396,N_3327);
or UO_612 (O_612,N_4258,N_4466);
nor UO_613 (O_613,N_3558,N_3811);
and UO_614 (O_614,N_4930,N_4965);
and UO_615 (O_615,N_4494,N_2538);
and UO_616 (O_616,N_4855,N_2902);
and UO_617 (O_617,N_4963,N_4547);
and UO_618 (O_618,N_3788,N_3082);
nand UO_619 (O_619,N_4376,N_4181);
nor UO_620 (O_620,N_2518,N_3974);
nand UO_621 (O_621,N_4095,N_4739);
or UO_622 (O_622,N_4743,N_4733);
nand UO_623 (O_623,N_2931,N_4643);
nand UO_624 (O_624,N_3942,N_2973);
nand UO_625 (O_625,N_3467,N_3320);
nor UO_626 (O_626,N_3616,N_3982);
nor UO_627 (O_627,N_4023,N_4110);
nor UO_628 (O_628,N_3534,N_3155);
nand UO_629 (O_629,N_4607,N_4559);
nor UO_630 (O_630,N_4211,N_3569);
nand UO_631 (O_631,N_2566,N_3718);
nor UO_632 (O_632,N_2933,N_3496);
and UO_633 (O_633,N_3809,N_4032);
nand UO_634 (O_634,N_2956,N_4990);
or UO_635 (O_635,N_2883,N_3064);
or UO_636 (O_636,N_4486,N_4601);
xnor UO_637 (O_637,N_3839,N_2569);
nand UO_638 (O_638,N_4270,N_3813);
or UO_639 (O_639,N_4149,N_4142);
nand UO_640 (O_640,N_4870,N_4121);
nor UO_641 (O_641,N_3509,N_3581);
xor UO_642 (O_642,N_4202,N_4236);
and UO_643 (O_643,N_2593,N_4644);
or UO_644 (O_644,N_3462,N_2834);
nor UO_645 (O_645,N_3921,N_4807);
and UO_646 (O_646,N_4495,N_4083);
nor UO_647 (O_647,N_4027,N_4544);
nor UO_648 (O_648,N_4238,N_3706);
nor UO_649 (O_649,N_3919,N_3400);
nor UO_650 (O_650,N_4351,N_3980);
nor UO_651 (O_651,N_4234,N_3319);
or UO_652 (O_652,N_4422,N_2892);
and UO_653 (O_653,N_4431,N_3356);
and UO_654 (O_654,N_2741,N_2535);
or UO_655 (O_655,N_3289,N_3844);
or UO_656 (O_656,N_4578,N_4529);
nor UO_657 (O_657,N_3967,N_4443);
and UO_658 (O_658,N_3636,N_2991);
nand UO_659 (O_659,N_2623,N_3033);
or UO_660 (O_660,N_4957,N_4724);
nor UO_661 (O_661,N_2971,N_3492);
nand UO_662 (O_662,N_3165,N_4105);
nand UO_663 (O_663,N_3073,N_4853);
nor UO_664 (O_664,N_3812,N_2756);
or UO_665 (O_665,N_4782,N_4152);
or UO_666 (O_666,N_4695,N_4012);
or UO_667 (O_667,N_3341,N_4620);
nor UO_668 (O_668,N_4629,N_2746);
nand UO_669 (O_669,N_3040,N_4690);
or UO_670 (O_670,N_3539,N_4478);
nor UO_671 (O_671,N_3702,N_4385);
nand UO_672 (O_672,N_3271,N_2651);
and UO_673 (O_673,N_3587,N_3032);
xor UO_674 (O_674,N_3822,N_3739);
nand UO_675 (O_675,N_4675,N_4439);
nand UO_676 (O_676,N_3370,N_2714);
nor UO_677 (O_677,N_3770,N_2626);
nor UO_678 (O_678,N_2710,N_3416);
and UO_679 (O_679,N_4010,N_4109);
and UO_680 (O_680,N_3645,N_4964);
or UO_681 (O_681,N_3725,N_3835);
nor UO_682 (O_682,N_3556,N_4143);
nand UO_683 (O_683,N_4700,N_4614);
nand UO_684 (O_684,N_3178,N_3038);
and UO_685 (O_685,N_4976,N_2705);
nor UO_686 (O_686,N_3528,N_3521);
nor UO_687 (O_687,N_2908,N_4340);
and UO_688 (O_688,N_4420,N_4479);
nand UO_689 (O_689,N_2676,N_3471);
and UO_690 (O_690,N_4185,N_4469);
and UO_691 (O_691,N_2641,N_4885);
nor UO_692 (O_692,N_4209,N_4207);
nor UO_693 (O_693,N_3656,N_2767);
nand UO_694 (O_694,N_3100,N_4277);
nand UO_695 (O_695,N_4689,N_3722);
nor UO_696 (O_696,N_3498,N_4646);
nand UO_697 (O_697,N_3837,N_2695);
or UO_698 (O_698,N_4517,N_2775);
nor UO_699 (O_699,N_3883,N_4276);
and UO_700 (O_700,N_4922,N_4368);
nand UO_701 (O_701,N_4300,N_2939);
and UO_702 (O_702,N_4709,N_4752);
or UO_703 (O_703,N_2875,N_2798);
xor UO_704 (O_704,N_4412,N_2534);
and UO_705 (O_705,N_3126,N_4346);
and UO_706 (O_706,N_4250,N_3299);
nor UO_707 (O_707,N_2634,N_3997);
nor UO_708 (O_708,N_3199,N_3891);
and UO_709 (O_709,N_3819,N_3960);
nor UO_710 (O_710,N_3051,N_4790);
and UO_711 (O_711,N_3247,N_3278);
nor UO_712 (O_712,N_3687,N_2863);
nand UO_713 (O_713,N_3382,N_4645);
and UO_714 (O_714,N_3252,N_3104);
or UO_715 (O_715,N_4793,N_4846);
or UO_716 (O_716,N_2700,N_3489);
and UO_717 (O_717,N_3697,N_4997);
or UO_718 (O_718,N_3745,N_3378);
and UO_719 (O_719,N_3174,N_3069);
nand UO_720 (O_720,N_4377,N_4072);
or UO_721 (O_721,N_4219,N_4735);
nor UO_722 (O_722,N_3371,N_2570);
or UO_723 (O_723,N_2555,N_3411);
nand UO_724 (O_724,N_4107,N_4949);
and UO_725 (O_725,N_2639,N_3388);
nand UO_726 (O_726,N_4167,N_4780);
or UO_727 (O_727,N_3754,N_3179);
and UO_728 (O_728,N_3747,N_4442);
or UO_729 (O_729,N_4119,N_3332);
nand UO_730 (O_730,N_3947,N_4133);
and UO_731 (O_731,N_2906,N_3907);
nor UO_732 (O_732,N_3004,N_3755);
nor UO_733 (O_733,N_3662,N_3729);
or UO_734 (O_734,N_3651,N_2983);
and UO_735 (O_735,N_4531,N_2904);
nand UO_736 (O_736,N_4379,N_2760);
and UO_737 (O_737,N_2561,N_2913);
or UO_738 (O_738,N_3432,N_2663);
nor UO_739 (O_739,N_3806,N_2692);
or UO_740 (O_740,N_3488,N_4115);
nand UO_741 (O_741,N_3904,N_3493);
nand UO_742 (O_742,N_3700,N_2864);
or UO_743 (O_743,N_3932,N_4849);
nand UO_744 (O_744,N_4047,N_3783);
or UO_745 (O_745,N_3985,N_3615);
nor UO_746 (O_746,N_4879,N_4210);
and UO_747 (O_747,N_2992,N_3477);
or UO_748 (O_748,N_3522,N_4177);
nand UO_749 (O_749,N_3407,N_3281);
nand UO_750 (O_750,N_2701,N_2643);
and UO_751 (O_751,N_3094,N_4186);
or UO_752 (O_752,N_4394,N_3535);
nor UO_753 (O_753,N_3006,N_4364);
nand UO_754 (O_754,N_2905,N_3846);
nand UO_755 (O_755,N_2635,N_3642);
nand UO_756 (O_756,N_3487,N_3564);
nor UO_757 (O_757,N_4488,N_2790);
nor UO_758 (O_758,N_4158,N_3941);
nor UO_759 (O_759,N_3961,N_3495);
or UO_760 (O_760,N_4310,N_4619);
or UO_761 (O_761,N_3450,N_4482);
nand UO_762 (O_762,N_4374,N_4939);
and UO_763 (O_763,N_2773,N_2605);
or UO_764 (O_764,N_2871,N_2850);
and UO_765 (O_765,N_4180,N_4847);
and UO_766 (O_766,N_2796,N_3709);
or UO_767 (O_767,N_3446,N_3661);
nor UO_768 (O_768,N_3297,N_4336);
or UO_769 (O_769,N_3666,N_2704);
nand UO_770 (O_770,N_4546,N_2608);
nor UO_771 (O_771,N_3034,N_4324);
nand UO_772 (O_772,N_4141,N_3675);
and UO_773 (O_773,N_4792,N_3920);
nand UO_774 (O_774,N_2504,N_3364);
nand UO_775 (O_775,N_3089,N_2821);
and UO_776 (O_776,N_4064,N_3649);
or UO_777 (O_777,N_3605,N_4691);
or UO_778 (O_778,N_4446,N_3428);
nand UO_779 (O_779,N_4842,N_4381);
or UO_780 (O_780,N_2709,N_2988);
or UO_781 (O_781,N_3540,N_3295);
and UO_782 (O_782,N_4920,N_3482);
xor UO_783 (O_783,N_4532,N_4278);
xor UO_784 (O_784,N_3775,N_2562);
and UO_785 (O_785,N_4281,N_4828);
nor UO_786 (O_786,N_3474,N_3231);
nor UO_787 (O_787,N_3353,N_3013);
nor UO_788 (O_788,N_2715,N_4682);
or UO_789 (O_789,N_2826,N_3372);
or UO_790 (O_790,N_4994,N_3129);
nand UO_791 (O_791,N_4670,N_4592);
and UO_792 (O_792,N_3081,N_3896);
nand UO_793 (O_793,N_3440,N_3635);
and UO_794 (O_794,N_3759,N_3671);
nor UO_795 (O_795,N_4137,N_3766);
nor UO_796 (O_796,N_4430,N_4903);
or UO_797 (O_797,N_4514,N_4656);
or UO_798 (O_798,N_3317,N_3499);
nor UO_799 (O_799,N_2565,N_2670);
or UO_800 (O_800,N_4818,N_4960);
nor UO_801 (O_801,N_4635,N_2680);
nor UO_802 (O_802,N_4008,N_3134);
and UO_803 (O_803,N_2806,N_4317);
nand UO_804 (O_804,N_2580,N_4472);
or UO_805 (O_805,N_3268,N_3712);
or UO_806 (O_806,N_3966,N_3560);
and UO_807 (O_807,N_3894,N_3067);
nand UO_808 (O_808,N_4425,N_2845);
nor UO_809 (O_809,N_4182,N_3047);
and UO_810 (O_810,N_4366,N_2537);
or UO_811 (O_811,N_4268,N_3028);
and UO_812 (O_812,N_4129,N_4533);
nor UO_813 (O_813,N_4067,N_3030);
and UO_814 (O_814,N_3173,N_2940);
nor UO_815 (O_815,N_4940,N_3461);
or UO_816 (O_816,N_4525,N_2571);
and UO_817 (O_817,N_4702,N_2514);
and UO_818 (O_818,N_4615,N_4117);
and UO_819 (O_819,N_3515,N_4352);
or UO_820 (O_820,N_3156,N_3826);
and UO_821 (O_821,N_4751,N_4102);
or UO_822 (O_822,N_3262,N_4062);
and UO_823 (O_823,N_4710,N_4059);
nand UO_824 (O_824,N_2591,N_3629);
nor UO_825 (O_825,N_3220,N_4623);
nor UO_826 (O_826,N_4353,N_3954);
nand UO_827 (O_827,N_4384,N_4314);
and UO_828 (O_828,N_4998,N_4073);
or UO_829 (O_829,N_3823,N_2897);
and UO_830 (O_830,N_2559,N_3197);
or UO_831 (O_831,N_3802,N_3369);
and UO_832 (O_832,N_2761,N_3956);
and UO_833 (O_833,N_3678,N_3176);
nor UO_834 (O_834,N_3085,N_4980);
or UO_835 (O_835,N_2590,N_3223);
nor UO_836 (O_836,N_2529,N_3996);
nand UO_837 (O_837,N_2870,N_4653);
and UO_838 (O_838,N_3274,N_4077);
and UO_839 (O_839,N_2894,N_4819);
nor UO_840 (O_840,N_4205,N_4981);
nor UO_841 (O_841,N_3767,N_4794);
nor UO_842 (O_842,N_3657,N_3989);
or UO_843 (O_843,N_4195,N_3029);
and UO_844 (O_844,N_4404,N_3715);
nor UO_845 (O_845,N_4033,N_4089);
xor UO_846 (O_846,N_4946,N_2573);
or UO_847 (O_847,N_2972,N_3441);
or UO_848 (O_848,N_2872,N_4116);
nand UO_849 (O_849,N_4657,N_3312);
nand UO_850 (O_850,N_3626,N_4825);
and UO_851 (O_851,N_3368,N_3592);
or UO_852 (O_852,N_3902,N_4440);
or UO_853 (O_853,N_3872,N_2926);
nor UO_854 (O_854,N_4130,N_3011);
nand UO_855 (O_855,N_3494,N_4246);
or UO_856 (O_856,N_3714,N_4820);
and UO_857 (O_857,N_4784,N_3175);
and UO_858 (O_858,N_2903,N_4396);
or UO_859 (O_859,N_3113,N_4315);
or UO_860 (O_860,N_4198,N_3916);
and UO_861 (O_861,N_4052,N_3465);
xnor UO_862 (O_862,N_3209,N_4470);
and UO_863 (O_863,N_4415,N_4919);
nor UO_864 (O_864,N_3043,N_2547);
nand UO_865 (O_865,N_2807,N_4956);
nand UO_866 (O_866,N_2928,N_4550);
nor UO_867 (O_867,N_3304,N_4383);
or UO_868 (O_868,N_4838,N_3154);
and UO_869 (O_869,N_4804,N_3442);
or UO_870 (O_870,N_3360,N_2678);
or UO_871 (O_871,N_4839,N_3923);
nor UO_872 (O_872,N_2677,N_3161);
and UO_873 (O_873,N_4071,N_2998);
nor UO_874 (O_874,N_3536,N_4433);
nand UO_875 (O_875,N_4512,N_3394);
or UO_876 (O_876,N_3971,N_3470);
or UO_877 (O_877,N_3772,N_4432);
and UO_878 (O_878,N_4279,N_4123);
xnor UO_879 (O_879,N_2942,N_4667);
and UO_880 (O_880,N_4542,N_3463);
nor UO_881 (O_881,N_4040,N_4654);
or UO_882 (O_882,N_2582,N_3672);
or UO_883 (O_883,N_4639,N_4093);
xor UO_884 (O_884,N_4749,N_4781);
and UO_885 (O_885,N_3915,N_3318);
or UO_886 (O_886,N_3734,N_3417);
nand UO_887 (O_887,N_3376,N_4954);
and UO_888 (O_888,N_4866,N_3897);
and UO_889 (O_889,N_4419,N_3832);
or UO_890 (O_890,N_3464,N_3553);
and UO_891 (O_891,N_3233,N_2895);
or UO_892 (O_892,N_3582,N_4038);
or UO_893 (O_893,N_4652,N_2750);
and UO_894 (O_894,N_2699,N_3552);
and UO_895 (O_895,N_3023,N_3738);
and UO_896 (O_896,N_4013,N_2653);
nor UO_897 (O_897,N_3251,N_2810);
and UO_898 (O_898,N_4628,N_3869);
nand UO_899 (O_899,N_3753,N_2674);
or UO_900 (O_900,N_2684,N_3938);
nand UO_901 (O_901,N_3351,N_3713);
nand UO_902 (O_902,N_4144,N_3455);
nand UO_903 (O_903,N_2519,N_2929);
and UO_904 (O_904,N_3138,N_3905);
nor UO_905 (O_905,N_4163,N_4208);
nor UO_906 (O_906,N_4507,N_2625);
and UO_907 (O_907,N_3917,N_2629);
nor UO_908 (O_908,N_3866,N_2739);
xor UO_909 (O_909,N_4128,N_2533);
nand UO_910 (O_910,N_3604,N_3401);
nand UO_911 (O_911,N_3010,N_4579);
nand UO_912 (O_912,N_3603,N_4666);
and UO_913 (O_913,N_3746,N_2531);
nor UO_914 (O_914,N_2627,N_4996);
or UO_915 (O_915,N_4280,N_3910);
nor UO_916 (O_916,N_3571,N_3935);
nand UO_917 (O_917,N_4999,N_4851);
and UO_918 (O_918,N_3692,N_4139);
or UO_919 (O_919,N_4237,N_4474);
or UO_920 (O_920,N_4910,N_4456);
xnor UO_921 (O_921,N_4344,N_3036);
nand UO_922 (O_922,N_2694,N_4018);
nor UO_923 (O_923,N_3912,N_3782);
and UO_924 (O_924,N_4160,N_3124);
or UO_925 (O_925,N_4041,N_3719);
or UO_926 (O_926,N_2659,N_4717);
nand UO_927 (O_927,N_3899,N_2769);
nor UO_928 (O_928,N_4603,N_4212);
nor UO_929 (O_929,N_4006,N_2735);
nor UO_930 (O_930,N_3760,N_3444);
nor UO_931 (O_931,N_3593,N_4391);
or UO_932 (O_932,N_2738,N_4557);
nor UO_933 (O_933,N_4294,N_3860);
and UO_934 (O_934,N_2812,N_4359);
nor UO_935 (O_935,N_4823,N_4566);
nand UO_936 (O_936,N_4705,N_4408);
or UO_937 (O_937,N_4543,N_4251);
and UO_938 (O_938,N_4706,N_4860);
and UO_939 (O_939,N_4704,N_3014);
nor UO_940 (O_940,N_3781,N_4173);
nor UO_941 (O_941,N_4231,N_3554);
nor UO_942 (O_942,N_3017,N_3395);
and UO_943 (O_943,N_2557,N_3768);
and UO_944 (O_944,N_4993,N_2501);
nand UO_945 (O_945,N_2876,N_4641);
or UO_946 (O_946,N_2900,N_4918);
nor UO_947 (O_947,N_3648,N_4975);
nor UO_948 (O_948,N_4081,N_3856);
nor UO_949 (O_949,N_3850,N_4009);
or UO_950 (O_950,N_3573,N_3828);
nor UO_951 (O_951,N_2707,N_4357);
and UO_952 (O_952,N_4627,N_2770);
nor UO_953 (O_953,N_3335,N_3752);
nor UO_954 (O_954,N_3950,N_2879);
nand UO_955 (O_955,N_4679,N_2838);
nand UO_956 (O_956,N_4007,N_4002);
or UO_957 (O_957,N_2583,N_4369);
and UO_958 (O_958,N_3668,N_3726);
nand UO_959 (O_959,N_4338,N_3701);
or UO_960 (O_960,N_2737,N_2743);
nor UO_961 (O_961,N_3227,N_3308);
and UO_962 (O_962,N_4971,N_3992);
and UO_963 (O_963,N_4151,N_4878);
and UO_964 (O_964,N_3049,N_3164);
or UO_965 (O_965,N_3674,N_4045);
xnor UO_966 (O_966,N_3092,N_3707);
nor UO_967 (O_967,N_2948,N_2606);
or UO_968 (O_968,N_4630,N_4613);
nand UO_969 (O_969,N_4240,N_2974);
nand UO_970 (O_970,N_4882,N_4655);
or UO_971 (O_971,N_4862,N_3538);
or UO_972 (O_972,N_4886,N_3250);
or UO_973 (O_973,N_2711,N_2717);
nor UO_974 (O_974,N_4606,N_3873);
or UO_975 (O_975,N_3381,N_2718);
and UO_976 (O_976,N_2712,N_3677);
and UO_977 (O_977,N_3435,N_3566);
nor UO_978 (O_978,N_3831,N_4938);
and UO_979 (O_979,N_2980,N_4348);
or UO_980 (O_980,N_4741,N_2795);
or UO_981 (O_981,N_3002,N_3096);
nand UO_982 (O_982,N_2754,N_4162);
or UO_983 (O_983,N_4053,N_3066);
nand UO_984 (O_984,N_4966,N_4555);
and UO_985 (O_985,N_3204,N_4464);
nand UO_986 (O_986,N_3083,N_3323);
nand UO_987 (O_987,N_4411,N_2652);
nor UO_988 (O_988,N_4104,N_2886);
nand UO_989 (O_989,N_3213,N_3514);
nor UO_990 (O_990,N_3940,N_4551);
xnor UO_991 (O_991,N_2999,N_3217);
or UO_992 (O_992,N_4485,N_4502);
nand UO_993 (O_993,N_3302,N_2616);
or UO_994 (O_994,N_2586,N_2815);
or UO_995 (O_995,N_4912,N_3230);
nand UO_996 (O_996,N_2861,N_3280);
nor UO_997 (O_997,N_4854,N_3512);
and UO_998 (O_998,N_4437,N_3848);
nand UO_999 (O_999,N_2527,N_4659);
endmodule