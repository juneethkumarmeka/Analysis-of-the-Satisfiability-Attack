module basic_2000_20000_2500_50_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xnor U0 (N_0,In_280,In_685);
nand U1 (N_1,In_897,In_1582);
nor U2 (N_2,In_1564,In_1643);
and U3 (N_3,In_533,In_484);
xor U4 (N_4,In_935,In_1362);
xnor U5 (N_5,In_1885,In_1878);
xor U6 (N_6,In_844,In_1673);
nor U7 (N_7,In_1559,In_63);
nand U8 (N_8,In_237,In_173);
nand U9 (N_9,In_1117,In_1932);
and U10 (N_10,In_116,In_1158);
nor U11 (N_11,In_1266,In_271);
xnor U12 (N_12,In_241,In_718);
and U13 (N_13,In_35,In_664);
nor U14 (N_14,In_1889,In_677);
or U15 (N_15,In_1585,In_1856);
and U16 (N_16,In_1935,In_1096);
xor U17 (N_17,In_44,In_1896);
or U18 (N_18,In_1906,In_146);
and U19 (N_19,In_700,In_1327);
nor U20 (N_20,In_185,In_1696);
and U21 (N_21,In_1799,In_776);
xor U22 (N_22,In_1299,In_164);
nand U23 (N_23,In_1404,In_1275);
and U24 (N_24,In_492,In_104);
nor U25 (N_25,In_495,In_569);
or U26 (N_26,In_707,In_435);
and U27 (N_27,In_628,In_208);
nor U28 (N_28,In_1430,In_141);
nor U29 (N_29,In_189,In_1229);
nand U30 (N_30,In_1520,In_1944);
nand U31 (N_31,In_1527,In_1899);
or U32 (N_32,In_1315,In_1674);
xnor U33 (N_33,In_1432,In_218);
nor U34 (N_34,In_420,In_801);
nor U35 (N_35,In_1057,In_295);
and U36 (N_36,In_265,In_1011);
or U37 (N_37,In_748,In_1152);
xor U38 (N_38,In_1713,In_1540);
xor U39 (N_39,In_268,In_1413);
and U40 (N_40,In_105,In_1610);
xor U41 (N_41,In_1496,In_1816);
xnor U42 (N_42,In_1340,In_927);
nand U43 (N_43,In_395,In_1341);
and U44 (N_44,In_1176,In_993);
xnor U45 (N_45,In_696,In_1184);
xnor U46 (N_46,In_527,In_1021);
nor U47 (N_47,In_544,In_1511);
xor U48 (N_48,In_1759,In_1730);
xor U49 (N_49,In_918,In_647);
nor U50 (N_50,In_1534,In_96);
nor U51 (N_51,In_1870,In_1181);
or U52 (N_52,In_670,In_60);
xor U53 (N_53,In_158,In_519);
xnor U54 (N_54,In_1571,In_656);
or U55 (N_55,In_1213,In_543);
xor U56 (N_56,In_1707,In_509);
nand U57 (N_57,In_247,In_631);
xor U58 (N_58,In_1918,In_1037);
nor U59 (N_59,In_402,In_1027);
and U60 (N_60,In_1798,In_950);
xor U61 (N_61,In_1784,In_600);
nor U62 (N_62,In_375,In_83);
xor U63 (N_63,In_1062,In_449);
nand U64 (N_64,In_709,In_592);
and U65 (N_65,In_756,In_1846);
and U66 (N_66,In_1562,In_1045);
nand U67 (N_67,In_360,In_1568);
and U68 (N_68,In_283,In_152);
nor U69 (N_69,In_223,In_1371);
and U70 (N_70,In_1143,In_1952);
xor U71 (N_71,In_673,In_1917);
nand U72 (N_72,In_318,In_1170);
and U73 (N_73,In_728,In_1701);
and U74 (N_74,In_1475,In_425);
and U75 (N_75,In_272,In_1531);
xor U76 (N_76,In_573,In_1063);
and U77 (N_77,In_1761,In_798);
nand U78 (N_78,In_1864,In_1958);
xor U79 (N_79,In_1907,In_303);
nor U80 (N_80,In_1159,In_846);
nor U81 (N_81,In_263,In_25);
xor U82 (N_82,In_292,In_373);
xnor U83 (N_83,In_1345,In_29);
nor U84 (N_84,In_1055,In_995);
and U85 (N_85,In_1734,In_1572);
or U86 (N_86,In_1904,In_1565);
nor U87 (N_87,In_1291,In_830);
and U88 (N_88,In_1853,In_741);
and U89 (N_89,In_396,In_1621);
xor U90 (N_90,In_558,In_1965);
and U91 (N_91,In_1136,In_1834);
and U92 (N_92,In_667,In_912);
xnor U93 (N_93,In_714,In_204);
or U94 (N_94,In_891,In_645);
nor U95 (N_95,In_1187,In_31);
nand U96 (N_96,In_1987,In_1156);
and U97 (N_97,In_1522,In_1548);
xor U98 (N_98,In_1635,In_1149);
nand U99 (N_99,In_190,In_1874);
nor U100 (N_100,In_749,In_1274);
or U101 (N_101,In_352,In_1589);
xnor U102 (N_102,In_1990,In_64);
or U103 (N_103,In_924,In_1733);
nand U104 (N_104,In_1429,In_938);
nor U105 (N_105,In_398,In_1480);
xnor U106 (N_106,In_1796,In_1352);
and U107 (N_107,In_90,In_553);
xnor U108 (N_108,In_1091,In_314);
or U109 (N_109,In_424,In_1975);
xor U110 (N_110,In_338,In_1479);
nor U111 (N_111,In_1431,In_674);
xnor U112 (N_112,In_811,In_883);
xor U113 (N_113,In_982,In_447);
xor U114 (N_114,In_925,In_605);
nor U115 (N_115,In_1766,In_1611);
or U116 (N_116,In_1836,In_1819);
xnor U117 (N_117,In_973,In_630);
nor U118 (N_118,In_1772,In_1344);
and U119 (N_119,In_277,In_1558);
or U120 (N_120,In_648,In_1203);
nand U121 (N_121,In_832,In_1214);
nor U122 (N_122,In_652,In_942);
or U123 (N_123,In_808,In_699);
or U124 (N_124,In_561,In_1485);
or U125 (N_125,In_1133,In_342);
xnor U126 (N_126,In_1793,In_1873);
or U127 (N_127,In_1619,In_1788);
nand U128 (N_128,In_366,In_165);
nand U129 (N_129,In_1258,In_568);
nor U130 (N_130,In_675,In_1460);
nor U131 (N_131,In_1105,In_1389);
and U132 (N_132,In_1415,In_646);
nand U133 (N_133,In_517,In_438);
nor U134 (N_134,In_1146,In_299);
nor U135 (N_135,In_1180,In_483);
xnor U136 (N_136,In_336,In_30);
nand U137 (N_137,In_1025,In_695);
and U138 (N_138,In_1546,In_802);
or U139 (N_139,In_1708,In_1338);
xor U140 (N_140,In_1403,In_1435);
or U141 (N_141,In_1523,In_287);
xor U142 (N_142,In_74,In_371);
or U143 (N_143,In_1791,In_273);
xnor U144 (N_144,In_1841,In_760);
xnor U145 (N_145,In_1882,In_1848);
and U146 (N_146,In_916,In_1252);
nand U147 (N_147,In_477,In_637);
nand U148 (N_148,In_551,In_1224);
xnor U149 (N_149,In_1646,In_1215);
nand U150 (N_150,In_1,In_822);
and U151 (N_151,In_722,In_160);
xor U152 (N_152,In_1456,In_242);
nand U153 (N_153,In_428,In_693);
and U154 (N_154,In_1519,In_1669);
nand U155 (N_155,In_493,In_1964);
or U156 (N_156,In_219,In_379);
nand U157 (N_157,In_1009,In_764);
nand U158 (N_158,In_170,In_1137);
xnor U159 (N_159,In_698,In_347);
or U160 (N_160,In_469,In_506);
nand U161 (N_161,In_1373,In_1951);
and U162 (N_162,In_15,In_412);
and U163 (N_163,In_1623,In_1634);
nand U164 (N_164,In_27,In_1428);
nor U165 (N_165,In_729,In_434);
xnor U166 (N_166,In_708,In_252);
or U167 (N_167,In_1075,In_818);
nor U168 (N_168,In_894,In_1116);
nor U169 (N_169,In_1406,In_977);
or U170 (N_170,In_1844,In_372);
and U171 (N_171,In_87,In_657);
and U172 (N_172,In_202,In_1263);
or U173 (N_173,In_1489,In_878);
or U174 (N_174,In_723,In_747);
nand U175 (N_175,In_1294,In_28);
and U176 (N_176,In_494,In_339);
xnor U177 (N_177,In_1241,In_381);
nand U178 (N_178,In_1207,In_1586);
or U179 (N_179,In_797,In_468);
nor U180 (N_180,In_632,In_1620);
or U181 (N_181,In_1378,In_1833);
xor U182 (N_182,In_1350,In_266);
xor U183 (N_183,In_1440,In_1061);
and U184 (N_184,In_1810,In_1545);
xor U185 (N_185,In_905,In_796);
xnor U186 (N_186,In_1386,In_1970);
nand U187 (N_187,In_515,In_1382);
xnor U188 (N_188,In_1065,In_1400);
or U189 (N_189,In_789,In_1992);
xnor U190 (N_190,In_1098,In_205);
or U191 (N_191,In_18,In_1962);
or U192 (N_192,In_1588,In_1043);
nand U193 (N_193,In_1238,In_979);
or U194 (N_194,In_1020,In_886);
and U195 (N_195,In_1677,In_1573);
xnor U196 (N_196,In_1078,In_458);
xor U197 (N_197,In_1265,In_124);
nand U198 (N_198,In_1804,In_545);
or U199 (N_199,In_731,In_279);
or U200 (N_200,In_36,In_680);
nor U201 (N_201,In_989,In_1938);
nor U202 (N_202,In_1821,In_1984);
and U203 (N_203,In_1245,In_431);
or U204 (N_204,In_650,In_301);
or U205 (N_205,In_1211,In_1459);
and U206 (N_206,In_1795,In_869);
and U207 (N_207,In_526,In_496);
or U208 (N_208,In_604,In_1463);
nor U209 (N_209,In_1337,In_1601);
xnor U210 (N_210,In_1943,In_1501);
nand U211 (N_211,In_996,In_625);
and U212 (N_212,In_964,In_121);
xnor U213 (N_213,In_1763,In_1441);
nand U214 (N_214,In_1495,In_365);
nand U215 (N_215,In_407,In_1416);
nor U216 (N_216,In_1609,In_459);
nor U217 (N_217,In_294,In_445);
nor U218 (N_218,In_1309,In_531);
and U219 (N_219,In_1687,In_833);
xor U220 (N_220,In_1838,In_1196);
nor U221 (N_221,In_1602,In_816);
and U222 (N_222,In_1250,In_1902);
and U223 (N_223,In_285,In_594);
xnor U224 (N_224,In_1201,In_195);
xnor U225 (N_225,In_1202,In_1538);
or U226 (N_226,In_1040,In_1805);
nor U227 (N_227,In_455,In_727);
xnor U228 (N_228,In_951,In_1410);
xnor U229 (N_229,In_1161,In_1825);
nand U230 (N_230,In_997,In_1458);
nor U231 (N_231,In_1753,In_70);
nor U232 (N_232,In_175,In_1569);
and U233 (N_233,In_1319,In_810);
nand U234 (N_234,In_1774,In_1281);
and U235 (N_235,In_1222,In_649);
nor U236 (N_236,In_1000,In_181);
xor U237 (N_237,In_1947,In_144);
nand U238 (N_238,In_1100,In_1705);
or U239 (N_239,In_1069,In_941);
or U240 (N_240,In_1018,In_274);
nand U241 (N_241,In_1731,In_1629);
xor U242 (N_242,In_1234,In_623);
and U243 (N_243,In_1038,In_1498);
or U244 (N_244,In_538,In_1064);
or U245 (N_245,In_1995,In_88);
nand U246 (N_246,In_1076,In_1505);
or U247 (N_247,In_726,In_1004);
nor U248 (N_248,In_143,In_1871);
nand U249 (N_249,In_1676,In_1304);
nand U250 (N_250,In_614,In_643);
or U251 (N_251,In_585,In_635);
or U252 (N_252,In_940,In_862);
or U253 (N_253,In_1886,In_991);
or U254 (N_254,In_762,In_583);
or U255 (N_255,In_203,In_159);
nor U256 (N_256,In_1636,In_467);
and U257 (N_257,In_453,In_1797);
nand U258 (N_258,In_1311,In_199);
nand U259 (N_259,In_1058,In_446);
xnor U260 (N_260,In_970,In_1127);
nand U261 (N_261,In_834,In_1271);
nand U262 (N_262,In_885,In_1112);
nand U263 (N_263,In_791,In_1614);
and U264 (N_264,In_489,In_82);
nand U265 (N_265,In_611,In_895);
nand U266 (N_266,In_906,In_1518);
xnor U267 (N_267,In_1849,In_1269);
nand U268 (N_268,In_860,In_1924);
nand U269 (N_269,In_1854,In_1684);
or U270 (N_270,In_1808,In_1320);
nand U271 (N_271,In_586,In_1926);
or U272 (N_272,In_873,In_1472);
and U273 (N_273,In_1749,In_1420);
and U274 (N_274,In_1289,In_1783);
nand U275 (N_275,In_1240,In_1380);
or U276 (N_276,In_331,In_236);
and U277 (N_277,In_1444,In_220);
and U278 (N_278,In_817,In_1008);
or U279 (N_279,In_1663,In_972);
or U280 (N_280,In_570,In_532);
nor U281 (N_281,In_397,In_1032);
nand U282 (N_282,In_884,In_409);
nor U283 (N_283,In_734,In_1462);
xnor U284 (N_284,In_787,In_478);
nor U285 (N_285,In_1433,In_300);
and U286 (N_286,In_686,In_1583);
nor U287 (N_287,In_575,In_1115);
and U288 (N_288,In_196,In_535);
xor U289 (N_289,In_1276,In_1244);
xor U290 (N_290,In_1054,In_546);
nor U291 (N_291,In_974,In_888);
nand U292 (N_292,In_472,In_1794);
nor U293 (N_293,In_779,In_1557);
xnor U294 (N_294,In_618,In_1171);
or U295 (N_295,In_1072,In_858);
xor U296 (N_296,In_240,In_1385);
xor U297 (N_297,In_689,In_394);
nor U298 (N_298,In_333,In_1515);
nor U299 (N_299,In_113,In_1724);
or U300 (N_300,In_1042,In_1991);
nor U301 (N_301,In_54,In_601);
or U302 (N_302,In_1357,In_317);
xnor U303 (N_303,In_1101,In_1030);
and U304 (N_304,In_1616,In_1827);
nor U305 (N_305,In_880,In_1603);
and U306 (N_306,In_10,In_1499);
xnor U307 (N_307,In_1384,In_307);
nand U308 (N_308,In_1887,In_1165);
nor U309 (N_309,In_403,In_244);
nand U310 (N_310,In_1913,In_430);
nor U311 (N_311,In_1561,In_38);
nor U312 (N_312,In_1931,In_1046);
xnor U313 (N_313,In_23,In_1948);
xor U314 (N_314,In_588,In_139);
xor U315 (N_315,In_854,In_59);
nand U316 (N_316,In_1418,In_933);
or U317 (N_317,In_1608,In_752);
nand U318 (N_318,In_740,In_1656);
nor U319 (N_319,In_476,In_1217);
or U320 (N_320,In_226,In_1706);
or U321 (N_321,In_1567,In_1323);
or U322 (N_322,In_1067,In_922);
or U323 (N_323,In_1082,In_1493);
and U324 (N_324,In_1086,In_177);
nand U325 (N_325,In_1039,In_1927);
nand U326 (N_326,In_217,In_634);
nand U327 (N_327,In_732,In_1197);
or U328 (N_328,In_1439,In_820);
or U329 (N_329,In_1711,In_1167);
nor U330 (N_330,In_421,In_1826);
xnor U331 (N_331,In_1925,In_960);
nand U332 (N_332,In_1405,In_259);
nor U333 (N_333,In_461,In_1736);
and U334 (N_334,In_201,In_427);
xor U335 (N_335,In_161,In_1090);
xor U336 (N_336,In_41,In_809);
or U337 (N_337,In_1070,In_1517);
xnor U338 (N_338,In_357,In_1551);
nor U339 (N_339,In_474,In_145);
and U340 (N_340,In_1452,In_275);
nand U341 (N_341,In_813,In_463);
nand U342 (N_342,In_669,In_914);
and U343 (N_343,In_1138,In_1750);
xor U344 (N_344,In_21,In_559);
nor U345 (N_345,In_865,In_1453);
and U346 (N_346,In_1273,In_311);
nor U347 (N_347,In_1071,In_815);
and U348 (N_348,In_929,In_313);
nand U349 (N_349,In_1892,In_1672);
nor U350 (N_350,In_824,In_1680);
xor U351 (N_351,In_861,In_382);
or U352 (N_352,In_1769,In_1381);
nand U353 (N_353,In_122,In_174);
nand U354 (N_354,In_856,In_1823);
nand U355 (N_355,In_857,In_1866);
or U356 (N_356,In_654,In_961);
or U357 (N_357,In_665,In_1477);
or U358 (N_358,In_1339,In_1175);
xor U359 (N_359,In_939,In_1120);
nand U360 (N_360,In_839,In_84);
or U361 (N_361,In_99,In_253);
or U362 (N_362,In_418,In_1879);
or U363 (N_363,In_1321,In_522);
and U364 (N_364,In_234,In_930);
nand U365 (N_365,In_1110,In_1504);
nor U366 (N_366,In_556,In_1660);
or U367 (N_367,In_1863,In_1461);
nor U368 (N_368,In_1876,In_389);
and U369 (N_369,In_1556,In_260);
nand U370 (N_370,In_1425,In_1737);
xnor U371 (N_371,In_786,In_98);
nor U372 (N_372,In_1929,In_1939);
xnor U373 (N_373,In_1328,In_1850);
nor U374 (N_374,In_1179,In_1638);
xnor U375 (N_375,In_1114,In_1348);
nor U376 (N_376,In_772,In_1738);
nand U377 (N_377,In_1858,In_1121);
or U378 (N_378,In_1284,In_1664);
xnor U379 (N_379,In_1637,In_1113);
or U380 (N_380,In_1861,In_1243);
nand U381 (N_381,In_516,In_1963);
xor U382 (N_382,In_42,In_1314);
nor U383 (N_383,In_1423,In_86);
and U384 (N_384,In_376,In_1683);
nor U385 (N_385,In_1366,In_1968);
nand U386 (N_386,In_539,In_1950);
nor U387 (N_387,In_1503,In_1698);
or U388 (N_388,In_140,In_1387);
xor U389 (N_389,In_480,In_1093);
nand U390 (N_390,In_123,In_1514);
xor U391 (N_391,In_1921,In_636);
nand U392 (N_392,In_902,In_485);
nand U393 (N_393,In_676,In_444);
and U394 (N_394,In_1194,In_1627);
xor U395 (N_395,In_1312,In_1442);
nor U396 (N_396,In_1059,In_1200);
xor U397 (N_397,In_549,In_1956);
or U398 (N_398,In_1754,In_1017);
or U399 (N_399,In_358,In_1164);
nand U400 (N_400,In_1144,In_37);
and U401 (N_401,In_871,In_481);
nor U402 (N_402,In_126,In_1288);
and U403 (N_403,In_1457,N_39);
or U404 (N_404,In_1219,In_1237);
and U405 (N_405,In_356,N_122);
nand U406 (N_406,In_131,In_1507);
or U407 (N_407,In_1625,In_1332);
and U408 (N_408,In_1331,In_804);
nand U409 (N_409,In_1729,N_164);
xnor U410 (N_410,In_994,In_1310);
or U411 (N_411,In_80,In_651);
nand U412 (N_412,In_191,In_829);
xor U413 (N_413,In_1712,N_367);
nor U414 (N_414,In_655,In_790);
or U415 (N_415,In_738,In_937);
or U416 (N_416,In_1450,In_163);
nand U417 (N_417,In_1407,In_1445);
and U418 (N_418,In_507,N_398);
xnor U419 (N_419,In_291,N_108);
xor U420 (N_420,In_1985,In_1957);
nand U421 (N_421,In_1139,In_875);
xor U422 (N_422,In_1688,In_1449);
or U423 (N_423,In_1399,In_510);
or U424 (N_424,N_248,N_273);
nor U425 (N_425,In_1806,In_1659);
xnor U426 (N_426,In_572,In_1437);
nor U427 (N_427,In_823,N_134);
or U428 (N_428,In_1376,In_715);
and U429 (N_429,N_81,In_1230);
nor U430 (N_430,In_442,In_1126);
nor U431 (N_431,In_1010,In_932);
and U432 (N_432,In_753,In_1108);
xor U433 (N_433,In_923,In_702);
nand U434 (N_434,In_255,In_1003);
or U435 (N_435,In_209,In_992);
nor U436 (N_436,In_20,In_1317);
or U437 (N_437,In_1154,In_475);
xor U438 (N_438,In_754,N_186);
xor U439 (N_439,In_392,N_175);
or U440 (N_440,In_337,In_155);
nor U441 (N_441,In_1893,N_365);
xor U442 (N_442,In_106,In_867);
nand U443 (N_443,N_98,In_390);
nor U444 (N_444,In_1700,In_1618);
or U445 (N_445,In_115,In_1443);
xnor U446 (N_446,In_1166,In_229);
nor U447 (N_447,In_264,In_745);
or U448 (N_448,N_204,In_943);
nand U449 (N_449,N_358,N_72);
nor U450 (N_450,N_174,N_369);
nand U451 (N_451,In_102,N_173);
nor U452 (N_452,In_641,N_243);
or U453 (N_453,In_755,In_1426);
nor U454 (N_454,In_1131,N_263);
nor U455 (N_455,In_843,In_1901);
nor U456 (N_456,In_1526,N_184);
nor U457 (N_457,In_1168,In_518);
and U458 (N_458,In_720,In_1102);
and U459 (N_459,In_8,In_50);
or U460 (N_460,In_1279,In_1820);
nand U461 (N_461,In_212,In_1591);
xnor U462 (N_462,In_842,N_396);
nor U463 (N_463,In_1360,In_1122);
nand U464 (N_464,In_1831,N_231);
nor U465 (N_465,In_1868,N_85);
and U466 (N_466,In_486,N_199);
or U467 (N_467,In_1624,In_946);
nor U468 (N_468,In_739,In_1414);
nor U469 (N_469,N_383,In_757);
xnor U470 (N_470,In_222,In_687);
nand U471 (N_471,N_202,N_285);
nand U472 (N_472,In_1272,N_114);
and U473 (N_473,In_1966,In_249);
or U474 (N_474,N_321,In_758);
nor U475 (N_475,In_111,N_86);
and U476 (N_476,In_777,N_247);
or U477 (N_477,In_450,N_298);
xnor U478 (N_478,In_821,In_348);
nor U479 (N_479,In_794,N_38);
or U480 (N_480,In_1728,In_855);
or U481 (N_481,N_178,N_107);
nand U482 (N_482,In_1257,In_1862);
nand U483 (N_483,N_337,In_286);
and U484 (N_484,In_1855,N_3);
nor U485 (N_485,In_184,N_141);
and U486 (N_486,In_58,N_293);
and U487 (N_487,In_419,In_1613);
xor U488 (N_488,In_206,In_1254);
nor U489 (N_489,In_975,In_1349);
or U490 (N_490,In_1290,N_262);
nor U491 (N_491,In_93,In_1095);
and U492 (N_492,N_308,In_1996);
and U493 (N_493,In_582,In_369);
or U494 (N_494,In_1424,In_591);
xnor U495 (N_495,In_759,In_1506);
and U496 (N_496,N_305,In_1394);
nand U497 (N_497,N_320,In_1811);
and U498 (N_498,N_6,In_1787);
or U499 (N_499,In_1605,N_348);
or U500 (N_500,N_209,In_1492);
and U501 (N_501,N_58,In_136);
nand U502 (N_502,In_1287,N_9);
xnor U503 (N_503,N_34,In_1693);
or U504 (N_504,In_387,In_848);
nand U505 (N_505,In_125,In_840);
nand U506 (N_506,In_383,In_1775);
xnor U507 (N_507,In_330,In_557);
or U508 (N_508,N_311,N_121);
nor U509 (N_509,In_1723,In_319);
nor U510 (N_510,N_257,In_43);
nand U511 (N_511,In_1411,In_34);
or U512 (N_512,In_130,In_1860);
nand U513 (N_513,N_316,In_1537);
nand U514 (N_514,In_1869,N_233);
xor U515 (N_515,In_114,In_1883);
nand U516 (N_516,In_595,In_1575);
xor U517 (N_517,N_310,In_440);
and U518 (N_518,In_1802,In_1818);
nand U519 (N_519,N_368,In_230);
or U520 (N_520,N_20,In_679);
and U521 (N_521,N_319,In_751);
and U522 (N_522,In_49,In_134);
nand U523 (N_523,In_1466,N_301);
or U524 (N_524,In_1598,In_788);
and U525 (N_525,In_1081,In_1747);
xnor U526 (N_526,In_1278,N_128);
nor U527 (N_527,In_1928,In_1976);
xor U528 (N_528,N_104,N_258);
nor U529 (N_529,N_132,N_42);
or U530 (N_530,In_503,N_222);
nand U531 (N_531,N_144,In_706);
nand U532 (N_532,N_296,In_1812);
or U533 (N_533,In_1270,In_828);
xor U534 (N_534,N_28,N_264);
xnor U535 (N_535,In_62,In_296);
or U536 (N_536,In_1584,In_1470);
or U537 (N_537,N_250,N_357);
and U538 (N_538,In_148,N_68);
nand U539 (N_539,In_990,In_520);
or U540 (N_540,In_1967,In_1313);
and U541 (N_541,In_1719,In_312);
xnor U542 (N_542,N_295,In_959);
xor U543 (N_543,In_1830,In_1118);
or U544 (N_544,In_448,N_56);
and U545 (N_545,In_683,In_1817);
nor U546 (N_546,N_194,In_849);
and U547 (N_547,In_1715,In_660);
nand U548 (N_548,N_143,In_1471);
or U549 (N_549,In_4,N_90);
or U550 (N_550,In_52,In_361);
nand U551 (N_551,In_1617,N_335);
xnor U552 (N_552,In_1727,In_1702);
xor U553 (N_553,In_1084,In_1367);
nor U554 (N_554,N_251,In_1186);
xor U555 (N_555,In_1773,In_1026);
xor U556 (N_556,N_7,N_78);
xor U557 (N_557,In_1232,In_1912);
or U558 (N_558,In_1668,In_694);
nand U559 (N_559,N_192,In_900);
nor U560 (N_560,In_1353,N_252);
or U561 (N_561,In_380,In_1395);
nor U562 (N_562,In_1735,In_845);
and U563 (N_563,N_2,In_926);
and U564 (N_564,N_29,In_1785);
nand U565 (N_565,N_271,In_917);
or U566 (N_566,In_7,In_1342);
nor U567 (N_567,In_24,In_1626);
nor U568 (N_568,In_769,In_17);
and U569 (N_569,In_351,In_1710);
or U570 (N_570,In_228,In_309);
nor U571 (N_571,In_795,In_1052);
xnor U572 (N_572,In_626,In_602);
and U573 (N_573,In_367,In_1125);
and U574 (N_574,In_498,In_919);
or U575 (N_575,In_998,In_1206);
xor U576 (N_576,In_92,In_550);
nand U577 (N_577,N_161,In_290);
nor U578 (N_578,In_1704,N_373);
nor U579 (N_579,In_451,N_347);
and U580 (N_580,In_956,In_1231);
and U581 (N_581,N_281,N_99);
xor U582 (N_582,In_1647,In_441);
xnor U583 (N_583,In_981,In_1752);
nand U584 (N_584,In_1322,In_1652);
nand U585 (N_585,In_501,In_1590);
nor U586 (N_586,In_1587,In_1541);
nor U587 (N_587,N_155,N_137);
nand U588 (N_588,In_644,In_213);
nor U589 (N_589,In_1822,In_1936);
or U590 (N_590,In_1694,N_236);
xnor U591 (N_591,In_1800,N_21);
nor U592 (N_592,In_653,In_1267);
xnor U593 (N_593,In_1083,In_250);
nand U594 (N_594,In_415,In_1890);
nor U595 (N_595,In_1756,In_335);
nor U596 (N_596,In_1661,In_710);
or U597 (N_597,In_774,In_370);
nand U598 (N_598,In_955,In_671);
nor U599 (N_599,In_103,In_1739);
or U600 (N_600,In_127,In_1370);
nor U601 (N_601,In_1358,N_185);
nand U602 (N_602,In_1140,In_837);
nand U603 (N_603,In_1767,In_1497);
and U604 (N_604,In_499,In_584);
xnor U605 (N_605,In_552,In_1262);
and U606 (N_606,N_322,In_1053);
and U607 (N_607,N_326,In_1451);
nand U608 (N_608,In_257,In_256);
nand U609 (N_609,In_1891,In_1365);
nor U610 (N_610,N_193,In_1532);
or U611 (N_611,N_172,N_254);
and U612 (N_612,In_1467,In_1024);
and U613 (N_613,In_1578,N_315);
and U614 (N_614,In_308,In_1779);
and U615 (N_615,In_954,N_381);
and U616 (N_616,N_70,N_215);
nand U617 (N_617,In_887,In_921);
and U618 (N_618,N_87,In_1780);
and U619 (N_619,In_293,In_1047);
or U620 (N_620,In_385,In_596);
xor U621 (N_621,In_1012,N_147);
nand U622 (N_622,In_712,In_1768);
and U623 (N_623,N_83,In_1336);
nor U624 (N_624,In_13,In_806);
xor U625 (N_625,In_1691,N_214);
or U626 (N_626,N_198,N_165);
or U627 (N_627,In_1671,N_292);
nand U628 (N_628,In_555,In_45);
nand U629 (N_629,In_108,N_24);
xnor U630 (N_630,In_1002,N_71);
xor U631 (N_631,In_1333,In_784);
nand U632 (N_632,In_1438,In_579);
nor U633 (N_633,In_40,In_471);
and U634 (N_634,In_1809,In_1190);
nand U635 (N_635,In_1665,In_1487);
nor U636 (N_636,In_194,In_1260);
nand U637 (N_637,In_1555,In_1725);
nand U638 (N_638,In_1920,N_14);
or U639 (N_639,N_385,N_168);
nor U640 (N_640,In_778,N_113);
or U641 (N_641,In_1840,In_1427);
and U642 (N_642,In_1130,In_1195);
xor U643 (N_643,In_1755,In_1482);
and U644 (N_644,In_71,In_1193);
or U645 (N_645,In_502,N_129);
or U646 (N_646,N_92,N_33);
nand U647 (N_647,In_1300,In_705);
nor U648 (N_648,N_79,In_1393);
or U649 (N_649,In_767,In_1644);
nor U650 (N_650,In_781,N_148);
and U651 (N_651,In_1955,In_1124);
nand U652 (N_652,In_1552,In_1296);
xor U653 (N_653,In_422,In_150);
xnor U654 (N_654,In_733,N_30);
and U655 (N_655,In_233,In_1954);
nand U656 (N_656,N_109,In_627);
or U657 (N_657,N_287,In_962);
and U658 (N_658,In_662,N_53);
and U659 (N_659,In_1436,In_51);
xnor U660 (N_660,In_1945,In_1894);
nor U661 (N_661,In_297,In_565);
and U662 (N_662,In_399,In_1953);
xnor U663 (N_663,In_0,In_761);
and U664 (N_664,In_898,N_390);
nor U665 (N_665,In_1553,In_785);
xor U666 (N_666,In_771,In_835);
xor U667 (N_667,N_256,In_304);
xnor U668 (N_668,In_1961,In_1248);
nor U669 (N_669,In_488,In_1801);
xnor U670 (N_670,In_1182,In_302);
nand U671 (N_671,In_39,In_903);
xor U672 (N_672,In_1839,In_1942);
nand U673 (N_673,In_872,In_542);
xor U674 (N_674,N_223,In_1392);
and U675 (N_675,N_290,N_366);
or U676 (N_676,In_1770,In_525);
xor U677 (N_677,In_207,In_1123);
and U678 (N_678,In_889,N_1);
xor U679 (N_679,In_345,N_270);
nor U680 (N_680,In_454,In_1228);
xor U681 (N_681,In_1221,N_370);
nor U682 (N_682,In_1989,In_350);
or U683 (N_683,In_521,In_1354);
nor U684 (N_684,In_1036,In_1742);
nor U685 (N_685,N_179,In_1079);
or U686 (N_686,In_1604,N_126);
and U687 (N_687,In_1977,In_1539);
or U688 (N_688,N_286,In_1689);
or U689 (N_689,In_807,N_156);
or U690 (N_690,N_210,In_1765);
nor U691 (N_691,N_300,N_115);
nand U692 (N_692,In_1740,N_282);
nand U693 (N_693,In_504,In_362);
or U694 (N_694,In_827,In_576);
or U695 (N_695,N_50,In_328);
xnor U696 (N_696,In_9,In_269);
and U697 (N_697,In_1550,In_1813);
and U698 (N_698,N_12,N_245);
xnor U699 (N_699,In_1104,In_1483);
nor U700 (N_700,N_226,N_22);
and U701 (N_701,In_215,N_59);
and U702 (N_702,In_183,N_304);
xnor U703 (N_703,N_283,In_1218);
and U704 (N_704,N_142,In_1094);
or U705 (N_705,N_201,In_765);
and U706 (N_706,In_1235,In_1363);
xnor U707 (N_707,N_313,In_172);
and U708 (N_708,In_640,In_590);
nor U709 (N_709,In_157,In_1593);
nor U710 (N_710,N_43,In_364);
nor U711 (N_711,In_1720,In_1316);
and U712 (N_712,In_746,In_1722);
nor U713 (N_713,N_5,N_218);
nand U714 (N_714,N_74,N_260);
xnor U715 (N_715,In_513,N_145);
xor U716 (N_716,In_270,In_587);
xnor U717 (N_717,In_1824,In_799);
or U718 (N_718,In_1516,In_1335);
and U719 (N_719,N_25,N_23);
nand U720 (N_720,In_464,In_1981);
xor U721 (N_721,N_125,In_391);
xnor U722 (N_722,In_432,In_200);
or U723 (N_723,N_61,In_547);
or U724 (N_724,N_361,In_1019);
nor U725 (N_725,In_368,N_160);
nor U726 (N_726,In_1361,In_1512);
or U727 (N_727,In_1703,In_1369);
nor U728 (N_728,N_206,N_157);
and U729 (N_729,In_439,In_78);
xor U730 (N_730,In_1283,In_19);
nor U731 (N_731,N_303,In_1383);
xnor U732 (N_732,In_1681,In_1484);
and U733 (N_733,In_1375,In_1226);
or U734 (N_734,In_1525,In_393);
xor U735 (N_735,In_1223,In_417);
or U736 (N_736,In_563,In_238);
nor U737 (N_737,In_1764,N_306);
and U738 (N_738,N_341,In_1909);
and U739 (N_739,In_1225,In_355);
nand U740 (N_740,In_879,In_863);
nor U741 (N_741,In_1216,In_1758);
and U742 (N_742,In_128,In_1973);
nor U743 (N_743,N_384,N_329);
and U744 (N_744,In_1872,In_678);
xor U745 (N_745,In_1209,In_968);
xor U746 (N_746,In_1402,N_36);
or U747 (N_747,In_1099,In_1421);
nor U748 (N_748,In_1915,In_404);
or U749 (N_749,In_703,In_188);
nand U750 (N_750,In_1993,In_341);
xor U751 (N_751,In_1111,In_814);
xor U752 (N_752,In_1191,N_177);
xnor U753 (N_753,N_41,In_167);
and U754 (N_754,In_332,In_1074);
nor U755 (N_755,In_1978,In_1757);
and U756 (N_756,In_684,N_242);
nand U757 (N_757,N_289,In_603);
or U758 (N_758,In_1141,In_736);
xor U759 (N_759,In_354,In_1377);
and U760 (N_760,N_388,In_1298);
nand U761 (N_761,In_523,N_124);
and U762 (N_762,In_1654,N_205);
or U763 (N_763,In_1745,In_742);
nand U764 (N_764,In_400,In_1277);
or U765 (N_765,In_1596,In_1986);
nand U766 (N_766,N_362,In_1264);
and U767 (N_767,In_1448,In_793);
and U768 (N_768,In_530,In_1163);
or U769 (N_769,In_298,N_220);
and U770 (N_770,In_1326,In_1227);
nand U771 (N_771,In_1088,In_608);
nand U772 (N_772,N_267,N_269);
or U773 (N_773,In_980,N_200);
and U774 (N_774,In_1031,N_324);
nor U775 (N_775,In_1845,In_540);
xor U776 (N_776,N_318,In_859);
and U777 (N_777,N_386,N_331);
nor U778 (N_778,In_1253,In_1542);
or U779 (N_779,In_243,In_1068);
xor U780 (N_780,N_102,In_899);
nand U781 (N_781,In_1060,In_1857);
nand U782 (N_782,In_987,N_64);
nand U783 (N_783,In_597,N_119);
nand U784 (N_784,In_711,In_619);
or U785 (N_785,In_1835,In_79);
nand U786 (N_786,N_212,In_100);
and U787 (N_787,In_536,In_717);
and U788 (N_788,In_831,N_120);
and U789 (N_789,In_16,In_1308);
nand U790 (N_790,In_2,N_73);
xor U791 (N_791,In_1692,In_1751);
or U792 (N_792,In_48,In_1303);
xor U793 (N_793,In_1259,In_639);
nor U794 (N_794,N_152,In_1923);
or U795 (N_795,In_882,In_1391);
nand U796 (N_796,In_1292,N_10);
and U797 (N_797,In_1771,In_1491);
nand U798 (N_798,In_1305,In_1576);
nand U799 (N_799,In_920,In_171);
and U800 (N_800,N_761,In_554);
and U801 (N_801,N_746,N_608);
and U802 (N_802,N_682,N_378);
xor U803 (N_803,In_246,N_353);
xnor U804 (N_804,In_1547,In_176);
or U805 (N_805,In_1560,In_1160);
nor U806 (N_806,N_783,N_330);
nand U807 (N_807,N_309,N_547);
nor U808 (N_808,In_151,In_690);
or U809 (N_809,N_8,N_60);
or U810 (N_810,N_560,N_635);
nor U811 (N_811,In_1210,In_193);
xor U812 (N_812,N_512,In_986);
and U813 (N_813,N_566,N_440);
nand U814 (N_814,N_438,In_66);
nand U815 (N_815,N_732,N_182);
nand U816 (N_816,In_95,In_907);
and U817 (N_817,N_589,In_560);
and U818 (N_818,In_512,In_142);
or U819 (N_819,In_944,N_768);
or U820 (N_820,In_1910,In_571);
or U821 (N_821,N_393,In_948);
xnor U822 (N_822,In_401,N_656);
nor U823 (N_823,N_374,N_437);
nand U824 (N_824,In_1398,N_342);
nand U825 (N_825,N_467,In_1468);
and U826 (N_826,In_359,N_711);
xnor U827 (N_827,In_1837,N_339);
xor U828 (N_828,In_1388,In_278);
or U829 (N_829,In_57,N_663);
nor U830 (N_830,In_1455,In_1500);
xor U831 (N_831,In_1446,In_1732);
xor U832 (N_832,In_187,N_687);
nand U833 (N_833,N_785,N_159);
and U834 (N_834,In_1911,N_670);
nor U835 (N_835,In_1325,N_601);
nor U836 (N_836,N_550,N_235);
xnor U837 (N_837,In_1877,In_1933);
or U838 (N_838,In_692,In_936);
nand U839 (N_839,In_1690,In_1183);
and U840 (N_840,N_268,In_1050);
xor U841 (N_841,In_26,In_284);
or U842 (N_842,In_374,In_1648);
nand U843 (N_843,In_999,In_564);
or U844 (N_844,N_739,N_688);
and U845 (N_845,N_536,In_1128);
nand U846 (N_846,In_537,N_425);
nand U847 (N_847,N_546,N_666);
xnor U848 (N_848,N_274,N_482);
nor U849 (N_849,N_94,In_1606);
or U850 (N_850,In_1106,In_1048);
or U851 (N_851,In_1726,In_1949);
or U852 (N_852,In_1151,In_378);
nor U853 (N_853,In_258,N_709);
nand U854 (N_854,In_1401,In_800);
nor U855 (N_855,In_1041,In_1530);
or U856 (N_856,N_492,In_322);
nand U857 (N_857,N_559,N_259);
and U858 (N_858,In_773,In_1174);
nand U859 (N_859,In_928,N_798);
xor U860 (N_860,N_435,N_190);
or U861 (N_861,N_54,In_276);
nand U862 (N_862,In_838,In_1033);
xor U863 (N_863,In_1346,N_707);
or U864 (N_864,In_1005,In_349);
or U865 (N_865,In_567,N_686);
and U866 (N_866,N_423,In_890);
nor U867 (N_867,N_238,N_776);
xnor U868 (N_868,In_254,N_532);
or U869 (N_869,N_577,In_1807);
xnor U870 (N_870,N_454,In_1937);
nand U871 (N_871,In_65,N_548);
and U872 (N_872,In_282,N_412);
nand U873 (N_873,N_579,N_502);
nand U874 (N_874,In_1107,In_1454);
xor U875 (N_875,In_154,In_1657);
xnor U876 (N_876,N_724,In_1494);
nor U877 (N_877,In_949,In_210);
or U878 (N_878,In_763,In_1628);
nor U879 (N_879,In_1474,N_680);
or U880 (N_880,In_913,In_599);
nor U881 (N_881,N_748,In_1464);
nand U882 (N_882,N_343,N_75);
nand U883 (N_883,In_1971,N_213);
xor U884 (N_884,N_409,N_728);
and U885 (N_885,In_110,In_852);
nor U886 (N_886,In_316,N_702);
or U887 (N_887,N_779,N_597);
or U888 (N_888,N_576,In_704);
or U889 (N_889,N_657,N_529);
nor U890 (N_890,N_510,In_168);
nand U891 (N_891,In_1188,N_653);
or U892 (N_892,In_69,In_221);
and U893 (N_893,N_745,N_784);
and U894 (N_894,In_984,In_1959);
nor U895 (N_895,In_881,N_508);
or U896 (N_896,In_46,In_659);
xnor U897 (N_897,In_1699,N_471);
xor U898 (N_898,In_1295,N_475);
or U899 (N_899,In_443,N_457);
or U900 (N_900,N_493,In_1655);
nand U901 (N_901,N_278,N_216);
xnor U902 (N_902,N_498,In_1633);
nor U903 (N_903,N_477,N_392);
xnor U904 (N_904,In_770,In_1709);
nand U905 (N_905,In_1044,In_224);
or U906 (N_906,N_698,In_910);
nand U907 (N_907,N_552,N_519);
and U908 (N_908,N_497,In_1409);
xnor U909 (N_909,In_724,In_406);
or U910 (N_910,In_1239,N_565);
and U911 (N_911,N_66,In_1828);
nand U912 (N_912,In_112,In_1946);
xnor U913 (N_913,N_360,In_668);
or U914 (N_914,N_443,N_534);
xor U915 (N_915,In_730,In_735);
or U916 (N_916,In_1285,In_251);
nand U917 (N_917,In_1748,In_1051);
or U918 (N_918,In_1829,In_76);
or U919 (N_919,In_1972,N_65);
nor U920 (N_920,In_1204,In_713);
and U921 (N_921,In_1178,In_1077);
nand U922 (N_922,In_5,N_414);
and U923 (N_923,N_752,N_708);
nor U924 (N_924,In_1236,In_850);
or U925 (N_925,N_727,In_1412);
xnor U926 (N_926,N_436,N_478);
or U927 (N_927,N_389,N_716);
nor U928 (N_928,In_682,In_931);
and U929 (N_929,N_693,N_465);
or U930 (N_930,In_1930,N_195);
nor U931 (N_931,N_578,N_541);
nor U932 (N_932,In_1508,N_648);
nand U933 (N_933,N_525,N_544);
nand U934 (N_934,N_227,N_356);
or U935 (N_935,In_766,In_620);
and U936 (N_936,In_178,N_659);
xor U937 (N_937,N_187,In_1577);
nor U938 (N_938,In_1640,N_617);
xnor U939 (N_939,In_1563,In_1645);
nor U940 (N_940,In_581,In_1073);
or U941 (N_941,N_594,In_953);
or U942 (N_942,N_614,N_564);
nor U943 (N_943,N_660,N_346);
or U944 (N_944,N_794,In_32);
nor U945 (N_945,In_429,N_787);
and U946 (N_946,In_1592,In_1481);
nand U947 (N_947,N_554,N_585);
nor U948 (N_948,In_346,N_453);
xnor U949 (N_949,In_149,N_461);
xnor U950 (N_950,N_382,In_988);
xnor U951 (N_951,In_1513,In_1622);
or U952 (N_952,In_1983,N_429);
or U953 (N_953,In_1922,In_3);
or U954 (N_954,N_13,N_332);
nand U955 (N_955,N_676,N_232);
or U956 (N_956,N_11,N_769);
or U957 (N_957,In_325,In_245);
nand U958 (N_958,In_1330,N_562);
or U959 (N_959,N_651,In_1686);
nand U960 (N_960,N_18,N_158);
nand U961 (N_961,In_688,N_522);
nand U962 (N_962,N_0,N_773);
and U963 (N_963,In_72,N_506);
nor U964 (N_964,In_624,N_399);
or U965 (N_965,N_420,In_1653);
nor U966 (N_966,In_231,In_1528);
or U967 (N_967,N_459,In_180);
or U968 (N_968,N_528,N_791);
xor U969 (N_969,In_958,N_613);
nand U970 (N_970,In_1129,N_630);
or U971 (N_971,N_416,N_89);
and U972 (N_972,In_768,N_751);
nor U973 (N_973,In_91,N_710);
or U974 (N_974,N_621,N_462);
nor U975 (N_975,N_116,In_1781);
or U976 (N_976,N_261,In_1760);
nand U977 (N_977,In_1544,In_1905);
xor U978 (N_978,In_22,In_1157);
or U979 (N_979,In_214,N_276);
nor U980 (N_980,N_49,In_120);
nor U981 (N_981,N_451,N_349);
xor U982 (N_982,N_225,In_47);
xnor U983 (N_983,In_1172,In_1842);
nor U984 (N_984,In_1974,N_249);
or U985 (N_985,N_394,In_1379);
nor U986 (N_986,N_67,In_466);
nor U987 (N_987,In_1599,N_640);
xnor U988 (N_988,N_405,N_444);
and U989 (N_989,In_153,In_1134);
xnor U990 (N_990,N_486,In_1465);
nor U991 (N_991,In_1233,N_183);
and U992 (N_992,N_44,N_755);
or U993 (N_993,N_759,In_976);
nand U994 (N_994,N_740,In_1594);
nor U995 (N_995,In_562,N_774);
nor U996 (N_996,In_1631,In_97);
nand U997 (N_997,N_427,In_1580);
or U998 (N_998,N_105,N_47);
or U999 (N_999,In_85,In_323);
nor U1000 (N_1000,In_1999,N_770);
or U1001 (N_1001,N_797,N_627);
or U1002 (N_1002,N_470,In_1478);
and U1003 (N_1003,In_411,In_452);
nor U1004 (N_1004,In_33,N_189);
or U1005 (N_1005,N_526,N_112);
xnor U1006 (N_1006,N_55,N_551);
nand U1007 (N_1007,N_569,N_151);
nand U1008 (N_1008,In_908,N_333);
or U1009 (N_1009,In_622,N_741);
or U1010 (N_1010,N_291,N_607);
or U1011 (N_1011,In_1119,N_489);
nand U1012 (N_1012,In_262,In_1035);
xor U1013 (N_1013,N_163,N_474);
and U1014 (N_1014,N_219,N_424);
and U1015 (N_1015,In_487,N_17);
or U1016 (N_1016,In_1148,N_644);
nor U1017 (N_1017,In_1607,In_721);
nor U1018 (N_1018,In_1908,N_790);
and U1019 (N_1019,In_1282,In_1741);
nor U1020 (N_1020,N_82,In_593);
nand U1021 (N_1021,In_963,In_1524);
nand U1022 (N_1022,In_534,N_775);
xnor U1023 (N_1023,N_480,N_224);
or U1024 (N_1024,N_312,N_344);
nor U1025 (N_1025,N_624,N_778);
nand U1026 (N_1026,In_893,N_234);
xnor U1027 (N_1027,N_391,N_530);
nor U1028 (N_1028,N_110,In_1001);
and U1029 (N_1029,In_598,In_1016);
and U1030 (N_1030,N_111,In_306);
nor U1031 (N_1031,N_265,In_1351);
nor U1032 (N_1032,In_1940,In_1396);
and U1033 (N_1033,N_679,In_1600);
or U1034 (N_1034,In_1597,N_208);
nor U1035 (N_1035,N_297,In_1147);
xor U1036 (N_1036,N_762,In_633);
nand U1037 (N_1037,N_32,N_138);
xor U1038 (N_1038,In_1261,N_169);
or U1039 (N_1039,In_896,N_556);
or U1040 (N_1040,In_1417,N_691);
or U1041 (N_1041,In_1502,N_623);
nand U1042 (N_1042,In_541,N_667);
or U1043 (N_1043,In_1080,In_225);
xor U1044 (N_1044,N_140,In_1847);
xnor U1045 (N_1045,N_596,N_266);
xnor U1046 (N_1046,N_504,In_1881);
and U1047 (N_1047,N_580,N_592);
and U1048 (N_1048,N_408,N_397);
nor U1049 (N_1049,In_107,In_1789);
and U1050 (N_1050,N_531,N_558);
xnor U1051 (N_1051,In_1867,N_230);
or U1052 (N_1052,In_1347,In_198);
xor U1053 (N_1053,N_618,N_641);
nor U1054 (N_1054,In_1132,In_1334);
and U1055 (N_1055,In_1815,N_520);
or U1056 (N_1056,N_314,In_261);
or U1057 (N_1057,N_355,In_851);
and U1058 (N_1058,N_722,N_729);
or U1059 (N_1059,In_410,In_353);
xor U1060 (N_1060,N_48,N_77);
nor U1061 (N_1061,In_1242,N_674);
xnor U1062 (N_1062,In_691,In_511);
or U1063 (N_1063,N_307,N_542);
xnor U1064 (N_1064,In_1408,N_413);
and U1065 (N_1065,N_507,In_1533);
or U1066 (N_1066,N_675,N_442);
nor U1067 (N_1067,In_162,N_448);
and U1068 (N_1068,N_696,In_983);
nor U1069 (N_1069,N_426,N_587);
nor U1070 (N_1070,N_328,N_117);
xnor U1071 (N_1071,In_966,N_197);
xnor U1072 (N_1072,In_775,N_673);
xor U1073 (N_1073,In_701,N_634);
or U1074 (N_1074,N_288,N_63);
nor U1075 (N_1075,N_524,N_26);
nand U1076 (N_1076,N_162,N_637);
and U1077 (N_1077,N_726,N_599);
nand U1078 (N_1078,N_272,In_1776);
xor U1079 (N_1079,In_1649,In_805);
nand U1080 (N_1080,In_334,N_628);
or U1081 (N_1081,In_1329,N_417);
xnor U1082 (N_1082,N_799,In_1851);
xor U1083 (N_1083,N_57,In_663);
nor U1084 (N_1084,In_934,N_725);
nand U1085 (N_1085,In_1642,N_433);
or U1086 (N_1086,In_1022,In_870);
or U1087 (N_1087,In_1198,In_56);
nand U1088 (N_1088,N_280,In_89);
xnor U1089 (N_1089,In_1066,N_136);
and U1090 (N_1090,N_422,In_1220);
xor U1091 (N_1091,In_1297,N_757);
nand U1092 (N_1092,In_186,In_473);
or U1093 (N_1093,In_566,N_620);
and U1094 (N_1094,In_179,In_1212);
nand U1095 (N_1095,N_180,N_539);
and U1096 (N_1096,N_655,N_167);
nand U1097 (N_1097,N_731,N_591);
nor U1098 (N_1098,In_1169,In_864);
nand U1099 (N_1099,In_1318,N_719);
nor U1100 (N_1100,N_733,In_812);
nand U1101 (N_1101,N_317,N_588);
xnor U1102 (N_1102,In_94,N_521);
nor U1103 (N_1103,N_501,In_343);
or U1104 (N_1104,N_284,N_466);
nor U1105 (N_1105,In_1150,N_154);
or U1106 (N_1106,In_1255,N_572);
and U1107 (N_1107,N_255,N_683);
nand U1108 (N_1108,In_81,In_1980);
nand U1109 (N_1109,In_1941,In_1029);
xor U1110 (N_1110,N_188,N_460);
and U1111 (N_1111,N_694,N_598);
nand U1112 (N_1112,N_730,In_892);
or U1113 (N_1113,In_1859,N_652);
and U1114 (N_1114,In_310,In_77);
nand U1115 (N_1115,In_68,N_777);
xor U1116 (N_1116,N_472,In_437);
nor U1117 (N_1117,N_221,In_876);
xnor U1118 (N_1118,N_407,N_352);
xnor U1119 (N_1119,In_281,N_713);
nor U1120 (N_1120,In_137,N_545);
nand U1121 (N_1121,In_138,In_1792);
nand U1122 (N_1122,N_153,In_14);
nand U1123 (N_1123,N_45,In_548);
nor U1124 (N_1124,N_91,N_571);
and U1125 (N_1125,In_117,In_1087);
xnor U1126 (N_1126,In_388,In_1884);
xor U1127 (N_1127,In_1013,N_518);
or U1128 (N_1128,In_6,In_969);
and U1129 (N_1129,N_712,N_35);
xor U1130 (N_1130,In_320,N_240);
xnor U1131 (N_1131,In_235,N_636);
nor U1132 (N_1132,N_495,N_734);
xnor U1133 (N_1133,N_611,In_1960);
xor U1134 (N_1134,In_819,In_456);
xor U1135 (N_1135,N_93,In_465);
or U1136 (N_1136,N_51,In_847);
nand U1137 (N_1137,In_55,N_354);
or U1138 (N_1138,N_455,N_796);
and U1139 (N_1139,N_609,In_1324);
nor U1140 (N_1140,N_780,In_135);
nor U1141 (N_1141,N_294,In_305);
nand U1142 (N_1142,In_133,In_508);
nor U1143 (N_1143,In_423,In_491);
or U1144 (N_1144,N_582,N_400);
and U1145 (N_1145,In_826,In_1177);
xnor U1146 (N_1146,In_947,In_1650);
and U1147 (N_1147,N_747,N_662);
xnor U1148 (N_1148,N_782,N_665);
or U1149 (N_1149,In_1529,N_253);
and U1150 (N_1150,N_754,In_1422);
xor U1151 (N_1151,In_156,In_524);
or U1152 (N_1152,N_650,N_468);
nand U1153 (N_1153,N_789,In_1919);
or U1154 (N_1154,N_431,N_714);
and U1155 (N_1155,In_329,In_12);
or U1156 (N_1156,In_227,In_1746);
or U1157 (N_1157,N_758,N_700);
xnor U1158 (N_1158,In_1302,In_1374);
or U1159 (N_1159,In_1612,N_469);
or U1160 (N_1160,N_441,N_481);
xnor U1161 (N_1161,In_1092,In_1307);
xor U1162 (N_1162,In_661,In_1251);
nor U1163 (N_1163,N_750,In_580);
or U1164 (N_1164,In_232,In_629);
nor U1165 (N_1165,N_661,In_462);
xnor U1166 (N_1166,In_288,In_101);
xor U1167 (N_1167,In_744,N_622);
nor U1168 (N_1168,In_1718,In_414);
or U1169 (N_1169,N_654,N_418);
or U1170 (N_1170,N_345,In_1574);
nor U1171 (N_1171,N_781,N_452);
or U1172 (N_1172,In_1085,In_505);
and U1173 (N_1173,In_1762,In_132);
and U1174 (N_1174,N_363,N_401);
or U1175 (N_1175,In_119,N_80);
or U1176 (N_1176,N_127,N_645);
and U1177 (N_1177,In_985,N_535);
xnor U1178 (N_1178,N_681,N_40);
nor U1179 (N_1179,In_719,N_487);
nand U1180 (N_1180,N_788,N_456);
xor U1181 (N_1181,N_513,In_1034);
xor U1182 (N_1182,N_323,In_1685);
and U1183 (N_1183,N_737,In_1249);
nor U1184 (N_1184,N_181,N_445);
and U1185 (N_1185,N_658,In_621);
and U1186 (N_1186,N_229,N_616);
xnor U1187 (N_1187,N_131,In_1006);
nor U1188 (N_1188,N_570,N_772);
and U1189 (N_1189,N_150,N_567);
nor U1190 (N_1190,N_606,In_836);
xor U1191 (N_1191,N_699,In_1142);
nor U1192 (N_1192,N_37,N_557);
xor U1193 (N_1193,N_146,N_351);
nor U1194 (N_1194,N_302,N_428);
xnor U1195 (N_1195,In_1988,N_239);
nor U1196 (N_1196,N_372,In_1486);
or U1197 (N_1197,In_1205,In_363);
nand U1198 (N_1198,In_326,N_246);
or U1199 (N_1199,N_689,N_96);
nor U1200 (N_1200,N_1106,In_1651);
nand U1201 (N_1201,N_850,N_1061);
nor U1202 (N_1202,In_61,N_997);
nor U1203 (N_1203,N_1089,N_753);
and U1204 (N_1204,In_1397,In_340);
xnor U1205 (N_1205,N_921,N_885);
xor U1206 (N_1206,In_874,In_169);
xnor U1207 (N_1207,N_804,N_533);
nand U1208 (N_1208,N_836,N_336);
xnor U1209 (N_1209,N_1005,N_473);
nand U1210 (N_1210,In_1109,N_1169);
nor U1211 (N_1211,N_1181,In_1155);
xnor U1212 (N_1212,N_923,N_170);
nand U1213 (N_1213,N_1029,N_900);
or U1214 (N_1214,N_1056,In_901);
xnor U1215 (N_1215,N_867,In_1979);
and U1216 (N_1216,N_1127,N_1085);
nor U1217 (N_1217,N_705,N_1126);
nand U1218 (N_1218,In_965,N_1063);
xor U1219 (N_1219,N_677,In_1570);
nand U1220 (N_1220,N_834,N_1151);
nor U1221 (N_1221,In_405,N_615);
nor U1222 (N_1222,N_1018,N_695);
or U1223 (N_1223,In_1716,N_1094);
nor U1224 (N_1224,N_1038,In_1998);
and U1225 (N_1225,N_802,N_1104);
xnor U1226 (N_1226,In_911,N_410);
nand U1227 (N_1227,In_1364,N_845);
or U1228 (N_1228,N_1194,N_977);
nor U1229 (N_1229,In_324,In_1247);
or U1230 (N_1230,N_1067,N_563);
nand U1231 (N_1231,N_511,N_505);
or U1232 (N_1232,N_1009,N_878);
nor U1233 (N_1233,N_1110,N_718);
nor U1234 (N_1234,N_237,N_1189);
nor U1235 (N_1235,N_955,N_926);
nand U1236 (N_1236,N_912,N_984);
or U1237 (N_1237,In_589,In_1089);
and U1238 (N_1238,N_1195,In_783);
or U1239 (N_1239,N_1052,In_1306);
nor U1240 (N_1240,N_950,N_866);
nor U1241 (N_1241,In_1786,N_888);
nand U1242 (N_1242,In_1682,In_267);
nand U1243 (N_1243,N_419,In_638);
xor U1244 (N_1244,In_1268,N_896);
xor U1245 (N_1245,N_792,In_697);
nand U1246 (N_1246,N_1191,N_31);
and U1247 (N_1247,N_643,In_1658);
and U1248 (N_1248,N_988,In_344);
nand U1249 (N_1249,In_606,In_1390);
nor U1250 (N_1250,In_1549,N_838);
and U1251 (N_1251,N_966,N_1123);
or U1252 (N_1252,N_947,N_865);
xor U1253 (N_1253,N_1032,N_924);
xnor U1254 (N_1254,N_1113,In_743);
nor U1255 (N_1255,N_857,N_359);
or U1256 (N_1256,N_911,N_1096);
and U1257 (N_1257,N_813,N_816);
and U1258 (N_1258,In_321,In_610);
nand U1259 (N_1259,N_364,In_1509);
xnor U1260 (N_1260,N_1115,N_756);
and U1261 (N_1261,N_721,In_792);
and U1262 (N_1262,N_820,In_1916);
or U1263 (N_1263,N_875,N_899);
nor U1264 (N_1264,N_938,N_893);
nand U1265 (N_1265,In_1843,N_843);
nand U1266 (N_1266,N_1058,N_1059);
and U1267 (N_1267,N_149,N_1073);
nand U1268 (N_1268,N_1003,N_908);
nor U1269 (N_1269,N_952,N_851);
nand U1270 (N_1270,N_1171,In_1007);
or U1271 (N_1271,N_583,N_1139);
nand U1272 (N_1272,N_494,N_1071);
xor U1273 (N_1273,N_678,N_350);
nor U1274 (N_1274,N_1015,In_868);
or U1275 (N_1275,N_999,N_1105);
nor U1276 (N_1276,In_1969,In_825);
nor U1277 (N_1277,N_479,N_1045);
nor U1278 (N_1278,N_1060,In_1343);
xor U1279 (N_1279,N_876,In_1280);
or U1280 (N_1280,N_825,N_987);
nand U1281 (N_1281,N_812,N_1008);
nor U1282 (N_1282,N_1155,N_603);
or U1283 (N_1283,N_1116,In_1666);
xnor U1284 (N_1284,N_959,N_1066);
nand U1285 (N_1285,N_1021,N_1124);
xor U1286 (N_1286,N_496,N_826);
or U1287 (N_1287,In_574,In_1595);
xor U1288 (N_1288,N_1174,In_500);
and U1289 (N_1289,N_509,N_800);
or U1290 (N_1290,N_720,N_856);
nand U1291 (N_1291,N_901,N_1054);
xor U1292 (N_1292,In_1566,N_1088);
and U1293 (N_1293,N_744,N_965);
nor U1294 (N_1294,In_877,In_658);
nor U1295 (N_1295,N_704,N_920);
nor U1296 (N_1296,N_973,N_1037);
nand U1297 (N_1297,In_1286,N_803);
nor U1298 (N_1298,N_593,N_862);
nand U1299 (N_1299,N_949,N_584);
nor U1300 (N_1300,In_479,In_1898);
nor U1301 (N_1301,N_928,N_1025);
nand U1302 (N_1302,N_786,N_1184);
or U1303 (N_1303,In_672,N_69);
and U1304 (N_1304,In_1023,N_1186);
and U1305 (N_1305,N_1142,N_922);
nand U1306 (N_1306,N_1095,In_1434);
and U1307 (N_1307,N_980,N_974);
nand U1308 (N_1308,N_1043,N_946);
nand U1309 (N_1309,N_805,N_824);
nand U1310 (N_1310,In_1803,N_1074);
nor U1311 (N_1311,In_1678,N_723);
or U1312 (N_1312,N_827,N_76);
nor U1313 (N_1313,N_1084,In_211);
and U1314 (N_1314,N_403,N_1010);
xor U1315 (N_1315,In_1476,N_595);
or U1316 (N_1316,In_612,N_819);
nor U1317 (N_1317,N_1107,N_815);
or U1318 (N_1318,N_275,N_629);
and U1319 (N_1319,N_685,N_421);
nor U1320 (N_1320,N_764,N_1079);
xnor U1321 (N_1321,In_1014,N_954);
nand U1322 (N_1322,N_1164,N_638);
xnor U1323 (N_1323,N_517,N_1097);
or U1324 (N_1324,In_1743,N_1093);
nand U1325 (N_1325,N_811,N_642);
nor U1326 (N_1326,N_1198,In_1199);
and U1327 (N_1327,N_1120,N_101);
or U1328 (N_1328,In_803,N_844);
nor U1329 (N_1329,N_996,N_602);
nand U1330 (N_1330,N_823,N_978);
xor U1331 (N_1331,N_1065,In_1368);
or U1332 (N_1332,N_1048,N_916);
nand U1333 (N_1333,N_166,In_1865);
xor U1334 (N_1334,N_887,N_1016);
and U1335 (N_1335,In_1667,N_228);
nand U1336 (N_1336,N_961,N_1128);
nor U1337 (N_1337,N_807,N_742);
nor U1338 (N_1338,In_1880,N_1149);
nand U1339 (N_1339,In_1778,N_4);
nand U1340 (N_1340,N_873,N_19);
xor U1341 (N_1341,N_945,In_118);
nor U1342 (N_1342,N_940,N_894);
nand U1343 (N_1343,N_1167,N_483);
nor U1344 (N_1344,N_877,N_573);
nor U1345 (N_1345,N_503,N_821);
xnor U1346 (N_1346,In_289,N_1047);
and U1347 (N_1347,N_1030,N_766);
nor U1348 (N_1348,In_1535,In_1777);
nor U1349 (N_1349,N_1178,N_1160);
and U1350 (N_1350,N_1082,N_1134);
nand U1351 (N_1351,N_1154,N_327);
and U1352 (N_1352,In_725,N_1119);
nand U1353 (N_1353,In_1982,N_860);
nor U1354 (N_1354,N_176,N_848);
and U1355 (N_1355,In_909,In_1717);
nand U1356 (N_1356,N_830,N_406);
xnor U1357 (N_1357,N_951,N_523);
and U1358 (N_1358,In_617,In_1355);
nand U1359 (N_1359,N_1137,In_1028);
or U1360 (N_1360,N_715,N_171);
or U1361 (N_1361,In_1488,N_1158);
and U1362 (N_1362,N_402,N_411);
or U1363 (N_1363,In_436,N_869);
nand U1364 (N_1364,N_1011,In_1639);
or U1365 (N_1365,N_994,N_818);
or U1366 (N_1366,In_1994,In_460);
nor U1367 (N_1367,In_1914,N_1004);
xor U1368 (N_1368,N_967,N_27);
nand U1369 (N_1369,N_749,N_806);
xnor U1370 (N_1370,In_497,N_1050);
xor U1371 (N_1371,N_325,In_681);
and U1372 (N_1372,In_182,N_1122);
xnor U1373 (N_1373,In_315,In_945);
nor U1374 (N_1374,N_1135,N_703);
xnor U1375 (N_1375,N_809,N_1017);
or U1376 (N_1376,N_874,In_1135);
and U1377 (N_1377,N_814,N_1068);
or U1378 (N_1378,In_197,N_972);
nor U1379 (N_1379,In_129,In_1301);
xnor U1380 (N_1380,N_537,N_853);
nor U1381 (N_1381,N_852,N_846);
and U1382 (N_1382,N_992,N_244);
nand U1383 (N_1383,N_910,N_1153);
xor U1384 (N_1384,N_100,N_1196);
nor U1385 (N_1385,N_902,In_327);
nor U1386 (N_1386,N_839,N_430);
nand U1387 (N_1387,In_1356,In_1662);
xor U1388 (N_1388,N_1078,N_932);
xnor U1389 (N_1389,N_586,N_612);
or U1390 (N_1390,In_577,In_1632);
nor U1391 (N_1391,N_817,N_871);
xor U1392 (N_1392,N_15,In_75);
or U1393 (N_1393,In_1049,N_879);
nand U1394 (N_1394,N_1042,N_488);
nor U1395 (N_1395,N_801,N_1019);
nand U1396 (N_1396,N_387,In_433);
or U1397 (N_1397,N_626,N_1111);
xor U1398 (N_1398,N_717,N_217);
nor U1399 (N_1399,In_470,N_991);
nor U1400 (N_1400,N_913,N_736);
nor U1401 (N_1401,N_968,N_130);
xor U1402 (N_1402,N_1132,N_1023);
and U1403 (N_1403,N_960,N_738);
nand U1404 (N_1404,In_1256,In_53);
and U1405 (N_1405,N_1118,N_767);
nand U1406 (N_1406,In_642,N_976);
and U1407 (N_1407,In_216,N_540);
nor U1408 (N_1408,N_485,N_863);
and U1409 (N_1409,N_376,N_1177);
or U1410 (N_1410,N_561,In_1790);
xor U1411 (N_1411,N_1041,N_1140);
and U1412 (N_1412,N_1121,N_633);
nor U1413 (N_1413,In_1581,In_1615);
nand U1414 (N_1414,N_1136,In_1103);
and U1415 (N_1415,N_277,In_514);
nand U1416 (N_1416,N_439,N_986);
and U1417 (N_1417,N_1165,In_1714);
xnor U1418 (N_1418,N_476,N_191);
xor U1419 (N_1419,N_918,N_1114);
nand U1420 (N_1420,N_931,N_998);
xnor U1421 (N_1421,N_684,N_574);
nor U1422 (N_1422,In_377,N_842);
or U1423 (N_1423,N_884,N_1193);
or U1424 (N_1424,In_1814,N_841);
nand U1425 (N_1425,N_697,N_1057);
nor U1426 (N_1426,N_203,In_166);
xnor U1427 (N_1427,N_516,N_549);
and U1428 (N_1428,N_1168,N_672);
or U1429 (N_1429,In_11,N_1012);
nand U1430 (N_1430,N_919,In_457);
or U1431 (N_1431,N_1125,N_970);
xor U1432 (N_1432,N_449,N_1112);
nand U1433 (N_1433,In_971,N_404);
and U1434 (N_1434,N_1080,N_1033);
xnor U1435 (N_1435,N_917,N_211);
and U1436 (N_1436,N_1157,N_925);
and U1437 (N_1437,N_432,N_625);
xnor U1438 (N_1438,N_858,N_1083);
xnor U1439 (N_1439,N_849,N_1062);
nand U1440 (N_1440,N_1000,In_239);
nor U1441 (N_1441,In_1782,N_1159);
nand U1442 (N_1442,N_1141,In_1721);
nor U1443 (N_1443,N_983,N_1090);
or U1444 (N_1444,N_1035,N_929);
or U1445 (N_1445,N_447,N_937);
nor U1446 (N_1446,N_1145,N_139);
or U1447 (N_1447,N_1086,N_133);
or U1448 (N_1448,In_957,N_944);
nor U1449 (N_1449,N_1002,N_1087);
or U1450 (N_1450,In_616,N_793);
nor U1451 (N_1451,N_600,In_1419);
and U1452 (N_1452,N_1197,N_957);
or U1453 (N_1453,N_958,In_1832);
or U1454 (N_1454,In_1447,In_578);
xnor U1455 (N_1455,N_334,N_969);
nor U1456 (N_1456,N_892,N_1138);
and U1457 (N_1457,N_95,N_88);
nor U1458 (N_1458,N_895,N_490);
or U1459 (N_1459,In_1903,N_971);
nand U1460 (N_1460,In_1695,In_1554);
xor U1461 (N_1461,N_765,N_904);
and U1462 (N_1462,N_377,N_907);
or U1463 (N_1463,N_632,N_1179);
xnor U1464 (N_1464,N_1108,In_607);
nor U1465 (N_1465,In_1359,N_1182);
and U1466 (N_1466,N_103,N_514);
or U1467 (N_1467,N_982,N_861);
or U1468 (N_1468,N_935,N_847);
and U1469 (N_1469,N_1192,N_905);
nand U1470 (N_1470,N_882,In_841);
and U1471 (N_1471,N_241,In_613);
nand U1472 (N_1472,N_1188,In_1208);
nor U1473 (N_1473,In_1641,In_1372);
or U1474 (N_1474,N_1183,N_897);
and U1475 (N_1475,N_375,N_1131);
nand U1476 (N_1476,N_1166,N_735);
and U1477 (N_1477,In_1543,N_16);
nor U1478 (N_1478,N_934,N_371);
or U1479 (N_1479,In_1162,In_1469);
xor U1480 (N_1480,In_482,N_499);
and U1481 (N_1481,In_384,N_62);
nor U1482 (N_1482,N_1049,N_299);
xnor U1483 (N_1483,N_883,N_664);
nand U1484 (N_1484,N_1053,N_568);
xnor U1485 (N_1485,N_1175,N_1176);
or U1486 (N_1486,In_73,N_1075);
and U1487 (N_1487,N_810,N_458);
xnor U1488 (N_1488,In_1189,N_639);
or U1489 (N_1489,N_279,In_750);
xnor U1490 (N_1490,N_962,N_943);
nor U1491 (N_1491,N_906,In_853);
nand U1492 (N_1492,In_490,N_1044);
nor U1493 (N_1493,In_1097,N_1133);
and U1494 (N_1494,N_1064,In_416);
nor U1495 (N_1495,N_1187,N_936);
or U1496 (N_1496,In_147,N_975);
nor U1497 (N_1497,N_575,N_463);
or U1498 (N_1498,N_1109,In_1145);
nand U1499 (N_1499,N_1069,In_716);
nand U1500 (N_1500,N_1161,N_1190);
and U1501 (N_1501,In_978,N_515);
nor U1502 (N_1502,N_1099,N_1006);
and U1503 (N_1503,N_671,N_1102);
nand U1504 (N_1504,N_979,In_248);
nand U1505 (N_1505,N_1055,In_967);
xor U1506 (N_1506,N_828,In_1744);
xor U1507 (N_1507,N_956,N_1031);
and U1508 (N_1508,N_859,N_771);
nor U1509 (N_1509,N_890,N_1040);
nor U1510 (N_1510,N_491,In_528);
nand U1511 (N_1511,N_692,N_379);
nor U1512 (N_1512,In_109,N_1070);
or U1513 (N_1513,In_1536,N_837);
or U1514 (N_1514,In_386,N_1092);
xnor U1515 (N_1515,N_808,N_484);
nor U1516 (N_1516,N_1180,N_868);
nor U1517 (N_1517,N_135,N_97);
or U1518 (N_1518,N_527,In_1670);
nand U1519 (N_1519,N_941,N_701);
xnor U1520 (N_1520,N_649,In_1192);
or U1521 (N_1521,N_1173,In_1293);
nor U1522 (N_1522,In_1934,N_123);
or U1523 (N_1523,N_891,N_46);
nor U1524 (N_1524,N_915,N_953);
xor U1525 (N_1525,N_647,N_1199);
and U1526 (N_1526,N_590,In_1888);
and U1527 (N_1527,N_870,In_904);
and U1528 (N_1528,In_1630,N_822);
or U1529 (N_1529,In_1510,N_1001);
xnor U1530 (N_1530,N_964,N_914);
xnor U1531 (N_1531,In_1875,In_1173);
xnor U1532 (N_1532,N_1156,In_408);
and U1533 (N_1533,In_413,N_1148);
nand U1534 (N_1534,In_1056,N_106);
nor U1535 (N_1535,N_881,N_1026);
or U1536 (N_1536,N_1013,N_446);
nor U1537 (N_1537,N_989,N_990);
nor U1538 (N_1538,N_610,N_1081);
nor U1539 (N_1539,In_866,N_1144);
xor U1540 (N_1540,In_1015,N_338);
nor U1541 (N_1541,N_760,N_829);
nor U1542 (N_1542,N_864,N_763);
nor U1543 (N_1543,N_604,N_985);
xor U1544 (N_1544,N_1162,N_795);
nand U1545 (N_1545,N_855,N_1072);
or U1546 (N_1546,N_415,N_903);
xnor U1547 (N_1547,N_927,N_948);
nor U1548 (N_1548,N_1117,In_609);
xor U1549 (N_1549,In_1185,In_192);
nor U1550 (N_1550,N_1147,In_666);
nand U1551 (N_1551,N_993,N_898);
nand U1552 (N_1552,In_1246,N_1077);
nand U1553 (N_1553,In_737,N_1091);
and U1554 (N_1554,In_915,N_207);
and U1555 (N_1555,In_1997,N_1036);
nand U1556 (N_1556,N_840,N_543);
xnor U1557 (N_1557,In_1900,N_1185);
nand U1558 (N_1558,In_1852,N_196);
nor U1559 (N_1559,N_380,N_605);
xor U1560 (N_1560,N_743,N_1024);
and U1561 (N_1561,N_646,N_1046);
nand U1562 (N_1562,N_1100,In_426);
nor U1563 (N_1563,In_782,In_1473);
xnor U1564 (N_1564,N_434,N_833);
xor U1565 (N_1565,N_981,In_1490);
or U1566 (N_1566,N_1150,In_1675);
and U1567 (N_1567,N_933,In_67);
and U1568 (N_1568,N_1039,N_854);
xnor U1569 (N_1569,N_1101,N_1028);
and U1570 (N_1570,N_52,In_529);
or U1571 (N_1571,N_1170,N_450);
xor U1572 (N_1572,N_669,N_118);
nor U1573 (N_1573,N_889,N_963);
nand U1574 (N_1574,N_581,N_538);
and U1575 (N_1575,N_619,N_1076);
xnor U1576 (N_1576,N_930,N_84);
or U1577 (N_1577,N_831,N_631);
or U1578 (N_1578,N_886,In_1697);
nand U1579 (N_1579,N_1146,N_1143);
or U1580 (N_1580,N_872,N_1034);
xor U1581 (N_1581,N_995,N_668);
nand U1582 (N_1582,In_1521,N_1103);
nor U1583 (N_1583,N_880,N_1027);
xor U1584 (N_1584,N_1007,N_464);
and U1585 (N_1585,N_1130,N_553);
and U1586 (N_1586,N_340,N_555);
or U1587 (N_1587,N_1020,In_615);
nor U1588 (N_1588,N_1129,N_500);
nor U1589 (N_1589,In_1895,N_942);
nand U1590 (N_1590,N_706,N_690);
xnor U1591 (N_1591,In_780,N_835);
or U1592 (N_1592,In_1153,N_1022);
or U1593 (N_1593,N_1014,N_1172);
nor U1594 (N_1594,In_1679,N_939);
nor U1595 (N_1595,N_1051,In_1579);
nand U1596 (N_1596,N_1098,N_1152);
or U1597 (N_1597,N_1163,In_1897);
nand U1598 (N_1598,N_909,N_832);
nand U1599 (N_1599,N_395,In_952);
nor U1600 (N_1600,N_1450,N_1404);
nand U1601 (N_1601,N_1228,N_1391);
nor U1602 (N_1602,N_1359,N_1216);
nand U1603 (N_1603,N_1380,N_1275);
and U1604 (N_1604,N_1203,N_1267);
nand U1605 (N_1605,N_1377,N_1438);
nor U1606 (N_1606,N_1400,N_1492);
nand U1607 (N_1607,N_1389,N_1313);
nand U1608 (N_1608,N_1514,N_1591);
and U1609 (N_1609,N_1394,N_1338);
or U1610 (N_1610,N_1234,N_1533);
nand U1611 (N_1611,N_1553,N_1350);
nand U1612 (N_1612,N_1596,N_1220);
xor U1613 (N_1613,N_1484,N_1333);
nor U1614 (N_1614,N_1419,N_1523);
and U1615 (N_1615,N_1520,N_1422);
nand U1616 (N_1616,N_1545,N_1204);
nand U1617 (N_1617,N_1294,N_1415);
or U1618 (N_1618,N_1347,N_1363);
and U1619 (N_1619,N_1326,N_1412);
nand U1620 (N_1620,N_1471,N_1570);
and U1621 (N_1621,N_1510,N_1232);
xor U1622 (N_1622,N_1386,N_1240);
nand U1623 (N_1623,N_1339,N_1369);
xor U1624 (N_1624,N_1429,N_1273);
and U1625 (N_1625,N_1399,N_1372);
xnor U1626 (N_1626,N_1513,N_1318);
and U1627 (N_1627,N_1451,N_1512);
xor U1628 (N_1628,N_1324,N_1455);
nand U1629 (N_1629,N_1534,N_1383);
or U1630 (N_1630,N_1280,N_1539);
xnor U1631 (N_1631,N_1327,N_1296);
xnor U1632 (N_1632,N_1384,N_1558);
nand U1633 (N_1633,N_1323,N_1238);
nand U1634 (N_1634,N_1443,N_1348);
nor U1635 (N_1635,N_1258,N_1542);
or U1636 (N_1636,N_1546,N_1241);
nor U1637 (N_1637,N_1448,N_1432);
nor U1638 (N_1638,N_1276,N_1373);
and U1639 (N_1639,N_1223,N_1552);
or U1640 (N_1640,N_1329,N_1571);
xor U1641 (N_1641,N_1439,N_1543);
and U1642 (N_1642,N_1403,N_1365);
and U1643 (N_1643,N_1592,N_1575);
and U1644 (N_1644,N_1544,N_1583);
nand U1645 (N_1645,N_1259,N_1444);
nand U1646 (N_1646,N_1499,N_1319);
nand U1647 (N_1647,N_1370,N_1330);
nand U1648 (N_1648,N_1505,N_1483);
nand U1649 (N_1649,N_1531,N_1494);
nor U1650 (N_1650,N_1222,N_1299);
nand U1651 (N_1651,N_1349,N_1224);
and U1652 (N_1652,N_1547,N_1239);
nor U1653 (N_1653,N_1374,N_1598);
xor U1654 (N_1654,N_1270,N_1581);
nor U1655 (N_1655,N_1211,N_1336);
nor U1656 (N_1656,N_1441,N_1242);
xor U1657 (N_1657,N_1453,N_1248);
nand U1658 (N_1658,N_1388,N_1298);
xnor U1659 (N_1659,N_1532,N_1378);
xor U1660 (N_1660,N_1381,N_1361);
nor U1661 (N_1661,N_1236,N_1507);
nand U1662 (N_1662,N_1231,N_1229);
nand U1663 (N_1663,N_1285,N_1511);
xor U1664 (N_1664,N_1521,N_1501);
xnor U1665 (N_1665,N_1593,N_1467);
xor U1666 (N_1666,N_1337,N_1251);
and U1667 (N_1667,N_1426,N_1564);
nand U1668 (N_1668,N_1476,N_1464);
or U1669 (N_1669,N_1358,N_1376);
nand U1670 (N_1670,N_1408,N_1246);
or U1671 (N_1671,N_1580,N_1207);
or U1672 (N_1672,N_1567,N_1262);
or U1673 (N_1673,N_1306,N_1459);
or U1674 (N_1674,N_1406,N_1230);
xnor U1675 (N_1675,N_1200,N_1456);
or U1676 (N_1676,N_1416,N_1500);
or U1677 (N_1677,N_1260,N_1482);
xor U1678 (N_1678,N_1586,N_1335);
xor U1679 (N_1679,N_1405,N_1574);
and U1680 (N_1680,N_1302,N_1291);
nand U1681 (N_1681,N_1562,N_1263);
or U1682 (N_1682,N_1409,N_1407);
xnor U1683 (N_1683,N_1309,N_1268);
nand U1684 (N_1684,N_1557,N_1414);
or U1685 (N_1685,N_1425,N_1402);
or U1686 (N_1686,N_1469,N_1496);
and U1687 (N_1687,N_1452,N_1588);
and U1688 (N_1688,N_1559,N_1478);
nand U1689 (N_1689,N_1488,N_1418);
or U1690 (N_1690,N_1289,N_1584);
and U1691 (N_1691,N_1481,N_1582);
and U1692 (N_1692,N_1247,N_1366);
and U1693 (N_1693,N_1221,N_1549);
and U1694 (N_1694,N_1274,N_1397);
nor U1695 (N_1695,N_1486,N_1357);
and U1696 (N_1696,N_1215,N_1528);
nand U1697 (N_1697,N_1423,N_1356);
nand U1698 (N_1698,N_1286,N_1340);
xor U1699 (N_1699,N_1427,N_1213);
or U1700 (N_1700,N_1310,N_1460);
nand U1701 (N_1701,N_1568,N_1205);
xor U1702 (N_1702,N_1250,N_1401);
or U1703 (N_1703,N_1487,N_1233);
and U1704 (N_1704,N_1212,N_1579);
xor U1705 (N_1705,N_1252,N_1244);
xnor U1706 (N_1706,N_1332,N_1392);
nor U1707 (N_1707,N_1364,N_1573);
nand U1708 (N_1708,N_1390,N_1504);
xnor U1709 (N_1709,N_1290,N_1410);
or U1710 (N_1710,N_1334,N_1227);
nand U1711 (N_1711,N_1519,N_1537);
and U1712 (N_1712,N_1517,N_1320);
nor U1713 (N_1713,N_1445,N_1555);
nor U1714 (N_1714,N_1253,N_1457);
and U1715 (N_1715,N_1292,N_1540);
and U1716 (N_1716,N_1561,N_1529);
nand U1717 (N_1717,N_1367,N_1526);
and U1718 (N_1718,N_1454,N_1442);
xor U1719 (N_1719,N_1503,N_1430);
and U1720 (N_1720,N_1278,N_1594);
or U1721 (N_1721,N_1282,N_1590);
nand U1722 (N_1722,N_1551,N_1490);
and U1723 (N_1723,N_1300,N_1254);
xor U1724 (N_1724,N_1431,N_1479);
nand U1725 (N_1725,N_1474,N_1465);
xor U1726 (N_1726,N_1343,N_1395);
and U1727 (N_1727,N_1225,N_1281);
or U1728 (N_1728,N_1325,N_1303);
and U1729 (N_1729,N_1345,N_1393);
xnor U1730 (N_1730,N_1530,N_1421);
and U1731 (N_1731,N_1473,N_1351);
nand U1732 (N_1732,N_1226,N_1256);
and U1733 (N_1733,N_1375,N_1447);
xnor U1734 (N_1734,N_1219,N_1498);
nor U1735 (N_1735,N_1209,N_1554);
nand U1736 (N_1736,N_1379,N_1489);
nor U1737 (N_1737,N_1566,N_1522);
xor U1738 (N_1738,N_1437,N_1360);
and U1739 (N_1739,N_1541,N_1560);
or U1740 (N_1740,N_1597,N_1265);
and U1741 (N_1741,N_1550,N_1577);
nor U1742 (N_1742,N_1202,N_1440);
nor U1743 (N_1743,N_1599,N_1536);
or U1744 (N_1744,N_1297,N_1411);
and U1745 (N_1745,N_1589,N_1353);
nand U1746 (N_1746,N_1518,N_1255);
nand U1747 (N_1747,N_1344,N_1436);
or U1748 (N_1748,N_1287,N_1508);
and U1749 (N_1749,N_1434,N_1461);
or U1750 (N_1750,N_1428,N_1527);
nor U1751 (N_1751,N_1271,N_1472);
and U1752 (N_1752,N_1525,N_1509);
and U1753 (N_1753,N_1371,N_1420);
or U1754 (N_1754,N_1572,N_1266);
nand U1755 (N_1755,N_1485,N_1458);
or U1756 (N_1756,N_1328,N_1368);
or U1757 (N_1757,N_1578,N_1214);
nor U1758 (N_1758,N_1516,N_1595);
nand U1759 (N_1759,N_1279,N_1470);
nor U1760 (N_1760,N_1396,N_1311);
xnor U1761 (N_1761,N_1331,N_1321);
or U1762 (N_1762,N_1295,N_1316);
nand U1763 (N_1763,N_1235,N_1312);
nand U1764 (N_1764,N_1283,N_1264);
nand U1765 (N_1765,N_1243,N_1315);
nand U1766 (N_1766,N_1515,N_1272);
nor U1767 (N_1767,N_1468,N_1433);
and U1768 (N_1768,N_1362,N_1210);
nor U1769 (N_1769,N_1317,N_1269);
and U1770 (N_1770,N_1354,N_1424);
nand U1771 (N_1771,N_1217,N_1502);
xnor U1772 (N_1772,N_1382,N_1308);
nor U1773 (N_1773,N_1385,N_1506);
nand U1774 (N_1774,N_1355,N_1304);
nor U1775 (N_1775,N_1206,N_1587);
nor U1776 (N_1776,N_1466,N_1497);
and U1777 (N_1777,N_1341,N_1245);
or U1778 (N_1778,N_1449,N_1462);
xnor U1779 (N_1779,N_1548,N_1352);
xor U1780 (N_1780,N_1565,N_1301);
nand U1781 (N_1781,N_1237,N_1307);
or U1782 (N_1782,N_1314,N_1342);
nor U1783 (N_1783,N_1417,N_1535);
and U1784 (N_1784,N_1463,N_1201);
xor U1785 (N_1785,N_1257,N_1538);
nand U1786 (N_1786,N_1480,N_1249);
nor U1787 (N_1787,N_1475,N_1556);
xor U1788 (N_1788,N_1346,N_1576);
xor U1789 (N_1789,N_1495,N_1446);
xor U1790 (N_1790,N_1293,N_1305);
and U1791 (N_1791,N_1261,N_1477);
xnor U1792 (N_1792,N_1322,N_1387);
nor U1793 (N_1793,N_1569,N_1284);
and U1794 (N_1794,N_1398,N_1277);
xor U1795 (N_1795,N_1413,N_1208);
nand U1796 (N_1796,N_1288,N_1218);
nand U1797 (N_1797,N_1493,N_1491);
and U1798 (N_1798,N_1563,N_1435);
xnor U1799 (N_1799,N_1524,N_1585);
or U1800 (N_1800,N_1363,N_1592);
nor U1801 (N_1801,N_1320,N_1456);
and U1802 (N_1802,N_1366,N_1495);
xor U1803 (N_1803,N_1369,N_1232);
xnor U1804 (N_1804,N_1285,N_1475);
and U1805 (N_1805,N_1477,N_1335);
nor U1806 (N_1806,N_1353,N_1411);
nor U1807 (N_1807,N_1523,N_1325);
xnor U1808 (N_1808,N_1292,N_1505);
nor U1809 (N_1809,N_1574,N_1492);
nor U1810 (N_1810,N_1359,N_1217);
xnor U1811 (N_1811,N_1566,N_1280);
xor U1812 (N_1812,N_1416,N_1552);
and U1813 (N_1813,N_1562,N_1415);
or U1814 (N_1814,N_1327,N_1263);
nor U1815 (N_1815,N_1571,N_1399);
or U1816 (N_1816,N_1343,N_1301);
nor U1817 (N_1817,N_1520,N_1312);
nor U1818 (N_1818,N_1215,N_1579);
nor U1819 (N_1819,N_1583,N_1248);
or U1820 (N_1820,N_1366,N_1540);
and U1821 (N_1821,N_1487,N_1227);
or U1822 (N_1822,N_1327,N_1407);
nor U1823 (N_1823,N_1598,N_1429);
nor U1824 (N_1824,N_1342,N_1489);
xor U1825 (N_1825,N_1456,N_1522);
nand U1826 (N_1826,N_1350,N_1216);
nor U1827 (N_1827,N_1396,N_1475);
and U1828 (N_1828,N_1547,N_1349);
xnor U1829 (N_1829,N_1492,N_1499);
nor U1830 (N_1830,N_1489,N_1454);
nand U1831 (N_1831,N_1519,N_1270);
nand U1832 (N_1832,N_1206,N_1295);
nor U1833 (N_1833,N_1430,N_1494);
nor U1834 (N_1834,N_1481,N_1592);
nor U1835 (N_1835,N_1300,N_1586);
nand U1836 (N_1836,N_1253,N_1586);
or U1837 (N_1837,N_1504,N_1345);
xor U1838 (N_1838,N_1298,N_1353);
xnor U1839 (N_1839,N_1268,N_1417);
xnor U1840 (N_1840,N_1256,N_1384);
or U1841 (N_1841,N_1394,N_1417);
nand U1842 (N_1842,N_1541,N_1256);
xnor U1843 (N_1843,N_1210,N_1527);
nand U1844 (N_1844,N_1435,N_1554);
xor U1845 (N_1845,N_1529,N_1471);
and U1846 (N_1846,N_1229,N_1448);
nand U1847 (N_1847,N_1576,N_1582);
nand U1848 (N_1848,N_1496,N_1296);
or U1849 (N_1849,N_1569,N_1281);
and U1850 (N_1850,N_1495,N_1227);
xnor U1851 (N_1851,N_1331,N_1560);
nor U1852 (N_1852,N_1447,N_1204);
xnor U1853 (N_1853,N_1402,N_1568);
or U1854 (N_1854,N_1299,N_1540);
nor U1855 (N_1855,N_1272,N_1535);
nor U1856 (N_1856,N_1524,N_1273);
xor U1857 (N_1857,N_1533,N_1448);
xnor U1858 (N_1858,N_1587,N_1403);
or U1859 (N_1859,N_1585,N_1440);
xnor U1860 (N_1860,N_1405,N_1507);
xor U1861 (N_1861,N_1231,N_1346);
and U1862 (N_1862,N_1214,N_1450);
or U1863 (N_1863,N_1580,N_1543);
or U1864 (N_1864,N_1348,N_1418);
or U1865 (N_1865,N_1597,N_1538);
xnor U1866 (N_1866,N_1447,N_1527);
and U1867 (N_1867,N_1374,N_1422);
nor U1868 (N_1868,N_1406,N_1413);
nor U1869 (N_1869,N_1231,N_1326);
xor U1870 (N_1870,N_1423,N_1347);
and U1871 (N_1871,N_1460,N_1518);
xnor U1872 (N_1872,N_1253,N_1420);
or U1873 (N_1873,N_1524,N_1261);
or U1874 (N_1874,N_1396,N_1357);
nor U1875 (N_1875,N_1315,N_1225);
and U1876 (N_1876,N_1361,N_1399);
nand U1877 (N_1877,N_1582,N_1595);
nand U1878 (N_1878,N_1328,N_1280);
xor U1879 (N_1879,N_1347,N_1508);
nor U1880 (N_1880,N_1520,N_1367);
and U1881 (N_1881,N_1572,N_1596);
xor U1882 (N_1882,N_1257,N_1450);
and U1883 (N_1883,N_1409,N_1504);
xor U1884 (N_1884,N_1492,N_1596);
and U1885 (N_1885,N_1235,N_1209);
xnor U1886 (N_1886,N_1455,N_1267);
nand U1887 (N_1887,N_1442,N_1345);
or U1888 (N_1888,N_1272,N_1556);
nand U1889 (N_1889,N_1304,N_1588);
and U1890 (N_1890,N_1228,N_1596);
xnor U1891 (N_1891,N_1321,N_1336);
nand U1892 (N_1892,N_1409,N_1404);
and U1893 (N_1893,N_1522,N_1311);
and U1894 (N_1894,N_1338,N_1353);
or U1895 (N_1895,N_1451,N_1516);
or U1896 (N_1896,N_1303,N_1291);
xnor U1897 (N_1897,N_1281,N_1385);
xor U1898 (N_1898,N_1377,N_1324);
or U1899 (N_1899,N_1576,N_1479);
nand U1900 (N_1900,N_1380,N_1225);
or U1901 (N_1901,N_1357,N_1531);
nand U1902 (N_1902,N_1357,N_1535);
xnor U1903 (N_1903,N_1434,N_1563);
nor U1904 (N_1904,N_1286,N_1542);
nand U1905 (N_1905,N_1276,N_1518);
nand U1906 (N_1906,N_1362,N_1217);
and U1907 (N_1907,N_1217,N_1516);
xnor U1908 (N_1908,N_1458,N_1362);
nor U1909 (N_1909,N_1227,N_1248);
nor U1910 (N_1910,N_1324,N_1234);
nor U1911 (N_1911,N_1219,N_1312);
xor U1912 (N_1912,N_1219,N_1434);
nand U1913 (N_1913,N_1271,N_1527);
and U1914 (N_1914,N_1555,N_1451);
and U1915 (N_1915,N_1234,N_1557);
xnor U1916 (N_1916,N_1302,N_1560);
xnor U1917 (N_1917,N_1468,N_1262);
xnor U1918 (N_1918,N_1551,N_1254);
or U1919 (N_1919,N_1377,N_1327);
or U1920 (N_1920,N_1221,N_1446);
and U1921 (N_1921,N_1517,N_1497);
nor U1922 (N_1922,N_1375,N_1318);
xor U1923 (N_1923,N_1581,N_1371);
xnor U1924 (N_1924,N_1228,N_1543);
xor U1925 (N_1925,N_1484,N_1429);
nand U1926 (N_1926,N_1574,N_1333);
xor U1927 (N_1927,N_1425,N_1235);
and U1928 (N_1928,N_1587,N_1529);
or U1929 (N_1929,N_1482,N_1483);
and U1930 (N_1930,N_1259,N_1500);
or U1931 (N_1931,N_1542,N_1516);
nand U1932 (N_1932,N_1244,N_1570);
or U1933 (N_1933,N_1457,N_1216);
and U1934 (N_1934,N_1303,N_1295);
and U1935 (N_1935,N_1398,N_1402);
and U1936 (N_1936,N_1412,N_1538);
nand U1937 (N_1937,N_1467,N_1381);
and U1938 (N_1938,N_1582,N_1291);
and U1939 (N_1939,N_1405,N_1563);
nor U1940 (N_1940,N_1363,N_1531);
nand U1941 (N_1941,N_1335,N_1543);
nor U1942 (N_1942,N_1427,N_1367);
and U1943 (N_1943,N_1423,N_1441);
and U1944 (N_1944,N_1219,N_1529);
nand U1945 (N_1945,N_1556,N_1225);
and U1946 (N_1946,N_1597,N_1315);
or U1947 (N_1947,N_1200,N_1392);
nand U1948 (N_1948,N_1515,N_1480);
and U1949 (N_1949,N_1300,N_1529);
and U1950 (N_1950,N_1456,N_1549);
and U1951 (N_1951,N_1314,N_1467);
or U1952 (N_1952,N_1259,N_1553);
or U1953 (N_1953,N_1453,N_1208);
or U1954 (N_1954,N_1531,N_1428);
nor U1955 (N_1955,N_1272,N_1483);
and U1956 (N_1956,N_1281,N_1221);
nor U1957 (N_1957,N_1282,N_1286);
xor U1958 (N_1958,N_1223,N_1489);
and U1959 (N_1959,N_1584,N_1526);
nor U1960 (N_1960,N_1424,N_1430);
nand U1961 (N_1961,N_1347,N_1553);
xor U1962 (N_1962,N_1247,N_1300);
and U1963 (N_1963,N_1487,N_1326);
xor U1964 (N_1964,N_1495,N_1413);
xnor U1965 (N_1965,N_1440,N_1223);
or U1966 (N_1966,N_1285,N_1351);
nand U1967 (N_1967,N_1449,N_1222);
and U1968 (N_1968,N_1485,N_1584);
or U1969 (N_1969,N_1365,N_1535);
nand U1970 (N_1970,N_1263,N_1381);
nor U1971 (N_1971,N_1206,N_1541);
xnor U1972 (N_1972,N_1299,N_1282);
and U1973 (N_1973,N_1319,N_1592);
and U1974 (N_1974,N_1318,N_1457);
and U1975 (N_1975,N_1349,N_1503);
and U1976 (N_1976,N_1247,N_1238);
nand U1977 (N_1977,N_1212,N_1528);
xor U1978 (N_1978,N_1394,N_1320);
nand U1979 (N_1979,N_1356,N_1340);
or U1980 (N_1980,N_1217,N_1349);
nand U1981 (N_1981,N_1503,N_1421);
and U1982 (N_1982,N_1529,N_1463);
or U1983 (N_1983,N_1499,N_1263);
nor U1984 (N_1984,N_1469,N_1234);
or U1985 (N_1985,N_1210,N_1399);
and U1986 (N_1986,N_1487,N_1388);
and U1987 (N_1987,N_1274,N_1480);
and U1988 (N_1988,N_1422,N_1569);
and U1989 (N_1989,N_1359,N_1563);
nand U1990 (N_1990,N_1408,N_1559);
xor U1991 (N_1991,N_1506,N_1326);
nand U1992 (N_1992,N_1445,N_1215);
nand U1993 (N_1993,N_1355,N_1558);
nor U1994 (N_1994,N_1231,N_1539);
nor U1995 (N_1995,N_1396,N_1477);
nand U1996 (N_1996,N_1426,N_1401);
nor U1997 (N_1997,N_1546,N_1354);
and U1998 (N_1998,N_1371,N_1466);
xnor U1999 (N_1999,N_1216,N_1569);
nor U2000 (N_2000,N_1751,N_1763);
and U2001 (N_2001,N_1645,N_1943);
nand U2002 (N_2002,N_1715,N_1723);
or U2003 (N_2003,N_1819,N_1953);
nor U2004 (N_2004,N_1849,N_1777);
nor U2005 (N_2005,N_1899,N_1983);
or U2006 (N_2006,N_1656,N_1750);
or U2007 (N_2007,N_1816,N_1684);
and U2008 (N_2008,N_1629,N_1818);
or U2009 (N_2009,N_1971,N_1725);
nor U2010 (N_2010,N_1604,N_1695);
or U2011 (N_2011,N_1927,N_1804);
and U2012 (N_2012,N_1749,N_1946);
and U2013 (N_2013,N_1958,N_1626);
xnor U2014 (N_2014,N_1766,N_1722);
and U2015 (N_2015,N_1982,N_1720);
or U2016 (N_2016,N_1920,N_1635);
nor U2017 (N_2017,N_1901,N_1637);
or U2018 (N_2018,N_1666,N_1970);
or U2019 (N_2019,N_1788,N_1783);
and U2020 (N_2020,N_1883,N_1906);
and U2021 (N_2021,N_1922,N_1713);
xnor U2022 (N_2022,N_1931,N_1634);
nor U2023 (N_2023,N_1960,N_1984);
and U2024 (N_2024,N_1974,N_1948);
xnor U2025 (N_2025,N_1782,N_1800);
or U2026 (N_2026,N_1916,N_1731);
nor U2027 (N_2027,N_1616,N_1888);
and U2028 (N_2028,N_1892,N_1738);
nand U2029 (N_2029,N_1843,N_1949);
or U2030 (N_2030,N_1900,N_1919);
and U2031 (N_2031,N_1620,N_1600);
nand U2032 (N_2032,N_1808,N_1878);
nor U2033 (N_2033,N_1833,N_1894);
and U2034 (N_2034,N_1654,N_1621);
or U2035 (N_2035,N_1796,N_1996);
xnor U2036 (N_2036,N_1700,N_1703);
nor U2037 (N_2037,N_1865,N_1895);
and U2038 (N_2038,N_1844,N_1602);
and U2039 (N_2039,N_1934,N_1679);
and U2040 (N_2040,N_1658,N_1813);
or U2041 (N_2041,N_1988,N_1893);
xor U2042 (N_2042,N_1753,N_1871);
or U2043 (N_2043,N_1968,N_1966);
xor U2044 (N_2044,N_1824,N_1923);
and U2045 (N_2045,N_1789,N_1936);
nand U2046 (N_2046,N_1908,N_1734);
and U2047 (N_2047,N_1730,N_1611);
or U2048 (N_2048,N_1683,N_1737);
nor U2049 (N_2049,N_1873,N_1719);
or U2050 (N_2050,N_1778,N_1647);
nor U2051 (N_2051,N_1619,N_1850);
or U2052 (N_2052,N_1852,N_1610);
or U2053 (N_2053,N_1907,N_1848);
nor U2054 (N_2054,N_1697,N_1925);
or U2055 (N_2055,N_1628,N_1864);
and U2056 (N_2056,N_1756,N_1685);
xnor U2057 (N_2057,N_1742,N_1969);
nor U2058 (N_2058,N_1680,N_1798);
and U2059 (N_2059,N_1729,N_1625);
xnor U2060 (N_2060,N_1929,N_1841);
or U2061 (N_2061,N_1917,N_1606);
nor U2062 (N_2062,N_1835,N_1912);
and U2063 (N_2063,N_1718,N_1909);
nor U2064 (N_2064,N_1743,N_1976);
or U2065 (N_2065,N_1829,N_1669);
nand U2066 (N_2066,N_1724,N_1866);
and U2067 (N_2067,N_1823,N_1915);
nand U2068 (N_2068,N_1839,N_1882);
xnor U2069 (N_2069,N_1964,N_1664);
or U2070 (N_2070,N_1986,N_1885);
nor U2071 (N_2071,N_1630,N_1999);
xnor U2072 (N_2072,N_1827,N_1608);
nor U2073 (N_2073,N_1639,N_1826);
nand U2074 (N_2074,N_1791,N_1998);
or U2075 (N_2075,N_1710,N_1601);
or U2076 (N_2076,N_1617,N_1614);
nor U2077 (N_2077,N_1972,N_1809);
or U2078 (N_2078,N_1633,N_1855);
nand U2079 (N_2079,N_1667,N_1913);
xor U2080 (N_2080,N_1759,N_1847);
xnor U2081 (N_2081,N_1653,N_1668);
or U2082 (N_2082,N_1784,N_1952);
xnor U2083 (N_2083,N_1631,N_1794);
nor U2084 (N_2084,N_1793,N_1812);
xor U2085 (N_2085,N_1940,N_1705);
nand U2086 (N_2086,N_1959,N_1837);
nand U2087 (N_2087,N_1941,N_1938);
and U2088 (N_2088,N_1762,N_1851);
and U2089 (N_2089,N_1661,N_1771);
nand U2090 (N_2090,N_1930,N_1609);
nand U2091 (N_2091,N_1854,N_1963);
or U2092 (N_2092,N_1859,N_1802);
and U2093 (N_2093,N_1896,N_1613);
and U2094 (N_2094,N_1698,N_1918);
nor U2095 (N_2095,N_1622,N_1775);
and U2096 (N_2096,N_1846,N_1961);
nand U2097 (N_2097,N_1772,N_1799);
xor U2098 (N_2098,N_1757,N_1921);
nor U2099 (N_2099,N_1662,N_1881);
xnor U2100 (N_2100,N_1954,N_1861);
and U2101 (N_2101,N_1735,N_1797);
xor U2102 (N_2102,N_1677,N_1997);
nor U2103 (N_2103,N_1675,N_1744);
xor U2104 (N_2104,N_1732,N_1646);
and U2105 (N_2105,N_1711,N_1615);
xnor U2106 (N_2106,N_1781,N_1678);
nand U2107 (N_2107,N_1761,N_1708);
xnor U2108 (N_2108,N_1696,N_1832);
nor U2109 (N_2109,N_1760,N_1649);
nor U2110 (N_2110,N_1728,N_1694);
and U2111 (N_2111,N_1785,N_1891);
nor U2112 (N_2112,N_1692,N_1754);
xor U2113 (N_2113,N_1636,N_1686);
nor U2114 (N_2114,N_1642,N_1942);
nor U2115 (N_2115,N_1682,N_1935);
or U2116 (N_2116,N_1672,N_1736);
xor U2117 (N_2117,N_1897,N_1657);
and U2118 (N_2118,N_1822,N_1856);
or U2119 (N_2119,N_1955,N_1945);
nand U2120 (N_2120,N_1928,N_1691);
or U2121 (N_2121,N_1877,N_1605);
or U2122 (N_2122,N_1659,N_1701);
xor U2123 (N_2123,N_1950,N_1787);
or U2124 (N_2124,N_1643,N_1932);
xnor U2125 (N_2125,N_1821,N_1977);
xor U2126 (N_2126,N_1801,N_1987);
and U2127 (N_2127,N_1674,N_1681);
nor U2128 (N_2128,N_1741,N_1648);
nor U2129 (N_2129,N_1924,N_1806);
and U2130 (N_2130,N_1830,N_1820);
and U2131 (N_2131,N_1687,N_1870);
or U2132 (N_2132,N_1768,N_1770);
nor U2133 (N_2133,N_1973,N_1879);
and U2134 (N_2134,N_1857,N_1814);
nand U2135 (N_2135,N_1979,N_1811);
and U2136 (N_2136,N_1769,N_1815);
and U2137 (N_2137,N_1962,N_1651);
xnor U2138 (N_2138,N_1624,N_1967);
and U2139 (N_2139,N_1795,N_1790);
nand U2140 (N_2140,N_1780,N_1985);
or U2141 (N_2141,N_1880,N_1714);
nand U2142 (N_2142,N_1956,N_1748);
nand U2143 (N_2143,N_1910,N_1623);
xnor U2144 (N_2144,N_1840,N_1644);
xor U2145 (N_2145,N_1740,N_1774);
and U2146 (N_2146,N_1926,N_1704);
nor U2147 (N_2147,N_1673,N_1957);
and U2148 (N_2148,N_1989,N_1746);
nand U2149 (N_2149,N_1699,N_1779);
and U2150 (N_2150,N_1872,N_1773);
or U2151 (N_2151,N_1805,N_1792);
and U2152 (N_2152,N_1721,N_1853);
and U2153 (N_2153,N_1867,N_1650);
nor U2154 (N_2154,N_1640,N_1810);
and U2155 (N_2155,N_1618,N_1693);
nor U2156 (N_2156,N_1905,N_1887);
nand U2157 (N_2157,N_1862,N_1764);
nor U2158 (N_2158,N_1911,N_1803);
nor U2159 (N_2159,N_1670,N_1706);
nand U2160 (N_2160,N_1876,N_1676);
or U2161 (N_2161,N_1632,N_1875);
and U2162 (N_2162,N_1995,N_1739);
or U2163 (N_2163,N_1991,N_1838);
and U2164 (N_2164,N_1755,N_1939);
or U2165 (N_2165,N_1869,N_1994);
nor U2166 (N_2166,N_1834,N_1655);
nand U2167 (N_2167,N_1980,N_1745);
and U2168 (N_2168,N_1993,N_1904);
nor U2169 (N_2169,N_1671,N_1828);
nand U2170 (N_2170,N_1690,N_1702);
or U2171 (N_2171,N_1652,N_1712);
and U2172 (N_2172,N_1689,N_1975);
nor U2173 (N_2173,N_1688,N_1845);
or U2174 (N_2174,N_1990,N_1914);
and U2175 (N_2175,N_1951,N_1874);
or U2176 (N_2176,N_1902,N_1992);
or U2177 (N_2177,N_1898,N_1858);
and U2178 (N_2178,N_1638,N_1727);
nor U2179 (N_2179,N_1627,N_1903);
nor U2180 (N_2180,N_1884,N_1944);
or U2181 (N_2181,N_1665,N_1660);
and U2182 (N_2182,N_1717,N_1707);
and U2183 (N_2183,N_1786,N_1767);
xor U2184 (N_2184,N_1758,N_1842);
nand U2185 (N_2185,N_1947,N_1825);
nand U2186 (N_2186,N_1937,N_1889);
xor U2187 (N_2187,N_1709,N_1860);
and U2188 (N_2188,N_1978,N_1836);
xor U2189 (N_2189,N_1890,N_1868);
nand U2190 (N_2190,N_1933,N_1965);
xor U2191 (N_2191,N_1716,N_1603);
xor U2192 (N_2192,N_1776,N_1612);
or U2193 (N_2193,N_1641,N_1726);
nor U2194 (N_2194,N_1807,N_1817);
nor U2195 (N_2195,N_1831,N_1863);
or U2196 (N_2196,N_1607,N_1752);
and U2197 (N_2197,N_1747,N_1886);
nand U2198 (N_2198,N_1733,N_1663);
or U2199 (N_2199,N_1981,N_1765);
and U2200 (N_2200,N_1675,N_1890);
and U2201 (N_2201,N_1910,N_1786);
and U2202 (N_2202,N_1710,N_1650);
or U2203 (N_2203,N_1687,N_1798);
and U2204 (N_2204,N_1827,N_1865);
or U2205 (N_2205,N_1730,N_1601);
xnor U2206 (N_2206,N_1834,N_1773);
nand U2207 (N_2207,N_1714,N_1858);
or U2208 (N_2208,N_1733,N_1979);
and U2209 (N_2209,N_1937,N_1771);
xor U2210 (N_2210,N_1619,N_1736);
or U2211 (N_2211,N_1828,N_1672);
nand U2212 (N_2212,N_1724,N_1977);
nand U2213 (N_2213,N_1993,N_1754);
xnor U2214 (N_2214,N_1918,N_1606);
xnor U2215 (N_2215,N_1654,N_1678);
xnor U2216 (N_2216,N_1739,N_1815);
xnor U2217 (N_2217,N_1636,N_1721);
or U2218 (N_2218,N_1605,N_1990);
xnor U2219 (N_2219,N_1646,N_1749);
nand U2220 (N_2220,N_1810,N_1792);
xnor U2221 (N_2221,N_1818,N_1774);
nor U2222 (N_2222,N_1722,N_1742);
nor U2223 (N_2223,N_1768,N_1713);
xnor U2224 (N_2224,N_1742,N_1950);
and U2225 (N_2225,N_1870,N_1988);
xnor U2226 (N_2226,N_1940,N_1811);
or U2227 (N_2227,N_1704,N_1844);
or U2228 (N_2228,N_1669,N_1653);
xnor U2229 (N_2229,N_1934,N_1622);
nand U2230 (N_2230,N_1872,N_1927);
nand U2231 (N_2231,N_1786,N_1707);
and U2232 (N_2232,N_1857,N_1621);
and U2233 (N_2233,N_1996,N_1716);
or U2234 (N_2234,N_1668,N_1775);
nor U2235 (N_2235,N_1631,N_1686);
or U2236 (N_2236,N_1664,N_1635);
nand U2237 (N_2237,N_1654,N_1663);
or U2238 (N_2238,N_1905,N_1953);
nor U2239 (N_2239,N_1993,N_1799);
nand U2240 (N_2240,N_1928,N_1824);
nor U2241 (N_2241,N_1667,N_1702);
nand U2242 (N_2242,N_1866,N_1607);
and U2243 (N_2243,N_1662,N_1740);
nand U2244 (N_2244,N_1906,N_1668);
nor U2245 (N_2245,N_1704,N_1947);
or U2246 (N_2246,N_1959,N_1988);
nand U2247 (N_2247,N_1680,N_1695);
or U2248 (N_2248,N_1679,N_1681);
nand U2249 (N_2249,N_1725,N_1980);
xnor U2250 (N_2250,N_1704,N_1974);
xor U2251 (N_2251,N_1975,N_1794);
and U2252 (N_2252,N_1732,N_1867);
or U2253 (N_2253,N_1819,N_1672);
nor U2254 (N_2254,N_1630,N_1655);
xor U2255 (N_2255,N_1662,N_1840);
nor U2256 (N_2256,N_1694,N_1789);
or U2257 (N_2257,N_1647,N_1688);
and U2258 (N_2258,N_1999,N_1796);
or U2259 (N_2259,N_1980,N_1675);
nand U2260 (N_2260,N_1965,N_1905);
and U2261 (N_2261,N_1600,N_1679);
nor U2262 (N_2262,N_1890,N_1709);
nor U2263 (N_2263,N_1903,N_1958);
xnor U2264 (N_2264,N_1781,N_1855);
nand U2265 (N_2265,N_1661,N_1821);
nor U2266 (N_2266,N_1816,N_1820);
xor U2267 (N_2267,N_1666,N_1852);
and U2268 (N_2268,N_1768,N_1722);
xor U2269 (N_2269,N_1621,N_1668);
and U2270 (N_2270,N_1927,N_1870);
or U2271 (N_2271,N_1679,N_1626);
nand U2272 (N_2272,N_1861,N_1695);
xnor U2273 (N_2273,N_1876,N_1661);
or U2274 (N_2274,N_1681,N_1630);
and U2275 (N_2275,N_1867,N_1887);
nand U2276 (N_2276,N_1907,N_1674);
nor U2277 (N_2277,N_1760,N_1782);
or U2278 (N_2278,N_1883,N_1848);
nor U2279 (N_2279,N_1919,N_1631);
nand U2280 (N_2280,N_1837,N_1768);
and U2281 (N_2281,N_1920,N_1742);
and U2282 (N_2282,N_1995,N_1917);
or U2283 (N_2283,N_1961,N_1912);
nor U2284 (N_2284,N_1633,N_1940);
nand U2285 (N_2285,N_1720,N_1818);
and U2286 (N_2286,N_1699,N_1909);
and U2287 (N_2287,N_1611,N_1909);
nand U2288 (N_2288,N_1776,N_1710);
or U2289 (N_2289,N_1651,N_1609);
nand U2290 (N_2290,N_1926,N_1874);
or U2291 (N_2291,N_1942,N_1794);
and U2292 (N_2292,N_1725,N_1601);
or U2293 (N_2293,N_1657,N_1705);
and U2294 (N_2294,N_1954,N_1851);
xor U2295 (N_2295,N_1633,N_1945);
nand U2296 (N_2296,N_1603,N_1959);
xor U2297 (N_2297,N_1735,N_1617);
or U2298 (N_2298,N_1710,N_1999);
nand U2299 (N_2299,N_1926,N_1789);
nand U2300 (N_2300,N_1776,N_1994);
and U2301 (N_2301,N_1995,N_1949);
xor U2302 (N_2302,N_1822,N_1716);
nand U2303 (N_2303,N_1850,N_1617);
xnor U2304 (N_2304,N_1797,N_1862);
nor U2305 (N_2305,N_1653,N_1811);
nand U2306 (N_2306,N_1694,N_1768);
nand U2307 (N_2307,N_1649,N_1725);
and U2308 (N_2308,N_1813,N_1761);
nor U2309 (N_2309,N_1610,N_1913);
or U2310 (N_2310,N_1789,N_1723);
and U2311 (N_2311,N_1618,N_1754);
or U2312 (N_2312,N_1999,N_1633);
nand U2313 (N_2313,N_1766,N_1946);
xor U2314 (N_2314,N_1899,N_1650);
nand U2315 (N_2315,N_1847,N_1838);
nor U2316 (N_2316,N_1612,N_1722);
nand U2317 (N_2317,N_1711,N_1827);
nor U2318 (N_2318,N_1948,N_1954);
nor U2319 (N_2319,N_1731,N_1834);
nor U2320 (N_2320,N_1743,N_1974);
or U2321 (N_2321,N_1818,N_1638);
nand U2322 (N_2322,N_1689,N_1967);
or U2323 (N_2323,N_1630,N_1629);
nand U2324 (N_2324,N_1970,N_1691);
nor U2325 (N_2325,N_1777,N_1808);
xor U2326 (N_2326,N_1944,N_1693);
nor U2327 (N_2327,N_1699,N_1880);
and U2328 (N_2328,N_1961,N_1904);
and U2329 (N_2329,N_1706,N_1765);
or U2330 (N_2330,N_1665,N_1808);
and U2331 (N_2331,N_1837,N_1809);
or U2332 (N_2332,N_1619,N_1680);
xor U2333 (N_2333,N_1715,N_1858);
and U2334 (N_2334,N_1873,N_1838);
xnor U2335 (N_2335,N_1718,N_1706);
nor U2336 (N_2336,N_1735,N_1968);
xnor U2337 (N_2337,N_1710,N_1797);
nor U2338 (N_2338,N_1840,N_1981);
nand U2339 (N_2339,N_1715,N_1770);
nand U2340 (N_2340,N_1938,N_1978);
or U2341 (N_2341,N_1681,N_1752);
xnor U2342 (N_2342,N_1858,N_1679);
nor U2343 (N_2343,N_1835,N_1727);
or U2344 (N_2344,N_1917,N_1971);
or U2345 (N_2345,N_1929,N_1824);
xnor U2346 (N_2346,N_1732,N_1665);
nor U2347 (N_2347,N_1845,N_1723);
or U2348 (N_2348,N_1946,N_1725);
nor U2349 (N_2349,N_1952,N_1768);
or U2350 (N_2350,N_1863,N_1754);
and U2351 (N_2351,N_1984,N_1726);
and U2352 (N_2352,N_1951,N_1829);
nor U2353 (N_2353,N_1949,N_1688);
nor U2354 (N_2354,N_1769,N_1729);
nand U2355 (N_2355,N_1755,N_1891);
or U2356 (N_2356,N_1951,N_1863);
nand U2357 (N_2357,N_1885,N_1642);
xnor U2358 (N_2358,N_1682,N_1891);
nand U2359 (N_2359,N_1782,N_1892);
and U2360 (N_2360,N_1625,N_1923);
or U2361 (N_2361,N_1793,N_1982);
and U2362 (N_2362,N_1723,N_1675);
and U2363 (N_2363,N_1865,N_1631);
or U2364 (N_2364,N_1861,N_1694);
or U2365 (N_2365,N_1631,N_1601);
nand U2366 (N_2366,N_1789,N_1893);
nand U2367 (N_2367,N_1970,N_1796);
xnor U2368 (N_2368,N_1678,N_1979);
xnor U2369 (N_2369,N_1705,N_1813);
or U2370 (N_2370,N_1813,N_1898);
nor U2371 (N_2371,N_1654,N_1634);
nand U2372 (N_2372,N_1712,N_1762);
xor U2373 (N_2373,N_1693,N_1884);
nand U2374 (N_2374,N_1660,N_1890);
xnor U2375 (N_2375,N_1702,N_1762);
xor U2376 (N_2376,N_1646,N_1980);
or U2377 (N_2377,N_1978,N_1800);
nand U2378 (N_2378,N_1868,N_1682);
nor U2379 (N_2379,N_1898,N_1618);
and U2380 (N_2380,N_1875,N_1697);
or U2381 (N_2381,N_1804,N_1753);
nor U2382 (N_2382,N_1622,N_1873);
nor U2383 (N_2383,N_1778,N_1785);
nand U2384 (N_2384,N_1929,N_1840);
nand U2385 (N_2385,N_1953,N_1758);
xor U2386 (N_2386,N_1738,N_1743);
and U2387 (N_2387,N_1905,N_1683);
xnor U2388 (N_2388,N_1920,N_1938);
nand U2389 (N_2389,N_1669,N_1955);
or U2390 (N_2390,N_1819,N_1857);
and U2391 (N_2391,N_1758,N_1666);
nor U2392 (N_2392,N_1779,N_1617);
or U2393 (N_2393,N_1924,N_1837);
nor U2394 (N_2394,N_1754,N_1868);
nand U2395 (N_2395,N_1923,N_1604);
xnor U2396 (N_2396,N_1733,N_1705);
or U2397 (N_2397,N_1733,N_1737);
xor U2398 (N_2398,N_1648,N_1830);
xor U2399 (N_2399,N_1957,N_1725);
nor U2400 (N_2400,N_2228,N_2172);
nand U2401 (N_2401,N_2353,N_2116);
and U2402 (N_2402,N_2373,N_2173);
nand U2403 (N_2403,N_2183,N_2186);
and U2404 (N_2404,N_2166,N_2355);
and U2405 (N_2405,N_2298,N_2255);
and U2406 (N_2406,N_2094,N_2220);
or U2407 (N_2407,N_2231,N_2117);
nand U2408 (N_2408,N_2306,N_2253);
nand U2409 (N_2409,N_2293,N_2018);
nand U2410 (N_2410,N_2140,N_2049);
nand U2411 (N_2411,N_2098,N_2167);
nand U2412 (N_2412,N_2267,N_2144);
and U2413 (N_2413,N_2350,N_2346);
xnor U2414 (N_2414,N_2130,N_2110);
nor U2415 (N_2415,N_2129,N_2349);
nand U2416 (N_2416,N_2342,N_2075);
xor U2417 (N_2417,N_2261,N_2056);
and U2418 (N_2418,N_2204,N_2371);
and U2419 (N_2419,N_2326,N_2364);
nor U2420 (N_2420,N_2099,N_2313);
nor U2421 (N_2421,N_2283,N_2196);
nor U2422 (N_2422,N_2202,N_2107);
and U2423 (N_2423,N_2042,N_2188);
or U2424 (N_2424,N_2125,N_2078);
nor U2425 (N_2425,N_2237,N_2064);
nand U2426 (N_2426,N_2041,N_2341);
nor U2427 (N_2427,N_2048,N_2126);
nand U2428 (N_2428,N_2396,N_2077);
and U2429 (N_2429,N_2068,N_2052);
nor U2430 (N_2430,N_2138,N_2055);
and U2431 (N_2431,N_2258,N_2175);
xor U2432 (N_2432,N_2023,N_2147);
nor U2433 (N_2433,N_2180,N_2376);
xor U2434 (N_2434,N_2359,N_2074);
or U2435 (N_2435,N_2395,N_2235);
nor U2436 (N_2436,N_2277,N_2141);
xnor U2437 (N_2437,N_2007,N_2020);
and U2438 (N_2438,N_2135,N_2027);
nand U2439 (N_2439,N_2134,N_2039);
nand U2440 (N_2440,N_2012,N_2321);
nor U2441 (N_2441,N_2272,N_2248);
nand U2442 (N_2442,N_2081,N_2307);
or U2443 (N_2443,N_2016,N_2392);
nand U2444 (N_2444,N_2150,N_2352);
and U2445 (N_2445,N_2105,N_2004);
and U2446 (N_2446,N_2148,N_2165);
xnor U2447 (N_2447,N_2066,N_2192);
nand U2448 (N_2448,N_2067,N_2312);
or U2449 (N_2449,N_2205,N_2224);
xnor U2450 (N_2450,N_2076,N_2325);
and U2451 (N_2451,N_2089,N_2333);
xor U2452 (N_2452,N_2337,N_2367);
nor U2453 (N_2453,N_2209,N_2361);
and U2454 (N_2454,N_2332,N_2390);
or U2455 (N_2455,N_2344,N_2327);
nor U2456 (N_2456,N_2374,N_2185);
nor U2457 (N_2457,N_2318,N_2245);
nor U2458 (N_2458,N_2159,N_2300);
or U2459 (N_2459,N_2137,N_2046);
and U2460 (N_2460,N_2132,N_2299);
and U2461 (N_2461,N_2028,N_2029);
nand U2462 (N_2462,N_2288,N_2223);
nor U2463 (N_2463,N_2314,N_2154);
nand U2464 (N_2464,N_2030,N_2351);
nand U2465 (N_2465,N_2254,N_2365);
nor U2466 (N_2466,N_2357,N_2251);
nand U2467 (N_2467,N_2241,N_2274);
and U2468 (N_2468,N_2397,N_2112);
and U2469 (N_2469,N_2229,N_2315);
xor U2470 (N_2470,N_2309,N_2133);
nand U2471 (N_2471,N_2026,N_2244);
xnor U2472 (N_2472,N_2174,N_2399);
and U2473 (N_2473,N_2247,N_2317);
and U2474 (N_2474,N_2304,N_2014);
nor U2475 (N_2475,N_2273,N_2032);
and U2476 (N_2476,N_2388,N_2389);
nor U2477 (N_2477,N_2122,N_2065);
and U2478 (N_2478,N_2363,N_2264);
xor U2479 (N_2479,N_2050,N_2003);
and U2480 (N_2480,N_2006,N_2128);
nand U2481 (N_2481,N_2013,N_2262);
and U2482 (N_2482,N_2278,N_2250);
nand U2483 (N_2483,N_2193,N_2215);
nor U2484 (N_2484,N_2249,N_2214);
nor U2485 (N_2485,N_2294,N_2222);
xnor U2486 (N_2486,N_2208,N_2162);
nand U2487 (N_2487,N_2015,N_2260);
or U2488 (N_2488,N_2211,N_2054);
nor U2489 (N_2489,N_2370,N_2292);
nor U2490 (N_2490,N_2009,N_2354);
and U2491 (N_2491,N_2275,N_2384);
or U2492 (N_2492,N_2328,N_2201);
or U2493 (N_2493,N_2316,N_2178);
xor U2494 (N_2494,N_2221,N_2071);
nor U2495 (N_2495,N_2335,N_2008);
and U2496 (N_2496,N_2149,N_2330);
nand U2497 (N_2497,N_2286,N_2198);
or U2498 (N_2498,N_2120,N_2219);
nor U2499 (N_2499,N_2197,N_2019);
or U2500 (N_2500,N_2142,N_2391);
and U2501 (N_2501,N_2072,N_2297);
nand U2502 (N_2502,N_2143,N_2232);
or U2503 (N_2503,N_2024,N_2338);
nand U2504 (N_2504,N_2000,N_2002);
or U2505 (N_2505,N_2043,N_2060);
xor U2506 (N_2506,N_2303,N_2073);
nor U2507 (N_2507,N_2001,N_2179);
nor U2508 (N_2508,N_2136,N_2123);
or U2509 (N_2509,N_2227,N_2115);
and U2510 (N_2510,N_2263,N_2119);
or U2511 (N_2511,N_2069,N_2289);
nand U2512 (N_2512,N_2238,N_2281);
xor U2513 (N_2513,N_2156,N_2284);
nand U2514 (N_2514,N_2190,N_2102);
xnor U2515 (N_2515,N_2182,N_2127);
xor U2516 (N_2516,N_2111,N_2213);
nand U2517 (N_2517,N_2096,N_2230);
and U2518 (N_2518,N_2381,N_2097);
nor U2519 (N_2519,N_2114,N_2170);
or U2520 (N_2520,N_2093,N_2017);
nor U2521 (N_2521,N_2080,N_2084);
or U2522 (N_2522,N_2011,N_2109);
nor U2523 (N_2523,N_2339,N_2082);
or U2524 (N_2524,N_2362,N_2319);
and U2525 (N_2525,N_2199,N_2394);
or U2526 (N_2526,N_2378,N_2021);
and U2527 (N_2527,N_2287,N_2160);
and U2528 (N_2528,N_2031,N_2345);
and U2529 (N_2529,N_2091,N_2369);
xor U2530 (N_2530,N_2379,N_2187);
or U2531 (N_2531,N_2225,N_2380);
and U2532 (N_2532,N_2265,N_2295);
xnor U2533 (N_2533,N_2377,N_2051);
and U2534 (N_2534,N_2386,N_2106);
or U2535 (N_2535,N_2382,N_2062);
nand U2536 (N_2536,N_2200,N_2372);
xor U2537 (N_2537,N_2393,N_2088);
and U2538 (N_2538,N_2025,N_2216);
xnor U2539 (N_2539,N_2087,N_2311);
nor U2540 (N_2540,N_2324,N_2385);
xor U2541 (N_2541,N_2058,N_2259);
nand U2542 (N_2542,N_2045,N_2206);
xor U2543 (N_2543,N_2336,N_2282);
or U2544 (N_2544,N_2005,N_2184);
nand U2545 (N_2545,N_2217,N_2358);
nand U2546 (N_2546,N_2153,N_2189);
nand U2547 (N_2547,N_2171,N_2104);
nor U2548 (N_2548,N_2079,N_2366);
nor U2549 (N_2549,N_2124,N_2296);
nor U2550 (N_2550,N_2177,N_2063);
xor U2551 (N_2551,N_2269,N_2329);
nor U2552 (N_2552,N_2279,N_2101);
and U2553 (N_2553,N_2323,N_2083);
nor U2554 (N_2554,N_2038,N_2322);
or U2555 (N_2555,N_2092,N_2059);
nand U2556 (N_2556,N_2061,N_2398);
and U2557 (N_2557,N_2085,N_2161);
xnor U2558 (N_2558,N_2191,N_2383);
xor U2559 (N_2559,N_2203,N_2040);
nand U2560 (N_2560,N_2164,N_2151);
nor U2561 (N_2561,N_2139,N_2207);
nor U2562 (N_2562,N_2010,N_2103);
nand U2563 (N_2563,N_2118,N_2131);
xor U2564 (N_2564,N_2152,N_2256);
and U2565 (N_2565,N_2053,N_2280);
nand U2566 (N_2566,N_2158,N_2121);
and U2567 (N_2567,N_2157,N_2168);
and U2568 (N_2568,N_2195,N_2194);
nand U2569 (N_2569,N_2348,N_2302);
and U2570 (N_2570,N_2305,N_2022);
nand U2571 (N_2571,N_2033,N_2240);
or U2572 (N_2572,N_2090,N_2290);
or U2573 (N_2573,N_2047,N_2239);
or U2574 (N_2574,N_2252,N_2113);
and U2575 (N_2575,N_2236,N_2095);
xor U2576 (N_2576,N_2176,N_2181);
xor U2577 (N_2577,N_2086,N_2268);
or U2578 (N_2578,N_2034,N_2057);
xnor U2579 (N_2579,N_2035,N_2340);
xnor U2580 (N_2580,N_2270,N_2285);
xnor U2581 (N_2581,N_2308,N_2037);
or U2582 (N_2582,N_2070,N_2387);
nor U2583 (N_2583,N_2276,N_2331);
xor U2584 (N_2584,N_2155,N_2246);
nor U2585 (N_2585,N_2347,N_2044);
nor U2586 (N_2586,N_2212,N_2036);
xnor U2587 (N_2587,N_2145,N_2226);
and U2588 (N_2588,N_2169,N_2375);
xor U2589 (N_2589,N_2266,N_2243);
or U2590 (N_2590,N_2360,N_2100);
and U2591 (N_2591,N_2356,N_2234);
xor U2592 (N_2592,N_2368,N_2271);
or U2593 (N_2593,N_2320,N_2334);
nor U2594 (N_2594,N_2146,N_2291);
nand U2595 (N_2595,N_2257,N_2108);
nand U2596 (N_2596,N_2218,N_2301);
or U2597 (N_2597,N_2210,N_2343);
and U2598 (N_2598,N_2310,N_2242);
and U2599 (N_2599,N_2233,N_2163);
xnor U2600 (N_2600,N_2199,N_2250);
and U2601 (N_2601,N_2141,N_2375);
nand U2602 (N_2602,N_2328,N_2232);
and U2603 (N_2603,N_2394,N_2193);
nand U2604 (N_2604,N_2228,N_2305);
and U2605 (N_2605,N_2112,N_2286);
or U2606 (N_2606,N_2081,N_2123);
and U2607 (N_2607,N_2114,N_2010);
and U2608 (N_2608,N_2261,N_2300);
or U2609 (N_2609,N_2086,N_2199);
xnor U2610 (N_2610,N_2290,N_2175);
nor U2611 (N_2611,N_2139,N_2104);
nand U2612 (N_2612,N_2142,N_2066);
xor U2613 (N_2613,N_2221,N_2189);
xor U2614 (N_2614,N_2046,N_2146);
xor U2615 (N_2615,N_2240,N_2037);
or U2616 (N_2616,N_2035,N_2233);
nor U2617 (N_2617,N_2155,N_2267);
and U2618 (N_2618,N_2361,N_2248);
and U2619 (N_2619,N_2196,N_2103);
and U2620 (N_2620,N_2247,N_2170);
and U2621 (N_2621,N_2049,N_2010);
xnor U2622 (N_2622,N_2002,N_2137);
and U2623 (N_2623,N_2342,N_2112);
xor U2624 (N_2624,N_2245,N_2360);
nand U2625 (N_2625,N_2245,N_2230);
nor U2626 (N_2626,N_2195,N_2358);
nor U2627 (N_2627,N_2069,N_2103);
xor U2628 (N_2628,N_2228,N_2396);
or U2629 (N_2629,N_2148,N_2344);
or U2630 (N_2630,N_2250,N_2249);
or U2631 (N_2631,N_2352,N_2060);
xnor U2632 (N_2632,N_2044,N_2344);
and U2633 (N_2633,N_2381,N_2397);
or U2634 (N_2634,N_2085,N_2291);
xor U2635 (N_2635,N_2205,N_2101);
and U2636 (N_2636,N_2057,N_2059);
or U2637 (N_2637,N_2081,N_2108);
xnor U2638 (N_2638,N_2104,N_2065);
or U2639 (N_2639,N_2084,N_2271);
or U2640 (N_2640,N_2063,N_2119);
nor U2641 (N_2641,N_2112,N_2014);
nand U2642 (N_2642,N_2295,N_2082);
or U2643 (N_2643,N_2233,N_2376);
xnor U2644 (N_2644,N_2163,N_2057);
nor U2645 (N_2645,N_2068,N_2323);
nand U2646 (N_2646,N_2335,N_2254);
nand U2647 (N_2647,N_2250,N_2369);
and U2648 (N_2648,N_2225,N_2106);
xnor U2649 (N_2649,N_2004,N_2289);
and U2650 (N_2650,N_2235,N_2012);
or U2651 (N_2651,N_2326,N_2395);
or U2652 (N_2652,N_2365,N_2361);
and U2653 (N_2653,N_2286,N_2248);
and U2654 (N_2654,N_2080,N_2192);
nand U2655 (N_2655,N_2210,N_2156);
and U2656 (N_2656,N_2218,N_2110);
xnor U2657 (N_2657,N_2365,N_2065);
nand U2658 (N_2658,N_2315,N_2123);
nor U2659 (N_2659,N_2320,N_2111);
nand U2660 (N_2660,N_2347,N_2312);
xnor U2661 (N_2661,N_2238,N_2179);
and U2662 (N_2662,N_2236,N_2063);
or U2663 (N_2663,N_2063,N_2137);
nand U2664 (N_2664,N_2229,N_2294);
xnor U2665 (N_2665,N_2063,N_2317);
nor U2666 (N_2666,N_2235,N_2377);
nor U2667 (N_2667,N_2014,N_2381);
nand U2668 (N_2668,N_2096,N_2393);
or U2669 (N_2669,N_2041,N_2376);
nand U2670 (N_2670,N_2137,N_2012);
nor U2671 (N_2671,N_2077,N_2104);
and U2672 (N_2672,N_2399,N_2389);
and U2673 (N_2673,N_2190,N_2301);
or U2674 (N_2674,N_2287,N_2149);
nand U2675 (N_2675,N_2198,N_2214);
xor U2676 (N_2676,N_2324,N_2105);
nand U2677 (N_2677,N_2021,N_2215);
nand U2678 (N_2678,N_2139,N_2222);
or U2679 (N_2679,N_2233,N_2155);
and U2680 (N_2680,N_2127,N_2282);
nand U2681 (N_2681,N_2177,N_2054);
and U2682 (N_2682,N_2011,N_2075);
or U2683 (N_2683,N_2002,N_2100);
xnor U2684 (N_2684,N_2228,N_2104);
or U2685 (N_2685,N_2208,N_2354);
and U2686 (N_2686,N_2244,N_2115);
and U2687 (N_2687,N_2387,N_2093);
xnor U2688 (N_2688,N_2172,N_2286);
xnor U2689 (N_2689,N_2288,N_2172);
and U2690 (N_2690,N_2071,N_2394);
nand U2691 (N_2691,N_2379,N_2352);
nand U2692 (N_2692,N_2153,N_2216);
nand U2693 (N_2693,N_2134,N_2260);
and U2694 (N_2694,N_2186,N_2120);
or U2695 (N_2695,N_2057,N_2070);
nor U2696 (N_2696,N_2128,N_2290);
and U2697 (N_2697,N_2131,N_2009);
nand U2698 (N_2698,N_2006,N_2182);
nand U2699 (N_2699,N_2320,N_2344);
nor U2700 (N_2700,N_2032,N_2084);
xnor U2701 (N_2701,N_2384,N_2383);
xnor U2702 (N_2702,N_2271,N_2292);
nor U2703 (N_2703,N_2311,N_2359);
xor U2704 (N_2704,N_2364,N_2024);
nand U2705 (N_2705,N_2062,N_2180);
or U2706 (N_2706,N_2171,N_2186);
and U2707 (N_2707,N_2261,N_2061);
nor U2708 (N_2708,N_2287,N_2305);
nand U2709 (N_2709,N_2399,N_2108);
xor U2710 (N_2710,N_2162,N_2050);
and U2711 (N_2711,N_2138,N_2068);
or U2712 (N_2712,N_2220,N_2207);
and U2713 (N_2713,N_2113,N_2357);
or U2714 (N_2714,N_2117,N_2380);
nand U2715 (N_2715,N_2258,N_2139);
or U2716 (N_2716,N_2188,N_2363);
nor U2717 (N_2717,N_2387,N_2202);
nand U2718 (N_2718,N_2164,N_2077);
or U2719 (N_2719,N_2017,N_2027);
xnor U2720 (N_2720,N_2277,N_2212);
nor U2721 (N_2721,N_2290,N_2181);
xor U2722 (N_2722,N_2148,N_2321);
or U2723 (N_2723,N_2070,N_2288);
nand U2724 (N_2724,N_2161,N_2310);
and U2725 (N_2725,N_2356,N_2129);
and U2726 (N_2726,N_2149,N_2140);
or U2727 (N_2727,N_2185,N_2273);
and U2728 (N_2728,N_2176,N_2018);
or U2729 (N_2729,N_2034,N_2209);
xnor U2730 (N_2730,N_2188,N_2270);
or U2731 (N_2731,N_2146,N_2274);
or U2732 (N_2732,N_2024,N_2280);
nor U2733 (N_2733,N_2000,N_2055);
xnor U2734 (N_2734,N_2309,N_2375);
xnor U2735 (N_2735,N_2179,N_2346);
xnor U2736 (N_2736,N_2126,N_2365);
nor U2737 (N_2737,N_2019,N_2290);
nand U2738 (N_2738,N_2290,N_2369);
nand U2739 (N_2739,N_2068,N_2027);
or U2740 (N_2740,N_2114,N_2133);
xor U2741 (N_2741,N_2148,N_2348);
nor U2742 (N_2742,N_2322,N_2113);
nand U2743 (N_2743,N_2345,N_2395);
or U2744 (N_2744,N_2351,N_2210);
and U2745 (N_2745,N_2347,N_2236);
or U2746 (N_2746,N_2018,N_2374);
nand U2747 (N_2747,N_2379,N_2285);
or U2748 (N_2748,N_2305,N_2037);
nand U2749 (N_2749,N_2285,N_2001);
or U2750 (N_2750,N_2036,N_2063);
nor U2751 (N_2751,N_2364,N_2167);
and U2752 (N_2752,N_2304,N_2276);
or U2753 (N_2753,N_2209,N_2370);
nor U2754 (N_2754,N_2035,N_2244);
nor U2755 (N_2755,N_2037,N_2307);
or U2756 (N_2756,N_2156,N_2126);
nor U2757 (N_2757,N_2358,N_2314);
or U2758 (N_2758,N_2159,N_2072);
and U2759 (N_2759,N_2195,N_2341);
nand U2760 (N_2760,N_2378,N_2220);
nor U2761 (N_2761,N_2084,N_2152);
and U2762 (N_2762,N_2165,N_2336);
and U2763 (N_2763,N_2164,N_2248);
or U2764 (N_2764,N_2309,N_2395);
nor U2765 (N_2765,N_2013,N_2071);
nand U2766 (N_2766,N_2326,N_2045);
nor U2767 (N_2767,N_2379,N_2325);
xnor U2768 (N_2768,N_2168,N_2000);
and U2769 (N_2769,N_2068,N_2097);
nand U2770 (N_2770,N_2012,N_2002);
nand U2771 (N_2771,N_2365,N_2232);
nand U2772 (N_2772,N_2301,N_2300);
and U2773 (N_2773,N_2018,N_2271);
or U2774 (N_2774,N_2081,N_2268);
or U2775 (N_2775,N_2301,N_2109);
xnor U2776 (N_2776,N_2232,N_2392);
nor U2777 (N_2777,N_2205,N_2052);
xnor U2778 (N_2778,N_2019,N_2051);
nor U2779 (N_2779,N_2202,N_2006);
xor U2780 (N_2780,N_2383,N_2019);
and U2781 (N_2781,N_2360,N_2378);
nand U2782 (N_2782,N_2125,N_2209);
nand U2783 (N_2783,N_2124,N_2334);
and U2784 (N_2784,N_2036,N_2055);
xor U2785 (N_2785,N_2282,N_2152);
nor U2786 (N_2786,N_2202,N_2119);
nand U2787 (N_2787,N_2351,N_2393);
xor U2788 (N_2788,N_2063,N_2318);
nor U2789 (N_2789,N_2013,N_2391);
or U2790 (N_2790,N_2310,N_2295);
nor U2791 (N_2791,N_2375,N_2156);
nand U2792 (N_2792,N_2271,N_2031);
nand U2793 (N_2793,N_2017,N_2135);
nand U2794 (N_2794,N_2248,N_2053);
nor U2795 (N_2795,N_2125,N_2192);
and U2796 (N_2796,N_2173,N_2384);
xnor U2797 (N_2797,N_2307,N_2156);
and U2798 (N_2798,N_2239,N_2354);
nor U2799 (N_2799,N_2068,N_2195);
xnor U2800 (N_2800,N_2631,N_2685);
nor U2801 (N_2801,N_2498,N_2656);
or U2802 (N_2802,N_2493,N_2652);
xor U2803 (N_2803,N_2437,N_2604);
xnor U2804 (N_2804,N_2785,N_2695);
xor U2805 (N_2805,N_2647,N_2427);
and U2806 (N_2806,N_2566,N_2738);
and U2807 (N_2807,N_2629,N_2408);
xor U2808 (N_2808,N_2414,N_2771);
xnor U2809 (N_2809,N_2732,N_2735);
xor U2810 (N_2810,N_2672,N_2727);
nand U2811 (N_2811,N_2488,N_2748);
nor U2812 (N_2812,N_2524,N_2676);
xor U2813 (N_2813,N_2556,N_2564);
or U2814 (N_2814,N_2623,N_2578);
or U2815 (N_2815,N_2753,N_2570);
nand U2816 (N_2816,N_2492,N_2412);
nor U2817 (N_2817,N_2441,N_2581);
and U2818 (N_2818,N_2466,N_2479);
or U2819 (N_2819,N_2596,N_2743);
xor U2820 (N_2820,N_2526,N_2595);
or U2821 (N_2821,N_2529,N_2590);
nor U2822 (N_2822,N_2776,N_2558);
nor U2823 (N_2823,N_2575,N_2605);
nor U2824 (N_2824,N_2431,N_2470);
nor U2825 (N_2825,N_2423,N_2523);
xor U2826 (N_2826,N_2615,N_2713);
or U2827 (N_2827,N_2537,N_2467);
or U2828 (N_2828,N_2769,N_2602);
xnor U2829 (N_2829,N_2746,N_2588);
and U2830 (N_2830,N_2795,N_2658);
or U2831 (N_2831,N_2799,N_2480);
or U2832 (N_2832,N_2786,N_2601);
xnor U2833 (N_2833,N_2563,N_2626);
and U2834 (N_2834,N_2597,N_2778);
or U2835 (N_2835,N_2677,N_2574);
xor U2836 (N_2836,N_2517,N_2620);
or U2837 (N_2837,N_2679,N_2712);
nor U2838 (N_2838,N_2411,N_2593);
or U2839 (N_2839,N_2547,N_2793);
nor U2840 (N_2840,N_2477,N_2619);
and U2841 (N_2841,N_2757,N_2459);
xor U2842 (N_2842,N_2462,N_2444);
nor U2843 (N_2843,N_2717,N_2664);
or U2844 (N_2844,N_2552,N_2463);
and U2845 (N_2845,N_2518,N_2538);
nor U2846 (N_2846,N_2555,N_2476);
nor U2847 (N_2847,N_2663,N_2460);
xnor U2848 (N_2848,N_2644,N_2469);
xnor U2849 (N_2849,N_2650,N_2780);
nor U2850 (N_2850,N_2797,N_2550);
nor U2851 (N_2851,N_2648,N_2655);
nor U2852 (N_2852,N_2584,N_2420);
xnor U2853 (N_2853,N_2554,N_2693);
nor U2854 (N_2854,N_2544,N_2495);
nor U2855 (N_2855,N_2768,N_2534);
and U2856 (N_2856,N_2761,N_2627);
xor U2857 (N_2857,N_2490,N_2452);
nand U2858 (N_2858,N_2752,N_2637);
or U2859 (N_2859,N_2458,N_2659);
nand U2860 (N_2860,N_2592,N_2763);
nor U2861 (N_2861,N_2496,N_2416);
nor U2862 (N_2862,N_2697,N_2454);
nor U2863 (N_2863,N_2511,N_2422);
and U2864 (N_2864,N_2440,N_2722);
and U2865 (N_2865,N_2653,N_2424);
xnor U2866 (N_2866,N_2600,N_2704);
nand U2867 (N_2867,N_2724,N_2583);
or U2868 (N_2868,N_2673,N_2782);
and U2869 (N_2869,N_2413,N_2791);
or U2870 (N_2870,N_2636,N_2472);
and U2871 (N_2871,N_2594,N_2429);
and U2872 (N_2872,N_2543,N_2505);
or U2873 (N_2873,N_2435,N_2551);
nor U2874 (N_2874,N_2450,N_2669);
and U2875 (N_2875,N_2775,N_2489);
or U2876 (N_2876,N_2535,N_2606);
nor U2877 (N_2877,N_2611,N_2609);
nand U2878 (N_2878,N_2504,N_2750);
and U2879 (N_2879,N_2443,N_2661);
or U2880 (N_2880,N_2789,N_2643);
nand U2881 (N_2881,N_2610,N_2635);
nor U2882 (N_2882,N_2709,N_2579);
xnor U2883 (N_2883,N_2740,N_2639);
xor U2884 (N_2884,N_2688,N_2777);
nand U2885 (N_2885,N_2720,N_2794);
and U2886 (N_2886,N_2621,N_2508);
and U2887 (N_2887,N_2756,N_2739);
or U2888 (N_2888,N_2560,N_2665);
or U2889 (N_2889,N_2478,N_2773);
nand U2890 (N_2890,N_2759,N_2487);
xnor U2891 (N_2891,N_2457,N_2783);
and U2892 (N_2892,N_2533,N_2714);
xnor U2893 (N_2893,N_2501,N_2696);
nand U2894 (N_2894,N_2521,N_2445);
nand U2895 (N_2895,N_2774,N_2497);
xnor U2896 (N_2896,N_2719,N_2401);
or U2897 (N_2897,N_2546,N_2787);
nor U2898 (N_2898,N_2474,N_2464);
xor U2899 (N_2899,N_2591,N_2528);
and U2900 (N_2900,N_2405,N_2772);
or U2901 (N_2901,N_2657,N_2607);
xnor U2902 (N_2902,N_2409,N_2660);
xnor U2903 (N_2903,N_2587,N_2725);
xnor U2904 (N_2904,N_2586,N_2475);
and U2905 (N_2905,N_2516,N_2421);
nor U2906 (N_2906,N_2402,N_2545);
nand U2907 (N_2907,N_2442,N_2567);
xnor U2908 (N_2908,N_2515,N_2674);
and U2909 (N_2909,N_2530,N_2744);
and U2910 (N_2910,N_2762,N_2539);
xor U2911 (N_2911,N_2668,N_2400);
nor U2912 (N_2912,N_2716,N_2404);
nor U2913 (N_2913,N_2519,N_2788);
nor U2914 (N_2914,N_2576,N_2749);
and U2915 (N_2915,N_2589,N_2766);
or U2916 (N_2916,N_2580,N_2760);
nor U2917 (N_2917,N_2747,N_2726);
nor U2918 (N_2918,N_2642,N_2666);
nor U2919 (N_2919,N_2682,N_2622);
and U2920 (N_2920,N_2430,N_2541);
or U2921 (N_2921,N_2540,N_2729);
nor U2922 (N_2922,N_2781,N_2485);
and U2923 (N_2923,N_2608,N_2751);
and U2924 (N_2924,N_2432,N_2667);
xor U2925 (N_2925,N_2755,N_2419);
nor U2926 (N_2926,N_2613,N_2557);
xnor U2927 (N_2927,N_2649,N_2486);
or U2928 (N_2928,N_2418,N_2569);
nor U2929 (N_2929,N_2765,N_2481);
xor U2930 (N_2930,N_2792,N_2630);
nand U2931 (N_2931,N_2572,N_2520);
or U2932 (N_2932,N_2506,N_2633);
nor U2933 (N_2933,N_2741,N_2625);
or U2934 (N_2934,N_2764,N_2767);
or U2935 (N_2935,N_2703,N_2745);
and U2936 (N_2936,N_2453,N_2721);
xnor U2937 (N_2937,N_2438,N_2436);
xor U2938 (N_2938,N_2730,N_2645);
and U2939 (N_2939,N_2684,N_2407);
nor U2940 (N_2940,N_2694,N_2417);
nor U2941 (N_2941,N_2565,N_2618);
or U2942 (N_2942,N_2582,N_2465);
nor U2943 (N_2943,N_2683,N_2707);
nor U2944 (N_2944,N_2553,N_2502);
nand U2945 (N_2945,N_2451,N_2705);
xor U2946 (N_2946,N_2692,N_2473);
xnor U2947 (N_2947,N_2603,N_2500);
nand U2948 (N_2948,N_2449,N_2455);
nor U2949 (N_2949,N_2691,N_2628);
nand U2950 (N_2950,N_2426,N_2651);
nor U2951 (N_2951,N_2571,N_2686);
nor U2952 (N_2952,N_2662,N_2503);
nand U2953 (N_2953,N_2448,N_2446);
xnor U2954 (N_2954,N_2728,N_2706);
and U2955 (N_2955,N_2568,N_2690);
or U2956 (N_2956,N_2507,N_2678);
xor U2957 (N_2957,N_2484,N_2447);
or U2958 (N_2958,N_2671,N_2532);
nor U2959 (N_2959,N_2784,N_2461);
nor U2960 (N_2960,N_2549,N_2562);
nor U2961 (N_2961,N_2681,N_2471);
nand U2962 (N_2962,N_2415,N_2612);
and U2963 (N_2963,N_2731,N_2710);
nand U2964 (N_2964,N_2509,N_2680);
and U2965 (N_2965,N_2654,N_2531);
and U2966 (N_2966,N_2456,N_2779);
nand U2967 (N_2967,N_2758,N_2510);
xor U2968 (N_2968,N_2718,N_2483);
nand U2969 (N_2969,N_2598,N_2499);
or U2970 (N_2970,N_2798,N_2770);
or U2971 (N_2971,N_2614,N_2577);
or U2972 (N_2972,N_2737,N_2711);
nor U2973 (N_2973,N_2754,N_2536);
xor U2974 (N_2974,N_2646,N_2670);
nand U2975 (N_2975,N_2616,N_2403);
xor U2976 (N_2976,N_2624,N_2701);
nor U2977 (N_2977,N_2736,N_2723);
and U2978 (N_2978,N_2425,N_2482);
or U2979 (N_2979,N_2638,N_2599);
nor U2980 (N_2980,N_2522,N_2634);
nor U2981 (N_2981,N_2491,N_2675);
and U2982 (N_2982,N_2700,N_2742);
xor U2983 (N_2983,N_2410,N_2617);
nor U2984 (N_2984,N_2734,N_2559);
or U2985 (N_2985,N_2641,N_2514);
nand U2986 (N_2986,N_2512,N_2428);
xor U2987 (N_2987,N_2433,N_2790);
nand U2988 (N_2988,N_2494,N_2525);
or U2989 (N_2989,N_2689,N_2708);
and U2990 (N_2990,N_2699,N_2573);
xor U2991 (N_2991,N_2640,N_2561);
nand U2992 (N_2992,N_2796,N_2698);
or U2993 (N_2993,N_2632,N_2585);
and U2994 (N_2994,N_2542,N_2406);
xnor U2995 (N_2995,N_2468,N_2548);
nor U2996 (N_2996,N_2439,N_2513);
and U2997 (N_2997,N_2715,N_2702);
or U2998 (N_2998,N_2527,N_2687);
xnor U2999 (N_2999,N_2434,N_2733);
nor U3000 (N_3000,N_2516,N_2617);
and U3001 (N_3001,N_2561,N_2700);
nor U3002 (N_3002,N_2418,N_2730);
xnor U3003 (N_3003,N_2536,N_2620);
nand U3004 (N_3004,N_2497,N_2765);
and U3005 (N_3005,N_2682,N_2576);
nor U3006 (N_3006,N_2616,N_2438);
xor U3007 (N_3007,N_2579,N_2713);
xnor U3008 (N_3008,N_2420,N_2795);
nor U3009 (N_3009,N_2780,N_2657);
and U3010 (N_3010,N_2712,N_2496);
and U3011 (N_3011,N_2494,N_2781);
or U3012 (N_3012,N_2527,N_2689);
xnor U3013 (N_3013,N_2415,N_2534);
or U3014 (N_3014,N_2693,N_2485);
nand U3015 (N_3015,N_2486,N_2622);
nor U3016 (N_3016,N_2724,N_2463);
nand U3017 (N_3017,N_2732,N_2672);
or U3018 (N_3018,N_2621,N_2671);
nor U3019 (N_3019,N_2569,N_2573);
xnor U3020 (N_3020,N_2680,N_2730);
nand U3021 (N_3021,N_2655,N_2565);
xnor U3022 (N_3022,N_2585,N_2757);
or U3023 (N_3023,N_2400,N_2575);
nor U3024 (N_3024,N_2516,N_2689);
or U3025 (N_3025,N_2531,N_2480);
nand U3026 (N_3026,N_2765,N_2558);
nand U3027 (N_3027,N_2531,N_2718);
nand U3028 (N_3028,N_2544,N_2691);
or U3029 (N_3029,N_2739,N_2400);
and U3030 (N_3030,N_2629,N_2777);
nor U3031 (N_3031,N_2401,N_2462);
xor U3032 (N_3032,N_2705,N_2462);
or U3033 (N_3033,N_2489,N_2682);
or U3034 (N_3034,N_2652,N_2786);
and U3035 (N_3035,N_2418,N_2706);
or U3036 (N_3036,N_2616,N_2622);
nor U3037 (N_3037,N_2512,N_2590);
nand U3038 (N_3038,N_2606,N_2708);
nand U3039 (N_3039,N_2444,N_2576);
nor U3040 (N_3040,N_2412,N_2675);
nor U3041 (N_3041,N_2538,N_2456);
nor U3042 (N_3042,N_2525,N_2797);
or U3043 (N_3043,N_2404,N_2748);
or U3044 (N_3044,N_2762,N_2449);
and U3045 (N_3045,N_2593,N_2476);
nand U3046 (N_3046,N_2665,N_2632);
nor U3047 (N_3047,N_2525,N_2435);
nor U3048 (N_3048,N_2532,N_2465);
nand U3049 (N_3049,N_2621,N_2633);
nor U3050 (N_3050,N_2508,N_2734);
nor U3051 (N_3051,N_2774,N_2417);
nor U3052 (N_3052,N_2646,N_2723);
xor U3053 (N_3053,N_2442,N_2663);
or U3054 (N_3054,N_2748,N_2613);
nor U3055 (N_3055,N_2779,N_2742);
or U3056 (N_3056,N_2523,N_2752);
and U3057 (N_3057,N_2634,N_2709);
xor U3058 (N_3058,N_2665,N_2656);
nor U3059 (N_3059,N_2733,N_2420);
and U3060 (N_3060,N_2739,N_2709);
nand U3061 (N_3061,N_2568,N_2692);
nand U3062 (N_3062,N_2667,N_2492);
and U3063 (N_3063,N_2735,N_2750);
xor U3064 (N_3064,N_2679,N_2429);
and U3065 (N_3065,N_2608,N_2657);
nand U3066 (N_3066,N_2456,N_2610);
and U3067 (N_3067,N_2623,N_2657);
nor U3068 (N_3068,N_2525,N_2718);
or U3069 (N_3069,N_2718,N_2642);
or U3070 (N_3070,N_2548,N_2756);
nand U3071 (N_3071,N_2458,N_2796);
nand U3072 (N_3072,N_2724,N_2460);
and U3073 (N_3073,N_2507,N_2455);
xnor U3074 (N_3074,N_2671,N_2650);
or U3075 (N_3075,N_2486,N_2723);
xnor U3076 (N_3076,N_2480,N_2461);
and U3077 (N_3077,N_2529,N_2479);
xnor U3078 (N_3078,N_2628,N_2484);
xnor U3079 (N_3079,N_2520,N_2582);
nand U3080 (N_3080,N_2464,N_2468);
xor U3081 (N_3081,N_2493,N_2694);
nand U3082 (N_3082,N_2476,N_2660);
xnor U3083 (N_3083,N_2653,N_2559);
and U3084 (N_3084,N_2732,N_2739);
or U3085 (N_3085,N_2671,N_2648);
xnor U3086 (N_3086,N_2582,N_2568);
or U3087 (N_3087,N_2752,N_2570);
nor U3088 (N_3088,N_2658,N_2508);
nand U3089 (N_3089,N_2499,N_2689);
xnor U3090 (N_3090,N_2703,N_2602);
xnor U3091 (N_3091,N_2541,N_2482);
or U3092 (N_3092,N_2445,N_2746);
or U3093 (N_3093,N_2781,N_2415);
or U3094 (N_3094,N_2751,N_2584);
nor U3095 (N_3095,N_2703,N_2458);
xor U3096 (N_3096,N_2537,N_2400);
and U3097 (N_3097,N_2772,N_2672);
or U3098 (N_3098,N_2695,N_2763);
xor U3099 (N_3099,N_2704,N_2514);
xnor U3100 (N_3100,N_2439,N_2444);
nor U3101 (N_3101,N_2448,N_2756);
nor U3102 (N_3102,N_2731,N_2782);
and U3103 (N_3103,N_2756,N_2719);
and U3104 (N_3104,N_2703,N_2570);
nor U3105 (N_3105,N_2593,N_2486);
and U3106 (N_3106,N_2414,N_2466);
or U3107 (N_3107,N_2610,N_2536);
nand U3108 (N_3108,N_2754,N_2745);
and U3109 (N_3109,N_2530,N_2775);
or U3110 (N_3110,N_2517,N_2771);
nand U3111 (N_3111,N_2770,N_2447);
nand U3112 (N_3112,N_2614,N_2765);
or U3113 (N_3113,N_2707,N_2421);
nor U3114 (N_3114,N_2652,N_2655);
xor U3115 (N_3115,N_2451,N_2654);
nand U3116 (N_3116,N_2492,N_2425);
and U3117 (N_3117,N_2775,N_2733);
xnor U3118 (N_3118,N_2456,N_2727);
nand U3119 (N_3119,N_2726,N_2716);
xor U3120 (N_3120,N_2640,N_2413);
nor U3121 (N_3121,N_2402,N_2421);
xnor U3122 (N_3122,N_2672,N_2763);
xnor U3123 (N_3123,N_2678,N_2509);
nand U3124 (N_3124,N_2670,N_2551);
nand U3125 (N_3125,N_2783,N_2538);
nand U3126 (N_3126,N_2610,N_2652);
nand U3127 (N_3127,N_2625,N_2737);
and U3128 (N_3128,N_2463,N_2405);
nand U3129 (N_3129,N_2644,N_2423);
or U3130 (N_3130,N_2671,N_2647);
or U3131 (N_3131,N_2560,N_2750);
or U3132 (N_3132,N_2756,N_2638);
nand U3133 (N_3133,N_2677,N_2553);
xnor U3134 (N_3134,N_2508,N_2704);
xor U3135 (N_3135,N_2497,N_2493);
nor U3136 (N_3136,N_2521,N_2524);
xor U3137 (N_3137,N_2650,N_2436);
and U3138 (N_3138,N_2438,N_2688);
nand U3139 (N_3139,N_2536,N_2556);
nand U3140 (N_3140,N_2524,N_2652);
or U3141 (N_3141,N_2661,N_2516);
or U3142 (N_3142,N_2706,N_2463);
and U3143 (N_3143,N_2410,N_2493);
xor U3144 (N_3144,N_2531,N_2476);
or U3145 (N_3145,N_2422,N_2545);
nor U3146 (N_3146,N_2633,N_2622);
nor U3147 (N_3147,N_2478,N_2749);
or U3148 (N_3148,N_2503,N_2588);
or U3149 (N_3149,N_2681,N_2506);
and U3150 (N_3150,N_2658,N_2628);
nor U3151 (N_3151,N_2600,N_2606);
and U3152 (N_3152,N_2611,N_2479);
nor U3153 (N_3153,N_2460,N_2774);
or U3154 (N_3154,N_2488,N_2451);
nand U3155 (N_3155,N_2427,N_2756);
or U3156 (N_3156,N_2722,N_2676);
xor U3157 (N_3157,N_2454,N_2634);
nand U3158 (N_3158,N_2710,N_2517);
xnor U3159 (N_3159,N_2685,N_2462);
or U3160 (N_3160,N_2714,N_2783);
nor U3161 (N_3161,N_2416,N_2504);
and U3162 (N_3162,N_2743,N_2577);
nor U3163 (N_3163,N_2718,N_2730);
or U3164 (N_3164,N_2577,N_2516);
nand U3165 (N_3165,N_2643,N_2467);
and U3166 (N_3166,N_2776,N_2574);
nand U3167 (N_3167,N_2626,N_2423);
nand U3168 (N_3168,N_2616,N_2662);
nor U3169 (N_3169,N_2567,N_2626);
or U3170 (N_3170,N_2781,N_2702);
and U3171 (N_3171,N_2723,N_2545);
nand U3172 (N_3172,N_2400,N_2509);
nand U3173 (N_3173,N_2764,N_2476);
and U3174 (N_3174,N_2680,N_2409);
nor U3175 (N_3175,N_2455,N_2667);
nand U3176 (N_3176,N_2778,N_2424);
and U3177 (N_3177,N_2678,N_2788);
nor U3178 (N_3178,N_2737,N_2750);
nor U3179 (N_3179,N_2569,N_2421);
nand U3180 (N_3180,N_2482,N_2587);
nor U3181 (N_3181,N_2449,N_2547);
and U3182 (N_3182,N_2629,N_2578);
nor U3183 (N_3183,N_2633,N_2521);
nand U3184 (N_3184,N_2775,N_2446);
and U3185 (N_3185,N_2497,N_2536);
nor U3186 (N_3186,N_2424,N_2631);
or U3187 (N_3187,N_2629,N_2657);
or U3188 (N_3188,N_2661,N_2558);
xnor U3189 (N_3189,N_2628,N_2480);
xor U3190 (N_3190,N_2485,N_2695);
and U3191 (N_3191,N_2737,N_2637);
or U3192 (N_3192,N_2560,N_2640);
or U3193 (N_3193,N_2562,N_2564);
or U3194 (N_3194,N_2568,N_2410);
and U3195 (N_3195,N_2594,N_2471);
and U3196 (N_3196,N_2780,N_2476);
or U3197 (N_3197,N_2716,N_2673);
nand U3198 (N_3198,N_2651,N_2703);
xor U3199 (N_3199,N_2784,N_2537);
or U3200 (N_3200,N_2964,N_3043);
nand U3201 (N_3201,N_3107,N_3181);
nand U3202 (N_3202,N_2802,N_3068);
or U3203 (N_3203,N_3103,N_2811);
nor U3204 (N_3204,N_3122,N_2924);
nor U3205 (N_3205,N_3047,N_2866);
nand U3206 (N_3206,N_3131,N_2949);
or U3207 (N_3207,N_2813,N_2872);
nor U3208 (N_3208,N_2932,N_2824);
nor U3209 (N_3209,N_3017,N_2886);
and U3210 (N_3210,N_3045,N_2981);
xnor U3211 (N_3211,N_3028,N_2898);
nand U3212 (N_3212,N_3033,N_2889);
or U3213 (N_3213,N_3167,N_3057);
and U3214 (N_3214,N_3083,N_3158);
nand U3215 (N_3215,N_2909,N_3048);
nand U3216 (N_3216,N_2925,N_3100);
or U3217 (N_3217,N_2881,N_3141);
xor U3218 (N_3218,N_2896,N_2833);
and U3219 (N_3219,N_2871,N_3104);
nor U3220 (N_3220,N_3007,N_2825);
and U3221 (N_3221,N_3012,N_2879);
nor U3222 (N_3222,N_3164,N_3024);
or U3223 (N_3223,N_3066,N_3003);
nor U3224 (N_3224,N_3002,N_3005);
nand U3225 (N_3225,N_2913,N_3163);
and U3226 (N_3226,N_2972,N_3187);
and U3227 (N_3227,N_2991,N_3172);
nand U3228 (N_3228,N_3199,N_2959);
or U3229 (N_3229,N_2857,N_2996);
or U3230 (N_3230,N_3085,N_3174);
nor U3231 (N_3231,N_2803,N_3123);
or U3232 (N_3232,N_2927,N_3064);
nor U3233 (N_3233,N_3126,N_2821);
and U3234 (N_3234,N_2910,N_3088);
xnor U3235 (N_3235,N_3050,N_3193);
and U3236 (N_3236,N_2890,N_2868);
nand U3237 (N_3237,N_3112,N_3188);
xor U3238 (N_3238,N_2990,N_3190);
and U3239 (N_3239,N_3102,N_3134);
and U3240 (N_3240,N_3150,N_2893);
nor U3241 (N_3241,N_2852,N_3159);
nand U3242 (N_3242,N_3145,N_3180);
xor U3243 (N_3243,N_2926,N_3095);
nor U3244 (N_3244,N_3021,N_2834);
xor U3245 (N_3245,N_3179,N_3069);
xor U3246 (N_3246,N_2930,N_2907);
or U3247 (N_3247,N_2837,N_2920);
or U3248 (N_3248,N_3182,N_3168);
and U3249 (N_3249,N_3132,N_3119);
and U3250 (N_3250,N_2812,N_2974);
xnor U3251 (N_3251,N_3004,N_3037);
nand U3252 (N_3252,N_3098,N_3053);
xnor U3253 (N_3253,N_3041,N_3177);
and U3254 (N_3254,N_2988,N_2903);
or U3255 (N_3255,N_3148,N_2955);
and U3256 (N_3256,N_2921,N_2846);
nand U3257 (N_3257,N_2801,N_3192);
nand U3258 (N_3258,N_2819,N_3097);
or U3259 (N_3259,N_3128,N_2968);
xnor U3260 (N_3260,N_3059,N_2978);
nor U3261 (N_3261,N_3061,N_3115);
xor U3262 (N_3262,N_3154,N_3042);
xnor U3263 (N_3263,N_3035,N_2912);
nor U3264 (N_3264,N_2805,N_3006);
xor U3265 (N_3265,N_3165,N_2975);
or U3266 (N_3266,N_3136,N_2832);
or U3267 (N_3267,N_2940,N_2993);
or U3268 (N_3268,N_2804,N_2947);
nand U3269 (N_3269,N_3087,N_2944);
nor U3270 (N_3270,N_3143,N_2841);
xor U3271 (N_3271,N_2830,N_2900);
nor U3272 (N_3272,N_3171,N_3118);
nor U3273 (N_3273,N_2800,N_2906);
and U3274 (N_3274,N_2863,N_3151);
or U3275 (N_3275,N_3025,N_3147);
and U3276 (N_3276,N_2983,N_2874);
or U3277 (N_3277,N_2885,N_2839);
nand U3278 (N_3278,N_3146,N_3133);
xnor U3279 (N_3279,N_3011,N_3170);
and U3280 (N_3280,N_2880,N_3065);
xor U3281 (N_3281,N_3009,N_2847);
or U3282 (N_3282,N_2862,N_2901);
and U3283 (N_3283,N_3022,N_3052);
nor U3284 (N_3284,N_2958,N_2894);
and U3285 (N_3285,N_2997,N_2922);
nor U3286 (N_3286,N_2979,N_2904);
or U3287 (N_3287,N_2814,N_3135);
nand U3288 (N_3288,N_2923,N_3081);
or U3289 (N_3289,N_2960,N_3078);
or U3290 (N_3290,N_2953,N_3054);
nand U3291 (N_3291,N_3157,N_3019);
xnor U3292 (N_3292,N_2992,N_3039);
and U3293 (N_3293,N_3176,N_2843);
and U3294 (N_3294,N_2838,N_2897);
nor U3295 (N_3295,N_3000,N_2938);
xnor U3296 (N_3296,N_2876,N_3169);
or U3297 (N_3297,N_3191,N_3178);
xor U3298 (N_3298,N_3189,N_3013);
nand U3299 (N_3299,N_2840,N_3055);
or U3300 (N_3300,N_3029,N_3092);
or U3301 (N_3301,N_3175,N_2963);
nand U3302 (N_3302,N_3138,N_3109);
xor U3303 (N_3303,N_3096,N_2877);
or U3304 (N_3304,N_3020,N_2809);
and U3305 (N_3305,N_3018,N_2845);
xor U3306 (N_3306,N_2956,N_3044);
xor U3307 (N_3307,N_2895,N_2854);
and U3308 (N_3308,N_3117,N_2950);
and U3309 (N_3309,N_2995,N_3183);
nor U3310 (N_3310,N_3070,N_3063);
or U3311 (N_3311,N_3166,N_2945);
and U3312 (N_3312,N_3086,N_2962);
nand U3313 (N_3313,N_2883,N_2977);
nand U3314 (N_3314,N_2954,N_3142);
or U3315 (N_3315,N_2858,N_3040);
and U3316 (N_3316,N_3038,N_2970);
or U3317 (N_3317,N_2861,N_3058);
nor U3318 (N_3318,N_3110,N_3030);
and U3319 (N_3319,N_2882,N_3160);
xnor U3320 (N_3320,N_3090,N_2943);
or U3321 (N_3321,N_3075,N_2929);
or U3322 (N_3322,N_2888,N_2859);
xor U3323 (N_3323,N_2986,N_2937);
and U3324 (N_3324,N_2931,N_3127);
nor U3325 (N_3325,N_2994,N_3010);
nor U3326 (N_3326,N_2965,N_2853);
nand U3327 (N_3327,N_2849,N_2817);
and U3328 (N_3328,N_3062,N_3162);
or U3329 (N_3329,N_2942,N_3089);
nor U3330 (N_3330,N_3111,N_2902);
or U3331 (N_3331,N_2869,N_3125);
xor U3332 (N_3332,N_2878,N_2915);
or U3333 (N_3333,N_2864,N_3108);
and U3334 (N_3334,N_2884,N_3140);
xnor U3335 (N_3335,N_3099,N_2916);
nand U3336 (N_3336,N_3144,N_3173);
or U3337 (N_3337,N_2820,N_2818);
and U3338 (N_3338,N_2939,N_2842);
and U3339 (N_3339,N_3080,N_2917);
or U3340 (N_3340,N_2957,N_2831);
and U3341 (N_3341,N_2999,N_3161);
nor U3342 (N_3342,N_2961,N_3027);
nand U3343 (N_3343,N_2850,N_3186);
nor U3344 (N_3344,N_2844,N_2856);
or U3345 (N_3345,N_3073,N_2985);
nand U3346 (N_3346,N_3184,N_3195);
xnor U3347 (N_3347,N_3032,N_3023);
nand U3348 (N_3348,N_3113,N_3077);
xnor U3349 (N_3349,N_2899,N_2976);
nand U3350 (N_3350,N_2836,N_2827);
xnor U3351 (N_3351,N_2865,N_2951);
xor U3352 (N_3352,N_3076,N_3001);
and U3353 (N_3353,N_3137,N_2969);
or U3354 (N_3354,N_2998,N_2914);
nand U3355 (N_3355,N_3079,N_2919);
and U3356 (N_3356,N_2918,N_3060);
nor U3357 (N_3357,N_2887,N_3049);
xor U3358 (N_3358,N_3056,N_3153);
or U3359 (N_3359,N_2891,N_2855);
or U3360 (N_3360,N_2806,N_3036);
nor U3361 (N_3361,N_2851,N_2870);
nand U3362 (N_3362,N_2908,N_2933);
or U3363 (N_3363,N_2816,N_3155);
or U3364 (N_3364,N_3198,N_3152);
xnor U3365 (N_3365,N_3106,N_3051);
and U3366 (N_3366,N_3026,N_2875);
or U3367 (N_3367,N_2807,N_2835);
nor U3368 (N_3368,N_3071,N_3031);
or U3369 (N_3369,N_2892,N_3129);
xnor U3370 (N_3370,N_3194,N_2810);
or U3371 (N_3371,N_2848,N_3105);
and U3372 (N_3372,N_2952,N_2823);
and U3373 (N_3373,N_3094,N_2905);
nor U3374 (N_3374,N_2867,N_2973);
or U3375 (N_3375,N_2948,N_3197);
nor U3376 (N_3376,N_2828,N_2934);
and U3377 (N_3377,N_2829,N_3084);
or U3378 (N_3378,N_3196,N_3072);
and U3379 (N_3379,N_2911,N_3121);
xnor U3380 (N_3380,N_2966,N_2808);
and U3381 (N_3381,N_3034,N_3082);
and U3382 (N_3382,N_2980,N_3014);
xor U3383 (N_3383,N_3074,N_3149);
xor U3384 (N_3384,N_3046,N_2982);
xnor U3385 (N_3385,N_2822,N_3015);
nand U3386 (N_3386,N_3114,N_2936);
xnor U3387 (N_3387,N_2984,N_3185);
nand U3388 (N_3388,N_2971,N_3120);
nand U3389 (N_3389,N_3016,N_3130);
and U3390 (N_3390,N_2873,N_2941);
nand U3391 (N_3391,N_2935,N_2815);
nand U3392 (N_3392,N_2946,N_2860);
and U3393 (N_3393,N_3116,N_2928);
nor U3394 (N_3394,N_3093,N_3156);
nor U3395 (N_3395,N_3124,N_3139);
xor U3396 (N_3396,N_2967,N_2987);
nand U3397 (N_3397,N_3067,N_3101);
or U3398 (N_3398,N_2826,N_2989);
and U3399 (N_3399,N_3091,N_3008);
nor U3400 (N_3400,N_3004,N_2878);
or U3401 (N_3401,N_3193,N_2866);
nor U3402 (N_3402,N_3079,N_2991);
nor U3403 (N_3403,N_3043,N_2849);
xor U3404 (N_3404,N_2951,N_3183);
or U3405 (N_3405,N_3017,N_3008);
xor U3406 (N_3406,N_2867,N_2948);
nand U3407 (N_3407,N_3112,N_3134);
nor U3408 (N_3408,N_3186,N_2959);
nand U3409 (N_3409,N_3033,N_2867);
nand U3410 (N_3410,N_3043,N_2951);
nor U3411 (N_3411,N_3062,N_2874);
xor U3412 (N_3412,N_2878,N_3185);
nor U3413 (N_3413,N_2809,N_3112);
nor U3414 (N_3414,N_3098,N_3116);
or U3415 (N_3415,N_2904,N_2870);
or U3416 (N_3416,N_2960,N_2946);
or U3417 (N_3417,N_3070,N_3051);
nand U3418 (N_3418,N_3018,N_2908);
nor U3419 (N_3419,N_2924,N_3107);
and U3420 (N_3420,N_2934,N_3127);
xnor U3421 (N_3421,N_2921,N_3133);
nand U3422 (N_3422,N_3083,N_3136);
nand U3423 (N_3423,N_3087,N_2827);
xor U3424 (N_3424,N_2802,N_2831);
nor U3425 (N_3425,N_3153,N_3100);
xnor U3426 (N_3426,N_3163,N_3073);
or U3427 (N_3427,N_3169,N_3127);
nand U3428 (N_3428,N_3185,N_2873);
and U3429 (N_3429,N_2964,N_2895);
xor U3430 (N_3430,N_3136,N_3166);
or U3431 (N_3431,N_2902,N_2847);
or U3432 (N_3432,N_3165,N_2968);
nand U3433 (N_3433,N_3036,N_3182);
or U3434 (N_3434,N_3069,N_2944);
and U3435 (N_3435,N_2848,N_3108);
nand U3436 (N_3436,N_2843,N_3081);
xnor U3437 (N_3437,N_3172,N_3179);
nor U3438 (N_3438,N_2970,N_2947);
nand U3439 (N_3439,N_2800,N_2808);
nor U3440 (N_3440,N_2904,N_3080);
nand U3441 (N_3441,N_2904,N_3162);
and U3442 (N_3442,N_2846,N_3119);
and U3443 (N_3443,N_2810,N_2886);
xnor U3444 (N_3444,N_2802,N_2891);
nand U3445 (N_3445,N_3069,N_3084);
xnor U3446 (N_3446,N_2985,N_2825);
and U3447 (N_3447,N_2836,N_3161);
or U3448 (N_3448,N_2830,N_3186);
nand U3449 (N_3449,N_3017,N_2844);
or U3450 (N_3450,N_2961,N_2935);
xor U3451 (N_3451,N_3074,N_2852);
or U3452 (N_3452,N_2990,N_3140);
and U3453 (N_3453,N_3165,N_2997);
or U3454 (N_3454,N_2919,N_2998);
and U3455 (N_3455,N_3098,N_3120);
nand U3456 (N_3456,N_3054,N_3019);
and U3457 (N_3457,N_3177,N_2928);
and U3458 (N_3458,N_3126,N_3089);
and U3459 (N_3459,N_2810,N_3198);
or U3460 (N_3460,N_2850,N_3111);
nor U3461 (N_3461,N_2815,N_2913);
xnor U3462 (N_3462,N_2936,N_3020);
or U3463 (N_3463,N_3184,N_2871);
nand U3464 (N_3464,N_3169,N_2937);
xnor U3465 (N_3465,N_3067,N_2960);
or U3466 (N_3466,N_3011,N_2901);
nand U3467 (N_3467,N_2954,N_3078);
and U3468 (N_3468,N_3084,N_2861);
nand U3469 (N_3469,N_2882,N_3168);
or U3470 (N_3470,N_3031,N_3129);
and U3471 (N_3471,N_2949,N_3111);
or U3472 (N_3472,N_3185,N_2817);
nand U3473 (N_3473,N_2832,N_3089);
or U3474 (N_3474,N_3060,N_3073);
nor U3475 (N_3475,N_2825,N_3181);
xor U3476 (N_3476,N_2810,N_3033);
xor U3477 (N_3477,N_3041,N_3186);
or U3478 (N_3478,N_2853,N_2892);
and U3479 (N_3479,N_3077,N_2943);
or U3480 (N_3480,N_2913,N_2859);
nand U3481 (N_3481,N_2822,N_2945);
nand U3482 (N_3482,N_2953,N_2853);
and U3483 (N_3483,N_2913,N_2892);
xnor U3484 (N_3484,N_2873,N_2864);
and U3485 (N_3485,N_2914,N_3153);
and U3486 (N_3486,N_3043,N_2916);
nor U3487 (N_3487,N_3088,N_2864);
or U3488 (N_3488,N_2811,N_2979);
and U3489 (N_3489,N_2993,N_2924);
and U3490 (N_3490,N_3040,N_3051);
or U3491 (N_3491,N_3040,N_3101);
nand U3492 (N_3492,N_2868,N_3141);
and U3493 (N_3493,N_2805,N_2858);
nor U3494 (N_3494,N_2841,N_3189);
nand U3495 (N_3495,N_3021,N_2824);
xor U3496 (N_3496,N_2920,N_2968);
nor U3497 (N_3497,N_2806,N_2981);
nor U3498 (N_3498,N_3193,N_3110);
nor U3499 (N_3499,N_3192,N_2863);
nor U3500 (N_3500,N_2899,N_2989);
nand U3501 (N_3501,N_3199,N_2917);
nand U3502 (N_3502,N_3090,N_3088);
nor U3503 (N_3503,N_2848,N_3158);
xnor U3504 (N_3504,N_2891,N_3003);
nor U3505 (N_3505,N_3025,N_3161);
nor U3506 (N_3506,N_3061,N_3105);
nor U3507 (N_3507,N_2855,N_2903);
or U3508 (N_3508,N_3088,N_2930);
nand U3509 (N_3509,N_2989,N_3078);
or U3510 (N_3510,N_2942,N_2940);
nor U3511 (N_3511,N_3146,N_3039);
nor U3512 (N_3512,N_2873,N_2841);
xnor U3513 (N_3513,N_3183,N_2996);
or U3514 (N_3514,N_2838,N_2878);
nand U3515 (N_3515,N_2878,N_3113);
nor U3516 (N_3516,N_3152,N_2859);
nand U3517 (N_3517,N_3046,N_2962);
and U3518 (N_3518,N_3090,N_2972);
nor U3519 (N_3519,N_3071,N_2876);
and U3520 (N_3520,N_3006,N_2817);
nor U3521 (N_3521,N_2980,N_2890);
and U3522 (N_3522,N_2813,N_2944);
or U3523 (N_3523,N_3020,N_2920);
xor U3524 (N_3524,N_3153,N_2939);
nor U3525 (N_3525,N_2916,N_3183);
xnor U3526 (N_3526,N_3141,N_2939);
or U3527 (N_3527,N_3162,N_3185);
and U3528 (N_3528,N_2875,N_2927);
or U3529 (N_3529,N_2849,N_2920);
xor U3530 (N_3530,N_2889,N_3024);
and U3531 (N_3531,N_3149,N_3053);
nand U3532 (N_3532,N_3083,N_3098);
xnor U3533 (N_3533,N_3198,N_3166);
xor U3534 (N_3534,N_2868,N_2804);
and U3535 (N_3535,N_3081,N_3047);
or U3536 (N_3536,N_2956,N_2894);
nand U3537 (N_3537,N_2881,N_3085);
xnor U3538 (N_3538,N_2842,N_3049);
xnor U3539 (N_3539,N_2958,N_2801);
or U3540 (N_3540,N_2801,N_2803);
nor U3541 (N_3541,N_2993,N_2920);
nor U3542 (N_3542,N_3184,N_3158);
nand U3543 (N_3543,N_3149,N_3034);
nand U3544 (N_3544,N_2928,N_3023);
xor U3545 (N_3545,N_3169,N_3158);
and U3546 (N_3546,N_2999,N_2946);
nor U3547 (N_3547,N_3080,N_2918);
nand U3548 (N_3548,N_3031,N_3015);
or U3549 (N_3549,N_2869,N_3157);
xnor U3550 (N_3550,N_3064,N_2836);
and U3551 (N_3551,N_2983,N_2945);
nor U3552 (N_3552,N_3156,N_2966);
or U3553 (N_3553,N_2938,N_2870);
nor U3554 (N_3554,N_3078,N_3157);
or U3555 (N_3555,N_3104,N_3019);
nor U3556 (N_3556,N_3010,N_2960);
and U3557 (N_3557,N_2947,N_3068);
and U3558 (N_3558,N_3036,N_3054);
nor U3559 (N_3559,N_3026,N_2814);
nand U3560 (N_3560,N_3107,N_2967);
xnor U3561 (N_3561,N_3192,N_2973);
nor U3562 (N_3562,N_2828,N_2866);
nand U3563 (N_3563,N_3137,N_2850);
nand U3564 (N_3564,N_2855,N_3069);
xnor U3565 (N_3565,N_2825,N_2824);
and U3566 (N_3566,N_2940,N_3052);
and U3567 (N_3567,N_2907,N_2867);
and U3568 (N_3568,N_2806,N_2989);
nor U3569 (N_3569,N_2881,N_2918);
nand U3570 (N_3570,N_3064,N_3099);
xor U3571 (N_3571,N_3004,N_3149);
nor U3572 (N_3572,N_3046,N_3159);
xnor U3573 (N_3573,N_3062,N_2817);
xor U3574 (N_3574,N_3093,N_3194);
nor U3575 (N_3575,N_3011,N_2971);
xor U3576 (N_3576,N_3085,N_3012);
nor U3577 (N_3577,N_3136,N_3137);
xnor U3578 (N_3578,N_3185,N_2994);
nor U3579 (N_3579,N_2901,N_3047);
nor U3580 (N_3580,N_3137,N_3069);
nand U3581 (N_3581,N_2815,N_2930);
nand U3582 (N_3582,N_3186,N_2871);
nor U3583 (N_3583,N_2870,N_2946);
nand U3584 (N_3584,N_3099,N_3013);
or U3585 (N_3585,N_2887,N_3012);
and U3586 (N_3586,N_3182,N_3065);
xnor U3587 (N_3587,N_3186,N_2836);
xnor U3588 (N_3588,N_2951,N_2893);
xnor U3589 (N_3589,N_3021,N_2973);
nand U3590 (N_3590,N_3119,N_2915);
xor U3591 (N_3591,N_2897,N_3022);
nor U3592 (N_3592,N_3013,N_3023);
nor U3593 (N_3593,N_3181,N_3017);
nand U3594 (N_3594,N_2811,N_2908);
or U3595 (N_3595,N_3075,N_3065);
nand U3596 (N_3596,N_2859,N_3098);
and U3597 (N_3597,N_2986,N_3091);
nor U3598 (N_3598,N_3121,N_2960);
nand U3599 (N_3599,N_2945,N_3129);
xor U3600 (N_3600,N_3492,N_3510);
nor U3601 (N_3601,N_3363,N_3581);
nor U3602 (N_3602,N_3205,N_3453);
or U3603 (N_3603,N_3253,N_3237);
and U3604 (N_3604,N_3270,N_3327);
or U3605 (N_3605,N_3257,N_3209);
xor U3606 (N_3606,N_3290,N_3494);
xnor U3607 (N_3607,N_3440,N_3439);
and U3608 (N_3608,N_3296,N_3304);
or U3609 (N_3609,N_3201,N_3335);
nand U3610 (N_3610,N_3218,N_3305);
nor U3611 (N_3611,N_3476,N_3558);
nor U3612 (N_3612,N_3544,N_3520);
or U3613 (N_3613,N_3217,N_3478);
nor U3614 (N_3614,N_3463,N_3405);
nor U3615 (N_3615,N_3452,N_3248);
or U3616 (N_3616,N_3243,N_3228);
nor U3617 (N_3617,N_3388,N_3281);
nand U3618 (N_3618,N_3576,N_3449);
nor U3619 (N_3619,N_3341,N_3414);
xnor U3620 (N_3620,N_3357,N_3545);
and U3621 (N_3621,N_3409,N_3344);
and U3622 (N_3622,N_3299,N_3391);
and U3623 (N_3623,N_3429,N_3285);
or U3624 (N_3624,N_3501,N_3559);
nand U3625 (N_3625,N_3435,N_3503);
nor U3626 (N_3626,N_3361,N_3508);
nand U3627 (N_3627,N_3204,N_3245);
and U3628 (N_3628,N_3360,N_3536);
or U3629 (N_3629,N_3365,N_3533);
or U3630 (N_3630,N_3460,N_3434);
or U3631 (N_3631,N_3423,N_3333);
xnor U3632 (N_3632,N_3349,N_3526);
or U3633 (N_3633,N_3548,N_3546);
xor U3634 (N_3634,N_3264,N_3272);
or U3635 (N_3635,N_3366,N_3359);
nor U3636 (N_3636,N_3597,N_3376);
and U3637 (N_3637,N_3256,N_3223);
and U3638 (N_3638,N_3258,N_3567);
and U3639 (N_3639,N_3455,N_3518);
xnor U3640 (N_3640,N_3266,N_3240);
or U3641 (N_3641,N_3332,N_3337);
nand U3642 (N_3642,N_3249,N_3527);
or U3643 (N_3643,N_3397,N_3324);
nor U3644 (N_3644,N_3474,N_3566);
or U3645 (N_3645,N_3431,N_3428);
nor U3646 (N_3646,N_3315,N_3417);
or U3647 (N_3647,N_3400,N_3513);
and U3648 (N_3648,N_3347,N_3499);
nand U3649 (N_3649,N_3459,N_3379);
nor U3650 (N_3650,N_3259,N_3458);
or U3651 (N_3651,N_3496,N_3557);
nand U3652 (N_3652,N_3252,N_3320);
nor U3653 (N_3653,N_3251,N_3308);
xor U3654 (N_3654,N_3580,N_3346);
and U3655 (N_3655,N_3437,N_3387);
nor U3656 (N_3656,N_3532,N_3329);
nor U3657 (N_3657,N_3396,N_3582);
nor U3658 (N_3658,N_3589,N_3464);
nand U3659 (N_3659,N_3512,N_3471);
xnor U3660 (N_3660,N_3301,N_3556);
or U3661 (N_3661,N_3490,N_3595);
nand U3662 (N_3662,N_3410,N_3331);
and U3663 (N_3663,N_3418,N_3424);
or U3664 (N_3664,N_3214,N_3554);
xor U3665 (N_3665,N_3367,N_3551);
xnor U3666 (N_3666,N_3506,N_3398);
and U3667 (N_3667,N_3489,N_3593);
nand U3668 (N_3668,N_3339,N_3383);
xor U3669 (N_3669,N_3528,N_3284);
xnor U3670 (N_3670,N_3564,N_3465);
and U3671 (N_3671,N_3336,N_3226);
nand U3672 (N_3672,N_3220,N_3571);
or U3673 (N_3673,N_3356,N_3411);
or U3674 (N_3674,N_3491,N_3416);
or U3675 (N_3675,N_3591,N_3210);
nor U3676 (N_3676,N_3487,N_3535);
xnor U3677 (N_3677,N_3403,N_3524);
or U3678 (N_3678,N_3280,N_3314);
nor U3679 (N_3679,N_3343,N_3294);
nor U3680 (N_3680,N_3348,N_3569);
nand U3681 (N_3681,N_3592,N_3594);
or U3682 (N_3682,N_3211,N_3541);
xor U3683 (N_3683,N_3234,N_3354);
nand U3684 (N_3684,N_3480,N_3224);
nor U3685 (N_3685,N_3547,N_3529);
xor U3686 (N_3686,N_3579,N_3374);
nand U3687 (N_3687,N_3488,N_3353);
xor U3688 (N_3688,N_3207,N_3586);
or U3689 (N_3689,N_3287,N_3511);
and U3690 (N_3690,N_3467,N_3275);
and U3691 (N_3691,N_3422,N_3380);
or U3692 (N_3692,N_3384,N_3202);
or U3693 (N_3693,N_3462,N_3229);
nand U3694 (N_3694,N_3330,N_3408);
nand U3695 (N_3695,N_3325,N_3441);
xnor U3696 (N_3696,N_3574,N_3382);
or U3697 (N_3697,N_3470,N_3230);
or U3698 (N_3698,N_3446,N_3369);
and U3699 (N_3699,N_3584,N_3454);
and U3700 (N_3700,N_3468,N_3427);
or U3701 (N_3701,N_3502,N_3432);
or U3702 (N_3702,N_3438,N_3246);
or U3703 (N_3703,N_3572,N_3260);
or U3704 (N_3704,N_3537,N_3568);
or U3705 (N_3705,N_3216,N_3504);
or U3706 (N_3706,N_3358,N_3412);
nand U3707 (N_3707,N_3406,N_3493);
and U3708 (N_3708,N_3451,N_3538);
or U3709 (N_3709,N_3507,N_3263);
and U3710 (N_3710,N_3552,N_3386);
xnor U3711 (N_3711,N_3231,N_3563);
nand U3712 (N_3712,N_3352,N_3222);
and U3713 (N_3713,N_3534,N_3485);
nor U3714 (N_3714,N_3543,N_3585);
nand U3715 (N_3715,N_3555,N_3312);
and U3716 (N_3716,N_3540,N_3262);
nand U3717 (N_3717,N_3522,N_3407);
or U3718 (N_3718,N_3283,N_3271);
and U3719 (N_3719,N_3241,N_3340);
and U3720 (N_3720,N_3447,N_3306);
xnor U3721 (N_3721,N_3461,N_3208);
nor U3722 (N_3722,N_3570,N_3292);
or U3723 (N_3723,N_3355,N_3206);
nor U3724 (N_3724,N_3390,N_3484);
xor U3725 (N_3725,N_3345,N_3255);
nand U3726 (N_3726,N_3531,N_3273);
xor U3727 (N_3727,N_3232,N_3278);
nor U3728 (N_3728,N_3368,N_3486);
or U3729 (N_3729,N_3542,N_3371);
nor U3730 (N_3730,N_3481,N_3268);
nand U3731 (N_3731,N_3338,N_3297);
and U3732 (N_3732,N_3415,N_3466);
nor U3733 (N_3733,N_3475,N_3575);
or U3734 (N_3734,N_3247,N_3307);
nand U3735 (N_3735,N_3373,N_3318);
nand U3736 (N_3736,N_3565,N_3221);
and U3737 (N_3737,N_3573,N_3239);
nand U3738 (N_3738,N_3291,N_3238);
nand U3739 (N_3739,N_3436,N_3514);
nand U3740 (N_3740,N_3378,N_3293);
nand U3741 (N_3741,N_3313,N_3517);
nand U3742 (N_3742,N_3413,N_3402);
nor U3743 (N_3743,N_3225,N_3394);
and U3744 (N_3744,N_3375,N_3300);
xnor U3745 (N_3745,N_3261,N_3482);
nor U3746 (N_3746,N_3203,N_3236);
xor U3747 (N_3747,N_3596,N_3500);
or U3748 (N_3748,N_3530,N_3473);
nor U3749 (N_3749,N_3282,N_3539);
and U3750 (N_3750,N_3242,N_3598);
and U3751 (N_3751,N_3560,N_3448);
nor U3752 (N_3752,N_3286,N_3381);
and U3753 (N_3753,N_3342,N_3497);
or U3754 (N_3754,N_3303,N_3350);
or U3755 (N_3755,N_3395,N_3421);
nor U3756 (N_3756,N_3515,N_3426);
and U3757 (N_3757,N_3457,N_3277);
nor U3758 (N_3758,N_3479,N_3495);
nand U3759 (N_3759,N_3254,N_3392);
and U3760 (N_3760,N_3279,N_3583);
xor U3761 (N_3761,N_3267,N_3445);
or U3762 (N_3762,N_3521,N_3235);
nor U3763 (N_3763,N_3227,N_3323);
nor U3764 (N_3764,N_3212,N_3433);
nor U3765 (N_3765,N_3483,N_3269);
xnor U3766 (N_3766,N_3276,N_3516);
and U3767 (N_3767,N_3334,N_3393);
xnor U3768 (N_3768,N_3364,N_3590);
and U3769 (N_3769,N_3523,N_3385);
nor U3770 (N_3770,N_3319,N_3244);
and U3771 (N_3771,N_3450,N_3509);
nand U3772 (N_3772,N_3311,N_3322);
nor U3773 (N_3773,N_3456,N_3389);
nor U3774 (N_3774,N_3250,N_3321);
and U3775 (N_3775,N_3498,N_3213);
and U3776 (N_3776,N_3309,N_3298);
and U3777 (N_3777,N_3351,N_3477);
nand U3778 (N_3778,N_3317,N_3362);
nor U3779 (N_3779,N_3550,N_3443);
nand U3780 (N_3780,N_3404,N_3587);
xor U3781 (N_3781,N_3549,N_3442);
or U3782 (N_3782,N_3316,N_3525);
or U3783 (N_3783,N_3233,N_3472);
xnor U3784 (N_3784,N_3430,N_3295);
xnor U3785 (N_3785,N_3577,N_3562);
or U3786 (N_3786,N_3328,N_3377);
or U3787 (N_3787,N_3370,N_3444);
and U3788 (N_3788,N_3310,N_3425);
or U3789 (N_3789,N_3505,N_3553);
and U3790 (N_3790,N_3469,N_3401);
xnor U3791 (N_3791,N_3399,N_3588);
nor U3792 (N_3792,N_3419,N_3200);
nand U3793 (N_3793,N_3420,N_3561);
or U3794 (N_3794,N_3265,N_3302);
or U3795 (N_3795,N_3599,N_3326);
nor U3796 (N_3796,N_3215,N_3274);
nor U3797 (N_3797,N_3219,N_3578);
nor U3798 (N_3798,N_3289,N_3372);
nor U3799 (N_3799,N_3288,N_3519);
xor U3800 (N_3800,N_3359,N_3321);
nor U3801 (N_3801,N_3265,N_3461);
or U3802 (N_3802,N_3496,N_3245);
or U3803 (N_3803,N_3460,N_3285);
xnor U3804 (N_3804,N_3250,N_3425);
or U3805 (N_3805,N_3567,N_3270);
xnor U3806 (N_3806,N_3333,N_3375);
nand U3807 (N_3807,N_3542,N_3415);
nand U3808 (N_3808,N_3273,N_3277);
nand U3809 (N_3809,N_3420,N_3488);
nor U3810 (N_3810,N_3384,N_3287);
nand U3811 (N_3811,N_3450,N_3559);
or U3812 (N_3812,N_3530,N_3534);
nand U3813 (N_3813,N_3370,N_3348);
nand U3814 (N_3814,N_3401,N_3279);
nand U3815 (N_3815,N_3341,N_3573);
nor U3816 (N_3816,N_3286,N_3516);
nor U3817 (N_3817,N_3594,N_3241);
and U3818 (N_3818,N_3293,N_3485);
nor U3819 (N_3819,N_3280,N_3294);
and U3820 (N_3820,N_3471,N_3208);
nand U3821 (N_3821,N_3321,N_3467);
nand U3822 (N_3822,N_3473,N_3429);
and U3823 (N_3823,N_3530,N_3445);
or U3824 (N_3824,N_3581,N_3226);
xor U3825 (N_3825,N_3264,N_3292);
nand U3826 (N_3826,N_3459,N_3558);
nor U3827 (N_3827,N_3297,N_3594);
xor U3828 (N_3828,N_3479,N_3285);
xor U3829 (N_3829,N_3425,N_3208);
or U3830 (N_3830,N_3218,N_3563);
nand U3831 (N_3831,N_3394,N_3248);
nor U3832 (N_3832,N_3202,N_3295);
nor U3833 (N_3833,N_3229,N_3562);
nor U3834 (N_3834,N_3541,N_3576);
nand U3835 (N_3835,N_3300,N_3279);
nor U3836 (N_3836,N_3543,N_3438);
and U3837 (N_3837,N_3577,N_3370);
and U3838 (N_3838,N_3247,N_3250);
nor U3839 (N_3839,N_3413,N_3450);
nor U3840 (N_3840,N_3497,N_3366);
nand U3841 (N_3841,N_3225,N_3592);
xor U3842 (N_3842,N_3480,N_3455);
and U3843 (N_3843,N_3378,N_3493);
nor U3844 (N_3844,N_3354,N_3357);
or U3845 (N_3845,N_3516,N_3243);
nand U3846 (N_3846,N_3241,N_3306);
xnor U3847 (N_3847,N_3353,N_3242);
xor U3848 (N_3848,N_3373,N_3441);
and U3849 (N_3849,N_3541,N_3547);
and U3850 (N_3850,N_3250,N_3551);
nor U3851 (N_3851,N_3499,N_3567);
and U3852 (N_3852,N_3357,N_3579);
xnor U3853 (N_3853,N_3559,N_3400);
nand U3854 (N_3854,N_3592,N_3387);
xnor U3855 (N_3855,N_3249,N_3285);
xor U3856 (N_3856,N_3200,N_3387);
nor U3857 (N_3857,N_3263,N_3579);
and U3858 (N_3858,N_3437,N_3405);
nor U3859 (N_3859,N_3413,N_3425);
xor U3860 (N_3860,N_3380,N_3451);
nor U3861 (N_3861,N_3435,N_3391);
xnor U3862 (N_3862,N_3378,N_3570);
and U3863 (N_3863,N_3589,N_3323);
and U3864 (N_3864,N_3489,N_3466);
nand U3865 (N_3865,N_3433,N_3497);
nor U3866 (N_3866,N_3227,N_3203);
nand U3867 (N_3867,N_3334,N_3217);
nor U3868 (N_3868,N_3291,N_3545);
xnor U3869 (N_3869,N_3578,N_3568);
and U3870 (N_3870,N_3338,N_3414);
nand U3871 (N_3871,N_3550,N_3409);
nor U3872 (N_3872,N_3281,N_3476);
and U3873 (N_3873,N_3567,N_3576);
nand U3874 (N_3874,N_3473,N_3267);
nor U3875 (N_3875,N_3244,N_3266);
and U3876 (N_3876,N_3239,N_3508);
nor U3877 (N_3877,N_3481,N_3457);
xor U3878 (N_3878,N_3316,N_3425);
or U3879 (N_3879,N_3572,N_3557);
xnor U3880 (N_3880,N_3588,N_3287);
nand U3881 (N_3881,N_3209,N_3294);
nor U3882 (N_3882,N_3298,N_3571);
and U3883 (N_3883,N_3580,N_3300);
nand U3884 (N_3884,N_3576,N_3271);
and U3885 (N_3885,N_3515,N_3312);
or U3886 (N_3886,N_3410,N_3552);
nand U3887 (N_3887,N_3499,N_3271);
and U3888 (N_3888,N_3404,N_3320);
nor U3889 (N_3889,N_3414,N_3394);
xor U3890 (N_3890,N_3529,N_3549);
nand U3891 (N_3891,N_3534,N_3256);
and U3892 (N_3892,N_3572,N_3291);
nor U3893 (N_3893,N_3295,N_3205);
and U3894 (N_3894,N_3575,N_3558);
xnor U3895 (N_3895,N_3527,N_3372);
and U3896 (N_3896,N_3400,N_3502);
and U3897 (N_3897,N_3562,N_3504);
nand U3898 (N_3898,N_3364,N_3353);
nand U3899 (N_3899,N_3498,N_3521);
and U3900 (N_3900,N_3501,N_3589);
nor U3901 (N_3901,N_3294,N_3382);
nor U3902 (N_3902,N_3504,N_3499);
or U3903 (N_3903,N_3510,N_3504);
xor U3904 (N_3904,N_3415,N_3227);
xor U3905 (N_3905,N_3474,N_3216);
nand U3906 (N_3906,N_3362,N_3405);
and U3907 (N_3907,N_3375,N_3274);
nand U3908 (N_3908,N_3351,N_3430);
nor U3909 (N_3909,N_3333,N_3428);
xnor U3910 (N_3910,N_3225,N_3345);
nand U3911 (N_3911,N_3321,N_3228);
or U3912 (N_3912,N_3320,N_3299);
xnor U3913 (N_3913,N_3331,N_3531);
xnor U3914 (N_3914,N_3411,N_3290);
or U3915 (N_3915,N_3341,N_3326);
nor U3916 (N_3916,N_3257,N_3340);
xnor U3917 (N_3917,N_3549,N_3396);
nand U3918 (N_3918,N_3507,N_3502);
xor U3919 (N_3919,N_3462,N_3584);
or U3920 (N_3920,N_3482,N_3500);
nor U3921 (N_3921,N_3543,N_3420);
xor U3922 (N_3922,N_3210,N_3426);
nor U3923 (N_3923,N_3204,N_3248);
nand U3924 (N_3924,N_3304,N_3490);
nand U3925 (N_3925,N_3522,N_3542);
nor U3926 (N_3926,N_3210,N_3340);
nor U3927 (N_3927,N_3492,N_3482);
nand U3928 (N_3928,N_3265,N_3286);
and U3929 (N_3929,N_3583,N_3387);
nor U3930 (N_3930,N_3327,N_3456);
xnor U3931 (N_3931,N_3323,N_3283);
and U3932 (N_3932,N_3212,N_3371);
nand U3933 (N_3933,N_3503,N_3452);
xnor U3934 (N_3934,N_3389,N_3461);
nor U3935 (N_3935,N_3370,N_3465);
nor U3936 (N_3936,N_3349,N_3441);
xor U3937 (N_3937,N_3254,N_3432);
nor U3938 (N_3938,N_3494,N_3439);
nor U3939 (N_3939,N_3326,N_3375);
and U3940 (N_3940,N_3515,N_3359);
nor U3941 (N_3941,N_3597,N_3225);
nor U3942 (N_3942,N_3338,N_3306);
nand U3943 (N_3943,N_3547,N_3456);
xor U3944 (N_3944,N_3538,N_3599);
xnor U3945 (N_3945,N_3427,N_3263);
xor U3946 (N_3946,N_3442,N_3580);
or U3947 (N_3947,N_3460,N_3503);
or U3948 (N_3948,N_3469,N_3327);
xor U3949 (N_3949,N_3407,N_3431);
nor U3950 (N_3950,N_3355,N_3235);
nor U3951 (N_3951,N_3344,N_3342);
nor U3952 (N_3952,N_3537,N_3395);
nor U3953 (N_3953,N_3530,N_3357);
nor U3954 (N_3954,N_3576,N_3590);
nand U3955 (N_3955,N_3427,N_3567);
nand U3956 (N_3956,N_3426,N_3364);
xor U3957 (N_3957,N_3591,N_3479);
and U3958 (N_3958,N_3213,N_3583);
xor U3959 (N_3959,N_3278,N_3492);
nand U3960 (N_3960,N_3237,N_3511);
xor U3961 (N_3961,N_3406,N_3564);
or U3962 (N_3962,N_3312,N_3330);
and U3963 (N_3963,N_3533,N_3530);
nand U3964 (N_3964,N_3241,N_3210);
nand U3965 (N_3965,N_3390,N_3320);
xnor U3966 (N_3966,N_3247,N_3395);
nand U3967 (N_3967,N_3235,N_3222);
xnor U3968 (N_3968,N_3202,N_3542);
nor U3969 (N_3969,N_3324,N_3203);
xor U3970 (N_3970,N_3355,N_3414);
xnor U3971 (N_3971,N_3272,N_3513);
xor U3972 (N_3972,N_3512,N_3542);
nand U3973 (N_3973,N_3273,N_3422);
nor U3974 (N_3974,N_3266,N_3506);
and U3975 (N_3975,N_3257,N_3442);
nand U3976 (N_3976,N_3531,N_3559);
and U3977 (N_3977,N_3353,N_3371);
or U3978 (N_3978,N_3422,N_3316);
and U3979 (N_3979,N_3226,N_3476);
xor U3980 (N_3980,N_3478,N_3243);
xnor U3981 (N_3981,N_3277,N_3202);
nand U3982 (N_3982,N_3305,N_3398);
or U3983 (N_3983,N_3453,N_3426);
or U3984 (N_3984,N_3577,N_3531);
or U3985 (N_3985,N_3543,N_3381);
and U3986 (N_3986,N_3543,N_3340);
xnor U3987 (N_3987,N_3228,N_3360);
xor U3988 (N_3988,N_3315,N_3454);
nor U3989 (N_3989,N_3541,N_3278);
xor U3990 (N_3990,N_3218,N_3385);
and U3991 (N_3991,N_3420,N_3287);
and U3992 (N_3992,N_3493,N_3477);
nand U3993 (N_3993,N_3436,N_3402);
and U3994 (N_3994,N_3481,N_3351);
nor U3995 (N_3995,N_3276,N_3485);
xor U3996 (N_3996,N_3268,N_3224);
xnor U3997 (N_3997,N_3423,N_3432);
nand U3998 (N_3998,N_3351,N_3313);
nand U3999 (N_3999,N_3275,N_3420);
nor U4000 (N_4000,N_3998,N_3766);
nand U4001 (N_4001,N_3620,N_3967);
nor U4002 (N_4002,N_3630,N_3736);
nor U4003 (N_4003,N_3695,N_3876);
nor U4004 (N_4004,N_3678,N_3790);
or U4005 (N_4005,N_3710,N_3794);
nor U4006 (N_4006,N_3791,N_3759);
nand U4007 (N_4007,N_3731,N_3920);
nand U4008 (N_4008,N_3768,N_3901);
or U4009 (N_4009,N_3732,N_3744);
or U4010 (N_4010,N_3764,N_3714);
xnor U4011 (N_4011,N_3979,N_3934);
and U4012 (N_4012,N_3716,N_3978);
or U4013 (N_4013,N_3958,N_3772);
nor U4014 (N_4014,N_3624,N_3812);
nor U4015 (N_4015,N_3820,N_3773);
nand U4016 (N_4016,N_3634,N_3676);
or U4017 (N_4017,N_3826,N_3842);
or U4018 (N_4018,N_3646,N_3844);
xnor U4019 (N_4019,N_3757,N_3957);
and U4020 (N_4020,N_3751,N_3765);
or U4021 (N_4021,N_3788,N_3718);
or U4022 (N_4022,N_3940,N_3739);
and U4023 (N_4023,N_3699,N_3662);
nor U4024 (N_4024,N_3918,N_3670);
or U4025 (N_4025,N_3825,N_3995);
or U4026 (N_4026,N_3947,N_3830);
nor U4027 (N_4027,N_3864,N_3980);
nand U4028 (N_4028,N_3805,N_3707);
and U4029 (N_4029,N_3720,N_3902);
and U4030 (N_4030,N_3972,N_3898);
xor U4031 (N_4031,N_3832,N_3996);
xnor U4032 (N_4032,N_3722,N_3660);
nand U4033 (N_4033,N_3908,N_3991);
or U4034 (N_4034,N_3795,N_3677);
nor U4035 (N_4035,N_3627,N_3784);
xor U4036 (N_4036,N_3877,N_3916);
nor U4037 (N_4037,N_3614,N_3973);
nor U4038 (N_4038,N_3692,N_3917);
nand U4039 (N_4039,N_3760,N_3609);
xnor U4040 (N_4040,N_3897,N_3645);
or U4041 (N_4041,N_3910,N_3850);
xnor U4042 (N_4042,N_3890,N_3956);
nand U4043 (N_4043,N_3709,N_3868);
nor U4044 (N_4044,N_3671,N_3623);
nor U4045 (N_4045,N_3726,N_3813);
nand U4046 (N_4046,N_3762,N_3841);
and U4047 (N_4047,N_3912,N_3665);
nand U4048 (N_4048,N_3892,N_3961);
or U4049 (N_4049,N_3666,N_3929);
nand U4050 (N_4050,N_3778,N_3856);
xnor U4051 (N_4051,N_3885,N_3834);
and U4052 (N_4052,N_3769,N_3811);
or U4053 (N_4053,N_3690,N_3870);
or U4054 (N_4054,N_3938,N_3983);
nand U4055 (N_4055,N_3734,N_3779);
xnor U4056 (N_4056,N_3700,N_3633);
or U4057 (N_4057,N_3982,N_3818);
and U4058 (N_4058,N_3889,N_3713);
and U4059 (N_4059,N_3796,N_3933);
or U4060 (N_4060,N_3988,N_3968);
nor U4061 (N_4061,N_3984,N_3786);
xor U4062 (N_4062,N_3815,N_3840);
nor U4063 (N_4063,N_3987,N_3895);
nor U4064 (N_4064,N_3869,N_3638);
and U4065 (N_4065,N_3730,N_3954);
and U4066 (N_4066,N_3680,N_3655);
xor U4067 (N_4067,N_3867,N_3833);
xor U4068 (N_4068,N_3927,N_3715);
xnor U4069 (N_4069,N_3611,N_3770);
nand U4070 (N_4070,N_3637,N_3792);
and U4071 (N_4071,N_3628,N_3802);
and U4072 (N_4072,N_3915,N_3740);
nand U4073 (N_4073,N_3657,N_3746);
nor U4074 (N_4074,N_3674,N_3724);
xnor U4075 (N_4075,N_3619,N_3754);
and U4076 (N_4076,N_3752,N_3787);
nor U4077 (N_4077,N_3774,N_3851);
or U4078 (N_4078,N_3937,N_3652);
and U4079 (N_4079,N_3650,N_3610);
xnor U4080 (N_4080,N_3992,N_3635);
nor U4081 (N_4081,N_3985,N_3862);
xnor U4082 (N_4082,N_3753,N_3741);
nand U4083 (N_4083,N_3697,N_3946);
or U4084 (N_4084,N_3698,N_3617);
and U4085 (N_4085,N_3612,N_3661);
nor U4086 (N_4086,N_3749,N_3807);
and U4087 (N_4087,N_3879,N_3828);
nor U4088 (N_4088,N_3848,N_3639);
xor U4089 (N_4089,N_3675,N_3643);
xor U4090 (N_4090,N_3663,N_3600);
nand U4091 (N_4091,N_3691,N_3816);
or U4092 (N_4092,N_3857,N_3728);
or U4093 (N_4093,N_3880,N_3944);
or U4094 (N_4094,N_3919,N_3603);
nor U4095 (N_4095,N_3893,N_3648);
or U4096 (N_4096,N_3706,N_3903);
nor U4097 (N_4097,N_3758,N_3939);
nor U4098 (N_4098,N_3708,N_3642);
xor U4099 (N_4099,N_3970,N_3763);
nor U4100 (N_4100,N_3785,N_3681);
xnor U4101 (N_4101,N_3965,N_3836);
nor U4102 (N_4102,N_3845,N_3647);
and U4103 (N_4103,N_3964,N_3953);
or U4104 (N_4104,N_3977,N_3814);
xnor U4105 (N_4105,N_3928,N_3911);
nor U4106 (N_4106,N_3727,N_3994);
nand U4107 (N_4107,N_3969,N_3712);
and U4108 (N_4108,N_3819,N_3997);
xnor U4109 (N_4109,N_3951,N_3881);
nor U4110 (N_4110,N_3952,N_3705);
and U4111 (N_4111,N_3669,N_3748);
and U4112 (N_4112,N_3673,N_3887);
nor U4113 (N_4113,N_3866,N_3755);
and U4114 (N_4114,N_3689,N_3914);
xor U4115 (N_4115,N_3629,N_3606);
nor U4116 (N_4116,N_3602,N_3899);
nor U4117 (N_4117,N_3960,N_3906);
or U4118 (N_4118,N_3696,N_3641);
and U4119 (N_4119,N_3658,N_3668);
xor U4120 (N_4120,N_3798,N_3806);
or U4121 (N_4121,N_3761,N_3835);
nor U4122 (N_4122,N_3839,N_3990);
nor U4123 (N_4123,N_3821,N_3687);
nor U4124 (N_4124,N_3659,N_3863);
or U4125 (N_4125,N_3962,N_3789);
xnor U4126 (N_4126,N_3966,N_3923);
and U4127 (N_4127,N_3986,N_3745);
nor U4128 (N_4128,N_3808,N_3809);
or U4129 (N_4129,N_3948,N_3604);
and U4130 (N_4130,N_3683,N_3804);
xnor U4131 (N_4131,N_3874,N_3636);
or U4132 (N_4132,N_3618,N_3613);
nor U4133 (N_4133,N_3737,N_3883);
xnor U4134 (N_4134,N_3651,N_3823);
nor U4135 (N_4135,N_3871,N_3931);
nand U4136 (N_4136,N_3608,N_3971);
nand U4137 (N_4137,N_3781,N_3886);
and U4138 (N_4138,N_3631,N_3626);
or U4139 (N_4139,N_3865,N_3756);
nor U4140 (N_4140,N_3838,N_3905);
or U4141 (N_4141,N_3738,N_3654);
nand U4142 (N_4142,N_3858,N_3777);
and U4143 (N_4143,N_3943,N_3974);
and U4144 (N_4144,N_3601,N_3801);
nand U4145 (N_4145,N_3733,N_3776);
nand U4146 (N_4146,N_3913,N_3930);
nor U4147 (N_4147,N_3797,N_3959);
nand U4148 (N_4148,N_3704,N_3942);
or U4149 (N_4149,N_3605,N_3932);
xnor U4150 (N_4150,N_3743,N_3843);
or U4151 (N_4151,N_3672,N_3803);
or U4152 (N_4152,N_3847,N_3644);
nand U4153 (N_4153,N_3949,N_3831);
and U4154 (N_4154,N_3701,N_3653);
or U4155 (N_4155,N_3615,N_3775);
nor U4156 (N_4156,N_3780,N_3926);
or U4157 (N_4157,N_3719,N_3860);
or U4158 (N_4158,N_3729,N_3925);
xnor U4159 (N_4159,N_3694,N_3935);
xnor U4160 (N_4160,N_3896,N_3684);
nor U4161 (N_4161,N_3667,N_3649);
and U4162 (N_4162,N_3922,N_3685);
xor U4163 (N_4163,N_3747,N_3829);
xor U4164 (N_4164,N_3625,N_3861);
or U4165 (N_4165,N_3981,N_3855);
nand U4166 (N_4166,N_3771,N_3621);
and U4167 (N_4167,N_3783,N_3999);
and U4168 (N_4168,N_3664,N_3921);
or U4169 (N_4169,N_3799,N_3872);
nor U4170 (N_4170,N_3742,N_3686);
and U4171 (N_4171,N_3976,N_3993);
and U4172 (N_4172,N_3725,N_3616);
xor U4173 (N_4173,N_3875,N_3682);
nor U4174 (N_4174,N_3882,N_3884);
and U4175 (N_4175,N_3817,N_3924);
xor U4176 (N_4176,N_3767,N_3793);
or U4177 (N_4177,N_3800,N_3703);
and U4178 (N_4178,N_3936,N_3632);
nor U4179 (N_4179,N_3782,N_3656);
and U4180 (N_4180,N_3975,N_3735);
nor U4181 (N_4181,N_3950,N_3622);
or U4182 (N_4182,N_3854,N_3852);
and U4183 (N_4183,N_3989,N_3750);
xor U4184 (N_4184,N_3878,N_3810);
nor U4185 (N_4185,N_3907,N_3904);
and U4186 (N_4186,N_3837,N_3900);
nor U4187 (N_4187,N_3822,N_3909);
or U4188 (N_4188,N_3891,N_3717);
or U4189 (N_4189,N_3702,N_3894);
or U4190 (N_4190,N_3945,N_3873);
nand U4191 (N_4191,N_3853,N_3849);
or U4192 (N_4192,N_3693,N_3888);
or U4193 (N_4193,N_3846,N_3688);
or U4194 (N_4194,N_3640,N_3941);
and U4195 (N_4195,N_3963,N_3723);
and U4196 (N_4196,N_3711,N_3721);
and U4197 (N_4197,N_3824,N_3679);
xor U4198 (N_4198,N_3859,N_3955);
nand U4199 (N_4199,N_3827,N_3607);
xnor U4200 (N_4200,N_3779,N_3750);
and U4201 (N_4201,N_3963,N_3865);
nand U4202 (N_4202,N_3777,N_3653);
nor U4203 (N_4203,N_3971,N_3840);
xor U4204 (N_4204,N_3908,N_3735);
nand U4205 (N_4205,N_3691,N_3855);
and U4206 (N_4206,N_3975,N_3952);
or U4207 (N_4207,N_3758,N_3668);
xor U4208 (N_4208,N_3629,N_3935);
xnor U4209 (N_4209,N_3951,N_3798);
or U4210 (N_4210,N_3970,N_3684);
and U4211 (N_4211,N_3618,N_3875);
or U4212 (N_4212,N_3862,N_3620);
and U4213 (N_4213,N_3998,N_3738);
or U4214 (N_4214,N_3907,N_3931);
nand U4215 (N_4215,N_3648,N_3800);
or U4216 (N_4216,N_3777,N_3908);
nor U4217 (N_4217,N_3734,N_3772);
and U4218 (N_4218,N_3638,N_3923);
nor U4219 (N_4219,N_3921,N_3918);
or U4220 (N_4220,N_3733,N_3975);
or U4221 (N_4221,N_3740,N_3865);
xnor U4222 (N_4222,N_3628,N_3745);
nand U4223 (N_4223,N_3994,N_3831);
nor U4224 (N_4224,N_3822,N_3717);
nor U4225 (N_4225,N_3922,N_3660);
xor U4226 (N_4226,N_3792,N_3665);
and U4227 (N_4227,N_3869,N_3771);
nand U4228 (N_4228,N_3891,N_3723);
xnor U4229 (N_4229,N_3689,N_3737);
and U4230 (N_4230,N_3826,N_3787);
or U4231 (N_4231,N_3610,N_3777);
nand U4232 (N_4232,N_3699,N_3942);
nor U4233 (N_4233,N_3805,N_3823);
nor U4234 (N_4234,N_3887,N_3718);
nand U4235 (N_4235,N_3811,N_3627);
xnor U4236 (N_4236,N_3817,N_3739);
xor U4237 (N_4237,N_3909,N_3660);
nand U4238 (N_4238,N_3855,N_3766);
nor U4239 (N_4239,N_3890,N_3840);
xor U4240 (N_4240,N_3686,N_3677);
nor U4241 (N_4241,N_3891,N_3781);
or U4242 (N_4242,N_3760,N_3971);
nand U4243 (N_4243,N_3869,N_3714);
or U4244 (N_4244,N_3993,N_3808);
xor U4245 (N_4245,N_3689,N_3975);
and U4246 (N_4246,N_3968,N_3679);
nor U4247 (N_4247,N_3720,N_3787);
or U4248 (N_4248,N_3847,N_3630);
and U4249 (N_4249,N_3697,N_3680);
or U4250 (N_4250,N_3907,N_3786);
nor U4251 (N_4251,N_3782,N_3681);
nand U4252 (N_4252,N_3854,N_3868);
and U4253 (N_4253,N_3632,N_3613);
or U4254 (N_4254,N_3793,N_3613);
xnor U4255 (N_4255,N_3779,N_3884);
nor U4256 (N_4256,N_3971,N_3614);
xor U4257 (N_4257,N_3987,N_3747);
nand U4258 (N_4258,N_3954,N_3964);
or U4259 (N_4259,N_3930,N_3925);
nor U4260 (N_4260,N_3994,N_3698);
or U4261 (N_4261,N_3862,N_3693);
nand U4262 (N_4262,N_3795,N_3988);
nor U4263 (N_4263,N_3836,N_3772);
xor U4264 (N_4264,N_3997,N_3634);
nand U4265 (N_4265,N_3917,N_3946);
xor U4266 (N_4266,N_3845,N_3895);
nor U4267 (N_4267,N_3935,N_3852);
or U4268 (N_4268,N_3982,N_3762);
nor U4269 (N_4269,N_3790,N_3635);
nand U4270 (N_4270,N_3638,N_3994);
or U4271 (N_4271,N_3834,N_3738);
nor U4272 (N_4272,N_3878,N_3766);
xnor U4273 (N_4273,N_3859,N_3978);
nand U4274 (N_4274,N_3912,N_3717);
xnor U4275 (N_4275,N_3801,N_3805);
xor U4276 (N_4276,N_3841,N_3712);
and U4277 (N_4277,N_3964,N_3794);
nor U4278 (N_4278,N_3808,N_3709);
nand U4279 (N_4279,N_3807,N_3675);
or U4280 (N_4280,N_3830,N_3917);
nand U4281 (N_4281,N_3738,N_3976);
nand U4282 (N_4282,N_3897,N_3846);
or U4283 (N_4283,N_3689,N_3693);
xor U4284 (N_4284,N_3947,N_3872);
and U4285 (N_4285,N_3923,N_3683);
and U4286 (N_4286,N_3633,N_3719);
nor U4287 (N_4287,N_3714,N_3760);
xnor U4288 (N_4288,N_3774,N_3877);
or U4289 (N_4289,N_3662,N_3792);
nand U4290 (N_4290,N_3842,N_3998);
nor U4291 (N_4291,N_3689,N_3928);
and U4292 (N_4292,N_3922,N_3870);
and U4293 (N_4293,N_3992,N_3772);
nand U4294 (N_4294,N_3614,N_3768);
or U4295 (N_4295,N_3904,N_3621);
xor U4296 (N_4296,N_3847,N_3863);
and U4297 (N_4297,N_3867,N_3987);
nand U4298 (N_4298,N_3814,N_3935);
nand U4299 (N_4299,N_3971,N_3745);
and U4300 (N_4300,N_3934,N_3709);
xor U4301 (N_4301,N_3820,N_3908);
xor U4302 (N_4302,N_3778,N_3854);
nor U4303 (N_4303,N_3746,N_3747);
nor U4304 (N_4304,N_3625,N_3885);
nor U4305 (N_4305,N_3690,N_3831);
xnor U4306 (N_4306,N_3738,N_3902);
xnor U4307 (N_4307,N_3809,N_3637);
xor U4308 (N_4308,N_3666,N_3763);
and U4309 (N_4309,N_3870,N_3831);
nor U4310 (N_4310,N_3835,N_3858);
xnor U4311 (N_4311,N_3665,N_3964);
or U4312 (N_4312,N_3849,N_3973);
or U4313 (N_4313,N_3721,N_3880);
xnor U4314 (N_4314,N_3983,N_3942);
nor U4315 (N_4315,N_3820,N_3848);
nand U4316 (N_4316,N_3910,N_3715);
xnor U4317 (N_4317,N_3680,N_3710);
nand U4318 (N_4318,N_3910,N_3932);
xnor U4319 (N_4319,N_3750,N_3602);
nand U4320 (N_4320,N_3983,N_3842);
nor U4321 (N_4321,N_3668,N_3630);
nand U4322 (N_4322,N_3820,N_3782);
and U4323 (N_4323,N_3943,N_3659);
xnor U4324 (N_4324,N_3724,N_3610);
nand U4325 (N_4325,N_3690,N_3798);
or U4326 (N_4326,N_3875,N_3850);
nand U4327 (N_4327,N_3667,N_3925);
nor U4328 (N_4328,N_3780,N_3742);
xnor U4329 (N_4329,N_3687,N_3816);
nor U4330 (N_4330,N_3896,N_3747);
nand U4331 (N_4331,N_3611,N_3814);
xor U4332 (N_4332,N_3798,N_3976);
and U4333 (N_4333,N_3778,N_3994);
nor U4334 (N_4334,N_3809,N_3702);
nand U4335 (N_4335,N_3929,N_3828);
nor U4336 (N_4336,N_3696,N_3871);
nor U4337 (N_4337,N_3942,N_3729);
nor U4338 (N_4338,N_3753,N_3708);
xnor U4339 (N_4339,N_3799,N_3935);
nand U4340 (N_4340,N_3837,N_3799);
or U4341 (N_4341,N_3866,N_3657);
or U4342 (N_4342,N_3865,N_3767);
and U4343 (N_4343,N_3876,N_3942);
nand U4344 (N_4344,N_3606,N_3892);
nor U4345 (N_4345,N_3893,N_3746);
nand U4346 (N_4346,N_3725,N_3617);
nor U4347 (N_4347,N_3688,N_3887);
and U4348 (N_4348,N_3649,N_3764);
or U4349 (N_4349,N_3753,N_3964);
and U4350 (N_4350,N_3840,N_3704);
nand U4351 (N_4351,N_3694,N_3607);
nand U4352 (N_4352,N_3938,N_3948);
or U4353 (N_4353,N_3733,N_3713);
nand U4354 (N_4354,N_3830,N_3874);
nand U4355 (N_4355,N_3989,N_3751);
nand U4356 (N_4356,N_3989,N_3637);
and U4357 (N_4357,N_3768,N_3823);
and U4358 (N_4358,N_3628,N_3612);
or U4359 (N_4359,N_3735,N_3945);
xnor U4360 (N_4360,N_3777,N_3971);
xnor U4361 (N_4361,N_3920,N_3753);
or U4362 (N_4362,N_3943,N_3627);
xor U4363 (N_4363,N_3983,N_3911);
nand U4364 (N_4364,N_3959,N_3771);
or U4365 (N_4365,N_3990,N_3819);
xor U4366 (N_4366,N_3796,N_3866);
or U4367 (N_4367,N_3855,N_3674);
xor U4368 (N_4368,N_3609,N_3796);
or U4369 (N_4369,N_3703,N_3746);
nand U4370 (N_4370,N_3722,N_3709);
xor U4371 (N_4371,N_3715,N_3934);
and U4372 (N_4372,N_3835,N_3995);
or U4373 (N_4373,N_3786,N_3785);
nand U4374 (N_4374,N_3971,N_3677);
and U4375 (N_4375,N_3934,N_3923);
xor U4376 (N_4376,N_3970,N_3691);
or U4377 (N_4377,N_3717,N_3698);
or U4378 (N_4378,N_3737,N_3775);
nand U4379 (N_4379,N_3812,N_3982);
nor U4380 (N_4380,N_3617,N_3768);
nand U4381 (N_4381,N_3785,N_3617);
and U4382 (N_4382,N_3842,N_3944);
and U4383 (N_4383,N_3691,N_3853);
or U4384 (N_4384,N_3733,N_3954);
nand U4385 (N_4385,N_3943,N_3892);
nor U4386 (N_4386,N_3659,N_3872);
and U4387 (N_4387,N_3766,N_3864);
xnor U4388 (N_4388,N_3914,N_3923);
or U4389 (N_4389,N_3900,N_3778);
nand U4390 (N_4390,N_3933,N_3769);
or U4391 (N_4391,N_3911,N_3772);
or U4392 (N_4392,N_3603,N_3872);
nand U4393 (N_4393,N_3672,N_3888);
xnor U4394 (N_4394,N_3817,N_3891);
nand U4395 (N_4395,N_3672,N_3873);
and U4396 (N_4396,N_3883,N_3924);
and U4397 (N_4397,N_3859,N_3948);
xnor U4398 (N_4398,N_3712,N_3718);
or U4399 (N_4399,N_3852,N_3657);
nor U4400 (N_4400,N_4123,N_4073);
xnor U4401 (N_4401,N_4204,N_4191);
and U4402 (N_4402,N_4292,N_4169);
or U4403 (N_4403,N_4274,N_4235);
nand U4404 (N_4404,N_4190,N_4384);
xnor U4405 (N_4405,N_4091,N_4245);
or U4406 (N_4406,N_4026,N_4134);
xor U4407 (N_4407,N_4342,N_4087);
and U4408 (N_4408,N_4156,N_4119);
nor U4409 (N_4409,N_4339,N_4271);
and U4410 (N_4410,N_4221,N_4198);
xnor U4411 (N_4411,N_4286,N_4149);
xnor U4412 (N_4412,N_4177,N_4267);
xor U4413 (N_4413,N_4047,N_4366);
nor U4414 (N_4414,N_4324,N_4142);
and U4415 (N_4415,N_4193,N_4275);
and U4416 (N_4416,N_4021,N_4211);
nor U4417 (N_4417,N_4037,N_4020);
nand U4418 (N_4418,N_4018,N_4337);
or U4419 (N_4419,N_4154,N_4290);
nor U4420 (N_4420,N_4242,N_4381);
or U4421 (N_4421,N_4048,N_4205);
nor U4422 (N_4422,N_4281,N_4196);
or U4423 (N_4423,N_4176,N_4171);
and U4424 (N_4424,N_4335,N_4078);
xor U4425 (N_4425,N_4210,N_4214);
and U4426 (N_4426,N_4302,N_4308);
nor U4427 (N_4427,N_4332,N_4365);
xor U4428 (N_4428,N_4028,N_4269);
or U4429 (N_4429,N_4257,N_4328);
or U4430 (N_4430,N_4092,N_4112);
xor U4431 (N_4431,N_4157,N_4340);
nand U4432 (N_4432,N_4170,N_4265);
and U4433 (N_4433,N_4166,N_4355);
xnor U4434 (N_4434,N_4317,N_4379);
nand U4435 (N_4435,N_4329,N_4293);
or U4436 (N_4436,N_4357,N_4122);
and U4437 (N_4437,N_4374,N_4377);
nand U4438 (N_4438,N_4255,N_4260);
nand U4439 (N_4439,N_4128,N_4225);
nor U4440 (N_4440,N_4007,N_4315);
nor U4441 (N_4441,N_4114,N_4129);
or U4442 (N_4442,N_4107,N_4035);
nand U4443 (N_4443,N_4354,N_4382);
nand U4444 (N_4444,N_4113,N_4179);
nor U4445 (N_4445,N_4227,N_4248);
xor U4446 (N_4446,N_4327,N_4015);
and U4447 (N_4447,N_4025,N_4017);
and U4448 (N_4448,N_4010,N_4059);
or U4449 (N_4449,N_4111,N_4163);
or U4450 (N_4450,N_4373,N_4061);
nor U4451 (N_4451,N_4124,N_4088);
and U4452 (N_4452,N_4361,N_4039);
xor U4453 (N_4453,N_4014,N_4063);
xnor U4454 (N_4454,N_4300,N_4385);
and U4455 (N_4455,N_4352,N_4116);
nor U4456 (N_4456,N_4239,N_4226);
nand U4457 (N_4457,N_4203,N_4273);
or U4458 (N_4458,N_4254,N_4282);
nor U4459 (N_4459,N_4206,N_4353);
xor U4460 (N_4460,N_4081,N_4053);
nand U4461 (N_4461,N_4098,N_4145);
or U4462 (N_4462,N_4362,N_4147);
or U4463 (N_4463,N_4049,N_4244);
nand U4464 (N_4464,N_4347,N_4238);
nand U4465 (N_4465,N_4234,N_4027);
nor U4466 (N_4466,N_4105,N_4005);
nand U4467 (N_4467,N_4256,N_4387);
xor U4468 (N_4468,N_4016,N_4033);
or U4469 (N_4469,N_4298,N_4000);
or U4470 (N_4470,N_4121,N_4249);
or U4471 (N_4471,N_4046,N_4164);
or U4472 (N_4472,N_4082,N_4294);
or U4473 (N_4473,N_4185,N_4189);
nand U4474 (N_4474,N_4133,N_4140);
and U4475 (N_4475,N_4022,N_4296);
or U4476 (N_4476,N_4085,N_4042);
xor U4477 (N_4477,N_4364,N_4303);
nand U4478 (N_4478,N_4103,N_4150);
and U4479 (N_4479,N_4371,N_4036);
or U4480 (N_4480,N_4330,N_4201);
or U4481 (N_4481,N_4218,N_4331);
or U4482 (N_4482,N_4029,N_4125);
and U4483 (N_4483,N_4104,N_4272);
or U4484 (N_4484,N_4158,N_4120);
nand U4485 (N_4485,N_4299,N_4212);
nand U4486 (N_4486,N_4322,N_4307);
and U4487 (N_4487,N_4376,N_4341);
xor U4488 (N_4488,N_4289,N_4208);
xnor U4489 (N_4489,N_4334,N_4323);
or U4490 (N_4490,N_4109,N_4174);
nor U4491 (N_4491,N_4052,N_4393);
and U4492 (N_4492,N_4161,N_4194);
nand U4493 (N_4493,N_4106,N_4181);
and U4494 (N_4494,N_4055,N_4146);
nor U4495 (N_4495,N_4222,N_4216);
and U4496 (N_4496,N_4153,N_4389);
xnor U4497 (N_4497,N_4396,N_4080);
xnor U4498 (N_4498,N_4162,N_4148);
nor U4499 (N_4499,N_4312,N_4251);
nand U4500 (N_4500,N_4001,N_4066);
or U4501 (N_4501,N_4187,N_4160);
or U4502 (N_4502,N_4363,N_4167);
xnor U4503 (N_4503,N_4350,N_4268);
or U4504 (N_4504,N_4011,N_4223);
and U4505 (N_4505,N_4285,N_4143);
nor U4506 (N_4506,N_4050,N_4057);
nand U4507 (N_4507,N_4391,N_4139);
or U4508 (N_4508,N_4084,N_4325);
nand U4509 (N_4509,N_4283,N_4338);
nand U4510 (N_4510,N_4390,N_4182);
and U4511 (N_4511,N_4388,N_4137);
or U4512 (N_4512,N_4392,N_4217);
nor U4513 (N_4513,N_4126,N_4310);
nor U4514 (N_4514,N_4056,N_4360);
xor U4515 (N_4515,N_4345,N_4183);
or U4516 (N_4516,N_4093,N_4110);
nand U4517 (N_4517,N_4266,N_4197);
and U4518 (N_4518,N_4200,N_4349);
nand U4519 (N_4519,N_4138,N_4368);
xnor U4520 (N_4520,N_4195,N_4395);
nand U4521 (N_4521,N_4358,N_4367);
or U4522 (N_4522,N_4030,N_4101);
nand U4523 (N_4523,N_4318,N_4241);
nor U4524 (N_4524,N_4250,N_4236);
nor U4525 (N_4525,N_4309,N_4165);
nor U4526 (N_4526,N_4263,N_4343);
nand U4527 (N_4527,N_4231,N_4279);
nand U4528 (N_4528,N_4058,N_4075);
xor U4529 (N_4529,N_4060,N_4144);
and U4530 (N_4530,N_4252,N_4253);
and U4531 (N_4531,N_4076,N_4288);
and U4532 (N_4532,N_4209,N_4024);
xor U4533 (N_4533,N_4168,N_4220);
xor U4534 (N_4534,N_4369,N_4259);
or U4535 (N_4535,N_4009,N_4213);
nand U4536 (N_4536,N_4192,N_4151);
nor U4537 (N_4537,N_4277,N_4013);
and U4538 (N_4538,N_4083,N_4270);
nor U4539 (N_4539,N_4043,N_4108);
nor U4540 (N_4540,N_4344,N_4135);
nor U4541 (N_4541,N_4321,N_4155);
xor U4542 (N_4542,N_4086,N_4115);
nor U4543 (N_4543,N_4316,N_4023);
xor U4544 (N_4544,N_4284,N_4247);
and U4545 (N_4545,N_4383,N_4090);
nand U4546 (N_4546,N_4258,N_4333);
xnor U4547 (N_4547,N_4041,N_4233);
xor U4548 (N_4548,N_4356,N_4032);
nor U4549 (N_4549,N_4399,N_4074);
nor U4550 (N_4550,N_4100,N_4054);
nand U4551 (N_4551,N_4261,N_4003);
nor U4552 (N_4552,N_4006,N_4243);
nand U4553 (N_4553,N_4240,N_4045);
or U4554 (N_4554,N_4040,N_4305);
and U4555 (N_4555,N_4178,N_4072);
or U4556 (N_4556,N_4351,N_4118);
and U4557 (N_4557,N_4172,N_4319);
or U4558 (N_4558,N_4065,N_4398);
xnor U4559 (N_4559,N_4008,N_4346);
nor U4560 (N_4560,N_4062,N_4099);
or U4561 (N_4561,N_4012,N_4068);
xor U4562 (N_4562,N_4287,N_4311);
and U4563 (N_4563,N_4199,N_4038);
xor U4564 (N_4564,N_4297,N_4394);
or U4565 (N_4565,N_4097,N_4291);
or U4566 (N_4566,N_4224,N_4102);
or U4567 (N_4567,N_4262,N_4127);
nor U4568 (N_4568,N_4246,N_4159);
or U4569 (N_4569,N_4348,N_4359);
nor U4570 (N_4570,N_4304,N_4370);
nand U4571 (N_4571,N_4077,N_4175);
nor U4572 (N_4572,N_4230,N_4079);
or U4573 (N_4573,N_4071,N_4219);
and U4574 (N_4574,N_4188,N_4131);
xnor U4575 (N_4575,N_4237,N_4044);
and U4576 (N_4576,N_4301,N_4180);
and U4577 (N_4577,N_4397,N_4152);
or U4578 (N_4578,N_4228,N_4207);
xnor U4579 (N_4579,N_4280,N_4031);
xor U4580 (N_4580,N_4141,N_4276);
nor U4581 (N_4581,N_4094,N_4136);
and U4582 (N_4582,N_4202,N_4264);
or U4583 (N_4583,N_4326,N_4320);
xnor U4584 (N_4584,N_4314,N_4336);
xor U4585 (N_4585,N_4173,N_4378);
and U4586 (N_4586,N_4278,N_4096);
or U4587 (N_4587,N_4386,N_4089);
and U4588 (N_4588,N_4019,N_4002);
xor U4589 (N_4589,N_4067,N_4295);
or U4590 (N_4590,N_4069,N_4004);
and U4591 (N_4591,N_4375,N_4070);
xor U4592 (N_4592,N_4380,N_4130);
or U4593 (N_4593,N_4064,N_4215);
nor U4594 (N_4594,N_4034,N_4184);
and U4595 (N_4595,N_4095,N_4232);
or U4596 (N_4596,N_4313,N_4132);
xnor U4597 (N_4597,N_4306,N_4117);
or U4598 (N_4598,N_4186,N_4372);
nor U4599 (N_4599,N_4229,N_4051);
nand U4600 (N_4600,N_4369,N_4169);
and U4601 (N_4601,N_4326,N_4270);
and U4602 (N_4602,N_4365,N_4213);
nor U4603 (N_4603,N_4162,N_4317);
or U4604 (N_4604,N_4307,N_4123);
or U4605 (N_4605,N_4354,N_4350);
or U4606 (N_4606,N_4239,N_4083);
and U4607 (N_4607,N_4237,N_4265);
xnor U4608 (N_4608,N_4211,N_4297);
nor U4609 (N_4609,N_4056,N_4030);
or U4610 (N_4610,N_4304,N_4150);
or U4611 (N_4611,N_4167,N_4200);
nor U4612 (N_4612,N_4002,N_4092);
nand U4613 (N_4613,N_4010,N_4340);
or U4614 (N_4614,N_4305,N_4117);
xnor U4615 (N_4615,N_4378,N_4092);
nor U4616 (N_4616,N_4162,N_4294);
or U4617 (N_4617,N_4150,N_4246);
and U4618 (N_4618,N_4090,N_4015);
nand U4619 (N_4619,N_4369,N_4364);
and U4620 (N_4620,N_4216,N_4070);
nand U4621 (N_4621,N_4363,N_4136);
nand U4622 (N_4622,N_4229,N_4213);
or U4623 (N_4623,N_4070,N_4276);
and U4624 (N_4624,N_4076,N_4184);
nand U4625 (N_4625,N_4195,N_4399);
or U4626 (N_4626,N_4213,N_4234);
nor U4627 (N_4627,N_4173,N_4105);
nor U4628 (N_4628,N_4028,N_4159);
nand U4629 (N_4629,N_4029,N_4199);
or U4630 (N_4630,N_4387,N_4371);
nor U4631 (N_4631,N_4351,N_4214);
nor U4632 (N_4632,N_4119,N_4178);
and U4633 (N_4633,N_4257,N_4264);
xor U4634 (N_4634,N_4151,N_4009);
and U4635 (N_4635,N_4007,N_4182);
and U4636 (N_4636,N_4307,N_4037);
nor U4637 (N_4637,N_4087,N_4246);
or U4638 (N_4638,N_4373,N_4031);
and U4639 (N_4639,N_4097,N_4371);
nor U4640 (N_4640,N_4264,N_4161);
or U4641 (N_4641,N_4157,N_4256);
nand U4642 (N_4642,N_4196,N_4000);
and U4643 (N_4643,N_4101,N_4315);
nand U4644 (N_4644,N_4086,N_4094);
nor U4645 (N_4645,N_4240,N_4298);
or U4646 (N_4646,N_4296,N_4061);
nand U4647 (N_4647,N_4260,N_4157);
nand U4648 (N_4648,N_4370,N_4274);
or U4649 (N_4649,N_4303,N_4361);
nand U4650 (N_4650,N_4195,N_4134);
or U4651 (N_4651,N_4169,N_4069);
and U4652 (N_4652,N_4065,N_4048);
and U4653 (N_4653,N_4226,N_4062);
or U4654 (N_4654,N_4086,N_4330);
xor U4655 (N_4655,N_4204,N_4219);
xnor U4656 (N_4656,N_4396,N_4384);
nand U4657 (N_4657,N_4293,N_4239);
nor U4658 (N_4658,N_4033,N_4000);
nand U4659 (N_4659,N_4392,N_4293);
or U4660 (N_4660,N_4192,N_4071);
or U4661 (N_4661,N_4396,N_4209);
xnor U4662 (N_4662,N_4191,N_4158);
or U4663 (N_4663,N_4113,N_4260);
nand U4664 (N_4664,N_4319,N_4001);
nor U4665 (N_4665,N_4000,N_4040);
xor U4666 (N_4666,N_4164,N_4109);
nor U4667 (N_4667,N_4200,N_4110);
or U4668 (N_4668,N_4094,N_4170);
xnor U4669 (N_4669,N_4178,N_4351);
nor U4670 (N_4670,N_4050,N_4210);
and U4671 (N_4671,N_4320,N_4100);
xnor U4672 (N_4672,N_4244,N_4354);
and U4673 (N_4673,N_4399,N_4141);
xor U4674 (N_4674,N_4091,N_4186);
nor U4675 (N_4675,N_4041,N_4185);
xor U4676 (N_4676,N_4063,N_4170);
or U4677 (N_4677,N_4066,N_4053);
nor U4678 (N_4678,N_4073,N_4362);
nor U4679 (N_4679,N_4072,N_4162);
nand U4680 (N_4680,N_4006,N_4070);
nor U4681 (N_4681,N_4347,N_4252);
xnor U4682 (N_4682,N_4151,N_4040);
nor U4683 (N_4683,N_4344,N_4114);
nor U4684 (N_4684,N_4053,N_4056);
nand U4685 (N_4685,N_4022,N_4016);
xor U4686 (N_4686,N_4223,N_4196);
and U4687 (N_4687,N_4394,N_4237);
xor U4688 (N_4688,N_4227,N_4371);
nand U4689 (N_4689,N_4001,N_4121);
xnor U4690 (N_4690,N_4362,N_4093);
xor U4691 (N_4691,N_4339,N_4346);
nand U4692 (N_4692,N_4394,N_4112);
and U4693 (N_4693,N_4315,N_4016);
xor U4694 (N_4694,N_4190,N_4350);
and U4695 (N_4695,N_4074,N_4048);
nand U4696 (N_4696,N_4107,N_4366);
nor U4697 (N_4697,N_4303,N_4043);
nand U4698 (N_4698,N_4147,N_4224);
or U4699 (N_4699,N_4274,N_4328);
nor U4700 (N_4700,N_4120,N_4176);
and U4701 (N_4701,N_4039,N_4073);
xor U4702 (N_4702,N_4331,N_4346);
nor U4703 (N_4703,N_4016,N_4059);
xnor U4704 (N_4704,N_4198,N_4054);
and U4705 (N_4705,N_4314,N_4109);
nand U4706 (N_4706,N_4116,N_4291);
nor U4707 (N_4707,N_4387,N_4217);
or U4708 (N_4708,N_4367,N_4148);
nor U4709 (N_4709,N_4246,N_4226);
and U4710 (N_4710,N_4093,N_4352);
xor U4711 (N_4711,N_4214,N_4386);
nor U4712 (N_4712,N_4290,N_4038);
and U4713 (N_4713,N_4297,N_4274);
and U4714 (N_4714,N_4079,N_4270);
and U4715 (N_4715,N_4125,N_4219);
or U4716 (N_4716,N_4015,N_4395);
nor U4717 (N_4717,N_4370,N_4076);
nand U4718 (N_4718,N_4050,N_4220);
nor U4719 (N_4719,N_4073,N_4019);
and U4720 (N_4720,N_4122,N_4043);
xor U4721 (N_4721,N_4243,N_4049);
nand U4722 (N_4722,N_4190,N_4202);
xor U4723 (N_4723,N_4080,N_4270);
nor U4724 (N_4724,N_4350,N_4077);
and U4725 (N_4725,N_4347,N_4300);
or U4726 (N_4726,N_4266,N_4229);
or U4727 (N_4727,N_4259,N_4268);
nor U4728 (N_4728,N_4166,N_4394);
nand U4729 (N_4729,N_4226,N_4170);
nor U4730 (N_4730,N_4202,N_4035);
nand U4731 (N_4731,N_4086,N_4238);
xnor U4732 (N_4732,N_4227,N_4223);
and U4733 (N_4733,N_4378,N_4153);
or U4734 (N_4734,N_4108,N_4147);
or U4735 (N_4735,N_4030,N_4367);
nand U4736 (N_4736,N_4201,N_4008);
nor U4737 (N_4737,N_4033,N_4119);
nand U4738 (N_4738,N_4224,N_4055);
nand U4739 (N_4739,N_4232,N_4043);
nor U4740 (N_4740,N_4325,N_4375);
nand U4741 (N_4741,N_4136,N_4317);
and U4742 (N_4742,N_4242,N_4278);
and U4743 (N_4743,N_4378,N_4199);
nor U4744 (N_4744,N_4140,N_4222);
or U4745 (N_4745,N_4388,N_4180);
or U4746 (N_4746,N_4011,N_4261);
nand U4747 (N_4747,N_4372,N_4241);
xor U4748 (N_4748,N_4230,N_4145);
and U4749 (N_4749,N_4303,N_4301);
nand U4750 (N_4750,N_4344,N_4017);
or U4751 (N_4751,N_4385,N_4290);
nor U4752 (N_4752,N_4144,N_4234);
and U4753 (N_4753,N_4358,N_4321);
nor U4754 (N_4754,N_4179,N_4002);
or U4755 (N_4755,N_4150,N_4228);
or U4756 (N_4756,N_4184,N_4397);
nor U4757 (N_4757,N_4352,N_4184);
and U4758 (N_4758,N_4020,N_4101);
nor U4759 (N_4759,N_4078,N_4383);
and U4760 (N_4760,N_4288,N_4005);
nand U4761 (N_4761,N_4048,N_4253);
nand U4762 (N_4762,N_4150,N_4356);
nand U4763 (N_4763,N_4091,N_4193);
nor U4764 (N_4764,N_4242,N_4311);
or U4765 (N_4765,N_4127,N_4197);
nor U4766 (N_4766,N_4073,N_4377);
nand U4767 (N_4767,N_4298,N_4246);
or U4768 (N_4768,N_4193,N_4081);
xor U4769 (N_4769,N_4210,N_4384);
xor U4770 (N_4770,N_4340,N_4266);
nand U4771 (N_4771,N_4083,N_4175);
nor U4772 (N_4772,N_4163,N_4236);
or U4773 (N_4773,N_4128,N_4042);
and U4774 (N_4774,N_4132,N_4035);
and U4775 (N_4775,N_4194,N_4124);
nand U4776 (N_4776,N_4031,N_4008);
xnor U4777 (N_4777,N_4090,N_4078);
and U4778 (N_4778,N_4255,N_4378);
xor U4779 (N_4779,N_4086,N_4163);
nor U4780 (N_4780,N_4022,N_4211);
xor U4781 (N_4781,N_4335,N_4048);
nand U4782 (N_4782,N_4093,N_4127);
nand U4783 (N_4783,N_4104,N_4234);
xnor U4784 (N_4784,N_4083,N_4298);
nand U4785 (N_4785,N_4051,N_4137);
nand U4786 (N_4786,N_4305,N_4362);
xnor U4787 (N_4787,N_4134,N_4038);
xor U4788 (N_4788,N_4082,N_4080);
and U4789 (N_4789,N_4104,N_4224);
nor U4790 (N_4790,N_4336,N_4287);
and U4791 (N_4791,N_4008,N_4087);
or U4792 (N_4792,N_4298,N_4097);
nand U4793 (N_4793,N_4240,N_4146);
or U4794 (N_4794,N_4346,N_4279);
nor U4795 (N_4795,N_4059,N_4035);
or U4796 (N_4796,N_4101,N_4003);
or U4797 (N_4797,N_4091,N_4259);
nor U4798 (N_4798,N_4242,N_4255);
or U4799 (N_4799,N_4252,N_4320);
nor U4800 (N_4800,N_4537,N_4402);
nor U4801 (N_4801,N_4531,N_4584);
and U4802 (N_4802,N_4629,N_4656);
or U4803 (N_4803,N_4796,N_4484);
nand U4804 (N_4804,N_4588,N_4503);
and U4805 (N_4805,N_4685,N_4785);
and U4806 (N_4806,N_4626,N_4706);
and U4807 (N_4807,N_4604,N_4623);
xnor U4808 (N_4808,N_4415,N_4699);
nand U4809 (N_4809,N_4433,N_4516);
or U4810 (N_4810,N_4659,N_4783);
xnor U4811 (N_4811,N_4747,N_4736);
xnor U4812 (N_4812,N_4671,N_4592);
or U4813 (N_4813,N_4709,N_4466);
nor U4814 (N_4814,N_4519,N_4478);
xnor U4815 (N_4815,N_4495,N_4674);
nand U4816 (N_4816,N_4406,N_4436);
nand U4817 (N_4817,N_4470,N_4493);
xnor U4818 (N_4818,N_4429,N_4556);
or U4819 (N_4819,N_4546,N_4549);
nand U4820 (N_4820,N_4514,N_4438);
nand U4821 (N_4821,N_4687,N_4780);
and U4822 (N_4822,N_4606,N_4455);
or U4823 (N_4823,N_4540,N_4536);
nor U4824 (N_4824,N_4797,N_4715);
nand U4825 (N_4825,N_4733,N_4424);
nand U4826 (N_4826,N_4748,N_4448);
nand U4827 (N_4827,N_4770,N_4467);
or U4828 (N_4828,N_4734,N_4427);
nand U4829 (N_4829,N_4670,N_4646);
or U4830 (N_4830,N_4459,N_4526);
or U4831 (N_4831,N_4698,N_4462);
nor U4832 (N_4832,N_4781,N_4614);
and U4833 (N_4833,N_4419,N_4430);
xor U4834 (N_4834,N_4653,N_4728);
nor U4835 (N_4835,N_4567,N_4724);
xnor U4836 (N_4836,N_4630,N_4764);
or U4837 (N_4837,N_4617,N_4644);
nand U4838 (N_4838,N_4517,N_4773);
or U4839 (N_4839,N_4663,N_4769);
and U4840 (N_4840,N_4654,N_4693);
and U4841 (N_4841,N_4635,N_4591);
xnor U4842 (N_4842,N_4515,N_4403);
and U4843 (N_4843,N_4413,N_4596);
nor U4844 (N_4844,N_4472,N_4689);
xor U4845 (N_4845,N_4662,N_4544);
xor U4846 (N_4846,N_4574,N_4759);
nand U4847 (N_4847,N_4795,N_4621);
xnor U4848 (N_4848,N_4707,N_4631);
nand U4849 (N_4849,N_4409,N_4624);
xor U4850 (N_4850,N_4774,N_4437);
xnor U4851 (N_4851,N_4502,N_4432);
or U4852 (N_4852,N_4586,N_4598);
xor U4853 (N_4853,N_4688,N_4739);
and U4854 (N_4854,N_4504,N_4562);
nor U4855 (N_4855,N_4593,N_4521);
xnor U4856 (N_4856,N_4657,N_4566);
nand U4857 (N_4857,N_4648,N_4690);
xnor U4858 (N_4858,N_4704,N_4440);
and U4859 (N_4859,N_4776,N_4771);
nor U4860 (N_4860,N_4702,N_4667);
xor U4861 (N_4861,N_4641,N_4552);
nand U4862 (N_4862,N_4603,N_4548);
xor U4863 (N_4863,N_4499,N_4420);
xnor U4864 (N_4864,N_4672,N_4608);
xor U4865 (N_4865,N_4425,N_4533);
or U4866 (N_4866,N_4510,N_4444);
nor U4867 (N_4867,N_4422,N_4511);
or U4868 (N_4868,N_4563,N_4465);
and U4869 (N_4869,N_4620,N_4611);
or U4870 (N_4870,N_4782,N_4528);
and U4871 (N_4871,N_4779,N_4730);
or U4872 (N_4872,N_4412,N_4692);
or U4873 (N_4873,N_4512,N_4453);
xor U4874 (N_4874,N_4754,N_4740);
nand U4875 (N_4875,N_4703,N_4579);
nor U4876 (N_4876,N_4560,N_4534);
nand U4877 (N_4877,N_4554,N_4557);
and U4878 (N_4878,N_4628,N_4778);
xor U4879 (N_4879,N_4655,N_4649);
or U4880 (N_4880,N_4650,N_4767);
xor U4881 (N_4881,N_4522,N_4445);
or U4882 (N_4882,N_4583,N_4542);
nor U4883 (N_4883,N_4460,N_4742);
or U4884 (N_4884,N_4675,N_4435);
nor U4885 (N_4885,N_4570,N_4575);
nand U4886 (N_4886,N_4483,N_4680);
and U4887 (N_4887,N_4716,N_4766);
and U4888 (N_4888,N_4523,N_4494);
or U4889 (N_4889,N_4463,N_4636);
nor U4890 (N_4890,N_4763,N_4558);
nor U4891 (N_4891,N_4561,N_4581);
and U4892 (N_4892,N_4505,N_4665);
nand U4893 (N_4893,N_4498,N_4696);
or U4894 (N_4894,N_4679,N_4513);
nand U4895 (N_4895,N_4551,N_4602);
nor U4896 (N_4896,N_4601,N_4666);
and U4897 (N_4897,N_4792,N_4589);
and U4898 (N_4898,N_4697,N_4594);
nor U4899 (N_4899,N_4597,N_4752);
or U4900 (N_4900,N_4652,N_4714);
nand U4901 (N_4901,N_4718,N_4788);
or U4902 (N_4902,N_4633,N_4743);
nor U4903 (N_4903,N_4417,N_4565);
and U4904 (N_4904,N_4684,N_4758);
nand U4905 (N_4905,N_4678,N_4447);
or U4906 (N_4906,N_4416,N_4789);
and U4907 (N_4907,N_4705,N_4725);
nor U4908 (N_4908,N_4737,N_4700);
nor U4909 (N_4909,N_4428,N_4553);
or U4910 (N_4910,N_4669,N_4787);
and U4911 (N_4911,N_4421,N_4410);
nor U4912 (N_4912,N_4691,N_4712);
or U4913 (N_4913,N_4547,N_4426);
nor U4914 (N_4914,N_4449,N_4423);
and U4915 (N_4915,N_4450,N_4527);
nor U4916 (N_4916,N_4580,N_4458);
nand U4917 (N_4917,N_4799,N_4468);
and U4918 (N_4918,N_4486,N_4695);
nor U4919 (N_4919,N_4744,N_4673);
or U4920 (N_4920,N_4474,N_4664);
xnor U4921 (N_4921,N_4480,N_4721);
and U4922 (N_4922,N_4595,N_4668);
or U4923 (N_4923,N_4681,N_4694);
or U4924 (N_4924,N_4590,N_4454);
or U4925 (N_4925,N_4572,N_4762);
xnor U4926 (N_4926,N_4701,N_4452);
nand U4927 (N_4927,N_4539,N_4755);
and U4928 (N_4928,N_4637,N_4622);
nor U4929 (N_4929,N_4461,N_4726);
nand U4930 (N_4930,N_4489,N_4405);
xnor U4931 (N_4931,N_4408,N_4757);
and U4932 (N_4932,N_4492,N_4543);
nand U4933 (N_4933,N_4686,N_4722);
nor U4934 (N_4934,N_4535,N_4576);
and U4935 (N_4935,N_4790,N_4645);
and U4936 (N_4936,N_4772,N_4711);
xor U4937 (N_4937,N_4497,N_4469);
nor U4938 (N_4938,N_4632,N_4569);
or U4939 (N_4939,N_4506,N_4634);
nand U4940 (N_4940,N_4676,N_4508);
and U4941 (N_4941,N_4476,N_4538);
and U4942 (N_4942,N_4488,N_4439);
nand U4943 (N_4943,N_4713,N_4609);
and U4944 (N_4944,N_4587,N_4477);
nand U4945 (N_4945,N_4451,N_4784);
and U4946 (N_4946,N_4793,N_4647);
nor U4947 (N_4947,N_4607,N_4509);
and U4948 (N_4948,N_4407,N_4446);
and U4949 (N_4949,N_4643,N_4442);
nand U4950 (N_4950,N_4525,N_4564);
nand U4951 (N_4951,N_4791,N_4616);
xnor U4952 (N_4952,N_4756,N_4431);
nand U4953 (N_4953,N_4582,N_4530);
or U4954 (N_4954,N_4500,N_4507);
xnor U4955 (N_4955,N_4418,N_4555);
and U4956 (N_4956,N_4717,N_4660);
or U4957 (N_4957,N_4559,N_4777);
and U4958 (N_4958,N_4571,N_4568);
nor U4959 (N_4959,N_4735,N_4414);
nand U4960 (N_4960,N_4481,N_4490);
nand U4961 (N_4961,N_4786,N_4751);
xor U4962 (N_4962,N_4750,N_4404);
or U4963 (N_4963,N_4677,N_4520);
nor U4964 (N_4964,N_4573,N_4610);
nor U4965 (N_4965,N_4727,N_4401);
nand U4966 (N_4966,N_4719,N_4487);
nor U4967 (N_4967,N_4471,N_4529);
and U4968 (N_4968,N_4794,N_4599);
xor U4969 (N_4969,N_4457,N_4798);
nand U4970 (N_4970,N_4491,N_4441);
or U4971 (N_4971,N_4639,N_4411);
or U4972 (N_4972,N_4753,N_4638);
nor U4973 (N_4973,N_4618,N_4485);
nor U4974 (N_4974,N_4746,N_4729);
and U4975 (N_4975,N_4640,N_4761);
nor U4976 (N_4976,N_4731,N_4464);
xor U4977 (N_4977,N_4745,N_4615);
and U4978 (N_4978,N_4578,N_4651);
or U4979 (N_4979,N_4585,N_4732);
xor U4980 (N_4980,N_4612,N_4456);
or U4981 (N_4981,N_4708,N_4738);
xnor U4982 (N_4982,N_4550,N_4768);
xnor U4983 (N_4983,N_4619,N_4479);
xor U4984 (N_4984,N_4658,N_4741);
and U4985 (N_4985,N_4473,N_4661);
nor U4986 (N_4986,N_4475,N_4524);
xnor U4987 (N_4987,N_4482,N_4600);
nor U4988 (N_4988,N_4760,N_4443);
and U4989 (N_4989,N_4710,N_4501);
xor U4990 (N_4990,N_4577,N_4541);
and U4991 (N_4991,N_4720,N_4496);
nor U4992 (N_4992,N_4434,N_4682);
and U4993 (N_4993,N_4605,N_4683);
xor U4994 (N_4994,N_4765,N_4749);
nor U4995 (N_4995,N_4775,N_4545);
or U4996 (N_4996,N_4613,N_4625);
and U4997 (N_4997,N_4642,N_4723);
nand U4998 (N_4998,N_4518,N_4627);
and U4999 (N_4999,N_4532,N_4400);
or U5000 (N_5000,N_4715,N_4613);
nand U5001 (N_5001,N_4756,N_4580);
and U5002 (N_5002,N_4506,N_4552);
xor U5003 (N_5003,N_4629,N_4531);
and U5004 (N_5004,N_4480,N_4720);
nor U5005 (N_5005,N_4460,N_4461);
xnor U5006 (N_5006,N_4630,N_4756);
nand U5007 (N_5007,N_4759,N_4756);
and U5008 (N_5008,N_4691,N_4548);
and U5009 (N_5009,N_4690,N_4462);
or U5010 (N_5010,N_4786,N_4525);
and U5011 (N_5011,N_4573,N_4684);
xnor U5012 (N_5012,N_4595,N_4559);
or U5013 (N_5013,N_4769,N_4799);
xor U5014 (N_5014,N_4571,N_4584);
or U5015 (N_5015,N_4479,N_4510);
nor U5016 (N_5016,N_4552,N_4587);
xnor U5017 (N_5017,N_4405,N_4654);
nor U5018 (N_5018,N_4729,N_4721);
nand U5019 (N_5019,N_4708,N_4432);
or U5020 (N_5020,N_4686,N_4576);
or U5021 (N_5021,N_4608,N_4668);
or U5022 (N_5022,N_4795,N_4606);
or U5023 (N_5023,N_4598,N_4745);
and U5024 (N_5024,N_4652,N_4441);
or U5025 (N_5025,N_4522,N_4426);
nand U5026 (N_5026,N_4653,N_4726);
nor U5027 (N_5027,N_4587,N_4701);
xor U5028 (N_5028,N_4582,N_4581);
and U5029 (N_5029,N_4490,N_4441);
nor U5030 (N_5030,N_4471,N_4741);
nand U5031 (N_5031,N_4714,N_4614);
nand U5032 (N_5032,N_4531,N_4648);
and U5033 (N_5033,N_4727,N_4560);
xor U5034 (N_5034,N_4699,N_4785);
nand U5035 (N_5035,N_4677,N_4627);
xor U5036 (N_5036,N_4735,N_4610);
nand U5037 (N_5037,N_4689,N_4454);
and U5038 (N_5038,N_4732,N_4638);
nor U5039 (N_5039,N_4440,N_4449);
xnor U5040 (N_5040,N_4519,N_4547);
nor U5041 (N_5041,N_4606,N_4755);
xnor U5042 (N_5042,N_4616,N_4545);
nor U5043 (N_5043,N_4768,N_4786);
or U5044 (N_5044,N_4541,N_4429);
xnor U5045 (N_5045,N_4400,N_4457);
nor U5046 (N_5046,N_4484,N_4641);
xor U5047 (N_5047,N_4670,N_4716);
and U5048 (N_5048,N_4688,N_4445);
nand U5049 (N_5049,N_4417,N_4746);
xnor U5050 (N_5050,N_4610,N_4619);
xnor U5051 (N_5051,N_4412,N_4462);
xnor U5052 (N_5052,N_4769,N_4705);
xor U5053 (N_5053,N_4487,N_4690);
or U5054 (N_5054,N_4666,N_4627);
xor U5055 (N_5055,N_4486,N_4440);
nand U5056 (N_5056,N_4417,N_4600);
nor U5057 (N_5057,N_4715,N_4425);
and U5058 (N_5058,N_4544,N_4530);
or U5059 (N_5059,N_4781,N_4516);
and U5060 (N_5060,N_4430,N_4491);
xnor U5061 (N_5061,N_4408,N_4785);
xor U5062 (N_5062,N_4781,N_4608);
nand U5063 (N_5063,N_4538,N_4746);
nand U5064 (N_5064,N_4611,N_4433);
nor U5065 (N_5065,N_4770,N_4473);
nor U5066 (N_5066,N_4535,N_4467);
nor U5067 (N_5067,N_4775,N_4454);
nand U5068 (N_5068,N_4612,N_4412);
nand U5069 (N_5069,N_4738,N_4583);
nor U5070 (N_5070,N_4449,N_4746);
or U5071 (N_5071,N_4618,N_4481);
xor U5072 (N_5072,N_4632,N_4655);
and U5073 (N_5073,N_4629,N_4529);
and U5074 (N_5074,N_4446,N_4515);
or U5075 (N_5075,N_4666,N_4722);
and U5076 (N_5076,N_4578,N_4774);
or U5077 (N_5077,N_4544,N_4649);
xnor U5078 (N_5078,N_4621,N_4602);
xor U5079 (N_5079,N_4668,N_4715);
nor U5080 (N_5080,N_4526,N_4790);
or U5081 (N_5081,N_4721,N_4481);
and U5082 (N_5082,N_4593,N_4652);
nor U5083 (N_5083,N_4548,N_4509);
or U5084 (N_5084,N_4488,N_4791);
nand U5085 (N_5085,N_4541,N_4486);
or U5086 (N_5086,N_4411,N_4444);
nand U5087 (N_5087,N_4545,N_4572);
and U5088 (N_5088,N_4790,N_4679);
xor U5089 (N_5089,N_4743,N_4767);
nand U5090 (N_5090,N_4780,N_4483);
xor U5091 (N_5091,N_4466,N_4467);
xor U5092 (N_5092,N_4752,N_4555);
xnor U5093 (N_5093,N_4714,N_4529);
nor U5094 (N_5094,N_4632,N_4758);
or U5095 (N_5095,N_4577,N_4473);
nor U5096 (N_5096,N_4445,N_4719);
xnor U5097 (N_5097,N_4608,N_4744);
nor U5098 (N_5098,N_4636,N_4569);
and U5099 (N_5099,N_4697,N_4692);
and U5100 (N_5100,N_4433,N_4799);
or U5101 (N_5101,N_4636,N_4625);
xor U5102 (N_5102,N_4562,N_4429);
nand U5103 (N_5103,N_4783,N_4572);
nand U5104 (N_5104,N_4731,N_4409);
nand U5105 (N_5105,N_4673,N_4516);
nand U5106 (N_5106,N_4794,N_4579);
nor U5107 (N_5107,N_4443,N_4722);
xor U5108 (N_5108,N_4423,N_4563);
and U5109 (N_5109,N_4736,N_4585);
and U5110 (N_5110,N_4780,N_4672);
nand U5111 (N_5111,N_4503,N_4518);
or U5112 (N_5112,N_4761,N_4462);
nor U5113 (N_5113,N_4439,N_4716);
or U5114 (N_5114,N_4594,N_4561);
nor U5115 (N_5115,N_4738,N_4506);
or U5116 (N_5116,N_4463,N_4470);
nor U5117 (N_5117,N_4477,N_4431);
or U5118 (N_5118,N_4649,N_4409);
nor U5119 (N_5119,N_4612,N_4562);
nor U5120 (N_5120,N_4732,N_4603);
nand U5121 (N_5121,N_4407,N_4571);
nor U5122 (N_5122,N_4567,N_4401);
or U5123 (N_5123,N_4798,N_4496);
nand U5124 (N_5124,N_4412,N_4532);
nand U5125 (N_5125,N_4571,N_4445);
nor U5126 (N_5126,N_4459,N_4681);
xor U5127 (N_5127,N_4733,N_4636);
xor U5128 (N_5128,N_4403,N_4674);
nor U5129 (N_5129,N_4714,N_4475);
and U5130 (N_5130,N_4606,N_4487);
and U5131 (N_5131,N_4536,N_4745);
xnor U5132 (N_5132,N_4645,N_4465);
nor U5133 (N_5133,N_4672,N_4733);
xor U5134 (N_5134,N_4707,N_4730);
and U5135 (N_5135,N_4536,N_4659);
or U5136 (N_5136,N_4765,N_4743);
nor U5137 (N_5137,N_4759,N_4755);
and U5138 (N_5138,N_4416,N_4722);
and U5139 (N_5139,N_4733,N_4593);
or U5140 (N_5140,N_4637,N_4507);
or U5141 (N_5141,N_4750,N_4577);
xor U5142 (N_5142,N_4482,N_4635);
xor U5143 (N_5143,N_4721,N_4798);
nor U5144 (N_5144,N_4625,N_4669);
nor U5145 (N_5145,N_4790,N_4762);
nor U5146 (N_5146,N_4401,N_4728);
or U5147 (N_5147,N_4642,N_4592);
and U5148 (N_5148,N_4441,N_4560);
or U5149 (N_5149,N_4675,N_4760);
nor U5150 (N_5150,N_4764,N_4729);
and U5151 (N_5151,N_4589,N_4771);
nand U5152 (N_5152,N_4577,N_4401);
nand U5153 (N_5153,N_4462,N_4592);
or U5154 (N_5154,N_4486,N_4427);
and U5155 (N_5155,N_4659,N_4535);
nor U5156 (N_5156,N_4589,N_4499);
and U5157 (N_5157,N_4768,N_4446);
nor U5158 (N_5158,N_4501,N_4562);
xor U5159 (N_5159,N_4723,N_4612);
and U5160 (N_5160,N_4752,N_4660);
nor U5161 (N_5161,N_4748,N_4609);
or U5162 (N_5162,N_4544,N_4480);
or U5163 (N_5163,N_4772,N_4721);
xnor U5164 (N_5164,N_4440,N_4650);
xor U5165 (N_5165,N_4778,N_4435);
or U5166 (N_5166,N_4402,N_4610);
and U5167 (N_5167,N_4761,N_4637);
xnor U5168 (N_5168,N_4780,N_4636);
nand U5169 (N_5169,N_4605,N_4533);
and U5170 (N_5170,N_4515,N_4505);
and U5171 (N_5171,N_4673,N_4423);
nor U5172 (N_5172,N_4558,N_4465);
nor U5173 (N_5173,N_4573,N_4661);
xnor U5174 (N_5174,N_4498,N_4542);
and U5175 (N_5175,N_4657,N_4671);
or U5176 (N_5176,N_4487,N_4581);
nor U5177 (N_5177,N_4423,N_4465);
nand U5178 (N_5178,N_4409,N_4621);
and U5179 (N_5179,N_4531,N_4748);
and U5180 (N_5180,N_4537,N_4623);
xor U5181 (N_5181,N_4607,N_4527);
nand U5182 (N_5182,N_4440,N_4612);
nor U5183 (N_5183,N_4580,N_4734);
nor U5184 (N_5184,N_4512,N_4694);
or U5185 (N_5185,N_4641,N_4569);
nor U5186 (N_5186,N_4656,N_4756);
or U5187 (N_5187,N_4624,N_4488);
xor U5188 (N_5188,N_4637,N_4572);
or U5189 (N_5189,N_4653,N_4753);
or U5190 (N_5190,N_4488,N_4744);
nor U5191 (N_5191,N_4745,N_4750);
nor U5192 (N_5192,N_4464,N_4529);
xnor U5193 (N_5193,N_4408,N_4577);
xnor U5194 (N_5194,N_4627,N_4629);
xnor U5195 (N_5195,N_4694,N_4622);
or U5196 (N_5196,N_4716,N_4667);
and U5197 (N_5197,N_4440,N_4490);
or U5198 (N_5198,N_4640,N_4468);
or U5199 (N_5199,N_4503,N_4657);
nor U5200 (N_5200,N_5139,N_4836);
nor U5201 (N_5201,N_5066,N_4884);
and U5202 (N_5202,N_5053,N_5142);
or U5203 (N_5203,N_5013,N_5118);
and U5204 (N_5204,N_5151,N_5011);
nor U5205 (N_5205,N_5137,N_4807);
or U5206 (N_5206,N_5140,N_4860);
nor U5207 (N_5207,N_5149,N_5076);
and U5208 (N_5208,N_5104,N_5070);
and U5209 (N_5209,N_5027,N_5133);
and U5210 (N_5210,N_5065,N_5183);
and U5211 (N_5211,N_5176,N_5044);
xor U5212 (N_5212,N_4985,N_4951);
xnor U5213 (N_5213,N_4847,N_5007);
xor U5214 (N_5214,N_5127,N_5086);
and U5215 (N_5215,N_4825,N_5000);
and U5216 (N_5216,N_4880,N_5004);
and U5217 (N_5217,N_5106,N_5023);
xor U5218 (N_5218,N_4958,N_4869);
or U5219 (N_5219,N_5016,N_4994);
xor U5220 (N_5220,N_5078,N_5052);
nand U5221 (N_5221,N_5006,N_4816);
nand U5222 (N_5222,N_4896,N_5074);
nand U5223 (N_5223,N_4840,N_4826);
nor U5224 (N_5224,N_5087,N_5085);
xor U5225 (N_5225,N_4913,N_5150);
nand U5226 (N_5226,N_5180,N_4843);
or U5227 (N_5227,N_4852,N_5042);
and U5228 (N_5228,N_5173,N_4982);
xnor U5229 (N_5229,N_5010,N_5162);
or U5230 (N_5230,N_5121,N_5136);
and U5231 (N_5231,N_4943,N_5100);
or U5232 (N_5232,N_4992,N_4952);
nand U5233 (N_5233,N_4933,N_4820);
nand U5234 (N_5234,N_4903,N_4802);
xnor U5235 (N_5235,N_5026,N_4881);
nand U5236 (N_5236,N_5029,N_4909);
and U5237 (N_5237,N_4928,N_5040);
or U5238 (N_5238,N_5194,N_4882);
nor U5239 (N_5239,N_4932,N_5135);
and U5240 (N_5240,N_4887,N_4835);
nor U5241 (N_5241,N_5167,N_4937);
and U5242 (N_5242,N_5037,N_4894);
nor U5243 (N_5243,N_4839,N_4904);
nor U5244 (N_5244,N_5071,N_4817);
and U5245 (N_5245,N_5148,N_4912);
or U5246 (N_5246,N_4968,N_4824);
nand U5247 (N_5247,N_4963,N_4919);
xor U5248 (N_5248,N_5022,N_5036);
nor U5249 (N_5249,N_5107,N_5034);
nor U5250 (N_5250,N_5064,N_5182);
and U5251 (N_5251,N_4845,N_5120);
nor U5252 (N_5252,N_4874,N_5166);
nand U5253 (N_5253,N_4871,N_5055);
xor U5254 (N_5254,N_5080,N_4953);
and U5255 (N_5255,N_5072,N_4828);
xor U5256 (N_5256,N_4853,N_5132);
xor U5257 (N_5257,N_4973,N_4892);
nor U5258 (N_5258,N_4942,N_4831);
nand U5259 (N_5259,N_5181,N_5169);
nor U5260 (N_5260,N_4927,N_4955);
nor U5261 (N_5261,N_5138,N_5122);
and U5262 (N_5262,N_4800,N_5110);
nand U5263 (N_5263,N_5081,N_4893);
and U5264 (N_5264,N_5045,N_4837);
or U5265 (N_5265,N_5189,N_5105);
and U5266 (N_5266,N_5184,N_5159);
and U5267 (N_5267,N_5021,N_5093);
xnor U5268 (N_5268,N_5198,N_5126);
or U5269 (N_5269,N_4987,N_5039);
xnor U5270 (N_5270,N_4944,N_4876);
nor U5271 (N_5271,N_5089,N_5079);
nor U5272 (N_5272,N_4939,N_5156);
or U5273 (N_5273,N_4935,N_4834);
xnor U5274 (N_5274,N_4849,N_5134);
xor U5275 (N_5275,N_5129,N_5157);
and U5276 (N_5276,N_5009,N_4812);
nand U5277 (N_5277,N_5090,N_5113);
nor U5278 (N_5278,N_4936,N_5188);
xor U5279 (N_5279,N_4901,N_5178);
nor U5280 (N_5280,N_4907,N_4844);
nor U5281 (N_5281,N_5197,N_4999);
and U5282 (N_5282,N_4854,N_4997);
nor U5283 (N_5283,N_5145,N_5082);
or U5284 (N_5284,N_5108,N_5175);
and U5285 (N_5285,N_5114,N_4917);
or U5286 (N_5286,N_4865,N_5047);
nor U5287 (N_5287,N_5186,N_5119);
or U5288 (N_5288,N_4855,N_4924);
or U5289 (N_5289,N_5060,N_5094);
nor U5290 (N_5290,N_4803,N_5024);
nand U5291 (N_5291,N_4851,N_5102);
nor U5292 (N_5292,N_4804,N_5141);
nand U5293 (N_5293,N_5192,N_5097);
nor U5294 (N_5294,N_5005,N_4883);
nand U5295 (N_5295,N_5112,N_5062);
nor U5296 (N_5296,N_5179,N_4988);
nor U5297 (N_5297,N_5038,N_5115);
nor U5298 (N_5298,N_5098,N_5050);
xnor U5299 (N_5299,N_4918,N_4940);
and U5300 (N_5300,N_4986,N_4885);
and U5301 (N_5301,N_5043,N_5172);
xor U5302 (N_5302,N_5031,N_4900);
nor U5303 (N_5303,N_4850,N_4926);
and U5304 (N_5304,N_5032,N_5155);
nand U5305 (N_5305,N_4878,N_5018);
nand U5306 (N_5306,N_5035,N_4947);
nand U5307 (N_5307,N_5091,N_4960);
or U5308 (N_5308,N_5161,N_5187);
or U5309 (N_5309,N_4975,N_5083);
xor U5310 (N_5310,N_4981,N_5163);
or U5311 (N_5311,N_4815,N_4827);
nand U5312 (N_5312,N_5067,N_4931);
nand U5313 (N_5313,N_5049,N_5130);
nor U5314 (N_5314,N_4964,N_4808);
xnor U5315 (N_5315,N_5077,N_4971);
nand U5316 (N_5316,N_4846,N_5111);
xnor U5317 (N_5317,N_5190,N_5058);
nand U5318 (N_5318,N_5088,N_4891);
nand U5319 (N_5319,N_5003,N_4866);
and U5320 (N_5320,N_4915,N_4864);
and U5321 (N_5321,N_5025,N_4923);
nor U5322 (N_5322,N_5041,N_5124);
or U5323 (N_5323,N_5061,N_5063);
or U5324 (N_5324,N_4862,N_5015);
or U5325 (N_5325,N_4910,N_5160);
xnor U5326 (N_5326,N_4821,N_5191);
and U5327 (N_5327,N_4967,N_4993);
nand U5328 (N_5328,N_4950,N_5158);
xnor U5329 (N_5329,N_4822,N_5057);
and U5330 (N_5330,N_4990,N_5103);
nor U5331 (N_5331,N_5084,N_4859);
and U5332 (N_5332,N_5146,N_4886);
or U5333 (N_5333,N_4823,N_5147);
nor U5334 (N_5334,N_5168,N_4945);
nand U5335 (N_5335,N_5030,N_4969);
nor U5336 (N_5336,N_5193,N_4956);
or U5337 (N_5337,N_4995,N_4830);
xor U5338 (N_5338,N_4929,N_5170);
and U5339 (N_5339,N_5095,N_4998);
xnor U5340 (N_5340,N_4813,N_5019);
or U5341 (N_5341,N_5154,N_4983);
nand U5342 (N_5342,N_4934,N_4962);
or U5343 (N_5343,N_4879,N_5012);
nor U5344 (N_5344,N_4925,N_4938);
nor U5345 (N_5345,N_5069,N_4957);
and U5346 (N_5346,N_4861,N_5131);
or U5347 (N_5347,N_5020,N_4970);
nor U5348 (N_5348,N_5068,N_5073);
and U5349 (N_5349,N_5092,N_4867);
and U5350 (N_5350,N_5056,N_5101);
nor U5351 (N_5351,N_4870,N_5117);
or U5352 (N_5352,N_4911,N_4902);
nand U5353 (N_5353,N_4805,N_4978);
nor U5354 (N_5354,N_4801,N_4991);
xor U5355 (N_5355,N_5075,N_5109);
nor U5356 (N_5356,N_4966,N_5196);
or U5357 (N_5357,N_4819,N_4806);
or U5358 (N_5358,N_5002,N_4890);
or U5359 (N_5359,N_4895,N_4946);
nor U5360 (N_5360,N_5143,N_4948);
and U5361 (N_5361,N_5096,N_4974);
nor U5362 (N_5362,N_4972,N_4941);
nand U5363 (N_5363,N_5017,N_4857);
nor U5364 (N_5364,N_5123,N_5128);
and U5365 (N_5365,N_4889,N_5152);
or U5366 (N_5366,N_4842,N_5028);
xor U5367 (N_5367,N_5054,N_5144);
nand U5368 (N_5368,N_4829,N_5014);
xnor U5369 (N_5369,N_5001,N_4921);
or U5370 (N_5370,N_5165,N_4809);
nor U5371 (N_5371,N_5171,N_4856);
and U5372 (N_5372,N_4872,N_5195);
nand U5373 (N_5373,N_4818,N_4961);
or U5374 (N_5374,N_4984,N_5048);
nand U5375 (N_5375,N_4848,N_4989);
nand U5376 (N_5376,N_5125,N_4908);
nor U5377 (N_5377,N_4877,N_5174);
nand U5378 (N_5378,N_5199,N_5059);
nand U5379 (N_5379,N_5033,N_4949);
xnor U5380 (N_5380,N_4838,N_5185);
or U5381 (N_5381,N_5046,N_5164);
nor U5382 (N_5382,N_4841,N_4954);
or U5383 (N_5383,N_4814,N_4977);
nor U5384 (N_5384,N_4965,N_4996);
nor U5385 (N_5385,N_4976,N_4930);
and U5386 (N_5386,N_4868,N_5008);
and U5387 (N_5387,N_5051,N_4833);
and U5388 (N_5388,N_4916,N_4811);
nand U5389 (N_5389,N_4875,N_4888);
xnor U5390 (N_5390,N_4810,N_4906);
nand U5391 (N_5391,N_5153,N_4980);
and U5392 (N_5392,N_4863,N_4832);
or U5393 (N_5393,N_4959,N_5177);
or U5394 (N_5394,N_4979,N_5099);
and U5395 (N_5395,N_4899,N_4905);
and U5396 (N_5396,N_4920,N_4873);
xor U5397 (N_5397,N_4858,N_4898);
nor U5398 (N_5398,N_4914,N_4922);
nand U5399 (N_5399,N_5116,N_4897);
or U5400 (N_5400,N_5029,N_5002);
nor U5401 (N_5401,N_4896,N_4917);
xor U5402 (N_5402,N_4890,N_5172);
xnor U5403 (N_5403,N_4936,N_4953);
or U5404 (N_5404,N_5060,N_5071);
nor U5405 (N_5405,N_4827,N_5083);
nand U5406 (N_5406,N_4965,N_5013);
or U5407 (N_5407,N_4991,N_4990);
xnor U5408 (N_5408,N_5030,N_4895);
nor U5409 (N_5409,N_5182,N_4914);
xnor U5410 (N_5410,N_5109,N_4920);
nor U5411 (N_5411,N_4981,N_5012);
xor U5412 (N_5412,N_5008,N_4855);
and U5413 (N_5413,N_5084,N_4817);
nor U5414 (N_5414,N_4886,N_5103);
nand U5415 (N_5415,N_5179,N_5144);
nand U5416 (N_5416,N_4824,N_4840);
and U5417 (N_5417,N_4892,N_5186);
xnor U5418 (N_5418,N_4825,N_4901);
xnor U5419 (N_5419,N_4851,N_5136);
and U5420 (N_5420,N_4993,N_5180);
xnor U5421 (N_5421,N_4905,N_5163);
xnor U5422 (N_5422,N_4896,N_4809);
nor U5423 (N_5423,N_5162,N_5054);
or U5424 (N_5424,N_4802,N_4927);
or U5425 (N_5425,N_5069,N_5043);
xnor U5426 (N_5426,N_4932,N_4849);
or U5427 (N_5427,N_4802,N_5146);
nand U5428 (N_5428,N_4882,N_5146);
or U5429 (N_5429,N_4809,N_4812);
or U5430 (N_5430,N_5170,N_4849);
nor U5431 (N_5431,N_4931,N_4861);
nand U5432 (N_5432,N_5113,N_4880);
and U5433 (N_5433,N_4946,N_4934);
and U5434 (N_5434,N_5172,N_5031);
nand U5435 (N_5435,N_4811,N_4880);
nor U5436 (N_5436,N_5032,N_5097);
and U5437 (N_5437,N_5150,N_4864);
nand U5438 (N_5438,N_5032,N_4846);
xnor U5439 (N_5439,N_4866,N_5172);
or U5440 (N_5440,N_4940,N_4812);
xor U5441 (N_5441,N_5063,N_5160);
nand U5442 (N_5442,N_4839,N_5142);
xor U5443 (N_5443,N_5148,N_4988);
or U5444 (N_5444,N_4837,N_4864);
xnor U5445 (N_5445,N_5113,N_4898);
and U5446 (N_5446,N_5001,N_5081);
xor U5447 (N_5447,N_5008,N_4940);
xor U5448 (N_5448,N_4802,N_4915);
nor U5449 (N_5449,N_5137,N_5190);
and U5450 (N_5450,N_4855,N_5187);
or U5451 (N_5451,N_5194,N_4801);
xnor U5452 (N_5452,N_4803,N_5038);
nor U5453 (N_5453,N_4896,N_5056);
and U5454 (N_5454,N_5121,N_5021);
xor U5455 (N_5455,N_4813,N_4959);
xor U5456 (N_5456,N_4816,N_5157);
nand U5457 (N_5457,N_5043,N_5135);
nor U5458 (N_5458,N_5194,N_4902);
xor U5459 (N_5459,N_5114,N_4806);
nand U5460 (N_5460,N_4803,N_5083);
nand U5461 (N_5461,N_5024,N_4839);
nand U5462 (N_5462,N_4933,N_5018);
nand U5463 (N_5463,N_5192,N_4850);
xor U5464 (N_5464,N_5134,N_4991);
or U5465 (N_5465,N_5045,N_5077);
nor U5466 (N_5466,N_4960,N_4945);
xnor U5467 (N_5467,N_4821,N_4985);
xnor U5468 (N_5468,N_5139,N_4977);
or U5469 (N_5469,N_4856,N_4816);
nand U5470 (N_5470,N_4809,N_4874);
and U5471 (N_5471,N_4879,N_5108);
and U5472 (N_5472,N_4848,N_4804);
nand U5473 (N_5473,N_4907,N_5171);
and U5474 (N_5474,N_4879,N_4947);
nand U5475 (N_5475,N_4843,N_5172);
nand U5476 (N_5476,N_4976,N_5139);
or U5477 (N_5477,N_5068,N_5156);
nor U5478 (N_5478,N_4949,N_5143);
xnor U5479 (N_5479,N_5042,N_4946);
nor U5480 (N_5480,N_5046,N_4945);
xor U5481 (N_5481,N_4965,N_4858);
or U5482 (N_5482,N_4904,N_4974);
or U5483 (N_5483,N_4830,N_4965);
xor U5484 (N_5484,N_5020,N_4892);
or U5485 (N_5485,N_4994,N_5152);
or U5486 (N_5486,N_4988,N_5163);
or U5487 (N_5487,N_5103,N_5040);
nor U5488 (N_5488,N_4905,N_5064);
xnor U5489 (N_5489,N_4931,N_5120);
and U5490 (N_5490,N_5025,N_5106);
xnor U5491 (N_5491,N_4958,N_5108);
nor U5492 (N_5492,N_5129,N_5192);
and U5493 (N_5493,N_5081,N_5054);
nor U5494 (N_5494,N_5007,N_4905);
and U5495 (N_5495,N_5047,N_5084);
nor U5496 (N_5496,N_5156,N_4839);
or U5497 (N_5497,N_4889,N_4936);
xnor U5498 (N_5498,N_5063,N_5001);
and U5499 (N_5499,N_4980,N_4802);
and U5500 (N_5500,N_4912,N_4926);
and U5501 (N_5501,N_5190,N_4898);
or U5502 (N_5502,N_4853,N_5064);
and U5503 (N_5503,N_4955,N_4905);
nand U5504 (N_5504,N_5163,N_5129);
xor U5505 (N_5505,N_4830,N_5150);
nand U5506 (N_5506,N_4882,N_4920);
xor U5507 (N_5507,N_5122,N_4916);
xnor U5508 (N_5508,N_5042,N_4889);
or U5509 (N_5509,N_4954,N_4863);
nand U5510 (N_5510,N_4987,N_4867);
nor U5511 (N_5511,N_4911,N_5043);
or U5512 (N_5512,N_5183,N_4965);
nand U5513 (N_5513,N_5089,N_5183);
xor U5514 (N_5514,N_4826,N_4835);
and U5515 (N_5515,N_5080,N_4866);
and U5516 (N_5516,N_5045,N_4892);
and U5517 (N_5517,N_5088,N_5074);
or U5518 (N_5518,N_4989,N_5060);
and U5519 (N_5519,N_5163,N_5108);
nor U5520 (N_5520,N_4867,N_4933);
or U5521 (N_5521,N_5160,N_4868);
nand U5522 (N_5522,N_4886,N_5129);
nand U5523 (N_5523,N_5182,N_4998);
and U5524 (N_5524,N_4873,N_5138);
or U5525 (N_5525,N_4931,N_5194);
nand U5526 (N_5526,N_5189,N_5112);
xnor U5527 (N_5527,N_4840,N_5088);
nand U5528 (N_5528,N_5033,N_5137);
and U5529 (N_5529,N_5124,N_4860);
or U5530 (N_5530,N_5024,N_5058);
xor U5531 (N_5531,N_4969,N_5173);
nand U5532 (N_5532,N_5032,N_5070);
nand U5533 (N_5533,N_5146,N_5085);
and U5534 (N_5534,N_5108,N_4867);
and U5535 (N_5535,N_5111,N_4836);
or U5536 (N_5536,N_5183,N_5134);
and U5537 (N_5537,N_5141,N_4887);
nor U5538 (N_5538,N_4819,N_5110);
nor U5539 (N_5539,N_4861,N_4970);
xnor U5540 (N_5540,N_5091,N_4822);
nand U5541 (N_5541,N_5109,N_4852);
nor U5542 (N_5542,N_4970,N_4984);
or U5543 (N_5543,N_4866,N_4975);
or U5544 (N_5544,N_5025,N_4833);
xnor U5545 (N_5545,N_5111,N_4894);
and U5546 (N_5546,N_5002,N_5177);
or U5547 (N_5547,N_5121,N_5071);
xor U5548 (N_5548,N_5140,N_5143);
xnor U5549 (N_5549,N_4807,N_5117);
and U5550 (N_5550,N_5020,N_5072);
nor U5551 (N_5551,N_5007,N_4943);
nand U5552 (N_5552,N_5100,N_4955);
xor U5553 (N_5553,N_5180,N_4918);
or U5554 (N_5554,N_5035,N_4982);
and U5555 (N_5555,N_5188,N_4970);
and U5556 (N_5556,N_5049,N_4815);
nand U5557 (N_5557,N_4928,N_4940);
and U5558 (N_5558,N_4950,N_5122);
nor U5559 (N_5559,N_4803,N_4912);
nand U5560 (N_5560,N_4834,N_5057);
nor U5561 (N_5561,N_4965,N_4980);
xor U5562 (N_5562,N_4996,N_4981);
or U5563 (N_5563,N_4993,N_5178);
nor U5564 (N_5564,N_5172,N_5120);
nand U5565 (N_5565,N_5100,N_5049);
nand U5566 (N_5566,N_4995,N_4832);
nor U5567 (N_5567,N_4828,N_4969);
nand U5568 (N_5568,N_5131,N_5035);
nand U5569 (N_5569,N_4895,N_4944);
nand U5570 (N_5570,N_5117,N_4844);
nor U5571 (N_5571,N_4815,N_4877);
and U5572 (N_5572,N_5125,N_4854);
nand U5573 (N_5573,N_5090,N_5130);
nor U5574 (N_5574,N_5085,N_5072);
and U5575 (N_5575,N_5180,N_5114);
xor U5576 (N_5576,N_4893,N_4811);
nor U5577 (N_5577,N_5123,N_5149);
xor U5578 (N_5578,N_5082,N_4803);
nand U5579 (N_5579,N_5162,N_5041);
and U5580 (N_5580,N_5118,N_4874);
and U5581 (N_5581,N_5145,N_5118);
nand U5582 (N_5582,N_4807,N_5056);
or U5583 (N_5583,N_4810,N_4840);
nand U5584 (N_5584,N_5003,N_4904);
xor U5585 (N_5585,N_4844,N_4996);
nor U5586 (N_5586,N_5152,N_4838);
xor U5587 (N_5587,N_4836,N_4928);
or U5588 (N_5588,N_4985,N_4823);
nand U5589 (N_5589,N_4860,N_4982);
or U5590 (N_5590,N_5009,N_5144);
and U5591 (N_5591,N_5080,N_5065);
or U5592 (N_5592,N_5155,N_4930);
nor U5593 (N_5593,N_4955,N_4972);
or U5594 (N_5594,N_4980,N_5166);
and U5595 (N_5595,N_5103,N_4805);
nand U5596 (N_5596,N_4991,N_5078);
nand U5597 (N_5597,N_4946,N_4953);
xor U5598 (N_5598,N_5007,N_4974);
xnor U5599 (N_5599,N_4829,N_5165);
and U5600 (N_5600,N_5513,N_5377);
or U5601 (N_5601,N_5353,N_5560);
nor U5602 (N_5602,N_5554,N_5271);
and U5603 (N_5603,N_5458,N_5260);
nand U5604 (N_5604,N_5504,N_5251);
or U5605 (N_5605,N_5323,N_5327);
xnor U5606 (N_5606,N_5390,N_5308);
nor U5607 (N_5607,N_5403,N_5439);
or U5608 (N_5608,N_5419,N_5510);
or U5609 (N_5609,N_5575,N_5384);
nor U5610 (N_5610,N_5380,N_5209);
nand U5611 (N_5611,N_5480,N_5434);
nand U5612 (N_5612,N_5290,N_5548);
xnor U5613 (N_5613,N_5282,N_5461);
nor U5614 (N_5614,N_5336,N_5596);
nand U5615 (N_5615,N_5404,N_5246);
nor U5616 (N_5616,N_5459,N_5597);
or U5617 (N_5617,N_5328,N_5430);
xnor U5618 (N_5618,N_5339,N_5495);
xnor U5619 (N_5619,N_5231,N_5499);
nand U5620 (N_5620,N_5526,N_5455);
or U5621 (N_5621,N_5305,N_5381);
nand U5622 (N_5622,N_5279,N_5393);
nand U5623 (N_5623,N_5345,N_5334);
or U5624 (N_5624,N_5230,N_5235);
nor U5625 (N_5625,N_5478,N_5340);
nor U5626 (N_5626,N_5262,N_5457);
nor U5627 (N_5627,N_5324,N_5483);
nor U5628 (N_5628,N_5268,N_5302);
nor U5629 (N_5629,N_5274,N_5201);
xor U5630 (N_5630,N_5446,N_5234);
nor U5631 (N_5631,N_5533,N_5202);
and U5632 (N_5632,N_5584,N_5438);
nand U5633 (N_5633,N_5476,N_5232);
nand U5634 (N_5634,N_5292,N_5316);
nand U5635 (N_5635,N_5304,N_5225);
and U5636 (N_5636,N_5501,N_5203);
nand U5637 (N_5637,N_5432,N_5307);
nor U5638 (N_5638,N_5433,N_5443);
xnor U5639 (N_5639,N_5357,N_5341);
and U5640 (N_5640,N_5352,N_5488);
and U5641 (N_5641,N_5534,N_5364);
xnor U5642 (N_5642,N_5583,N_5541);
or U5643 (N_5643,N_5485,N_5423);
or U5644 (N_5644,N_5374,N_5589);
nand U5645 (N_5645,N_5417,N_5227);
nand U5646 (N_5646,N_5278,N_5372);
and U5647 (N_5647,N_5286,N_5591);
xor U5648 (N_5648,N_5537,N_5369);
xor U5649 (N_5649,N_5284,N_5317);
nand U5650 (N_5650,N_5294,N_5378);
or U5651 (N_5651,N_5258,N_5545);
xnor U5652 (N_5652,N_5303,N_5330);
xor U5653 (N_5653,N_5517,N_5261);
nand U5654 (N_5654,N_5557,N_5590);
or U5655 (N_5655,N_5358,N_5559);
xnor U5656 (N_5656,N_5578,N_5579);
and U5657 (N_5657,N_5204,N_5542);
and U5658 (N_5658,N_5319,N_5418);
xor U5659 (N_5659,N_5569,N_5530);
nor U5660 (N_5660,N_5572,N_5405);
nand U5661 (N_5661,N_5524,N_5255);
and U5662 (N_5662,N_5528,N_5257);
nor U5663 (N_5663,N_5344,N_5347);
nor U5664 (N_5664,N_5426,N_5506);
nor U5665 (N_5665,N_5291,N_5587);
or U5666 (N_5666,N_5211,N_5236);
or U5667 (N_5667,N_5566,N_5332);
xnor U5668 (N_5668,N_5217,N_5472);
xnor U5669 (N_5669,N_5402,N_5277);
nand U5670 (N_5670,N_5266,N_5376);
nand U5671 (N_5671,N_5555,N_5571);
and U5672 (N_5672,N_5422,N_5233);
nand U5673 (N_5673,N_5318,N_5539);
nand U5674 (N_5674,N_5300,N_5360);
and U5675 (N_5675,N_5511,N_5259);
nand U5676 (N_5676,N_5296,N_5482);
nand U5677 (N_5677,N_5490,N_5410);
nand U5678 (N_5678,N_5283,N_5370);
nor U5679 (N_5679,N_5514,N_5315);
nor U5680 (N_5680,N_5264,N_5212);
xor U5681 (N_5681,N_5200,N_5391);
xor U5682 (N_5682,N_5523,N_5582);
xor U5683 (N_5683,N_5289,N_5263);
nor U5684 (N_5684,N_5320,N_5500);
xor U5685 (N_5685,N_5245,N_5564);
and U5686 (N_5686,N_5389,N_5301);
and U5687 (N_5687,N_5477,N_5536);
or U5688 (N_5688,N_5313,N_5428);
nand U5689 (N_5689,N_5348,N_5516);
or U5690 (N_5690,N_5474,N_5210);
and U5691 (N_5691,N_5363,N_5208);
and U5692 (N_5692,N_5576,N_5242);
or U5693 (N_5693,N_5414,N_5401);
xor U5694 (N_5694,N_5355,N_5333);
or U5695 (N_5695,N_5558,N_5385);
and U5696 (N_5696,N_5416,N_5522);
and U5697 (N_5697,N_5529,N_5441);
xnor U5698 (N_5698,N_5415,N_5365);
and U5699 (N_5699,N_5281,N_5598);
nand U5700 (N_5700,N_5429,N_5409);
nor U5701 (N_5701,N_5437,N_5556);
xnor U5702 (N_5702,N_5270,N_5399);
nand U5703 (N_5703,N_5435,N_5407);
nor U5704 (N_5704,N_5465,N_5521);
nor U5705 (N_5705,N_5525,N_5487);
and U5706 (N_5706,N_5505,N_5585);
or U5707 (N_5707,N_5515,N_5354);
and U5708 (N_5708,N_5386,N_5400);
and U5709 (N_5709,N_5338,N_5295);
nor U5710 (N_5710,N_5244,N_5298);
nand U5711 (N_5711,N_5420,N_5456);
nand U5712 (N_5712,N_5498,N_5322);
and U5713 (N_5713,N_5509,N_5469);
nand U5714 (N_5714,N_5253,N_5594);
xor U5715 (N_5715,N_5563,N_5512);
xnor U5716 (N_5716,N_5468,N_5481);
nand U5717 (N_5717,N_5342,N_5424);
or U5718 (N_5718,N_5220,N_5215);
nor U5719 (N_5719,N_5224,N_5392);
and U5720 (N_5720,N_5273,N_5275);
nor U5721 (N_5721,N_5249,N_5346);
or U5722 (N_5722,N_5361,N_5207);
nand U5723 (N_5723,N_5586,N_5466);
or U5724 (N_5724,N_5219,N_5397);
nand U5725 (N_5725,N_5454,N_5460);
or U5726 (N_5726,N_5494,N_5535);
and U5727 (N_5727,N_5497,N_5412);
and U5728 (N_5728,N_5350,N_5240);
and U5729 (N_5729,N_5321,N_5272);
or U5730 (N_5730,N_5565,N_5206);
or U5731 (N_5731,N_5444,N_5508);
nand U5732 (N_5732,N_5570,N_5577);
or U5733 (N_5733,N_5551,N_5593);
xor U5734 (N_5734,N_5507,N_5337);
nand U5735 (N_5735,N_5213,N_5451);
xor U5736 (N_5736,N_5568,N_5371);
xnor U5737 (N_5737,N_5325,N_5285);
xnor U5738 (N_5738,N_5309,N_5448);
nand U5739 (N_5739,N_5373,N_5493);
and U5740 (N_5740,N_5408,N_5229);
or U5741 (N_5741,N_5398,N_5519);
nor U5742 (N_5742,N_5248,N_5595);
or U5743 (N_5743,N_5351,N_5237);
or U5744 (N_5744,N_5543,N_5411);
or U5745 (N_5745,N_5561,N_5449);
and U5746 (N_5746,N_5471,N_5254);
and U5747 (N_5747,N_5581,N_5310);
xnor U5748 (N_5748,N_5427,N_5395);
and U5749 (N_5749,N_5492,N_5574);
xor U5750 (N_5750,N_5226,N_5531);
nor U5751 (N_5751,N_5463,N_5479);
nor U5752 (N_5752,N_5383,N_5518);
and U5753 (N_5753,N_5573,N_5238);
nand U5754 (N_5754,N_5440,N_5221);
nand U5755 (N_5755,N_5538,N_5445);
and U5756 (N_5756,N_5314,N_5484);
nor U5757 (N_5757,N_5382,N_5306);
nor U5758 (N_5758,N_5567,N_5367);
nor U5759 (N_5759,N_5413,N_5205);
and U5760 (N_5760,N_5216,N_5239);
and U5761 (N_5761,N_5243,N_5450);
xor U5762 (N_5762,N_5362,N_5228);
xnor U5763 (N_5763,N_5288,N_5540);
xor U5764 (N_5764,N_5452,N_5502);
xnor U5765 (N_5765,N_5553,N_5475);
and U5766 (N_5766,N_5467,N_5599);
and U5767 (N_5767,N_5473,N_5247);
and U5768 (N_5768,N_5326,N_5453);
or U5769 (N_5769,N_5470,N_5375);
xor U5770 (N_5770,N_5520,N_5588);
and U5771 (N_5771,N_5241,N_5256);
nor U5772 (N_5772,N_5299,N_5267);
and U5773 (N_5773,N_5287,N_5464);
or U5774 (N_5774,N_5486,N_5368);
nor U5775 (N_5775,N_5343,N_5222);
or U5776 (N_5776,N_5544,N_5552);
nor U5777 (N_5777,N_5447,N_5218);
nor U5778 (N_5778,N_5546,N_5388);
nand U5779 (N_5779,N_5462,N_5312);
nor U5780 (N_5780,N_5379,N_5293);
nor U5781 (N_5781,N_5562,N_5265);
nand U5782 (N_5782,N_5387,N_5406);
or U5783 (N_5783,N_5214,N_5550);
nor U5784 (N_5784,N_5366,N_5252);
xor U5785 (N_5785,N_5394,N_5335);
or U5786 (N_5786,N_5297,N_5356);
and U5787 (N_5787,N_5532,N_5580);
or U5788 (N_5788,N_5496,N_5549);
and U5789 (N_5789,N_5503,N_5359);
nor U5790 (N_5790,N_5442,N_5592);
nand U5791 (N_5791,N_5311,N_5436);
nor U5792 (N_5792,N_5331,N_5431);
nand U5793 (N_5793,N_5269,N_5421);
nand U5794 (N_5794,N_5223,N_5396);
nand U5795 (N_5795,N_5250,N_5491);
nor U5796 (N_5796,N_5547,N_5276);
and U5797 (N_5797,N_5280,N_5425);
nor U5798 (N_5798,N_5329,N_5489);
nor U5799 (N_5799,N_5349,N_5527);
nand U5800 (N_5800,N_5594,N_5451);
nor U5801 (N_5801,N_5355,N_5283);
nor U5802 (N_5802,N_5392,N_5315);
xnor U5803 (N_5803,N_5393,N_5500);
and U5804 (N_5804,N_5284,N_5312);
nand U5805 (N_5805,N_5336,N_5266);
or U5806 (N_5806,N_5437,N_5301);
xor U5807 (N_5807,N_5305,N_5454);
and U5808 (N_5808,N_5297,N_5428);
nand U5809 (N_5809,N_5339,N_5257);
xnor U5810 (N_5810,N_5578,N_5473);
or U5811 (N_5811,N_5291,N_5558);
or U5812 (N_5812,N_5583,N_5528);
or U5813 (N_5813,N_5265,N_5202);
xor U5814 (N_5814,N_5242,N_5328);
nand U5815 (N_5815,N_5443,N_5487);
or U5816 (N_5816,N_5266,N_5508);
or U5817 (N_5817,N_5483,N_5550);
and U5818 (N_5818,N_5575,N_5407);
and U5819 (N_5819,N_5248,N_5214);
nor U5820 (N_5820,N_5252,N_5494);
nand U5821 (N_5821,N_5588,N_5318);
xnor U5822 (N_5822,N_5223,N_5273);
xor U5823 (N_5823,N_5462,N_5244);
nand U5824 (N_5824,N_5213,N_5592);
xor U5825 (N_5825,N_5595,N_5347);
or U5826 (N_5826,N_5269,N_5243);
xor U5827 (N_5827,N_5321,N_5546);
nor U5828 (N_5828,N_5400,N_5398);
nand U5829 (N_5829,N_5599,N_5365);
nor U5830 (N_5830,N_5317,N_5497);
nor U5831 (N_5831,N_5232,N_5404);
nand U5832 (N_5832,N_5222,N_5487);
nor U5833 (N_5833,N_5562,N_5394);
or U5834 (N_5834,N_5438,N_5583);
nor U5835 (N_5835,N_5373,N_5267);
and U5836 (N_5836,N_5290,N_5585);
nand U5837 (N_5837,N_5218,N_5473);
nand U5838 (N_5838,N_5371,N_5507);
xor U5839 (N_5839,N_5253,N_5299);
or U5840 (N_5840,N_5233,N_5389);
nand U5841 (N_5841,N_5468,N_5586);
xor U5842 (N_5842,N_5487,N_5582);
or U5843 (N_5843,N_5249,N_5504);
or U5844 (N_5844,N_5497,N_5496);
and U5845 (N_5845,N_5562,N_5364);
nand U5846 (N_5846,N_5244,N_5517);
nand U5847 (N_5847,N_5465,N_5291);
nor U5848 (N_5848,N_5201,N_5325);
nand U5849 (N_5849,N_5477,N_5412);
or U5850 (N_5850,N_5587,N_5435);
xnor U5851 (N_5851,N_5458,N_5432);
nand U5852 (N_5852,N_5586,N_5203);
and U5853 (N_5853,N_5252,N_5419);
and U5854 (N_5854,N_5205,N_5262);
xor U5855 (N_5855,N_5536,N_5351);
or U5856 (N_5856,N_5239,N_5428);
and U5857 (N_5857,N_5418,N_5261);
nor U5858 (N_5858,N_5571,N_5249);
nor U5859 (N_5859,N_5426,N_5597);
nand U5860 (N_5860,N_5396,N_5343);
xnor U5861 (N_5861,N_5374,N_5514);
nor U5862 (N_5862,N_5302,N_5446);
or U5863 (N_5863,N_5466,N_5592);
or U5864 (N_5864,N_5317,N_5238);
and U5865 (N_5865,N_5527,N_5486);
xor U5866 (N_5866,N_5200,N_5402);
nor U5867 (N_5867,N_5570,N_5575);
xnor U5868 (N_5868,N_5593,N_5465);
nand U5869 (N_5869,N_5554,N_5267);
nand U5870 (N_5870,N_5239,N_5322);
or U5871 (N_5871,N_5371,N_5499);
nand U5872 (N_5872,N_5344,N_5296);
or U5873 (N_5873,N_5281,N_5432);
xor U5874 (N_5874,N_5566,N_5471);
xnor U5875 (N_5875,N_5332,N_5558);
or U5876 (N_5876,N_5452,N_5302);
nor U5877 (N_5877,N_5561,N_5417);
nor U5878 (N_5878,N_5503,N_5374);
nor U5879 (N_5879,N_5459,N_5493);
nor U5880 (N_5880,N_5557,N_5364);
xor U5881 (N_5881,N_5554,N_5218);
or U5882 (N_5882,N_5379,N_5519);
or U5883 (N_5883,N_5483,N_5372);
nor U5884 (N_5884,N_5452,N_5402);
or U5885 (N_5885,N_5280,N_5553);
nor U5886 (N_5886,N_5580,N_5423);
nand U5887 (N_5887,N_5469,N_5376);
nand U5888 (N_5888,N_5204,N_5328);
or U5889 (N_5889,N_5265,N_5405);
nand U5890 (N_5890,N_5323,N_5452);
nand U5891 (N_5891,N_5268,N_5381);
xnor U5892 (N_5892,N_5421,N_5324);
xor U5893 (N_5893,N_5274,N_5361);
and U5894 (N_5894,N_5444,N_5455);
or U5895 (N_5895,N_5228,N_5590);
nand U5896 (N_5896,N_5377,N_5356);
nor U5897 (N_5897,N_5355,N_5320);
nand U5898 (N_5898,N_5440,N_5279);
xnor U5899 (N_5899,N_5569,N_5238);
or U5900 (N_5900,N_5275,N_5587);
nand U5901 (N_5901,N_5570,N_5588);
and U5902 (N_5902,N_5532,N_5392);
nand U5903 (N_5903,N_5345,N_5487);
or U5904 (N_5904,N_5340,N_5531);
and U5905 (N_5905,N_5563,N_5264);
and U5906 (N_5906,N_5245,N_5271);
and U5907 (N_5907,N_5256,N_5226);
xor U5908 (N_5908,N_5354,N_5444);
xnor U5909 (N_5909,N_5437,N_5232);
and U5910 (N_5910,N_5250,N_5408);
nand U5911 (N_5911,N_5456,N_5205);
xor U5912 (N_5912,N_5217,N_5434);
and U5913 (N_5913,N_5498,N_5220);
xnor U5914 (N_5914,N_5507,N_5487);
or U5915 (N_5915,N_5411,N_5348);
nand U5916 (N_5916,N_5293,N_5492);
nor U5917 (N_5917,N_5329,N_5501);
and U5918 (N_5918,N_5250,N_5490);
and U5919 (N_5919,N_5393,N_5592);
nor U5920 (N_5920,N_5548,N_5297);
and U5921 (N_5921,N_5200,N_5525);
or U5922 (N_5922,N_5455,N_5492);
nand U5923 (N_5923,N_5239,N_5248);
nand U5924 (N_5924,N_5248,N_5564);
and U5925 (N_5925,N_5342,N_5545);
nor U5926 (N_5926,N_5444,N_5487);
and U5927 (N_5927,N_5372,N_5284);
nand U5928 (N_5928,N_5532,N_5408);
nand U5929 (N_5929,N_5358,N_5459);
xnor U5930 (N_5930,N_5474,N_5451);
and U5931 (N_5931,N_5286,N_5560);
nor U5932 (N_5932,N_5463,N_5207);
nand U5933 (N_5933,N_5496,N_5426);
xnor U5934 (N_5934,N_5458,N_5553);
nand U5935 (N_5935,N_5380,N_5496);
and U5936 (N_5936,N_5441,N_5255);
nand U5937 (N_5937,N_5438,N_5236);
nand U5938 (N_5938,N_5472,N_5348);
and U5939 (N_5939,N_5409,N_5439);
nand U5940 (N_5940,N_5206,N_5535);
nor U5941 (N_5941,N_5376,N_5480);
nor U5942 (N_5942,N_5236,N_5486);
xnor U5943 (N_5943,N_5485,N_5437);
nand U5944 (N_5944,N_5580,N_5395);
nand U5945 (N_5945,N_5457,N_5554);
or U5946 (N_5946,N_5444,N_5494);
and U5947 (N_5947,N_5567,N_5517);
xor U5948 (N_5948,N_5374,N_5534);
xnor U5949 (N_5949,N_5526,N_5234);
xnor U5950 (N_5950,N_5564,N_5403);
and U5951 (N_5951,N_5384,N_5428);
xnor U5952 (N_5952,N_5516,N_5233);
nor U5953 (N_5953,N_5560,N_5201);
xor U5954 (N_5954,N_5472,N_5389);
xnor U5955 (N_5955,N_5362,N_5285);
or U5956 (N_5956,N_5215,N_5564);
or U5957 (N_5957,N_5557,N_5465);
nor U5958 (N_5958,N_5491,N_5362);
xnor U5959 (N_5959,N_5511,N_5435);
nor U5960 (N_5960,N_5347,N_5318);
nor U5961 (N_5961,N_5249,N_5221);
nor U5962 (N_5962,N_5335,N_5463);
and U5963 (N_5963,N_5318,N_5505);
xor U5964 (N_5964,N_5239,N_5599);
xnor U5965 (N_5965,N_5492,N_5435);
nand U5966 (N_5966,N_5358,N_5580);
and U5967 (N_5967,N_5576,N_5244);
or U5968 (N_5968,N_5224,N_5483);
xor U5969 (N_5969,N_5450,N_5272);
or U5970 (N_5970,N_5428,N_5271);
xor U5971 (N_5971,N_5518,N_5463);
nor U5972 (N_5972,N_5332,N_5315);
or U5973 (N_5973,N_5544,N_5511);
or U5974 (N_5974,N_5295,N_5481);
or U5975 (N_5975,N_5268,N_5261);
and U5976 (N_5976,N_5250,N_5460);
and U5977 (N_5977,N_5595,N_5530);
nand U5978 (N_5978,N_5549,N_5213);
or U5979 (N_5979,N_5232,N_5593);
or U5980 (N_5980,N_5445,N_5433);
nand U5981 (N_5981,N_5438,N_5265);
nand U5982 (N_5982,N_5584,N_5492);
and U5983 (N_5983,N_5599,N_5376);
and U5984 (N_5984,N_5494,N_5334);
nand U5985 (N_5985,N_5579,N_5543);
xnor U5986 (N_5986,N_5514,N_5400);
nand U5987 (N_5987,N_5599,N_5438);
xnor U5988 (N_5988,N_5425,N_5408);
xnor U5989 (N_5989,N_5252,N_5522);
or U5990 (N_5990,N_5335,N_5554);
and U5991 (N_5991,N_5262,N_5279);
xnor U5992 (N_5992,N_5535,N_5567);
nand U5993 (N_5993,N_5366,N_5434);
or U5994 (N_5994,N_5349,N_5202);
and U5995 (N_5995,N_5515,N_5287);
nor U5996 (N_5996,N_5335,N_5409);
or U5997 (N_5997,N_5573,N_5233);
and U5998 (N_5998,N_5377,N_5574);
nor U5999 (N_5999,N_5560,N_5591);
or U6000 (N_6000,N_5678,N_5960);
nor U6001 (N_6001,N_5823,N_5987);
nand U6002 (N_6002,N_5821,N_5742);
xnor U6003 (N_6003,N_5639,N_5635);
nor U6004 (N_6004,N_5619,N_5829);
and U6005 (N_6005,N_5764,N_5672);
nor U6006 (N_6006,N_5618,N_5658);
or U6007 (N_6007,N_5758,N_5608);
nand U6008 (N_6008,N_5709,N_5941);
nand U6009 (N_6009,N_5693,N_5780);
nor U6010 (N_6010,N_5889,N_5686);
nand U6011 (N_6011,N_5797,N_5803);
nor U6012 (N_6012,N_5975,N_5757);
xor U6013 (N_6013,N_5971,N_5914);
nand U6014 (N_6014,N_5982,N_5876);
nor U6015 (N_6015,N_5657,N_5673);
nor U6016 (N_6016,N_5951,N_5827);
nand U6017 (N_6017,N_5986,N_5683);
nand U6018 (N_6018,N_5974,N_5631);
and U6019 (N_6019,N_5706,N_5826);
xnor U6020 (N_6020,N_5893,N_5769);
nand U6021 (N_6021,N_5981,N_5944);
nor U6022 (N_6022,N_5988,N_5729);
and U6023 (N_6023,N_5952,N_5864);
or U6024 (N_6024,N_5701,N_5647);
and U6025 (N_6025,N_5967,N_5909);
or U6026 (N_6026,N_5902,N_5809);
and U6027 (N_6027,N_5853,N_5861);
nor U6028 (N_6028,N_5659,N_5749);
xor U6029 (N_6029,N_5750,N_5817);
or U6030 (N_6030,N_5989,N_5883);
nand U6031 (N_6031,N_5763,N_5807);
or U6032 (N_6032,N_5995,N_5779);
nor U6033 (N_6033,N_5689,N_5910);
nor U6034 (N_6034,N_5813,N_5980);
xnor U6035 (N_6035,N_5816,N_5743);
nor U6036 (N_6036,N_5613,N_5677);
nand U6037 (N_6037,N_5973,N_5945);
nor U6038 (N_6038,N_5690,N_5851);
xnor U6039 (N_6039,N_5640,N_5898);
or U6040 (N_6040,N_5983,N_5928);
nand U6041 (N_6041,N_5887,N_5993);
nand U6042 (N_6042,N_5692,N_5771);
nor U6043 (N_6043,N_5671,N_5783);
nand U6044 (N_6044,N_5992,N_5860);
nor U6045 (N_6045,N_5790,N_5630);
nor U6046 (N_6046,N_5710,N_5832);
nor U6047 (N_6047,N_5956,N_5705);
xor U6048 (N_6048,N_5725,N_5990);
nand U6049 (N_6049,N_5999,N_5994);
xor U6050 (N_6050,N_5962,N_5949);
nand U6051 (N_6051,N_5906,N_5805);
and U6052 (N_6052,N_5676,N_5932);
nand U6053 (N_6053,N_5760,N_5859);
or U6054 (N_6054,N_5824,N_5814);
nor U6055 (N_6055,N_5753,N_5746);
or U6056 (N_6056,N_5789,N_5615);
or U6057 (N_6057,N_5917,N_5822);
nor U6058 (N_6058,N_5724,N_5795);
xor U6059 (N_6059,N_5674,N_5921);
nand U6060 (N_6060,N_5642,N_5651);
and U6061 (N_6061,N_5698,N_5874);
and U6062 (N_6062,N_5890,N_5722);
and U6063 (N_6063,N_5863,N_5648);
xor U6064 (N_6064,N_5935,N_5963);
or U6065 (N_6065,N_5785,N_5804);
nand U6066 (N_6066,N_5778,N_5937);
nand U6067 (N_6067,N_5800,N_5741);
nand U6068 (N_6068,N_5748,N_5977);
or U6069 (N_6069,N_5765,N_5682);
and U6070 (N_6070,N_5793,N_5784);
and U6071 (N_6071,N_5830,N_5633);
xnor U6072 (N_6072,N_5802,N_5862);
and U6073 (N_6073,N_5879,N_5782);
nor U6074 (N_6074,N_5794,N_5601);
or U6075 (N_6075,N_5856,N_5612);
nand U6076 (N_6076,N_5735,N_5786);
nand U6077 (N_6077,N_5711,N_5970);
nor U6078 (N_6078,N_5798,N_5675);
xor U6079 (N_6079,N_5978,N_5972);
nand U6080 (N_6080,N_5926,N_5896);
nor U6081 (N_6081,N_5919,N_5903);
and U6082 (N_6082,N_5702,N_5838);
nand U6083 (N_6083,N_5623,N_5828);
or U6084 (N_6084,N_5628,N_5911);
nand U6085 (N_6085,N_5728,N_5787);
or U6086 (N_6086,N_5907,N_5738);
nor U6087 (N_6087,N_5684,N_5810);
and U6088 (N_6088,N_5607,N_5820);
or U6089 (N_6089,N_5846,N_5897);
xnor U6090 (N_6090,N_5772,N_5718);
and U6091 (N_6091,N_5716,N_5873);
nand U6092 (N_6092,N_5997,N_5894);
xor U6093 (N_6093,N_5913,N_5720);
and U6094 (N_6094,N_5654,N_5609);
xnor U6095 (N_6095,N_5646,N_5842);
nand U6096 (N_6096,N_5796,N_5744);
and U6097 (N_6097,N_5899,N_5708);
xnor U6098 (N_6098,N_5717,N_5611);
xor U6099 (N_6099,N_5695,N_5884);
and U6100 (N_6100,N_5755,N_5959);
nand U6101 (N_6101,N_5957,N_5877);
nand U6102 (N_6102,N_5931,N_5865);
or U6103 (N_6103,N_5681,N_5918);
or U6104 (N_6104,N_5660,N_5900);
and U6105 (N_6105,N_5996,N_5767);
nor U6106 (N_6106,N_5811,N_5621);
nand U6107 (N_6107,N_5691,N_5745);
or U6108 (N_6108,N_5852,N_5979);
or U6109 (N_6109,N_5847,N_5934);
and U6110 (N_6110,N_5849,N_5806);
nand U6111 (N_6111,N_5943,N_5892);
nor U6112 (N_6112,N_5868,N_5948);
nand U6113 (N_6113,N_5679,N_5882);
nor U6114 (N_6114,N_5685,N_5940);
or U6115 (N_6115,N_5662,N_5632);
and U6116 (N_6116,N_5904,N_5819);
and U6117 (N_6117,N_5837,N_5694);
nand U6118 (N_6118,N_5984,N_5953);
nand U6119 (N_6119,N_5622,N_5688);
nand U6120 (N_6120,N_5699,N_5670);
xnor U6121 (N_6121,N_5707,N_5886);
xor U6122 (N_6122,N_5620,N_5704);
or U6123 (N_6123,N_5627,N_5661);
xnor U6124 (N_6124,N_5600,N_5930);
nor U6125 (N_6125,N_5626,N_5730);
and U6126 (N_6126,N_5740,N_5799);
nand U6127 (N_6127,N_5696,N_5713);
or U6128 (N_6128,N_5936,N_5857);
and U6129 (N_6129,N_5650,N_5969);
nor U6130 (N_6130,N_5697,N_5845);
nor U6131 (N_6131,N_5655,N_5739);
or U6132 (N_6132,N_5920,N_5629);
nor U6133 (N_6133,N_5922,N_5766);
or U6134 (N_6134,N_5942,N_5732);
nor U6135 (N_6135,N_5625,N_5715);
and U6136 (N_6136,N_5638,N_5946);
and U6137 (N_6137,N_5924,N_5726);
xnor U6138 (N_6138,N_5666,N_5700);
nor U6139 (N_6139,N_5916,N_5754);
nand U6140 (N_6140,N_5835,N_5881);
xnor U6141 (N_6141,N_5808,N_5653);
nor U6142 (N_6142,N_5905,N_5727);
xnor U6143 (N_6143,N_5938,N_5774);
nor U6144 (N_6144,N_5895,N_5901);
or U6145 (N_6145,N_5850,N_5875);
nor U6146 (N_6146,N_5756,N_5610);
xnor U6147 (N_6147,N_5602,N_5665);
nor U6148 (N_6148,N_5915,N_5663);
or U6149 (N_6149,N_5652,N_5752);
nand U6150 (N_6150,N_5624,N_5606);
or U6151 (N_6151,N_5844,N_5751);
nand U6152 (N_6152,N_5762,N_5954);
nor U6153 (N_6153,N_5734,N_5637);
nand U6154 (N_6154,N_5634,N_5836);
or U6155 (N_6155,N_5761,N_5605);
or U6156 (N_6156,N_5812,N_5776);
xor U6157 (N_6157,N_5645,N_5768);
xnor U6158 (N_6158,N_5891,N_5616);
nand U6159 (N_6159,N_5643,N_5801);
nand U6160 (N_6160,N_5791,N_5933);
nor U6161 (N_6161,N_5719,N_5991);
or U6162 (N_6162,N_5818,N_5976);
nor U6163 (N_6163,N_5964,N_5770);
and U6164 (N_6164,N_5656,N_5958);
nor U6165 (N_6165,N_5733,N_5998);
nand U6166 (N_6166,N_5908,N_5721);
nand U6167 (N_6167,N_5878,N_5888);
and U6168 (N_6168,N_5866,N_5747);
nor U6169 (N_6169,N_5927,N_5985);
or U6170 (N_6170,N_5885,N_5723);
nor U6171 (N_6171,N_5923,N_5736);
or U6172 (N_6172,N_5834,N_5871);
nand U6173 (N_6173,N_5867,N_5870);
nand U6174 (N_6174,N_5947,N_5668);
nor U6175 (N_6175,N_5855,N_5872);
or U6176 (N_6176,N_5703,N_5839);
xnor U6177 (N_6177,N_5649,N_5848);
nor U6178 (N_6178,N_5687,N_5604);
nand U6179 (N_6179,N_5955,N_5667);
nand U6180 (N_6180,N_5759,N_5664);
nand U6181 (N_6181,N_5950,N_5965);
xor U6182 (N_6182,N_5843,N_5788);
or U6183 (N_6183,N_5968,N_5912);
xor U6184 (N_6184,N_5669,N_5731);
and U6185 (N_6185,N_5966,N_5880);
nand U6186 (N_6186,N_5831,N_5636);
or U6187 (N_6187,N_5939,N_5781);
nand U6188 (N_6188,N_5854,N_5617);
or U6189 (N_6189,N_5737,N_5644);
and U6190 (N_6190,N_5714,N_5833);
and U6191 (N_6191,N_5825,N_5858);
or U6192 (N_6192,N_5712,N_5929);
or U6193 (N_6193,N_5603,N_5792);
nand U6194 (N_6194,N_5680,N_5815);
and U6195 (N_6195,N_5775,N_5841);
nand U6196 (N_6196,N_5773,N_5840);
nand U6197 (N_6197,N_5961,N_5869);
or U6198 (N_6198,N_5641,N_5614);
and U6199 (N_6199,N_5777,N_5925);
and U6200 (N_6200,N_5682,N_5779);
or U6201 (N_6201,N_5775,N_5903);
and U6202 (N_6202,N_5957,N_5961);
nand U6203 (N_6203,N_5698,N_5897);
or U6204 (N_6204,N_5909,N_5987);
nor U6205 (N_6205,N_5782,N_5952);
or U6206 (N_6206,N_5932,N_5952);
and U6207 (N_6207,N_5731,N_5941);
xnor U6208 (N_6208,N_5724,N_5679);
nand U6209 (N_6209,N_5932,N_5620);
nor U6210 (N_6210,N_5922,N_5754);
nor U6211 (N_6211,N_5734,N_5738);
or U6212 (N_6212,N_5648,N_5830);
and U6213 (N_6213,N_5707,N_5620);
xor U6214 (N_6214,N_5737,N_5857);
nor U6215 (N_6215,N_5815,N_5771);
and U6216 (N_6216,N_5829,N_5876);
or U6217 (N_6217,N_5745,N_5854);
xor U6218 (N_6218,N_5603,N_5915);
or U6219 (N_6219,N_5868,N_5749);
nor U6220 (N_6220,N_5671,N_5819);
and U6221 (N_6221,N_5678,N_5937);
nor U6222 (N_6222,N_5636,N_5655);
nand U6223 (N_6223,N_5816,N_5846);
nand U6224 (N_6224,N_5763,N_5879);
xor U6225 (N_6225,N_5631,N_5886);
or U6226 (N_6226,N_5824,N_5617);
xor U6227 (N_6227,N_5922,N_5782);
nor U6228 (N_6228,N_5895,N_5890);
nand U6229 (N_6229,N_5934,N_5911);
or U6230 (N_6230,N_5737,N_5944);
xor U6231 (N_6231,N_5961,N_5674);
xnor U6232 (N_6232,N_5890,N_5766);
xor U6233 (N_6233,N_5975,N_5730);
nand U6234 (N_6234,N_5816,N_5833);
xnor U6235 (N_6235,N_5836,N_5614);
nor U6236 (N_6236,N_5869,N_5689);
and U6237 (N_6237,N_5982,N_5774);
xor U6238 (N_6238,N_5905,N_5663);
nor U6239 (N_6239,N_5615,N_5929);
or U6240 (N_6240,N_5904,N_5952);
xor U6241 (N_6241,N_5958,N_5724);
nor U6242 (N_6242,N_5943,N_5940);
nor U6243 (N_6243,N_5895,N_5648);
nand U6244 (N_6244,N_5719,N_5726);
or U6245 (N_6245,N_5702,N_5726);
or U6246 (N_6246,N_5976,N_5754);
xor U6247 (N_6247,N_5617,N_5932);
nor U6248 (N_6248,N_5635,N_5709);
and U6249 (N_6249,N_5876,N_5874);
nand U6250 (N_6250,N_5894,N_5928);
nand U6251 (N_6251,N_5909,N_5682);
and U6252 (N_6252,N_5671,N_5645);
xor U6253 (N_6253,N_5821,N_5612);
nand U6254 (N_6254,N_5748,N_5608);
and U6255 (N_6255,N_5984,N_5977);
nand U6256 (N_6256,N_5966,N_5738);
and U6257 (N_6257,N_5716,N_5905);
xor U6258 (N_6258,N_5676,N_5704);
xor U6259 (N_6259,N_5906,N_5715);
or U6260 (N_6260,N_5778,N_5978);
nand U6261 (N_6261,N_5781,N_5609);
xor U6262 (N_6262,N_5881,N_5938);
nand U6263 (N_6263,N_5726,N_5652);
or U6264 (N_6264,N_5977,N_5738);
nor U6265 (N_6265,N_5775,N_5635);
nor U6266 (N_6266,N_5891,N_5996);
and U6267 (N_6267,N_5835,N_5782);
nand U6268 (N_6268,N_5671,N_5879);
nor U6269 (N_6269,N_5705,N_5788);
or U6270 (N_6270,N_5634,N_5768);
nor U6271 (N_6271,N_5876,N_5760);
and U6272 (N_6272,N_5902,N_5794);
and U6273 (N_6273,N_5641,N_5798);
or U6274 (N_6274,N_5733,N_5610);
and U6275 (N_6275,N_5647,N_5763);
or U6276 (N_6276,N_5918,N_5877);
xnor U6277 (N_6277,N_5611,N_5799);
and U6278 (N_6278,N_5605,N_5620);
or U6279 (N_6279,N_5668,N_5788);
xnor U6280 (N_6280,N_5661,N_5878);
or U6281 (N_6281,N_5981,N_5956);
or U6282 (N_6282,N_5753,N_5745);
nor U6283 (N_6283,N_5963,N_5746);
or U6284 (N_6284,N_5722,N_5800);
nand U6285 (N_6285,N_5704,N_5666);
nor U6286 (N_6286,N_5944,N_5615);
and U6287 (N_6287,N_5797,N_5777);
and U6288 (N_6288,N_5715,N_5984);
or U6289 (N_6289,N_5833,N_5899);
nor U6290 (N_6290,N_5889,N_5655);
or U6291 (N_6291,N_5863,N_5986);
or U6292 (N_6292,N_5869,N_5896);
nand U6293 (N_6293,N_5896,N_5667);
and U6294 (N_6294,N_5685,N_5820);
or U6295 (N_6295,N_5717,N_5884);
nor U6296 (N_6296,N_5992,N_5918);
or U6297 (N_6297,N_5816,N_5651);
and U6298 (N_6298,N_5785,N_5746);
nand U6299 (N_6299,N_5694,N_5867);
or U6300 (N_6300,N_5841,N_5646);
nand U6301 (N_6301,N_5659,N_5877);
xnor U6302 (N_6302,N_5734,N_5858);
nor U6303 (N_6303,N_5658,N_5637);
and U6304 (N_6304,N_5954,N_5850);
nand U6305 (N_6305,N_5674,N_5698);
or U6306 (N_6306,N_5880,N_5663);
xnor U6307 (N_6307,N_5912,N_5995);
xnor U6308 (N_6308,N_5664,N_5836);
xnor U6309 (N_6309,N_5925,N_5749);
nor U6310 (N_6310,N_5894,N_5909);
or U6311 (N_6311,N_5757,N_5725);
or U6312 (N_6312,N_5606,N_5858);
xor U6313 (N_6313,N_5802,N_5956);
nor U6314 (N_6314,N_5981,N_5894);
and U6315 (N_6315,N_5905,N_5855);
nand U6316 (N_6316,N_5678,N_5755);
xor U6317 (N_6317,N_5932,N_5957);
nor U6318 (N_6318,N_5736,N_5948);
nand U6319 (N_6319,N_5941,N_5632);
and U6320 (N_6320,N_5809,N_5832);
nor U6321 (N_6321,N_5635,N_5618);
or U6322 (N_6322,N_5850,N_5751);
or U6323 (N_6323,N_5775,N_5883);
nand U6324 (N_6324,N_5682,N_5676);
and U6325 (N_6325,N_5616,N_5858);
or U6326 (N_6326,N_5915,N_5617);
xor U6327 (N_6327,N_5648,N_5981);
or U6328 (N_6328,N_5802,N_5831);
nand U6329 (N_6329,N_5895,N_5923);
nor U6330 (N_6330,N_5647,N_5640);
nand U6331 (N_6331,N_5848,N_5883);
xnor U6332 (N_6332,N_5886,N_5863);
or U6333 (N_6333,N_5981,N_5821);
or U6334 (N_6334,N_5774,N_5821);
or U6335 (N_6335,N_5995,N_5775);
nand U6336 (N_6336,N_5635,N_5973);
nor U6337 (N_6337,N_5982,N_5742);
and U6338 (N_6338,N_5697,N_5702);
xnor U6339 (N_6339,N_5683,N_5735);
and U6340 (N_6340,N_5715,N_5704);
xor U6341 (N_6341,N_5894,N_5671);
or U6342 (N_6342,N_5768,N_5865);
nand U6343 (N_6343,N_5689,N_5871);
nand U6344 (N_6344,N_5868,N_5865);
or U6345 (N_6345,N_5795,N_5721);
nand U6346 (N_6346,N_5619,N_5902);
or U6347 (N_6347,N_5720,N_5779);
or U6348 (N_6348,N_5779,N_5726);
and U6349 (N_6349,N_5743,N_5923);
nor U6350 (N_6350,N_5638,N_5709);
nand U6351 (N_6351,N_5948,N_5651);
nor U6352 (N_6352,N_5782,N_5681);
nor U6353 (N_6353,N_5859,N_5677);
xor U6354 (N_6354,N_5909,N_5734);
xor U6355 (N_6355,N_5931,N_5899);
and U6356 (N_6356,N_5829,N_5817);
xnor U6357 (N_6357,N_5948,N_5850);
and U6358 (N_6358,N_5925,N_5848);
xnor U6359 (N_6359,N_5689,N_5715);
and U6360 (N_6360,N_5635,N_5628);
nand U6361 (N_6361,N_5727,N_5900);
nor U6362 (N_6362,N_5936,N_5657);
xnor U6363 (N_6363,N_5615,N_5753);
nand U6364 (N_6364,N_5783,N_5745);
or U6365 (N_6365,N_5695,N_5904);
and U6366 (N_6366,N_5814,N_5683);
nor U6367 (N_6367,N_5874,N_5867);
and U6368 (N_6368,N_5947,N_5619);
nand U6369 (N_6369,N_5782,N_5763);
xor U6370 (N_6370,N_5753,N_5712);
and U6371 (N_6371,N_5652,N_5888);
nor U6372 (N_6372,N_5897,N_5619);
nand U6373 (N_6373,N_5622,N_5916);
xnor U6374 (N_6374,N_5661,N_5717);
or U6375 (N_6375,N_5837,N_5904);
nor U6376 (N_6376,N_5839,N_5894);
nand U6377 (N_6377,N_5817,N_5891);
or U6378 (N_6378,N_5697,N_5768);
and U6379 (N_6379,N_5650,N_5628);
and U6380 (N_6380,N_5784,N_5677);
xnor U6381 (N_6381,N_5733,N_5839);
nand U6382 (N_6382,N_5837,N_5878);
nor U6383 (N_6383,N_5726,N_5642);
and U6384 (N_6384,N_5943,N_5977);
or U6385 (N_6385,N_5896,N_5664);
nand U6386 (N_6386,N_5821,N_5654);
nand U6387 (N_6387,N_5769,N_5793);
nand U6388 (N_6388,N_5810,N_5920);
nor U6389 (N_6389,N_5758,N_5737);
or U6390 (N_6390,N_5758,N_5921);
nand U6391 (N_6391,N_5691,N_5847);
and U6392 (N_6392,N_5985,N_5949);
nand U6393 (N_6393,N_5703,N_5773);
xor U6394 (N_6394,N_5941,N_5783);
nand U6395 (N_6395,N_5679,N_5631);
nor U6396 (N_6396,N_5660,N_5724);
nand U6397 (N_6397,N_5877,N_5771);
and U6398 (N_6398,N_5883,N_5717);
nand U6399 (N_6399,N_5989,N_5709);
nor U6400 (N_6400,N_6399,N_6122);
nand U6401 (N_6401,N_6214,N_6375);
xnor U6402 (N_6402,N_6204,N_6275);
nor U6403 (N_6403,N_6007,N_6180);
nand U6404 (N_6404,N_6132,N_6077);
xnor U6405 (N_6405,N_6222,N_6338);
nand U6406 (N_6406,N_6070,N_6333);
nor U6407 (N_6407,N_6182,N_6276);
nand U6408 (N_6408,N_6289,N_6095);
nand U6409 (N_6409,N_6252,N_6133);
or U6410 (N_6410,N_6201,N_6361);
nor U6411 (N_6411,N_6346,N_6358);
nor U6412 (N_6412,N_6374,N_6256);
nor U6413 (N_6413,N_6176,N_6093);
and U6414 (N_6414,N_6061,N_6145);
nor U6415 (N_6415,N_6281,N_6271);
or U6416 (N_6416,N_6000,N_6161);
or U6417 (N_6417,N_6292,N_6310);
and U6418 (N_6418,N_6034,N_6035);
nand U6419 (N_6419,N_6126,N_6384);
nand U6420 (N_6420,N_6189,N_6109);
xnor U6421 (N_6421,N_6187,N_6159);
xnor U6422 (N_6422,N_6389,N_6247);
nor U6423 (N_6423,N_6391,N_6055);
or U6424 (N_6424,N_6112,N_6149);
xnor U6425 (N_6425,N_6316,N_6115);
nor U6426 (N_6426,N_6368,N_6045);
nor U6427 (N_6427,N_6286,N_6010);
xor U6428 (N_6428,N_6359,N_6129);
or U6429 (N_6429,N_6366,N_6317);
and U6430 (N_6430,N_6341,N_6396);
xnor U6431 (N_6431,N_6261,N_6282);
xnor U6432 (N_6432,N_6002,N_6325);
and U6433 (N_6433,N_6337,N_6297);
nor U6434 (N_6434,N_6227,N_6137);
and U6435 (N_6435,N_6198,N_6185);
nand U6436 (N_6436,N_6178,N_6099);
xor U6437 (N_6437,N_6342,N_6335);
nand U6438 (N_6438,N_6081,N_6230);
nand U6439 (N_6439,N_6170,N_6380);
or U6440 (N_6440,N_6283,N_6372);
nand U6441 (N_6441,N_6304,N_6344);
xnor U6442 (N_6442,N_6251,N_6388);
xnor U6443 (N_6443,N_6387,N_6215);
and U6444 (N_6444,N_6195,N_6296);
or U6445 (N_6445,N_6142,N_6078);
xor U6446 (N_6446,N_6197,N_6378);
xor U6447 (N_6447,N_6158,N_6037);
xor U6448 (N_6448,N_6111,N_6280);
or U6449 (N_6449,N_6305,N_6246);
nand U6450 (N_6450,N_6324,N_6373);
nor U6451 (N_6451,N_6011,N_6328);
nand U6452 (N_6452,N_6269,N_6308);
xor U6453 (N_6453,N_6143,N_6274);
nor U6454 (N_6454,N_6021,N_6302);
xor U6455 (N_6455,N_6015,N_6057);
and U6456 (N_6456,N_6395,N_6196);
or U6457 (N_6457,N_6257,N_6311);
and U6458 (N_6458,N_6221,N_6354);
xnor U6459 (N_6459,N_6031,N_6117);
xnor U6460 (N_6460,N_6089,N_6242);
and U6461 (N_6461,N_6295,N_6004);
or U6462 (N_6462,N_6028,N_6082);
nor U6463 (N_6463,N_6014,N_6124);
and U6464 (N_6464,N_6177,N_6162);
xor U6465 (N_6465,N_6160,N_6075);
or U6466 (N_6466,N_6024,N_6234);
or U6467 (N_6467,N_6345,N_6125);
nor U6468 (N_6468,N_6350,N_6202);
xnor U6469 (N_6469,N_6179,N_6226);
and U6470 (N_6470,N_6118,N_6394);
and U6471 (N_6471,N_6138,N_6259);
xor U6472 (N_6472,N_6113,N_6284);
nor U6473 (N_6473,N_6266,N_6065);
and U6474 (N_6474,N_6206,N_6013);
or U6475 (N_6475,N_6131,N_6244);
nor U6476 (N_6476,N_6017,N_6232);
and U6477 (N_6477,N_6123,N_6166);
nor U6478 (N_6478,N_6155,N_6058);
nand U6479 (N_6479,N_6085,N_6083);
and U6480 (N_6480,N_6036,N_6051);
and U6481 (N_6481,N_6139,N_6397);
xnor U6482 (N_6482,N_6285,N_6119);
xnor U6483 (N_6483,N_6114,N_6104);
nand U6484 (N_6484,N_6369,N_6192);
nand U6485 (N_6485,N_6336,N_6249);
and U6486 (N_6486,N_6044,N_6235);
nand U6487 (N_6487,N_6224,N_6025);
and U6488 (N_6488,N_6029,N_6184);
nand U6489 (N_6489,N_6216,N_6203);
and U6490 (N_6490,N_6194,N_6313);
or U6491 (N_6491,N_6248,N_6175);
nor U6492 (N_6492,N_6066,N_6121);
or U6493 (N_6493,N_6091,N_6237);
and U6494 (N_6494,N_6087,N_6217);
or U6495 (N_6495,N_6032,N_6026);
nand U6496 (N_6496,N_6174,N_6183);
or U6497 (N_6497,N_6363,N_6277);
or U6498 (N_6498,N_6098,N_6319);
and U6499 (N_6499,N_6225,N_6103);
nor U6500 (N_6500,N_6233,N_6008);
or U6501 (N_6501,N_6006,N_6127);
nand U6502 (N_6502,N_6146,N_6188);
xor U6503 (N_6503,N_6240,N_6278);
nand U6504 (N_6504,N_6299,N_6253);
nand U6505 (N_6505,N_6339,N_6038);
and U6506 (N_6506,N_6144,N_6264);
nand U6507 (N_6507,N_6209,N_6154);
nor U6508 (N_6508,N_6329,N_6049);
or U6509 (N_6509,N_6043,N_6294);
or U6510 (N_6510,N_6245,N_6106);
and U6511 (N_6511,N_6080,N_6360);
xor U6512 (N_6512,N_6056,N_6054);
nor U6513 (N_6513,N_6268,N_6381);
and U6514 (N_6514,N_6140,N_6067);
nand U6515 (N_6515,N_6348,N_6218);
or U6516 (N_6516,N_6300,N_6063);
or U6517 (N_6517,N_6330,N_6072);
or U6518 (N_6518,N_6255,N_6064);
nor U6519 (N_6519,N_6377,N_6102);
or U6520 (N_6520,N_6150,N_6236);
and U6521 (N_6521,N_6105,N_6141);
and U6522 (N_6522,N_6379,N_6263);
and U6523 (N_6523,N_6041,N_6096);
and U6524 (N_6524,N_6084,N_6211);
and U6525 (N_6525,N_6016,N_6100);
nand U6526 (N_6526,N_6321,N_6207);
xor U6527 (N_6527,N_6250,N_6205);
and U6528 (N_6528,N_6392,N_6301);
nor U6529 (N_6529,N_6241,N_6101);
nand U6530 (N_6530,N_6136,N_6306);
or U6531 (N_6531,N_6298,N_6326);
nor U6532 (N_6532,N_6071,N_6191);
and U6533 (N_6533,N_6092,N_6018);
nand U6534 (N_6534,N_6199,N_6370);
nand U6535 (N_6535,N_6332,N_6110);
nor U6536 (N_6536,N_6398,N_6314);
xnor U6537 (N_6537,N_6153,N_6027);
nand U6538 (N_6538,N_6307,N_6288);
xor U6539 (N_6539,N_6390,N_6164);
and U6540 (N_6540,N_6009,N_6340);
xnor U6541 (N_6541,N_6047,N_6385);
and U6542 (N_6542,N_6135,N_6130);
nand U6543 (N_6543,N_6386,N_6068);
or U6544 (N_6544,N_6267,N_6273);
and U6545 (N_6545,N_6003,N_6254);
nand U6546 (N_6546,N_6312,N_6351);
or U6547 (N_6547,N_6367,N_6291);
and U6548 (N_6548,N_6239,N_6094);
or U6549 (N_6549,N_6327,N_6347);
xor U6550 (N_6550,N_6073,N_6069);
nand U6551 (N_6551,N_6148,N_6362);
or U6552 (N_6552,N_6157,N_6053);
or U6553 (N_6553,N_6005,N_6156);
and U6554 (N_6554,N_6079,N_6279);
xnor U6555 (N_6555,N_6200,N_6076);
or U6556 (N_6556,N_6040,N_6383);
or U6557 (N_6557,N_6393,N_6062);
nor U6558 (N_6558,N_6128,N_6090);
or U6559 (N_6559,N_6356,N_6097);
and U6560 (N_6560,N_6231,N_6039);
and U6561 (N_6561,N_6238,N_6030);
xor U6562 (N_6562,N_6186,N_6376);
nand U6563 (N_6563,N_6151,N_6108);
nand U6564 (N_6564,N_6019,N_6152);
xor U6565 (N_6565,N_6167,N_6318);
nand U6566 (N_6566,N_6220,N_6033);
xor U6567 (N_6567,N_6352,N_6258);
nor U6568 (N_6568,N_6303,N_6213);
nor U6569 (N_6569,N_6353,N_6365);
xnor U6570 (N_6570,N_6042,N_6290);
and U6571 (N_6571,N_6181,N_6208);
xor U6572 (N_6572,N_6270,N_6193);
nor U6573 (N_6573,N_6020,N_6223);
xor U6574 (N_6574,N_6147,N_6371);
and U6575 (N_6575,N_6046,N_6320);
or U6576 (N_6576,N_6265,N_6134);
nor U6577 (N_6577,N_6052,N_6120);
nand U6578 (N_6578,N_6168,N_6169);
nor U6579 (N_6579,N_6364,N_6243);
or U6580 (N_6580,N_6088,N_6229);
nand U6581 (N_6581,N_6001,N_6190);
or U6582 (N_6582,N_6086,N_6309);
or U6583 (N_6583,N_6212,N_6074);
nand U6584 (N_6584,N_6382,N_6323);
or U6585 (N_6585,N_6357,N_6022);
or U6586 (N_6586,N_6272,N_6023);
xnor U6587 (N_6587,N_6260,N_6315);
nor U6588 (N_6588,N_6349,N_6228);
nand U6589 (N_6589,N_6322,N_6171);
nor U6590 (N_6590,N_6163,N_6219);
xor U6591 (N_6591,N_6107,N_6050);
or U6592 (N_6592,N_6343,N_6012);
and U6593 (N_6593,N_6334,N_6172);
or U6594 (N_6594,N_6262,N_6173);
nand U6595 (N_6595,N_6355,N_6287);
or U6596 (N_6596,N_6331,N_6165);
nor U6597 (N_6597,N_6048,N_6059);
nor U6598 (N_6598,N_6116,N_6060);
or U6599 (N_6599,N_6210,N_6293);
or U6600 (N_6600,N_6341,N_6261);
nand U6601 (N_6601,N_6241,N_6214);
nor U6602 (N_6602,N_6262,N_6264);
and U6603 (N_6603,N_6154,N_6057);
nand U6604 (N_6604,N_6343,N_6236);
nand U6605 (N_6605,N_6139,N_6372);
nor U6606 (N_6606,N_6060,N_6098);
and U6607 (N_6607,N_6021,N_6124);
nand U6608 (N_6608,N_6132,N_6330);
xor U6609 (N_6609,N_6176,N_6041);
or U6610 (N_6610,N_6316,N_6399);
or U6611 (N_6611,N_6119,N_6003);
nand U6612 (N_6612,N_6304,N_6033);
or U6613 (N_6613,N_6303,N_6161);
or U6614 (N_6614,N_6041,N_6022);
nor U6615 (N_6615,N_6286,N_6055);
or U6616 (N_6616,N_6342,N_6219);
nand U6617 (N_6617,N_6311,N_6101);
nor U6618 (N_6618,N_6109,N_6267);
nand U6619 (N_6619,N_6168,N_6335);
and U6620 (N_6620,N_6300,N_6254);
xor U6621 (N_6621,N_6277,N_6025);
nor U6622 (N_6622,N_6329,N_6178);
xor U6623 (N_6623,N_6169,N_6277);
nand U6624 (N_6624,N_6024,N_6116);
and U6625 (N_6625,N_6097,N_6398);
xor U6626 (N_6626,N_6355,N_6331);
xnor U6627 (N_6627,N_6244,N_6279);
or U6628 (N_6628,N_6018,N_6012);
or U6629 (N_6629,N_6091,N_6284);
or U6630 (N_6630,N_6093,N_6083);
and U6631 (N_6631,N_6063,N_6082);
nand U6632 (N_6632,N_6171,N_6140);
and U6633 (N_6633,N_6270,N_6272);
nand U6634 (N_6634,N_6287,N_6025);
xnor U6635 (N_6635,N_6320,N_6001);
nor U6636 (N_6636,N_6264,N_6374);
or U6637 (N_6637,N_6349,N_6347);
nor U6638 (N_6638,N_6350,N_6209);
nor U6639 (N_6639,N_6173,N_6167);
or U6640 (N_6640,N_6308,N_6367);
nor U6641 (N_6641,N_6040,N_6368);
and U6642 (N_6642,N_6310,N_6280);
nor U6643 (N_6643,N_6302,N_6244);
nand U6644 (N_6644,N_6045,N_6134);
nor U6645 (N_6645,N_6114,N_6186);
and U6646 (N_6646,N_6287,N_6248);
and U6647 (N_6647,N_6247,N_6268);
and U6648 (N_6648,N_6331,N_6197);
and U6649 (N_6649,N_6193,N_6328);
xnor U6650 (N_6650,N_6127,N_6379);
nand U6651 (N_6651,N_6325,N_6030);
nor U6652 (N_6652,N_6231,N_6340);
and U6653 (N_6653,N_6060,N_6145);
and U6654 (N_6654,N_6237,N_6031);
nor U6655 (N_6655,N_6251,N_6225);
xor U6656 (N_6656,N_6258,N_6194);
or U6657 (N_6657,N_6022,N_6102);
and U6658 (N_6658,N_6161,N_6270);
and U6659 (N_6659,N_6012,N_6387);
or U6660 (N_6660,N_6206,N_6363);
nand U6661 (N_6661,N_6266,N_6396);
xor U6662 (N_6662,N_6223,N_6048);
and U6663 (N_6663,N_6288,N_6366);
and U6664 (N_6664,N_6055,N_6049);
and U6665 (N_6665,N_6289,N_6261);
and U6666 (N_6666,N_6349,N_6243);
or U6667 (N_6667,N_6301,N_6289);
and U6668 (N_6668,N_6329,N_6135);
nand U6669 (N_6669,N_6221,N_6306);
or U6670 (N_6670,N_6275,N_6368);
and U6671 (N_6671,N_6166,N_6249);
nand U6672 (N_6672,N_6296,N_6222);
xor U6673 (N_6673,N_6138,N_6058);
nand U6674 (N_6674,N_6202,N_6329);
and U6675 (N_6675,N_6381,N_6143);
nand U6676 (N_6676,N_6260,N_6214);
xnor U6677 (N_6677,N_6283,N_6245);
and U6678 (N_6678,N_6141,N_6293);
and U6679 (N_6679,N_6115,N_6296);
nand U6680 (N_6680,N_6331,N_6381);
nor U6681 (N_6681,N_6227,N_6251);
nor U6682 (N_6682,N_6045,N_6234);
or U6683 (N_6683,N_6280,N_6253);
or U6684 (N_6684,N_6320,N_6157);
xor U6685 (N_6685,N_6263,N_6082);
nor U6686 (N_6686,N_6395,N_6242);
nor U6687 (N_6687,N_6053,N_6342);
xnor U6688 (N_6688,N_6264,N_6216);
nor U6689 (N_6689,N_6273,N_6184);
nand U6690 (N_6690,N_6079,N_6110);
nor U6691 (N_6691,N_6166,N_6189);
or U6692 (N_6692,N_6283,N_6318);
or U6693 (N_6693,N_6343,N_6009);
nand U6694 (N_6694,N_6304,N_6166);
or U6695 (N_6695,N_6040,N_6180);
nor U6696 (N_6696,N_6239,N_6281);
or U6697 (N_6697,N_6285,N_6334);
and U6698 (N_6698,N_6227,N_6276);
and U6699 (N_6699,N_6231,N_6305);
xor U6700 (N_6700,N_6267,N_6151);
nor U6701 (N_6701,N_6186,N_6380);
nand U6702 (N_6702,N_6288,N_6328);
nor U6703 (N_6703,N_6108,N_6334);
nor U6704 (N_6704,N_6170,N_6335);
xor U6705 (N_6705,N_6324,N_6193);
nor U6706 (N_6706,N_6169,N_6021);
xnor U6707 (N_6707,N_6189,N_6055);
nand U6708 (N_6708,N_6370,N_6284);
or U6709 (N_6709,N_6059,N_6206);
or U6710 (N_6710,N_6296,N_6253);
or U6711 (N_6711,N_6315,N_6030);
nor U6712 (N_6712,N_6182,N_6194);
xnor U6713 (N_6713,N_6213,N_6138);
or U6714 (N_6714,N_6228,N_6130);
and U6715 (N_6715,N_6242,N_6000);
or U6716 (N_6716,N_6060,N_6146);
nor U6717 (N_6717,N_6309,N_6352);
and U6718 (N_6718,N_6134,N_6050);
nand U6719 (N_6719,N_6129,N_6372);
xor U6720 (N_6720,N_6239,N_6152);
nor U6721 (N_6721,N_6385,N_6102);
or U6722 (N_6722,N_6330,N_6198);
and U6723 (N_6723,N_6313,N_6100);
nand U6724 (N_6724,N_6242,N_6262);
and U6725 (N_6725,N_6094,N_6126);
nor U6726 (N_6726,N_6173,N_6104);
nor U6727 (N_6727,N_6102,N_6103);
or U6728 (N_6728,N_6060,N_6261);
nor U6729 (N_6729,N_6204,N_6000);
xor U6730 (N_6730,N_6375,N_6350);
nor U6731 (N_6731,N_6131,N_6114);
or U6732 (N_6732,N_6331,N_6249);
and U6733 (N_6733,N_6167,N_6053);
and U6734 (N_6734,N_6302,N_6223);
or U6735 (N_6735,N_6149,N_6293);
nand U6736 (N_6736,N_6272,N_6003);
xor U6737 (N_6737,N_6215,N_6121);
and U6738 (N_6738,N_6373,N_6332);
nor U6739 (N_6739,N_6283,N_6107);
nor U6740 (N_6740,N_6011,N_6062);
or U6741 (N_6741,N_6323,N_6127);
nand U6742 (N_6742,N_6390,N_6300);
nand U6743 (N_6743,N_6194,N_6041);
xor U6744 (N_6744,N_6312,N_6000);
and U6745 (N_6745,N_6128,N_6359);
nor U6746 (N_6746,N_6027,N_6043);
xor U6747 (N_6747,N_6364,N_6310);
xor U6748 (N_6748,N_6223,N_6060);
xor U6749 (N_6749,N_6378,N_6394);
xnor U6750 (N_6750,N_6377,N_6330);
and U6751 (N_6751,N_6308,N_6154);
nor U6752 (N_6752,N_6104,N_6291);
and U6753 (N_6753,N_6354,N_6397);
nor U6754 (N_6754,N_6124,N_6244);
nand U6755 (N_6755,N_6388,N_6051);
or U6756 (N_6756,N_6273,N_6383);
xnor U6757 (N_6757,N_6296,N_6368);
nand U6758 (N_6758,N_6071,N_6379);
nor U6759 (N_6759,N_6101,N_6350);
xor U6760 (N_6760,N_6167,N_6399);
xnor U6761 (N_6761,N_6127,N_6363);
nand U6762 (N_6762,N_6027,N_6392);
nand U6763 (N_6763,N_6124,N_6051);
xnor U6764 (N_6764,N_6042,N_6071);
nor U6765 (N_6765,N_6097,N_6110);
or U6766 (N_6766,N_6150,N_6282);
xor U6767 (N_6767,N_6063,N_6269);
nor U6768 (N_6768,N_6296,N_6118);
or U6769 (N_6769,N_6196,N_6398);
nand U6770 (N_6770,N_6015,N_6350);
xnor U6771 (N_6771,N_6186,N_6389);
and U6772 (N_6772,N_6150,N_6109);
nand U6773 (N_6773,N_6346,N_6344);
or U6774 (N_6774,N_6176,N_6284);
and U6775 (N_6775,N_6058,N_6031);
xor U6776 (N_6776,N_6271,N_6232);
nand U6777 (N_6777,N_6134,N_6136);
nor U6778 (N_6778,N_6229,N_6398);
or U6779 (N_6779,N_6187,N_6161);
and U6780 (N_6780,N_6261,N_6065);
xor U6781 (N_6781,N_6290,N_6261);
nand U6782 (N_6782,N_6157,N_6044);
nor U6783 (N_6783,N_6266,N_6225);
xor U6784 (N_6784,N_6313,N_6358);
or U6785 (N_6785,N_6178,N_6054);
or U6786 (N_6786,N_6207,N_6299);
and U6787 (N_6787,N_6255,N_6173);
nand U6788 (N_6788,N_6218,N_6129);
or U6789 (N_6789,N_6172,N_6113);
or U6790 (N_6790,N_6030,N_6080);
nand U6791 (N_6791,N_6058,N_6246);
and U6792 (N_6792,N_6342,N_6331);
xnor U6793 (N_6793,N_6220,N_6016);
nand U6794 (N_6794,N_6322,N_6116);
xor U6795 (N_6795,N_6316,N_6251);
nor U6796 (N_6796,N_6083,N_6069);
xnor U6797 (N_6797,N_6347,N_6053);
nor U6798 (N_6798,N_6267,N_6078);
xnor U6799 (N_6799,N_6047,N_6096);
and U6800 (N_6800,N_6526,N_6433);
or U6801 (N_6801,N_6589,N_6746);
nand U6802 (N_6802,N_6451,N_6727);
and U6803 (N_6803,N_6584,N_6464);
nand U6804 (N_6804,N_6428,N_6674);
or U6805 (N_6805,N_6681,N_6752);
and U6806 (N_6806,N_6569,N_6778);
and U6807 (N_6807,N_6643,N_6436);
nand U6808 (N_6808,N_6583,N_6705);
and U6809 (N_6809,N_6521,N_6505);
nor U6810 (N_6810,N_6604,N_6517);
nand U6811 (N_6811,N_6599,N_6425);
or U6812 (N_6812,N_6788,N_6651);
or U6813 (N_6813,N_6603,N_6668);
or U6814 (N_6814,N_6633,N_6733);
xnor U6815 (N_6815,N_6795,N_6781);
xor U6816 (N_6816,N_6424,N_6406);
and U6817 (N_6817,N_6680,N_6468);
or U6818 (N_6818,N_6774,N_6782);
or U6819 (N_6819,N_6528,N_6465);
and U6820 (N_6820,N_6435,N_6707);
nor U6821 (N_6821,N_6783,N_6462);
and U6822 (N_6822,N_6459,N_6729);
and U6823 (N_6823,N_6497,N_6485);
nand U6824 (N_6824,N_6504,N_6749);
xor U6825 (N_6825,N_6780,N_6500);
and U6826 (N_6826,N_6514,N_6690);
and U6827 (N_6827,N_6540,N_6760);
nor U6828 (N_6828,N_6405,N_6686);
or U6829 (N_6829,N_6693,N_6565);
nor U6830 (N_6830,N_6796,N_6522);
xor U6831 (N_6831,N_6562,N_6661);
nor U6832 (N_6832,N_6732,N_6560);
nand U6833 (N_6833,N_6445,N_6508);
or U6834 (N_6834,N_6620,N_6640);
nor U6835 (N_6835,N_6775,N_6646);
xor U6836 (N_6836,N_6726,N_6506);
or U6837 (N_6837,N_6471,N_6472);
xor U6838 (N_6838,N_6502,N_6558);
xnor U6839 (N_6839,N_6654,N_6607);
or U6840 (N_6840,N_6738,N_6568);
nand U6841 (N_6841,N_6722,N_6701);
and U6842 (N_6842,N_6615,N_6657);
or U6843 (N_6843,N_6402,N_6757);
nor U6844 (N_6844,N_6717,N_6623);
and U6845 (N_6845,N_6437,N_6688);
nor U6846 (N_6846,N_6422,N_6696);
nand U6847 (N_6847,N_6564,N_6672);
xnor U6848 (N_6848,N_6684,N_6475);
nor U6849 (N_6849,N_6700,N_6789);
and U6850 (N_6850,N_6546,N_6534);
and U6851 (N_6851,N_6751,N_6593);
nand U6852 (N_6852,N_6638,N_6682);
nor U6853 (N_6853,N_6737,N_6404);
xor U6854 (N_6854,N_6645,N_6531);
nand U6855 (N_6855,N_6659,N_6578);
or U6856 (N_6856,N_6719,N_6739);
nor U6857 (N_6857,N_6523,N_6588);
or U6858 (N_6858,N_6652,N_6592);
nor U6859 (N_6859,N_6618,N_6772);
and U6860 (N_6860,N_6622,N_6755);
nand U6861 (N_6861,N_6676,N_6527);
and U6862 (N_6862,N_6694,N_6456);
or U6863 (N_6863,N_6492,N_6720);
xnor U6864 (N_6864,N_6476,N_6799);
xnor U6865 (N_6865,N_6455,N_6725);
nand U6866 (N_6866,N_6621,N_6577);
nor U6867 (N_6867,N_6642,N_6488);
nor U6868 (N_6868,N_6677,N_6709);
nor U6869 (N_6869,N_6473,N_6625);
xor U6870 (N_6870,N_6596,N_6634);
nor U6871 (N_6871,N_6703,N_6450);
xnor U6872 (N_6872,N_6507,N_6552);
nor U6873 (N_6873,N_6470,N_6770);
xnor U6874 (N_6874,N_6605,N_6617);
or U6875 (N_6875,N_6535,N_6417);
and U6876 (N_6876,N_6484,N_6438);
and U6877 (N_6877,N_6594,N_6670);
and U6878 (N_6878,N_6411,N_6637);
nor U6879 (N_6879,N_6478,N_6763);
nand U6880 (N_6880,N_6667,N_6631);
or U6881 (N_6881,N_6793,N_6499);
and U6882 (N_6882,N_6481,N_6415);
xnor U6883 (N_6883,N_6699,N_6792);
xnor U6884 (N_6884,N_6443,N_6414);
nand U6885 (N_6885,N_6477,N_6590);
or U6886 (N_6886,N_6446,N_6791);
nand U6887 (N_6887,N_6786,N_6734);
nand U6888 (N_6888,N_6754,N_6427);
xor U6889 (N_6889,N_6494,N_6773);
xor U6890 (N_6890,N_6602,N_6544);
nand U6891 (N_6891,N_6479,N_6591);
and U6892 (N_6892,N_6495,N_6416);
nand U6893 (N_6893,N_6610,N_6624);
xnor U6894 (N_6894,N_6745,N_6660);
xnor U6895 (N_6895,N_6777,N_6553);
nor U6896 (N_6896,N_6491,N_6790);
and U6897 (N_6897,N_6431,N_6794);
nor U6898 (N_6898,N_6650,N_6413);
or U6899 (N_6899,N_6410,N_6501);
and U6900 (N_6900,N_6766,N_6555);
xor U6901 (N_6901,N_6718,N_6515);
and U6902 (N_6902,N_6665,N_6741);
xor U6903 (N_6903,N_6616,N_6639);
nor U6904 (N_6904,N_6430,N_6510);
nand U6905 (N_6905,N_6635,N_6641);
xnor U6906 (N_6906,N_6532,N_6440);
nand U6907 (N_6907,N_6750,N_6454);
nand U6908 (N_6908,N_6611,N_6708);
nor U6909 (N_6909,N_6776,N_6675);
or U6910 (N_6910,N_6669,N_6606);
nand U6911 (N_6911,N_6516,N_6697);
and U6912 (N_6912,N_6715,N_6600);
and U6913 (N_6913,N_6758,N_6448);
nor U6914 (N_6914,N_6740,N_6408);
nor U6915 (N_6915,N_6647,N_6545);
xnor U6916 (N_6916,N_6573,N_6664);
nor U6917 (N_6917,N_6487,N_6711);
and U6918 (N_6918,N_6762,N_6756);
and U6919 (N_6919,N_6539,N_6743);
and U6920 (N_6920,N_6530,N_6721);
or U6921 (N_6921,N_6400,N_6561);
xnor U6922 (N_6922,N_6649,N_6550);
and U6923 (N_6923,N_6666,N_6679);
xor U6924 (N_6924,N_6689,N_6761);
or U6925 (N_6925,N_6627,N_6458);
or U6926 (N_6926,N_6768,N_6582);
xor U6927 (N_6927,N_6467,N_6630);
nor U6928 (N_6928,N_6662,N_6658);
and U6929 (N_6929,N_6636,N_6538);
nand U6930 (N_6930,N_6798,N_6692);
nand U6931 (N_6931,N_6695,N_6403);
nand U6932 (N_6932,N_6572,N_6742);
xor U6933 (N_6933,N_6779,N_6629);
xor U6934 (N_6934,N_6432,N_6595);
and U6935 (N_6935,N_6698,N_6714);
and U6936 (N_6936,N_6576,N_6784);
nand U6937 (N_6937,N_6482,N_6736);
or U6938 (N_6938,N_6673,N_6469);
or U6939 (N_6939,N_6614,N_6474);
nand U6940 (N_6940,N_6656,N_6712);
or U6941 (N_6941,N_6747,N_6765);
xnor U6942 (N_6942,N_6575,N_6567);
and U6943 (N_6943,N_6483,N_6529);
xnor U6944 (N_6944,N_6728,N_6498);
nor U6945 (N_6945,N_6524,N_6628);
nor U6946 (N_6946,N_6493,N_6644);
xnor U6947 (N_6947,N_6759,N_6787);
nand U6948 (N_6948,N_6706,N_6547);
or U6949 (N_6949,N_6574,N_6556);
nor U6950 (N_6950,N_6587,N_6519);
or U6951 (N_6951,N_6449,N_6598);
xor U6952 (N_6952,N_6678,N_6511);
nor U6953 (N_6953,N_6426,N_6581);
or U6954 (N_6954,N_6585,N_6429);
and U6955 (N_6955,N_6542,N_6533);
xnor U6956 (N_6956,N_6744,N_6580);
or U6957 (N_6957,N_6608,N_6704);
xor U6958 (N_6958,N_6723,N_6730);
nor U6959 (N_6959,N_6420,N_6683);
and U6960 (N_6960,N_6549,N_6489);
and U6961 (N_6961,N_6586,N_6518);
xnor U6962 (N_6962,N_6447,N_6653);
and U6963 (N_6963,N_6626,N_6543);
xor U6964 (N_6964,N_6563,N_6566);
nor U6965 (N_6965,N_6655,N_6771);
nand U6966 (N_6966,N_6444,N_6503);
nand U6967 (N_6967,N_6731,N_6724);
nand U6968 (N_6968,N_6463,N_6579);
nor U6969 (N_6969,N_6466,N_6713);
nand U6970 (N_6970,N_6513,N_6486);
nand U6971 (N_6971,N_6496,N_6439);
or U6972 (N_6972,N_6559,N_6612);
nor U6973 (N_6973,N_6434,N_6457);
and U6974 (N_6974,N_6442,N_6460);
nor U6975 (N_6975,N_6785,N_6702);
and U6976 (N_6976,N_6548,N_6419);
nand U6977 (N_6977,N_6541,N_6480);
and U6978 (N_6978,N_6648,N_6797);
nand U6979 (N_6979,N_6452,N_6418);
nand U6980 (N_6980,N_6710,N_6537);
nand U6981 (N_6981,N_6685,N_6735);
nor U6982 (N_6982,N_6716,N_6409);
nor U6983 (N_6983,N_6609,N_6570);
and U6984 (N_6984,N_6401,N_6571);
nor U6985 (N_6985,N_6554,N_6421);
or U6986 (N_6986,N_6490,N_6767);
nand U6987 (N_6987,N_6441,N_6619);
and U6988 (N_6988,N_6525,N_6764);
or U6989 (N_6989,N_6663,N_6407);
or U6990 (N_6990,N_6748,N_6632);
nor U6991 (N_6991,N_6691,N_6551);
or U6992 (N_6992,N_6512,N_6601);
or U6993 (N_6993,N_6597,N_6557);
and U6994 (N_6994,N_6687,N_6461);
nor U6995 (N_6995,N_6753,N_6536);
or U6996 (N_6996,N_6412,N_6423);
and U6997 (N_6997,N_6769,N_6671);
nand U6998 (N_6998,N_6509,N_6520);
xnor U6999 (N_6999,N_6453,N_6613);
or U7000 (N_7000,N_6424,N_6774);
and U7001 (N_7001,N_6584,N_6478);
xor U7002 (N_7002,N_6799,N_6781);
nand U7003 (N_7003,N_6770,N_6600);
xnor U7004 (N_7004,N_6469,N_6773);
nor U7005 (N_7005,N_6733,N_6657);
nor U7006 (N_7006,N_6548,N_6445);
nand U7007 (N_7007,N_6793,N_6789);
or U7008 (N_7008,N_6785,N_6787);
and U7009 (N_7009,N_6526,N_6558);
xnor U7010 (N_7010,N_6694,N_6761);
or U7011 (N_7011,N_6685,N_6773);
and U7012 (N_7012,N_6751,N_6753);
xnor U7013 (N_7013,N_6528,N_6478);
xor U7014 (N_7014,N_6444,N_6471);
xnor U7015 (N_7015,N_6662,N_6558);
nor U7016 (N_7016,N_6752,N_6709);
nor U7017 (N_7017,N_6459,N_6565);
xor U7018 (N_7018,N_6401,N_6788);
xor U7019 (N_7019,N_6473,N_6471);
and U7020 (N_7020,N_6649,N_6646);
xnor U7021 (N_7021,N_6758,N_6530);
or U7022 (N_7022,N_6420,N_6481);
xor U7023 (N_7023,N_6733,N_6715);
nor U7024 (N_7024,N_6606,N_6565);
nor U7025 (N_7025,N_6510,N_6764);
or U7026 (N_7026,N_6438,N_6756);
xnor U7027 (N_7027,N_6575,N_6660);
nand U7028 (N_7028,N_6748,N_6656);
xor U7029 (N_7029,N_6480,N_6537);
xnor U7030 (N_7030,N_6428,N_6608);
or U7031 (N_7031,N_6564,N_6431);
or U7032 (N_7032,N_6658,N_6735);
and U7033 (N_7033,N_6665,N_6539);
xor U7034 (N_7034,N_6795,N_6771);
nand U7035 (N_7035,N_6491,N_6468);
or U7036 (N_7036,N_6454,N_6549);
and U7037 (N_7037,N_6548,N_6494);
nand U7038 (N_7038,N_6596,N_6754);
nand U7039 (N_7039,N_6520,N_6484);
nand U7040 (N_7040,N_6680,N_6588);
nand U7041 (N_7041,N_6617,N_6753);
nor U7042 (N_7042,N_6659,N_6586);
and U7043 (N_7043,N_6471,N_6468);
nand U7044 (N_7044,N_6481,N_6697);
and U7045 (N_7045,N_6795,N_6445);
nor U7046 (N_7046,N_6772,N_6420);
nand U7047 (N_7047,N_6507,N_6524);
and U7048 (N_7048,N_6508,N_6434);
and U7049 (N_7049,N_6638,N_6599);
and U7050 (N_7050,N_6548,N_6541);
xnor U7051 (N_7051,N_6659,N_6753);
and U7052 (N_7052,N_6766,N_6601);
or U7053 (N_7053,N_6488,N_6593);
xnor U7054 (N_7054,N_6551,N_6451);
or U7055 (N_7055,N_6711,N_6413);
nor U7056 (N_7056,N_6771,N_6686);
or U7057 (N_7057,N_6521,N_6768);
or U7058 (N_7058,N_6764,N_6707);
nor U7059 (N_7059,N_6498,N_6612);
nand U7060 (N_7060,N_6728,N_6677);
or U7061 (N_7061,N_6551,N_6502);
nor U7062 (N_7062,N_6478,N_6448);
xor U7063 (N_7063,N_6521,N_6734);
or U7064 (N_7064,N_6621,N_6473);
xor U7065 (N_7065,N_6789,N_6564);
nor U7066 (N_7066,N_6689,N_6724);
and U7067 (N_7067,N_6615,N_6720);
nand U7068 (N_7068,N_6505,N_6403);
nand U7069 (N_7069,N_6463,N_6646);
or U7070 (N_7070,N_6446,N_6569);
and U7071 (N_7071,N_6664,N_6670);
nand U7072 (N_7072,N_6604,N_6502);
nor U7073 (N_7073,N_6723,N_6606);
xnor U7074 (N_7074,N_6403,N_6749);
nand U7075 (N_7075,N_6610,N_6628);
nor U7076 (N_7076,N_6736,N_6429);
nand U7077 (N_7077,N_6669,N_6524);
nor U7078 (N_7078,N_6658,N_6497);
xnor U7079 (N_7079,N_6622,N_6490);
nor U7080 (N_7080,N_6683,N_6546);
and U7081 (N_7081,N_6758,N_6450);
nor U7082 (N_7082,N_6461,N_6718);
or U7083 (N_7083,N_6699,N_6683);
xnor U7084 (N_7084,N_6532,N_6645);
or U7085 (N_7085,N_6577,N_6589);
nand U7086 (N_7086,N_6670,N_6435);
or U7087 (N_7087,N_6478,N_6693);
nor U7088 (N_7088,N_6733,N_6680);
or U7089 (N_7089,N_6750,N_6680);
and U7090 (N_7090,N_6779,N_6543);
nor U7091 (N_7091,N_6500,N_6448);
nor U7092 (N_7092,N_6673,N_6604);
or U7093 (N_7093,N_6475,N_6498);
and U7094 (N_7094,N_6649,N_6777);
or U7095 (N_7095,N_6572,N_6588);
and U7096 (N_7096,N_6523,N_6791);
nand U7097 (N_7097,N_6422,N_6599);
and U7098 (N_7098,N_6472,N_6631);
xor U7099 (N_7099,N_6485,N_6618);
xor U7100 (N_7100,N_6762,N_6523);
nand U7101 (N_7101,N_6419,N_6400);
or U7102 (N_7102,N_6649,N_6753);
nand U7103 (N_7103,N_6710,N_6463);
nand U7104 (N_7104,N_6574,N_6455);
or U7105 (N_7105,N_6790,N_6486);
nor U7106 (N_7106,N_6615,N_6675);
nor U7107 (N_7107,N_6799,N_6410);
and U7108 (N_7108,N_6660,N_6673);
nor U7109 (N_7109,N_6546,N_6780);
nor U7110 (N_7110,N_6710,N_6566);
and U7111 (N_7111,N_6509,N_6449);
nor U7112 (N_7112,N_6687,N_6647);
or U7113 (N_7113,N_6490,N_6713);
nor U7114 (N_7114,N_6521,N_6451);
nor U7115 (N_7115,N_6779,N_6588);
and U7116 (N_7116,N_6401,N_6789);
xor U7117 (N_7117,N_6534,N_6568);
nor U7118 (N_7118,N_6543,N_6466);
nor U7119 (N_7119,N_6669,N_6487);
nand U7120 (N_7120,N_6755,N_6726);
nand U7121 (N_7121,N_6773,N_6544);
and U7122 (N_7122,N_6658,N_6580);
xnor U7123 (N_7123,N_6555,N_6496);
and U7124 (N_7124,N_6666,N_6639);
and U7125 (N_7125,N_6470,N_6416);
nand U7126 (N_7126,N_6733,N_6735);
or U7127 (N_7127,N_6526,N_6506);
or U7128 (N_7128,N_6780,N_6482);
nor U7129 (N_7129,N_6665,N_6739);
nand U7130 (N_7130,N_6481,N_6540);
and U7131 (N_7131,N_6770,N_6579);
or U7132 (N_7132,N_6619,N_6643);
xnor U7133 (N_7133,N_6633,N_6663);
xor U7134 (N_7134,N_6640,N_6416);
and U7135 (N_7135,N_6604,N_6647);
nand U7136 (N_7136,N_6456,N_6670);
xor U7137 (N_7137,N_6613,N_6591);
and U7138 (N_7138,N_6425,N_6716);
nand U7139 (N_7139,N_6789,N_6460);
xnor U7140 (N_7140,N_6553,N_6722);
and U7141 (N_7141,N_6791,N_6425);
xnor U7142 (N_7142,N_6604,N_6675);
xnor U7143 (N_7143,N_6744,N_6445);
or U7144 (N_7144,N_6554,N_6592);
xnor U7145 (N_7145,N_6604,N_6639);
nor U7146 (N_7146,N_6754,N_6749);
nand U7147 (N_7147,N_6648,N_6763);
xor U7148 (N_7148,N_6573,N_6770);
or U7149 (N_7149,N_6643,N_6705);
and U7150 (N_7150,N_6466,N_6456);
nand U7151 (N_7151,N_6522,N_6737);
nor U7152 (N_7152,N_6500,N_6457);
nor U7153 (N_7153,N_6542,N_6532);
nor U7154 (N_7154,N_6513,N_6745);
and U7155 (N_7155,N_6659,N_6521);
nand U7156 (N_7156,N_6437,N_6776);
nor U7157 (N_7157,N_6689,N_6785);
nor U7158 (N_7158,N_6415,N_6783);
xor U7159 (N_7159,N_6577,N_6669);
and U7160 (N_7160,N_6786,N_6559);
nor U7161 (N_7161,N_6527,N_6473);
nor U7162 (N_7162,N_6675,N_6750);
nor U7163 (N_7163,N_6623,N_6755);
and U7164 (N_7164,N_6621,N_6439);
or U7165 (N_7165,N_6740,N_6778);
and U7166 (N_7166,N_6732,N_6725);
or U7167 (N_7167,N_6773,N_6550);
or U7168 (N_7168,N_6440,N_6408);
and U7169 (N_7169,N_6706,N_6778);
and U7170 (N_7170,N_6578,N_6454);
xnor U7171 (N_7171,N_6443,N_6698);
nor U7172 (N_7172,N_6605,N_6742);
xnor U7173 (N_7173,N_6630,N_6549);
nor U7174 (N_7174,N_6508,N_6794);
nand U7175 (N_7175,N_6789,N_6729);
or U7176 (N_7176,N_6637,N_6709);
and U7177 (N_7177,N_6658,N_6561);
nor U7178 (N_7178,N_6653,N_6545);
or U7179 (N_7179,N_6511,N_6642);
or U7180 (N_7180,N_6577,N_6620);
nand U7181 (N_7181,N_6415,N_6689);
or U7182 (N_7182,N_6469,N_6489);
nand U7183 (N_7183,N_6672,N_6778);
xor U7184 (N_7184,N_6735,N_6631);
or U7185 (N_7185,N_6407,N_6550);
or U7186 (N_7186,N_6508,N_6590);
xnor U7187 (N_7187,N_6792,N_6697);
xor U7188 (N_7188,N_6501,N_6489);
xor U7189 (N_7189,N_6667,N_6421);
nor U7190 (N_7190,N_6704,N_6493);
and U7191 (N_7191,N_6737,N_6722);
xnor U7192 (N_7192,N_6656,N_6670);
xnor U7193 (N_7193,N_6762,N_6522);
nor U7194 (N_7194,N_6694,N_6562);
xor U7195 (N_7195,N_6635,N_6728);
nand U7196 (N_7196,N_6778,N_6654);
or U7197 (N_7197,N_6761,N_6492);
or U7198 (N_7198,N_6775,N_6562);
or U7199 (N_7199,N_6692,N_6540);
nand U7200 (N_7200,N_6857,N_7071);
or U7201 (N_7201,N_6994,N_6827);
or U7202 (N_7202,N_7085,N_6880);
nor U7203 (N_7203,N_6872,N_6839);
and U7204 (N_7204,N_6978,N_7082);
nand U7205 (N_7205,N_6855,N_6930);
nor U7206 (N_7206,N_7099,N_6992);
nor U7207 (N_7207,N_7007,N_6884);
and U7208 (N_7208,N_7077,N_7027);
and U7209 (N_7209,N_6902,N_6996);
nor U7210 (N_7210,N_7095,N_7135);
nor U7211 (N_7211,N_6854,N_6966);
nand U7212 (N_7212,N_6892,N_7032);
nand U7213 (N_7213,N_6981,N_7106);
and U7214 (N_7214,N_7115,N_7096);
xnor U7215 (N_7215,N_7014,N_7100);
or U7216 (N_7216,N_6985,N_7010);
and U7217 (N_7217,N_7108,N_6976);
or U7218 (N_7218,N_7046,N_7073);
nand U7219 (N_7219,N_7044,N_7145);
nor U7220 (N_7220,N_6899,N_6968);
and U7221 (N_7221,N_6943,N_7016);
nor U7222 (N_7222,N_6871,N_6831);
nand U7223 (N_7223,N_7158,N_6998);
or U7224 (N_7224,N_7024,N_6832);
nor U7225 (N_7225,N_6838,N_7191);
nand U7226 (N_7226,N_7011,N_7107);
xnor U7227 (N_7227,N_7043,N_6882);
and U7228 (N_7228,N_7150,N_7171);
and U7229 (N_7229,N_6819,N_7136);
xnor U7230 (N_7230,N_7009,N_7058);
xnor U7231 (N_7231,N_7002,N_7160);
xnor U7232 (N_7232,N_7003,N_6843);
and U7233 (N_7233,N_7091,N_7086);
nand U7234 (N_7234,N_7124,N_7176);
and U7235 (N_7235,N_7051,N_6970);
and U7236 (N_7236,N_6858,N_6807);
or U7237 (N_7237,N_7035,N_6802);
and U7238 (N_7238,N_7052,N_6964);
or U7239 (N_7239,N_7164,N_7156);
nand U7240 (N_7240,N_7129,N_6864);
nor U7241 (N_7241,N_7074,N_7159);
nand U7242 (N_7242,N_7059,N_7126);
nor U7243 (N_7243,N_7199,N_6820);
nor U7244 (N_7244,N_7192,N_6954);
nor U7245 (N_7245,N_6979,N_7036);
and U7246 (N_7246,N_6921,N_7012);
or U7247 (N_7247,N_7087,N_7068);
and U7248 (N_7248,N_7019,N_6801);
nand U7249 (N_7249,N_6957,N_6849);
nor U7250 (N_7250,N_6949,N_7110);
or U7251 (N_7251,N_6861,N_6947);
nor U7252 (N_7252,N_7067,N_7081);
nand U7253 (N_7253,N_6823,N_7170);
or U7254 (N_7254,N_7195,N_6980);
or U7255 (N_7255,N_7064,N_7181);
or U7256 (N_7256,N_7113,N_7117);
and U7257 (N_7257,N_6893,N_7182);
nor U7258 (N_7258,N_6983,N_7013);
and U7259 (N_7259,N_6973,N_7188);
and U7260 (N_7260,N_6925,N_6960);
nand U7261 (N_7261,N_6920,N_7140);
nand U7262 (N_7262,N_6805,N_7193);
or U7263 (N_7263,N_6800,N_6837);
xnor U7264 (N_7264,N_7054,N_6876);
nand U7265 (N_7265,N_6944,N_7139);
nand U7266 (N_7266,N_6900,N_6914);
or U7267 (N_7267,N_6834,N_7184);
xor U7268 (N_7268,N_6886,N_6939);
and U7269 (N_7269,N_7090,N_6821);
nor U7270 (N_7270,N_7190,N_6896);
nand U7271 (N_7271,N_7093,N_6905);
nand U7272 (N_7272,N_7165,N_7120);
nor U7273 (N_7273,N_7174,N_6867);
and U7274 (N_7274,N_6847,N_6895);
and U7275 (N_7275,N_7157,N_7004);
nor U7276 (N_7276,N_6814,N_7080);
and U7277 (N_7277,N_7050,N_6803);
and U7278 (N_7278,N_6956,N_6937);
and U7279 (N_7279,N_6917,N_6927);
and U7280 (N_7280,N_6863,N_6933);
nor U7281 (N_7281,N_6824,N_6915);
or U7282 (N_7282,N_6999,N_7161);
nor U7283 (N_7283,N_7154,N_6894);
nand U7284 (N_7284,N_6975,N_6942);
nand U7285 (N_7285,N_7057,N_7053);
xor U7286 (N_7286,N_7178,N_7006);
xor U7287 (N_7287,N_7169,N_7063);
nor U7288 (N_7288,N_7127,N_6878);
nor U7289 (N_7289,N_6963,N_6989);
nand U7290 (N_7290,N_7076,N_6918);
and U7291 (N_7291,N_6982,N_7128);
nand U7292 (N_7292,N_6815,N_7103);
nand U7293 (N_7293,N_7070,N_7065);
and U7294 (N_7294,N_6889,N_7196);
nand U7295 (N_7295,N_6868,N_7062);
and U7296 (N_7296,N_6840,N_6959);
and U7297 (N_7297,N_7031,N_6833);
nor U7298 (N_7298,N_6897,N_6935);
or U7299 (N_7299,N_6919,N_7029);
or U7300 (N_7300,N_7147,N_6958);
and U7301 (N_7301,N_7079,N_6859);
xor U7302 (N_7302,N_7055,N_7026);
or U7303 (N_7303,N_7000,N_6810);
and U7304 (N_7304,N_7021,N_6940);
xor U7305 (N_7305,N_6852,N_7069);
nor U7306 (N_7306,N_7134,N_6813);
or U7307 (N_7307,N_6997,N_6984);
xnor U7308 (N_7308,N_7109,N_6865);
nor U7309 (N_7309,N_7123,N_7111);
and U7310 (N_7310,N_7173,N_7001);
or U7311 (N_7311,N_7028,N_7149);
or U7312 (N_7312,N_6869,N_7179);
and U7313 (N_7313,N_7125,N_6913);
nor U7314 (N_7314,N_7180,N_6846);
xor U7315 (N_7315,N_6866,N_6931);
xnor U7316 (N_7316,N_6906,N_6951);
and U7317 (N_7317,N_6990,N_7017);
xor U7318 (N_7318,N_6972,N_6853);
nor U7319 (N_7319,N_6928,N_7133);
or U7320 (N_7320,N_7020,N_6946);
or U7321 (N_7321,N_7039,N_7097);
or U7322 (N_7322,N_6829,N_7137);
nor U7323 (N_7323,N_7033,N_6874);
nand U7324 (N_7324,N_6808,N_6873);
or U7325 (N_7325,N_6870,N_6890);
or U7326 (N_7326,N_7185,N_6862);
or U7327 (N_7327,N_6850,N_6883);
nor U7328 (N_7328,N_7018,N_7121);
xor U7329 (N_7329,N_6891,N_6887);
nor U7330 (N_7330,N_6825,N_7116);
nor U7331 (N_7331,N_6811,N_7198);
xnor U7332 (N_7332,N_6877,N_6822);
and U7333 (N_7333,N_6961,N_7155);
nor U7334 (N_7334,N_7168,N_6851);
nor U7335 (N_7335,N_6948,N_6924);
xnor U7336 (N_7336,N_7061,N_6836);
nand U7337 (N_7337,N_7008,N_6929);
or U7338 (N_7338,N_7166,N_7092);
xnor U7339 (N_7339,N_6845,N_7060);
and U7340 (N_7340,N_6817,N_6945);
xnor U7341 (N_7341,N_7119,N_6991);
or U7342 (N_7342,N_7152,N_6922);
and U7343 (N_7343,N_6860,N_6856);
xnor U7344 (N_7344,N_7104,N_7048);
xor U7345 (N_7345,N_6941,N_6916);
or U7346 (N_7346,N_7005,N_6977);
nor U7347 (N_7347,N_6936,N_7189);
nand U7348 (N_7348,N_7056,N_7041);
nor U7349 (N_7349,N_6911,N_7132);
nor U7350 (N_7350,N_7118,N_7131);
and U7351 (N_7351,N_6898,N_7037);
and U7352 (N_7352,N_6923,N_7177);
nor U7353 (N_7353,N_6879,N_7122);
or U7354 (N_7354,N_7072,N_6988);
nor U7355 (N_7355,N_6885,N_6962);
or U7356 (N_7356,N_7047,N_6926);
nor U7357 (N_7357,N_6993,N_7130);
nand U7358 (N_7358,N_6974,N_7084);
or U7359 (N_7359,N_7172,N_6842);
nand U7360 (N_7360,N_6953,N_6901);
xnor U7361 (N_7361,N_7141,N_6816);
and U7362 (N_7362,N_7197,N_7040);
and U7363 (N_7363,N_7030,N_6934);
nand U7364 (N_7364,N_6995,N_7015);
and U7365 (N_7365,N_7148,N_6806);
xor U7366 (N_7366,N_7066,N_7112);
and U7367 (N_7367,N_6841,N_7078);
or U7368 (N_7368,N_7187,N_7163);
or U7369 (N_7369,N_6909,N_7025);
nand U7370 (N_7370,N_6907,N_6826);
xnor U7371 (N_7371,N_6818,N_7098);
or U7372 (N_7372,N_6967,N_7023);
xor U7373 (N_7373,N_6912,N_6950);
nand U7374 (N_7374,N_7162,N_7022);
nand U7375 (N_7375,N_7083,N_7142);
xnor U7376 (N_7376,N_6828,N_6938);
nand U7377 (N_7377,N_7094,N_7114);
or U7378 (N_7378,N_7045,N_7183);
nor U7379 (N_7379,N_7144,N_7102);
xor U7380 (N_7380,N_6969,N_7151);
nor U7381 (N_7381,N_6965,N_6932);
xor U7382 (N_7382,N_6809,N_6830);
nor U7383 (N_7383,N_6971,N_6910);
nor U7384 (N_7384,N_7089,N_7101);
or U7385 (N_7385,N_7088,N_6804);
nor U7386 (N_7386,N_7153,N_7167);
or U7387 (N_7387,N_7034,N_6812);
nand U7388 (N_7388,N_6881,N_7146);
xor U7389 (N_7389,N_7186,N_7194);
or U7390 (N_7390,N_6908,N_7042);
nor U7391 (N_7391,N_6875,N_6848);
nand U7392 (N_7392,N_7049,N_6904);
nand U7393 (N_7393,N_6888,N_7038);
nor U7394 (N_7394,N_7175,N_6986);
xor U7395 (N_7395,N_6955,N_6844);
xnor U7396 (N_7396,N_7138,N_7075);
xnor U7397 (N_7397,N_6835,N_6987);
nand U7398 (N_7398,N_6903,N_6952);
nor U7399 (N_7399,N_7105,N_7143);
nand U7400 (N_7400,N_7078,N_6963);
xor U7401 (N_7401,N_6879,N_6811);
nand U7402 (N_7402,N_6962,N_7184);
or U7403 (N_7403,N_6887,N_6924);
nand U7404 (N_7404,N_6902,N_7138);
nand U7405 (N_7405,N_6881,N_7061);
or U7406 (N_7406,N_7027,N_7056);
nand U7407 (N_7407,N_7023,N_6907);
xor U7408 (N_7408,N_7076,N_6864);
or U7409 (N_7409,N_7046,N_6807);
or U7410 (N_7410,N_7023,N_6961);
xor U7411 (N_7411,N_7086,N_6895);
and U7412 (N_7412,N_7018,N_6802);
and U7413 (N_7413,N_7190,N_7124);
xor U7414 (N_7414,N_6880,N_7060);
nor U7415 (N_7415,N_6810,N_6867);
xor U7416 (N_7416,N_7020,N_6916);
nor U7417 (N_7417,N_6932,N_7004);
and U7418 (N_7418,N_6905,N_6998);
and U7419 (N_7419,N_7064,N_7018);
and U7420 (N_7420,N_6959,N_6901);
xor U7421 (N_7421,N_7094,N_7103);
and U7422 (N_7422,N_6900,N_6835);
or U7423 (N_7423,N_7010,N_7183);
and U7424 (N_7424,N_7039,N_6921);
nand U7425 (N_7425,N_7015,N_7136);
nor U7426 (N_7426,N_6901,N_6999);
and U7427 (N_7427,N_7113,N_6931);
xor U7428 (N_7428,N_7085,N_7103);
or U7429 (N_7429,N_7031,N_7167);
and U7430 (N_7430,N_7133,N_7073);
or U7431 (N_7431,N_6970,N_7159);
and U7432 (N_7432,N_6812,N_7137);
and U7433 (N_7433,N_6828,N_6874);
xnor U7434 (N_7434,N_6944,N_6881);
and U7435 (N_7435,N_6992,N_6924);
nand U7436 (N_7436,N_6991,N_7035);
xor U7437 (N_7437,N_7078,N_7033);
xor U7438 (N_7438,N_7044,N_6957);
nor U7439 (N_7439,N_7054,N_7195);
nand U7440 (N_7440,N_6805,N_7182);
xnor U7441 (N_7441,N_7138,N_7035);
or U7442 (N_7442,N_6936,N_7133);
and U7443 (N_7443,N_6939,N_7084);
xnor U7444 (N_7444,N_6940,N_6835);
and U7445 (N_7445,N_7039,N_7122);
xnor U7446 (N_7446,N_7110,N_6950);
nor U7447 (N_7447,N_7002,N_7089);
nand U7448 (N_7448,N_6998,N_6945);
xor U7449 (N_7449,N_7046,N_6988);
or U7450 (N_7450,N_7199,N_7084);
nor U7451 (N_7451,N_6919,N_6936);
nand U7452 (N_7452,N_7018,N_6825);
or U7453 (N_7453,N_6992,N_7094);
xnor U7454 (N_7454,N_7104,N_7178);
or U7455 (N_7455,N_7165,N_7033);
nand U7456 (N_7456,N_7140,N_7145);
nor U7457 (N_7457,N_6837,N_6951);
and U7458 (N_7458,N_6873,N_6807);
nor U7459 (N_7459,N_7144,N_6891);
and U7460 (N_7460,N_6834,N_7068);
nand U7461 (N_7461,N_7140,N_7000);
and U7462 (N_7462,N_6921,N_6811);
or U7463 (N_7463,N_7155,N_6958);
and U7464 (N_7464,N_6877,N_7010);
or U7465 (N_7465,N_7064,N_6923);
or U7466 (N_7466,N_7111,N_7084);
nand U7467 (N_7467,N_6801,N_7095);
nor U7468 (N_7468,N_7103,N_6807);
xor U7469 (N_7469,N_7183,N_6940);
nor U7470 (N_7470,N_7132,N_6882);
nand U7471 (N_7471,N_6911,N_7026);
xnor U7472 (N_7472,N_6827,N_7114);
nor U7473 (N_7473,N_6920,N_6932);
nor U7474 (N_7474,N_6849,N_7086);
and U7475 (N_7475,N_7166,N_7140);
and U7476 (N_7476,N_6909,N_7099);
nor U7477 (N_7477,N_6989,N_6952);
and U7478 (N_7478,N_7153,N_6938);
or U7479 (N_7479,N_7176,N_7157);
nor U7480 (N_7480,N_6979,N_7048);
or U7481 (N_7481,N_6915,N_7001);
nor U7482 (N_7482,N_7022,N_7091);
nor U7483 (N_7483,N_7085,N_6965);
nor U7484 (N_7484,N_7105,N_7137);
xnor U7485 (N_7485,N_6920,N_7033);
xor U7486 (N_7486,N_6966,N_6892);
or U7487 (N_7487,N_6932,N_6977);
xor U7488 (N_7488,N_7047,N_7048);
and U7489 (N_7489,N_6881,N_7011);
nor U7490 (N_7490,N_7024,N_6990);
xor U7491 (N_7491,N_7193,N_6933);
nor U7492 (N_7492,N_7074,N_7123);
xor U7493 (N_7493,N_6804,N_7168);
nand U7494 (N_7494,N_7178,N_6802);
nand U7495 (N_7495,N_6880,N_7184);
or U7496 (N_7496,N_6958,N_6834);
nor U7497 (N_7497,N_6831,N_6855);
nor U7498 (N_7498,N_6988,N_6957);
xor U7499 (N_7499,N_7136,N_6872);
nand U7500 (N_7500,N_7055,N_6856);
nor U7501 (N_7501,N_6827,N_6899);
nand U7502 (N_7502,N_6883,N_6995);
and U7503 (N_7503,N_6825,N_6834);
nand U7504 (N_7504,N_7163,N_7025);
nor U7505 (N_7505,N_7145,N_7137);
nand U7506 (N_7506,N_6954,N_6853);
nand U7507 (N_7507,N_6939,N_7114);
nand U7508 (N_7508,N_6987,N_7032);
or U7509 (N_7509,N_7193,N_7102);
or U7510 (N_7510,N_7109,N_7131);
and U7511 (N_7511,N_6864,N_6976);
xnor U7512 (N_7512,N_7177,N_7091);
nor U7513 (N_7513,N_6913,N_6945);
or U7514 (N_7514,N_7070,N_7080);
nand U7515 (N_7515,N_7060,N_7048);
and U7516 (N_7516,N_7164,N_7163);
nand U7517 (N_7517,N_6969,N_6952);
nand U7518 (N_7518,N_6973,N_6828);
or U7519 (N_7519,N_6988,N_6928);
xnor U7520 (N_7520,N_7074,N_7004);
and U7521 (N_7521,N_6953,N_7137);
xnor U7522 (N_7522,N_6825,N_7146);
nor U7523 (N_7523,N_7003,N_6896);
nor U7524 (N_7524,N_6812,N_7199);
or U7525 (N_7525,N_7073,N_7025);
nor U7526 (N_7526,N_7149,N_7053);
or U7527 (N_7527,N_7063,N_6879);
or U7528 (N_7528,N_6874,N_7132);
nor U7529 (N_7529,N_6890,N_7177);
and U7530 (N_7530,N_6941,N_6898);
xnor U7531 (N_7531,N_6907,N_7157);
and U7532 (N_7532,N_7029,N_7147);
nor U7533 (N_7533,N_6948,N_7142);
and U7534 (N_7534,N_7129,N_6884);
nor U7535 (N_7535,N_7130,N_7080);
xnor U7536 (N_7536,N_7081,N_7043);
nand U7537 (N_7537,N_7166,N_7057);
or U7538 (N_7538,N_7015,N_6873);
nand U7539 (N_7539,N_6942,N_6995);
and U7540 (N_7540,N_7038,N_6833);
nor U7541 (N_7541,N_6893,N_6915);
nor U7542 (N_7542,N_6800,N_6964);
and U7543 (N_7543,N_7023,N_7113);
and U7544 (N_7544,N_6977,N_6802);
nor U7545 (N_7545,N_7070,N_7158);
nand U7546 (N_7546,N_7058,N_7165);
nor U7547 (N_7547,N_6976,N_7055);
xnor U7548 (N_7548,N_7056,N_7128);
nor U7549 (N_7549,N_7002,N_6967);
nand U7550 (N_7550,N_7026,N_6897);
or U7551 (N_7551,N_6979,N_6829);
nand U7552 (N_7552,N_7020,N_6978);
xnor U7553 (N_7553,N_6987,N_6996);
nand U7554 (N_7554,N_6924,N_6902);
nand U7555 (N_7555,N_6872,N_7117);
or U7556 (N_7556,N_6916,N_6963);
nor U7557 (N_7557,N_7111,N_7036);
nor U7558 (N_7558,N_6928,N_6804);
xnor U7559 (N_7559,N_6802,N_7148);
and U7560 (N_7560,N_7163,N_6988);
xor U7561 (N_7561,N_7006,N_7121);
and U7562 (N_7562,N_6926,N_7053);
nand U7563 (N_7563,N_6868,N_7146);
nor U7564 (N_7564,N_6959,N_7076);
xor U7565 (N_7565,N_7109,N_7119);
nand U7566 (N_7566,N_7176,N_7174);
nand U7567 (N_7567,N_6808,N_6843);
and U7568 (N_7568,N_6874,N_7082);
nor U7569 (N_7569,N_7123,N_7039);
nand U7570 (N_7570,N_6910,N_6995);
or U7571 (N_7571,N_7179,N_6849);
or U7572 (N_7572,N_6817,N_7042);
or U7573 (N_7573,N_6812,N_6927);
xor U7574 (N_7574,N_7103,N_6935);
xor U7575 (N_7575,N_6900,N_7175);
nor U7576 (N_7576,N_6842,N_6957);
nor U7577 (N_7577,N_7021,N_7011);
xnor U7578 (N_7578,N_6920,N_7188);
nand U7579 (N_7579,N_7023,N_7136);
or U7580 (N_7580,N_6957,N_6835);
xnor U7581 (N_7581,N_7110,N_7162);
and U7582 (N_7582,N_7177,N_6806);
or U7583 (N_7583,N_6957,N_7018);
nor U7584 (N_7584,N_6944,N_7082);
xnor U7585 (N_7585,N_7149,N_6874);
or U7586 (N_7586,N_7074,N_6993);
or U7587 (N_7587,N_6934,N_7166);
xnor U7588 (N_7588,N_7086,N_7185);
or U7589 (N_7589,N_7041,N_7194);
nor U7590 (N_7590,N_7020,N_6974);
nand U7591 (N_7591,N_7077,N_7142);
or U7592 (N_7592,N_7130,N_6930);
nand U7593 (N_7593,N_7138,N_7165);
xnor U7594 (N_7594,N_7094,N_7151);
nor U7595 (N_7595,N_7021,N_6882);
and U7596 (N_7596,N_7008,N_6819);
nor U7597 (N_7597,N_6980,N_7071);
xnor U7598 (N_7598,N_6980,N_7139);
or U7599 (N_7599,N_6811,N_7161);
and U7600 (N_7600,N_7380,N_7551);
or U7601 (N_7601,N_7245,N_7446);
xnor U7602 (N_7602,N_7499,N_7349);
nor U7603 (N_7603,N_7597,N_7405);
nor U7604 (N_7604,N_7215,N_7583);
xor U7605 (N_7605,N_7352,N_7284);
or U7606 (N_7606,N_7233,N_7267);
and U7607 (N_7607,N_7547,N_7275);
nor U7608 (N_7608,N_7502,N_7249);
xor U7609 (N_7609,N_7252,N_7508);
or U7610 (N_7610,N_7419,N_7390);
nor U7611 (N_7611,N_7479,N_7332);
and U7612 (N_7612,N_7598,N_7202);
xnor U7613 (N_7613,N_7384,N_7437);
nor U7614 (N_7614,N_7457,N_7507);
xor U7615 (N_7615,N_7316,N_7262);
xor U7616 (N_7616,N_7595,N_7473);
xnor U7617 (N_7617,N_7451,N_7448);
or U7618 (N_7618,N_7381,N_7206);
nand U7619 (N_7619,N_7219,N_7357);
nor U7620 (N_7620,N_7310,N_7331);
and U7621 (N_7621,N_7368,N_7234);
nand U7622 (N_7622,N_7476,N_7366);
or U7623 (N_7623,N_7226,N_7225);
and U7624 (N_7624,N_7420,N_7238);
nand U7625 (N_7625,N_7548,N_7318);
nor U7626 (N_7626,N_7577,N_7305);
xnor U7627 (N_7627,N_7271,N_7328);
and U7628 (N_7628,N_7312,N_7445);
nand U7629 (N_7629,N_7309,N_7397);
nand U7630 (N_7630,N_7415,N_7570);
or U7631 (N_7631,N_7295,N_7425);
nand U7632 (N_7632,N_7486,N_7336);
nor U7633 (N_7633,N_7520,N_7385);
or U7634 (N_7634,N_7562,N_7356);
nand U7635 (N_7635,N_7201,N_7449);
and U7636 (N_7636,N_7535,N_7247);
xor U7637 (N_7637,N_7365,N_7589);
nand U7638 (N_7638,N_7463,N_7335);
nor U7639 (N_7639,N_7418,N_7475);
or U7640 (N_7640,N_7441,N_7421);
xnor U7641 (N_7641,N_7599,N_7574);
nor U7642 (N_7642,N_7416,N_7253);
nand U7643 (N_7643,N_7319,N_7558);
nand U7644 (N_7644,N_7423,N_7593);
nand U7645 (N_7645,N_7491,N_7340);
nand U7646 (N_7646,N_7343,N_7452);
nor U7647 (N_7647,N_7469,N_7263);
and U7648 (N_7648,N_7532,N_7482);
or U7649 (N_7649,N_7321,N_7293);
nand U7650 (N_7650,N_7382,N_7325);
nor U7651 (N_7651,N_7587,N_7314);
xnor U7652 (N_7652,N_7200,N_7408);
nand U7653 (N_7653,N_7460,N_7229);
and U7654 (N_7654,N_7212,N_7265);
nand U7655 (N_7655,N_7334,N_7303);
or U7656 (N_7656,N_7531,N_7232);
xor U7657 (N_7657,N_7487,N_7203);
or U7658 (N_7658,N_7484,N_7306);
nand U7659 (N_7659,N_7403,N_7584);
xnor U7660 (N_7660,N_7243,N_7566);
nand U7661 (N_7661,N_7269,N_7470);
and U7662 (N_7662,N_7259,N_7376);
nand U7663 (N_7663,N_7355,N_7521);
or U7664 (N_7664,N_7542,N_7485);
and U7665 (N_7665,N_7501,N_7431);
and U7666 (N_7666,N_7354,N_7468);
xor U7667 (N_7667,N_7594,N_7515);
nand U7668 (N_7668,N_7523,N_7281);
xnor U7669 (N_7669,N_7285,N_7237);
nand U7670 (N_7670,N_7579,N_7311);
nand U7671 (N_7671,N_7456,N_7218);
or U7672 (N_7672,N_7315,N_7545);
nor U7673 (N_7673,N_7533,N_7294);
or U7674 (N_7674,N_7276,N_7373);
and U7675 (N_7675,N_7224,N_7563);
or U7676 (N_7676,N_7537,N_7514);
xor U7677 (N_7677,N_7436,N_7369);
or U7678 (N_7678,N_7304,N_7287);
nand U7679 (N_7679,N_7258,N_7555);
and U7680 (N_7680,N_7517,N_7346);
and U7681 (N_7681,N_7400,N_7498);
nand U7682 (N_7682,N_7454,N_7512);
xnor U7683 (N_7683,N_7550,N_7227);
nor U7684 (N_7684,N_7344,N_7274);
nand U7685 (N_7685,N_7573,N_7527);
or U7686 (N_7686,N_7513,N_7273);
nor U7687 (N_7687,N_7526,N_7544);
or U7688 (N_7688,N_7244,N_7364);
and U7689 (N_7689,N_7474,N_7270);
or U7690 (N_7690,N_7239,N_7223);
nand U7691 (N_7691,N_7472,N_7511);
or U7692 (N_7692,N_7552,N_7255);
or U7693 (N_7693,N_7278,N_7289);
and U7694 (N_7694,N_7268,N_7353);
nand U7695 (N_7695,N_7298,N_7455);
nand U7696 (N_7696,N_7447,N_7337);
nand U7697 (N_7697,N_7481,N_7444);
xor U7698 (N_7698,N_7500,N_7586);
xnor U7699 (N_7699,N_7327,N_7489);
and U7700 (N_7700,N_7559,N_7488);
xor U7701 (N_7701,N_7401,N_7288);
nand U7702 (N_7702,N_7308,N_7264);
xnor U7703 (N_7703,N_7497,N_7326);
and U7704 (N_7704,N_7464,N_7291);
or U7705 (N_7705,N_7217,N_7588);
nor U7706 (N_7706,N_7280,N_7414);
nor U7707 (N_7707,N_7338,N_7393);
or U7708 (N_7708,N_7266,N_7462);
nor U7709 (N_7709,N_7525,N_7216);
or U7710 (N_7710,N_7543,N_7211);
nand U7711 (N_7711,N_7467,N_7461);
and U7712 (N_7712,N_7493,N_7496);
xnor U7713 (N_7713,N_7568,N_7323);
nor U7714 (N_7714,N_7471,N_7580);
nor U7715 (N_7715,N_7534,N_7221);
nor U7716 (N_7716,N_7509,N_7541);
xnor U7717 (N_7717,N_7490,N_7510);
xnor U7718 (N_7718,N_7596,N_7313);
or U7719 (N_7719,N_7299,N_7363);
and U7720 (N_7720,N_7554,N_7411);
xnor U7721 (N_7721,N_7504,N_7450);
or U7722 (N_7722,N_7297,N_7427);
and U7723 (N_7723,N_7240,N_7248);
and U7724 (N_7724,N_7495,N_7214);
nor U7725 (N_7725,N_7430,N_7567);
or U7726 (N_7726,N_7370,N_7459);
nand U7727 (N_7727,N_7296,N_7389);
and U7728 (N_7728,N_7359,N_7205);
nor U7729 (N_7729,N_7553,N_7417);
nor U7730 (N_7730,N_7372,N_7342);
or U7731 (N_7731,N_7506,N_7591);
and U7732 (N_7732,N_7522,N_7569);
xor U7733 (N_7733,N_7560,N_7518);
nor U7734 (N_7734,N_7379,N_7329);
xor U7735 (N_7735,N_7348,N_7465);
and U7736 (N_7736,N_7432,N_7286);
nand U7737 (N_7737,N_7375,N_7387);
or U7738 (N_7738,N_7367,N_7442);
nor U7739 (N_7739,N_7426,N_7261);
and U7740 (N_7740,N_7402,N_7483);
nor U7741 (N_7741,N_7571,N_7204);
nor U7742 (N_7742,N_7235,N_7561);
nand U7743 (N_7743,N_7433,N_7422);
or U7744 (N_7744,N_7307,N_7578);
or U7745 (N_7745,N_7404,N_7440);
and U7746 (N_7746,N_7590,N_7396);
xnor U7747 (N_7747,N_7524,N_7413);
or U7748 (N_7748,N_7351,N_7333);
xor U7749 (N_7749,N_7505,N_7207);
nor U7750 (N_7750,N_7539,N_7383);
and U7751 (N_7751,N_7208,N_7477);
xnor U7752 (N_7752,N_7209,N_7302);
nand U7753 (N_7753,N_7242,N_7429);
and U7754 (N_7754,N_7536,N_7581);
nor U7755 (N_7755,N_7516,N_7210);
nor U7756 (N_7756,N_7478,N_7546);
nand U7757 (N_7757,N_7453,N_7439);
and U7758 (N_7758,N_7222,N_7582);
nor U7759 (N_7759,N_7435,N_7528);
nor U7760 (N_7760,N_7256,N_7374);
nand U7761 (N_7761,N_7330,N_7395);
or U7762 (N_7762,N_7236,N_7360);
nor U7763 (N_7763,N_7228,N_7350);
or U7764 (N_7764,N_7251,N_7361);
nor U7765 (N_7765,N_7407,N_7377);
nor U7766 (N_7766,N_7576,N_7378);
and U7767 (N_7767,N_7388,N_7260);
nor U7768 (N_7768,N_7530,N_7592);
or U7769 (N_7769,N_7339,N_7322);
xor U7770 (N_7770,N_7434,N_7503);
xor U7771 (N_7771,N_7443,N_7399);
or U7772 (N_7772,N_7386,N_7540);
or U7773 (N_7773,N_7277,N_7572);
nand U7774 (N_7774,N_7272,N_7231);
or U7775 (N_7775,N_7292,N_7341);
nand U7776 (N_7776,N_7347,N_7250);
and U7777 (N_7777,N_7279,N_7317);
or U7778 (N_7778,N_7362,N_7492);
nand U7779 (N_7779,N_7257,N_7428);
nor U7780 (N_7780,N_7345,N_7282);
and U7781 (N_7781,N_7358,N_7424);
or U7782 (N_7782,N_7254,N_7529);
nand U7783 (N_7783,N_7301,N_7290);
nor U7784 (N_7784,N_7466,N_7230);
xor U7785 (N_7785,N_7300,N_7557);
xor U7786 (N_7786,N_7519,N_7220);
or U7787 (N_7787,N_7213,N_7458);
nand U7788 (N_7788,N_7410,N_7575);
or U7789 (N_7789,N_7480,N_7438);
nand U7790 (N_7790,N_7565,N_7324);
and U7791 (N_7791,N_7371,N_7585);
or U7792 (N_7792,N_7398,N_7392);
and U7793 (N_7793,N_7564,N_7394);
or U7794 (N_7794,N_7494,N_7549);
or U7795 (N_7795,N_7241,N_7406);
nor U7796 (N_7796,N_7320,N_7556);
or U7797 (N_7797,N_7412,N_7538);
xnor U7798 (N_7798,N_7283,N_7391);
xor U7799 (N_7799,N_7246,N_7409);
or U7800 (N_7800,N_7322,N_7381);
or U7801 (N_7801,N_7314,N_7237);
nand U7802 (N_7802,N_7379,N_7598);
xor U7803 (N_7803,N_7499,N_7567);
xor U7804 (N_7804,N_7596,N_7556);
and U7805 (N_7805,N_7560,N_7349);
nand U7806 (N_7806,N_7211,N_7296);
nand U7807 (N_7807,N_7554,N_7319);
nand U7808 (N_7808,N_7345,N_7578);
and U7809 (N_7809,N_7451,N_7316);
and U7810 (N_7810,N_7458,N_7566);
nand U7811 (N_7811,N_7333,N_7577);
nor U7812 (N_7812,N_7561,N_7557);
or U7813 (N_7813,N_7453,N_7205);
xnor U7814 (N_7814,N_7377,N_7334);
nor U7815 (N_7815,N_7326,N_7350);
nor U7816 (N_7816,N_7512,N_7568);
and U7817 (N_7817,N_7489,N_7460);
nor U7818 (N_7818,N_7453,N_7235);
and U7819 (N_7819,N_7533,N_7321);
nor U7820 (N_7820,N_7298,N_7511);
or U7821 (N_7821,N_7500,N_7598);
nor U7822 (N_7822,N_7507,N_7404);
and U7823 (N_7823,N_7234,N_7395);
or U7824 (N_7824,N_7472,N_7257);
nand U7825 (N_7825,N_7552,N_7318);
nand U7826 (N_7826,N_7434,N_7579);
nor U7827 (N_7827,N_7531,N_7583);
nor U7828 (N_7828,N_7207,N_7538);
xor U7829 (N_7829,N_7430,N_7324);
xor U7830 (N_7830,N_7558,N_7226);
nor U7831 (N_7831,N_7206,N_7288);
and U7832 (N_7832,N_7297,N_7502);
and U7833 (N_7833,N_7203,N_7336);
or U7834 (N_7834,N_7396,N_7516);
nand U7835 (N_7835,N_7330,N_7414);
and U7836 (N_7836,N_7404,N_7542);
or U7837 (N_7837,N_7240,N_7430);
nand U7838 (N_7838,N_7453,N_7278);
nand U7839 (N_7839,N_7329,N_7263);
xnor U7840 (N_7840,N_7334,N_7285);
xor U7841 (N_7841,N_7471,N_7313);
nor U7842 (N_7842,N_7297,N_7597);
or U7843 (N_7843,N_7381,N_7432);
or U7844 (N_7844,N_7221,N_7357);
nor U7845 (N_7845,N_7535,N_7484);
xnor U7846 (N_7846,N_7385,N_7222);
xnor U7847 (N_7847,N_7540,N_7471);
or U7848 (N_7848,N_7438,N_7426);
xor U7849 (N_7849,N_7565,N_7295);
nor U7850 (N_7850,N_7291,N_7409);
xor U7851 (N_7851,N_7487,N_7561);
nand U7852 (N_7852,N_7308,N_7590);
or U7853 (N_7853,N_7522,N_7287);
xnor U7854 (N_7854,N_7348,N_7529);
or U7855 (N_7855,N_7280,N_7271);
xor U7856 (N_7856,N_7245,N_7454);
xnor U7857 (N_7857,N_7494,N_7294);
nand U7858 (N_7858,N_7511,N_7313);
or U7859 (N_7859,N_7397,N_7571);
nor U7860 (N_7860,N_7218,N_7254);
or U7861 (N_7861,N_7570,N_7382);
nand U7862 (N_7862,N_7403,N_7393);
or U7863 (N_7863,N_7337,N_7227);
and U7864 (N_7864,N_7499,N_7451);
nand U7865 (N_7865,N_7319,N_7330);
nor U7866 (N_7866,N_7581,N_7554);
nand U7867 (N_7867,N_7504,N_7512);
xnor U7868 (N_7868,N_7589,N_7489);
xnor U7869 (N_7869,N_7352,N_7230);
xor U7870 (N_7870,N_7420,N_7243);
nand U7871 (N_7871,N_7232,N_7415);
or U7872 (N_7872,N_7398,N_7530);
nor U7873 (N_7873,N_7304,N_7503);
and U7874 (N_7874,N_7361,N_7464);
nand U7875 (N_7875,N_7429,N_7527);
nor U7876 (N_7876,N_7574,N_7326);
nand U7877 (N_7877,N_7228,N_7524);
nor U7878 (N_7878,N_7307,N_7444);
xor U7879 (N_7879,N_7487,N_7264);
or U7880 (N_7880,N_7455,N_7363);
and U7881 (N_7881,N_7335,N_7408);
xor U7882 (N_7882,N_7543,N_7437);
nand U7883 (N_7883,N_7351,N_7225);
nand U7884 (N_7884,N_7514,N_7375);
and U7885 (N_7885,N_7226,N_7327);
xor U7886 (N_7886,N_7528,N_7395);
xor U7887 (N_7887,N_7253,N_7336);
or U7888 (N_7888,N_7220,N_7372);
or U7889 (N_7889,N_7352,N_7317);
xnor U7890 (N_7890,N_7493,N_7456);
nor U7891 (N_7891,N_7546,N_7458);
and U7892 (N_7892,N_7284,N_7354);
nand U7893 (N_7893,N_7486,N_7362);
or U7894 (N_7894,N_7465,N_7599);
xor U7895 (N_7895,N_7437,N_7395);
or U7896 (N_7896,N_7213,N_7294);
or U7897 (N_7897,N_7571,N_7245);
nor U7898 (N_7898,N_7253,N_7559);
or U7899 (N_7899,N_7353,N_7207);
or U7900 (N_7900,N_7585,N_7271);
or U7901 (N_7901,N_7230,N_7414);
xor U7902 (N_7902,N_7564,N_7309);
and U7903 (N_7903,N_7494,N_7550);
nor U7904 (N_7904,N_7497,N_7594);
and U7905 (N_7905,N_7399,N_7336);
and U7906 (N_7906,N_7249,N_7582);
nor U7907 (N_7907,N_7520,N_7475);
or U7908 (N_7908,N_7353,N_7564);
or U7909 (N_7909,N_7526,N_7390);
and U7910 (N_7910,N_7467,N_7357);
xor U7911 (N_7911,N_7591,N_7437);
or U7912 (N_7912,N_7266,N_7235);
and U7913 (N_7913,N_7458,N_7241);
or U7914 (N_7914,N_7362,N_7503);
nor U7915 (N_7915,N_7380,N_7455);
or U7916 (N_7916,N_7375,N_7398);
nand U7917 (N_7917,N_7459,N_7554);
xnor U7918 (N_7918,N_7528,N_7231);
and U7919 (N_7919,N_7416,N_7247);
or U7920 (N_7920,N_7412,N_7257);
nor U7921 (N_7921,N_7502,N_7355);
and U7922 (N_7922,N_7264,N_7412);
nor U7923 (N_7923,N_7408,N_7225);
and U7924 (N_7924,N_7273,N_7584);
nor U7925 (N_7925,N_7570,N_7214);
nor U7926 (N_7926,N_7276,N_7227);
xor U7927 (N_7927,N_7225,N_7336);
or U7928 (N_7928,N_7495,N_7371);
nor U7929 (N_7929,N_7413,N_7218);
and U7930 (N_7930,N_7248,N_7418);
nor U7931 (N_7931,N_7487,N_7298);
or U7932 (N_7932,N_7485,N_7556);
nor U7933 (N_7933,N_7267,N_7414);
and U7934 (N_7934,N_7208,N_7353);
and U7935 (N_7935,N_7440,N_7214);
and U7936 (N_7936,N_7522,N_7236);
nor U7937 (N_7937,N_7548,N_7343);
xor U7938 (N_7938,N_7310,N_7225);
nand U7939 (N_7939,N_7521,N_7347);
xnor U7940 (N_7940,N_7530,N_7568);
nor U7941 (N_7941,N_7253,N_7573);
nand U7942 (N_7942,N_7561,N_7343);
xor U7943 (N_7943,N_7587,N_7225);
nor U7944 (N_7944,N_7442,N_7421);
nor U7945 (N_7945,N_7307,N_7249);
nand U7946 (N_7946,N_7511,N_7466);
and U7947 (N_7947,N_7583,N_7233);
nor U7948 (N_7948,N_7536,N_7565);
nor U7949 (N_7949,N_7463,N_7563);
or U7950 (N_7950,N_7360,N_7566);
nand U7951 (N_7951,N_7505,N_7322);
nor U7952 (N_7952,N_7526,N_7580);
or U7953 (N_7953,N_7285,N_7577);
nor U7954 (N_7954,N_7278,N_7207);
or U7955 (N_7955,N_7550,N_7318);
xnor U7956 (N_7956,N_7561,N_7513);
or U7957 (N_7957,N_7453,N_7416);
nor U7958 (N_7958,N_7299,N_7476);
or U7959 (N_7959,N_7515,N_7347);
and U7960 (N_7960,N_7202,N_7222);
xnor U7961 (N_7961,N_7317,N_7518);
nand U7962 (N_7962,N_7512,N_7230);
nand U7963 (N_7963,N_7392,N_7474);
xnor U7964 (N_7964,N_7250,N_7314);
or U7965 (N_7965,N_7467,N_7472);
and U7966 (N_7966,N_7229,N_7241);
and U7967 (N_7967,N_7563,N_7402);
xnor U7968 (N_7968,N_7510,N_7258);
or U7969 (N_7969,N_7204,N_7338);
nand U7970 (N_7970,N_7512,N_7580);
and U7971 (N_7971,N_7501,N_7263);
or U7972 (N_7972,N_7287,N_7242);
nand U7973 (N_7973,N_7425,N_7339);
xor U7974 (N_7974,N_7377,N_7565);
xnor U7975 (N_7975,N_7351,N_7394);
nor U7976 (N_7976,N_7291,N_7381);
nand U7977 (N_7977,N_7231,N_7300);
xor U7978 (N_7978,N_7298,N_7465);
nor U7979 (N_7979,N_7564,N_7231);
xor U7980 (N_7980,N_7471,N_7349);
or U7981 (N_7981,N_7367,N_7350);
nand U7982 (N_7982,N_7439,N_7373);
or U7983 (N_7983,N_7487,N_7263);
and U7984 (N_7984,N_7205,N_7494);
or U7985 (N_7985,N_7220,N_7273);
nor U7986 (N_7986,N_7578,N_7438);
nor U7987 (N_7987,N_7377,N_7532);
and U7988 (N_7988,N_7411,N_7472);
nor U7989 (N_7989,N_7460,N_7342);
and U7990 (N_7990,N_7534,N_7261);
nor U7991 (N_7991,N_7241,N_7282);
and U7992 (N_7992,N_7233,N_7225);
nor U7993 (N_7993,N_7349,N_7541);
or U7994 (N_7994,N_7402,N_7260);
and U7995 (N_7995,N_7519,N_7346);
and U7996 (N_7996,N_7201,N_7462);
and U7997 (N_7997,N_7525,N_7273);
nand U7998 (N_7998,N_7535,N_7362);
or U7999 (N_7999,N_7500,N_7380);
and U8000 (N_8000,N_7676,N_7766);
nand U8001 (N_8001,N_7790,N_7685);
and U8002 (N_8002,N_7610,N_7930);
and U8003 (N_8003,N_7828,N_7735);
and U8004 (N_8004,N_7670,N_7955);
and U8005 (N_8005,N_7633,N_7797);
or U8006 (N_8006,N_7748,N_7872);
nand U8007 (N_8007,N_7689,N_7983);
and U8008 (N_8008,N_7961,N_7687);
nor U8009 (N_8009,N_7860,N_7706);
nand U8010 (N_8010,N_7924,N_7900);
nand U8011 (N_8011,N_7656,N_7700);
xor U8012 (N_8012,N_7720,N_7767);
or U8013 (N_8013,N_7732,N_7614);
xnor U8014 (N_8014,N_7885,N_7972);
nor U8015 (N_8015,N_7840,N_7819);
nand U8016 (N_8016,N_7897,N_7631);
or U8017 (N_8017,N_7753,N_7811);
and U8018 (N_8018,N_7902,N_7803);
nand U8019 (N_8019,N_7665,N_7867);
and U8020 (N_8020,N_7931,N_7745);
xnor U8021 (N_8021,N_7603,N_7796);
and U8022 (N_8022,N_7761,N_7786);
nand U8023 (N_8023,N_7815,N_7939);
xor U8024 (N_8024,N_7878,N_7801);
and U8025 (N_8025,N_7929,N_7742);
xnor U8026 (N_8026,N_7770,N_7870);
nand U8027 (N_8027,N_7859,N_7608);
nor U8028 (N_8028,N_7919,N_7952);
nor U8029 (N_8029,N_7994,N_7727);
or U8030 (N_8030,N_7873,N_7768);
nor U8031 (N_8031,N_7917,N_7731);
nand U8032 (N_8032,N_7818,N_7776);
xor U8033 (N_8033,N_7830,N_7901);
xnor U8034 (N_8034,N_7975,N_7705);
nor U8035 (N_8035,N_7949,N_7852);
or U8036 (N_8036,N_7711,N_7658);
nand U8037 (N_8037,N_7984,N_7707);
and U8038 (N_8038,N_7691,N_7607);
and U8039 (N_8039,N_7978,N_7789);
nor U8040 (N_8040,N_7916,N_7947);
nand U8041 (N_8041,N_7954,N_7673);
xor U8042 (N_8042,N_7773,N_7999);
nand U8043 (N_8043,N_7764,N_7646);
or U8044 (N_8044,N_7765,N_7798);
and U8045 (N_8045,N_7617,N_7960);
xor U8046 (N_8046,N_7654,N_7849);
xnor U8047 (N_8047,N_7688,N_7835);
or U8048 (N_8048,N_7925,N_7667);
and U8049 (N_8049,N_7683,N_7788);
or U8050 (N_8050,N_7616,N_7655);
xnor U8051 (N_8051,N_7934,N_7751);
nor U8052 (N_8052,N_7845,N_7879);
nand U8053 (N_8053,N_7956,N_7805);
xor U8054 (N_8054,N_7958,N_7906);
nor U8055 (N_8055,N_7998,N_7693);
or U8056 (N_8056,N_7836,N_7716);
or U8057 (N_8057,N_7756,N_7923);
or U8058 (N_8058,N_7605,N_7883);
xnor U8059 (N_8059,N_7963,N_7992);
nor U8060 (N_8060,N_7944,N_7965);
xor U8061 (N_8061,N_7825,N_7936);
and U8062 (N_8062,N_7675,N_7663);
nand U8063 (N_8063,N_7813,N_7821);
and U8064 (N_8064,N_7838,N_7785);
nand U8065 (N_8065,N_7857,N_7635);
or U8066 (N_8066,N_7717,N_7697);
nor U8067 (N_8067,N_7793,N_7908);
and U8068 (N_8068,N_7943,N_7772);
or U8069 (N_8069,N_7971,N_7846);
xnor U8070 (N_8070,N_7854,N_7666);
nor U8071 (N_8071,N_7763,N_7953);
xnor U8072 (N_8072,N_7771,N_7973);
or U8073 (N_8073,N_7966,N_7841);
or U8074 (N_8074,N_7853,N_7649);
xnor U8075 (N_8075,N_7913,N_7634);
nor U8076 (N_8076,N_7833,N_7938);
nand U8077 (N_8077,N_7699,N_7904);
nand U8078 (N_8078,N_7777,N_7792);
or U8079 (N_8079,N_7969,N_7782);
or U8080 (N_8080,N_7834,N_7737);
xor U8081 (N_8081,N_7628,N_7613);
xnor U8082 (N_8082,N_7847,N_7632);
or U8083 (N_8083,N_7645,N_7886);
nand U8084 (N_8084,N_7807,N_7875);
or U8085 (N_8085,N_7881,N_7642);
and U8086 (N_8086,N_7743,N_7657);
nand U8087 (N_8087,N_7890,N_7959);
xor U8088 (N_8088,N_7866,N_7621);
or U8089 (N_8089,N_7714,N_7868);
nand U8090 (N_8090,N_7606,N_7730);
nand U8091 (N_8091,N_7639,N_7620);
and U8092 (N_8092,N_7827,N_7750);
or U8093 (N_8093,N_7692,N_7848);
and U8094 (N_8094,N_7874,N_7888);
and U8095 (N_8095,N_7744,N_7704);
xnor U8096 (N_8096,N_7668,N_7967);
nor U8097 (N_8097,N_7957,N_7926);
nor U8098 (N_8098,N_7802,N_7880);
xor U8099 (N_8099,N_7661,N_7829);
and U8100 (N_8100,N_7903,N_7659);
nand U8101 (N_8101,N_7783,N_7701);
nand U8102 (N_8102,N_7647,N_7612);
nand U8103 (N_8103,N_7914,N_7774);
and U8104 (N_8104,N_7889,N_7991);
or U8105 (N_8105,N_7652,N_7780);
and U8106 (N_8106,N_7945,N_7862);
or U8107 (N_8107,N_7600,N_7909);
or U8108 (N_8108,N_7970,N_7746);
nand U8109 (N_8109,N_7951,N_7712);
or U8110 (N_8110,N_7725,N_7723);
xnor U8111 (N_8111,N_7976,N_7740);
nor U8112 (N_8112,N_7648,N_7899);
nand U8113 (N_8113,N_7898,N_7602);
nor U8114 (N_8114,N_7722,N_7993);
nand U8115 (N_8115,N_7625,N_7709);
and U8116 (N_8116,N_7907,N_7912);
nor U8117 (N_8117,N_7988,N_7942);
nor U8118 (N_8118,N_7817,N_7824);
nor U8119 (N_8119,N_7794,N_7877);
nor U8120 (N_8120,N_7618,N_7671);
xor U8121 (N_8121,N_7921,N_7987);
or U8122 (N_8122,N_7703,N_7922);
or U8123 (N_8123,N_7686,N_7747);
and U8124 (N_8124,N_7651,N_7630);
nor U8125 (N_8125,N_7762,N_7749);
and U8126 (N_8126,N_7791,N_7968);
and U8127 (N_8127,N_7678,N_7941);
nand U8128 (N_8128,N_7604,N_7626);
and U8129 (N_8129,N_7719,N_7660);
or U8130 (N_8130,N_7644,N_7728);
nor U8131 (N_8131,N_7698,N_7804);
or U8132 (N_8132,N_7911,N_7869);
xnor U8133 (N_8133,N_7808,N_7726);
or U8134 (N_8134,N_7876,N_7641);
nor U8135 (N_8135,N_7812,N_7609);
nor U8136 (N_8136,N_7729,N_7850);
or U8137 (N_8137,N_7778,N_7640);
xnor U8138 (N_8138,N_7871,N_7674);
xnor U8139 (N_8139,N_7864,N_7769);
xor U8140 (N_8140,N_7855,N_7781);
or U8141 (N_8141,N_7733,N_7893);
and U8142 (N_8142,N_7682,N_7928);
and U8143 (N_8143,N_7891,N_7806);
xnor U8144 (N_8144,N_7964,N_7927);
nand U8145 (N_8145,N_7800,N_7843);
or U8146 (N_8146,N_7933,N_7882);
nor U8147 (N_8147,N_7977,N_7937);
xor U8148 (N_8148,N_7643,N_7662);
nand U8149 (N_8149,N_7851,N_7915);
nand U8150 (N_8150,N_7837,N_7677);
nor U8151 (N_8151,N_7861,N_7996);
nand U8152 (N_8152,N_7680,N_7946);
nand U8153 (N_8153,N_7974,N_7995);
nand U8154 (N_8154,N_7787,N_7816);
nand U8155 (N_8155,N_7831,N_7636);
nor U8156 (N_8156,N_7810,N_7950);
and U8157 (N_8157,N_7601,N_7684);
nand U8158 (N_8158,N_7695,N_7624);
xor U8159 (N_8159,N_7638,N_7962);
nand U8160 (N_8160,N_7611,N_7989);
and U8161 (N_8161,N_7724,N_7759);
nand U8162 (N_8162,N_7814,N_7681);
nor U8163 (N_8163,N_7894,N_7884);
nand U8164 (N_8164,N_7760,N_7905);
nand U8165 (N_8165,N_7948,N_7755);
nor U8166 (N_8166,N_7650,N_7826);
xor U8167 (N_8167,N_7910,N_7754);
nor U8168 (N_8168,N_7887,N_7739);
nor U8169 (N_8169,N_7896,N_7920);
nand U8170 (N_8170,N_7710,N_7997);
xor U8171 (N_8171,N_7981,N_7820);
xor U8172 (N_8172,N_7736,N_7713);
or U8173 (N_8173,N_7795,N_7892);
and U8174 (N_8174,N_7856,N_7822);
nand U8175 (N_8175,N_7932,N_7979);
nor U8176 (N_8176,N_7741,N_7799);
or U8177 (N_8177,N_7694,N_7775);
xnor U8178 (N_8178,N_7986,N_7863);
or U8179 (N_8179,N_7734,N_7637);
xnor U8180 (N_8180,N_7752,N_7779);
and U8181 (N_8181,N_7715,N_7935);
xnor U8182 (N_8182,N_7858,N_7619);
xor U8183 (N_8183,N_7718,N_7844);
xor U8184 (N_8184,N_7895,N_7918);
xnor U8185 (N_8185,N_7980,N_7664);
xor U8186 (N_8186,N_7721,N_7823);
nand U8187 (N_8187,N_7672,N_7622);
nand U8188 (N_8188,N_7623,N_7629);
xnor U8189 (N_8189,N_7738,N_7627);
and U8190 (N_8190,N_7708,N_7990);
nor U8191 (N_8191,N_7839,N_7809);
nand U8192 (N_8192,N_7758,N_7784);
nor U8193 (N_8193,N_7832,N_7757);
and U8194 (N_8194,N_7696,N_7669);
nand U8195 (N_8195,N_7690,N_7615);
xnor U8196 (N_8196,N_7940,N_7842);
nor U8197 (N_8197,N_7865,N_7679);
nand U8198 (N_8198,N_7985,N_7982);
or U8199 (N_8199,N_7702,N_7653);
and U8200 (N_8200,N_7985,N_7919);
nor U8201 (N_8201,N_7972,N_7975);
xnor U8202 (N_8202,N_7605,N_7668);
or U8203 (N_8203,N_7743,N_7661);
and U8204 (N_8204,N_7979,N_7836);
and U8205 (N_8205,N_7604,N_7730);
nor U8206 (N_8206,N_7635,N_7983);
nor U8207 (N_8207,N_7865,N_7757);
nand U8208 (N_8208,N_7957,N_7748);
and U8209 (N_8209,N_7998,N_7904);
or U8210 (N_8210,N_7790,N_7832);
or U8211 (N_8211,N_7895,N_7625);
nand U8212 (N_8212,N_7933,N_7828);
or U8213 (N_8213,N_7616,N_7722);
or U8214 (N_8214,N_7862,N_7834);
xnor U8215 (N_8215,N_7700,N_7600);
and U8216 (N_8216,N_7940,N_7708);
and U8217 (N_8217,N_7709,N_7881);
or U8218 (N_8218,N_7615,N_7952);
nand U8219 (N_8219,N_7899,N_7952);
nand U8220 (N_8220,N_7622,N_7707);
or U8221 (N_8221,N_7816,N_7633);
nand U8222 (N_8222,N_7810,N_7927);
nor U8223 (N_8223,N_7871,N_7916);
nor U8224 (N_8224,N_7817,N_7983);
and U8225 (N_8225,N_7888,N_7762);
nand U8226 (N_8226,N_7750,N_7969);
nor U8227 (N_8227,N_7843,N_7789);
nand U8228 (N_8228,N_7928,N_7825);
or U8229 (N_8229,N_7837,N_7922);
nor U8230 (N_8230,N_7994,N_7785);
and U8231 (N_8231,N_7615,N_7798);
xnor U8232 (N_8232,N_7724,N_7960);
and U8233 (N_8233,N_7936,N_7711);
or U8234 (N_8234,N_7753,N_7747);
nand U8235 (N_8235,N_7845,N_7776);
and U8236 (N_8236,N_7866,N_7943);
nand U8237 (N_8237,N_7624,N_7858);
or U8238 (N_8238,N_7829,N_7773);
or U8239 (N_8239,N_7705,N_7618);
or U8240 (N_8240,N_7768,N_7898);
and U8241 (N_8241,N_7844,N_7796);
nand U8242 (N_8242,N_7907,N_7680);
nand U8243 (N_8243,N_7793,N_7827);
and U8244 (N_8244,N_7958,N_7827);
or U8245 (N_8245,N_7747,N_7667);
nand U8246 (N_8246,N_7629,N_7865);
nor U8247 (N_8247,N_7830,N_7809);
xor U8248 (N_8248,N_7604,N_7813);
nand U8249 (N_8249,N_7701,N_7997);
nor U8250 (N_8250,N_7632,N_7794);
and U8251 (N_8251,N_7757,N_7732);
xnor U8252 (N_8252,N_7990,N_7865);
and U8253 (N_8253,N_7941,N_7927);
and U8254 (N_8254,N_7828,N_7920);
nor U8255 (N_8255,N_7978,N_7889);
nand U8256 (N_8256,N_7930,N_7941);
nand U8257 (N_8257,N_7792,N_7786);
nand U8258 (N_8258,N_7668,N_7736);
nand U8259 (N_8259,N_7704,N_7721);
or U8260 (N_8260,N_7894,N_7899);
xnor U8261 (N_8261,N_7850,N_7773);
nand U8262 (N_8262,N_7961,N_7989);
xor U8263 (N_8263,N_7716,N_7745);
xor U8264 (N_8264,N_7726,N_7772);
or U8265 (N_8265,N_7972,N_7847);
xor U8266 (N_8266,N_7957,N_7734);
nor U8267 (N_8267,N_7842,N_7880);
nand U8268 (N_8268,N_7925,N_7875);
nand U8269 (N_8269,N_7820,N_7997);
xor U8270 (N_8270,N_7692,N_7735);
nor U8271 (N_8271,N_7848,N_7905);
xnor U8272 (N_8272,N_7878,N_7769);
nor U8273 (N_8273,N_7908,N_7829);
nand U8274 (N_8274,N_7654,N_7848);
or U8275 (N_8275,N_7941,N_7898);
nor U8276 (N_8276,N_7721,N_7647);
nor U8277 (N_8277,N_7880,N_7613);
nor U8278 (N_8278,N_7921,N_7676);
or U8279 (N_8279,N_7610,N_7956);
and U8280 (N_8280,N_7762,N_7981);
nor U8281 (N_8281,N_7832,N_7700);
nand U8282 (N_8282,N_7652,N_7870);
and U8283 (N_8283,N_7851,N_7991);
nor U8284 (N_8284,N_7934,N_7707);
and U8285 (N_8285,N_7900,N_7684);
or U8286 (N_8286,N_7769,N_7737);
nor U8287 (N_8287,N_7951,N_7636);
or U8288 (N_8288,N_7821,N_7755);
and U8289 (N_8289,N_7666,N_7768);
xnor U8290 (N_8290,N_7741,N_7996);
xnor U8291 (N_8291,N_7987,N_7802);
nor U8292 (N_8292,N_7831,N_7803);
and U8293 (N_8293,N_7947,N_7982);
xnor U8294 (N_8294,N_7853,N_7627);
and U8295 (N_8295,N_7618,N_7870);
xor U8296 (N_8296,N_7800,N_7639);
xor U8297 (N_8297,N_7838,N_7752);
nand U8298 (N_8298,N_7783,N_7672);
or U8299 (N_8299,N_7851,N_7602);
xnor U8300 (N_8300,N_7979,N_7769);
and U8301 (N_8301,N_7602,N_7670);
nor U8302 (N_8302,N_7865,N_7870);
and U8303 (N_8303,N_7657,N_7883);
or U8304 (N_8304,N_7875,N_7750);
xor U8305 (N_8305,N_7678,N_7923);
and U8306 (N_8306,N_7962,N_7841);
nand U8307 (N_8307,N_7909,N_7860);
nand U8308 (N_8308,N_7843,N_7744);
or U8309 (N_8309,N_7796,N_7877);
nand U8310 (N_8310,N_7628,N_7974);
and U8311 (N_8311,N_7631,N_7961);
nand U8312 (N_8312,N_7881,N_7685);
xor U8313 (N_8313,N_7720,N_7764);
nor U8314 (N_8314,N_7728,N_7782);
or U8315 (N_8315,N_7981,N_7906);
xnor U8316 (N_8316,N_7603,N_7727);
nand U8317 (N_8317,N_7959,N_7723);
or U8318 (N_8318,N_7665,N_7764);
nand U8319 (N_8319,N_7961,N_7723);
nor U8320 (N_8320,N_7797,N_7788);
nor U8321 (N_8321,N_7998,N_7736);
or U8322 (N_8322,N_7637,N_7607);
or U8323 (N_8323,N_7755,N_7998);
xnor U8324 (N_8324,N_7628,N_7715);
and U8325 (N_8325,N_7830,N_7639);
and U8326 (N_8326,N_7612,N_7799);
nand U8327 (N_8327,N_7681,N_7680);
or U8328 (N_8328,N_7918,N_7825);
nor U8329 (N_8329,N_7881,N_7684);
and U8330 (N_8330,N_7968,N_7944);
and U8331 (N_8331,N_7719,N_7680);
nand U8332 (N_8332,N_7680,N_7899);
and U8333 (N_8333,N_7890,N_7770);
xor U8334 (N_8334,N_7798,N_7659);
and U8335 (N_8335,N_7880,N_7717);
and U8336 (N_8336,N_7898,N_7681);
xnor U8337 (N_8337,N_7941,N_7650);
and U8338 (N_8338,N_7665,N_7866);
or U8339 (N_8339,N_7917,N_7876);
nand U8340 (N_8340,N_7610,N_7724);
nand U8341 (N_8341,N_7789,N_7661);
or U8342 (N_8342,N_7912,N_7816);
or U8343 (N_8343,N_7897,N_7642);
or U8344 (N_8344,N_7618,N_7977);
and U8345 (N_8345,N_7822,N_7980);
nand U8346 (N_8346,N_7926,N_7911);
nand U8347 (N_8347,N_7735,N_7982);
nand U8348 (N_8348,N_7792,N_7816);
xor U8349 (N_8349,N_7705,N_7672);
xor U8350 (N_8350,N_7642,N_7973);
xnor U8351 (N_8351,N_7646,N_7634);
and U8352 (N_8352,N_7612,N_7908);
nor U8353 (N_8353,N_7943,N_7792);
nand U8354 (N_8354,N_7914,N_7959);
and U8355 (N_8355,N_7915,N_7777);
or U8356 (N_8356,N_7624,N_7937);
nand U8357 (N_8357,N_7764,N_7975);
and U8358 (N_8358,N_7691,N_7785);
or U8359 (N_8359,N_7610,N_7794);
nor U8360 (N_8360,N_7795,N_7989);
nand U8361 (N_8361,N_7737,N_7867);
and U8362 (N_8362,N_7699,N_7934);
nor U8363 (N_8363,N_7695,N_7629);
and U8364 (N_8364,N_7625,N_7921);
nor U8365 (N_8365,N_7680,N_7872);
nor U8366 (N_8366,N_7939,N_7837);
and U8367 (N_8367,N_7966,N_7905);
nor U8368 (N_8368,N_7665,N_7674);
nor U8369 (N_8369,N_7841,N_7637);
nor U8370 (N_8370,N_7618,N_7900);
nand U8371 (N_8371,N_7819,N_7914);
and U8372 (N_8372,N_7766,N_7753);
or U8373 (N_8373,N_7650,N_7736);
or U8374 (N_8374,N_7636,N_7858);
and U8375 (N_8375,N_7831,N_7914);
nand U8376 (N_8376,N_7887,N_7696);
and U8377 (N_8377,N_7779,N_7729);
or U8378 (N_8378,N_7765,N_7927);
or U8379 (N_8379,N_7882,N_7820);
or U8380 (N_8380,N_7907,N_7944);
and U8381 (N_8381,N_7854,N_7992);
nor U8382 (N_8382,N_7767,N_7778);
nor U8383 (N_8383,N_7600,N_7810);
or U8384 (N_8384,N_7735,N_7906);
nor U8385 (N_8385,N_7990,N_7779);
and U8386 (N_8386,N_7876,N_7873);
nor U8387 (N_8387,N_7694,N_7953);
nor U8388 (N_8388,N_7791,N_7751);
and U8389 (N_8389,N_7906,N_7663);
nand U8390 (N_8390,N_7938,N_7718);
nor U8391 (N_8391,N_7774,N_7842);
or U8392 (N_8392,N_7611,N_7912);
nor U8393 (N_8393,N_7750,N_7882);
nand U8394 (N_8394,N_7741,N_7780);
and U8395 (N_8395,N_7974,N_7757);
or U8396 (N_8396,N_7815,N_7824);
xor U8397 (N_8397,N_7693,N_7735);
xnor U8398 (N_8398,N_7635,N_7862);
nor U8399 (N_8399,N_7974,N_7703);
xor U8400 (N_8400,N_8170,N_8296);
and U8401 (N_8401,N_8267,N_8057);
and U8402 (N_8402,N_8372,N_8060);
nor U8403 (N_8403,N_8245,N_8302);
nor U8404 (N_8404,N_8384,N_8225);
or U8405 (N_8405,N_8256,N_8163);
or U8406 (N_8406,N_8089,N_8120);
nand U8407 (N_8407,N_8326,N_8152);
xnor U8408 (N_8408,N_8050,N_8025);
nor U8409 (N_8409,N_8146,N_8123);
nor U8410 (N_8410,N_8046,N_8385);
and U8411 (N_8411,N_8353,N_8012);
or U8412 (N_8412,N_8017,N_8303);
nor U8413 (N_8413,N_8139,N_8233);
nor U8414 (N_8414,N_8086,N_8249);
and U8415 (N_8415,N_8186,N_8076);
and U8416 (N_8416,N_8305,N_8125);
nand U8417 (N_8417,N_8237,N_8119);
xor U8418 (N_8418,N_8390,N_8301);
and U8419 (N_8419,N_8315,N_8395);
nor U8420 (N_8420,N_8009,N_8295);
and U8421 (N_8421,N_8355,N_8199);
xor U8422 (N_8422,N_8065,N_8091);
or U8423 (N_8423,N_8298,N_8087);
nand U8424 (N_8424,N_8354,N_8068);
nand U8425 (N_8425,N_8138,N_8192);
or U8426 (N_8426,N_8160,N_8378);
and U8427 (N_8427,N_8329,N_8097);
xor U8428 (N_8428,N_8211,N_8083);
and U8429 (N_8429,N_8345,N_8039);
nor U8430 (N_8430,N_8197,N_8351);
and U8431 (N_8431,N_8389,N_8277);
nand U8432 (N_8432,N_8208,N_8055);
nand U8433 (N_8433,N_8288,N_8201);
or U8434 (N_8434,N_8275,N_8387);
xnor U8435 (N_8435,N_8085,N_8168);
or U8436 (N_8436,N_8118,N_8052);
nor U8437 (N_8437,N_8343,N_8191);
nand U8438 (N_8438,N_8193,N_8321);
nor U8439 (N_8439,N_8010,N_8143);
and U8440 (N_8440,N_8058,N_8096);
and U8441 (N_8441,N_8350,N_8364);
and U8442 (N_8442,N_8289,N_8374);
or U8443 (N_8443,N_8113,N_8394);
or U8444 (N_8444,N_8373,N_8126);
nand U8445 (N_8445,N_8397,N_8136);
and U8446 (N_8446,N_8260,N_8024);
nor U8447 (N_8447,N_8176,N_8279);
and U8448 (N_8448,N_8034,N_8051);
or U8449 (N_8449,N_8259,N_8239);
nor U8450 (N_8450,N_8070,N_8377);
xor U8451 (N_8451,N_8347,N_8011);
nor U8452 (N_8452,N_8336,N_8367);
xnor U8453 (N_8453,N_8099,N_8227);
xor U8454 (N_8454,N_8338,N_8100);
nand U8455 (N_8455,N_8348,N_8150);
nor U8456 (N_8456,N_8036,N_8151);
nand U8457 (N_8457,N_8229,N_8314);
nand U8458 (N_8458,N_8098,N_8200);
nand U8459 (N_8459,N_8081,N_8077);
nor U8460 (N_8460,N_8148,N_8327);
xor U8461 (N_8461,N_8287,N_8272);
or U8462 (N_8462,N_8244,N_8021);
or U8463 (N_8463,N_8171,N_8383);
and U8464 (N_8464,N_8381,N_8088);
nor U8465 (N_8465,N_8035,N_8334);
nor U8466 (N_8466,N_8221,N_8231);
nand U8467 (N_8467,N_8264,N_8273);
nand U8468 (N_8468,N_8331,N_8155);
and U8469 (N_8469,N_8323,N_8268);
nand U8470 (N_8470,N_8014,N_8142);
nand U8471 (N_8471,N_8369,N_8167);
nand U8472 (N_8472,N_8356,N_8174);
xnor U8473 (N_8473,N_8319,N_8008);
nor U8474 (N_8474,N_8101,N_8175);
xor U8475 (N_8475,N_8145,N_8242);
xnor U8476 (N_8476,N_8324,N_8005);
nand U8477 (N_8477,N_8306,N_8198);
nor U8478 (N_8478,N_8311,N_8222);
nor U8479 (N_8479,N_8019,N_8308);
nand U8480 (N_8480,N_8206,N_8335);
nor U8481 (N_8481,N_8153,N_8004);
xor U8482 (N_8482,N_8165,N_8210);
xor U8483 (N_8483,N_8299,N_8195);
and U8484 (N_8484,N_8094,N_8283);
nor U8485 (N_8485,N_8031,N_8263);
xor U8486 (N_8486,N_8341,N_8149);
or U8487 (N_8487,N_8161,N_8013);
xnor U8488 (N_8488,N_8183,N_8300);
xnor U8489 (N_8489,N_8207,N_8320);
xnor U8490 (N_8490,N_8379,N_8205);
nor U8491 (N_8491,N_8059,N_8217);
xnor U8492 (N_8492,N_8223,N_8074);
nand U8493 (N_8493,N_8003,N_8002);
xor U8494 (N_8494,N_8307,N_8023);
xnor U8495 (N_8495,N_8238,N_8292);
nor U8496 (N_8496,N_8339,N_8213);
and U8497 (N_8497,N_8262,N_8360);
or U8498 (N_8498,N_8173,N_8116);
nor U8499 (N_8499,N_8376,N_8038);
nor U8500 (N_8500,N_8284,N_8026);
and U8501 (N_8501,N_8228,N_8093);
xnor U8502 (N_8502,N_8215,N_8140);
nor U8503 (N_8503,N_8258,N_8234);
and U8504 (N_8504,N_8240,N_8265);
xnor U8505 (N_8505,N_8007,N_8015);
nor U8506 (N_8506,N_8110,N_8117);
and U8507 (N_8507,N_8122,N_8092);
xor U8508 (N_8508,N_8037,N_8020);
xnor U8509 (N_8509,N_8157,N_8181);
nor U8510 (N_8510,N_8203,N_8134);
nand U8511 (N_8511,N_8224,N_8269);
nor U8512 (N_8512,N_8169,N_8281);
or U8513 (N_8513,N_8090,N_8297);
or U8514 (N_8514,N_8349,N_8000);
xnor U8515 (N_8515,N_8182,N_8166);
nor U8516 (N_8516,N_8131,N_8078);
xnor U8517 (N_8517,N_8040,N_8187);
nor U8518 (N_8518,N_8212,N_8084);
and U8519 (N_8519,N_8340,N_8274);
nand U8520 (N_8520,N_8184,N_8112);
nor U8521 (N_8521,N_8032,N_8313);
xnor U8522 (N_8522,N_8346,N_8371);
and U8523 (N_8523,N_8177,N_8178);
and U8524 (N_8524,N_8042,N_8130);
and U8525 (N_8525,N_8105,N_8066);
xor U8526 (N_8526,N_8393,N_8016);
or U8527 (N_8527,N_8018,N_8333);
and U8528 (N_8528,N_8214,N_8115);
xnor U8529 (N_8529,N_8337,N_8188);
nand U8530 (N_8530,N_8361,N_8382);
or U8531 (N_8531,N_8332,N_8294);
and U8532 (N_8532,N_8330,N_8255);
xnor U8533 (N_8533,N_8365,N_8022);
nand U8534 (N_8534,N_8127,N_8250);
or U8535 (N_8535,N_8043,N_8396);
nand U8536 (N_8536,N_8128,N_8135);
nor U8537 (N_8537,N_8104,N_8209);
nor U8538 (N_8538,N_8073,N_8072);
nand U8539 (N_8539,N_8106,N_8271);
and U8540 (N_8540,N_8129,N_8309);
xor U8541 (N_8541,N_8102,N_8103);
nand U8542 (N_8542,N_8082,N_8322);
or U8543 (N_8543,N_8114,N_8156);
or U8544 (N_8544,N_8179,N_8001);
nand U8545 (N_8545,N_8352,N_8154);
and U8546 (N_8546,N_8063,N_8218);
nor U8547 (N_8547,N_8044,N_8285);
or U8548 (N_8548,N_8276,N_8318);
or U8549 (N_8549,N_8252,N_8029);
nand U8550 (N_8550,N_8121,N_8241);
and U8551 (N_8551,N_8194,N_8164);
nand U8552 (N_8552,N_8049,N_8282);
nand U8553 (N_8553,N_8048,N_8235);
or U8554 (N_8554,N_8366,N_8219);
xnor U8555 (N_8555,N_8030,N_8278);
xor U8556 (N_8556,N_8261,N_8312);
nand U8557 (N_8557,N_8028,N_8061);
nor U8558 (N_8558,N_8254,N_8247);
nand U8559 (N_8559,N_8226,N_8147);
xor U8560 (N_8560,N_8041,N_8248);
or U8561 (N_8561,N_8375,N_8236);
nor U8562 (N_8562,N_8180,N_8033);
nand U8563 (N_8563,N_8251,N_8391);
nand U8564 (N_8564,N_8079,N_8270);
or U8565 (N_8565,N_8291,N_8399);
xor U8566 (N_8566,N_8342,N_8246);
xnor U8567 (N_8567,N_8133,N_8137);
nor U8568 (N_8568,N_8216,N_8053);
nand U8569 (N_8569,N_8310,N_8124);
and U8570 (N_8570,N_8232,N_8054);
xor U8571 (N_8571,N_8280,N_8243);
nand U8572 (N_8572,N_8253,N_8095);
nand U8573 (N_8573,N_8172,N_8071);
nor U8574 (N_8574,N_8304,N_8362);
nor U8575 (N_8575,N_8045,N_8380);
nor U8576 (N_8576,N_8359,N_8075);
or U8577 (N_8577,N_8316,N_8358);
nand U8578 (N_8578,N_8185,N_8317);
xnor U8579 (N_8579,N_8220,N_8067);
or U8580 (N_8580,N_8257,N_8196);
or U8581 (N_8581,N_8162,N_8363);
xnor U8582 (N_8582,N_8286,N_8370);
and U8583 (N_8583,N_8047,N_8368);
or U8584 (N_8584,N_8290,N_8111);
or U8585 (N_8585,N_8144,N_8266);
nand U8586 (N_8586,N_8080,N_8159);
xor U8587 (N_8587,N_8204,N_8158);
or U8588 (N_8588,N_8293,N_8344);
nor U8589 (N_8589,N_8141,N_8069);
or U8590 (N_8590,N_8189,N_8398);
or U8591 (N_8591,N_8107,N_8202);
and U8592 (N_8592,N_8132,N_8388);
xor U8593 (N_8593,N_8006,N_8056);
xor U8594 (N_8594,N_8027,N_8064);
xor U8595 (N_8595,N_8108,N_8392);
xnor U8596 (N_8596,N_8386,N_8357);
nand U8597 (N_8597,N_8328,N_8062);
and U8598 (N_8598,N_8190,N_8325);
nand U8599 (N_8599,N_8109,N_8230);
xnor U8600 (N_8600,N_8100,N_8095);
or U8601 (N_8601,N_8252,N_8242);
xor U8602 (N_8602,N_8150,N_8254);
or U8603 (N_8603,N_8384,N_8235);
nand U8604 (N_8604,N_8221,N_8225);
xor U8605 (N_8605,N_8046,N_8304);
or U8606 (N_8606,N_8018,N_8251);
and U8607 (N_8607,N_8224,N_8102);
and U8608 (N_8608,N_8383,N_8373);
and U8609 (N_8609,N_8127,N_8225);
xnor U8610 (N_8610,N_8393,N_8125);
and U8611 (N_8611,N_8139,N_8099);
and U8612 (N_8612,N_8007,N_8331);
or U8613 (N_8613,N_8042,N_8378);
nor U8614 (N_8614,N_8346,N_8328);
and U8615 (N_8615,N_8225,N_8390);
nor U8616 (N_8616,N_8338,N_8140);
xor U8617 (N_8617,N_8106,N_8363);
or U8618 (N_8618,N_8087,N_8252);
nor U8619 (N_8619,N_8131,N_8120);
nor U8620 (N_8620,N_8357,N_8124);
xnor U8621 (N_8621,N_8328,N_8297);
xnor U8622 (N_8622,N_8375,N_8294);
nor U8623 (N_8623,N_8055,N_8346);
nor U8624 (N_8624,N_8242,N_8011);
xnor U8625 (N_8625,N_8142,N_8255);
nand U8626 (N_8626,N_8166,N_8318);
and U8627 (N_8627,N_8118,N_8117);
and U8628 (N_8628,N_8346,N_8043);
or U8629 (N_8629,N_8256,N_8069);
xor U8630 (N_8630,N_8240,N_8158);
and U8631 (N_8631,N_8243,N_8232);
or U8632 (N_8632,N_8245,N_8395);
xnor U8633 (N_8633,N_8090,N_8088);
or U8634 (N_8634,N_8240,N_8165);
nor U8635 (N_8635,N_8262,N_8087);
nand U8636 (N_8636,N_8144,N_8175);
nand U8637 (N_8637,N_8127,N_8022);
xnor U8638 (N_8638,N_8238,N_8184);
nor U8639 (N_8639,N_8185,N_8150);
nand U8640 (N_8640,N_8028,N_8196);
xnor U8641 (N_8641,N_8192,N_8370);
or U8642 (N_8642,N_8057,N_8184);
xor U8643 (N_8643,N_8326,N_8066);
nand U8644 (N_8644,N_8051,N_8366);
or U8645 (N_8645,N_8175,N_8336);
nor U8646 (N_8646,N_8007,N_8339);
nor U8647 (N_8647,N_8030,N_8111);
xnor U8648 (N_8648,N_8057,N_8264);
xnor U8649 (N_8649,N_8312,N_8147);
nor U8650 (N_8650,N_8298,N_8320);
nor U8651 (N_8651,N_8296,N_8191);
xnor U8652 (N_8652,N_8354,N_8290);
or U8653 (N_8653,N_8343,N_8265);
nor U8654 (N_8654,N_8304,N_8257);
and U8655 (N_8655,N_8006,N_8210);
and U8656 (N_8656,N_8019,N_8383);
and U8657 (N_8657,N_8164,N_8131);
xor U8658 (N_8658,N_8311,N_8324);
nor U8659 (N_8659,N_8300,N_8026);
xor U8660 (N_8660,N_8221,N_8079);
and U8661 (N_8661,N_8079,N_8052);
xnor U8662 (N_8662,N_8268,N_8146);
or U8663 (N_8663,N_8371,N_8263);
and U8664 (N_8664,N_8002,N_8314);
nand U8665 (N_8665,N_8311,N_8036);
or U8666 (N_8666,N_8348,N_8390);
nor U8667 (N_8667,N_8187,N_8356);
nor U8668 (N_8668,N_8022,N_8186);
nand U8669 (N_8669,N_8147,N_8194);
nand U8670 (N_8670,N_8235,N_8378);
or U8671 (N_8671,N_8141,N_8152);
nor U8672 (N_8672,N_8382,N_8323);
and U8673 (N_8673,N_8199,N_8204);
and U8674 (N_8674,N_8120,N_8048);
xnor U8675 (N_8675,N_8050,N_8216);
and U8676 (N_8676,N_8128,N_8015);
nand U8677 (N_8677,N_8026,N_8108);
xor U8678 (N_8678,N_8187,N_8206);
or U8679 (N_8679,N_8144,N_8107);
xnor U8680 (N_8680,N_8182,N_8130);
xor U8681 (N_8681,N_8049,N_8396);
xnor U8682 (N_8682,N_8317,N_8104);
nand U8683 (N_8683,N_8064,N_8303);
nor U8684 (N_8684,N_8143,N_8024);
and U8685 (N_8685,N_8139,N_8019);
or U8686 (N_8686,N_8236,N_8040);
nor U8687 (N_8687,N_8162,N_8214);
nor U8688 (N_8688,N_8217,N_8290);
or U8689 (N_8689,N_8323,N_8003);
nor U8690 (N_8690,N_8012,N_8054);
nand U8691 (N_8691,N_8332,N_8123);
and U8692 (N_8692,N_8166,N_8073);
or U8693 (N_8693,N_8292,N_8105);
nand U8694 (N_8694,N_8017,N_8367);
nor U8695 (N_8695,N_8342,N_8022);
or U8696 (N_8696,N_8096,N_8178);
and U8697 (N_8697,N_8374,N_8071);
xnor U8698 (N_8698,N_8194,N_8080);
nor U8699 (N_8699,N_8226,N_8369);
and U8700 (N_8700,N_8370,N_8217);
nand U8701 (N_8701,N_8396,N_8273);
nand U8702 (N_8702,N_8214,N_8074);
nand U8703 (N_8703,N_8142,N_8325);
nand U8704 (N_8704,N_8178,N_8395);
nor U8705 (N_8705,N_8353,N_8066);
or U8706 (N_8706,N_8297,N_8227);
and U8707 (N_8707,N_8098,N_8276);
and U8708 (N_8708,N_8103,N_8069);
xor U8709 (N_8709,N_8043,N_8048);
or U8710 (N_8710,N_8313,N_8316);
nand U8711 (N_8711,N_8098,N_8131);
or U8712 (N_8712,N_8007,N_8201);
or U8713 (N_8713,N_8249,N_8376);
xor U8714 (N_8714,N_8364,N_8331);
or U8715 (N_8715,N_8193,N_8028);
or U8716 (N_8716,N_8083,N_8016);
or U8717 (N_8717,N_8270,N_8369);
and U8718 (N_8718,N_8052,N_8140);
nor U8719 (N_8719,N_8021,N_8180);
nor U8720 (N_8720,N_8360,N_8204);
or U8721 (N_8721,N_8273,N_8279);
nand U8722 (N_8722,N_8014,N_8316);
nor U8723 (N_8723,N_8071,N_8328);
nor U8724 (N_8724,N_8051,N_8013);
nand U8725 (N_8725,N_8042,N_8218);
nor U8726 (N_8726,N_8390,N_8332);
xor U8727 (N_8727,N_8190,N_8197);
or U8728 (N_8728,N_8190,N_8021);
nand U8729 (N_8729,N_8199,N_8061);
or U8730 (N_8730,N_8153,N_8284);
or U8731 (N_8731,N_8162,N_8079);
and U8732 (N_8732,N_8204,N_8082);
nand U8733 (N_8733,N_8111,N_8075);
nor U8734 (N_8734,N_8184,N_8356);
and U8735 (N_8735,N_8153,N_8228);
xnor U8736 (N_8736,N_8010,N_8064);
and U8737 (N_8737,N_8255,N_8079);
xor U8738 (N_8738,N_8110,N_8087);
nor U8739 (N_8739,N_8112,N_8208);
nor U8740 (N_8740,N_8203,N_8048);
nor U8741 (N_8741,N_8364,N_8227);
or U8742 (N_8742,N_8344,N_8051);
nand U8743 (N_8743,N_8174,N_8007);
xor U8744 (N_8744,N_8290,N_8220);
xor U8745 (N_8745,N_8080,N_8296);
nor U8746 (N_8746,N_8377,N_8277);
and U8747 (N_8747,N_8042,N_8007);
xor U8748 (N_8748,N_8123,N_8141);
and U8749 (N_8749,N_8279,N_8190);
nand U8750 (N_8750,N_8298,N_8219);
and U8751 (N_8751,N_8207,N_8346);
xor U8752 (N_8752,N_8239,N_8129);
or U8753 (N_8753,N_8220,N_8358);
nand U8754 (N_8754,N_8187,N_8318);
xnor U8755 (N_8755,N_8302,N_8380);
and U8756 (N_8756,N_8120,N_8335);
nor U8757 (N_8757,N_8035,N_8104);
nand U8758 (N_8758,N_8235,N_8294);
xnor U8759 (N_8759,N_8065,N_8130);
nor U8760 (N_8760,N_8214,N_8167);
and U8761 (N_8761,N_8248,N_8384);
nand U8762 (N_8762,N_8080,N_8344);
and U8763 (N_8763,N_8200,N_8082);
xnor U8764 (N_8764,N_8245,N_8065);
xor U8765 (N_8765,N_8023,N_8155);
nand U8766 (N_8766,N_8068,N_8072);
nor U8767 (N_8767,N_8069,N_8051);
and U8768 (N_8768,N_8340,N_8193);
nor U8769 (N_8769,N_8099,N_8337);
or U8770 (N_8770,N_8390,N_8058);
or U8771 (N_8771,N_8007,N_8053);
xor U8772 (N_8772,N_8214,N_8139);
nand U8773 (N_8773,N_8253,N_8039);
or U8774 (N_8774,N_8325,N_8130);
nand U8775 (N_8775,N_8033,N_8068);
xor U8776 (N_8776,N_8031,N_8094);
or U8777 (N_8777,N_8173,N_8204);
xnor U8778 (N_8778,N_8341,N_8152);
or U8779 (N_8779,N_8186,N_8181);
xor U8780 (N_8780,N_8121,N_8075);
and U8781 (N_8781,N_8068,N_8009);
or U8782 (N_8782,N_8178,N_8086);
xor U8783 (N_8783,N_8396,N_8270);
xnor U8784 (N_8784,N_8164,N_8373);
and U8785 (N_8785,N_8327,N_8005);
nor U8786 (N_8786,N_8187,N_8342);
or U8787 (N_8787,N_8343,N_8272);
xor U8788 (N_8788,N_8043,N_8159);
nor U8789 (N_8789,N_8338,N_8390);
nand U8790 (N_8790,N_8328,N_8093);
nand U8791 (N_8791,N_8180,N_8288);
or U8792 (N_8792,N_8391,N_8030);
and U8793 (N_8793,N_8029,N_8058);
and U8794 (N_8794,N_8089,N_8261);
xnor U8795 (N_8795,N_8390,N_8093);
nor U8796 (N_8796,N_8388,N_8164);
xnor U8797 (N_8797,N_8282,N_8261);
nor U8798 (N_8798,N_8104,N_8008);
and U8799 (N_8799,N_8360,N_8260);
or U8800 (N_8800,N_8633,N_8629);
nor U8801 (N_8801,N_8702,N_8603);
nor U8802 (N_8802,N_8609,N_8585);
and U8803 (N_8803,N_8599,N_8761);
or U8804 (N_8804,N_8671,N_8708);
and U8805 (N_8805,N_8605,N_8455);
xnor U8806 (N_8806,N_8524,N_8746);
nand U8807 (N_8807,N_8411,N_8622);
xor U8808 (N_8808,N_8707,N_8744);
xnor U8809 (N_8809,N_8548,N_8688);
xnor U8810 (N_8810,N_8793,N_8491);
nor U8811 (N_8811,N_8578,N_8695);
or U8812 (N_8812,N_8452,N_8525);
and U8813 (N_8813,N_8617,N_8598);
xor U8814 (N_8814,N_8677,N_8637);
or U8815 (N_8815,N_8409,N_8659);
and U8816 (N_8816,N_8780,N_8459);
xor U8817 (N_8817,N_8626,N_8787);
xnor U8818 (N_8818,N_8588,N_8748);
nor U8819 (N_8819,N_8709,N_8541);
nor U8820 (N_8820,N_8571,N_8697);
and U8821 (N_8821,N_8631,N_8667);
and U8822 (N_8822,N_8754,N_8500);
or U8823 (N_8823,N_8757,N_8597);
nor U8824 (N_8824,N_8489,N_8447);
nand U8825 (N_8825,N_8666,N_8435);
xor U8826 (N_8826,N_8678,N_8503);
and U8827 (N_8827,N_8621,N_8612);
and U8828 (N_8828,N_8499,N_8451);
nor U8829 (N_8829,N_8798,N_8574);
nand U8830 (N_8830,N_8752,N_8508);
nor U8831 (N_8831,N_8795,N_8649);
xnor U8832 (N_8832,N_8783,N_8657);
and U8833 (N_8833,N_8547,N_8774);
nor U8834 (N_8834,N_8786,N_8427);
nor U8835 (N_8835,N_8497,N_8521);
nor U8836 (N_8836,N_8410,N_8462);
nand U8837 (N_8837,N_8767,N_8401);
xor U8838 (N_8838,N_8660,N_8593);
xor U8839 (N_8839,N_8737,N_8625);
xor U8840 (N_8840,N_8782,N_8791);
nor U8841 (N_8841,N_8794,N_8572);
nor U8842 (N_8842,N_8444,N_8797);
nand U8843 (N_8843,N_8472,N_8400);
nand U8844 (N_8844,N_8712,N_8681);
nand U8845 (N_8845,N_8454,N_8670);
and U8846 (N_8846,N_8556,N_8747);
nand U8847 (N_8847,N_8422,N_8638);
xnor U8848 (N_8848,N_8545,N_8537);
or U8849 (N_8849,N_8762,N_8564);
or U8850 (N_8850,N_8724,N_8692);
or U8851 (N_8851,N_8531,N_8604);
nor U8852 (N_8852,N_8554,N_8471);
and U8853 (N_8853,N_8720,N_8738);
xnor U8854 (N_8854,N_8779,N_8650);
nand U8855 (N_8855,N_8705,N_8716);
and U8856 (N_8856,N_8769,N_8680);
nand U8857 (N_8857,N_8778,N_8546);
and U8858 (N_8858,N_8682,N_8684);
nand U8859 (N_8859,N_8405,N_8492);
or U8860 (N_8860,N_8421,N_8674);
xnor U8861 (N_8861,N_8721,N_8723);
or U8862 (N_8862,N_8656,N_8696);
or U8863 (N_8863,N_8713,N_8763);
or U8864 (N_8864,N_8628,N_8504);
xnor U8865 (N_8865,N_8490,N_8722);
nand U8866 (N_8866,N_8466,N_8602);
nor U8867 (N_8867,N_8557,N_8408);
nand U8868 (N_8868,N_8461,N_8584);
and U8869 (N_8869,N_8523,N_8542);
nand U8870 (N_8870,N_8736,N_8594);
nor U8871 (N_8871,N_8469,N_8580);
or U8872 (N_8872,N_8544,N_8683);
nor U8873 (N_8873,N_8424,N_8648);
xor U8874 (N_8874,N_8474,N_8565);
nor U8875 (N_8875,N_8570,N_8642);
nor U8876 (N_8876,N_8618,N_8507);
nor U8877 (N_8877,N_8442,N_8481);
xor U8878 (N_8878,N_8776,N_8620);
nor U8879 (N_8879,N_8711,N_8479);
and U8880 (N_8880,N_8669,N_8511);
or U8881 (N_8881,N_8536,N_8607);
xor U8882 (N_8882,N_8627,N_8581);
nor U8883 (N_8883,N_8756,N_8413);
or U8884 (N_8884,N_8645,N_8549);
nor U8885 (N_8885,N_8520,N_8687);
and U8886 (N_8886,N_8781,N_8750);
xnor U8887 (N_8887,N_8543,N_8784);
or U8888 (N_8888,N_8582,N_8733);
xnor U8889 (N_8889,N_8701,N_8575);
and U8890 (N_8890,N_8509,N_8691);
nor U8891 (N_8891,N_8475,N_8426);
or U8892 (N_8892,N_8792,N_8685);
nand U8893 (N_8893,N_8694,N_8495);
xnor U8894 (N_8894,N_8592,N_8486);
nand U8895 (N_8895,N_8600,N_8505);
and U8896 (N_8896,N_8601,N_8415);
nand U8897 (N_8897,N_8457,N_8640);
and U8898 (N_8898,N_8758,N_8412);
or U8899 (N_8899,N_8676,N_8653);
or U8900 (N_8900,N_8573,N_8577);
xnor U8901 (N_8901,N_8539,N_8561);
nor U8902 (N_8902,N_8477,N_8689);
nor U8903 (N_8903,N_8519,N_8552);
nand U8904 (N_8904,N_8773,N_8587);
nor U8905 (N_8905,N_8501,N_8586);
nand U8906 (N_8906,N_8624,N_8726);
nor U8907 (N_8907,N_8514,N_8406);
nand U8908 (N_8908,N_8460,N_8432);
nand U8909 (N_8909,N_8735,N_8517);
or U8910 (N_8910,N_8772,N_8731);
nand U8911 (N_8911,N_8483,N_8465);
xor U8912 (N_8912,N_8771,N_8431);
nand U8913 (N_8913,N_8765,N_8510);
xnor U8914 (N_8914,N_8550,N_8576);
xor U8915 (N_8915,N_8743,N_8718);
nor U8916 (N_8916,N_8560,N_8438);
nand U8917 (N_8917,N_8568,N_8799);
or U8918 (N_8918,N_8567,N_8518);
nor U8919 (N_8919,N_8719,N_8698);
xor U8920 (N_8920,N_8608,N_8533);
or U8921 (N_8921,N_8606,N_8555);
nand U8922 (N_8922,N_8796,N_8652);
xor U8923 (N_8923,N_8651,N_8591);
xor U8924 (N_8924,N_8615,N_8540);
or U8925 (N_8925,N_8703,N_8407);
and U8926 (N_8926,N_8453,N_8436);
nor U8927 (N_8927,N_8636,N_8693);
or U8928 (N_8928,N_8589,N_8535);
nor U8929 (N_8929,N_8704,N_8751);
and U8930 (N_8930,N_8727,N_8498);
or U8931 (N_8931,N_8528,N_8658);
and U8932 (N_8932,N_8742,N_8429);
or U8933 (N_8933,N_8428,N_8732);
and U8934 (N_8934,N_8714,N_8632);
xnor U8935 (N_8935,N_8559,N_8595);
xnor U8936 (N_8936,N_8663,N_8473);
and U8937 (N_8937,N_8450,N_8423);
xor U8938 (N_8938,N_8506,N_8513);
xor U8939 (N_8939,N_8641,N_8488);
nor U8940 (N_8940,N_8686,N_8456);
nor U8941 (N_8941,N_8515,N_8777);
nor U8942 (N_8942,N_8614,N_8467);
xor U8943 (N_8943,N_8458,N_8534);
nand U8944 (N_8944,N_8749,N_8646);
nand U8945 (N_8945,N_8527,N_8717);
or U8946 (N_8946,N_8635,N_8416);
nand U8947 (N_8947,N_8404,N_8654);
and U8948 (N_8948,N_8493,N_8643);
nor U8949 (N_8949,N_8664,N_8482);
nand U8950 (N_8950,N_8553,N_8430);
and U8951 (N_8951,N_8433,N_8579);
and U8952 (N_8952,N_8526,N_8655);
xor U8953 (N_8953,N_8496,N_8502);
xor U8954 (N_8954,N_8419,N_8788);
or U8955 (N_8955,N_8484,N_8785);
and U8956 (N_8956,N_8741,N_8789);
xor U8957 (N_8957,N_8672,N_8730);
or U8958 (N_8958,N_8437,N_8449);
or U8959 (N_8959,N_8690,N_8480);
nand U8960 (N_8960,N_8764,N_8468);
and U8961 (N_8961,N_8700,N_8661);
nand U8962 (N_8962,N_8551,N_8558);
nand U8963 (N_8963,N_8522,N_8734);
or U8964 (N_8964,N_8699,N_8745);
or U8965 (N_8965,N_8464,N_8402);
nor U8966 (N_8966,N_8644,N_8538);
nor U8967 (N_8967,N_8770,N_8446);
xnor U8968 (N_8968,N_8619,N_8755);
nand U8969 (N_8969,N_8706,N_8403);
and U8970 (N_8970,N_8616,N_8476);
and U8971 (N_8971,N_8417,N_8739);
nor U8972 (N_8972,N_8566,N_8516);
nand U8973 (N_8973,N_8441,N_8434);
nor U8974 (N_8974,N_8532,N_8775);
xor U8975 (N_8975,N_8759,N_8463);
or U8976 (N_8976,N_8443,N_8665);
and U8977 (N_8977,N_8623,N_8647);
nor U8978 (N_8978,N_8418,N_8611);
nand U8979 (N_8979,N_8420,N_8583);
xor U8980 (N_8980,N_8448,N_8679);
or U8981 (N_8981,N_8753,N_8610);
nor U8982 (N_8982,N_8414,N_8662);
xnor U8983 (N_8983,N_8439,N_8634);
or U8984 (N_8984,N_8760,N_8639);
xor U8985 (N_8985,N_8725,N_8729);
xnor U8986 (N_8986,N_8494,N_8512);
xor U8987 (N_8987,N_8740,N_8529);
nand U8988 (N_8988,N_8766,N_8728);
nor U8989 (N_8989,N_8445,N_8485);
nor U8990 (N_8990,N_8569,N_8530);
and U8991 (N_8991,N_8562,N_8790);
xnor U8992 (N_8992,N_8613,N_8470);
xor U8993 (N_8993,N_8563,N_8710);
nor U8994 (N_8994,N_8425,N_8596);
nor U8995 (N_8995,N_8673,N_8590);
xor U8996 (N_8996,N_8715,N_8768);
or U8997 (N_8997,N_8440,N_8630);
or U8998 (N_8998,N_8478,N_8668);
or U8999 (N_8999,N_8675,N_8487);
xnor U9000 (N_9000,N_8616,N_8584);
nor U9001 (N_9001,N_8693,N_8611);
xor U9002 (N_9002,N_8492,N_8783);
xor U9003 (N_9003,N_8648,N_8772);
and U9004 (N_9004,N_8668,N_8463);
and U9005 (N_9005,N_8500,N_8682);
nor U9006 (N_9006,N_8588,N_8405);
xor U9007 (N_9007,N_8747,N_8624);
nor U9008 (N_9008,N_8468,N_8558);
xnor U9009 (N_9009,N_8415,N_8687);
xnor U9010 (N_9010,N_8556,N_8735);
xor U9011 (N_9011,N_8652,N_8547);
nor U9012 (N_9012,N_8751,N_8640);
xor U9013 (N_9013,N_8511,N_8448);
or U9014 (N_9014,N_8688,N_8476);
and U9015 (N_9015,N_8661,N_8507);
nand U9016 (N_9016,N_8404,N_8602);
nand U9017 (N_9017,N_8770,N_8430);
or U9018 (N_9018,N_8667,N_8648);
or U9019 (N_9019,N_8643,N_8451);
xor U9020 (N_9020,N_8773,N_8438);
nand U9021 (N_9021,N_8456,N_8592);
xor U9022 (N_9022,N_8597,N_8633);
nor U9023 (N_9023,N_8534,N_8473);
and U9024 (N_9024,N_8511,N_8657);
and U9025 (N_9025,N_8693,N_8676);
nor U9026 (N_9026,N_8480,N_8638);
xor U9027 (N_9027,N_8444,N_8547);
nand U9028 (N_9028,N_8748,N_8517);
xor U9029 (N_9029,N_8464,N_8530);
xor U9030 (N_9030,N_8760,N_8656);
xor U9031 (N_9031,N_8479,N_8701);
and U9032 (N_9032,N_8543,N_8771);
and U9033 (N_9033,N_8578,N_8677);
nand U9034 (N_9034,N_8702,N_8573);
xor U9035 (N_9035,N_8428,N_8635);
nor U9036 (N_9036,N_8658,N_8752);
or U9037 (N_9037,N_8440,N_8532);
nor U9038 (N_9038,N_8748,N_8413);
xor U9039 (N_9039,N_8465,N_8732);
nor U9040 (N_9040,N_8758,N_8541);
nor U9041 (N_9041,N_8769,N_8484);
nand U9042 (N_9042,N_8724,N_8661);
xnor U9043 (N_9043,N_8471,N_8715);
xnor U9044 (N_9044,N_8769,N_8566);
nor U9045 (N_9045,N_8671,N_8698);
and U9046 (N_9046,N_8573,N_8604);
and U9047 (N_9047,N_8759,N_8612);
nor U9048 (N_9048,N_8559,N_8543);
and U9049 (N_9049,N_8669,N_8718);
nand U9050 (N_9050,N_8737,N_8751);
nand U9051 (N_9051,N_8527,N_8431);
or U9052 (N_9052,N_8797,N_8507);
nand U9053 (N_9053,N_8606,N_8785);
xnor U9054 (N_9054,N_8489,N_8683);
nand U9055 (N_9055,N_8711,N_8702);
nand U9056 (N_9056,N_8739,N_8580);
and U9057 (N_9057,N_8734,N_8753);
and U9058 (N_9058,N_8541,N_8677);
xor U9059 (N_9059,N_8400,N_8538);
xor U9060 (N_9060,N_8400,N_8754);
nor U9061 (N_9061,N_8707,N_8779);
nand U9062 (N_9062,N_8446,N_8468);
or U9063 (N_9063,N_8614,N_8443);
or U9064 (N_9064,N_8519,N_8631);
nand U9065 (N_9065,N_8588,N_8694);
and U9066 (N_9066,N_8754,N_8511);
xnor U9067 (N_9067,N_8481,N_8477);
or U9068 (N_9068,N_8756,N_8677);
xor U9069 (N_9069,N_8653,N_8670);
nand U9070 (N_9070,N_8505,N_8723);
xnor U9071 (N_9071,N_8430,N_8660);
or U9072 (N_9072,N_8658,N_8471);
and U9073 (N_9073,N_8721,N_8774);
nand U9074 (N_9074,N_8603,N_8470);
nand U9075 (N_9075,N_8574,N_8781);
or U9076 (N_9076,N_8539,N_8460);
and U9077 (N_9077,N_8416,N_8655);
xnor U9078 (N_9078,N_8455,N_8743);
xor U9079 (N_9079,N_8677,N_8454);
or U9080 (N_9080,N_8536,N_8690);
nand U9081 (N_9081,N_8531,N_8754);
or U9082 (N_9082,N_8404,N_8790);
xnor U9083 (N_9083,N_8440,N_8679);
nand U9084 (N_9084,N_8607,N_8581);
xor U9085 (N_9085,N_8469,N_8799);
and U9086 (N_9086,N_8616,N_8582);
nor U9087 (N_9087,N_8402,N_8509);
nand U9088 (N_9088,N_8762,N_8771);
nand U9089 (N_9089,N_8441,N_8781);
and U9090 (N_9090,N_8421,N_8574);
nor U9091 (N_9091,N_8615,N_8531);
nor U9092 (N_9092,N_8477,N_8421);
nand U9093 (N_9093,N_8415,N_8525);
nand U9094 (N_9094,N_8443,N_8515);
or U9095 (N_9095,N_8562,N_8703);
nand U9096 (N_9096,N_8548,N_8658);
or U9097 (N_9097,N_8656,N_8551);
and U9098 (N_9098,N_8737,N_8427);
nand U9099 (N_9099,N_8694,N_8607);
or U9100 (N_9100,N_8623,N_8515);
nand U9101 (N_9101,N_8669,N_8404);
xnor U9102 (N_9102,N_8470,N_8731);
nor U9103 (N_9103,N_8730,N_8732);
nor U9104 (N_9104,N_8540,N_8754);
and U9105 (N_9105,N_8711,N_8474);
nor U9106 (N_9106,N_8429,N_8790);
and U9107 (N_9107,N_8610,N_8724);
xor U9108 (N_9108,N_8422,N_8652);
or U9109 (N_9109,N_8402,N_8403);
nand U9110 (N_9110,N_8755,N_8613);
or U9111 (N_9111,N_8775,N_8707);
or U9112 (N_9112,N_8605,N_8405);
nand U9113 (N_9113,N_8682,N_8521);
nand U9114 (N_9114,N_8729,N_8400);
or U9115 (N_9115,N_8764,N_8553);
and U9116 (N_9116,N_8662,N_8783);
xor U9117 (N_9117,N_8758,N_8621);
and U9118 (N_9118,N_8634,N_8550);
nand U9119 (N_9119,N_8417,N_8494);
and U9120 (N_9120,N_8550,N_8623);
xor U9121 (N_9121,N_8714,N_8588);
xor U9122 (N_9122,N_8751,N_8602);
nand U9123 (N_9123,N_8544,N_8466);
or U9124 (N_9124,N_8731,N_8528);
nor U9125 (N_9125,N_8747,N_8679);
nand U9126 (N_9126,N_8644,N_8659);
nand U9127 (N_9127,N_8588,N_8629);
or U9128 (N_9128,N_8732,N_8784);
nor U9129 (N_9129,N_8616,N_8679);
nand U9130 (N_9130,N_8740,N_8542);
nor U9131 (N_9131,N_8741,N_8528);
nand U9132 (N_9132,N_8674,N_8784);
or U9133 (N_9133,N_8717,N_8707);
or U9134 (N_9134,N_8774,N_8703);
xor U9135 (N_9135,N_8531,N_8493);
xor U9136 (N_9136,N_8640,N_8403);
nor U9137 (N_9137,N_8571,N_8515);
or U9138 (N_9138,N_8477,N_8480);
or U9139 (N_9139,N_8549,N_8451);
nand U9140 (N_9140,N_8682,N_8574);
or U9141 (N_9141,N_8663,N_8637);
or U9142 (N_9142,N_8449,N_8789);
xor U9143 (N_9143,N_8790,N_8581);
and U9144 (N_9144,N_8553,N_8450);
nand U9145 (N_9145,N_8745,N_8407);
xor U9146 (N_9146,N_8743,N_8692);
and U9147 (N_9147,N_8430,N_8455);
or U9148 (N_9148,N_8494,N_8778);
nor U9149 (N_9149,N_8537,N_8690);
and U9150 (N_9150,N_8406,N_8717);
or U9151 (N_9151,N_8714,N_8761);
nand U9152 (N_9152,N_8704,N_8667);
xor U9153 (N_9153,N_8411,N_8429);
nor U9154 (N_9154,N_8583,N_8452);
or U9155 (N_9155,N_8454,N_8613);
and U9156 (N_9156,N_8583,N_8472);
xor U9157 (N_9157,N_8495,N_8731);
nor U9158 (N_9158,N_8616,N_8461);
xnor U9159 (N_9159,N_8603,N_8782);
or U9160 (N_9160,N_8756,N_8500);
xnor U9161 (N_9161,N_8440,N_8677);
nor U9162 (N_9162,N_8537,N_8561);
nor U9163 (N_9163,N_8637,N_8679);
and U9164 (N_9164,N_8776,N_8772);
nand U9165 (N_9165,N_8448,N_8760);
or U9166 (N_9166,N_8498,N_8635);
and U9167 (N_9167,N_8773,N_8607);
or U9168 (N_9168,N_8445,N_8469);
and U9169 (N_9169,N_8500,N_8577);
or U9170 (N_9170,N_8414,N_8517);
nor U9171 (N_9171,N_8403,N_8661);
and U9172 (N_9172,N_8407,N_8573);
and U9173 (N_9173,N_8529,N_8572);
xor U9174 (N_9174,N_8592,N_8692);
nor U9175 (N_9175,N_8519,N_8490);
nand U9176 (N_9176,N_8607,N_8652);
xor U9177 (N_9177,N_8502,N_8504);
nand U9178 (N_9178,N_8533,N_8536);
xor U9179 (N_9179,N_8628,N_8797);
or U9180 (N_9180,N_8645,N_8474);
xnor U9181 (N_9181,N_8758,N_8655);
nor U9182 (N_9182,N_8556,N_8669);
or U9183 (N_9183,N_8466,N_8748);
xnor U9184 (N_9184,N_8556,N_8745);
nand U9185 (N_9185,N_8656,N_8783);
or U9186 (N_9186,N_8645,N_8484);
and U9187 (N_9187,N_8640,N_8590);
and U9188 (N_9188,N_8570,N_8579);
nand U9189 (N_9189,N_8594,N_8758);
xor U9190 (N_9190,N_8789,N_8683);
xor U9191 (N_9191,N_8740,N_8410);
nor U9192 (N_9192,N_8434,N_8427);
or U9193 (N_9193,N_8568,N_8407);
nor U9194 (N_9194,N_8765,N_8577);
nor U9195 (N_9195,N_8557,N_8423);
xor U9196 (N_9196,N_8687,N_8796);
xor U9197 (N_9197,N_8652,N_8795);
xnor U9198 (N_9198,N_8760,N_8459);
and U9199 (N_9199,N_8529,N_8536);
nand U9200 (N_9200,N_8807,N_8829);
nor U9201 (N_9201,N_8822,N_9156);
nand U9202 (N_9202,N_8948,N_9005);
xnor U9203 (N_9203,N_9189,N_9131);
nor U9204 (N_9204,N_9122,N_9089);
and U9205 (N_9205,N_8811,N_9107);
or U9206 (N_9206,N_9153,N_9094);
or U9207 (N_9207,N_8824,N_8989);
and U9208 (N_9208,N_8936,N_9025);
nand U9209 (N_9209,N_9098,N_9178);
nand U9210 (N_9210,N_8944,N_8814);
nor U9211 (N_9211,N_8970,N_9149);
nor U9212 (N_9212,N_9069,N_9195);
and U9213 (N_9213,N_9079,N_8832);
nor U9214 (N_9214,N_9148,N_9150);
and U9215 (N_9215,N_8867,N_9099);
nand U9216 (N_9216,N_9046,N_8966);
nand U9217 (N_9217,N_8837,N_8841);
xnor U9218 (N_9218,N_9001,N_9093);
or U9219 (N_9219,N_8945,N_9115);
nor U9220 (N_9220,N_8800,N_8911);
and U9221 (N_9221,N_8886,N_9187);
nor U9222 (N_9222,N_8958,N_9143);
and U9223 (N_9223,N_9038,N_8889);
or U9224 (N_9224,N_9108,N_9052);
and U9225 (N_9225,N_9063,N_9049);
xor U9226 (N_9226,N_9065,N_8918);
xnor U9227 (N_9227,N_9197,N_9062);
and U9228 (N_9228,N_9152,N_9003);
nor U9229 (N_9229,N_9169,N_9088);
and U9230 (N_9230,N_9196,N_8981);
and U9231 (N_9231,N_9092,N_8825);
and U9232 (N_9232,N_9199,N_8879);
or U9233 (N_9233,N_9112,N_8977);
nand U9234 (N_9234,N_8908,N_8852);
xnor U9235 (N_9235,N_9055,N_8940);
or U9236 (N_9236,N_8850,N_8969);
xnor U9237 (N_9237,N_8866,N_9004);
nand U9238 (N_9238,N_9159,N_8872);
nand U9239 (N_9239,N_9076,N_8817);
xnor U9240 (N_9240,N_9000,N_9158);
xnor U9241 (N_9241,N_8952,N_9124);
nand U9242 (N_9242,N_8818,N_8883);
or U9243 (N_9243,N_9028,N_8968);
nor U9244 (N_9244,N_9032,N_8967);
and U9245 (N_9245,N_8845,N_9100);
or U9246 (N_9246,N_8954,N_9043);
or U9247 (N_9247,N_8887,N_8991);
or U9248 (N_9248,N_9194,N_8890);
xnor U9249 (N_9249,N_9192,N_9008);
or U9250 (N_9250,N_8942,N_9014);
xnor U9251 (N_9251,N_8851,N_8869);
nand U9252 (N_9252,N_8858,N_9177);
xor U9253 (N_9253,N_9051,N_8894);
nand U9254 (N_9254,N_8877,N_9030);
xor U9255 (N_9255,N_9012,N_9002);
xor U9256 (N_9256,N_8934,N_8881);
nor U9257 (N_9257,N_9050,N_8932);
nor U9258 (N_9258,N_8802,N_8979);
nand U9259 (N_9259,N_8855,N_9132);
nand U9260 (N_9260,N_8860,N_8861);
or U9261 (N_9261,N_9072,N_9057);
nand U9262 (N_9262,N_8836,N_9058);
and U9263 (N_9263,N_8900,N_8997);
nand U9264 (N_9264,N_8804,N_9091);
xnor U9265 (N_9265,N_8941,N_8904);
nand U9266 (N_9266,N_9070,N_8957);
and U9267 (N_9267,N_8853,N_8835);
nand U9268 (N_9268,N_9027,N_8924);
xnor U9269 (N_9269,N_8930,N_8923);
nor U9270 (N_9270,N_8986,N_9162);
nor U9271 (N_9271,N_8812,N_9024);
or U9272 (N_9272,N_9082,N_9154);
or U9273 (N_9273,N_9193,N_9142);
nor U9274 (N_9274,N_9133,N_8976);
or U9275 (N_9275,N_9015,N_8990);
nor U9276 (N_9276,N_9114,N_8899);
and U9277 (N_9277,N_9117,N_9116);
nor U9278 (N_9278,N_8959,N_9085);
xor U9279 (N_9279,N_8839,N_9007);
nor U9280 (N_9280,N_8819,N_8913);
or U9281 (N_9281,N_8999,N_8985);
nand U9282 (N_9282,N_8917,N_8947);
nor U9283 (N_9283,N_8992,N_8928);
or U9284 (N_9284,N_8865,N_9066);
nor U9285 (N_9285,N_9145,N_8809);
nor U9286 (N_9286,N_8826,N_8823);
and U9287 (N_9287,N_9056,N_9119);
or U9288 (N_9288,N_9184,N_8962);
xor U9289 (N_9289,N_8854,N_8827);
nor U9290 (N_9290,N_8916,N_9134);
nand U9291 (N_9291,N_9101,N_8974);
xnor U9292 (N_9292,N_8975,N_9074);
or U9293 (N_9293,N_8933,N_9037);
xnor U9294 (N_9294,N_8960,N_9035);
nand U9295 (N_9295,N_8920,N_8840);
and U9296 (N_9296,N_9160,N_9110);
or U9297 (N_9297,N_8888,N_8863);
nor U9298 (N_9298,N_9047,N_9186);
or U9299 (N_9299,N_8963,N_8983);
and U9300 (N_9300,N_8898,N_9164);
and U9301 (N_9301,N_9054,N_9146);
xnor U9302 (N_9302,N_9044,N_8955);
and U9303 (N_9303,N_8856,N_9073);
nor U9304 (N_9304,N_8919,N_9176);
nor U9305 (N_9305,N_8998,N_9022);
xor U9306 (N_9306,N_8939,N_9118);
xor U9307 (N_9307,N_8834,N_8831);
nand U9308 (N_9308,N_9060,N_9151);
xnor U9309 (N_9309,N_9139,N_8864);
and U9310 (N_9310,N_8956,N_8874);
xnor U9311 (N_9311,N_9130,N_8922);
xor U9312 (N_9312,N_9041,N_9109);
nor U9313 (N_9313,N_8891,N_9053);
or U9314 (N_9314,N_9113,N_9059);
and U9315 (N_9315,N_9147,N_8984);
xor U9316 (N_9316,N_8805,N_9067);
nand U9317 (N_9317,N_8848,N_8878);
or U9318 (N_9318,N_9077,N_9080);
and U9319 (N_9319,N_9026,N_8849);
nor U9320 (N_9320,N_9031,N_8902);
nand U9321 (N_9321,N_9138,N_9182);
and U9322 (N_9322,N_8870,N_9157);
nand U9323 (N_9323,N_8915,N_9121);
xnor U9324 (N_9324,N_8843,N_8830);
nor U9325 (N_9325,N_9048,N_8921);
or U9326 (N_9326,N_9165,N_8876);
xnor U9327 (N_9327,N_9068,N_9128);
nor U9328 (N_9328,N_8808,N_8821);
nand U9329 (N_9329,N_8972,N_9102);
nor U9330 (N_9330,N_8816,N_8885);
and U9331 (N_9331,N_9111,N_8906);
and U9332 (N_9332,N_9135,N_9191);
xor U9333 (N_9333,N_8937,N_8842);
nor U9334 (N_9334,N_8912,N_9009);
nand U9335 (N_9335,N_9019,N_8910);
nand U9336 (N_9336,N_9020,N_8896);
or U9337 (N_9337,N_8873,N_9179);
and U9338 (N_9338,N_9161,N_8938);
or U9339 (N_9339,N_8995,N_9140);
or U9340 (N_9340,N_9018,N_8844);
xor U9341 (N_9341,N_9011,N_8961);
xor U9342 (N_9342,N_9181,N_9075);
and U9343 (N_9343,N_9084,N_8838);
and U9344 (N_9344,N_8965,N_9125);
xor U9345 (N_9345,N_9104,N_9010);
or U9346 (N_9346,N_8880,N_9036);
xnor U9347 (N_9347,N_8857,N_8813);
nand U9348 (N_9348,N_8982,N_9168);
or U9349 (N_9349,N_8994,N_8914);
or U9350 (N_9350,N_9120,N_9144);
nor U9351 (N_9351,N_8806,N_9172);
and U9352 (N_9352,N_9061,N_8949);
and U9353 (N_9353,N_8895,N_9166);
or U9354 (N_9354,N_9174,N_8847);
or U9355 (N_9355,N_9126,N_9180);
and U9356 (N_9356,N_8901,N_9090);
nor U9357 (N_9357,N_9123,N_8882);
or U9358 (N_9358,N_9083,N_8996);
nor U9359 (N_9359,N_8993,N_8892);
and U9360 (N_9360,N_9029,N_8801);
nor U9361 (N_9361,N_9033,N_9006);
nand U9362 (N_9362,N_9127,N_8846);
nand U9363 (N_9363,N_9190,N_9167);
xor U9364 (N_9364,N_9034,N_9171);
and U9365 (N_9365,N_8978,N_8871);
xnor U9366 (N_9366,N_8935,N_9013);
nand U9367 (N_9367,N_9173,N_8951);
and U9368 (N_9368,N_9086,N_8950);
and U9369 (N_9369,N_9040,N_9021);
and U9370 (N_9370,N_9017,N_9064);
and U9371 (N_9371,N_8931,N_9078);
nor U9372 (N_9372,N_8980,N_9106);
and U9373 (N_9373,N_8803,N_8943);
or U9374 (N_9374,N_9163,N_8903);
xnor U9375 (N_9375,N_9129,N_8925);
nor U9376 (N_9376,N_8897,N_9087);
and U9377 (N_9377,N_8810,N_9175);
or U9378 (N_9378,N_9023,N_8905);
nor U9379 (N_9379,N_9016,N_9198);
or U9380 (N_9380,N_9141,N_9103);
nor U9381 (N_9381,N_8868,N_9105);
xor U9382 (N_9382,N_9185,N_8953);
nand U9383 (N_9383,N_9042,N_9045);
and U9384 (N_9384,N_8987,N_8884);
nand U9385 (N_9385,N_8973,N_9095);
nor U9386 (N_9386,N_8815,N_8971);
nand U9387 (N_9387,N_9155,N_8909);
or U9388 (N_9388,N_8926,N_9071);
nor U9389 (N_9389,N_8828,N_9188);
or U9390 (N_9390,N_8833,N_8820);
xor U9391 (N_9391,N_9170,N_8964);
and U9392 (N_9392,N_8929,N_8927);
xnor U9393 (N_9393,N_9183,N_9096);
nand U9394 (N_9394,N_9039,N_8859);
xnor U9395 (N_9395,N_8946,N_8893);
nor U9396 (N_9396,N_8988,N_9136);
and U9397 (N_9397,N_8907,N_9081);
or U9398 (N_9398,N_8862,N_8875);
or U9399 (N_9399,N_9097,N_9137);
and U9400 (N_9400,N_8949,N_9135);
xor U9401 (N_9401,N_9162,N_9158);
and U9402 (N_9402,N_9031,N_8881);
and U9403 (N_9403,N_8920,N_8852);
and U9404 (N_9404,N_8947,N_8976);
and U9405 (N_9405,N_9194,N_9166);
nand U9406 (N_9406,N_8860,N_9086);
or U9407 (N_9407,N_8950,N_8901);
nor U9408 (N_9408,N_8959,N_8827);
nand U9409 (N_9409,N_9012,N_9197);
and U9410 (N_9410,N_8850,N_8834);
xnor U9411 (N_9411,N_8829,N_9104);
and U9412 (N_9412,N_8963,N_8834);
nor U9413 (N_9413,N_8975,N_9002);
nand U9414 (N_9414,N_8985,N_8911);
nand U9415 (N_9415,N_8981,N_9117);
and U9416 (N_9416,N_8803,N_9102);
or U9417 (N_9417,N_8979,N_8807);
nor U9418 (N_9418,N_8889,N_8945);
and U9419 (N_9419,N_9110,N_9033);
xnor U9420 (N_9420,N_8840,N_8959);
nor U9421 (N_9421,N_8825,N_8855);
or U9422 (N_9422,N_8947,N_9045);
nor U9423 (N_9423,N_8884,N_9116);
nand U9424 (N_9424,N_9151,N_8970);
nor U9425 (N_9425,N_9045,N_8948);
and U9426 (N_9426,N_8881,N_9088);
xnor U9427 (N_9427,N_9133,N_8954);
nor U9428 (N_9428,N_9053,N_8817);
and U9429 (N_9429,N_9014,N_9105);
nand U9430 (N_9430,N_8864,N_9059);
and U9431 (N_9431,N_9124,N_8981);
or U9432 (N_9432,N_8995,N_8886);
and U9433 (N_9433,N_9193,N_8876);
nand U9434 (N_9434,N_8967,N_8852);
xor U9435 (N_9435,N_9027,N_8897);
nand U9436 (N_9436,N_9034,N_8833);
or U9437 (N_9437,N_8940,N_9041);
nor U9438 (N_9438,N_9021,N_8950);
xnor U9439 (N_9439,N_9010,N_8969);
or U9440 (N_9440,N_8802,N_9125);
nand U9441 (N_9441,N_8988,N_9181);
nand U9442 (N_9442,N_9120,N_8830);
or U9443 (N_9443,N_9047,N_8985);
nand U9444 (N_9444,N_9065,N_8971);
nor U9445 (N_9445,N_9003,N_9137);
and U9446 (N_9446,N_9001,N_9166);
xor U9447 (N_9447,N_9054,N_9190);
xor U9448 (N_9448,N_8870,N_9026);
or U9449 (N_9449,N_8841,N_8947);
or U9450 (N_9450,N_9131,N_9067);
xor U9451 (N_9451,N_8818,N_8938);
and U9452 (N_9452,N_9016,N_9197);
nand U9453 (N_9453,N_9048,N_9085);
nor U9454 (N_9454,N_9016,N_8994);
and U9455 (N_9455,N_9011,N_9112);
nor U9456 (N_9456,N_9163,N_9174);
nand U9457 (N_9457,N_8987,N_9119);
xnor U9458 (N_9458,N_9010,N_8864);
and U9459 (N_9459,N_8814,N_9130);
and U9460 (N_9460,N_9101,N_9022);
nor U9461 (N_9461,N_8858,N_8830);
nor U9462 (N_9462,N_9037,N_8948);
or U9463 (N_9463,N_8805,N_9164);
or U9464 (N_9464,N_9117,N_9063);
or U9465 (N_9465,N_9006,N_8811);
nor U9466 (N_9466,N_9023,N_9169);
nand U9467 (N_9467,N_8831,N_9059);
nand U9468 (N_9468,N_8926,N_8866);
or U9469 (N_9469,N_8806,N_9063);
or U9470 (N_9470,N_8884,N_9038);
and U9471 (N_9471,N_9012,N_9132);
nand U9472 (N_9472,N_9076,N_9110);
nor U9473 (N_9473,N_9014,N_9145);
xor U9474 (N_9474,N_9085,N_8837);
xnor U9475 (N_9475,N_9060,N_9058);
xor U9476 (N_9476,N_9071,N_9115);
and U9477 (N_9477,N_8889,N_8905);
nand U9478 (N_9478,N_8982,N_8907);
nand U9479 (N_9479,N_9064,N_8921);
nor U9480 (N_9480,N_8876,N_8991);
or U9481 (N_9481,N_9025,N_8865);
and U9482 (N_9482,N_8985,N_8874);
or U9483 (N_9483,N_8956,N_9045);
nand U9484 (N_9484,N_9088,N_9080);
or U9485 (N_9485,N_9165,N_8807);
nand U9486 (N_9486,N_8903,N_8955);
or U9487 (N_9487,N_8905,N_9020);
or U9488 (N_9488,N_9054,N_8831);
nand U9489 (N_9489,N_8883,N_8949);
or U9490 (N_9490,N_9190,N_8800);
xor U9491 (N_9491,N_9087,N_8942);
nand U9492 (N_9492,N_9023,N_8959);
xor U9493 (N_9493,N_8875,N_9178);
nand U9494 (N_9494,N_8870,N_9070);
nor U9495 (N_9495,N_9021,N_9156);
xor U9496 (N_9496,N_9113,N_8802);
xnor U9497 (N_9497,N_8919,N_9147);
xor U9498 (N_9498,N_8908,N_8930);
and U9499 (N_9499,N_9011,N_9158);
nor U9500 (N_9500,N_8992,N_9159);
or U9501 (N_9501,N_8979,N_9057);
nor U9502 (N_9502,N_9117,N_9095);
and U9503 (N_9503,N_8916,N_8865);
xnor U9504 (N_9504,N_8893,N_9003);
or U9505 (N_9505,N_8950,N_9001);
nand U9506 (N_9506,N_9119,N_9190);
nor U9507 (N_9507,N_9079,N_9096);
xnor U9508 (N_9508,N_8977,N_9006);
and U9509 (N_9509,N_9199,N_8841);
nand U9510 (N_9510,N_8961,N_8811);
nand U9511 (N_9511,N_8905,N_9196);
and U9512 (N_9512,N_8855,N_8845);
xnor U9513 (N_9513,N_8898,N_9161);
nand U9514 (N_9514,N_8806,N_9050);
and U9515 (N_9515,N_8949,N_8989);
or U9516 (N_9516,N_9192,N_8959);
nand U9517 (N_9517,N_8866,N_9120);
or U9518 (N_9518,N_9009,N_8965);
xor U9519 (N_9519,N_8832,N_9177);
xor U9520 (N_9520,N_9005,N_8918);
and U9521 (N_9521,N_8861,N_8844);
and U9522 (N_9522,N_9017,N_9050);
nand U9523 (N_9523,N_8842,N_8976);
nor U9524 (N_9524,N_9017,N_9052);
nand U9525 (N_9525,N_9122,N_8894);
nor U9526 (N_9526,N_8816,N_8842);
nor U9527 (N_9527,N_9147,N_8816);
xor U9528 (N_9528,N_8895,N_8997);
nor U9529 (N_9529,N_8839,N_9056);
xnor U9530 (N_9530,N_9051,N_9146);
xor U9531 (N_9531,N_8835,N_8826);
xnor U9532 (N_9532,N_9147,N_9023);
and U9533 (N_9533,N_8970,N_8916);
nand U9534 (N_9534,N_8849,N_9126);
nand U9535 (N_9535,N_9170,N_8843);
and U9536 (N_9536,N_9104,N_8809);
nand U9537 (N_9537,N_8803,N_8880);
and U9538 (N_9538,N_9068,N_9039);
nand U9539 (N_9539,N_9165,N_8894);
xor U9540 (N_9540,N_8947,N_8968);
nand U9541 (N_9541,N_9108,N_9174);
or U9542 (N_9542,N_9000,N_9073);
nand U9543 (N_9543,N_8852,N_9115);
nor U9544 (N_9544,N_9157,N_8834);
xnor U9545 (N_9545,N_9104,N_8921);
or U9546 (N_9546,N_8939,N_8958);
nor U9547 (N_9547,N_9001,N_8978);
or U9548 (N_9548,N_9141,N_9059);
nor U9549 (N_9549,N_9141,N_9161);
nand U9550 (N_9550,N_9160,N_8801);
and U9551 (N_9551,N_9009,N_9120);
and U9552 (N_9552,N_8909,N_8883);
nand U9553 (N_9553,N_8982,N_8994);
nand U9554 (N_9554,N_9195,N_9022);
and U9555 (N_9555,N_9076,N_9125);
nor U9556 (N_9556,N_8981,N_9194);
xnor U9557 (N_9557,N_8931,N_8900);
or U9558 (N_9558,N_9141,N_9124);
xor U9559 (N_9559,N_8893,N_9066);
or U9560 (N_9560,N_8818,N_9041);
nor U9561 (N_9561,N_8994,N_8978);
nor U9562 (N_9562,N_9140,N_8913);
nor U9563 (N_9563,N_8932,N_8820);
nor U9564 (N_9564,N_9137,N_9098);
and U9565 (N_9565,N_9122,N_9124);
xor U9566 (N_9566,N_9136,N_8894);
nor U9567 (N_9567,N_9017,N_9138);
or U9568 (N_9568,N_9066,N_8981);
or U9569 (N_9569,N_9059,N_9170);
nand U9570 (N_9570,N_8856,N_9150);
xor U9571 (N_9571,N_8864,N_9150);
nand U9572 (N_9572,N_9108,N_9093);
xnor U9573 (N_9573,N_8862,N_9124);
xnor U9574 (N_9574,N_8811,N_9171);
and U9575 (N_9575,N_9025,N_9135);
and U9576 (N_9576,N_8998,N_9053);
or U9577 (N_9577,N_8942,N_8953);
xnor U9578 (N_9578,N_8974,N_8891);
nor U9579 (N_9579,N_8919,N_9034);
and U9580 (N_9580,N_8926,N_9066);
or U9581 (N_9581,N_9095,N_9055);
nand U9582 (N_9582,N_9198,N_8990);
and U9583 (N_9583,N_9174,N_9044);
nor U9584 (N_9584,N_8965,N_9111);
nand U9585 (N_9585,N_9129,N_9123);
and U9586 (N_9586,N_9071,N_8971);
or U9587 (N_9587,N_8838,N_9191);
nand U9588 (N_9588,N_8945,N_8877);
xor U9589 (N_9589,N_9000,N_8990);
xor U9590 (N_9590,N_9108,N_8836);
and U9591 (N_9591,N_9079,N_9041);
and U9592 (N_9592,N_8983,N_8856);
and U9593 (N_9593,N_8908,N_8992);
nor U9594 (N_9594,N_8888,N_9088);
or U9595 (N_9595,N_9011,N_8980);
or U9596 (N_9596,N_8967,N_9064);
nor U9597 (N_9597,N_8885,N_9183);
nand U9598 (N_9598,N_9015,N_9073);
nor U9599 (N_9599,N_9108,N_9014);
nor U9600 (N_9600,N_9355,N_9304);
nor U9601 (N_9601,N_9352,N_9565);
or U9602 (N_9602,N_9209,N_9598);
and U9603 (N_9603,N_9523,N_9286);
or U9604 (N_9604,N_9596,N_9587);
nand U9605 (N_9605,N_9445,N_9368);
xnor U9606 (N_9606,N_9345,N_9595);
nand U9607 (N_9607,N_9379,N_9257);
or U9608 (N_9608,N_9211,N_9437);
nor U9609 (N_9609,N_9366,N_9435);
xor U9610 (N_9610,N_9444,N_9513);
xnor U9611 (N_9611,N_9338,N_9436);
and U9612 (N_9612,N_9305,N_9446);
or U9613 (N_9613,N_9458,N_9325);
xor U9614 (N_9614,N_9291,N_9389);
nand U9615 (N_9615,N_9224,N_9205);
nor U9616 (N_9616,N_9510,N_9512);
and U9617 (N_9617,N_9433,N_9397);
nand U9618 (N_9618,N_9400,N_9360);
or U9619 (N_9619,N_9200,N_9482);
xnor U9620 (N_9620,N_9315,N_9295);
xnor U9621 (N_9621,N_9330,N_9550);
xor U9622 (N_9622,N_9216,N_9331);
or U9623 (N_9623,N_9522,N_9532);
nor U9624 (N_9624,N_9229,N_9395);
nor U9625 (N_9625,N_9329,N_9278);
and U9626 (N_9626,N_9254,N_9393);
xnor U9627 (N_9627,N_9577,N_9378);
or U9628 (N_9628,N_9594,N_9206);
xnor U9629 (N_9629,N_9471,N_9493);
or U9630 (N_9630,N_9496,N_9407);
or U9631 (N_9631,N_9293,N_9237);
nand U9632 (N_9632,N_9528,N_9574);
and U9633 (N_9633,N_9374,N_9362);
xnor U9634 (N_9634,N_9571,N_9261);
xor U9635 (N_9635,N_9544,N_9251);
xor U9636 (N_9636,N_9385,N_9466);
nor U9637 (N_9637,N_9258,N_9236);
nand U9638 (N_9638,N_9202,N_9572);
xnor U9639 (N_9639,N_9451,N_9369);
nor U9640 (N_9640,N_9396,N_9506);
nand U9641 (N_9641,N_9307,N_9343);
or U9642 (N_9642,N_9241,N_9204);
xor U9643 (N_9643,N_9421,N_9452);
nor U9644 (N_9644,N_9408,N_9275);
nor U9645 (N_9645,N_9511,N_9464);
and U9646 (N_9646,N_9226,N_9414);
nor U9647 (N_9647,N_9423,N_9288);
or U9648 (N_9648,N_9339,N_9590);
nand U9649 (N_9649,N_9575,N_9539);
nor U9650 (N_9650,N_9592,N_9542);
or U9651 (N_9651,N_9246,N_9581);
or U9652 (N_9652,N_9490,N_9336);
and U9653 (N_9653,N_9322,N_9440);
xor U9654 (N_9654,N_9386,N_9468);
and U9655 (N_9655,N_9530,N_9248);
and U9656 (N_9656,N_9457,N_9504);
or U9657 (N_9657,N_9399,N_9370);
nor U9658 (N_9658,N_9431,N_9289);
and U9659 (N_9659,N_9350,N_9357);
and U9660 (N_9660,N_9524,N_9533);
or U9661 (N_9661,N_9300,N_9459);
or U9662 (N_9662,N_9364,N_9240);
and U9663 (N_9663,N_9526,N_9463);
nor U9664 (N_9664,N_9384,N_9208);
or U9665 (N_9665,N_9551,N_9243);
xnor U9666 (N_9666,N_9447,N_9376);
nor U9667 (N_9667,N_9372,N_9221);
xnor U9668 (N_9668,N_9486,N_9543);
nor U9669 (N_9669,N_9280,N_9439);
nor U9670 (N_9670,N_9567,N_9425);
nor U9671 (N_9671,N_9245,N_9568);
nand U9672 (N_9672,N_9515,N_9277);
and U9673 (N_9673,N_9525,N_9502);
or U9674 (N_9674,N_9273,N_9579);
and U9675 (N_9675,N_9474,N_9531);
or U9676 (N_9676,N_9546,N_9485);
nor U9677 (N_9677,N_9298,N_9207);
nor U9678 (N_9678,N_9538,N_9456);
nor U9679 (N_9679,N_9497,N_9349);
nand U9680 (N_9680,N_9301,N_9472);
xnor U9681 (N_9681,N_9244,N_9235);
nand U9682 (N_9682,N_9255,N_9401);
nor U9683 (N_9683,N_9308,N_9210);
or U9684 (N_9684,N_9488,N_9266);
or U9685 (N_9685,N_9487,N_9317);
nor U9686 (N_9686,N_9358,N_9274);
nand U9687 (N_9687,N_9316,N_9292);
and U9688 (N_9688,N_9230,N_9409);
or U9689 (N_9689,N_9553,N_9453);
xor U9690 (N_9690,N_9501,N_9247);
xnor U9691 (N_9691,N_9265,N_9503);
xor U9692 (N_9692,N_9563,N_9227);
nor U9693 (N_9693,N_9371,N_9297);
or U9694 (N_9694,N_9483,N_9271);
or U9695 (N_9695,N_9570,N_9561);
xor U9696 (N_9696,N_9517,N_9420);
xor U9697 (N_9697,N_9249,N_9489);
nand U9698 (N_9698,N_9537,N_9259);
and U9699 (N_9699,N_9333,N_9545);
or U9700 (N_9700,N_9494,N_9593);
xnor U9701 (N_9701,N_9250,N_9541);
nor U9702 (N_9702,N_9552,N_9521);
or U9703 (N_9703,N_9467,N_9282);
or U9704 (N_9704,N_9377,N_9225);
xnor U9705 (N_9705,N_9335,N_9302);
nand U9706 (N_9706,N_9529,N_9536);
nand U9707 (N_9707,N_9215,N_9281);
and U9708 (N_9708,N_9426,N_9262);
xnor U9709 (N_9709,N_9564,N_9448);
nor U9710 (N_9710,N_9213,N_9422);
nor U9711 (N_9711,N_9242,N_9394);
nor U9712 (N_9712,N_9231,N_9573);
xnor U9713 (N_9713,N_9558,N_9268);
and U9714 (N_9714,N_9388,N_9450);
nand U9715 (N_9715,N_9212,N_9228);
xor U9716 (N_9716,N_9264,N_9356);
and U9717 (N_9717,N_9419,N_9363);
nor U9718 (N_9718,N_9219,N_9365);
or U9719 (N_9719,N_9578,N_9582);
nand U9720 (N_9720,N_9585,N_9500);
nand U9721 (N_9721,N_9424,N_9406);
nand U9722 (N_9722,N_9346,N_9432);
nor U9723 (N_9723,N_9566,N_9354);
or U9724 (N_9724,N_9320,N_9465);
nor U9725 (N_9725,N_9238,N_9390);
xor U9726 (N_9726,N_9287,N_9548);
and U9727 (N_9727,N_9481,N_9284);
nor U9728 (N_9728,N_9410,N_9359);
nand U9729 (N_9729,N_9233,N_9392);
xor U9730 (N_9730,N_9491,N_9220);
nand U9731 (N_9731,N_9344,N_9239);
nor U9732 (N_9732,N_9516,N_9584);
xor U9733 (N_9733,N_9222,N_9441);
xor U9734 (N_9734,N_9310,N_9480);
xnor U9735 (N_9735,N_9381,N_9256);
nor U9736 (N_9736,N_9234,N_9417);
nor U9737 (N_9737,N_9427,N_9518);
or U9738 (N_9738,N_9527,N_9323);
and U9739 (N_9739,N_9294,N_9442);
or U9740 (N_9740,N_9554,N_9462);
xor U9741 (N_9741,N_9285,N_9398);
or U9742 (N_9742,N_9473,N_9520);
xnor U9743 (N_9743,N_9404,N_9560);
nand U9744 (N_9744,N_9270,N_9290);
nand U9745 (N_9745,N_9597,N_9557);
xor U9746 (N_9746,N_9555,N_9413);
xnor U9747 (N_9747,N_9469,N_9498);
and U9748 (N_9748,N_9319,N_9253);
xnor U9749 (N_9749,N_9547,N_9387);
xor U9750 (N_9750,N_9283,N_9492);
nor U9751 (N_9751,N_9223,N_9430);
and U9752 (N_9752,N_9303,N_9509);
nor U9753 (N_9753,N_9382,N_9272);
xor U9754 (N_9754,N_9267,N_9218);
nand U9755 (N_9755,N_9334,N_9296);
nand U9756 (N_9756,N_9321,N_9309);
nor U9757 (N_9757,N_9434,N_9332);
nand U9758 (N_9758,N_9449,N_9351);
xor U9759 (N_9759,N_9232,N_9591);
nor U9760 (N_9760,N_9562,N_9324);
nor U9761 (N_9761,N_9475,N_9438);
or U9762 (N_9762,N_9540,N_9361);
nand U9763 (N_9763,N_9380,N_9580);
xnor U9764 (N_9764,N_9589,N_9314);
nand U9765 (N_9765,N_9263,N_9318);
nor U9766 (N_9766,N_9416,N_9383);
nand U9767 (N_9767,N_9507,N_9535);
xor U9768 (N_9768,N_9429,N_9375);
nand U9769 (N_9769,N_9299,N_9412);
or U9770 (N_9770,N_9478,N_9326);
nand U9771 (N_9771,N_9411,N_9279);
and U9772 (N_9772,N_9328,N_9477);
or U9773 (N_9773,N_9269,N_9549);
nor U9774 (N_9774,N_9534,N_9476);
xor U9775 (N_9775,N_9313,N_9599);
or U9776 (N_9776,N_9217,N_9252);
nor U9777 (N_9777,N_9327,N_9418);
and U9778 (N_9778,N_9454,N_9402);
nand U9779 (N_9779,N_9260,N_9337);
nand U9780 (N_9780,N_9455,N_9484);
and U9781 (N_9781,N_9519,N_9470);
nand U9782 (N_9782,N_9556,N_9348);
nand U9783 (N_9783,N_9576,N_9559);
xor U9784 (N_9784,N_9569,N_9583);
xor U9785 (N_9785,N_9312,N_9508);
nor U9786 (N_9786,N_9588,N_9391);
nand U9787 (N_9787,N_9342,N_9214);
xnor U9788 (N_9788,N_9373,N_9461);
nor U9789 (N_9789,N_9367,N_9347);
nand U9790 (N_9790,N_9479,N_9340);
nor U9791 (N_9791,N_9201,N_9276);
nor U9792 (N_9792,N_9203,N_9428);
or U9793 (N_9793,N_9353,N_9499);
and U9794 (N_9794,N_9415,N_9403);
nor U9795 (N_9795,N_9505,N_9460);
nand U9796 (N_9796,N_9306,N_9311);
nor U9797 (N_9797,N_9586,N_9341);
xnor U9798 (N_9798,N_9443,N_9514);
nand U9799 (N_9799,N_9495,N_9405);
or U9800 (N_9800,N_9202,N_9430);
nand U9801 (N_9801,N_9389,N_9497);
xnor U9802 (N_9802,N_9443,N_9240);
nand U9803 (N_9803,N_9238,N_9281);
and U9804 (N_9804,N_9522,N_9331);
nand U9805 (N_9805,N_9284,N_9365);
nor U9806 (N_9806,N_9241,N_9495);
and U9807 (N_9807,N_9277,N_9472);
nor U9808 (N_9808,N_9506,N_9239);
and U9809 (N_9809,N_9345,N_9295);
xor U9810 (N_9810,N_9488,N_9249);
and U9811 (N_9811,N_9292,N_9537);
nand U9812 (N_9812,N_9323,N_9461);
nand U9813 (N_9813,N_9386,N_9509);
or U9814 (N_9814,N_9532,N_9204);
or U9815 (N_9815,N_9384,N_9447);
or U9816 (N_9816,N_9304,N_9483);
xor U9817 (N_9817,N_9209,N_9336);
or U9818 (N_9818,N_9312,N_9559);
and U9819 (N_9819,N_9587,N_9544);
or U9820 (N_9820,N_9435,N_9411);
and U9821 (N_9821,N_9290,N_9446);
nand U9822 (N_9822,N_9200,N_9556);
xor U9823 (N_9823,N_9365,N_9345);
or U9824 (N_9824,N_9413,N_9521);
nor U9825 (N_9825,N_9449,N_9395);
nand U9826 (N_9826,N_9493,N_9441);
xor U9827 (N_9827,N_9285,N_9452);
xor U9828 (N_9828,N_9268,N_9346);
and U9829 (N_9829,N_9520,N_9206);
or U9830 (N_9830,N_9263,N_9569);
xnor U9831 (N_9831,N_9507,N_9553);
nor U9832 (N_9832,N_9278,N_9342);
xor U9833 (N_9833,N_9299,N_9362);
nand U9834 (N_9834,N_9219,N_9596);
or U9835 (N_9835,N_9471,N_9291);
nand U9836 (N_9836,N_9220,N_9597);
nor U9837 (N_9837,N_9575,N_9415);
nand U9838 (N_9838,N_9495,N_9343);
nand U9839 (N_9839,N_9427,N_9339);
or U9840 (N_9840,N_9485,N_9308);
nand U9841 (N_9841,N_9475,N_9342);
and U9842 (N_9842,N_9373,N_9387);
and U9843 (N_9843,N_9398,N_9554);
and U9844 (N_9844,N_9242,N_9237);
and U9845 (N_9845,N_9482,N_9260);
xnor U9846 (N_9846,N_9425,N_9478);
nand U9847 (N_9847,N_9302,N_9483);
xnor U9848 (N_9848,N_9218,N_9312);
and U9849 (N_9849,N_9434,N_9562);
nor U9850 (N_9850,N_9501,N_9230);
xor U9851 (N_9851,N_9279,N_9383);
nor U9852 (N_9852,N_9539,N_9318);
nand U9853 (N_9853,N_9369,N_9394);
or U9854 (N_9854,N_9327,N_9288);
nand U9855 (N_9855,N_9416,N_9329);
nor U9856 (N_9856,N_9551,N_9541);
xnor U9857 (N_9857,N_9215,N_9315);
xnor U9858 (N_9858,N_9246,N_9525);
and U9859 (N_9859,N_9501,N_9323);
nor U9860 (N_9860,N_9310,N_9309);
nor U9861 (N_9861,N_9236,N_9326);
or U9862 (N_9862,N_9246,N_9527);
or U9863 (N_9863,N_9308,N_9331);
nand U9864 (N_9864,N_9310,N_9449);
xnor U9865 (N_9865,N_9473,N_9572);
nor U9866 (N_9866,N_9361,N_9565);
and U9867 (N_9867,N_9272,N_9434);
nand U9868 (N_9868,N_9388,N_9547);
nor U9869 (N_9869,N_9406,N_9540);
and U9870 (N_9870,N_9352,N_9258);
or U9871 (N_9871,N_9401,N_9596);
and U9872 (N_9872,N_9206,N_9473);
and U9873 (N_9873,N_9514,N_9263);
or U9874 (N_9874,N_9269,N_9322);
and U9875 (N_9875,N_9205,N_9299);
or U9876 (N_9876,N_9540,N_9437);
nor U9877 (N_9877,N_9270,N_9323);
nor U9878 (N_9878,N_9319,N_9303);
nand U9879 (N_9879,N_9535,N_9377);
nand U9880 (N_9880,N_9596,N_9304);
and U9881 (N_9881,N_9514,N_9372);
nand U9882 (N_9882,N_9273,N_9462);
nand U9883 (N_9883,N_9545,N_9378);
or U9884 (N_9884,N_9411,N_9200);
nor U9885 (N_9885,N_9403,N_9269);
and U9886 (N_9886,N_9326,N_9536);
nor U9887 (N_9887,N_9294,N_9208);
nand U9888 (N_9888,N_9332,N_9349);
nand U9889 (N_9889,N_9338,N_9209);
nand U9890 (N_9890,N_9543,N_9460);
and U9891 (N_9891,N_9309,N_9404);
or U9892 (N_9892,N_9347,N_9467);
or U9893 (N_9893,N_9583,N_9314);
nand U9894 (N_9894,N_9392,N_9485);
nand U9895 (N_9895,N_9352,N_9404);
and U9896 (N_9896,N_9289,N_9248);
nand U9897 (N_9897,N_9492,N_9211);
nor U9898 (N_9898,N_9583,N_9471);
and U9899 (N_9899,N_9229,N_9488);
nor U9900 (N_9900,N_9309,N_9246);
or U9901 (N_9901,N_9312,N_9305);
and U9902 (N_9902,N_9230,N_9485);
nor U9903 (N_9903,N_9551,N_9437);
xnor U9904 (N_9904,N_9366,N_9229);
or U9905 (N_9905,N_9473,N_9274);
and U9906 (N_9906,N_9510,N_9421);
nand U9907 (N_9907,N_9349,N_9445);
nor U9908 (N_9908,N_9467,N_9492);
xnor U9909 (N_9909,N_9261,N_9468);
nand U9910 (N_9910,N_9482,N_9465);
or U9911 (N_9911,N_9496,N_9239);
xnor U9912 (N_9912,N_9219,N_9301);
and U9913 (N_9913,N_9337,N_9367);
xor U9914 (N_9914,N_9281,N_9269);
or U9915 (N_9915,N_9485,N_9437);
nand U9916 (N_9916,N_9512,N_9355);
nor U9917 (N_9917,N_9300,N_9228);
and U9918 (N_9918,N_9480,N_9481);
or U9919 (N_9919,N_9432,N_9216);
xor U9920 (N_9920,N_9584,N_9358);
nor U9921 (N_9921,N_9591,N_9554);
nor U9922 (N_9922,N_9481,N_9587);
nor U9923 (N_9923,N_9307,N_9553);
nor U9924 (N_9924,N_9227,N_9347);
nand U9925 (N_9925,N_9410,N_9578);
nor U9926 (N_9926,N_9239,N_9203);
nand U9927 (N_9927,N_9428,N_9340);
nor U9928 (N_9928,N_9417,N_9565);
nand U9929 (N_9929,N_9268,N_9361);
nand U9930 (N_9930,N_9564,N_9325);
nor U9931 (N_9931,N_9579,N_9234);
xnor U9932 (N_9932,N_9253,N_9358);
xnor U9933 (N_9933,N_9449,N_9492);
or U9934 (N_9934,N_9569,N_9407);
or U9935 (N_9935,N_9598,N_9321);
or U9936 (N_9936,N_9397,N_9287);
xnor U9937 (N_9937,N_9582,N_9224);
or U9938 (N_9938,N_9505,N_9538);
and U9939 (N_9939,N_9385,N_9391);
xnor U9940 (N_9940,N_9341,N_9485);
nor U9941 (N_9941,N_9587,N_9343);
nand U9942 (N_9942,N_9592,N_9486);
or U9943 (N_9943,N_9412,N_9356);
nand U9944 (N_9944,N_9526,N_9296);
or U9945 (N_9945,N_9461,N_9226);
nand U9946 (N_9946,N_9213,N_9290);
nor U9947 (N_9947,N_9468,N_9599);
and U9948 (N_9948,N_9413,N_9320);
and U9949 (N_9949,N_9381,N_9557);
or U9950 (N_9950,N_9568,N_9399);
or U9951 (N_9951,N_9201,N_9316);
nor U9952 (N_9952,N_9508,N_9465);
and U9953 (N_9953,N_9325,N_9570);
nand U9954 (N_9954,N_9271,N_9512);
xor U9955 (N_9955,N_9552,N_9536);
xnor U9956 (N_9956,N_9272,N_9360);
nand U9957 (N_9957,N_9272,N_9423);
and U9958 (N_9958,N_9327,N_9438);
nor U9959 (N_9959,N_9498,N_9217);
or U9960 (N_9960,N_9453,N_9295);
nand U9961 (N_9961,N_9211,N_9267);
nor U9962 (N_9962,N_9211,N_9330);
and U9963 (N_9963,N_9452,N_9471);
or U9964 (N_9964,N_9419,N_9273);
xor U9965 (N_9965,N_9238,N_9318);
or U9966 (N_9966,N_9561,N_9294);
or U9967 (N_9967,N_9448,N_9245);
nand U9968 (N_9968,N_9372,N_9237);
nand U9969 (N_9969,N_9341,N_9369);
nand U9970 (N_9970,N_9220,N_9293);
xnor U9971 (N_9971,N_9350,N_9540);
nor U9972 (N_9972,N_9451,N_9228);
nor U9973 (N_9973,N_9497,N_9462);
xor U9974 (N_9974,N_9594,N_9409);
xnor U9975 (N_9975,N_9296,N_9454);
xnor U9976 (N_9976,N_9254,N_9564);
xnor U9977 (N_9977,N_9319,N_9501);
nand U9978 (N_9978,N_9236,N_9265);
xnor U9979 (N_9979,N_9432,N_9428);
or U9980 (N_9980,N_9258,N_9280);
xor U9981 (N_9981,N_9222,N_9231);
nor U9982 (N_9982,N_9245,N_9589);
nor U9983 (N_9983,N_9531,N_9239);
nand U9984 (N_9984,N_9354,N_9416);
nor U9985 (N_9985,N_9495,N_9504);
nor U9986 (N_9986,N_9566,N_9234);
nor U9987 (N_9987,N_9307,N_9557);
or U9988 (N_9988,N_9290,N_9215);
and U9989 (N_9989,N_9418,N_9453);
and U9990 (N_9990,N_9492,N_9541);
nor U9991 (N_9991,N_9215,N_9252);
nor U9992 (N_9992,N_9539,N_9541);
and U9993 (N_9993,N_9320,N_9403);
nand U9994 (N_9994,N_9269,N_9406);
xnor U9995 (N_9995,N_9571,N_9551);
xnor U9996 (N_9996,N_9381,N_9460);
nor U9997 (N_9997,N_9372,N_9347);
nand U9998 (N_9998,N_9356,N_9500);
or U9999 (N_9999,N_9599,N_9328);
xnor U10000 (N_10000,N_9658,N_9922);
and U10001 (N_10001,N_9877,N_9974);
nor U10002 (N_10002,N_9622,N_9775);
xnor U10003 (N_10003,N_9838,N_9923);
nor U10004 (N_10004,N_9740,N_9819);
and U10005 (N_10005,N_9713,N_9681);
nor U10006 (N_10006,N_9771,N_9892);
xor U10007 (N_10007,N_9600,N_9940);
nand U10008 (N_10008,N_9620,N_9730);
and U10009 (N_10009,N_9711,N_9635);
or U10010 (N_10010,N_9610,N_9844);
xor U10011 (N_10011,N_9677,N_9686);
and U10012 (N_10012,N_9993,N_9723);
xor U10013 (N_10013,N_9830,N_9800);
nor U10014 (N_10014,N_9815,N_9864);
or U10015 (N_10015,N_9665,N_9774);
or U10016 (N_10016,N_9908,N_9631);
and U10017 (N_10017,N_9884,N_9885);
and U10018 (N_10018,N_9925,N_9679);
nor U10019 (N_10019,N_9987,N_9700);
or U10020 (N_10020,N_9789,N_9797);
nor U10021 (N_10021,N_9847,N_9882);
nor U10022 (N_10022,N_9707,N_9902);
nand U10023 (N_10023,N_9957,N_9672);
nand U10024 (N_10024,N_9655,N_9788);
nor U10025 (N_10025,N_9968,N_9924);
nand U10026 (N_10026,N_9701,N_9613);
xnor U10027 (N_10027,N_9856,N_9778);
and U10028 (N_10028,N_9917,N_9971);
and U10029 (N_10029,N_9854,N_9979);
nand U10030 (N_10030,N_9870,N_9629);
nor U10031 (N_10031,N_9688,N_9717);
or U10032 (N_10032,N_9732,N_9961);
nand U10033 (N_10033,N_9805,N_9669);
nand U10034 (N_10034,N_9855,N_9947);
nand U10035 (N_10035,N_9764,N_9733);
xnor U10036 (N_10036,N_9958,N_9822);
and U10037 (N_10037,N_9663,N_9779);
or U10038 (N_10038,N_9801,N_9934);
xor U10039 (N_10039,N_9953,N_9683);
nand U10040 (N_10040,N_9682,N_9921);
or U10041 (N_10041,N_9736,N_9799);
and U10042 (N_10042,N_9770,N_9706);
nand U10043 (N_10043,N_9816,N_9731);
xnor U10044 (N_10044,N_9914,N_9916);
xor U10045 (N_10045,N_9603,N_9929);
nor U10046 (N_10046,N_9959,N_9840);
nor U10047 (N_10047,N_9752,N_9963);
and U10048 (N_10048,N_9633,N_9738);
nor U10049 (N_10049,N_9932,N_9605);
and U10050 (N_10050,N_9754,N_9980);
or U10051 (N_10051,N_9909,N_9767);
or U10052 (N_10052,N_9760,N_9915);
or U10053 (N_10053,N_9810,N_9868);
or U10054 (N_10054,N_9858,N_9790);
nor U10055 (N_10055,N_9849,N_9966);
nand U10056 (N_10056,N_9865,N_9803);
or U10057 (N_10057,N_9699,N_9689);
nor U10058 (N_10058,N_9920,N_9601);
or U10059 (N_10059,N_9741,N_9626);
nor U10060 (N_10060,N_9606,N_9793);
nand U10061 (N_10061,N_9883,N_9956);
and U10062 (N_10062,N_9808,N_9937);
and U10063 (N_10063,N_9895,N_9654);
xnor U10064 (N_10064,N_9604,N_9728);
xnor U10065 (N_10065,N_9724,N_9725);
nor U10066 (N_10066,N_9964,N_9696);
nand U10067 (N_10067,N_9852,N_9656);
nand U10068 (N_10068,N_9969,N_9662);
nand U10069 (N_10069,N_9640,N_9893);
and U10070 (N_10070,N_9933,N_9988);
and U10071 (N_10071,N_9863,N_9650);
or U10072 (N_10072,N_9862,N_9950);
nor U10073 (N_10073,N_9763,N_9729);
nand U10074 (N_10074,N_9755,N_9753);
or U10075 (N_10075,N_9829,N_9674);
nor U10076 (N_10076,N_9942,N_9714);
and U10077 (N_10077,N_9873,N_9625);
or U10078 (N_10078,N_9690,N_9794);
nand U10079 (N_10079,N_9667,N_9802);
or U10080 (N_10080,N_9617,N_9871);
nand U10081 (N_10081,N_9692,N_9630);
or U10082 (N_10082,N_9765,N_9996);
xor U10083 (N_10083,N_9680,N_9685);
and U10084 (N_10084,N_9670,N_9879);
nor U10085 (N_10085,N_9842,N_9967);
nor U10086 (N_10086,N_9716,N_9911);
nor U10087 (N_10087,N_9703,N_9995);
nand U10088 (N_10088,N_9839,N_9621);
xnor U10089 (N_10089,N_9935,N_9825);
or U10090 (N_10090,N_9850,N_9919);
xor U10091 (N_10091,N_9787,N_9983);
and U10092 (N_10092,N_9820,N_9989);
nand U10093 (N_10093,N_9901,N_9756);
or U10094 (N_10094,N_9647,N_9811);
nand U10095 (N_10095,N_9960,N_9894);
or U10096 (N_10096,N_9627,N_9824);
xnor U10097 (N_10097,N_9628,N_9876);
and U10098 (N_10098,N_9990,N_9936);
nand U10099 (N_10099,N_9722,N_9719);
or U10100 (N_10100,N_9757,N_9768);
nand U10101 (N_10101,N_9761,N_9708);
and U10102 (N_10102,N_9737,N_9782);
and U10103 (N_10103,N_9720,N_9972);
nor U10104 (N_10104,N_9931,N_9661);
or U10105 (N_10105,N_9821,N_9702);
xor U10106 (N_10106,N_9848,N_9780);
nor U10107 (N_10107,N_9886,N_9607);
nand U10108 (N_10108,N_9875,N_9938);
and U10109 (N_10109,N_9860,N_9785);
or U10110 (N_10110,N_9612,N_9673);
nor U10111 (N_10111,N_9747,N_9618);
xnor U10112 (N_10112,N_9712,N_9837);
and U10113 (N_10113,N_9889,N_9927);
or U10114 (N_10114,N_9982,N_9671);
nor U10115 (N_10115,N_9851,N_9695);
nand U10116 (N_10116,N_9833,N_9639);
and U10117 (N_10117,N_9866,N_9634);
or U10118 (N_10118,N_9910,N_9898);
nand U10119 (N_10119,N_9726,N_9943);
xor U10120 (N_10120,N_9999,N_9691);
nor U10121 (N_10121,N_9985,N_9945);
and U10122 (N_10122,N_9928,N_9951);
and U10123 (N_10123,N_9687,N_9704);
and U10124 (N_10124,N_9872,N_9705);
xor U10125 (N_10125,N_9795,N_9721);
xnor U10126 (N_10126,N_9874,N_9666);
or U10127 (N_10127,N_9694,N_9739);
nor U10128 (N_10128,N_9818,N_9745);
xor U10129 (N_10129,N_9759,N_9727);
and U10130 (N_10130,N_9975,N_9749);
nor U10131 (N_10131,N_9913,N_9867);
nand U10132 (N_10132,N_9616,N_9637);
and U10133 (N_10133,N_9984,N_9792);
nand U10134 (N_10134,N_9698,N_9976);
nand U10135 (N_10135,N_9978,N_9676);
or U10136 (N_10136,N_9948,N_9977);
xnor U10137 (N_10137,N_9715,N_9807);
nand U10138 (N_10138,N_9817,N_9773);
and U10139 (N_10139,N_9939,N_9880);
or U10140 (N_10140,N_9997,N_9904);
and U10141 (N_10141,N_9742,N_9944);
or U10142 (N_10142,N_9841,N_9831);
nor U10143 (N_10143,N_9697,N_9709);
nor U10144 (N_10144,N_9602,N_9784);
or U10145 (N_10145,N_9887,N_9614);
or U10146 (N_10146,N_9869,N_9734);
nor U10147 (N_10147,N_9965,N_9632);
nand U10148 (N_10148,N_9828,N_9918);
or U10149 (N_10149,N_9970,N_9891);
and U10150 (N_10150,N_9623,N_9641);
and U10151 (N_10151,N_9660,N_9861);
nand U10152 (N_10152,N_9651,N_9798);
nor U10153 (N_10153,N_9907,N_9645);
nand U10154 (N_10154,N_9718,N_9648);
nor U10155 (N_10155,N_9710,N_9649);
xnor U10156 (N_10156,N_9735,N_9777);
and U10157 (N_10157,N_9846,N_9878);
or U10158 (N_10158,N_9845,N_9653);
and U10159 (N_10159,N_9812,N_9624);
or U10160 (N_10160,N_9832,N_9946);
xnor U10161 (N_10161,N_9952,N_9748);
xnor U10162 (N_10162,N_9991,N_9643);
nand U10163 (N_10163,N_9834,N_9664);
and U10164 (N_10164,N_9659,N_9758);
and U10165 (N_10165,N_9684,N_9783);
and U10166 (N_10166,N_9857,N_9890);
nand U10167 (N_10167,N_9744,N_9804);
nand U10168 (N_10168,N_9823,N_9678);
or U10169 (N_10169,N_9992,N_9646);
nand U10170 (N_10170,N_9611,N_9642);
or U10171 (N_10171,N_9608,N_9781);
nand U10172 (N_10172,N_9644,N_9981);
or U10173 (N_10173,N_9994,N_9881);
nor U10174 (N_10174,N_9668,N_9652);
nor U10175 (N_10175,N_9843,N_9796);
and U10176 (N_10176,N_9638,N_9809);
and U10177 (N_10177,N_9973,N_9806);
xor U10178 (N_10178,N_9905,N_9930);
nand U10179 (N_10179,N_9998,N_9888);
and U10180 (N_10180,N_9609,N_9750);
nor U10181 (N_10181,N_9772,N_9903);
or U10182 (N_10182,N_9693,N_9813);
nor U10183 (N_10183,N_9826,N_9743);
xor U10184 (N_10184,N_9751,N_9859);
or U10185 (N_10185,N_9776,N_9900);
xnor U10186 (N_10186,N_9675,N_9941);
nand U10187 (N_10187,N_9912,N_9955);
xor U10188 (N_10188,N_9896,N_9853);
nand U10189 (N_10189,N_9786,N_9986);
or U10190 (N_10190,N_9746,N_9762);
nand U10191 (N_10191,N_9791,N_9906);
nor U10192 (N_10192,N_9836,N_9766);
or U10193 (N_10193,N_9615,N_9949);
nor U10194 (N_10194,N_9619,N_9814);
xnor U10195 (N_10195,N_9954,N_9962);
nand U10196 (N_10196,N_9827,N_9835);
nor U10197 (N_10197,N_9926,N_9657);
nand U10198 (N_10198,N_9899,N_9636);
nor U10199 (N_10199,N_9897,N_9769);
and U10200 (N_10200,N_9649,N_9822);
or U10201 (N_10201,N_9714,N_9621);
nand U10202 (N_10202,N_9625,N_9842);
nor U10203 (N_10203,N_9998,N_9933);
xnor U10204 (N_10204,N_9845,N_9702);
nand U10205 (N_10205,N_9681,N_9696);
or U10206 (N_10206,N_9991,N_9908);
or U10207 (N_10207,N_9799,N_9820);
or U10208 (N_10208,N_9811,N_9908);
xor U10209 (N_10209,N_9685,N_9973);
nor U10210 (N_10210,N_9931,N_9840);
and U10211 (N_10211,N_9840,N_9982);
xnor U10212 (N_10212,N_9601,N_9871);
or U10213 (N_10213,N_9975,N_9977);
nor U10214 (N_10214,N_9783,N_9952);
nor U10215 (N_10215,N_9966,N_9610);
nor U10216 (N_10216,N_9639,N_9736);
nor U10217 (N_10217,N_9895,N_9617);
nand U10218 (N_10218,N_9733,N_9709);
xnor U10219 (N_10219,N_9868,N_9653);
or U10220 (N_10220,N_9948,N_9886);
and U10221 (N_10221,N_9784,N_9614);
or U10222 (N_10222,N_9667,N_9876);
nand U10223 (N_10223,N_9964,N_9993);
or U10224 (N_10224,N_9853,N_9646);
and U10225 (N_10225,N_9656,N_9611);
nor U10226 (N_10226,N_9630,N_9783);
nor U10227 (N_10227,N_9742,N_9603);
and U10228 (N_10228,N_9825,N_9700);
and U10229 (N_10229,N_9703,N_9958);
nor U10230 (N_10230,N_9976,N_9830);
nor U10231 (N_10231,N_9656,N_9693);
xor U10232 (N_10232,N_9859,N_9680);
or U10233 (N_10233,N_9988,N_9952);
xnor U10234 (N_10234,N_9739,N_9730);
nand U10235 (N_10235,N_9830,N_9741);
and U10236 (N_10236,N_9699,N_9686);
and U10237 (N_10237,N_9991,N_9896);
or U10238 (N_10238,N_9756,N_9728);
nand U10239 (N_10239,N_9863,N_9961);
or U10240 (N_10240,N_9797,N_9615);
nor U10241 (N_10241,N_9711,N_9883);
xnor U10242 (N_10242,N_9761,N_9829);
xnor U10243 (N_10243,N_9880,N_9787);
and U10244 (N_10244,N_9642,N_9873);
nand U10245 (N_10245,N_9840,N_9603);
nor U10246 (N_10246,N_9900,N_9848);
nor U10247 (N_10247,N_9895,N_9708);
nand U10248 (N_10248,N_9608,N_9685);
xnor U10249 (N_10249,N_9929,N_9881);
nand U10250 (N_10250,N_9785,N_9859);
and U10251 (N_10251,N_9922,N_9641);
nand U10252 (N_10252,N_9867,N_9627);
or U10253 (N_10253,N_9720,N_9954);
or U10254 (N_10254,N_9783,N_9915);
xnor U10255 (N_10255,N_9751,N_9683);
nor U10256 (N_10256,N_9952,N_9853);
xnor U10257 (N_10257,N_9621,N_9977);
nand U10258 (N_10258,N_9658,N_9710);
and U10259 (N_10259,N_9707,N_9864);
or U10260 (N_10260,N_9956,N_9822);
xor U10261 (N_10261,N_9966,N_9799);
xor U10262 (N_10262,N_9688,N_9660);
or U10263 (N_10263,N_9906,N_9822);
xor U10264 (N_10264,N_9969,N_9977);
nor U10265 (N_10265,N_9835,N_9660);
or U10266 (N_10266,N_9852,N_9904);
xnor U10267 (N_10267,N_9811,N_9936);
xor U10268 (N_10268,N_9987,N_9991);
and U10269 (N_10269,N_9668,N_9735);
or U10270 (N_10270,N_9767,N_9856);
and U10271 (N_10271,N_9651,N_9641);
xor U10272 (N_10272,N_9893,N_9657);
and U10273 (N_10273,N_9838,N_9666);
and U10274 (N_10274,N_9812,N_9620);
or U10275 (N_10275,N_9925,N_9675);
nor U10276 (N_10276,N_9825,N_9828);
nor U10277 (N_10277,N_9783,N_9835);
nor U10278 (N_10278,N_9690,N_9716);
nor U10279 (N_10279,N_9740,N_9639);
or U10280 (N_10280,N_9629,N_9682);
xor U10281 (N_10281,N_9931,N_9837);
xnor U10282 (N_10282,N_9900,N_9915);
nand U10283 (N_10283,N_9833,N_9847);
xnor U10284 (N_10284,N_9995,N_9653);
and U10285 (N_10285,N_9763,N_9970);
nor U10286 (N_10286,N_9703,N_9627);
xor U10287 (N_10287,N_9769,N_9737);
and U10288 (N_10288,N_9764,N_9984);
xnor U10289 (N_10289,N_9964,N_9856);
and U10290 (N_10290,N_9847,N_9642);
or U10291 (N_10291,N_9884,N_9632);
or U10292 (N_10292,N_9738,N_9926);
and U10293 (N_10293,N_9815,N_9924);
xor U10294 (N_10294,N_9786,N_9766);
nor U10295 (N_10295,N_9776,N_9816);
nand U10296 (N_10296,N_9735,N_9966);
xnor U10297 (N_10297,N_9756,N_9631);
or U10298 (N_10298,N_9657,N_9976);
or U10299 (N_10299,N_9863,N_9923);
xnor U10300 (N_10300,N_9613,N_9944);
nor U10301 (N_10301,N_9954,N_9788);
or U10302 (N_10302,N_9809,N_9991);
xnor U10303 (N_10303,N_9646,N_9960);
nor U10304 (N_10304,N_9729,N_9926);
xnor U10305 (N_10305,N_9665,N_9879);
or U10306 (N_10306,N_9850,N_9873);
or U10307 (N_10307,N_9998,N_9697);
or U10308 (N_10308,N_9936,N_9601);
nand U10309 (N_10309,N_9671,N_9610);
nand U10310 (N_10310,N_9778,N_9997);
xor U10311 (N_10311,N_9959,N_9709);
and U10312 (N_10312,N_9903,N_9927);
nand U10313 (N_10313,N_9755,N_9729);
nand U10314 (N_10314,N_9605,N_9744);
nand U10315 (N_10315,N_9774,N_9663);
xnor U10316 (N_10316,N_9690,N_9800);
and U10317 (N_10317,N_9818,N_9837);
nor U10318 (N_10318,N_9710,N_9703);
and U10319 (N_10319,N_9889,N_9968);
or U10320 (N_10320,N_9704,N_9937);
or U10321 (N_10321,N_9724,N_9772);
nand U10322 (N_10322,N_9966,N_9770);
nor U10323 (N_10323,N_9966,N_9857);
xnor U10324 (N_10324,N_9670,N_9967);
and U10325 (N_10325,N_9984,N_9755);
nand U10326 (N_10326,N_9859,N_9691);
xor U10327 (N_10327,N_9749,N_9669);
and U10328 (N_10328,N_9609,N_9616);
nor U10329 (N_10329,N_9648,N_9692);
or U10330 (N_10330,N_9978,N_9893);
or U10331 (N_10331,N_9818,N_9936);
xor U10332 (N_10332,N_9740,N_9753);
or U10333 (N_10333,N_9668,N_9971);
nor U10334 (N_10334,N_9689,N_9807);
nand U10335 (N_10335,N_9919,N_9897);
nand U10336 (N_10336,N_9767,N_9838);
nor U10337 (N_10337,N_9931,N_9639);
or U10338 (N_10338,N_9667,N_9611);
or U10339 (N_10339,N_9890,N_9928);
nand U10340 (N_10340,N_9953,N_9654);
xnor U10341 (N_10341,N_9876,N_9715);
nor U10342 (N_10342,N_9901,N_9714);
nor U10343 (N_10343,N_9677,N_9960);
and U10344 (N_10344,N_9723,N_9641);
nor U10345 (N_10345,N_9847,N_9678);
nor U10346 (N_10346,N_9956,N_9809);
xnor U10347 (N_10347,N_9938,N_9743);
nand U10348 (N_10348,N_9955,N_9977);
nand U10349 (N_10349,N_9940,N_9735);
and U10350 (N_10350,N_9676,N_9785);
nor U10351 (N_10351,N_9874,N_9832);
or U10352 (N_10352,N_9763,N_9633);
nor U10353 (N_10353,N_9684,N_9661);
and U10354 (N_10354,N_9922,N_9815);
xor U10355 (N_10355,N_9933,N_9706);
and U10356 (N_10356,N_9869,N_9710);
and U10357 (N_10357,N_9722,N_9982);
nand U10358 (N_10358,N_9764,N_9843);
or U10359 (N_10359,N_9686,N_9681);
nor U10360 (N_10360,N_9905,N_9856);
and U10361 (N_10361,N_9966,N_9689);
or U10362 (N_10362,N_9915,N_9721);
and U10363 (N_10363,N_9890,N_9910);
and U10364 (N_10364,N_9724,N_9703);
xor U10365 (N_10365,N_9957,N_9991);
nand U10366 (N_10366,N_9984,N_9697);
nor U10367 (N_10367,N_9865,N_9748);
xnor U10368 (N_10368,N_9973,N_9737);
nand U10369 (N_10369,N_9714,N_9697);
nor U10370 (N_10370,N_9960,N_9929);
and U10371 (N_10371,N_9846,N_9899);
and U10372 (N_10372,N_9691,N_9981);
nor U10373 (N_10373,N_9707,N_9797);
or U10374 (N_10374,N_9704,N_9693);
or U10375 (N_10375,N_9746,N_9934);
and U10376 (N_10376,N_9809,N_9844);
nand U10377 (N_10377,N_9826,N_9671);
or U10378 (N_10378,N_9903,N_9954);
xnor U10379 (N_10379,N_9843,N_9929);
nor U10380 (N_10380,N_9656,N_9630);
or U10381 (N_10381,N_9829,N_9632);
nor U10382 (N_10382,N_9878,N_9799);
and U10383 (N_10383,N_9626,N_9766);
and U10384 (N_10384,N_9839,N_9957);
nor U10385 (N_10385,N_9806,N_9970);
nor U10386 (N_10386,N_9739,N_9776);
nand U10387 (N_10387,N_9876,N_9676);
and U10388 (N_10388,N_9746,N_9766);
and U10389 (N_10389,N_9745,N_9947);
or U10390 (N_10390,N_9632,N_9798);
or U10391 (N_10391,N_9826,N_9635);
or U10392 (N_10392,N_9777,N_9716);
or U10393 (N_10393,N_9620,N_9874);
and U10394 (N_10394,N_9694,N_9707);
or U10395 (N_10395,N_9634,N_9982);
nor U10396 (N_10396,N_9985,N_9627);
nor U10397 (N_10397,N_9875,N_9865);
nor U10398 (N_10398,N_9664,N_9895);
nand U10399 (N_10399,N_9805,N_9631);
nor U10400 (N_10400,N_10219,N_10258);
nand U10401 (N_10401,N_10051,N_10004);
nor U10402 (N_10402,N_10373,N_10358);
nor U10403 (N_10403,N_10244,N_10098);
or U10404 (N_10404,N_10111,N_10361);
and U10405 (N_10405,N_10251,N_10276);
and U10406 (N_10406,N_10049,N_10288);
and U10407 (N_10407,N_10372,N_10313);
and U10408 (N_10408,N_10337,N_10307);
or U10409 (N_10409,N_10318,N_10001);
or U10410 (N_10410,N_10347,N_10142);
and U10411 (N_10411,N_10390,N_10026);
nor U10412 (N_10412,N_10332,N_10386);
or U10413 (N_10413,N_10343,N_10385);
nand U10414 (N_10414,N_10353,N_10212);
or U10415 (N_10415,N_10223,N_10235);
xor U10416 (N_10416,N_10189,N_10155);
nor U10417 (N_10417,N_10099,N_10114);
and U10418 (N_10418,N_10160,N_10342);
xor U10419 (N_10419,N_10246,N_10222);
nand U10420 (N_10420,N_10133,N_10165);
and U10421 (N_10421,N_10330,N_10256);
xnor U10422 (N_10422,N_10170,N_10397);
xnor U10423 (N_10423,N_10064,N_10089);
nand U10424 (N_10424,N_10265,N_10029);
xor U10425 (N_10425,N_10094,N_10214);
xnor U10426 (N_10426,N_10243,N_10323);
or U10427 (N_10427,N_10032,N_10322);
and U10428 (N_10428,N_10125,N_10087);
or U10429 (N_10429,N_10270,N_10028);
or U10430 (N_10430,N_10017,N_10168);
xnor U10431 (N_10431,N_10092,N_10338);
xnor U10432 (N_10432,N_10317,N_10232);
or U10433 (N_10433,N_10305,N_10078);
and U10434 (N_10434,N_10107,N_10171);
xnor U10435 (N_10435,N_10069,N_10056);
and U10436 (N_10436,N_10203,N_10110);
xor U10437 (N_10437,N_10135,N_10269);
and U10438 (N_10438,N_10312,N_10309);
nor U10439 (N_10439,N_10197,N_10122);
nand U10440 (N_10440,N_10070,N_10082);
or U10441 (N_10441,N_10253,N_10341);
or U10442 (N_10442,N_10231,N_10134);
or U10443 (N_10443,N_10395,N_10141);
nand U10444 (N_10444,N_10228,N_10351);
and U10445 (N_10445,N_10040,N_10211);
nor U10446 (N_10446,N_10393,N_10076);
and U10447 (N_10447,N_10301,N_10140);
and U10448 (N_10448,N_10375,N_10149);
nand U10449 (N_10449,N_10006,N_10097);
and U10450 (N_10450,N_10195,N_10384);
nor U10451 (N_10451,N_10057,N_10349);
nand U10452 (N_10452,N_10273,N_10113);
or U10453 (N_10453,N_10013,N_10052);
and U10454 (N_10454,N_10039,N_10316);
xor U10455 (N_10455,N_10020,N_10396);
nand U10456 (N_10456,N_10074,N_10352);
nand U10457 (N_10457,N_10162,N_10234);
or U10458 (N_10458,N_10005,N_10216);
nor U10459 (N_10459,N_10024,N_10339);
xor U10460 (N_10460,N_10072,N_10278);
nand U10461 (N_10461,N_10310,N_10363);
nor U10462 (N_10462,N_10240,N_10146);
nor U10463 (N_10463,N_10055,N_10277);
and U10464 (N_10464,N_10043,N_10184);
and U10465 (N_10465,N_10311,N_10132);
nand U10466 (N_10466,N_10180,N_10178);
xnor U10467 (N_10467,N_10192,N_10071);
nand U10468 (N_10468,N_10336,N_10241);
nor U10469 (N_10469,N_10066,N_10002);
xnor U10470 (N_10470,N_10102,N_10209);
nand U10471 (N_10471,N_10117,N_10105);
xor U10472 (N_10472,N_10289,N_10210);
and U10473 (N_10473,N_10095,N_10154);
and U10474 (N_10474,N_10213,N_10166);
nor U10475 (N_10475,N_10164,N_10199);
nor U10476 (N_10476,N_10227,N_10088);
nor U10477 (N_10477,N_10255,N_10348);
or U10478 (N_10478,N_10179,N_10392);
and U10479 (N_10479,N_10237,N_10045);
nand U10480 (N_10480,N_10328,N_10290);
xnor U10481 (N_10481,N_10126,N_10294);
or U10482 (N_10482,N_10249,N_10173);
nor U10483 (N_10483,N_10371,N_10308);
and U10484 (N_10484,N_10297,N_10283);
or U10485 (N_10485,N_10137,N_10163);
or U10486 (N_10486,N_10370,N_10296);
or U10487 (N_10487,N_10355,N_10083);
and U10488 (N_10488,N_10100,N_10009);
and U10489 (N_10489,N_10226,N_10053);
xnor U10490 (N_10490,N_10200,N_10007);
nand U10491 (N_10491,N_10172,N_10067);
nand U10492 (N_10492,N_10127,N_10207);
and U10493 (N_10493,N_10236,N_10292);
or U10494 (N_10494,N_10389,N_10109);
and U10495 (N_10495,N_10187,N_10198);
and U10496 (N_10496,N_10048,N_10280);
xnor U10497 (N_10497,N_10224,N_10174);
nor U10498 (N_10498,N_10275,N_10248);
nand U10499 (N_10499,N_10144,N_10264);
or U10500 (N_10500,N_10383,N_10156);
or U10501 (N_10501,N_10181,N_10364);
nor U10502 (N_10502,N_10081,N_10038);
and U10503 (N_10503,N_10041,N_10027);
nor U10504 (N_10504,N_10357,N_10010);
nand U10505 (N_10505,N_10018,N_10217);
and U10506 (N_10506,N_10382,N_10016);
nor U10507 (N_10507,N_10025,N_10073);
xor U10508 (N_10508,N_10131,N_10194);
or U10509 (N_10509,N_10042,N_10011);
or U10510 (N_10510,N_10157,N_10360);
nand U10511 (N_10511,N_10138,N_10128);
or U10512 (N_10512,N_10037,N_10119);
nor U10513 (N_10513,N_10003,N_10334);
nor U10514 (N_10514,N_10115,N_10084);
and U10515 (N_10515,N_10359,N_10093);
nor U10516 (N_10516,N_10242,N_10054);
nand U10517 (N_10517,N_10201,N_10106);
nor U10518 (N_10518,N_10369,N_10065);
nor U10519 (N_10519,N_10196,N_10378);
or U10520 (N_10520,N_10143,N_10302);
nor U10521 (N_10521,N_10188,N_10077);
xor U10522 (N_10522,N_10068,N_10252);
nor U10523 (N_10523,N_10215,N_10233);
or U10524 (N_10524,N_10019,N_10285);
nand U10525 (N_10525,N_10368,N_10175);
or U10526 (N_10526,N_10101,N_10177);
or U10527 (N_10527,N_10075,N_10367);
xor U10528 (N_10528,N_10250,N_10014);
xor U10529 (N_10529,N_10298,N_10350);
nand U10530 (N_10530,N_10123,N_10022);
xor U10531 (N_10531,N_10379,N_10191);
or U10532 (N_10532,N_10090,N_10304);
nand U10533 (N_10533,N_10152,N_10345);
nand U10534 (N_10534,N_10047,N_10012);
xnor U10535 (N_10535,N_10259,N_10182);
and U10536 (N_10536,N_10186,N_10208);
nor U10537 (N_10537,N_10060,N_10169);
xnor U10538 (N_10538,N_10272,N_10079);
or U10539 (N_10539,N_10021,N_10116);
nor U10540 (N_10540,N_10120,N_10023);
nand U10541 (N_10541,N_10058,N_10033);
nand U10542 (N_10542,N_10303,N_10036);
nor U10543 (N_10543,N_10150,N_10254);
nand U10544 (N_10544,N_10377,N_10206);
or U10545 (N_10545,N_10324,N_10282);
xor U10546 (N_10546,N_10015,N_10085);
and U10547 (N_10547,N_10086,N_10333);
xnor U10548 (N_10548,N_10374,N_10391);
and U10549 (N_10549,N_10031,N_10221);
or U10550 (N_10550,N_10112,N_10262);
or U10551 (N_10551,N_10118,N_10096);
xnor U10552 (N_10552,N_10279,N_10145);
nor U10553 (N_10553,N_10387,N_10286);
or U10554 (N_10554,N_10062,N_10204);
and U10555 (N_10555,N_10121,N_10245);
nand U10556 (N_10556,N_10151,N_10108);
nor U10557 (N_10557,N_10176,N_10147);
nand U10558 (N_10558,N_10320,N_10356);
nand U10559 (N_10559,N_10329,N_10261);
or U10560 (N_10560,N_10291,N_10271);
nor U10561 (N_10561,N_10008,N_10319);
nor U10562 (N_10562,N_10344,N_10331);
and U10563 (N_10563,N_10394,N_10388);
and U10564 (N_10564,N_10340,N_10103);
xnor U10565 (N_10565,N_10354,N_10063);
or U10566 (N_10566,N_10030,N_10299);
and U10567 (N_10567,N_10185,N_10130);
and U10568 (N_10568,N_10284,N_10274);
and U10569 (N_10569,N_10000,N_10295);
or U10570 (N_10570,N_10193,N_10129);
and U10571 (N_10571,N_10380,N_10161);
or U10572 (N_10572,N_10266,N_10202);
and U10573 (N_10573,N_10326,N_10381);
nor U10574 (N_10574,N_10260,N_10050);
or U10575 (N_10575,N_10080,N_10238);
nand U10576 (N_10576,N_10239,N_10306);
or U10577 (N_10577,N_10281,N_10325);
xnor U10578 (N_10578,N_10225,N_10335);
or U10579 (N_10579,N_10139,N_10300);
nand U10580 (N_10580,N_10104,N_10293);
and U10581 (N_10581,N_10366,N_10321);
nand U10582 (N_10582,N_10314,N_10263);
or U10583 (N_10583,N_10376,N_10218);
and U10584 (N_10584,N_10190,N_10159);
nand U10585 (N_10585,N_10167,N_10044);
and U10586 (N_10586,N_10034,N_10148);
or U10587 (N_10587,N_10035,N_10158);
and U10588 (N_10588,N_10205,N_10183);
and U10589 (N_10589,N_10267,N_10136);
nor U10590 (N_10590,N_10230,N_10124);
nor U10591 (N_10591,N_10399,N_10268);
nand U10592 (N_10592,N_10220,N_10153);
nand U10593 (N_10593,N_10315,N_10362);
and U10594 (N_10594,N_10091,N_10346);
nand U10595 (N_10595,N_10061,N_10287);
or U10596 (N_10596,N_10365,N_10257);
nor U10597 (N_10597,N_10046,N_10398);
or U10598 (N_10598,N_10327,N_10229);
nand U10599 (N_10599,N_10247,N_10059);
or U10600 (N_10600,N_10136,N_10384);
nor U10601 (N_10601,N_10228,N_10018);
and U10602 (N_10602,N_10257,N_10154);
xnor U10603 (N_10603,N_10028,N_10393);
nor U10604 (N_10604,N_10300,N_10082);
or U10605 (N_10605,N_10385,N_10379);
or U10606 (N_10606,N_10262,N_10367);
xnor U10607 (N_10607,N_10340,N_10315);
nand U10608 (N_10608,N_10222,N_10144);
nand U10609 (N_10609,N_10230,N_10309);
nor U10610 (N_10610,N_10197,N_10117);
xor U10611 (N_10611,N_10393,N_10189);
xnor U10612 (N_10612,N_10056,N_10177);
nand U10613 (N_10613,N_10316,N_10090);
or U10614 (N_10614,N_10350,N_10132);
xor U10615 (N_10615,N_10295,N_10247);
xor U10616 (N_10616,N_10107,N_10258);
and U10617 (N_10617,N_10189,N_10033);
xnor U10618 (N_10618,N_10016,N_10229);
and U10619 (N_10619,N_10306,N_10140);
nand U10620 (N_10620,N_10287,N_10098);
nor U10621 (N_10621,N_10247,N_10183);
or U10622 (N_10622,N_10200,N_10337);
or U10623 (N_10623,N_10190,N_10000);
xnor U10624 (N_10624,N_10126,N_10183);
nor U10625 (N_10625,N_10244,N_10012);
xor U10626 (N_10626,N_10300,N_10054);
nor U10627 (N_10627,N_10051,N_10211);
nor U10628 (N_10628,N_10272,N_10055);
and U10629 (N_10629,N_10277,N_10366);
xnor U10630 (N_10630,N_10134,N_10261);
nand U10631 (N_10631,N_10348,N_10322);
xnor U10632 (N_10632,N_10017,N_10100);
or U10633 (N_10633,N_10250,N_10346);
nand U10634 (N_10634,N_10366,N_10185);
xnor U10635 (N_10635,N_10170,N_10001);
nor U10636 (N_10636,N_10368,N_10147);
nand U10637 (N_10637,N_10338,N_10011);
or U10638 (N_10638,N_10225,N_10185);
nand U10639 (N_10639,N_10352,N_10368);
nor U10640 (N_10640,N_10263,N_10362);
nand U10641 (N_10641,N_10395,N_10306);
xor U10642 (N_10642,N_10004,N_10398);
nand U10643 (N_10643,N_10326,N_10103);
or U10644 (N_10644,N_10165,N_10232);
xnor U10645 (N_10645,N_10360,N_10347);
xor U10646 (N_10646,N_10176,N_10343);
xor U10647 (N_10647,N_10023,N_10148);
and U10648 (N_10648,N_10003,N_10046);
nor U10649 (N_10649,N_10293,N_10225);
nor U10650 (N_10650,N_10008,N_10361);
nand U10651 (N_10651,N_10308,N_10352);
nand U10652 (N_10652,N_10143,N_10317);
xor U10653 (N_10653,N_10374,N_10161);
nand U10654 (N_10654,N_10065,N_10340);
nor U10655 (N_10655,N_10232,N_10023);
xnor U10656 (N_10656,N_10180,N_10117);
nor U10657 (N_10657,N_10257,N_10104);
nand U10658 (N_10658,N_10253,N_10169);
and U10659 (N_10659,N_10076,N_10130);
nor U10660 (N_10660,N_10245,N_10277);
and U10661 (N_10661,N_10101,N_10276);
nor U10662 (N_10662,N_10125,N_10311);
nand U10663 (N_10663,N_10008,N_10189);
xnor U10664 (N_10664,N_10097,N_10278);
nor U10665 (N_10665,N_10125,N_10369);
or U10666 (N_10666,N_10325,N_10023);
xnor U10667 (N_10667,N_10374,N_10319);
and U10668 (N_10668,N_10293,N_10159);
nor U10669 (N_10669,N_10165,N_10296);
or U10670 (N_10670,N_10079,N_10141);
and U10671 (N_10671,N_10203,N_10272);
or U10672 (N_10672,N_10380,N_10333);
or U10673 (N_10673,N_10196,N_10073);
xor U10674 (N_10674,N_10294,N_10132);
nor U10675 (N_10675,N_10322,N_10057);
or U10676 (N_10676,N_10232,N_10088);
nand U10677 (N_10677,N_10111,N_10162);
nand U10678 (N_10678,N_10251,N_10040);
nand U10679 (N_10679,N_10121,N_10332);
nor U10680 (N_10680,N_10220,N_10147);
nand U10681 (N_10681,N_10067,N_10298);
xnor U10682 (N_10682,N_10376,N_10154);
nand U10683 (N_10683,N_10123,N_10008);
or U10684 (N_10684,N_10310,N_10376);
and U10685 (N_10685,N_10354,N_10281);
nand U10686 (N_10686,N_10291,N_10305);
or U10687 (N_10687,N_10113,N_10119);
and U10688 (N_10688,N_10240,N_10363);
nor U10689 (N_10689,N_10103,N_10207);
and U10690 (N_10690,N_10020,N_10054);
nand U10691 (N_10691,N_10300,N_10173);
and U10692 (N_10692,N_10318,N_10280);
or U10693 (N_10693,N_10215,N_10296);
xor U10694 (N_10694,N_10099,N_10095);
and U10695 (N_10695,N_10378,N_10140);
nand U10696 (N_10696,N_10228,N_10074);
xor U10697 (N_10697,N_10186,N_10131);
and U10698 (N_10698,N_10279,N_10073);
and U10699 (N_10699,N_10157,N_10049);
or U10700 (N_10700,N_10294,N_10044);
xnor U10701 (N_10701,N_10272,N_10082);
or U10702 (N_10702,N_10073,N_10112);
or U10703 (N_10703,N_10265,N_10311);
xnor U10704 (N_10704,N_10217,N_10130);
and U10705 (N_10705,N_10288,N_10116);
or U10706 (N_10706,N_10021,N_10185);
and U10707 (N_10707,N_10233,N_10360);
and U10708 (N_10708,N_10008,N_10386);
or U10709 (N_10709,N_10114,N_10330);
or U10710 (N_10710,N_10002,N_10081);
nor U10711 (N_10711,N_10196,N_10101);
nand U10712 (N_10712,N_10111,N_10061);
nor U10713 (N_10713,N_10300,N_10276);
and U10714 (N_10714,N_10341,N_10344);
or U10715 (N_10715,N_10198,N_10072);
nand U10716 (N_10716,N_10095,N_10055);
or U10717 (N_10717,N_10247,N_10363);
nor U10718 (N_10718,N_10120,N_10280);
nor U10719 (N_10719,N_10259,N_10114);
xnor U10720 (N_10720,N_10354,N_10233);
or U10721 (N_10721,N_10140,N_10202);
nor U10722 (N_10722,N_10142,N_10093);
and U10723 (N_10723,N_10060,N_10035);
or U10724 (N_10724,N_10115,N_10029);
or U10725 (N_10725,N_10399,N_10047);
or U10726 (N_10726,N_10034,N_10302);
nor U10727 (N_10727,N_10045,N_10200);
xor U10728 (N_10728,N_10291,N_10292);
and U10729 (N_10729,N_10096,N_10237);
nor U10730 (N_10730,N_10362,N_10346);
and U10731 (N_10731,N_10088,N_10244);
nand U10732 (N_10732,N_10140,N_10165);
nor U10733 (N_10733,N_10179,N_10116);
or U10734 (N_10734,N_10021,N_10352);
xnor U10735 (N_10735,N_10252,N_10370);
nand U10736 (N_10736,N_10077,N_10057);
and U10737 (N_10737,N_10305,N_10221);
xnor U10738 (N_10738,N_10154,N_10204);
xor U10739 (N_10739,N_10108,N_10097);
xor U10740 (N_10740,N_10292,N_10132);
and U10741 (N_10741,N_10015,N_10395);
nor U10742 (N_10742,N_10258,N_10271);
or U10743 (N_10743,N_10012,N_10324);
nor U10744 (N_10744,N_10007,N_10186);
or U10745 (N_10745,N_10156,N_10186);
or U10746 (N_10746,N_10330,N_10312);
or U10747 (N_10747,N_10336,N_10259);
xnor U10748 (N_10748,N_10393,N_10101);
nor U10749 (N_10749,N_10043,N_10142);
nand U10750 (N_10750,N_10327,N_10002);
nand U10751 (N_10751,N_10156,N_10054);
nand U10752 (N_10752,N_10393,N_10172);
nor U10753 (N_10753,N_10053,N_10396);
or U10754 (N_10754,N_10167,N_10282);
and U10755 (N_10755,N_10072,N_10381);
and U10756 (N_10756,N_10007,N_10181);
xnor U10757 (N_10757,N_10023,N_10136);
or U10758 (N_10758,N_10123,N_10356);
or U10759 (N_10759,N_10127,N_10107);
and U10760 (N_10760,N_10087,N_10162);
or U10761 (N_10761,N_10065,N_10155);
nand U10762 (N_10762,N_10209,N_10274);
and U10763 (N_10763,N_10366,N_10183);
nor U10764 (N_10764,N_10288,N_10291);
and U10765 (N_10765,N_10152,N_10308);
xnor U10766 (N_10766,N_10104,N_10097);
nor U10767 (N_10767,N_10238,N_10027);
nor U10768 (N_10768,N_10018,N_10121);
nand U10769 (N_10769,N_10172,N_10236);
nand U10770 (N_10770,N_10382,N_10048);
nand U10771 (N_10771,N_10389,N_10229);
nor U10772 (N_10772,N_10013,N_10271);
xor U10773 (N_10773,N_10275,N_10198);
xor U10774 (N_10774,N_10278,N_10258);
xor U10775 (N_10775,N_10344,N_10095);
or U10776 (N_10776,N_10263,N_10262);
nand U10777 (N_10777,N_10125,N_10386);
or U10778 (N_10778,N_10381,N_10062);
nand U10779 (N_10779,N_10104,N_10388);
or U10780 (N_10780,N_10167,N_10185);
nor U10781 (N_10781,N_10126,N_10306);
or U10782 (N_10782,N_10262,N_10212);
and U10783 (N_10783,N_10384,N_10087);
nand U10784 (N_10784,N_10038,N_10196);
nor U10785 (N_10785,N_10281,N_10184);
nor U10786 (N_10786,N_10325,N_10085);
nand U10787 (N_10787,N_10288,N_10009);
nor U10788 (N_10788,N_10207,N_10327);
nand U10789 (N_10789,N_10252,N_10331);
nor U10790 (N_10790,N_10236,N_10075);
nand U10791 (N_10791,N_10352,N_10178);
nor U10792 (N_10792,N_10250,N_10372);
or U10793 (N_10793,N_10115,N_10092);
xnor U10794 (N_10794,N_10054,N_10174);
and U10795 (N_10795,N_10103,N_10208);
and U10796 (N_10796,N_10053,N_10166);
and U10797 (N_10797,N_10306,N_10320);
nand U10798 (N_10798,N_10178,N_10384);
or U10799 (N_10799,N_10368,N_10386);
and U10800 (N_10800,N_10452,N_10710);
or U10801 (N_10801,N_10423,N_10700);
nand U10802 (N_10802,N_10416,N_10497);
nor U10803 (N_10803,N_10521,N_10559);
nand U10804 (N_10804,N_10544,N_10421);
xnor U10805 (N_10805,N_10788,N_10750);
xor U10806 (N_10806,N_10549,N_10543);
nor U10807 (N_10807,N_10512,N_10786);
nor U10808 (N_10808,N_10688,N_10578);
and U10809 (N_10809,N_10432,N_10552);
nor U10810 (N_10810,N_10734,N_10517);
xnor U10811 (N_10811,N_10585,N_10584);
or U10812 (N_10812,N_10437,N_10637);
xnor U10813 (N_10813,N_10694,N_10796);
nand U10814 (N_10814,N_10611,N_10696);
or U10815 (N_10815,N_10771,N_10422);
xnor U10816 (N_10816,N_10539,N_10572);
nor U10817 (N_10817,N_10442,N_10516);
xor U10818 (N_10818,N_10684,N_10769);
xnor U10819 (N_10819,N_10547,N_10441);
nand U10820 (N_10820,N_10460,N_10721);
and U10821 (N_10821,N_10486,N_10733);
nor U10822 (N_10822,N_10480,N_10514);
nand U10823 (N_10823,N_10557,N_10616);
or U10824 (N_10824,N_10610,N_10476);
or U10825 (N_10825,N_10618,N_10551);
or U10826 (N_10826,N_10400,N_10474);
or U10827 (N_10827,N_10609,N_10785);
nor U10828 (N_10828,N_10711,N_10633);
and U10829 (N_10829,N_10670,N_10523);
and U10830 (N_10830,N_10504,N_10573);
xnor U10831 (N_10831,N_10406,N_10493);
or U10832 (N_10832,N_10770,N_10553);
nand U10833 (N_10833,N_10583,N_10600);
or U10834 (N_10834,N_10653,N_10648);
and U10835 (N_10835,N_10424,N_10625);
xnor U10836 (N_10836,N_10703,N_10628);
xor U10837 (N_10837,N_10784,N_10768);
or U10838 (N_10838,N_10562,N_10759);
nor U10839 (N_10839,N_10465,N_10425);
or U10840 (N_10840,N_10738,N_10530);
nor U10841 (N_10841,N_10753,N_10718);
xor U10842 (N_10842,N_10494,N_10613);
or U10843 (N_10843,N_10459,N_10495);
and U10844 (N_10844,N_10436,N_10720);
or U10845 (N_10845,N_10498,N_10568);
nor U10846 (N_10846,N_10443,N_10751);
nor U10847 (N_10847,N_10579,N_10636);
and U10848 (N_10848,N_10640,N_10737);
xor U10849 (N_10849,N_10453,N_10566);
nand U10850 (N_10850,N_10415,N_10546);
and U10851 (N_10851,N_10524,N_10657);
or U10852 (N_10852,N_10508,N_10499);
nor U10853 (N_10853,N_10599,N_10799);
nor U10854 (N_10854,N_10680,N_10775);
xor U10855 (N_10855,N_10575,N_10622);
and U10856 (N_10856,N_10596,N_10463);
or U10857 (N_10857,N_10627,N_10590);
and U10858 (N_10858,N_10492,N_10401);
xor U10859 (N_10859,N_10438,N_10444);
xor U10860 (N_10860,N_10647,N_10763);
and U10861 (N_10861,N_10540,N_10686);
nand U10862 (N_10862,N_10532,N_10794);
nand U10863 (N_10863,N_10702,N_10467);
or U10864 (N_10864,N_10764,N_10761);
xnor U10865 (N_10865,N_10665,N_10780);
nand U10866 (N_10866,N_10748,N_10526);
nand U10867 (N_10867,N_10477,N_10587);
and U10868 (N_10868,N_10614,N_10560);
nand U10869 (N_10869,N_10687,N_10715);
or U10870 (N_10870,N_10663,N_10740);
xor U10871 (N_10871,N_10722,N_10773);
or U10872 (N_10872,N_10791,N_10641);
nand U10873 (N_10873,N_10440,N_10458);
nor U10874 (N_10874,N_10790,N_10746);
nor U10875 (N_10875,N_10732,N_10659);
xnor U10876 (N_10876,N_10669,N_10646);
xor U10877 (N_10877,N_10515,N_10554);
xor U10878 (N_10878,N_10541,N_10760);
xnor U10879 (N_10879,N_10623,N_10581);
xor U10880 (N_10880,N_10472,N_10586);
or U10881 (N_10881,N_10531,N_10548);
nand U10882 (N_10882,N_10608,N_10580);
nand U10883 (N_10883,N_10419,N_10409);
and U10884 (N_10884,N_10466,N_10735);
and U10885 (N_10885,N_10707,N_10675);
or U10886 (N_10886,N_10448,N_10709);
nor U10887 (N_10887,N_10783,N_10428);
and U10888 (N_10888,N_10676,N_10781);
xnor U10889 (N_10889,N_10471,N_10574);
nand U10890 (N_10890,N_10649,N_10506);
and U10891 (N_10891,N_10723,N_10536);
xnor U10892 (N_10892,N_10408,N_10542);
nor U10893 (N_10893,N_10652,N_10749);
xor U10894 (N_10894,N_10456,N_10643);
and U10895 (N_10895,N_10435,N_10538);
or U10896 (N_10896,N_10565,N_10621);
and U10897 (N_10897,N_10682,N_10741);
and U10898 (N_10898,N_10602,N_10489);
and U10899 (N_10899,N_10752,N_10607);
nand U10900 (N_10900,N_10658,N_10561);
nor U10901 (N_10901,N_10569,N_10550);
and U10902 (N_10902,N_10701,N_10592);
nor U10903 (N_10903,N_10782,N_10606);
nand U10904 (N_10904,N_10772,N_10555);
and U10905 (N_10905,N_10427,N_10457);
or U10906 (N_10906,N_10582,N_10730);
nand U10907 (N_10907,N_10545,N_10470);
nand U10908 (N_10908,N_10713,N_10413);
xnor U10909 (N_10909,N_10520,N_10511);
and U10910 (N_10910,N_10513,N_10449);
nand U10911 (N_10911,N_10671,N_10434);
or U10912 (N_10912,N_10402,N_10431);
nor U10913 (N_10913,N_10795,N_10525);
nor U10914 (N_10914,N_10461,N_10447);
and U10915 (N_10915,N_10655,N_10726);
nor U10916 (N_10916,N_10482,N_10484);
or U10917 (N_10917,N_10635,N_10598);
nand U10918 (N_10918,N_10535,N_10660);
nand U10919 (N_10919,N_10507,N_10510);
or U10920 (N_10920,N_10464,N_10604);
nor U10921 (N_10921,N_10481,N_10755);
or U10922 (N_10922,N_10490,N_10639);
and U10923 (N_10923,N_10736,N_10527);
nor U10924 (N_10924,N_10757,N_10597);
and U10925 (N_10925,N_10762,N_10570);
or U10926 (N_10926,N_10681,N_10727);
xnor U10927 (N_10927,N_10758,N_10689);
xnor U10928 (N_10928,N_10767,N_10411);
or U10929 (N_10929,N_10468,N_10792);
and U10930 (N_10930,N_10629,N_10414);
nand U10931 (N_10931,N_10712,N_10503);
or U10932 (N_10932,N_10704,N_10430);
nand U10933 (N_10933,N_10502,N_10673);
nor U10934 (N_10934,N_10487,N_10403);
or U10935 (N_10935,N_10674,N_10683);
nand U10936 (N_10936,N_10473,N_10787);
nand U10937 (N_10937,N_10619,N_10743);
xor U10938 (N_10938,N_10501,N_10708);
and U10939 (N_10939,N_10651,N_10693);
nand U10940 (N_10940,N_10500,N_10601);
nand U10941 (N_10941,N_10667,N_10631);
nand U10942 (N_10942,N_10662,N_10634);
xor U10943 (N_10943,N_10410,N_10603);
xor U10944 (N_10944,N_10698,N_10563);
nand U10945 (N_10945,N_10576,N_10479);
nor U10946 (N_10946,N_10699,N_10446);
nor U10947 (N_10947,N_10672,N_10725);
nor U10948 (N_10948,N_10778,N_10462);
nand U10949 (N_10949,N_10505,N_10685);
xor U10950 (N_10950,N_10417,N_10533);
xor U10951 (N_10951,N_10776,N_10588);
nand U10952 (N_10952,N_10638,N_10656);
nor U10953 (N_10953,N_10766,N_10529);
xnor U10954 (N_10954,N_10678,N_10626);
nor U10955 (N_10955,N_10666,N_10595);
nand U10956 (N_10956,N_10624,N_10668);
nor U10957 (N_10957,N_10528,N_10691);
and U10958 (N_10958,N_10729,N_10793);
nor U10959 (N_10959,N_10485,N_10483);
xor U10960 (N_10960,N_10605,N_10612);
nand U10961 (N_10961,N_10742,N_10577);
or U10962 (N_10962,N_10519,N_10739);
nand U10963 (N_10963,N_10664,N_10779);
or U10964 (N_10964,N_10469,N_10537);
xnor U10965 (N_10965,N_10717,N_10589);
and U10966 (N_10966,N_10426,N_10714);
and U10967 (N_10967,N_10747,N_10439);
xor U10968 (N_10968,N_10744,N_10455);
or U10969 (N_10969,N_10650,N_10774);
nand U10970 (N_10970,N_10496,N_10491);
and U10971 (N_10971,N_10690,N_10642);
and U10972 (N_10972,N_10420,N_10522);
and U10973 (N_10973,N_10591,N_10475);
and U10974 (N_10974,N_10719,N_10412);
nand U10975 (N_10975,N_10478,N_10797);
or U10976 (N_10976,N_10620,N_10556);
or U10977 (N_10977,N_10756,N_10404);
nor U10978 (N_10978,N_10765,N_10567);
nor U10979 (N_10979,N_10754,N_10644);
nand U10980 (N_10980,N_10558,N_10445);
nor U10981 (N_10981,N_10617,N_10645);
nand U10982 (N_10982,N_10509,N_10593);
or U10983 (N_10983,N_10488,N_10654);
nand U10984 (N_10984,N_10789,N_10728);
nand U10985 (N_10985,N_10705,N_10777);
xnor U10986 (N_10986,N_10632,N_10407);
nor U10987 (N_10987,N_10716,N_10534);
nand U10988 (N_10988,N_10706,N_10692);
or U10989 (N_10989,N_10450,N_10731);
nand U10990 (N_10990,N_10571,N_10451);
xor U10991 (N_10991,N_10615,N_10518);
nand U10992 (N_10992,N_10679,N_10697);
and U10993 (N_10993,N_10564,N_10724);
or U10994 (N_10994,N_10405,N_10630);
xor U10995 (N_10995,N_10695,N_10429);
nor U10996 (N_10996,N_10677,N_10433);
nand U10997 (N_10997,N_10594,N_10661);
nor U10998 (N_10998,N_10745,N_10418);
nor U10999 (N_10999,N_10798,N_10454);
xor U11000 (N_11000,N_10559,N_10650);
nor U11001 (N_11001,N_10649,N_10454);
nand U11002 (N_11002,N_10735,N_10471);
and U11003 (N_11003,N_10610,N_10620);
or U11004 (N_11004,N_10762,N_10401);
and U11005 (N_11005,N_10673,N_10482);
xor U11006 (N_11006,N_10725,N_10768);
xor U11007 (N_11007,N_10518,N_10500);
nand U11008 (N_11008,N_10674,N_10762);
xnor U11009 (N_11009,N_10493,N_10514);
and U11010 (N_11010,N_10776,N_10698);
nor U11011 (N_11011,N_10688,N_10536);
nor U11012 (N_11012,N_10674,N_10495);
nand U11013 (N_11013,N_10432,N_10741);
nand U11014 (N_11014,N_10593,N_10516);
or U11015 (N_11015,N_10706,N_10477);
and U11016 (N_11016,N_10509,N_10791);
nor U11017 (N_11017,N_10531,N_10484);
xor U11018 (N_11018,N_10595,N_10407);
and U11019 (N_11019,N_10700,N_10588);
xor U11020 (N_11020,N_10684,N_10637);
nand U11021 (N_11021,N_10449,N_10401);
xor U11022 (N_11022,N_10594,N_10671);
nor U11023 (N_11023,N_10726,N_10546);
xnor U11024 (N_11024,N_10527,N_10626);
xor U11025 (N_11025,N_10655,N_10466);
and U11026 (N_11026,N_10441,N_10691);
nand U11027 (N_11027,N_10567,N_10420);
xor U11028 (N_11028,N_10634,N_10517);
nor U11029 (N_11029,N_10461,N_10453);
nand U11030 (N_11030,N_10440,N_10759);
nor U11031 (N_11031,N_10474,N_10783);
nand U11032 (N_11032,N_10710,N_10409);
xor U11033 (N_11033,N_10633,N_10477);
nand U11034 (N_11034,N_10518,N_10496);
nand U11035 (N_11035,N_10616,N_10405);
and U11036 (N_11036,N_10696,N_10562);
or U11037 (N_11037,N_10650,N_10482);
nand U11038 (N_11038,N_10442,N_10607);
or U11039 (N_11039,N_10467,N_10412);
nand U11040 (N_11040,N_10494,N_10752);
or U11041 (N_11041,N_10431,N_10596);
nand U11042 (N_11042,N_10458,N_10727);
or U11043 (N_11043,N_10400,N_10673);
xnor U11044 (N_11044,N_10718,N_10798);
and U11045 (N_11045,N_10646,N_10737);
or U11046 (N_11046,N_10737,N_10632);
nor U11047 (N_11047,N_10516,N_10597);
and U11048 (N_11048,N_10773,N_10632);
or U11049 (N_11049,N_10787,N_10765);
or U11050 (N_11050,N_10562,N_10545);
xnor U11051 (N_11051,N_10513,N_10699);
nand U11052 (N_11052,N_10465,N_10574);
or U11053 (N_11053,N_10780,N_10634);
nand U11054 (N_11054,N_10452,N_10794);
and U11055 (N_11055,N_10516,N_10729);
nand U11056 (N_11056,N_10685,N_10495);
xnor U11057 (N_11057,N_10799,N_10504);
and U11058 (N_11058,N_10426,N_10785);
and U11059 (N_11059,N_10630,N_10494);
or U11060 (N_11060,N_10422,N_10656);
xnor U11061 (N_11061,N_10413,N_10749);
or U11062 (N_11062,N_10493,N_10694);
and U11063 (N_11063,N_10776,N_10710);
nand U11064 (N_11064,N_10401,N_10703);
and U11065 (N_11065,N_10410,N_10426);
nor U11066 (N_11066,N_10649,N_10788);
or U11067 (N_11067,N_10687,N_10642);
nor U11068 (N_11068,N_10469,N_10687);
and U11069 (N_11069,N_10600,N_10705);
or U11070 (N_11070,N_10762,N_10520);
and U11071 (N_11071,N_10624,N_10578);
nor U11072 (N_11072,N_10530,N_10625);
and U11073 (N_11073,N_10570,N_10723);
nor U11074 (N_11074,N_10566,N_10491);
and U11075 (N_11075,N_10583,N_10640);
or U11076 (N_11076,N_10613,N_10437);
nor U11077 (N_11077,N_10571,N_10642);
or U11078 (N_11078,N_10736,N_10752);
nand U11079 (N_11079,N_10770,N_10402);
xor U11080 (N_11080,N_10775,N_10504);
or U11081 (N_11081,N_10743,N_10657);
or U11082 (N_11082,N_10552,N_10672);
xnor U11083 (N_11083,N_10466,N_10639);
and U11084 (N_11084,N_10668,N_10778);
or U11085 (N_11085,N_10501,N_10443);
or U11086 (N_11086,N_10506,N_10624);
or U11087 (N_11087,N_10603,N_10583);
or U11088 (N_11088,N_10502,N_10719);
nand U11089 (N_11089,N_10740,N_10632);
nand U11090 (N_11090,N_10532,N_10475);
or U11091 (N_11091,N_10558,N_10410);
or U11092 (N_11092,N_10528,N_10517);
nor U11093 (N_11093,N_10671,N_10418);
nand U11094 (N_11094,N_10765,N_10591);
nor U11095 (N_11095,N_10415,N_10562);
nand U11096 (N_11096,N_10485,N_10567);
and U11097 (N_11097,N_10512,N_10441);
nand U11098 (N_11098,N_10788,N_10748);
nand U11099 (N_11099,N_10508,N_10486);
xnor U11100 (N_11100,N_10606,N_10564);
xnor U11101 (N_11101,N_10483,N_10449);
nor U11102 (N_11102,N_10697,N_10471);
or U11103 (N_11103,N_10541,N_10749);
and U11104 (N_11104,N_10648,N_10675);
nand U11105 (N_11105,N_10660,N_10714);
and U11106 (N_11106,N_10482,N_10699);
nor U11107 (N_11107,N_10686,N_10798);
xnor U11108 (N_11108,N_10767,N_10599);
nor U11109 (N_11109,N_10555,N_10658);
nand U11110 (N_11110,N_10691,N_10651);
and U11111 (N_11111,N_10523,N_10450);
nor U11112 (N_11112,N_10459,N_10597);
nor U11113 (N_11113,N_10628,N_10531);
nand U11114 (N_11114,N_10699,N_10757);
or U11115 (N_11115,N_10529,N_10505);
or U11116 (N_11116,N_10454,N_10438);
or U11117 (N_11117,N_10594,N_10600);
nand U11118 (N_11118,N_10599,N_10704);
nor U11119 (N_11119,N_10636,N_10587);
nand U11120 (N_11120,N_10675,N_10551);
and U11121 (N_11121,N_10776,N_10633);
xor U11122 (N_11122,N_10612,N_10721);
or U11123 (N_11123,N_10633,N_10703);
nand U11124 (N_11124,N_10635,N_10455);
nor U11125 (N_11125,N_10619,N_10723);
or U11126 (N_11126,N_10549,N_10408);
or U11127 (N_11127,N_10747,N_10665);
nand U11128 (N_11128,N_10767,N_10522);
or U11129 (N_11129,N_10534,N_10732);
xnor U11130 (N_11130,N_10416,N_10514);
and U11131 (N_11131,N_10688,N_10730);
nor U11132 (N_11132,N_10625,N_10453);
and U11133 (N_11133,N_10664,N_10417);
xor U11134 (N_11134,N_10703,N_10533);
xor U11135 (N_11135,N_10711,N_10726);
nand U11136 (N_11136,N_10665,N_10488);
and U11137 (N_11137,N_10650,N_10448);
or U11138 (N_11138,N_10693,N_10505);
or U11139 (N_11139,N_10659,N_10685);
xor U11140 (N_11140,N_10650,N_10541);
xor U11141 (N_11141,N_10620,N_10628);
xnor U11142 (N_11142,N_10584,N_10552);
nand U11143 (N_11143,N_10609,N_10403);
xor U11144 (N_11144,N_10531,N_10403);
and U11145 (N_11145,N_10449,N_10746);
nor U11146 (N_11146,N_10640,N_10659);
and U11147 (N_11147,N_10755,N_10596);
nor U11148 (N_11148,N_10598,N_10540);
nor U11149 (N_11149,N_10418,N_10679);
nor U11150 (N_11150,N_10541,N_10757);
nor U11151 (N_11151,N_10429,N_10440);
xnor U11152 (N_11152,N_10563,N_10706);
nor U11153 (N_11153,N_10527,N_10542);
or U11154 (N_11154,N_10581,N_10610);
xnor U11155 (N_11155,N_10445,N_10573);
xor U11156 (N_11156,N_10671,N_10604);
nor U11157 (N_11157,N_10571,N_10639);
or U11158 (N_11158,N_10605,N_10781);
xnor U11159 (N_11159,N_10758,N_10416);
and U11160 (N_11160,N_10753,N_10549);
and U11161 (N_11161,N_10681,N_10466);
xor U11162 (N_11162,N_10716,N_10410);
xnor U11163 (N_11163,N_10680,N_10773);
or U11164 (N_11164,N_10520,N_10614);
xor U11165 (N_11165,N_10733,N_10769);
and U11166 (N_11166,N_10494,N_10749);
nand U11167 (N_11167,N_10627,N_10541);
nand U11168 (N_11168,N_10452,N_10703);
and U11169 (N_11169,N_10776,N_10502);
or U11170 (N_11170,N_10580,N_10533);
xnor U11171 (N_11171,N_10576,N_10631);
nor U11172 (N_11172,N_10713,N_10727);
and U11173 (N_11173,N_10791,N_10739);
nor U11174 (N_11174,N_10715,N_10470);
or U11175 (N_11175,N_10690,N_10468);
and U11176 (N_11176,N_10783,N_10623);
or U11177 (N_11177,N_10532,N_10520);
nand U11178 (N_11178,N_10559,N_10550);
xor U11179 (N_11179,N_10528,N_10728);
xor U11180 (N_11180,N_10431,N_10775);
and U11181 (N_11181,N_10413,N_10536);
nor U11182 (N_11182,N_10582,N_10510);
nor U11183 (N_11183,N_10659,N_10528);
nor U11184 (N_11184,N_10611,N_10498);
nand U11185 (N_11185,N_10650,N_10529);
and U11186 (N_11186,N_10736,N_10732);
nor U11187 (N_11187,N_10547,N_10644);
nand U11188 (N_11188,N_10544,N_10493);
and U11189 (N_11189,N_10457,N_10546);
xor U11190 (N_11190,N_10419,N_10696);
or U11191 (N_11191,N_10466,N_10607);
or U11192 (N_11192,N_10769,N_10595);
nand U11193 (N_11193,N_10666,N_10463);
or U11194 (N_11194,N_10744,N_10735);
nand U11195 (N_11195,N_10679,N_10740);
or U11196 (N_11196,N_10728,N_10766);
or U11197 (N_11197,N_10742,N_10422);
and U11198 (N_11198,N_10505,N_10497);
and U11199 (N_11199,N_10765,N_10709);
and U11200 (N_11200,N_11063,N_11105);
nand U11201 (N_11201,N_11068,N_10859);
xnor U11202 (N_11202,N_10897,N_10885);
nor U11203 (N_11203,N_11128,N_10836);
nor U11204 (N_11204,N_11053,N_10888);
xnor U11205 (N_11205,N_11048,N_11189);
xor U11206 (N_11206,N_11121,N_10866);
or U11207 (N_11207,N_11066,N_11170);
or U11208 (N_11208,N_11138,N_10861);
or U11209 (N_11209,N_10921,N_11113);
nor U11210 (N_11210,N_10907,N_11158);
or U11211 (N_11211,N_10905,N_11093);
xor U11212 (N_11212,N_10973,N_10972);
or U11213 (N_11213,N_11036,N_11132);
and U11214 (N_11214,N_11007,N_11012);
nor U11215 (N_11215,N_11051,N_11155);
or U11216 (N_11216,N_10954,N_10994);
xor U11217 (N_11217,N_10842,N_10804);
xor U11218 (N_11218,N_10814,N_11035);
nor U11219 (N_11219,N_10989,N_11139);
or U11220 (N_11220,N_11116,N_10943);
nand U11221 (N_11221,N_11129,N_11074);
xor U11222 (N_11222,N_11131,N_10818);
nand U11223 (N_11223,N_10813,N_11173);
xor U11224 (N_11224,N_11145,N_10961);
or U11225 (N_11225,N_10894,N_11147);
nand U11226 (N_11226,N_11161,N_10987);
xor U11227 (N_11227,N_10940,N_10979);
nand U11228 (N_11228,N_10837,N_11049);
nor U11229 (N_11229,N_10909,N_10832);
and U11230 (N_11230,N_11032,N_10857);
or U11231 (N_11231,N_10974,N_10852);
nor U11232 (N_11232,N_11187,N_10957);
and U11233 (N_11233,N_11120,N_10944);
nor U11234 (N_11234,N_10945,N_10825);
or U11235 (N_11235,N_11125,N_11033);
nor U11236 (N_11236,N_10868,N_11015);
xnor U11237 (N_11237,N_10838,N_10934);
nor U11238 (N_11238,N_10995,N_11002);
or U11239 (N_11239,N_10926,N_10935);
or U11240 (N_11240,N_10819,N_10924);
and U11241 (N_11241,N_10920,N_10919);
xor U11242 (N_11242,N_10906,N_10850);
or U11243 (N_11243,N_10834,N_11045);
or U11244 (N_11244,N_10878,N_10965);
and U11245 (N_11245,N_11117,N_11114);
nor U11246 (N_11246,N_10928,N_11110);
xor U11247 (N_11247,N_11177,N_10848);
and U11248 (N_11248,N_10996,N_11008);
xnor U11249 (N_11249,N_10922,N_11169);
or U11250 (N_11250,N_10830,N_11181);
and U11251 (N_11251,N_10964,N_10971);
nor U11252 (N_11252,N_11119,N_11106);
xor U11253 (N_11253,N_10929,N_10820);
or U11254 (N_11254,N_11149,N_10948);
and U11255 (N_11255,N_10843,N_10821);
nor U11256 (N_11256,N_11148,N_10913);
nor U11257 (N_11257,N_11054,N_11073);
or U11258 (N_11258,N_11030,N_10895);
or U11259 (N_11259,N_10982,N_10882);
or U11260 (N_11260,N_11004,N_11141);
or U11261 (N_11261,N_10855,N_11070);
nand U11262 (N_11262,N_11182,N_11130);
nand U11263 (N_11263,N_11183,N_11099);
nand U11264 (N_11264,N_11024,N_11025);
or U11265 (N_11265,N_11162,N_10846);
nand U11266 (N_11266,N_10849,N_11082);
or U11267 (N_11267,N_11018,N_10997);
nand U11268 (N_11268,N_11014,N_11109);
or U11269 (N_11269,N_10899,N_10839);
or U11270 (N_11270,N_11151,N_10864);
xnor U11271 (N_11271,N_10962,N_10931);
and U11272 (N_11272,N_11010,N_10960);
and U11273 (N_11273,N_11076,N_10952);
nor U11274 (N_11274,N_10941,N_11056);
or U11275 (N_11275,N_11194,N_11091);
and U11276 (N_11276,N_11192,N_10956);
nand U11277 (N_11277,N_10873,N_11188);
or U11278 (N_11278,N_11159,N_10817);
nand U11279 (N_11279,N_11026,N_11034);
xnor U11280 (N_11280,N_11011,N_11016);
xor U11281 (N_11281,N_11152,N_11174);
and U11282 (N_11282,N_10917,N_11107);
or U11283 (N_11283,N_11031,N_11144);
xor U11284 (N_11284,N_10884,N_11175);
nor U11285 (N_11285,N_10865,N_11085);
nor U11286 (N_11286,N_10910,N_11153);
xor U11287 (N_11287,N_10851,N_10876);
xor U11288 (N_11288,N_11111,N_11124);
nor U11289 (N_11289,N_11084,N_10985);
and U11290 (N_11290,N_10856,N_11042);
nand U11291 (N_11291,N_10992,N_10886);
nor U11292 (N_11292,N_10988,N_10900);
and U11293 (N_11293,N_10875,N_11087);
and U11294 (N_11294,N_11058,N_10806);
nor U11295 (N_11295,N_10959,N_11140);
nand U11296 (N_11296,N_10809,N_10808);
nor U11297 (N_11297,N_11083,N_11168);
or U11298 (N_11298,N_10860,N_10918);
xor U11299 (N_11299,N_11071,N_10903);
or U11300 (N_11300,N_11143,N_10984);
nand U11301 (N_11301,N_10999,N_10896);
nor U11302 (N_11302,N_10932,N_11134);
xor U11303 (N_11303,N_10829,N_11163);
or U11304 (N_11304,N_10841,N_11092);
nand U11305 (N_11305,N_10863,N_11179);
or U11306 (N_11306,N_10810,N_11061);
xnor U11307 (N_11307,N_11190,N_10807);
xor U11308 (N_11308,N_11052,N_11006);
or U11309 (N_11309,N_10822,N_10862);
xnor U11310 (N_11310,N_11046,N_10923);
nor U11311 (N_11311,N_11003,N_11047);
nor U11312 (N_11312,N_11127,N_10847);
xor U11313 (N_11313,N_10812,N_11167);
and U11314 (N_11314,N_11094,N_11098);
or U11315 (N_11315,N_10904,N_10950);
nand U11316 (N_11316,N_11199,N_11081);
nor U11317 (N_11317,N_11044,N_10867);
nand U11318 (N_11318,N_10916,N_11009);
xor U11319 (N_11319,N_10898,N_11108);
or U11320 (N_11320,N_11126,N_11089);
and U11321 (N_11321,N_11193,N_11095);
and U11322 (N_11322,N_11112,N_10975);
and U11323 (N_11323,N_10854,N_10968);
or U11324 (N_11324,N_11028,N_11135);
xnor U11325 (N_11325,N_10811,N_10815);
nor U11326 (N_11326,N_10976,N_10990);
xor U11327 (N_11327,N_10933,N_10947);
and U11328 (N_11328,N_10883,N_10823);
and U11329 (N_11329,N_11022,N_11029);
xor U11330 (N_11330,N_10936,N_11078);
and U11331 (N_11331,N_11180,N_11186);
nand U11332 (N_11332,N_10998,N_11142);
xnor U11333 (N_11333,N_11137,N_11017);
nand U11334 (N_11334,N_10893,N_11039);
or U11335 (N_11335,N_11164,N_11103);
or U11336 (N_11336,N_11069,N_10833);
and U11337 (N_11337,N_11096,N_10914);
xor U11338 (N_11338,N_11156,N_10970);
and U11339 (N_11339,N_10872,N_10844);
or U11340 (N_11340,N_11086,N_10892);
xnor U11341 (N_11341,N_10958,N_10966);
or U11342 (N_11342,N_10963,N_11020);
or U11343 (N_11343,N_11037,N_10912);
nand U11344 (N_11344,N_10889,N_10942);
and U11345 (N_11345,N_10877,N_11057);
xnor U11346 (N_11346,N_10800,N_11185);
nand U11347 (N_11347,N_10927,N_10993);
nor U11348 (N_11348,N_10828,N_11067);
xor U11349 (N_11349,N_10802,N_11100);
xnor U11350 (N_11350,N_10840,N_11178);
nor U11351 (N_11351,N_10801,N_10967);
nor U11352 (N_11352,N_10953,N_11040);
and U11353 (N_11353,N_10890,N_10930);
and U11354 (N_11354,N_10949,N_10925);
and U11355 (N_11355,N_11133,N_10835);
or U11356 (N_11356,N_10858,N_11005);
xor U11357 (N_11357,N_10938,N_10880);
nor U11358 (N_11358,N_11088,N_10939);
or U11359 (N_11359,N_10845,N_10853);
and U11360 (N_11360,N_10827,N_11171);
nand U11361 (N_11361,N_10955,N_11176);
nor U11362 (N_11362,N_11072,N_11050);
nor U11363 (N_11363,N_10911,N_11136);
nand U11364 (N_11364,N_10937,N_11001);
xnor U11365 (N_11365,N_11097,N_11165);
nand U11366 (N_11366,N_11080,N_10969);
xnor U11367 (N_11367,N_11184,N_11019);
nor U11368 (N_11368,N_11023,N_10915);
xnor U11369 (N_11369,N_11059,N_10977);
or U11370 (N_11370,N_11191,N_11043);
or U11371 (N_11371,N_10983,N_11077);
xor U11372 (N_11372,N_11123,N_11075);
nand U11373 (N_11373,N_11196,N_11195);
nand U11374 (N_11374,N_11150,N_11090);
nor U11375 (N_11375,N_10908,N_11038);
or U11376 (N_11376,N_10986,N_10816);
xnor U11377 (N_11377,N_10831,N_10980);
or U11378 (N_11378,N_10879,N_10824);
nor U11379 (N_11379,N_11122,N_11157);
nor U11380 (N_11380,N_10901,N_10887);
nand U11381 (N_11381,N_11102,N_10946);
nor U11382 (N_11382,N_11198,N_10871);
nor U11383 (N_11383,N_10902,N_11064);
and U11384 (N_11384,N_11027,N_11065);
nand U11385 (N_11385,N_11041,N_10869);
nor U11386 (N_11386,N_10874,N_11079);
nor U11387 (N_11387,N_11062,N_11060);
xor U11388 (N_11388,N_11172,N_11000);
xnor U11389 (N_11389,N_10978,N_10991);
or U11390 (N_11390,N_10803,N_11118);
xor U11391 (N_11391,N_11115,N_11146);
nand U11392 (N_11392,N_10951,N_10826);
or U11393 (N_11393,N_11055,N_11101);
xnor U11394 (N_11394,N_10891,N_11013);
nand U11395 (N_11395,N_10881,N_10981);
nand U11396 (N_11396,N_11154,N_11021);
nand U11397 (N_11397,N_11160,N_10805);
xor U11398 (N_11398,N_10870,N_11197);
or U11399 (N_11399,N_11166,N_11104);
xnor U11400 (N_11400,N_11031,N_11156);
or U11401 (N_11401,N_11106,N_10947);
nor U11402 (N_11402,N_10928,N_11076);
nand U11403 (N_11403,N_11060,N_11055);
xnor U11404 (N_11404,N_11031,N_10828);
nor U11405 (N_11405,N_10933,N_11084);
and U11406 (N_11406,N_10907,N_10993);
and U11407 (N_11407,N_11108,N_11050);
or U11408 (N_11408,N_11159,N_10858);
or U11409 (N_11409,N_10988,N_10868);
and U11410 (N_11410,N_11062,N_11034);
nor U11411 (N_11411,N_11034,N_10893);
nor U11412 (N_11412,N_11112,N_11172);
nor U11413 (N_11413,N_10929,N_11110);
xor U11414 (N_11414,N_11086,N_11024);
nand U11415 (N_11415,N_11181,N_10855);
nor U11416 (N_11416,N_10900,N_10849);
nor U11417 (N_11417,N_11063,N_10871);
and U11418 (N_11418,N_10972,N_10861);
and U11419 (N_11419,N_10979,N_10876);
xnor U11420 (N_11420,N_10920,N_11152);
and U11421 (N_11421,N_11085,N_11010);
and U11422 (N_11422,N_11007,N_10822);
nand U11423 (N_11423,N_10887,N_10824);
and U11424 (N_11424,N_10820,N_10995);
or U11425 (N_11425,N_10823,N_10849);
xnor U11426 (N_11426,N_10805,N_10950);
xnor U11427 (N_11427,N_10950,N_11042);
and U11428 (N_11428,N_11178,N_11124);
nor U11429 (N_11429,N_11112,N_10989);
and U11430 (N_11430,N_10819,N_11054);
or U11431 (N_11431,N_10910,N_10975);
nor U11432 (N_11432,N_11101,N_11157);
and U11433 (N_11433,N_11051,N_10991);
or U11434 (N_11434,N_10833,N_10884);
nor U11435 (N_11435,N_11055,N_11085);
and U11436 (N_11436,N_11181,N_10884);
nor U11437 (N_11437,N_10869,N_10801);
or U11438 (N_11438,N_11131,N_10947);
and U11439 (N_11439,N_10950,N_10872);
or U11440 (N_11440,N_11035,N_10963);
or U11441 (N_11441,N_11118,N_10927);
nor U11442 (N_11442,N_11052,N_10920);
nand U11443 (N_11443,N_10852,N_10924);
and U11444 (N_11444,N_10939,N_11081);
or U11445 (N_11445,N_11143,N_11171);
nor U11446 (N_11446,N_11192,N_11139);
nor U11447 (N_11447,N_10869,N_11119);
nor U11448 (N_11448,N_10991,N_11187);
or U11449 (N_11449,N_10846,N_10888);
nand U11450 (N_11450,N_10813,N_11078);
or U11451 (N_11451,N_11119,N_10873);
nand U11452 (N_11452,N_11177,N_11083);
or U11453 (N_11453,N_10946,N_11013);
and U11454 (N_11454,N_11043,N_11153);
xor U11455 (N_11455,N_10836,N_10938);
nand U11456 (N_11456,N_10821,N_11094);
nor U11457 (N_11457,N_11163,N_11141);
nor U11458 (N_11458,N_11064,N_11152);
nor U11459 (N_11459,N_10816,N_11029);
or U11460 (N_11460,N_10898,N_11121);
and U11461 (N_11461,N_10838,N_10904);
and U11462 (N_11462,N_11194,N_11139);
nor U11463 (N_11463,N_11134,N_10889);
xor U11464 (N_11464,N_10966,N_10804);
nor U11465 (N_11465,N_11158,N_10941);
nand U11466 (N_11466,N_11006,N_11144);
and U11467 (N_11467,N_11094,N_10921);
or U11468 (N_11468,N_11100,N_11052);
nor U11469 (N_11469,N_10995,N_11023);
and U11470 (N_11470,N_11093,N_10834);
nand U11471 (N_11471,N_11034,N_11004);
xor U11472 (N_11472,N_11182,N_10992);
nand U11473 (N_11473,N_11057,N_11147);
xnor U11474 (N_11474,N_11031,N_10926);
or U11475 (N_11475,N_11122,N_10823);
or U11476 (N_11476,N_10944,N_10825);
or U11477 (N_11477,N_10974,N_11190);
nand U11478 (N_11478,N_11035,N_10946);
nand U11479 (N_11479,N_10957,N_11107);
nand U11480 (N_11480,N_11040,N_10865);
nor U11481 (N_11481,N_11091,N_10884);
nand U11482 (N_11482,N_10930,N_11100);
or U11483 (N_11483,N_11118,N_11177);
xnor U11484 (N_11484,N_10873,N_10880);
and U11485 (N_11485,N_11130,N_11092);
or U11486 (N_11486,N_11108,N_10964);
nor U11487 (N_11487,N_11162,N_11091);
xor U11488 (N_11488,N_10927,N_11152);
nor U11489 (N_11489,N_11160,N_10891);
nand U11490 (N_11490,N_10983,N_11193);
or U11491 (N_11491,N_10944,N_11187);
or U11492 (N_11492,N_10885,N_10965);
or U11493 (N_11493,N_10874,N_11070);
nor U11494 (N_11494,N_10830,N_10804);
xor U11495 (N_11495,N_11003,N_10861);
and U11496 (N_11496,N_11083,N_10866);
or U11497 (N_11497,N_10921,N_10932);
nor U11498 (N_11498,N_10886,N_11190);
xor U11499 (N_11499,N_10824,N_11088);
nand U11500 (N_11500,N_10821,N_11043);
nand U11501 (N_11501,N_10978,N_10897);
nand U11502 (N_11502,N_10905,N_11003);
nand U11503 (N_11503,N_11077,N_10956);
nand U11504 (N_11504,N_11003,N_11040);
nor U11505 (N_11505,N_11018,N_11147);
and U11506 (N_11506,N_11001,N_10802);
nand U11507 (N_11507,N_11142,N_11077);
or U11508 (N_11508,N_11196,N_11162);
nor U11509 (N_11509,N_11069,N_11079);
nand U11510 (N_11510,N_10956,N_10959);
nand U11511 (N_11511,N_11129,N_10859);
or U11512 (N_11512,N_11063,N_10856);
or U11513 (N_11513,N_11120,N_11033);
or U11514 (N_11514,N_10863,N_11082);
xnor U11515 (N_11515,N_11048,N_11123);
and U11516 (N_11516,N_10886,N_11106);
nand U11517 (N_11517,N_11197,N_11075);
nand U11518 (N_11518,N_10902,N_11152);
or U11519 (N_11519,N_10901,N_10941);
xor U11520 (N_11520,N_10888,N_10942);
or U11521 (N_11521,N_11100,N_10863);
and U11522 (N_11522,N_10994,N_10876);
and U11523 (N_11523,N_11068,N_10888);
xor U11524 (N_11524,N_10853,N_10983);
nor U11525 (N_11525,N_10846,N_11102);
nor U11526 (N_11526,N_11138,N_11167);
or U11527 (N_11527,N_10861,N_10845);
or U11528 (N_11528,N_10864,N_11153);
nor U11529 (N_11529,N_11131,N_11190);
or U11530 (N_11530,N_10852,N_10869);
nand U11531 (N_11531,N_10879,N_10888);
nand U11532 (N_11532,N_11079,N_10964);
xor U11533 (N_11533,N_10870,N_11106);
xnor U11534 (N_11534,N_11083,N_11096);
or U11535 (N_11535,N_10828,N_10943);
nand U11536 (N_11536,N_11072,N_10941);
nand U11537 (N_11537,N_10919,N_11065);
xor U11538 (N_11538,N_10975,N_10926);
nor U11539 (N_11539,N_11113,N_10849);
nor U11540 (N_11540,N_10908,N_10973);
nor U11541 (N_11541,N_10963,N_11083);
or U11542 (N_11542,N_11078,N_10825);
nor U11543 (N_11543,N_11189,N_11192);
nor U11544 (N_11544,N_11075,N_11155);
and U11545 (N_11545,N_11032,N_10955);
nor U11546 (N_11546,N_10996,N_10845);
and U11547 (N_11547,N_10814,N_11067);
xor U11548 (N_11548,N_10818,N_10933);
or U11549 (N_11549,N_10930,N_11079);
nor U11550 (N_11550,N_10931,N_11184);
and U11551 (N_11551,N_11013,N_10842);
or U11552 (N_11552,N_11056,N_10825);
or U11553 (N_11553,N_10875,N_11081);
xnor U11554 (N_11554,N_10833,N_11046);
nor U11555 (N_11555,N_11120,N_10883);
and U11556 (N_11556,N_10876,N_10886);
nor U11557 (N_11557,N_10966,N_11060);
or U11558 (N_11558,N_10976,N_11118);
nor U11559 (N_11559,N_11162,N_11161);
nor U11560 (N_11560,N_11185,N_11176);
xor U11561 (N_11561,N_11178,N_11019);
and U11562 (N_11562,N_11081,N_10933);
nand U11563 (N_11563,N_11112,N_10827);
nand U11564 (N_11564,N_11163,N_10821);
and U11565 (N_11565,N_10841,N_11153);
or U11566 (N_11566,N_11020,N_11166);
or U11567 (N_11567,N_11187,N_11134);
and U11568 (N_11568,N_11155,N_10803);
nand U11569 (N_11569,N_11056,N_10926);
nor U11570 (N_11570,N_10936,N_10908);
xor U11571 (N_11571,N_11030,N_11185);
nor U11572 (N_11572,N_11135,N_11042);
xnor U11573 (N_11573,N_10899,N_10919);
and U11574 (N_11574,N_11149,N_10996);
nor U11575 (N_11575,N_11007,N_10802);
xnor U11576 (N_11576,N_11089,N_11142);
xor U11577 (N_11577,N_10996,N_10977);
xnor U11578 (N_11578,N_10956,N_11024);
and U11579 (N_11579,N_11118,N_11078);
nand U11580 (N_11580,N_11114,N_10921);
and U11581 (N_11581,N_11027,N_10879);
or U11582 (N_11582,N_10971,N_11188);
and U11583 (N_11583,N_10943,N_10903);
nand U11584 (N_11584,N_11144,N_10898);
and U11585 (N_11585,N_10976,N_11106);
or U11586 (N_11586,N_10852,N_11054);
or U11587 (N_11587,N_11186,N_11071);
xor U11588 (N_11588,N_10911,N_10963);
or U11589 (N_11589,N_10816,N_11001);
and U11590 (N_11590,N_11024,N_10841);
nor U11591 (N_11591,N_10892,N_11004);
and U11592 (N_11592,N_11161,N_10968);
and U11593 (N_11593,N_11180,N_10861);
or U11594 (N_11594,N_10977,N_10932);
and U11595 (N_11595,N_11189,N_11196);
nor U11596 (N_11596,N_10934,N_10979);
xnor U11597 (N_11597,N_11124,N_10933);
nor U11598 (N_11598,N_11035,N_11053);
nand U11599 (N_11599,N_11065,N_10923);
xnor U11600 (N_11600,N_11222,N_11578);
xor U11601 (N_11601,N_11372,N_11221);
and U11602 (N_11602,N_11486,N_11492);
nand U11603 (N_11603,N_11467,N_11510);
nor U11604 (N_11604,N_11526,N_11546);
xnor U11605 (N_11605,N_11333,N_11200);
and U11606 (N_11606,N_11208,N_11588);
xor U11607 (N_11607,N_11274,N_11584);
xor U11608 (N_11608,N_11566,N_11388);
and U11609 (N_11609,N_11214,N_11408);
or U11610 (N_11610,N_11521,N_11548);
and U11611 (N_11611,N_11480,N_11218);
and U11612 (N_11612,N_11284,N_11577);
nand U11613 (N_11613,N_11213,N_11359);
xor U11614 (N_11614,N_11361,N_11367);
and U11615 (N_11615,N_11565,N_11438);
nand U11616 (N_11616,N_11316,N_11471);
nor U11617 (N_11617,N_11369,N_11423);
nand U11618 (N_11618,N_11335,N_11580);
or U11619 (N_11619,N_11234,N_11466);
nor U11620 (N_11620,N_11394,N_11539);
and U11621 (N_11621,N_11528,N_11329);
or U11622 (N_11622,N_11445,N_11331);
nor U11623 (N_11623,N_11449,N_11468);
or U11624 (N_11624,N_11383,N_11243);
nor U11625 (N_11625,N_11490,N_11550);
nand U11626 (N_11626,N_11594,N_11227);
nand U11627 (N_11627,N_11502,N_11259);
nor U11628 (N_11628,N_11436,N_11235);
and U11629 (N_11629,N_11419,N_11231);
and U11630 (N_11630,N_11410,N_11322);
xor U11631 (N_11631,N_11413,N_11385);
nand U11632 (N_11632,N_11448,N_11389);
or U11633 (N_11633,N_11248,N_11533);
xnor U11634 (N_11634,N_11304,N_11292);
nor U11635 (N_11635,N_11344,N_11209);
or U11636 (N_11636,N_11277,N_11444);
or U11637 (N_11637,N_11576,N_11404);
and U11638 (N_11638,N_11430,N_11545);
and U11639 (N_11639,N_11543,N_11527);
and U11640 (N_11640,N_11593,N_11422);
nand U11641 (N_11641,N_11224,N_11400);
nor U11642 (N_11642,N_11523,N_11267);
and U11643 (N_11643,N_11461,N_11379);
nor U11644 (N_11644,N_11290,N_11247);
and U11645 (N_11645,N_11371,N_11441);
nor U11646 (N_11646,N_11559,N_11253);
nor U11647 (N_11647,N_11210,N_11348);
and U11648 (N_11648,N_11515,N_11206);
or U11649 (N_11649,N_11317,N_11555);
nand U11650 (N_11650,N_11479,N_11340);
nor U11651 (N_11651,N_11308,N_11332);
or U11652 (N_11652,N_11350,N_11249);
and U11653 (N_11653,N_11437,N_11525);
xor U11654 (N_11654,N_11431,N_11396);
nor U11655 (N_11655,N_11498,N_11399);
xor U11656 (N_11656,N_11226,N_11228);
and U11657 (N_11657,N_11244,N_11553);
nand U11658 (N_11658,N_11509,N_11428);
xor U11659 (N_11659,N_11382,N_11390);
nand U11660 (N_11660,N_11363,N_11517);
xnor U11661 (N_11661,N_11551,N_11263);
xnor U11662 (N_11662,N_11307,N_11564);
or U11663 (N_11663,N_11392,N_11387);
nor U11664 (N_11664,N_11567,N_11429);
nor U11665 (N_11665,N_11417,N_11421);
xnor U11666 (N_11666,N_11572,N_11531);
nand U11667 (N_11667,N_11241,N_11415);
nand U11668 (N_11668,N_11460,N_11301);
nor U11669 (N_11669,N_11395,N_11286);
and U11670 (N_11670,N_11411,N_11475);
nor U11671 (N_11671,N_11434,N_11465);
nand U11672 (N_11672,N_11268,N_11405);
nand U11673 (N_11673,N_11416,N_11433);
and U11674 (N_11674,N_11435,N_11477);
nand U11675 (N_11675,N_11570,N_11450);
nand U11676 (N_11676,N_11314,N_11522);
nor U11677 (N_11677,N_11534,N_11302);
and U11678 (N_11678,N_11356,N_11542);
xnor U11679 (N_11679,N_11452,N_11457);
nor U11680 (N_11680,N_11325,N_11571);
xnor U11681 (N_11681,N_11455,N_11575);
and U11682 (N_11682,N_11473,N_11380);
nor U11683 (N_11683,N_11552,N_11326);
xor U11684 (N_11684,N_11362,N_11532);
nor U11685 (N_11685,N_11512,N_11454);
nor U11686 (N_11686,N_11251,N_11469);
nor U11687 (N_11687,N_11425,N_11557);
and U11688 (N_11688,N_11544,N_11393);
xor U11689 (N_11689,N_11318,N_11530);
nand U11690 (N_11690,N_11412,N_11586);
or U11691 (N_11691,N_11260,N_11403);
nor U11692 (N_11692,N_11491,N_11484);
nand U11693 (N_11693,N_11289,N_11319);
nand U11694 (N_11694,N_11511,N_11574);
nor U11695 (N_11695,N_11494,N_11309);
nor U11696 (N_11696,N_11245,N_11300);
or U11697 (N_11697,N_11352,N_11269);
and U11698 (N_11698,N_11374,N_11589);
or U11699 (N_11699,N_11424,N_11513);
nand U11700 (N_11700,N_11398,N_11556);
xnor U11701 (N_11701,N_11500,N_11219);
nand U11702 (N_11702,N_11489,N_11229);
nand U11703 (N_11703,N_11323,N_11585);
xor U11704 (N_11704,N_11485,N_11558);
nand U11705 (N_11705,N_11217,N_11560);
xnor U11706 (N_11706,N_11474,N_11216);
nand U11707 (N_11707,N_11265,N_11418);
or U11708 (N_11708,N_11347,N_11339);
or U11709 (N_11709,N_11293,N_11296);
or U11710 (N_11710,N_11481,N_11569);
nor U11711 (N_11711,N_11598,N_11368);
xor U11712 (N_11712,N_11375,N_11257);
nor U11713 (N_11713,N_11239,N_11328);
nand U11714 (N_11714,N_11281,N_11282);
nand U11715 (N_11715,N_11495,N_11355);
xor U11716 (N_11716,N_11414,N_11358);
xor U11717 (N_11717,N_11581,N_11201);
xnor U11718 (N_11718,N_11298,N_11315);
nand U11719 (N_11719,N_11327,N_11261);
and U11720 (N_11720,N_11223,N_11204);
nor U11721 (N_11721,N_11205,N_11202);
or U11722 (N_11722,N_11288,N_11280);
nand U11723 (N_11723,N_11295,N_11391);
nor U11724 (N_11724,N_11285,N_11233);
nand U11725 (N_11725,N_11346,N_11341);
xor U11726 (N_11726,N_11464,N_11587);
xnor U11727 (N_11727,N_11518,N_11312);
and U11728 (N_11728,N_11562,N_11272);
nand U11729 (N_11729,N_11357,N_11462);
or U11730 (N_11730,N_11520,N_11561);
xor U11731 (N_11731,N_11456,N_11573);
nand U11732 (N_11732,N_11493,N_11440);
xor U11733 (N_11733,N_11255,N_11264);
xor U11734 (N_11734,N_11351,N_11488);
xor U11735 (N_11735,N_11311,N_11386);
nand U11736 (N_11736,N_11426,N_11501);
nand U11737 (N_11737,N_11366,N_11225);
or U11738 (N_11738,N_11294,N_11409);
and U11739 (N_11739,N_11373,N_11563);
xnor U11740 (N_11740,N_11483,N_11353);
or U11741 (N_11741,N_11376,N_11443);
and U11742 (N_11742,N_11271,N_11478);
xnor U11743 (N_11743,N_11299,N_11338);
xnor U11744 (N_11744,N_11275,N_11579);
or U11745 (N_11745,N_11591,N_11303);
xnor U11746 (N_11746,N_11583,N_11207);
nand U11747 (N_11747,N_11279,N_11599);
xnor U11748 (N_11748,N_11597,N_11273);
or U11749 (N_11749,N_11401,N_11212);
nand U11750 (N_11750,N_11453,N_11549);
xor U11751 (N_11751,N_11291,N_11305);
xor U11752 (N_11752,N_11506,N_11536);
or U11753 (N_11753,N_11497,N_11370);
or U11754 (N_11754,N_11297,N_11378);
nand U11755 (N_11755,N_11278,N_11582);
xnor U11756 (N_11756,N_11321,N_11310);
xor U11757 (N_11757,N_11236,N_11343);
nand U11758 (N_11758,N_11406,N_11215);
nand U11759 (N_11759,N_11258,N_11407);
nand U11760 (N_11760,N_11220,N_11287);
or U11761 (N_11761,N_11342,N_11540);
or U11762 (N_11762,N_11592,N_11320);
or U11763 (N_11763,N_11472,N_11313);
xnor U11764 (N_11764,N_11337,N_11504);
or U11765 (N_11765,N_11237,N_11487);
nor U11766 (N_11766,N_11330,N_11254);
or U11767 (N_11767,N_11324,N_11252);
xor U11768 (N_11768,N_11503,N_11496);
nand U11769 (N_11769,N_11427,N_11334);
nand U11770 (N_11770,N_11349,N_11365);
xor U11771 (N_11771,N_11538,N_11442);
xnor U11772 (N_11772,N_11519,N_11508);
nand U11773 (N_11773,N_11240,N_11381);
and U11774 (N_11774,N_11439,N_11451);
and U11775 (N_11775,N_11507,N_11541);
or U11776 (N_11776,N_11232,N_11596);
and U11777 (N_11777,N_11432,N_11537);
nor U11778 (N_11778,N_11470,N_11246);
or U11779 (N_11779,N_11458,N_11595);
nand U11780 (N_11780,N_11238,N_11364);
or U11781 (N_11781,N_11402,N_11529);
and U11782 (N_11782,N_11250,N_11384);
nor U11783 (N_11783,N_11516,N_11211);
nand U11784 (N_11784,N_11459,N_11499);
nand U11785 (N_11785,N_11446,N_11270);
or U11786 (N_11786,N_11360,N_11524);
or U11787 (N_11787,N_11354,N_11377);
and U11788 (N_11788,N_11547,N_11283);
nand U11789 (N_11789,N_11420,N_11262);
or U11790 (N_11790,N_11568,N_11447);
nand U11791 (N_11791,N_11554,N_11203);
xnor U11792 (N_11792,N_11397,N_11590);
nor U11793 (N_11793,N_11463,N_11505);
xnor U11794 (N_11794,N_11345,N_11336);
nor U11795 (N_11795,N_11535,N_11256);
and U11796 (N_11796,N_11482,N_11276);
xor U11797 (N_11797,N_11476,N_11266);
or U11798 (N_11798,N_11230,N_11514);
nor U11799 (N_11799,N_11306,N_11242);
and U11800 (N_11800,N_11403,N_11490);
xor U11801 (N_11801,N_11332,N_11303);
or U11802 (N_11802,N_11540,N_11310);
and U11803 (N_11803,N_11474,N_11254);
nor U11804 (N_11804,N_11385,N_11461);
xor U11805 (N_11805,N_11308,N_11514);
nor U11806 (N_11806,N_11394,N_11423);
xnor U11807 (N_11807,N_11352,N_11239);
nand U11808 (N_11808,N_11248,N_11508);
nand U11809 (N_11809,N_11284,N_11227);
and U11810 (N_11810,N_11201,N_11406);
xor U11811 (N_11811,N_11583,N_11562);
nor U11812 (N_11812,N_11263,N_11462);
nor U11813 (N_11813,N_11450,N_11515);
and U11814 (N_11814,N_11447,N_11229);
and U11815 (N_11815,N_11203,N_11252);
nor U11816 (N_11816,N_11353,N_11282);
and U11817 (N_11817,N_11542,N_11308);
xor U11818 (N_11818,N_11450,N_11349);
nor U11819 (N_11819,N_11285,N_11407);
nand U11820 (N_11820,N_11214,N_11279);
nand U11821 (N_11821,N_11251,N_11579);
nand U11822 (N_11822,N_11504,N_11401);
or U11823 (N_11823,N_11481,N_11267);
nor U11824 (N_11824,N_11415,N_11277);
xor U11825 (N_11825,N_11394,N_11264);
xnor U11826 (N_11826,N_11222,N_11506);
or U11827 (N_11827,N_11257,N_11215);
or U11828 (N_11828,N_11415,N_11515);
nand U11829 (N_11829,N_11408,N_11244);
xnor U11830 (N_11830,N_11226,N_11430);
xnor U11831 (N_11831,N_11448,N_11599);
nor U11832 (N_11832,N_11295,N_11270);
or U11833 (N_11833,N_11227,N_11462);
nor U11834 (N_11834,N_11312,N_11381);
nand U11835 (N_11835,N_11384,N_11349);
xnor U11836 (N_11836,N_11451,N_11262);
and U11837 (N_11837,N_11500,N_11329);
xnor U11838 (N_11838,N_11557,N_11597);
xnor U11839 (N_11839,N_11366,N_11244);
or U11840 (N_11840,N_11293,N_11528);
and U11841 (N_11841,N_11496,N_11439);
or U11842 (N_11842,N_11212,N_11306);
or U11843 (N_11843,N_11483,N_11331);
or U11844 (N_11844,N_11229,N_11390);
nor U11845 (N_11845,N_11499,N_11218);
xnor U11846 (N_11846,N_11401,N_11391);
nor U11847 (N_11847,N_11445,N_11243);
and U11848 (N_11848,N_11499,N_11537);
or U11849 (N_11849,N_11248,N_11294);
nand U11850 (N_11850,N_11382,N_11234);
and U11851 (N_11851,N_11397,N_11484);
or U11852 (N_11852,N_11297,N_11238);
nor U11853 (N_11853,N_11439,N_11547);
nor U11854 (N_11854,N_11458,N_11363);
or U11855 (N_11855,N_11511,N_11330);
and U11856 (N_11856,N_11298,N_11454);
xor U11857 (N_11857,N_11585,N_11502);
nand U11858 (N_11858,N_11272,N_11317);
nor U11859 (N_11859,N_11525,N_11234);
or U11860 (N_11860,N_11292,N_11487);
xor U11861 (N_11861,N_11483,N_11574);
nor U11862 (N_11862,N_11326,N_11444);
nor U11863 (N_11863,N_11575,N_11261);
xnor U11864 (N_11864,N_11484,N_11243);
xor U11865 (N_11865,N_11299,N_11215);
xnor U11866 (N_11866,N_11592,N_11246);
nor U11867 (N_11867,N_11572,N_11399);
and U11868 (N_11868,N_11410,N_11390);
nor U11869 (N_11869,N_11460,N_11544);
and U11870 (N_11870,N_11565,N_11470);
nand U11871 (N_11871,N_11599,N_11347);
nor U11872 (N_11872,N_11528,N_11500);
or U11873 (N_11873,N_11583,N_11227);
nor U11874 (N_11874,N_11490,N_11301);
nand U11875 (N_11875,N_11336,N_11264);
and U11876 (N_11876,N_11231,N_11217);
nand U11877 (N_11877,N_11593,N_11549);
or U11878 (N_11878,N_11368,N_11388);
and U11879 (N_11879,N_11359,N_11550);
and U11880 (N_11880,N_11355,N_11243);
or U11881 (N_11881,N_11204,N_11455);
nor U11882 (N_11882,N_11250,N_11540);
xnor U11883 (N_11883,N_11592,N_11284);
nor U11884 (N_11884,N_11554,N_11265);
nor U11885 (N_11885,N_11498,N_11458);
xor U11886 (N_11886,N_11561,N_11224);
or U11887 (N_11887,N_11298,N_11209);
or U11888 (N_11888,N_11302,N_11482);
or U11889 (N_11889,N_11269,N_11393);
nand U11890 (N_11890,N_11407,N_11265);
and U11891 (N_11891,N_11566,N_11296);
and U11892 (N_11892,N_11594,N_11252);
and U11893 (N_11893,N_11567,N_11471);
xnor U11894 (N_11894,N_11320,N_11597);
and U11895 (N_11895,N_11543,N_11489);
xor U11896 (N_11896,N_11237,N_11463);
and U11897 (N_11897,N_11360,N_11435);
nand U11898 (N_11898,N_11572,N_11419);
nor U11899 (N_11899,N_11326,N_11465);
and U11900 (N_11900,N_11450,N_11563);
nand U11901 (N_11901,N_11563,N_11530);
or U11902 (N_11902,N_11375,N_11579);
and U11903 (N_11903,N_11550,N_11533);
and U11904 (N_11904,N_11589,N_11411);
xnor U11905 (N_11905,N_11381,N_11253);
or U11906 (N_11906,N_11403,N_11373);
nand U11907 (N_11907,N_11346,N_11304);
and U11908 (N_11908,N_11486,N_11226);
and U11909 (N_11909,N_11521,N_11300);
nand U11910 (N_11910,N_11260,N_11385);
and U11911 (N_11911,N_11477,N_11536);
or U11912 (N_11912,N_11549,N_11382);
nor U11913 (N_11913,N_11270,N_11271);
nor U11914 (N_11914,N_11346,N_11585);
or U11915 (N_11915,N_11395,N_11319);
xor U11916 (N_11916,N_11417,N_11230);
or U11917 (N_11917,N_11287,N_11572);
nand U11918 (N_11918,N_11504,N_11362);
nor U11919 (N_11919,N_11340,N_11391);
nand U11920 (N_11920,N_11313,N_11273);
and U11921 (N_11921,N_11512,N_11451);
nor U11922 (N_11922,N_11296,N_11256);
or U11923 (N_11923,N_11251,N_11471);
nor U11924 (N_11924,N_11361,N_11436);
and U11925 (N_11925,N_11388,N_11296);
xor U11926 (N_11926,N_11267,N_11379);
xor U11927 (N_11927,N_11388,N_11593);
nor U11928 (N_11928,N_11330,N_11322);
nor U11929 (N_11929,N_11272,N_11462);
or U11930 (N_11930,N_11409,N_11291);
nor U11931 (N_11931,N_11302,N_11546);
xnor U11932 (N_11932,N_11580,N_11589);
nand U11933 (N_11933,N_11230,N_11299);
nand U11934 (N_11934,N_11311,N_11456);
and U11935 (N_11935,N_11353,N_11508);
nor U11936 (N_11936,N_11471,N_11411);
nor U11937 (N_11937,N_11233,N_11333);
nor U11938 (N_11938,N_11519,N_11261);
xor U11939 (N_11939,N_11466,N_11586);
and U11940 (N_11940,N_11525,N_11562);
xnor U11941 (N_11941,N_11419,N_11584);
nand U11942 (N_11942,N_11278,N_11405);
nand U11943 (N_11943,N_11597,N_11237);
nor U11944 (N_11944,N_11267,N_11521);
nor U11945 (N_11945,N_11473,N_11498);
and U11946 (N_11946,N_11552,N_11573);
nand U11947 (N_11947,N_11576,N_11231);
or U11948 (N_11948,N_11370,N_11572);
and U11949 (N_11949,N_11386,N_11265);
and U11950 (N_11950,N_11497,N_11277);
xnor U11951 (N_11951,N_11282,N_11521);
nand U11952 (N_11952,N_11295,N_11253);
and U11953 (N_11953,N_11542,N_11296);
nor U11954 (N_11954,N_11448,N_11257);
nor U11955 (N_11955,N_11433,N_11335);
or U11956 (N_11956,N_11270,N_11418);
or U11957 (N_11957,N_11346,N_11397);
nand U11958 (N_11958,N_11330,N_11348);
or U11959 (N_11959,N_11422,N_11455);
nor U11960 (N_11960,N_11559,N_11392);
xnor U11961 (N_11961,N_11201,N_11208);
nand U11962 (N_11962,N_11314,N_11533);
xor U11963 (N_11963,N_11478,N_11438);
xnor U11964 (N_11964,N_11208,N_11304);
or U11965 (N_11965,N_11213,N_11350);
nor U11966 (N_11966,N_11244,N_11236);
and U11967 (N_11967,N_11332,N_11444);
or U11968 (N_11968,N_11270,N_11537);
xor U11969 (N_11969,N_11259,N_11509);
nor U11970 (N_11970,N_11233,N_11266);
nand U11971 (N_11971,N_11305,N_11557);
xor U11972 (N_11972,N_11221,N_11454);
or U11973 (N_11973,N_11515,N_11487);
nor U11974 (N_11974,N_11563,N_11568);
nand U11975 (N_11975,N_11331,N_11309);
nand U11976 (N_11976,N_11276,N_11319);
and U11977 (N_11977,N_11234,N_11509);
and U11978 (N_11978,N_11565,N_11365);
nor U11979 (N_11979,N_11283,N_11237);
or U11980 (N_11980,N_11508,N_11242);
and U11981 (N_11981,N_11348,N_11338);
and U11982 (N_11982,N_11337,N_11446);
or U11983 (N_11983,N_11260,N_11413);
xnor U11984 (N_11984,N_11505,N_11557);
xor U11985 (N_11985,N_11491,N_11524);
and U11986 (N_11986,N_11237,N_11312);
or U11987 (N_11987,N_11481,N_11407);
nor U11988 (N_11988,N_11431,N_11291);
nand U11989 (N_11989,N_11524,N_11388);
nor U11990 (N_11990,N_11529,N_11449);
xnor U11991 (N_11991,N_11513,N_11435);
and U11992 (N_11992,N_11238,N_11373);
xnor U11993 (N_11993,N_11382,N_11539);
or U11994 (N_11994,N_11491,N_11257);
xor U11995 (N_11995,N_11516,N_11295);
nand U11996 (N_11996,N_11249,N_11344);
nor U11997 (N_11997,N_11212,N_11567);
or U11998 (N_11998,N_11488,N_11292);
nand U11999 (N_11999,N_11333,N_11407);
nand U12000 (N_12000,N_11838,N_11723);
xnor U12001 (N_12001,N_11703,N_11681);
and U12002 (N_12002,N_11721,N_11618);
xnor U12003 (N_12003,N_11648,N_11919);
nand U12004 (N_12004,N_11988,N_11717);
or U12005 (N_12005,N_11792,N_11659);
nor U12006 (N_12006,N_11674,N_11960);
nand U12007 (N_12007,N_11977,N_11600);
nand U12008 (N_12008,N_11900,N_11682);
nor U12009 (N_12009,N_11661,N_11733);
xor U12010 (N_12010,N_11821,N_11641);
nand U12011 (N_12011,N_11754,N_11625);
or U12012 (N_12012,N_11958,N_11795);
nor U12013 (N_12013,N_11980,N_11999);
nor U12014 (N_12014,N_11832,N_11653);
nor U12015 (N_12015,N_11780,N_11987);
or U12016 (N_12016,N_11727,N_11891);
xor U12017 (N_12017,N_11956,N_11728);
nand U12018 (N_12018,N_11679,N_11798);
and U12019 (N_12019,N_11668,N_11881);
or U12020 (N_12020,N_11730,N_11797);
or U12021 (N_12021,N_11812,N_11862);
and U12022 (N_12022,N_11697,N_11803);
and U12023 (N_12023,N_11811,N_11612);
xnor U12024 (N_12024,N_11870,N_11745);
nand U12025 (N_12025,N_11722,N_11781);
xnor U12026 (N_12026,N_11864,N_11649);
xnor U12027 (N_12027,N_11757,N_11732);
xor U12028 (N_12028,N_11946,N_11741);
or U12029 (N_12029,N_11913,N_11859);
nor U12030 (N_12030,N_11850,N_11950);
xor U12031 (N_12031,N_11675,N_11710);
nor U12032 (N_12032,N_11607,N_11922);
xnor U12033 (N_12033,N_11673,N_11655);
or U12034 (N_12034,N_11963,N_11790);
xnor U12035 (N_12035,N_11796,N_11689);
and U12036 (N_12036,N_11845,N_11925);
or U12037 (N_12037,N_11662,N_11895);
and U12038 (N_12038,N_11942,N_11753);
nor U12039 (N_12039,N_11635,N_11606);
nor U12040 (N_12040,N_11636,N_11678);
xnor U12041 (N_12041,N_11914,N_11983);
nand U12042 (N_12042,N_11973,N_11769);
or U12043 (N_12043,N_11959,N_11844);
xor U12044 (N_12044,N_11670,N_11885);
nand U12045 (N_12045,N_11691,N_11755);
xnor U12046 (N_12046,N_11667,N_11645);
xnor U12047 (N_12047,N_11970,N_11601);
xor U12048 (N_12048,N_11837,N_11809);
nor U12049 (N_12049,N_11647,N_11929);
xnor U12050 (N_12050,N_11897,N_11948);
xnor U12051 (N_12051,N_11715,N_11969);
xnor U12052 (N_12052,N_11957,N_11768);
and U12053 (N_12053,N_11773,N_11704);
and U12054 (N_12054,N_11737,N_11799);
nand U12055 (N_12055,N_11979,N_11941);
or U12056 (N_12056,N_11813,N_11990);
nand U12057 (N_12057,N_11763,N_11751);
and U12058 (N_12058,N_11971,N_11991);
or U12059 (N_12059,N_11716,N_11713);
nor U12060 (N_12060,N_11793,N_11714);
nor U12061 (N_12061,N_11924,N_11967);
xor U12062 (N_12062,N_11756,N_11794);
and U12063 (N_12063,N_11605,N_11752);
nand U12064 (N_12064,N_11746,N_11829);
or U12065 (N_12065,N_11886,N_11677);
nand U12066 (N_12066,N_11731,N_11939);
xor U12067 (N_12067,N_11921,N_11724);
xnor U12068 (N_12068,N_11616,N_11611);
nor U12069 (N_12069,N_11863,N_11861);
xor U12070 (N_12070,N_11726,N_11962);
nand U12071 (N_12071,N_11966,N_11742);
xnor U12072 (N_12072,N_11857,N_11765);
xor U12073 (N_12073,N_11748,N_11938);
or U12074 (N_12074,N_11855,N_11986);
nand U12075 (N_12075,N_11693,N_11774);
nand U12076 (N_12076,N_11851,N_11627);
nand U12077 (N_12077,N_11676,N_11998);
nand U12078 (N_12078,N_11631,N_11981);
nand U12079 (N_12079,N_11909,N_11712);
and U12080 (N_12080,N_11615,N_11603);
nand U12081 (N_12081,N_11873,N_11906);
nor U12082 (N_12082,N_11978,N_11974);
or U12083 (N_12083,N_11869,N_11623);
or U12084 (N_12084,N_11652,N_11935);
nand U12085 (N_12085,N_11918,N_11690);
and U12086 (N_12086,N_11894,N_11638);
nor U12087 (N_12087,N_11608,N_11672);
nand U12088 (N_12088,N_11776,N_11660);
and U12089 (N_12089,N_11740,N_11688);
and U12090 (N_12090,N_11878,N_11833);
xnor U12091 (N_12091,N_11734,N_11743);
or U12092 (N_12092,N_11617,N_11646);
nor U12093 (N_12093,N_11802,N_11854);
or U12094 (N_12094,N_11828,N_11898);
xnor U12095 (N_12095,N_11739,N_11815);
nor U12096 (N_12096,N_11788,N_11842);
nor U12097 (N_12097,N_11666,N_11772);
xnor U12098 (N_12098,N_11849,N_11830);
xnor U12099 (N_12099,N_11985,N_11926);
and U12100 (N_12100,N_11917,N_11620);
and U12101 (N_12101,N_11887,N_11778);
and U12102 (N_12102,N_11651,N_11902);
and U12103 (N_12103,N_11928,N_11949);
xnor U12104 (N_12104,N_11867,N_11968);
xor U12105 (N_12105,N_11718,N_11656);
and U12106 (N_12106,N_11705,N_11927);
nand U12107 (N_12107,N_11910,N_11791);
or U12108 (N_12108,N_11684,N_11953);
xnor U12109 (N_12109,N_11901,N_11642);
nand U12110 (N_12110,N_11884,N_11860);
nand U12111 (N_12111,N_11804,N_11976);
nand U12112 (N_12112,N_11916,N_11801);
and U12113 (N_12113,N_11945,N_11955);
nand U12114 (N_12114,N_11643,N_11671);
nand U12115 (N_12115,N_11633,N_11852);
and U12116 (N_12116,N_11896,N_11800);
nand U12117 (N_12117,N_11984,N_11814);
and U12118 (N_12118,N_11709,N_11808);
or U12119 (N_12119,N_11997,N_11771);
xnor U12120 (N_12120,N_11747,N_11858);
xor U12121 (N_12121,N_11698,N_11882);
xnor U12122 (N_12122,N_11706,N_11818);
or U12123 (N_12123,N_11729,N_11604);
or U12124 (N_12124,N_11911,N_11629);
nand U12125 (N_12125,N_11866,N_11915);
nand U12126 (N_12126,N_11719,N_11836);
or U12127 (N_12127,N_11784,N_11764);
nand U12128 (N_12128,N_11687,N_11694);
and U12129 (N_12129,N_11750,N_11904);
or U12130 (N_12130,N_11626,N_11826);
nor U12131 (N_12131,N_11879,N_11680);
nor U12132 (N_12132,N_11965,N_11699);
nor U12133 (N_12133,N_11868,N_11890);
xor U12134 (N_12134,N_11657,N_11664);
and U12135 (N_12135,N_11806,N_11923);
or U12136 (N_12136,N_11669,N_11903);
nand U12137 (N_12137,N_11760,N_11759);
nand U12138 (N_12138,N_11936,N_11650);
or U12139 (N_12139,N_11841,N_11665);
or U12140 (N_12140,N_11692,N_11619);
or U12141 (N_12141,N_11943,N_11920);
nor U12142 (N_12142,N_11735,N_11761);
nand U12143 (N_12143,N_11634,N_11762);
nand U12144 (N_12144,N_11610,N_11621);
xnor U12145 (N_12145,N_11865,N_11810);
xnor U12146 (N_12146,N_11964,N_11933);
xnor U12147 (N_12147,N_11622,N_11785);
nand U12148 (N_12148,N_11695,N_11930);
xnor U12149 (N_12149,N_11874,N_11834);
nand U12150 (N_12150,N_11817,N_11843);
or U12151 (N_12151,N_11972,N_11807);
nand U12152 (N_12152,N_11663,N_11877);
nor U12153 (N_12153,N_11982,N_11995);
xnor U12154 (N_12154,N_11839,N_11816);
or U12155 (N_12155,N_11853,N_11934);
nor U12156 (N_12156,N_11823,N_11848);
nand U12157 (N_12157,N_11614,N_11912);
xor U12158 (N_12158,N_11872,N_11820);
xnor U12159 (N_12159,N_11613,N_11822);
nand U12160 (N_12160,N_11947,N_11686);
or U12161 (N_12161,N_11779,N_11944);
nor U12162 (N_12162,N_11954,N_11892);
and U12163 (N_12163,N_11951,N_11871);
or U12164 (N_12164,N_11707,N_11883);
or U12165 (N_12165,N_11819,N_11893);
nor U12166 (N_12166,N_11840,N_11630);
and U12167 (N_12167,N_11696,N_11628);
xor U12168 (N_12168,N_11789,N_11993);
nor U12169 (N_12169,N_11766,N_11783);
or U12170 (N_12170,N_11989,N_11758);
nor U12171 (N_12171,N_11787,N_11846);
or U12172 (N_12172,N_11637,N_11700);
or U12173 (N_12173,N_11711,N_11888);
nor U12174 (N_12174,N_11708,N_11624);
nor U12175 (N_12175,N_11889,N_11876);
nor U12176 (N_12176,N_11825,N_11880);
nor U12177 (N_12177,N_11952,N_11786);
nor U12178 (N_12178,N_11905,N_11899);
nor U12179 (N_12179,N_11736,N_11775);
and U12180 (N_12180,N_11658,N_11831);
nor U12181 (N_12181,N_11940,N_11609);
nor U12182 (N_12182,N_11961,N_11701);
nand U12183 (N_12183,N_11937,N_11685);
nand U12184 (N_12184,N_11847,N_11805);
nor U12185 (N_12185,N_11639,N_11749);
nor U12186 (N_12186,N_11640,N_11770);
and U12187 (N_12187,N_11702,N_11644);
xnor U12188 (N_12188,N_11992,N_11996);
nor U12189 (N_12189,N_11994,N_11908);
nand U12190 (N_12190,N_11975,N_11725);
xor U12191 (N_12191,N_11931,N_11720);
xnor U12192 (N_12192,N_11827,N_11654);
nand U12193 (N_12193,N_11767,N_11782);
and U12194 (N_12194,N_11744,N_11907);
and U12195 (N_12195,N_11932,N_11602);
nand U12196 (N_12196,N_11738,N_11777);
nand U12197 (N_12197,N_11824,N_11856);
nor U12198 (N_12198,N_11875,N_11632);
nand U12199 (N_12199,N_11683,N_11835);
and U12200 (N_12200,N_11950,N_11608);
xor U12201 (N_12201,N_11985,N_11992);
or U12202 (N_12202,N_11957,N_11911);
xnor U12203 (N_12203,N_11948,N_11818);
nor U12204 (N_12204,N_11693,N_11796);
xor U12205 (N_12205,N_11870,N_11775);
and U12206 (N_12206,N_11654,N_11961);
and U12207 (N_12207,N_11737,N_11603);
or U12208 (N_12208,N_11918,N_11803);
nand U12209 (N_12209,N_11739,N_11805);
nand U12210 (N_12210,N_11939,N_11852);
and U12211 (N_12211,N_11997,N_11947);
nand U12212 (N_12212,N_11921,N_11910);
nand U12213 (N_12213,N_11858,N_11895);
xor U12214 (N_12214,N_11728,N_11776);
and U12215 (N_12215,N_11786,N_11668);
and U12216 (N_12216,N_11897,N_11699);
and U12217 (N_12217,N_11923,N_11953);
or U12218 (N_12218,N_11786,N_11891);
or U12219 (N_12219,N_11755,N_11721);
nand U12220 (N_12220,N_11726,N_11602);
or U12221 (N_12221,N_11666,N_11880);
or U12222 (N_12222,N_11835,N_11938);
xnor U12223 (N_12223,N_11864,N_11623);
nor U12224 (N_12224,N_11744,N_11619);
or U12225 (N_12225,N_11890,N_11836);
xnor U12226 (N_12226,N_11781,N_11646);
nor U12227 (N_12227,N_11735,N_11767);
nor U12228 (N_12228,N_11962,N_11868);
nor U12229 (N_12229,N_11943,N_11627);
xor U12230 (N_12230,N_11981,N_11782);
nand U12231 (N_12231,N_11658,N_11827);
or U12232 (N_12232,N_11619,N_11972);
or U12233 (N_12233,N_11612,N_11716);
nand U12234 (N_12234,N_11834,N_11770);
nand U12235 (N_12235,N_11642,N_11654);
nand U12236 (N_12236,N_11847,N_11817);
xnor U12237 (N_12237,N_11945,N_11932);
nand U12238 (N_12238,N_11753,N_11840);
nand U12239 (N_12239,N_11804,N_11617);
xor U12240 (N_12240,N_11830,N_11814);
xnor U12241 (N_12241,N_11616,N_11767);
or U12242 (N_12242,N_11705,N_11973);
xor U12243 (N_12243,N_11779,N_11984);
or U12244 (N_12244,N_11864,N_11660);
or U12245 (N_12245,N_11983,N_11836);
nand U12246 (N_12246,N_11975,N_11886);
nor U12247 (N_12247,N_11602,N_11977);
nand U12248 (N_12248,N_11901,N_11967);
xnor U12249 (N_12249,N_11799,N_11925);
xnor U12250 (N_12250,N_11724,N_11905);
nand U12251 (N_12251,N_11842,N_11827);
nor U12252 (N_12252,N_11890,N_11947);
and U12253 (N_12253,N_11894,N_11754);
nand U12254 (N_12254,N_11945,N_11870);
xnor U12255 (N_12255,N_11793,N_11695);
and U12256 (N_12256,N_11876,N_11948);
and U12257 (N_12257,N_11615,N_11793);
and U12258 (N_12258,N_11855,N_11702);
and U12259 (N_12259,N_11825,N_11738);
nor U12260 (N_12260,N_11810,N_11914);
and U12261 (N_12261,N_11984,N_11880);
nand U12262 (N_12262,N_11973,N_11979);
and U12263 (N_12263,N_11755,N_11889);
nor U12264 (N_12264,N_11983,N_11859);
nor U12265 (N_12265,N_11617,N_11951);
or U12266 (N_12266,N_11942,N_11813);
xor U12267 (N_12267,N_11669,N_11601);
and U12268 (N_12268,N_11817,N_11614);
nor U12269 (N_12269,N_11856,N_11790);
nand U12270 (N_12270,N_11941,N_11949);
xnor U12271 (N_12271,N_11999,N_11620);
or U12272 (N_12272,N_11732,N_11633);
and U12273 (N_12273,N_11752,N_11837);
and U12274 (N_12274,N_11952,N_11767);
and U12275 (N_12275,N_11857,N_11934);
and U12276 (N_12276,N_11647,N_11809);
and U12277 (N_12277,N_11933,N_11693);
nand U12278 (N_12278,N_11927,N_11930);
nand U12279 (N_12279,N_11860,N_11783);
and U12280 (N_12280,N_11967,N_11912);
or U12281 (N_12281,N_11731,N_11615);
nand U12282 (N_12282,N_11934,N_11684);
nand U12283 (N_12283,N_11818,N_11787);
and U12284 (N_12284,N_11641,N_11926);
xor U12285 (N_12285,N_11813,N_11850);
xor U12286 (N_12286,N_11666,N_11623);
nor U12287 (N_12287,N_11782,N_11891);
xnor U12288 (N_12288,N_11731,N_11612);
xor U12289 (N_12289,N_11662,N_11783);
nor U12290 (N_12290,N_11780,N_11718);
nor U12291 (N_12291,N_11899,N_11660);
nand U12292 (N_12292,N_11636,N_11915);
or U12293 (N_12293,N_11838,N_11971);
nor U12294 (N_12294,N_11873,N_11645);
nand U12295 (N_12295,N_11856,N_11627);
and U12296 (N_12296,N_11830,N_11845);
or U12297 (N_12297,N_11990,N_11654);
or U12298 (N_12298,N_11823,N_11888);
xnor U12299 (N_12299,N_11748,N_11954);
or U12300 (N_12300,N_11784,N_11661);
and U12301 (N_12301,N_11957,N_11802);
nor U12302 (N_12302,N_11722,N_11751);
and U12303 (N_12303,N_11791,N_11960);
and U12304 (N_12304,N_11745,N_11851);
nand U12305 (N_12305,N_11793,N_11994);
and U12306 (N_12306,N_11954,N_11833);
or U12307 (N_12307,N_11825,N_11646);
and U12308 (N_12308,N_11770,N_11942);
xnor U12309 (N_12309,N_11941,N_11733);
nor U12310 (N_12310,N_11904,N_11601);
nor U12311 (N_12311,N_11780,N_11954);
nor U12312 (N_12312,N_11886,N_11957);
or U12313 (N_12313,N_11845,N_11836);
xnor U12314 (N_12314,N_11767,N_11763);
and U12315 (N_12315,N_11704,N_11734);
or U12316 (N_12316,N_11680,N_11960);
and U12317 (N_12317,N_11629,N_11762);
and U12318 (N_12318,N_11774,N_11785);
and U12319 (N_12319,N_11886,N_11611);
nor U12320 (N_12320,N_11706,N_11698);
nor U12321 (N_12321,N_11707,N_11972);
or U12322 (N_12322,N_11651,N_11837);
nand U12323 (N_12323,N_11631,N_11833);
and U12324 (N_12324,N_11956,N_11752);
and U12325 (N_12325,N_11718,N_11805);
nand U12326 (N_12326,N_11655,N_11897);
xor U12327 (N_12327,N_11830,N_11971);
nand U12328 (N_12328,N_11961,N_11662);
nand U12329 (N_12329,N_11671,N_11952);
or U12330 (N_12330,N_11834,N_11926);
xnor U12331 (N_12331,N_11609,N_11757);
nor U12332 (N_12332,N_11750,N_11644);
xor U12333 (N_12333,N_11895,N_11997);
nor U12334 (N_12334,N_11603,N_11609);
xor U12335 (N_12335,N_11943,N_11875);
nand U12336 (N_12336,N_11901,N_11858);
and U12337 (N_12337,N_11831,N_11985);
nand U12338 (N_12338,N_11645,N_11729);
and U12339 (N_12339,N_11675,N_11891);
and U12340 (N_12340,N_11769,N_11782);
or U12341 (N_12341,N_11853,N_11613);
nand U12342 (N_12342,N_11980,N_11955);
and U12343 (N_12343,N_11734,N_11957);
and U12344 (N_12344,N_11820,N_11646);
and U12345 (N_12345,N_11860,N_11804);
nand U12346 (N_12346,N_11744,N_11640);
or U12347 (N_12347,N_11606,N_11649);
nor U12348 (N_12348,N_11655,N_11971);
xor U12349 (N_12349,N_11692,N_11955);
nand U12350 (N_12350,N_11611,N_11986);
nand U12351 (N_12351,N_11654,N_11683);
nand U12352 (N_12352,N_11600,N_11643);
nand U12353 (N_12353,N_11775,N_11980);
and U12354 (N_12354,N_11861,N_11970);
nand U12355 (N_12355,N_11893,N_11672);
and U12356 (N_12356,N_11911,N_11819);
nor U12357 (N_12357,N_11980,N_11774);
and U12358 (N_12358,N_11945,N_11630);
nand U12359 (N_12359,N_11997,N_11607);
and U12360 (N_12360,N_11970,N_11816);
nor U12361 (N_12361,N_11913,N_11935);
or U12362 (N_12362,N_11854,N_11921);
or U12363 (N_12363,N_11724,N_11991);
xnor U12364 (N_12364,N_11743,N_11934);
and U12365 (N_12365,N_11711,N_11962);
and U12366 (N_12366,N_11635,N_11701);
xor U12367 (N_12367,N_11889,N_11603);
xnor U12368 (N_12368,N_11958,N_11749);
or U12369 (N_12369,N_11898,N_11981);
nand U12370 (N_12370,N_11904,N_11628);
and U12371 (N_12371,N_11715,N_11631);
or U12372 (N_12372,N_11626,N_11685);
nand U12373 (N_12373,N_11983,N_11949);
nor U12374 (N_12374,N_11932,N_11907);
nand U12375 (N_12375,N_11760,N_11774);
or U12376 (N_12376,N_11705,N_11977);
nand U12377 (N_12377,N_11882,N_11870);
or U12378 (N_12378,N_11819,N_11766);
and U12379 (N_12379,N_11746,N_11919);
or U12380 (N_12380,N_11892,N_11859);
or U12381 (N_12381,N_11972,N_11644);
or U12382 (N_12382,N_11804,N_11972);
xnor U12383 (N_12383,N_11705,N_11962);
xnor U12384 (N_12384,N_11669,N_11731);
nor U12385 (N_12385,N_11835,N_11648);
nand U12386 (N_12386,N_11941,N_11747);
xor U12387 (N_12387,N_11745,N_11985);
nand U12388 (N_12388,N_11618,N_11842);
or U12389 (N_12389,N_11919,N_11938);
nand U12390 (N_12390,N_11912,N_11796);
xnor U12391 (N_12391,N_11605,N_11900);
and U12392 (N_12392,N_11752,N_11855);
or U12393 (N_12393,N_11803,N_11745);
and U12394 (N_12394,N_11711,N_11693);
nor U12395 (N_12395,N_11611,N_11758);
or U12396 (N_12396,N_11993,N_11774);
and U12397 (N_12397,N_11661,N_11602);
nand U12398 (N_12398,N_11938,N_11621);
or U12399 (N_12399,N_11745,N_11979);
and U12400 (N_12400,N_12096,N_12029);
and U12401 (N_12401,N_12392,N_12195);
nor U12402 (N_12402,N_12156,N_12199);
xnor U12403 (N_12403,N_12024,N_12163);
nor U12404 (N_12404,N_12296,N_12311);
nand U12405 (N_12405,N_12299,N_12042);
xnor U12406 (N_12406,N_12372,N_12216);
nand U12407 (N_12407,N_12355,N_12119);
nand U12408 (N_12408,N_12356,N_12287);
nor U12409 (N_12409,N_12185,N_12089);
or U12410 (N_12410,N_12290,N_12208);
xor U12411 (N_12411,N_12159,N_12212);
nor U12412 (N_12412,N_12055,N_12080);
nor U12413 (N_12413,N_12245,N_12386);
xor U12414 (N_12414,N_12368,N_12016);
or U12415 (N_12415,N_12142,N_12230);
nand U12416 (N_12416,N_12031,N_12121);
and U12417 (N_12417,N_12277,N_12380);
or U12418 (N_12418,N_12072,N_12394);
and U12419 (N_12419,N_12381,N_12207);
xor U12420 (N_12420,N_12047,N_12065);
nor U12421 (N_12421,N_12345,N_12048);
nor U12422 (N_12422,N_12340,N_12013);
and U12423 (N_12423,N_12050,N_12218);
nor U12424 (N_12424,N_12330,N_12169);
xor U12425 (N_12425,N_12187,N_12382);
xnor U12426 (N_12426,N_12081,N_12348);
nor U12427 (N_12427,N_12360,N_12113);
xnor U12428 (N_12428,N_12166,N_12133);
or U12429 (N_12429,N_12030,N_12231);
nand U12430 (N_12430,N_12160,N_12061);
nand U12431 (N_12431,N_12329,N_12312);
nor U12432 (N_12432,N_12366,N_12377);
and U12433 (N_12433,N_12399,N_12017);
xnor U12434 (N_12434,N_12197,N_12250);
nor U12435 (N_12435,N_12173,N_12075);
nand U12436 (N_12436,N_12052,N_12153);
or U12437 (N_12437,N_12229,N_12264);
or U12438 (N_12438,N_12064,N_12182);
and U12439 (N_12439,N_12371,N_12379);
nor U12440 (N_12440,N_12301,N_12375);
nand U12441 (N_12441,N_12053,N_12391);
nor U12442 (N_12442,N_12200,N_12083);
and U12443 (N_12443,N_12023,N_12003);
or U12444 (N_12444,N_12222,N_12140);
and U12445 (N_12445,N_12210,N_12268);
and U12446 (N_12446,N_12148,N_12398);
nand U12447 (N_12447,N_12190,N_12221);
xor U12448 (N_12448,N_12035,N_12079);
or U12449 (N_12449,N_12135,N_12337);
or U12450 (N_12450,N_12165,N_12309);
or U12451 (N_12451,N_12105,N_12331);
xnor U12452 (N_12452,N_12044,N_12223);
nand U12453 (N_12453,N_12178,N_12102);
or U12454 (N_12454,N_12319,N_12383);
or U12455 (N_12455,N_12149,N_12310);
and U12456 (N_12456,N_12009,N_12155);
nor U12457 (N_12457,N_12300,N_12070);
xnor U12458 (N_12458,N_12120,N_12193);
nor U12459 (N_12459,N_12302,N_12320);
nor U12460 (N_12460,N_12242,N_12104);
xnor U12461 (N_12461,N_12201,N_12339);
xnor U12462 (N_12462,N_12059,N_12248);
or U12463 (N_12463,N_12343,N_12184);
or U12464 (N_12464,N_12077,N_12293);
xor U12465 (N_12465,N_12259,N_12332);
xor U12466 (N_12466,N_12137,N_12114);
and U12467 (N_12467,N_12313,N_12060);
and U12468 (N_12468,N_12385,N_12316);
xnor U12469 (N_12469,N_12269,N_12097);
and U12470 (N_12470,N_12349,N_12361);
and U12471 (N_12471,N_12235,N_12007);
xnor U12472 (N_12472,N_12325,N_12327);
and U12473 (N_12473,N_12188,N_12006);
nor U12474 (N_12474,N_12227,N_12074);
or U12475 (N_12475,N_12134,N_12344);
nand U12476 (N_12476,N_12132,N_12046);
or U12477 (N_12477,N_12298,N_12295);
nand U12478 (N_12478,N_12318,N_12352);
and U12479 (N_12479,N_12037,N_12236);
or U12480 (N_12480,N_12151,N_12004);
or U12481 (N_12481,N_12014,N_12239);
nor U12482 (N_12482,N_12001,N_12334);
or U12483 (N_12483,N_12261,N_12171);
nand U12484 (N_12484,N_12333,N_12143);
nand U12485 (N_12485,N_12049,N_12198);
and U12486 (N_12486,N_12373,N_12152);
or U12487 (N_12487,N_12091,N_12365);
nor U12488 (N_12488,N_12186,N_12088);
nor U12489 (N_12489,N_12246,N_12018);
nand U12490 (N_12490,N_12280,N_12128);
nand U12491 (N_12491,N_12021,N_12043);
nand U12492 (N_12492,N_12226,N_12283);
or U12493 (N_12493,N_12191,N_12202);
xnor U12494 (N_12494,N_12034,N_12117);
nor U12495 (N_12495,N_12328,N_12095);
or U12496 (N_12496,N_12374,N_12336);
or U12497 (N_12497,N_12051,N_12346);
and U12498 (N_12498,N_12350,N_12291);
nand U12499 (N_12499,N_12256,N_12127);
and U12500 (N_12500,N_12292,N_12110);
nand U12501 (N_12501,N_12270,N_12157);
and U12502 (N_12502,N_12168,N_12285);
xnor U12503 (N_12503,N_12063,N_12158);
or U12504 (N_12504,N_12090,N_12251);
xnor U12505 (N_12505,N_12179,N_12122);
and U12506 (N_12506,N_12136,N_12062);
nor U12507 (N_12507,N_12196,N_12027);
and U12508 (N_12508,N_12303,N_12111);
nor U12509 (N_12509,N_12278,N_12359);
xor U12510 (N_12510,N_12369,N_12323);
nand U12511 (N_12511,N_12150,N_12289);
xor U12512 (N_12512,N_12262,N_12011);
nor U12513 (N_12513,N_12162,N_12306);
or U12514 (N_12514,N_12315,N_12396);
or U12515 (N_12515,N_12177,N_12321);
and U12516 (N_12516,N_12008,N_12108);
xnor U12517 (N_12517,N_12214,N_12260);
and U12518 (N_12518,N_12294,N_12267);
nor U12519 (N_12519,N_12025,N_12351);
nor U12520 (N_12520,N_12005,N_12286);
nand U12521 (N_12521,N_12341,N_12039);
or U12522 (N_12522,N_12206,N_12237);
nor U12523 (N_12523,N_12228,N_12305);
and U12524 (N_12524,N_12068,N_12271);
xnor U12525 (N_12525,N_12357,N_12161);
or U12526 (N_12526,N_12066,N_12106);
nand U12527 (N_12527,N_12279,N_12189);
or U12528 (N_12528,N_12205,N_12054);
nand U12529 (N_12529,N_12243,N_12308);
nor U12530 (N_12530,N_12093,N_12082);
xnor U12531 (N_12531,N_12026,N_12194);
and U12532 (N_12532,N_12376,N_12232);
nand U12533 (N_12533,N_12086,N_12087);
xnor U12534 (N_12534,N_12238,N_12304);
nor U12535 (N_12535,N_12322,N_12020);
nand U12536 (N_12536,N_12130,N_12022);
nor U12537 (N_12537,N_12118,N_12126);
and U12538 (N_12538,N_12183,N_12220);
or U12539 (N_12539,N_12019,N_12213);
xor U12540 (N_12540,N_12098,N_12273);
or U12541 (N_12541,N_12266,N_12378);
or U12542 (N_12542,N_12367,N_12254);
and U12543 (N_12543,N_12056,N_12028);
and U12544 (N_12544,N_12057,N_12099);
nor U12545 (N_12545,N_12282,N_12275);
nor U12546 (N_12546,N_12129,N_12107);
nor U12547 (N_12547,N_12180,N_12170);
and U12548 (N_12548,N_12146,N_12244);
nand U12549 (N_12549,N_12217,N_12347);
nand U12550 (N_12550,N_12253,N_12094);
or U12551 (N_12551,N_12116,N_12307);
nand U12552 (N_12552,N_12085,N_12125);
nor U12553 (N_12553,N_12233,N_12384);
nand U12554 (N_12554,N_12058,N_12138);
xor U12555 (N_12555,N_12224,N_12076);
and U12556 (N_12556,N_12203,N_12247);
xnor U12557 (N_12557,N_12390,N_12338);
and U12558 (N_12558,N_12240,N_12326);
nor U12559 (N_12559,N_12387,N_12252);
or U12560 (N_12560,N_12175,N_12219);
xnor U12561 (N_12561,N_12147,N_12272);
nand U12562 (N_12562,N_12032,N_12274);
nand U12563 (N_12563,N_12015,N_12265);
nand U12564 (N_12564,N_12036,N_12362);
xnor U12565 (N_12565,N_12174,N_12364);
nand U12566 (N_12566,N_12389,N_12172);
and U12567 (N_12567,N_12144,N_12314);
xor U12568 (N_12568,N_12281,N_12354);
xor U12569 (N_12569,N_12012,N_12234);
nand U12570 (N_12570,N_12215,N_12045);
nand U12571 (N_12571,N_12363,N_12033);
nor U12572 (N_12572,N_12154,N_12209);
xnor U12573 (N_12573,N_12257,N_12204);
and U12574 (N_12574,N_12258,N_12071);
xor U12575 (N_12575,N_12288,N_12353);
nor U12576 (N_12576,N_12040,N_12284);
and U12577 (N_12577,N_12176,N_12109);
and U12578 (N_12578,N_12112,N_12241);
and U12579 (N_12579,N_12010,N_12002);
and U12580 (N_12580,N_12000,N_12370);
xnor U12581 (N_12581,N_12092,N_12041);
and U12582 (N_12582,N_12255,N_12141);
nand U12583 (N_12583,N_12167,N_12324);
or U12584 (N_12584,N_12139,N_12103);
and U12585 (N_12585,N_12225,N_12073);
nor U12586 (N_12586,N_12395,N_12115);
and U12587 (N_12587,N_12100,N_12069);
nor U12588 (N_12588,N_12145,N_12342);
nor U12589 (N_12589,N_12276,N_12078);
nor U12590 (N_12590,N_12124,N_12263);
xor U12591 (N_12591,N_12131,N_12211);
xor U12592 (N_12592,N_12192,N_12335);
xor U12593 (N_12593,N_12123,N_12038);
xnor U12594 (N_12594,N_12317,N_12084);
or U12595 (N_12595,N_12393,N_12358);
or U12596 (N_12596,N_12249,N_12397);
nand U12597 (N_12597,N_12164,N_12388);
nand U12598 (N_12598,N_12067,N_12181);
or U12599 (N_12599,N_12297,N_12101);
nor U12600 (N_12600,N_12316,N_12366);
and U12601 (N_12601,N_12013,N_12273);
nor U12602 (N_12602,N_12391,N_12201);
or U12603 (N_12603,N_12247,N_12069);
or U12604 (N_12604,N_12213,N_12276);
nand U12605 (N_12605,N_12163,N_12138);
xor U12606 (N_12606,N_12148,N_12263);
or U12607 (N_12607,N_12113,N_12106);
nor U12608 (N_12608,N_12170,N_12119);
xor U12609 (N_12609,N_12038,N_12324);
or U12610 (N_12610,N_12211,N_12266);
or U12611 (N_12611,N_12149,N_12355);
xor U12612 (N_12612,N_12294,N_12158);
nand U12613 (N_12613,N_12315,N_12127);
nor U12614 (N_12614,N_12119,N_12389);
xor U12615 (N_12615,N_12104,N_12287);
and U12616 (N_12616,N_12355,N_12378);
or U12617 (N_12617,N_12107,N_12147);
or U12618 (N_12618,N_12022,N_12039);
or U12619 (N_12619,N_12106,N_12387);
and U12620 (N_12620,N_12030,N_12312);
nor U12621 (N_12621,N_12119,N_12130);
nand U12622 (N_12622,N_12333,N_12368);
and U12623 (N_12623,N_12286,N_12048);
xor U12624 (N_12624,N_12044,N_12249);
xnor U12625 (N_12625,N_12024,N_12170);
xor U12626 (N_12626,N_12148,N_12240);
nor U12627 (N_12627,N_12364,N_12021);
xnor U12628 (N_12628,N_12195,N_12296);
nand U12629 (N_12629,N_12217,N_12215);
or U12630 (N_12630,N_12346,N_12159);
nor U12631 (N_12631,N_12167,N_12329);
or U12632 (N_12632,N_12017,N_12389);
nand U12633 (N_12633,N_12026,N_12035);
and U12634 (N_12634,N_12370,N_12238);
or U12635 (N_12635,N_12238,N_12369);
and U12636 (N_12636,N_12171,N_12276);
and U12637 (N_12637,N_12184,N_12242);
and U12638 (N_12638,N_12223,N_12201);
and U12639 (N_12639,N_12208,N_12120);
nand U12640 (N_12640,N_12175,N_12253);
nand U12641 (N_12641,N_12150,N_12042);
xnor U12642 (N_12642,N_12260,N_12251);
or U12643 (N_12643,N_12075,N_12389);
nand U12644 (N_12644,N_12040,N_12004);
nor U12645 (N_12645,N_12364,N_12212);
or U12646 (N_12646,N_12168,N_12275);
and U12647 (N_12647,N_12013,N_12139);
and U12648 (N_12648,N_12064,N_12005);
nand U12649 (N_12649,N_12257,N_12136);
or U12650 (N_12650,N_12335,N_12170);
or U12651 (N_12651,N_12299,N_12072);
xnor U12652 (N_12652,N_12322,N_12329);
nand U12653 (N_12653,N_12271,N_12150);
xor U12654 (N_12654,N_12333,N_12209);
or U12655 (N_12655,N_12239,N_12055);
and U12656 (N_12656,N_12315,N_12250);
nand U12657 (N_12657,N_12125,N_12213);
xnor U12658 (N_12658,N_12034,N_12241);
xor U12659 (N_12659,N_12087,N_12174);
or U12660 (N_12660,N_12177,N_12217);
nor U12661 (N_12661,N_12319,N_12314);
xnor U12662 (N_12662,N_12005,N_12172);
nand U12663 (N_12663,N_12393,N_12382);
nand U12664 (N_12664,N_12206,N_12374);
nand U12665 (N_12665,N_12362,N_12380);
or U12666 (N_12666,N_12188,N_12082);
and U12667 (N_12667,N_12260,N_12381);
nand U12668 (N_12668,N_12173,N_12175);
nand U12669 (N_12669,N_12101,N_12202);
or U12670 (N_12670,N_12266,N_12385);
nand U12671 (N_12671,N_12017,N_12286);
nor U12672 (N_12672,N_12014,N_12104);
nand U12673 (N_12673,N_12238,N_12146);
or U12674 (N_12674,N_12350,N_12027);
nor U12675 (N_12675,N_12001,N_12122);
and U12676 (N_12676,N_12209,N_12114);
and U12677 (N_12677,N_12322,N_12369);
nand U12678 (N_12678,N_12127,N_12034);
nand U12679 (N_12679,N_12117,N_12247);
nand U12680 (N_12680,N_12229,N_12142);
nor U12681 (N_12681,N_12276,N_12227);
nor U12682 (N_12682,N_12041,N_12222);
nand U12683 (N_12683,N_12191,N_12068);
nor U12684 (N_12684,N_12112,N_12238);
and U12685 (N_12685,N_12286,N_12318);
and U12686 (N_12686,N_12365,N_12264);
nand U12687 (N_12687,N_12392,N_12102);
xor U12688 (N_12688,N_12173,N_12162);
nor U12689 (N_12689,N_12321,N_12037);
xnor U12690 (N_12690,N_12204,N_12102);
nand U12691 (N_12691,N_12345,N_12302);
and U12692 (N_12692,N_12201,N_12110);
or U12693 (N_12693,N_12096,N_12109);
nand U12694 (N_12694,N_12058,N_12381);
xor U12695 (N_12695,N_12208,N_12279);
or U12696 (N_12696,N_12112,N_12374);
xor U12697 (N_12697,N_12117,N_12006);
nor U12698 (N_12698,N_12161,N_12321);
xor U12699 (N_12699,N_12163,N_12144);
nand U12700 (N_12700,N_12146,N_12276);
and U12701 (N_12701,N_12224,N_12327);
nor U12702 (N_12702,N_12146,N_12174);
nor U12703 (N_12703,N_12227,N_12041);
nand U12704 (N_12704,N_12191,N_12016);
nor U12705 (N_12705,N_12043,N_12266);
nor U12706 (N_12706,N_12097,N_12256);
or U12707 (N_12707,N_12349,N_12351);
nand U12708 (N_12708,N_12180,N_12227);
and U12709 (N_12709,N_12148,N_12282);
and U12710 (N_12710,N_12346,N_12178);
or U12711 (N_12711,N_12369,N_12331);
or U12712 (N_12712,N_12134,N_12175);
and U12713 (N_12713,N_12026,N_12109);
or U12714 (N_12714,N_12220,N_12246);
or U12715 (N_12715,N_12387,N_12386);
or U12716 (N_12716,N_12325,N_12356);
and U12717 (N_12717,N_12224,N_12259);
and U12718 (N_12718,N_12018,N_12387);
nand U12719 (N_12719,N_12288,N_12043);
nor U12720 (N_12720,N_12037,N_12012);
and U12721 (N_12721,N_12177,N_12073);
nor U12722 (N_12722,N_12330,N_12306);
nand U12723 (N_12723,N_12247,N_12202);
xor U12724 (N_12724,N_12214,N_12074);
nand U12725 (N_12725,N_12209,N_12198);
or U12726 (N_12726,N_12157,N_12234);
nor U12727 (N_12727,N_12350,N_12352);
nor U12728 (N_12728,N_12185,N_12260);
nand U12729 (N_12729,N_12108,N_12062);
or U12730 (N_12730,N_12294,N_12313);
and U12731 (N_12731,N_12241,N_12396);
and U12732 (N_12732,N_12123,N_12242);
nand U12733 (N_12733,N_12314,N_12218);
or U12734 (N_12734,N_12170,N_12138);
nor U12735 (N_12735,N_12119,N_12016);
and U12736 (N_12736,N_12124,N_12194);
nor U12737 (N_12737,N_12070,N_12071);
nor U12738 (N_12738,N_12050,N_12353);
xnor U12739 (N_12739,N_12305,N_12158);
nand U12740 (N_12740,N_12340,N_12115);
xnor U12741 (N_12741,N_12272,N_12105);
and U12742 (N_12742,N_12146,N_12162);
xor U12743 (N_12743,N_12056,N_12063);
or U12744 (N_12744,N_12104,N_12093);
and U12745 (N_12745,N_12399,N_12287);
and U12746 (N_12746,N_12189,N_12327);
nand U12747 (N_12747,N_12111,N_12215);
and U12748 (N_12748,N_12325,N_12182);
and U12749 (N_12749,N_12032,N_12118);
nor U12750 (N_12750,N_12363,N_12128);
nor U12751 (N_12751,N_12060,N_12016);
and U12752 (N_12752,N_12198,N_12073);
xnor U12753 (N_12753,N_12395,N_12373);
and U12754 (N_12754,N_12399,N_12098);
nand U12755 (N_12755,N_12224,N_12101);
xor U12756 (N_12756,N_12288,N_12100);
nand U12757 (N_12757,N_12318,N_12285);
or U12758 (N_12758,N_12235,N_12239);
nand U12759 (N_12759,N_12220,N_12088);
xnor U12760 (N_12760,N_12060,N_12339);
and U12761 (N_12761,N_12218,N_12259);
and U12762 (N_12762,N_12266,N_12391);
or U12763 (N_12763,N_12226,N_12299);
or U12764 (N_12764,N_12306,N_12049);
nor U12765 (N_12765,N_12307,N_12301);
xnor U12766 (N_12766,N_12245,N_12184);
xor U12767 (N_12767,N_12202,N_12089);
nand U12768 (N_12768,N_12213,N_12249);
or U12769 (N_12769,N_12096,N_12161);
nand U12770 (N_12770,N_12046,N_12202);
nand U12771 (N_12771,N_12094,N_12157);
nand U12772 (N_12772,N_12380,N_12325);
nand U12773 (N_12773,N_12177,N_12294);
and U12774 (N_12774,N_12068,N_12177);
and U12775 (N_12775,N_12182,N_12021);
xnor U12776 (N_12776,N_12384,N_12019);
or U12777 (N_12777,N_12311,N_12114);
and U12778 (N_12778,N_12170,N_12347);
nand U12779 (N_12779,N_12294,N_12076);
or U12780 (N_12780,N_12287,N_12142);
nor U12781 (N_12781,N_12173,N_12119);
xor U12782 (N_12782,N_12243,N_12269);
or U12783 (N_12783,N_12387,N_12308);
nor U12784 (N_12784,N_12088,N_12201);
xnor U12785 (N_12785,N_12149,N_12030);
nand U12786 (N_12786,N_12113,N_12005);
nor U12787 (N_12787,N_12219,N_12028);
xnor U12788 (N_12788,N_12174,N_12093);
nor U12789 (N_12789,N_12007,N_12045);
and U12790 (N_12790,N_12035,N_12370);
nor U12791 (N_12791,N_12246,N_12024);
and U12792 (N_12792,N_12246,N_12268);
nand U12793 (N_12793,N_12253,N_12364);
and U12794 (N_12794,N_12149,N_12083);
nor U12795 (N_12795,N_12327,N_12374);
and U12796 (N_12796,N_12000,N_12228);
or U12797 (N_12797,N_12231,N_12162);
nand U12798 (N_12798,N_12329,N_12382);
and U12799 (N_12799,N_12180,N_12109);
nand U12800 (N_12800,N_12672,N_12670);
and U12801 (N_12801,N_12702,N_12738);
and U12802 (N_12802,N_12606,N_12709);
and U12803 (N_12803,N_12425,N_12525);
nand U12804 (N_12804,N_12778,N_12576);
xnor U12805 (N_12805,N_12611,N_12724);
xor U12806 (N_12806,N_12439,N_12695);
xor U12807 (N_12807,N_12733,N_12698);
or U12808 (N_12808,N_12661,N_12686);
or U12809 (N_12809,N_12510,N_12448);
nand U12810 (N_12810,N_12496,N_12572);
nand U12811 (N_12811,N_12538,N_12453);
and U12812 (N_12812,N_12789,N_12684);
xor U12813 (N_12813,N_12430,N_12776);
xor U12814 (N_12814,N_12527,N_12402);
and U12815 (N_12815,N_12557,N_12751);
nor U12816 (N_12816,N_12436,N_12750);
or U12817 (N_12817,N_12705,N_12495);
nor U12818 (N_12818,N_12762,N_12506);
xnor U12819 (N_12819,N_12437,N_12563);
and U12820 (N_12820,N_12679,N_12416);
or U12821 (N_12821,N_12536,N_12788);
nand U12822 (N_12822,N_12450,N_12467);
or U12823 (N_12823,N_12619,N_12405);
xnor U12824 (N_12824,N_12745,N_12499);
and U12825 (N_12825,N_12498,N_12432);
or U12826 (N_12826,N_12710,N_12683);
nor U12827 (N_12827,N_12719,N_12647);
nor U12828 (N_12828,N_12784,N_12526);
and U12829 (N_12829,N_12799,N_12642);
and U12830 (N_12830,N_12452,N_12478);
xor U12831 (N_12831,N_12463,N_12699);
xor U12832 (N_12832,N_12424,N_12616);
xnor U12833 (N_12833,N_12585,N_12404);
or U12834 (N_12834,N_12484,N_12598);
nand U12835 (N_12835,N_12435,N_12791);
nor U12836 (N_12836,N_12515,N_12420);
nor U12837 (N_12837,N_12639,N_12769);
nor U12838 (N_12838,N_12730,N_12549);
xnor U12839 (N_12839,N_12472,N_12663);
and U12840 (N_12840,N_12595,N_12792);
or U12841 (N_12841,N_12537,N_12741);
nand U12842 (N_12842,N_12466,N_12521);
and U12843 (N_12843,N_12516,N_12423);
or U12844 (N_12844,N_12440,N_12454);
and U12845 (N_12845,N_12600,N_12480);
and U12846 (N_12846,N_12421,N_12594);
nand U12847 (N_12847,N_12651,N_12685);
nand U12848 (N_12848,N_12773,N_12471);
nor U12849 (N_12849,N_12566,N_12654);
nor U12850 (N_12850,N_12414,N_12535);
and U12851 (N_12851,N_12697,N_12485);
nor U12852 (N_12852,N_12748,N_12599);
xnor U12853 (N_12853,N_12627,N_12446);
and U12854 (N_12854,N_12785,N_12715);
and U12855 (N_12855,N_12579,N_12665);
and U12856 (N_12856,N_12490,N_12575);
nand U12857 (N_12857,N_12509,N_12468);
and U12858 (N_12858,N_12633,N_12637);
xor U12859 (N_12859,N_12507,N_12584);
or U12860 (N_12860,N_12671,N_12641);
and U12861 (N_12861,N_12754,N_12489);
nor U12862 (N_12862,N_12529,N_12434);
or U12863 (N_12863,N_12593,N_12493);
and U12864 (N_12864,N_12483,N_12708);
nor U12865 (N_12865,N_12532,N_12588);
xor U12866 (N_12866,N_12429,N_12644);
and U12867 (N_12867,N_12765,N_12638);
and U12868 (N_12868,N_12486,N_12624);
xor U12869 (N_12869,N_12722,N_12597);
and U12870 (N_12870,N_12688,N_12592);
or U12871 (N_12871,N_12550,N_12634);
or U12872 (N_12872,N_12564,N_12504);
or U12873 (N_12873,N_12796,N_12479);
or U12874 (N_12874,N_12407,N_12548);
or U12875 (N_12875,N_12497,N_12590);
nor U12876 (N_12876,N_12691,N_12706);
nand U12877 (N_12877,N_12739,N_12519);
nor U12878 (N_12878,N_12607,N_12441);
and U12879 (N_12879,N_12783,N_12712);
nand U12880 (N_12880,N_12674,N_12682);
nor U12881 (N_12881,N_12613,N_12426);
or U12882 (N_12882,N_12676,N_12621);
nand U12883 (N_12883,N_12793,N_12689);
or U12884 (N_12884,N_12657,N_12492);
xor U12885 (N_12885,N_12401,N_12523);
nand U12886 (N_12886,N_12469,N_12562);
or U12887 (N_12887,N_12589,N_12675);
nor U12888 (N_12888,N_12797,N_12617);
and U12889 (N_12889,N_12474,N_12544);
or U12890 (N_12890,N_12727,N_12666);
or U12891 (N_12891,N_12707,N_12481);
nand U12892 (N_12892,N_12455,N_12664);
nand U12893 (N_12893,N_12615,N_12582);
nor U12894 (N_12894,N_12512,N_12626);
nor U12895 (N_12895,N_12655,N_12763);
and U12896 (N_12896,N_12703,N_12458);
or U12897 (N_12897,N_12660,N_12410);
and U12898 (N_12898,N_12648,N_12723);
and U12899 (N_12899,N_12746,N_12462);
or U12900 (N_12900,N_12524,N_12400);
and U12901 (N_12901,N_12444,N_12629);
or U12902 (N_12902,N_12780,N_12500);
xor U12903 (N_12903,N_12596,N_12716);
nor U12904 (N_12904,N_12680,N_12728);
and U12905 (N_12905,N_12650,N_12687);
nand U12906 (N_12906,N_12749,N_12764);
and U12907 (N_12907,N_12692,N_12412);
and U12908 (N_12908,N_12678,N_12605);
or U12909 (N_12909,N_12554,N_12438);
and U12910 (N_12910,N_12726,N_12433);
or U12911 (N_12911,N_12658,N_12758);
nor U12912 (N_12912,N_12417,N_12587);
or U12913 (N_12913,N_12561,N_12571);
nor U12914 (N_12914,N_12476,N_12568);
xor U12915 (N_12915,N_12591,N_12623);
nor U12916 (N_12916,N_12503,N_12413);
nor U12917 (N_12917,N_12445,N_12461);
and U12918 (N_12918,N_12668,N_12431);
nand U12919 (N_12919,N_12403,N_12772);
or U12920 (N_12920,N_12681,N_12477);
and U12921 (N_12921,N_12517,N_12761);
nor U12922 (N_12922,N_12694,N_12505);
or U12923 (N_12923,N_12736,N_12570);
or U12924 (N_12924,N_12636,N_12534);
and U12925 (N_12925,N_12714,N_12742);
and U12926 (N_12926,N_12408,N_12482);
nand U12927 (N_12927,N_12622,N_12475);
nor U12928 (N_12928,N_12552,N_12625);
xor U12929 (N_12929,N_12720,N_12774);
or U12930 (N_12930,N_12460,N_12643);
nand U12931 (N_12931,N_12555,N_12604);
nor U12932 (N_12932,N_12649,N_12620);
nor U12933 (N_12933,N_12646,N_12528);
nor U12934 (N_12934,N_12752,N_12545);
xor U12935 (N_12935,N_12508,N_12721);
and U12936 (N_12936,N_12560,N_12565);
xor U12937 (N_12937,N_12464,N_12608);
or U12938 (N_12938,N_12418,N_12669);
nor U12939 (N_12939,N_12744,N_12511);
or U12940 (N_12940,N_12795,N_12574);
nand U12941 (N_12941,N_12770,N_12662);
nor U12942 (N_12942,N_12737,N_12541);
and U12943 (N_12943,N_12547,N_12558);
nand U12944 (N_12944,N_12743,N_12757);
and U12945 (N_12945,N_12533,N_12735);
and U12946 (N_12946,N_12630,N_12777);
xnor U12947 (N_12947,N_12488,N_12411);
nor U12948 (N_12948,N_12614,N_12790);
or U12949 (N_12949,N_12696,N_12610);
or U12950 (N_12950,N_12732,N_12518);
or U12951 (N_12951,N_12768,N_12456);
xnor U12952 (N_12952,N_12766,N_12711);
xor U12953 (N_12953,N_12580,N_12406);
and U12954 (N_12954,N_12618,N_12451);
or U12955 (N_12955,N_12567,N_12546);
xor U12956 (N_12956,N_12577,N_12559);
nand U12957 (N_12957,N_12513,N_12573);
nand U12958 (N_12958,N_12794,N_12428);
nor U12959 (N_12959,N_12427,N_12640);
or U12960 (N_12960,N_12470,N_12656);
xor U12961 (N_12961,N_12586,N_12457);
or U12962 (N_12962,N_12449,N_12731);
and U12963 (N_12963,N_12540,N_12539);
nand U12964 (N_12964,N_12601,N_12422);
nor U12965 (N_12965,N_12781,N_12583);
and U12966 (N_12966,N_12522,N_12747);
or U12967 (N_12967,N_12659,N_12775);
xnor U12968 (N_12968,N_12415,N_12631);
nor U12969 (N_12969,N_12556,N_12713);
xor U12970 (N_12970,N_12612,N_12779);
xor U12971 (N_12971,N_12494,N_12419);
nand U12972 (N_12972,N_12442,N_12628);
nor U12973 (N_12973,N_12645,N_12798);
xnor U12974 (N_12974,N_12531,N_12514);
nand U12975 (N_12975,N_12447,N_12690);
and U12976 (N_12976,N_12473,N_12786);
and U12977 (N_12977,N_12725,N_12653);
or U12978 (N_12978,N_12782,N_12581);
nor U12979 (N_12979,N_12491,N_12465);
and U12980 (N_12980,N_12704,N_12569);
and U12981 (N_12981,N_12502,N_12767);
nor U12982 (N_12982,N_12701,N_12771);
and U12983 (N_12983,N_12755,N_12520);
xor U12984 (N_12984,N_12667,N_12693);
or U12985 (N_12985,N_12635,N_12718);
nor U12986 (N_12986,N_12787,N_12543);
nand U12987 (N_12987,N_12530,N_12443);
xor U12988 (N_12988,N_12578,N_12632);
nand U12989 (N_12989,N_12459,N_12753);
or U12990 (N_12990,N_12717,N_12609);
nor U12991 (N_12991,N_12603,N_12551);
xor U12992 (N_12992,N_12700,N_12729);
or U12993 (N_12993,N_12602,N_12734);
nor U12994 (N_12994,N_12487,N_12760);
nor U12995 (N_12995,N_12501,N_12677);
and U12996 (N_12996,N_12756,N_12652);
nand U12997 (N_12997,N_12759,N_12673);
or U12998 (N_12998,N_12553,N_12409);
and U12999 (N_12999,N_12740,N_12542);
nor U13000 (N_13000,N_12668,N_12649);
or U13001 (N_13001,N_12683,N_12640);
or U13002 (N_13002,N_12649,N_12408);
and U13003 (N_13003,N_12497,N_12409);
or U13004 (N_13004,N_12663,N_12485);
xnor U13005 (N_13005,N_12736,N_12716);
and U13006 (N_13006,N_12454,N_12678);
xor U13007 (N_13007,N_12620,N_12625);
and U13008 (N_13008,N_12712,N_12694);
and U13009 (N_13009,N_12565,N_12541);
nand U13010 (N_13010,N_12680,N_12797);
or U13011 (N_13011,N_12529,N_12584);
xor U13012 (N_13012,N_12657,N_12497);
nand U13013 (N_13013,N_12783,N_12736);
nand U13014 (N_13014,N_12744,N_12493);
nor U13015 (N_13015,N_12420,N_12444);
nor U13016 (N_13016,N_12749,N_12677);
xor U13017 (N_13017,N_12644,N_12560);
nor U13018 (N_13018,N_12589,N_12625);
nor U13019 (N_13019,N_12614,N_12725);
and U13020 (N_13020,N_12435,N_12585);
nor U13021 (N_13021,N_12769,N_12576);
xnor U13022 (N_13022,N_12476,N_12644);
nand U13023 (N_13023,N_12453,N_12778);
or U13024 (N_13024,N_12564,N_12559);
xor U13025 (N_13025,N_12755,N_12596);
nand U13026 (N_13026,N_12678,N_12739);
nand U13027 (N_13027,N_12544,N_12457);
nand U13028 (N_13028,N_12488,N_12537);
and U13029 (N_13029,N_12794,N_12412);
nor U13030 (N_13030,N_12719,N_12624);
or U13031 (N_13031,N_12754,N_12446);
xor U13032 (N_13032,N_12533,N_12630);
xor U13033 (N_13033,N_12690,N_12600);
and U13034 (N_13034,N_12771,N_12447);
or U13035 (N_13035,N_12400,N_12495);
and U13036 (N_13036,N_12688,N_12537);
nand U13037 (N_13037,N_12524,N_12765);
or U13038 (N_13038,N_12518,N_12719);
nand U13039 (N_13039,N_12531,N_12724);
or U13040 (N_13040,N_12665,N_12499);
xnor U13041 (N_13041,N_12561,N_12430);
nor U13042 (N_13042,N_12545,N_12706);
xor U13043 (N_13043,N_12534,N_12467);
or U13044 (N_13044,N_12760,N_12567);
xnor U13045 (N_13045,N_12708,N_12401);
nor U13046 (N_13046,N_12485,N_12514);
xnor U13047 (N_13047,N_12688,N_12671);
and U13048 (N_13048,N_12627,N_12517);
and U13049 (N_13049,N_12542,N_12787);
or U13050 (N_13050,N_12492,N_12464);
and U13051 (N_13051,N_12683,N_12734);
or U13052 (N_13052,N_12777,N_12591);
nand U13053 (N_13053,N_12783,N_12606);
nor U13054 (N_13054,N_12503,N_12614);
nor U13055 (N_13055,N_12656,N_12492);
nand U13056 (N_13056,N_12742,N_12786);
nand U13057 (N_13057,N_12719,N_12691);
or U13058 (N_13058,N_12539,N_12498);
nand U13059 (N_13059,N_12510,N_12787);
xor U13060 (N_13060,N_12537,N_12565);
and U13061 (N_13061,N_12516,N_12474);
nand U13062 (N_13062,N_12406,N_12683);
and U13063 (N_13063,N_12596,N_12477);
nor U13064 (N_13064,N_12728,N_12552);
nand U13065 (N_13065,N_12587,N_12734);
nand U13066 (N_13066,N_12559,N_12703);
or U13067 (N_13067,N_12682,N_12418);
and U13068 (N_13068,N_12428,N_12470);
and U13069 (N_13069,N_12460,N_12697);
nor U13070 (N_13070,N_12402,N_12572);
nor U13071 (N_13071,N_12722,N_12609);
xnor U13072 (N_13072,N_12734,N_12637);
nand U13073 (N_13073,N_12442,N_12684);
and U13074 (N_13074,N_12680,N_12574);
or U13075 (N_13075,N_12651,N_12701);
or U13076 (N_13076,N_12402,N_12646);
and U13077 (N_13077,N_12516,N_12453);
nor U13078 (N_13078,N_12445,N_12528);
or U13079 (N_13079,N_12595,N_12515);
nor U13080 (N_13080,N_12488,N_12640);
and U13081 (N_13081,N_12402,N_12756);
and U13082 (N_13082,N_12615,N_12767);
or U13083 (N_13083,N_12414,N_12558);
nand U13084 (N_13084,N_12679,N_12561);
xnor U13085 (N_13085,N_12450,N_12669);
and U13086 (N_13086,N_12650,N_12786);
and U13087 (N_13087,N_12463,N_12691);
nand U13088 (N_13088,N_12783,N_12571);
nor U13089 (N_13089,N_12701,N_12615);
and U13090 (N_13090,N_12635,N_12497);
nand U13091 (N_13091,N_12635,N_12751);
xor U13092 (N_13092,N_12543,N_12771);
nor U13093 (N_13093,N_12644,N_12716);
and U13094 (N_13094,N_12731,N_12594);
xor U13095 (N_13095,N_12513,N_12470);
nand U13096 (N_13096,N_12657,N_12697);
and U13097 (N_13097,N_12633,N_12427);
nor U13098 (N_13098,N_12675,N_12799);
nor U13099 (N_13099,N_12608,N_12442);
and U13100 (N_13100,N_12432,N_12536);
nand U13101 (N_13101,N_12542,N_12454);
xor U13102 (N_13102,N_12569,N_12630);
and U13103 (N_13103,N_12681,N_12434);
nor U13104 (N_13104,N_12574,N_12457);
and U13105 (N_13105,N_12683,N_12634);
or U13106 (N_13106,N_12796,N_12501);
or U13107 (N_13107,N_12754,N_12554);
nand U13108 (N_13108,N_12672,N_12454);
and U13109 (N_13109,N_12682,N_12410);
xnor U13110 (N_13110,N_12716,N_12631);
nand U13111 (N_13111,N_12455,N_12554);
and U13112 (N_13112,N_12621,N_12582);
nand U13113 (N_13113,N_12659,N_12494);
or U13114 (N_13114,N_12772,N_12794);
nor U13115 (N_13115,N_12667,N_12735);
xor U13116 (N_13116,N_12524,N_12671);
and U13117 (N_13117,N_12520,N_12794);
xor U13118 (N_13118,N_12599,N_12485);
xor U13119 (N_13119,N_12707,N_12464);
and U13120 (N_13120,N_12696,N_12612);
or U13121 (N_13121,N_12785,N_12480);
nor U13122 (N_13122,N_12475,N_12451);
and U13123 (N_13123,N_12683,N_12779);
xor U13124 (N_13124,N_12542,N_12690);
and U13125 (N_13125,N_12683,N_12530);
or U13126 (N_13126,N_12620,N_12527);
or U13127 (N_13127,N_12513,N_12499);
xnor U13128 (N_13128,N_12549,N_12496);
and U13129 (N_13129,N_12595,N_12423);
nand U13130 (N_13130,N_12521,N_12453);
nand U13131 (N_13131,N_12517,N_12767);
or U13132 (N_13132,N_12470,N_12441);
nor U13133 (N_13133,N_12755,N_12705);
or U13134 (N_13134,N_12537,N_12736);
nor U13135 (N_13135,N_12474,N_12412);
nand U13136 (N_13136,N_12709,N_12470);
xor U13137 (N_13137,N_12482,N_12775);
nand U13138 (N_13138,N_12433,N_12520);
nor U13139 (N_13139,N_12658,N_12499);
nor U13140 (N_13140,N_12731,N_12418);
nor U13141 (N_13141,N_12686,N_12755);
xor U13142 (N_13142,N_12414,N_12676);
or U13143 (N_13143,N_12794,N_12789);
nand U13144 (N_13144,N_12637,N_12481);
nor U13145 (N_13145,N_12624,N_12691);
xor U13146 (N_13146,N_12439,N_12502);
nand U13147 (N_13147,N_12460,N_12549);
and U13148 (N_13148,N_12491,N_12785);
and U13149 (N_13149,N_12467,N_12638);
xor U13150 (N_13150,N_12562,N_12483);
or U13151 (N_13151,N_12719,N_12726);
xnor U13152 (N_13152,N_12537,N_12585);
nand U13153 (N_13153,N_12552,N_12646);
nor U13154 (N_13154,N_12551,N_12774);
xor U13155 (N_13155,N_12737,N_12501);
and U13156 (N_13156,N_12485,N_12641);
or U13157 (N_13157,N_12714,N_12419);
or U13158 (N_13158,N_12511,N_12690);
and U13159 (N_13159,N_12794,N_12444);
xnor U13160 (N_13160,N_12528,N_12641);
nor U13161 (N_13161,N_12638,N_12687);
xnor U13162 (N_13162,N_12506,N_12572);
nor U13163 (N_13163,N_12637,N_12706);
nor U13164 (N_13164,N_12617,N_12656);
and U13165 (N_13165,N_12569,N_12696);
xor U13166 (N_13166,N_12684,N_12522);
nor U13167 (N_13167,N_12432,N_12439);
and U13168 (N_13168,N_12425,N_12604);
nand U13169 (N_13169,N_12460,N_12545);
nor U13170 (N_13170,N_12687,N_12441);
and U13171 (N_13171,N_12428,N_12721);
and U13172 (N_13172,N_12698,N_12447);
and U13173 (N_13173,N_12492,N_12403);
xnor U13174 (N_13174,N_12546,N_12441);
or U13175 (N_13175,N_12637,N_12492);
and U13176 (N_13176,N_12764,N_12758);
or U13177 (N_13177,N_12671,N_12775);
xor U13178 (N_13178,N_12522,N_12543);
or U13179 (N_13179,N_12558,N_12798);
and U13180 (N_13180,N_12482,N_12656);
xnor U13181 (N_13181,N_12565,N_12650);
xnor U13182 (N_13182,N_12405,N_12437);
or U13183 (N_13183,N_12484,N_12732);
nand U13184 (N_13184,N_12639,N_12487);
or U13185 (N_13185,N_12752,N_12617);
xnor U13186 (N_13186,N_12787,N_12412);
nor U13187 (N_13187,N_12427,N_12441);
nor U13188 (N_13188,N_12755,N_12536);
xnor U13189 (N_13189,N_12531,N_12445);
nor U13190 (N_13190,N_12746,N_12711);
nand U13191 (N_13191,N_12758,N_12645);
nor U13192 (N_13192,N_12575,N_12677);
nand U13193 (N_13193,N_12679,N_12756);
and U13194 (N_13194,N_12523,N_12694);
nand U13195 (N_13195,N_12455,N_12563);
xor U13196 (N_13196,N_12684,N_12599);
nand U13197 (N_13197,N_12408,N_12647);
xor U13198 (N_13198,N_12684,N_12729);
nand U13199 (N_13199,N_12540,N_12754);
and U13200 (N_13200,N_12966,N_13028);
nor U13201 (N_13201,N_13088,N_12981);
nor U13202 (N_13202,N_12957,N_13037);
and U13203 (N_13203,N_13084,N_12924);
xor U13204 (N_13204,N_13188,N_13151);
or U13205 (N_13205,N_12994,N_12881);
xnor U13206 (N_13206,N_13081,N_12896);
nor U13207 (N_13207,N_13092,N_12891);
or U13208 (N_13208,N_13123,N_13101);
nor U13209 (N_13209,N_13046,N_13180);
and U13210 (N_13210,N_13022,N_13069);
nand U13211 (N_13211,N_12855,N_12802);
nand U13212 (N_13212,N_12932,N_12805);
nor U13213 (N_13213,N_13042,N_12913);
or U13214 (N_13214,N_13119,N_13172);
nor U13215 (N_13215,N_12955,N_12937);
or U13216 (N_13216,N_12817,N_12916);
and U13217 (N_13217,N_12845,N_13168);
or U13218 (N_13218,N_12972,N_12959);
nand U13219 (N_13219,N_12840,N_13135);
xnor U13220 (N_13220,N_12970,N_12879);
xor U13221 (N_13221,N_12919,N_12854);
and U13222 (N_13222,N_13139,N_13107);
nand U13223 (N_13223,N_12998,N_13045);
xnor U13224 (N_13224,N_13128,N_12943);
nand U13225 (N_13225,N_13083,N_12939);
xnor U13226 (N_13226,N_12894,N_13087);
and U13227 (N_13227,N_13072,N_13029);
or U13228 (N_13228,N_13016,N_13142);
nand U13229 (N_13229,N_13183,N_13075);
nand U13230 (N_13230,N_13059,N_13194);
and U13231 (N_13231,N_13167,N_12814);
nor U13232 (N_13232,N_13019,N_12931);
or U13233 (N_13233,N_12909,N_13140);
xor U13234 (N_13234,N_12857,N_13147);
nor U13235 (N_13235,N_13157,N_13031);
xor U13236 (N_13236,N_12942,N_13171);
nor U13237 (N_13237,N_12829,N_13114);
or U13238 (N_13238,N_12818,N_12899);
xnor U13239 (N_13239,N_12827,N_12807);
and U13240 (N_13240,N_12884,N_13111);
or U13241 (N_13241,N_12984,N_12882);
nand U13242 (N_13242,N_12858,N_12834);
nand U13243 (N_13243,N_12934,N_12800);
nand U13244 (N_13244,N_13163,N_12833);
and U13245 (N_13245,N_12904,N_13179);
xnor U13246 (N_13246,N_13047,N_12999);
nand U13247 (N_13247,N_12963,N_13152);
and U13248 (N_13248,N_12869,N_13025);
nand U13249 (N_13249,N_13121,N_13093);
and U13250 (N_13250,N_13080,N_12867);
nand U13251 (N_13251,N_12940,N_13078);
or U13252 (N_13252,N_13010,N_13043);
or U13253 (N_13253,N_13155,N_13000);
nor U13254 (N_13254,N_12996,N_12828);
xnor U13255 (N_13255,N_12961,N_13017);
and U13256 (N_13256,N_12809,N_13091);
and U13257 (N_13257,N_13174,N_13074);
or U13258 (N_13258,N_12822,N_12841);
nand U13259 (N_13259,N_13001,N_12908);
xor U13260 (N_13260,N_12836,N_12976);
and U13261 (N_13261,N_13076,N_12893);
nand U13262 (N_13262,N_13054,N_12941);
and U13263 (N_13263,N_13090,N_13098);
and U13264 (N_13264,N_12997,N_13041);
nor U13265 (N_13265,N_12946,N_12975);
or U13266 (N_13266,N_13064,N_12803);
xor U13267 (N_13267,N_12923,N_12987);
xnor U13268 (N_13268,N_13071,N_13068);
xnor U13269 (N_13269,N_13131,N_13053);
xor U13270 (N_13270,N_13013,N_12907);
or U13271 (N_13271,N_12830,N_13035);
and U13272 (N_13272,N_12826,N_12985);
or U13273 (N_13273,N_12849,N_13165);
nor U13274 (N_13274,N_12848,N_13170);
and U13275 (N_13275,N_13120,N_12842);
and U13276 (N_13276,N_13136,N_12921);
or U13277 (N_13277,N_12812,N_13097);
nor U13278 (N_13278,N_13115,N_13094);
xnor U13279 (N_13279,N_13106,N_12948);
xnor U13280 (N_13280,N_12917,N_12851);
nor U13281 (N_13281,N_13039,N_13026);
and U13282 (N_13282,N_12898,N_13061);
nand U13283 (N_13283,N_13187,N_13024);
nor U13284 (N_13284,N_13146,N_13021);
nor U13285 (N_13285,N_13138,N_13100);
or U13286 (N_13286,N_13181,N_12971);
and U13287 (N_13287,N_12837,N_12878);
and U13288 (N_13288,N_13030,N_13085);
nand U13289 (N_13289,N_13148,N_12873);
and U13290 (N_13290,N_12960,N_12969);
xnor U13291 (N_13291,N_12801,N_12962);
and U13292 (N_13292,N_12965,N_13175);
or U13293 (N_13293,N_12905,N_13133);
or U13294 (N_13294,N_13102,N_13050);
or U13295 (N_13295,N_12995,N_13004);
or U13296 (N_13296,N_13118,N_13158);
nand U13297 (N_13297,N_12925,N_12968);
xor U13298 (N_13298,N_13130,N_13190);
and U13299 (N_13299,N_12922,N_13011);
nand U13300 (N_13300,N_12936,N_13073);
or U13301 (N_13301,N_12821,N_12811);
nand U13302 (N_13302,N_12868,N_13143);
nand U13303 (N_13303,N_13186,N_13185);
or U13304 (N_13304,N_13062,N_13018);
or U13305 (N_13305,N_12918,N_13058);
or U13306 (N_13306,N_12831,N_13198);
nor U13307 (N_13307,N_12846,N_12986);
xor U13308 (N_13308,N_12928,N_12886);
xor U13309 (N_13309,N_12982,N_13012);
nand U13310 (N_13310,N_13132,N_13003);
nor U13311 (N_13311,N_13020,N_12804);
xnor U13312 (N_13312,N_13199,N_12863);
or U13313 (N_13313,N_12877,N_12875);
nor U13314 (N_13314,N_12983,N_13150);
nor U13315 (N_13315,N_13145,N_13056);
or U13316 (N_13316,N_12990,N_12926);
nor U13317 (N_13317,N_13060,N_13116);
nand U13318 (N_13318,N_13154,N_12864);
or U13319 (N_13319,N_13014,N_13095);
or U13320 (N_13320,N_12810,N_12911);
xnor U13321 (N_13321,N_12870,N_12856);
xnor U13322 (N_13322,N_12992,N_13177);
or U13323 (N_13323,N_12892,N_13079);
nor U13324 (N_13324,N_13169,N_12947);
and U13325 (N_13325,N_13027,N_12993);
nand U13326 (N_13326,N_13166,N_13196);
xnor U13327 (N_13327,N_13040,N_12808);
nor U13328 (N_13328,N_12903,N_13164);
xnor U13329 (N_13329,N_13160,N_12927);
nor U13330 (N_13330,N_13178,N_12880);
nand U13331 (N_13331,N_12953,N_12823);
xor U13332 (N_13332,N_12954,N_13193);
or U13333 (N_13333,N_13002,N_12978);
nand U13334 (N_13334,N_13007,N_13159);
or U13335 (N_13335,N_12860,N_13070);
or U13336 (N_13336,N_13161,N_12895);
nor U13337 (N_13337,N_12910,N_12951);
nand U13338 (N_13338,N_12874,N_12847);
nor U13339 (N_13339,N_13057,N_13162);
or U13340 (N_13340,N_12871,N_13117);
and U13341 (N_13341,N_12887,N_12952);
or U13342 (N_13342,N_13032,N_12825);
xor U13343 (N_13343,N_13105,N_12956);
nand U13344 (N_13344,N_13191,N_13182);
nand U13345 (N_13345,N_13006,N_12885);
nand U13346 (N_13346,N_12958,N_13051);
nand U13347 (N_13347,N_13048,N_13125);
nor U13348 (N_13348,N_13063,N_12852);
xnor U13349 (N_13349,N_13036,N_12813);
xor U13350 (N_13350,N_13124,N_13044);
nor U13351 (N_13351,N_12865,N_12989);
xnor U13352 (N_13352,N_13034,N_12980);
and U13353 (N_13353,N_13008,N_13144);
xor U13354 (N_13354,N_12872,N_13038);
nand U13355 (N_13355,N_13149,N_13052);
or U13356 (N_13356,N_12915,N_13195);
xor U13357 (N_13357,N_12974,N_12973);
xnor U13358 (N_13358,N_12824,N_13089);
or U13359 (N_13359,N_12832,N_12933);
or U13360 (N_13360,N_12889,N_13055);
nor U13361 (N_13361,N_12862,N_12991);
xnor U13362 (N_13362,N_13015,N_13126);
xor U13363 (N_13363,N_13110,N_13096);
and U13364 (N_13364,N_13049,N_12914);
and U13365 (N_13365,N_13184,N_12897);
and U13366 (N_13366,N_12888,N_13127);
or U13367 (N_13367,N_13129,N_12861);
and U13368 (N_13368,N_13077,N_13023);
xor U13369 (N_13369,N_12944,N_13082);
nor U13370 (N_13370,N_13173,N_13189);
nand U13371 (N_13371,N_12935,N_13156);
xor U13372 (N_13372,N_12866,N_12929);
xor U13373 (N_13373,N_12890,N_12853);
xor U13374 (N_13374,N_12967,N_12901);
xor U13375 (N_13375,N_12945,N_13103);
and U13376 (N_13376,N_13009,N_12820);
or U13377 (N_13377,N_12815,N_13113);
xor U13378 (N_13378,N_13086,N_12977);
nand U13379 (N_13379,N_12843,N_13065);
or U13380 (N_13380,N_12883,N_12988);
and U13381 (N_13381,N_13067,N_12839);
xnor U13382 (N_13382,N_13104,N_13005);
nor U13383 (N_13383,N_12816,N_12876);
nor U13384 (N_13384,N_12838,N_13176);
nand U13385 (N_13385,N_12906,N_12835);
xnor U13386 (N_13386,N_12949,N_12950);
or U13387 (N_13387,N_13108,N_12859);
or U13388 (N_13388,N_13033,N_12930);
xor U13389 (N_13389,N_13122,N_13153);
nand U13390 (N_13390,N_13099,N_13197);
or U13391 (N_13391,N_13134,N_12920);
and U13392 (N_13392,N_13109,N_12902);
xnor U13393 (N_13393,N_12819,N_13137);
nand U13394 (N_13394,N_13192,N_12938);
or U13395 (N_13395,N_12850,N_13066);
nor U13396 (N_13396,N_12806,N_12979);
and U13397 (N_13397,N_12844,N_12912);
nand U13398 (N_13398,N_13141,N_12900);
xor U13399 (N_13399,N_12964,N_13112);
nand U13400 (N_13400,N_12956,N_12849);
or U13401 (N_13401,N_12850,N_13132);
and U13402 (N_13402,N_13013,N_12868);
and U13403 (N_13403,N_12811,N_13108);
and U13404 (N_13404,N_13132,N_12961);
xor U13405 (N_13405,N_12921,N_12938);
xnor U13406 (N_13406,N_12904,N_13106);
nand U13407 (N_13407,N_13033,N_13056);
or U13408 (N_13408,N_13183,N_12989);
and U13409 (N_13409,N_13142,N_13009);
nand U13410 (N_13410,N_12841,N_12981);
nand U13411 (N_13411,N_12865,N_13171);
nor U13412 (N_13412,N_12853,N_12921);
and U13413 (N_13413,N_12865,N_12803);
xor U13414 (N_13414,N_13124,N_13061);
or U13415 (N_13415,N_13084,N_13075);
nand U13416 (N_13416,N_12826,N_13080);
or U13417 (N_13417,N_12943,N_12950);
nand U13418 (N_13418,N_12887,N_12825);
nand U13419 (N_13419,N_13040,N_12820);
nor U13420 (N_13420,N_12847,N_13117);
or U13421 (N_13421,N_13141,N_12912);
nand U13422 (N_13422,N_12940,N_13064);
xnor U13423 (N_13423,N_13161,N_12932);
nor U13424 (N_13424,N_13059,N_13081);
and U13425 (N_13425,N_13030,N_12873);
or U13426 (N_13426,N_13016,N_13167);
xnor U13427 (N_13427,N_13143,N_12844);
and U13428 (N_13428,N_13004,N_13018);
xnor U13429 (N_13429,N_13175,N_13007);
nor U13430 (N_13430,N_12821,N_12946);
and U13431 (N_13431,N_13140,N_13003);
nor U13432 (N_13432,N_13080,N_12809);
xor U13433 (N_13433,N_12873,N_13169);
nand U13434 (N_13434,N_12877,N_12918);
or U13435 (N_13435,N_13045,N_13177);
nor U13436 (N_13436,N_13183,N_13051);
and U13437 (N_13437,N_12968,N_12906);
or U13438 (N_13438,N_13047,N_13068);
and U13439 (N_13439,N_13126,N_13007);
nor U13440 (N_13440,N_12966,N_12829);
nor U13441 (N_13441,N_12980,N_13179);
xor U13442 (N_13442,N_12966,N_12801);
and U13443 (N_13443,N_12891,N_13079);
or U13444 (N_13444,N_12944,N_13189);
nor U13445 (N_13445,N_12810,N_13051);
nor U13446 (N_13446,N_12992,N_13159);
nand U13447 (N_13447,N_13164,N_12875);
xor U13448 (N_13448,N_13128,N_12930);
or U13449 (N_13449,N_13006,N_13082);
nand U13450 (N_13450,N_12808,N_13005);
xor U13451 (N_13451,N_13170,N_12857);
and U13452 (N_13452,N_12854,N_13189);
or U13453 (N_13453,N_13172,N_13106);
nand U13454 (N_13454,N_13019,N_12812);
nor U13455 (N_13455,N_13070,N_12986);
and U13456 (N_13456,N_12980,N_12942);
nand U13457 (N_13457,N_12985,N_12852);
or U13458 (N_13458,N_13155,N_13176);
xnor U13459 (N_13459,N_13071,N_12996);
or U13460 (N_13460,N_12999,N_13011);
xnor U13461 (N_13461,N_12876,N_12885);
nor U13462 (N_13462,N_12971,N_12941);
xor U13463 (N_13463,N_12808,N_13148);
or U13464 (N_13464,N_13087,N_12812);
or U13465 (N_13465,N_12918,N_13158);
or U13466 (N_13466,N_12976,N_13000);
and U13467 (N_13467,N_13063,N_13114);
xnor U13468 (N_13468,N_13110,N_13078);
or U13469 (N_13469,N_13150,N_13151);
or U13470 (N_13470,N_13151,N_12814);
xor U13471 (N_13471,N_13123,N_12888);
or U13472 (N_13472,N_12987,N_12952);
xnor U13473 (N_13473,N_13090,N_13155);
nor U13474 (N_13474,N_12873,N_12926);
nor U13475 (N_13475,N_13050,N_13181);
nor U13476 (N_13476,N_13079,N_12840);
nor U13477 (N_13477,N_13165,N_13071);
xnor U13478 (N_13478,N_12997,N_12992);
and U13479 (N_13479,N_13182,N_12959);
or U13480 (N_13480,N_12966,N_12936);
nor U13481 (N_13481,N_12819,N_12878);
nand U13482 (N_13482,N_13081,N_12943);
nand U13483 (N_13483,N_12977,N_13153);
xnor U13484 (N_13484,N_13118,N_12872);
nand U13485 (N_13485,N_13183,N_13149);
xnor U13486 (N_13486,N_13153,N_12902);
nand U13487 (N_13487,N_13163,N_13088);
nand U13488 (N_13488,N_12941,N_13092);
xnor U13489 (N_13489,N_13111,N_12981);
or U13490 (N_13490,N_12944,N_13006);
nand U13491 (N_13491,N_13065,N_12803);
xnor U13492 (N_13492,N_12974,N_13049);
and U13493 (N_13493,N_13057,N_13166);
xor U13494 (N_13494,N_13154,N_12966);
nor U13495 (N_13495,N_13080,N_13065);
or U13496 (N_13496,N_13151,N_12934);
xor U13497 (N_13497,N_12813,N_12840);
nand U13498 (N_13498,N_13029,N_13154);
and U13499 (N_13499,N_12901,N_12991);
nand U13500 (N_13500,N_13152,N_13030);
nor U13501 (N_13501,N_13132,N_13125);
and U13502 (N_13502,N_13126,N_13028);
or U13503 (N_13503,N_12917,N_13189);
and U13504 (N_13504,N_13174,N_12896);
or U13505 (N_13505,N_12891,N_12953);
xor U13506 (N_13506,N_12928,N_13022);
or U13507 (N_13507,N_12960,N_12988);
nor U13508 (N_13508,N_13025,N_12874);
nor U13509 (N_13509,N_13049,N_13003);
xnor U13510 (N_13510,N_12932,N_13083);
or U13511 (N_13511,N_13098,N_13045);
and U13512 (N_13512,N_13041,N_13021);
xnor U13513 (N_13513,N_12890,N_13047);
or U13514 (N_13514,N_12914,N_12888);
xnor U13515 (N_13515,N_12867,N_12906);
or U13516 (N_13516,N_13028,N_13065);
and U13517 (N_13517,N_13158,N_12943);
nor U13518 (N_13518,N_12812,N_13031);
nand U13519 (N_13519,N_12841,N_13005);
and U13520 (N_13520,N_12808,N_13032);
nor U13521 (N_13521,N_12938,N_13006);
or U13522 (N_13522,N_12890,N_13157);
xor U13523 (N_13523,N_13116,N_12885);
nand U13524 (N_13524,N_12839,N_12925);
or U13525 (N_13525,N_12984,N_12925);
nand U13526 (N_13526,N_12877,N_13118);
nand U13527 (N_13527,N_12989,N_12828);
and U13528 (N_13528,N_13198,N_12951);
and U13529 (N_13529,N_13182,N_12839);
or U13530 (N_13530,N_13111,N_12826);
xnor U13531 (N_13531,N_13062,N_13198);
and U13532 (N_13532,N_13040,N_13121);
and U13533 (N_13533,N_13091,N_12972);
and U13534 (N_13534,N_13070,N_13170);
nand U13535 (N_13535,N_13177,N_12951);
xor U13536 (N_13536,N_12822,N_12866);
nand U13537 (N_13537,N_13048,N_12876);
nand U13538 (N_13538,N_12951,N_13082);
nor U13539 (N_13539,N_13182,N_13144);
nand U13540 (N_13540,N_12831,N_12998);
and U13541 (N_13541,N_13193,N_12905);
or U13542 (N_13542,N_12988,N_13167);
nand U13543 (N_13543,N_13013,N_13018);
or U13544 (N_13544,N_13159,N_12847);
and U13545 (N_13545,N_13136,N_13024);
or U13546 (N_13546,N_12969,N_12883);
nand U13547 (N_13547,N_13033,N_13057);
or U13548 (N_13548,N_12951,N_13042);
xor U13549 (N_13549,N_13114,N_13127);
nor U13550 (N_13550,N_13164,N_13028);
and U13551 (N_13551,N_12838,N_12936);
and U13552 (N_13552,N_13150,N_13128);
nand U13553 (N_13553,N_13174,N_12908);
or U13554 (N_13554,N_13025,N_13167);
or U13555 (N_13555,N_12980,N_12907);
and U13556 (N_13556,N_12997,N_13129);
xor U13557 (N_13557,N_13077,N_13062);
xor U13558 (N_13558,N_13198,N_12820);
xor U13559 (N_13559,N_12901,N_12871);
and U13560 (N_13560,N_13154,N_12805);
nand U13561 (N_13561,N_13125,N_12890);
xor U13562 (N_13562,N_13041,N_12853);
or U13563 (N_13563,N_12852,N_12906);
nand U13564 (N_13564,N_12903,N_12906);
and U13565 (N_13565,N_12832,N_13190);
or U13566 (N_13566,N_12825,N_12998);
xnor U13567 (N_13567,N_12899,N_12801);
nor U13568 (N_13568,N_12891,N_13198);
nor U13569 (N_13569,N_12838,N_12960);
and U13570 (N_13570,N_12849,N_13193);
xnor U13571 (N_13571,N_12849,N_13039);
and U13572 (N_13572,N_12823,N_13016);
nand U13573 (N_13573,N_13137,N_13160);
nand U13574 (N_13574,N_12988,N_13186);
xnor U13575 (N_13575,N_12876,N_13178);
or U13576 (N_13576,N_13192,N_12906);
nand U13577 (N_13577,N_12826,N_13192);
or U13578 (N_13578,N_13159,N_12872);
xnor U13579 (N_13579,N_12903,N_12881);
nand U13580 (N_13580,N_13129,N_13142);
nand U13581 (N_13581,N_13037,N_13035);
or U13582 (N_13582,N_12907,N_12941);
or U13583 (N_13583,N_13182,N_13159);
and U13584 (N_13584,N_13197,N_12929);
and U13585 (N_13585,N_13038,N_13126);
or U13586 (N_13586,N_13110,N_13189);
xor U13587 (N_13587,N_13187,N_13146);
xnor U13588 (N_13588,N_13136,N_13008);
nor U13589 (N_13589,N_13050,N_13063);
or U13590 (N_13590,N_12879,N_12825);
xnor U13591 (N_13591,N_13198,N_12804);
and U13592 (N_13592,N_12995,N_12945);
and U13593 (N_13593,N_13041,N_13163);
nand U13594 (N_13594,N_13063,N_13077);
or U13595 (N_13595,N_12844,N_13156);
nand U13596 (N_13596,N_13113,N_12971);
and U13597 (N_13597,N_12904,N_12909);
xnor U13598 (N_13598,N_13125,N_13056);
xor U13599 (N_13599,N_12981,N_13061);
and U13600 (N_13600,N_13494,N_13314);
nor U13601 (N_13601,N_13414,N_13293);
and U13602 (N_13602,N_13589,N_13592);
nand U13603 (N_13603,N_13391,N_13245);
nor U13604 (N_13604,N_13450,N_13436);
nor U13605 (N_13605,N_13231,N_13473);
and U13606 (N_13606,N_13484,N_13270);
or U13607 (N_13607,N_13254,N_13580);
nand U13608 (N_13608,N_13476,N_13407);
nor U13609 (N_13609,N_13576,N_13572);
nor U13610 (N_13610,N_13218,N_13405);
nor U13611 (N_13611,N_13243,N_13328);
nor U13612 (N_13612,N_13297,N_13581);
or U13613 (N_13613,N_13275,N_13377);
xnor U13614 (N_13614,N_13406,N_13345);
and U13615 (N_13615,N_13442,N_13499);
nor U13616 (N_13616,N_13444,N_13514);
xor U13617 (N_13617,N_13467,N_13493);
nor U13618 (N_13618,N_13252,N_13353);
or U13619 (N_13619,N_13224,N_13417);
or U13620 (N_13620,N_13479,N_13287);
nand U13621 (N_13621,N_13438,N_13336);
xnor U13622 (N_13622,N_13378,N_13472);
nand U13623 (N_13623,N_13273,N_13216);
xor U13624 (N_13624,N_13430,N_13382);
nor U13625 (N_13625,N_13540,N_13329);
or U13626 (N_13626,N_13221,N_13244);
and U13627 (N_13627,N_13211,N_13453);
or U13628 (N_13628,N_13352,N_13338);
nor U13629 (N_13629,N_13300,N_13586);
and U13630 (N_13630,N_13209,N_13385);
and U13631 (N_13631,N_13542,N_13400);
nand U13632 (N_13632,N_13319,N_13220);
xnor U13633 (N_13633,N_13529,N_13236);
xnor U13634 (N_13634,N_13553,N_13272);
xor U13635 (N_13635,N_13262,N_13235);
nand U13636 (N_13636,N_13390,N_13585);
xnor U13637 (N_13637,N_13298,N_13375);
nor U13638 (N_13638,N_13555,N_13266);
xor U13639 (N_13639,N_13426,N_13452);
and U13640 (N_13640,N_13318,N_13461);
or U13641 (N_13641,N_13348,N_13276);
and U13642 (N_13642,N_13310,N_13408);
xnor U13643 (N_13643,N_13441,N_13564);
or U13644 (N_13644,N_13487,N_13501);
or U13645 (N_13645,N_13371,N_13360);
and U13646 (N_13646,N_13343,N_13420);
and U13647 (N_13647,N_13474,N_13544);
nor U13648 (N_13648,N_13491,N_13361);
xnor U13649 (N_13649,N_13478,N_13289);
nand U13650 (N_13650,N_13448,N_13306);
and U13651 (N_13651,N_13471,N_13554);
xnor U13652 (N_13652,N_13323,N_13455);
or U13653 (N_13653,N_13446,N_13296);
and U13654 (N_13654,N_13206,N_13295);
and U13655 (N_13655,N_13340,N_13435);
or U13656 (N_13656,N_13324,N_13258);
nor U13657 (N_13657,N_13482,N_13409);
and U13658 (N_13658,N_13341,N_13590);
xnor U13659 (N_13659,N_13237,N_13480);
xnor U13660 (N_13660,N_13278,N_13233);
xnor U13661 (N_13661,N_13366,N_13465);
nor U13662 (N_13662,N_13519,N_13508);
and U13663 (N_13663,N_13416,N_13239);
and U13664 (N_13664,N_13565,N_13412);
nand U13665 (N_13665,N_13477,N_13264);
xor U13666 (N_13666,N_13546,N_13411);
nor U13667 (N_13667,N_13528,N_13563);
xnor U13668 (N_13668,N_13304,N_13517);
nand U13669 (N_13669,N_13434,N_13463);
and U13670 (N_13670,N_13315,N_13579);
and U13671 (N_13671,N_13305,N_13568);
and U13672 (N_13672,N_13432,N_13227);
and U13673 (N_13673,N_13556,N_13200);
nor U13674 (N_13674,N_13202,N_13561);
xnor U13675 (N_13675,N_13303,N_13279);
or U13676 (N_13676,N_13524,N_13458);
and U13677 (N_13677,N_13373,N_13204);
xor U13678 (N_13678,N_13531,N_13316);
and U13679 (N_13679,N_13368,N_13380);
and U13680 (N_13680,N_13357,N_13515);
nor U13681 (N_13681,N_13466,N_13229);
xor U13682 (N_13682,N_13427,N_13238);
nor U13683 (N_13683,N_13285,N_13331);
nor U13684 (N_13684,N_13396,N_13267);
or U13685 (N_13685,N_13538,N_13386);
nand U13686 (N_13686,N_13381,N_13510);
or U13687 (N_13687,N_13559,N_13313);
nand U13688 (N_13688,N_13212,N_13440);
nor U13689 (N_13689,N_13454,N_13537);
nor U13690 (N_13690,N_13376,N_13349);
or U13691 (N_13691,N_13443,N_13261);
nor U13692 (N_13692,N_13469,N_13549);
xnor U13693 (N_13693,N_13251,N_13277);
nor U13694 (N_13694,N_13535,N_13219);
and U13695 (N_13695,N_13367,N_13523);
xnor U13696 (N_13696,N_13439,N_13288);
and U13697 (N_13697,N_13370,N_13397);
nand U13698 (N_13698,N_13228,N_13525);
xor U13699 (N_13699,N_13225,N_13539);
nor U13700 (N_13700,N_13424,N_13560);
nand U13701 (N_13701,N_13398,N_13488);
xor U13702 (N_13702,N_13223,N_13240);
and U13703 (N_13703,N_13207,N_13203);
nor U13704 (N_13704,N_13536,N_13374);
and U13705 (N_13705,N_13392,N_13337);
nand U13706 (N_13706,N_13363,N_13326);
xnor U13707 (N_13707,N_13583,N_13505);
nand U13708 (N_13708,N_13595,N_13578);
nand U13709 (N_13709,N_13246,N_13299);
and U13710 (N_13710,N_13213,N_13317);
and U13711 (N_13711,N_13460,N_13507);
or U13712 (N_13712,N_13489,N_13372);
or U13713 (N_13713,N_13562,N_13521);
and U13714 (N_13714,N_13362,N_13445);
nand U13715 (N_13715,N_13526,N_13567);
nor U13716 (N_13716,N_13545,N_13513);
xnor U13717 (N_13717,N_13571,N_13419);
xnor U13718 (N_13718,N_13355,N_13551);
nand U13719 (N_13719,N_13451,N_13506);
or U13720 (N_13720,N_13543,N_13350);
xnor U13721 (N_13721,N_13587,N_13573);
xor U13722 (N_13722,N_13201,N_13582);
xnor U13723 (N_13723,N_13271,N_13259);
xor U13724 (N_13724,N_13230,N_13500);
nor U13725 (N_13725,N_13599,N_13558);
or U13726 (N_13726,N_13356,N_13344);
nand U13727 (N_13727,N_13394,N_13308);
or U13728 (N_13728,N_13403,N_13208);
xnor U13729 (N_13729,N_13301,N_13257);
nor U13730 (N_13730,N_13312,N_13292);
or U13731 (N_13731,N_13483,N_13512);
or U13732 (N_13732,N_13268,N_13459);
and U13733 (N_13733,N_13541,N_13332);
nor U13734 (N_13734,N_13504,N_13388);
nand U13735 (N_13735,N_13234,N_13548);
xnor U13736 (N_13736,N_13418,N_13214);
and U13737 (N_13737,N_13347,N_13248);
nand U13738 (N_13738,N_13509,N_13522);
or U13739 (N_13739,N_13263,N_13247);
or U13740 (N_13740,N_13456,N_13596);
or U13741 (N_13741,N_13311,N_13335);
nand U13742 (N_13742,N_13320,N_13433);
nor U13743 (N_13743,N_13282,N_13333);
xor U13744 (N_13744,N_13379,N_13395);
and U13745 (N_13745,N_13401,N_13533);
nand U13746 (N_13746,N_13283,N_13250);
nor U13747 (N_13747,N_13413,N_13294);
or U13748 (N_13748,N_13437,N_13410);
xnor U13749 (N_13749,N_13232,N_13569);
xnor U13750 (N_13750,N_13428,N_13475);
nand U13751 (N_13751,N_13566,N_13534);
nor U13752 (N_13752,N_13364,N_13217);
and U13753 (N_13753,N_13584,N_13346);
or U13754 (N_13754,N_13286,N_13389);
or U13755 (N_13755,N_13290,N_13594);
and U13756 (N_13756,N_13518,N_13342);
nand U13757 (N_13757,N_13325,N_13485);
nand U13758 (N_13758,N_13447,N_13574);
xor U13759 (N_13759,N_13492,N_13423);
and U13760 (N_13760,N_13253,N_13365);
or U13761 (N_13761,N_13588,N_13557);
nor U13762 (N_13762,N_13486,N_13511);
or U13763 (N_13763,N_13280,N_13242);
xor U13764 (N_13764,N_13358,N_13498);
or U13765 (N_13765,N_13481,N_13383);
nor U13766 (N_13766,N_13321,N_13520);
and U13767 (N_13767,N_13496,N_13334);
nor U13768 (N_13768,N_13330,N_13291);
and U13769 (N_13769,N_13393,N_13402);
nand U13770 (N_13770,N_13449,N_13265);
nor U13771 (N_13771,N_13249,N_13339);
or U13772 (N_13772,N_13577,N_13547);
or U13773 (N_13773,N_13255,N_13597);
or U13774 (N_13774,N_13495,N_13354);
nand U13775 (N_13775,N_13274,N_13415);
nand U13776 (N_13776,N_13470,N_13490);
and U13777 (N_13777,N_13497,N_13302);
nor U13778 (N_13778,N_13241,N_13205);
and U13779 (N_13779,N_13256,N_13457);
xnor U13780 (N_13780,N_13550,N_13421);
nand U13781 (N_13781,N_13269,N_13322);
or U13782 (N_13782,N_13307,N_13575);
nand U13783 (N_13783,N_13351,N_13260);
xnor U13784 (N_13784,N_13210,N_13359);
nand U13785 (N_13785,N_13384,N_13399);
or U13786 (N_13786,N_13502,N_13570);
nor U13787 (N_13787,N_13222,N_13281);
nand U13788 (N_13788,N_13425,N_13429);
or U13789 (N_13789,N_13462,N_13369);
xnor U13790 (N_13790,N_13284,N_13591);
and U13791 (N_13791,N_13226,N_13552);
nor U13792 (N_13792,N_13464,N_13530);
nand U13793 (N_13793,N_13215,N_13598);
nor U13794 (N_13794,N_13309,N_13327);
and U13795 (N_13795,N_13503,N_13387);
nor U13796 (N_13796,N_13431,N_13404);
or U13797 (N_13797,N_13593,N_13532);
nor U13798 (N_13798,N_13516,N_13422);
or U13799 (N_13799,N_13468,N_13527);
nand U13800 (N_13800,N_13543,N_13303);
and U13801 (N_13801,N_13279,N_13560);
nor U13802 (N_13802,N_13395,N_13214);
and U13803 (N_13803,N_13543,N_13330);
xor U13804 (N_13804,N_13235,N_13596);
xor U13805 (N_13805,N_13487,N_13267);
and U13806 (N_13806,N_13266,N_13564);
nor U13807 (N_13807,N_13212,N_13510);
nor U13808 (N_13808,N_13387,N_13392);
or U13809 (N_13809,N_13489,N_13339);
xnor U13810 (N_13810,N_13314,N_13335);
or U13811 (N_13811,N_13303,N_13338);
or U13812 (N_13812,N_13538,N_13360);
xor U13813 (N_13813,N_13386,N_13432);
nor U13814 (N_13814,N_13280,N_13532);
nand U13815 (N_13815,N_13257,N_13559);
xor U13816 (N_13816,N_13315,N_13484);
and U13817 (N_13817,N_13461,N_13201);
nor U13818 (N_13818,N_13261,N_13338);
nor U13819 (N_13819,N_13308,N_13435);
xor U13820 (N_13820,N_13374,N_13223);
or U13821 (N_13821,N_13223,N_13408);
nor U13822 (N_13822,N_13359,N_13227);
and U13823 (N_13823,N_13356,N_13515);
nor U13824 (N_13824,N_13570,N_13568);
and U13825 (N_13825,N_13572,N_13499);
xor U13826 (N_13826,N_13228,N_13572);
xnor U13827 (N_13827,N_13502,N_13488);
or U13828 (N_13828,N_13462,N_13263);
and U13829 (N_13829,N_13294,N_13550);
and U13830 (N_13830,N_13515,N_13376);
nand U13831 (N_13831,N_13222,N_13217);
xnor U13832 (N_13832,N_13426,N_13598);
or U13833 (N_13833,N_13216,N_13435);
nor U13834 (N_13834,N_13440,N_13377);
or U13835 (N_13835,N_13448,N_13336);
nor U13836 (N_13836,N_13296,N_13524);
or U13837 (N_13837,N_13200,N_13555);
and U13838 (N_13838,N_13311,N_13426);
or U13839 (N_13839,N_13510,N_13452);
xnor U13840 (N_13840,N_13482,N_13282);
and U13841 (N_13841,N_13577,N_13484);
nor U13842 (N_13842,N_13599,N_13483);
xnor U13843 (N_13843,N_13386,N_13340);
nand U13844 (N_13844,N_13372,N_13555);
nor U13845 (N_13845,N_13478,N_13551);
xnor U13846 (N_13846,N_13408,N_13339);
or U13847 (N_13847,N_13364,N_13427);
or U13848 (N_13848,N_13416,N_13231);
nand U13849 (N_13849,N_13500,N_13579);
or U13850 (N_13850,N_13384,N_13469);
nor U13851 (N_13851,N_13481,N_13405);
xnor U13852 (N_13852,N_13220,N_13340);
nand U13853 (N_13853,N_13395,N_13264);
and U13854 (N_13854,N_13335,N_13493);
and U13855 (N_13855,N_13398,N_13227);
xnor U13856 (N_13856,N_13344,N_13387);
or U13857 (N_13857,N_13537,N_13382);
xor U13858 (N_13858,N_13473,N_13212);
and U13859 (N_13859,N_13308,N_13319);
nand U13860 (N_13860,N_13539,N_13320);
nor U13861 (N_13861,N_13353,N_13571);
nand U13862 (N_13862,N_13578,N_13486);
or U13863 (N_13863,N_13318,N_13433);
xnor U13864 (N_13864,N_13525,N_13259);
nand U13865 (N_13865,N_13348,N_13223);
or U13866 (N_13866,N_13474,N_13577);
and U13867 (N_13867,N_13526,N_13204);
xnor U13868 (N_13868,N_13568,N_13282);
or U13869 (N_13869,N_13267,N_13456);
and U13870 (N_13870,N_13242,N_13269);
xnor U13871 (N_13871,N_13266,N_13228);
nand U13872 (N_13872,N_13272,N_13238);
nand U13873 (N_13873,N_13496,N_13500);
nor U13874 (N_13874,N_13341,N_13524);
xor U13875 (N_13875,N_13441,N_13439);
and U13876 (N_13876,N_13350,N_13267);
and U13877 (N_13877,N_13429,N_13375);
xor U13878 (N_13878,N_13239,N_13465);
nor U13879 (N_13879,N_13403,N_13418);
nand U13880 (N_13880,N_13276,N_13254);
or U13881 (N_13881,N_13439,N_13307);
or U13882 (N_13882,N_13343,N_13583);
xnor U13883 (N_13883,N_13550,N_13248);
and U13884 (N_13884,N_13401,N_13555);
and U13885 (N_13885,N_13212,N_13481);
or U13886 (N_13886,N_13259,N_13505);
xnor U13887 (N_13887,N_13409,N_13475);
and U13888 (N_13888,N_13306,N_13345);
xor U13889 (N_13889,N_13597,N_13535);
and U13890 (N_13890,N_13362,N_13475);
or U13891 (N_13891,N_13358,N_13260);
nand U13892 (N_13892,N_13562,N_13441);
nand U13893 (N_13893,N_13561,N_13346);
or U13894 (N_13894,N_13488,N_13357);
and U13895 (N_13895,N_13345,N_13224);
nor U13896 (N_13896,N_13398,N_13505);
nand U13897 (N_13897,N_13269,N_13550);
nand U13898 (N_13898,N_13491,N_13397);
xor U13899 (N_13899,N_13415,N_13303);
and U13900 (N_13900,N_13486,N_13537);
and U13901 (N_13901,N_13305,N_13253);
nand U13902 (N_13902,N_13249,N_13235);
xnor U13903 (N_13903,N_13440,N_13328);
nand U13904 (N_13904,N_13493,N_13286);
nor U13905 (N_13905,N_13237,N_13549);
and U13906 (N_13906,N_13515,N_13355);
and U13907 (N_13907,N_13587,N_13325);
and U13908 (N_13908,N_13522,N_13389);
nor U13909 (N_13909,N_13239,N_13364);
nand U13910 (N_13910,N_13291,N_13451);
and U13911 (N_13911,N_13226,N_13314);
and U13912 (N_13912,N_13278,N_13434);
xor U13913 (N_13913,N_13375,N_13407);
xnor U13914 (N_13914,N_13557,N_13567);
or U13915 (N_13915,N_13567,N_13298);
nor U13916 (N_13916,N_13281,N_13408);
xnor U13917 (N_13917,N_13309,N_13405);
nor U13918 (N_13918,N_13564,N_13419);
and U13919 (N_13919,N_13255,N_13317);
nand U13920 (N_13920,N_13357,N_13312);
or U13921 (N_13921,N_13249,N_13322);
and U13922 (N_13922,N_13456,N_13539);
xor U13923 (N_13923,N_13266,N_13417);
nand U13924 (N_13924,N_13274,N_13506);
xor U13925 (N_13925,N_13322,N_13398);
or U13926 (N_13926,N_13284,N_13397);
or U13927 (N_13927,N_13584,N_13447);
nand U13928 (N_13928,N_13236,N_13526);
xnor U13929 (N_13929,N_13408,N_13446);
or U13930 (N_13930,N_13201,N_13332);
nor U13931 (N_13931,N_13353,N_13549);
xnor U13932 (N_13932,N_13312,N_13572);
or U13933 (N_13933,N_13341,N_13516);
nor U13934 (N_13934,N_13576,N_13304);
nor U13935 (N_13935,N_13506,N_13351);
nand U13936 (N_13936,N_13523,N_13211);
or U13937 (N_13937,N_13471,N_13319);
or U13938 (N_13938,N_13446,N_13280);
nand U13939 (N_13939,N_13261,N_13572);
or U13940 (N_13940,N_13573,N_13456);
nor U13941 (N_13941,N_13315,N_13221);
nor U13942 (N_13942,N_13411,N_13208);
and U13943 (N_13943,N_13231,N_13314);
nand U13944 (N_13944,N_13352,N_13444);
nand U13945 (N_13945,N_13287,N_13504);
and U13946 (N_13946,N_13414,N_13555);
nor U13947 (N_13947,N_13354,N_13223);
nor U13948 (N_13948,N_13549,N_13413);
and U13949 (N_13949,N_13244,N_13251);
nand U13950 (N_13950,N_13249,N_13410);
xnor U13951 (N_13951,N_13352,N_13579);
and U13952 (N_13952,N_13557,N_13521);
nand U13953 (N_13953,N_13530,N_13502);
nor U13954 (N_13954,N_13426,N_13475);
or U13955 (N_13955,N_13591,N_13581);
or U13956 (N_13956,N_13411,N_13353);
xor U13957 (N_13957,N_13491,N_13221);
and U13958 (N_13958,N_13522,N_13395);
nor U13959 (N_13959,N_13282,N_13403);
nor U13960 (N_13960,N_13275,N_13578);
xnor U13961 (N_13961,N_13394,N_13339);
nor U13962 (N_13962,N_13206,N_13501);
or U13963 (N_13963,N_13550,N_13501);
nor U13964 (N_13964,N_13235,N_13311);
or U13965 (N_13965,N_13533,N_13590);
xnor U13966 (N_13966,N_13225,N_13462);
xor U13967 (N_13967,N_13450,N_13400);
and U13968 (N_13968,N_13500,N_13382);
nor U13969 (N_13969,N_13384,N_13574);
nor U13970 (N_13970,N_13312,N_13406);
or U13971 (N_13971,N_13428,N_13286);
or U13972 (N_13972,N_13506,N_13516);
or U13973 (N_13973,N_13540,N_13328);
xor U13974 (N_13974,N_13353,N_13516);
or U13975 (N_13975,N_13466,N_13308);
nand U13976 (N_13976,N_13222,N_13504);
nor U13977 (N_13977,N_13585,N_13317);
and U13978 (N_13978,N_13446,N_13397);
xor U13979 (N_13979,N_13473,N_13478);
nor U13980 (N_13980,N_13504,N_13488);
or U13981 (N_13981,N_13452,N_13291);
xor U13982 (N_13982,N_13258,N_13373);
nand U13983 (N_13983,N_13349,N_13368);
nor U13984 (N_13984,N_13260,N_13314);
xor U13985 (N_13985,N_13402,N_13583);
nand U13986 (N_13986,N_13208,N_13372);
or U13987 (N_13987,N_13349,N_13458);
nand U13988 (N_13988,N_13562,N_13327);
or U13989 (N_13989,N_13225,N_13262);
or U13990 (N_13990,N_13510,N_13400);
or U13991 (N_13991,N_13575,N_13362);
xor U13992 (N_13992,N_13279,N_13238);
nand U13993 (N_13993,N_13539,N_13415);
nand U13994 (N_13994,N_13537,N_13433);
and U13995 (N_13995,N_13347,N_13228);
and U13996 (N_13996,N_13288,N_13410);
and U13997 (N_13997,N_13408,N_13257);
and U13998 (N_13998,N_13423,N_13548);
and U13999 (N_13999,N_13526,N_13469);
or U14000 (N_14000,N_13939,N_13987);
xor U14001 (N_14001,N_13941,N_13846);
nor U14002 (N_14002,N_13782,N_13823);
nand U14003 (N_14003,N_13955,N_13871);
nor U14004 (N_14004,N_13947,N_13818);
or U14005 (N_14005,N_13933,N_13935);
xor U14006 (N_14006,N_13805,N_13901);
nor U14007 (N_14007,N_13815,N_13793);
and U14008 (N_14008,N_13698,N_13876);
xnor U14009 (N_14009,N_13624,N_13739);
nor U14010 (N_14010,N_13796,N_13748);
nor U14011 (N_14011,N_13853,N_13865);
nor U14012 (N_14012,N_13714,N_13753);
nand U14013 (N_14013,N_13887,N_13663);
and U14014 (N_14014,N_13812,N_13828);
xnor U14015 (N_14015,N_13743,N_13689);
nand U14016 (N_14016,N_13655,N_13697);
and U14017 (N_14017,N_13731,N_13838);
xor U14018 (N_14018,N_13914,N_13756);
nand U14019 (N_14019,N_13958,N_13999);
xor U14020 (N_14020,N_13819,N_13722);
and U14021 (N_14021,N_13848,N_13826);
and U14022 (N_14022,N_13681,N_13735);
and U14023 (N_14023,N_13951,N_13686);
or U14024 (N_14024,N_13842,N_13621);
and U14025 (N_14025,N_13737,N_13769);
or U14026 (N_14026,N_13776,N_13789);
xnor U14027 (N_14027,N_13639,N_13705);
or U14028 (N_14028,N_13648,N_13626);
xnor U14029 (N_14029,N_13728,N_13924);
or U14030 (N_14030,N_13992,N_13725);
or U14031 (N_14031,N_13784,N_13980);
and U14032 (N_14032,N_13817,N_13618);
and U14033 (N_14033,N_13936,N_13970);
xor U14034 (N_14034,N_13844,N_13647);
and U14035 (N_14035,N_13858,N_13963);
nor U14036 (N_14036,N_13872,N_13931);
nor U14037 (N_14037,N_13726,N_13959);
nand U14038 (N_14038,N_13640,N_13813);
nand U14039 (N_14039,N_13800,N_13612);
or U14040 (N_14040,N_13617,N_13835);
and U14041 (N_14041,N_13915,N_13650);
nand U14042 (N_14042,N_13679,N_13688);
and U14043 (N_14043,N_13966,N_13710);
xnor U14044 (N_14044,N_13905,N_13913);
xor U14045 (N_14045,N_13691,N_13623);
xor U14046 (N_14046,N_13998,N_13867);
or U14047 (N_14047,N_13785,N_13696);
or U14048 (N_14048,N_13642,N_13934);
nand U14049 (N_14049,N_13615,N_13797);
xor U14050 (N_14050,N_13707,N_13897);
nand U14051 (N_14051,N_13600,N_13968);
xnor U14052 (N_14052,N_13902,N_13693);
and U14053 (N_14053,N_13699,N_13918);
and U14054 (N_14054,N_13669,N_13656);
and U14055 (N_14055,N_13622,N_13717);
xnor U14056 (N_14056,N_13795,N_13733);
and U14057 (N_14057,N_13907,N_13889);
nor U14058 (N_14058,N_13954,N_13984);
nor U14059 (N_14059,N_13874,N_13929);
nor U14060 (N_14060,N_13777,N_13685);
or U14061 (N_14061,N_13757,N_13709);
nand U14062 (N_14062,N_13940,N_13811);
or U14063 (N_14063,N_13899,N_13791);
xor U14064 (N_14064,N_13809,N_13900);
xor U14065 (N_14065,N_13744,N_13630);
nand U14066 (N_14066,N_13875,N_13896);
xor U14067 (N_14067,N_13781,N_13862);
xor U14068 (N_14068,N_13891,N_13657);
xnor U14069 (N_14069,N_13926,N_13711);
and U14070 (N_14070,N_13892,N_13943);
nor U14071 (N_14071,N_13879,N_13960);
nor U14072 (N_14072,N_13682,N_13665);
and U14073 (N_14073,N_13652,N_13773);
or U14074 (N_14074,N_13868,N_13917);
xor U14075 (N_14075,N_13834,N_13921);
nor U14076 (N_14076,N_13859,N_13604);
or U14077 (N_14077,N_13982,N_13827);
nor U14078 (N_14078,N_13990,N_13765);
xor U14079 (N_14079,N_13692,N_13856);
nand U14080 (N_14080,N_13978,N_13767);
or U14081 (N_14081,N_13863,N_13839);
or U14082 (N_14082,N_13690,N_13836);
xnor U14083 (N_14083,N_13830,N_13822);
nor U14084 (N_14084,N_13806,N_13721);
and U14085 (N_14085,N_13886,N_13677);
xnor U14086 (N_14086,N_13794,N_13651);
nand U14087 (N_14087,N_13723,N_13895);
xor U14088 (N_14088,N_13849,N_13649);
or U14089 (N_14089,N_13957,N_13882);
nand U14090 (N_14090,N_13625,N_13994);
nand U14091 (N_14091,N_13614,N_13755);
or U14092 (N_14092,N_13979,N_13949);
nand U14093 (N_14093,N_13798,N_13606);
nor U14094 (N_14094,N_13780,N_13724);
or U14095 (N_14095,N_13790,N_13802);
nor U14096 (N_14096,N_13973,N_13703);
or U14097 (N_14097,N_13683,N_13964);
nor U14098 (N_14098,N_13706,N_13734);
nor U14099 (N_14099,N_13632,N_13729);
xnor U14100 (N_14100,N_13909,N_13851);
or U14101 (N_14101,N_13713,N_13962);
xor U14102 (N_14102,N_13634,N_13788);
and U14103 (N_14103,N_13619,N_13991);
or U14104 (N_14104,N_13736,N_13730);
xor U14105 (N_14105,N_13923,N_13824);
xor U14106 (N_14106,N_13668,N_13661);
nand U14107 (N_14107,N_13602,N_13888);
or U14108 (N_14108,N_13832,N_13654);
nor U14109 (N_14109,N_13953,N_13814);
or U14110 (N_14110,N_13803,N_13673);
or U14111 (N_14111,N_13742,N_13660);
xnor U14112 (N_14112,N_13928,N_13760);
xor U14113 (N_14113,N_13870,N_13667);
xor U14114 (N_14114,N_13774,N_13631);
and U14115 (N_14115,N_13927,N_13971);
xnor U14116 (N_14116,N_13825,N_13873);
or U14117 (N_14117,N_13837,N_13976);
nor U14118 (N_14118,N_13664,N_13770);
nand U14119 (N_14119,N_13904,N_13993);
xor U14120 (N_14120,N_13855,N_13911);
nand U14121 (N_14121,N_13611,N_13629);
nand U14122 (N_14122,N_13799,N_13866);
xnor U14123 (N_14123,N_13861,N_13704);
nor U14124 (N_14124,N_13745,N_13759);
nand U14125 (N_14125,N_13845,N_13857);
nand U14126 (N_14126,N_13877,N_13938);
or U14127 (N_14127,N_13944,N_13718);
and U14128 (N_14128,N_13783,N_13792);
and U14129 (N_14129,N_13662,N_13684);
and U14130 (N_14130,N_13910,N_13981);
xor U14131 (N_14131,N_13620,N_13772);
and U14132 (N_14132,N_13658,N_13750);
and U14133 (N_14133,N_13925,N_13995);
and U14134 (N_14134,N_13674,N_13645);
nor U14135 (N_14135,N_13840,N_13961);
or U14136 (N_14136,N_13787,N_13956);
and U14137 (N_14137,N_13678,N_13820);
nand U14138 (N_14138,N_13860,N_13719);
or U14139 (N_14139,N_13628,N_13869);
or U14140 (N_14140,N_13644,N_13633);
nand U14141 (N_14141,N_13740,N_13680);
xnor U14142 (N_14142,N_13764,N_13942);
nor U14143 (N_14143,N_13930,N_13603);
and U14144 (N_14144,N_13779,N_13912);
and U14145 (N_14145,N_13808,N_13919);
nand U14146 (N_14146,N_13920,N_13937);
nand U14147 (N_14147,N_13771,N_13903);
nor U14148 (N_14148,N_13763,N_13701);
nor U14149 (N_14149,N_13786,N_13746);
xor U14150 (N_14150,N_13676,N_13801);
xor U14151 (N_14151,N_13885,N_13643);
xnor U14152 (N_14152,N_13616,N_13727);
xnor U14153 (N_14153,N_13670,N_13997);
nand U14154 (N_14154,N_13715,N_13607);
nor U14155 (N_14155,N_13945,N_13922);
nand U14156 (N_14156,N_13880,N_13687);
nor U14157 (N_14157,N_13601,N_13768);
nand U14158 (N_14158,N_13810,N_13636);
nand U14159 (N_14159,N_13653,N_13969);
xor U14160 (N_14160,N_13841,N_13666);
nor U14161 (N_14161,N_13738,N_13752);
nand U14162 (N_14162,N_13766,N_13878);
nor U14163 (N_14163,N_13850,N_13988);
nor U14164 (N_14164,N_13807,N_13831);
and U14165 (N_14165,N_13635,N_13948);
and U14166 (N_14166,N_13672,N_13986);
and U14167 (N_14167,N_13821,N_13605);
and U14168 (N_14168,N_13712,N_13847);
and U14169 (N_14169,N_13854,N_13829);
xor U14170 (N_14170,N_13695,N_13761);
xor U14171 (N_14171,N_13778,N_13996);
xnor U14172 (N_14172,N_13747,N_13833);
nor U14173 (N_14173,N_13977,N_13916);
xnor U14174 (N_14174,N_13758,N_13893);
nor U14175 (N_14175,N_13610,N_13694);
nand U14176 (N_14176,N_13890,N_13804);
nor U14177 (N_14177,N_13608,N_13720);
nor U14178 (N_14178,N_13716,N_13975);
xnor U14179 (N_14179,N_13609,N_13932);
or U14180 (N_14180,N_13637,N_13972);
or U14181 (N_14181,N_13884,N_13751);
nor U14182 (N_14182,N_13627,N_13843);
xor U14183 (N_14183,N_13641,N_13646);
xor U14184 (N_14184,N_13952,N_13675);
and U14185 (N_14185,N_13908,N_13906);
xnor U14186 (N_14186,N_13732,N_13983);
and U14187 (N_14187,N_13965,N_13775);
or U14188 (N_14188,N_13894,N_13700);
or U14189 (N_14189,N_13946,N_13754);
nor U14190 (N_14190,N_13881,N_13967);
or U14191 (N_14191,N_13816,N_13898);
xnor U14192 (N_14192,N_13671,N_13749);
nand U14193 (N_14193,N_13659,N_13974);
nand U14194 (N_14194,N_13708,N_13762);
xor U14195 (N_14195,N_13852,N_13702);
nand U14196 (N_14196,N_13950,N_13864);
and U14197 (N_14197,N_13741,N_13989);
xnor U14198 (N_14198,N_13883,N_13613);
and U14199 (N_14199,N_13985,N_13638);
nor U14200 (N_14200,N_13922,N_13825);
and U14201 (N_14201,N_13985,N_13853);
nor U14202 (N_14202,N_13833,N_13895);
or U14203 (N_14203,N_13945,N_13889);
nand U14204 (N_14204,N_13702,N_13770);
or U14205 (N_14205,N_13851,N_13942);
and U14206 (N_14206,N_13768,N_13871);
and U14207 (N_14207,N_13656,N_13613);
nor U14208 (N_14208,N_13768,N_13660);
nor U14209 (N_14209,N_13740,N_13679);
or U14210 (N_14210,N_13790,N_13795);
nand U14211 (N_14211,N_13803,N_13863);
nand U14212 (N_14212,N_13919,N_13667);
nor U14213 (N_14213,N_13881,N_13965);
and U14214 (N_14214,N_13865,N_13756);
or U14215 (N_14215,N_13742,N_13827);
nor U14216 (N_14216,N_13767,N_13667);
nor U14217 (N_14217,N_13743,N_13757);
nand U14218 (N_14218,N_13894,N_13617);
nand U14219 (N_14219,N_13672,N_13734);
nor U14220 (N_14220,N_13901,N_13929);
or U14221 (N_14221,N_13765,N_13807);
and U14222 (N_14222,N_13841,N_13723);
xor U14223 (N_14223,N_13828,N_13958);
and U14224 (N_14224,N_13658,N_13609);
nor U14225 (N_14225,N_13644,N_13807);
or U14226 (N_14226,N_13625,N_13669);
xor U14227 (N_14227,N_13614,N_13760);
nor U14228 (N_14228,N_13926,N_13870);
or U14229 (N_14229,N_13637,N_13849);
nor U14230 (N_14230,N_13655,N_13796);
xnor U14231 (N_14231,N_13799,N_13654);
nand U14232 (N_14232,N_13682,N_13633);
or U14233 (N_14233,N_13674,N_13705);
or U14234 (N_14234,N_13829,N_13749);
nand U14235 (N_14235,N_13960,N_13935);
or U14236 (N_14236,N_13896,N_13831);
or U14237 (N_14237,N_13711,N_13905);
nor U14238 (N_14238,N_13668,N_13732);
xor U14239 (N_14239,N_13901,N_13734);
nand U14240 (N_14240,N_13682,N_13999);
nor U14241 (N_14241,N_13630,N_13988);
xor U14242 (N_14242,N_13907,N_13921);
nand U14243 (N_14243,N_13708,N_13844);
xnor U14244 (N_14244,N_13694,N_13873);
nor U14245 (N_14245,N_13966,N_13878);
nor U14246 (N_14246,N_13809,N_13881);
or U14247 (N_14247,N_13798,N_13727);
nor U14248 (N_14248,N_13922,N_13731);
nand U14249 (N_14249,N_13878,N_13655);
xnor U14250 (N_14250,N_13645,N_13762);
nor U14251 (N_14251,N_13788,N_13696);
nor U14252 (N_14252,N_13942,N_13902);
nor U14253 (N_14253,N_13972,N_13913);
nand U14254 (N_14254,N_13947,N_13906);
nor U14255 (N_14255,N_13860,N_13918);
and U14256 (N_14256,N_13667,N_13886);
nor U14257 (N_14257,N_13984,N_13708);
nand U14258 (N_14258,N_13737,N_13809);
and U14259 (N_14259,N_13603,N_13947);
and U14260 (N_14260,N_13696,N_13979);
nand U14261 (N_14261,N_13793,N_13857);
nor U14262 (N_14262,N_13719,N_13746);
or U14263 (N_14263,N_13716,N_13884);
nor U14264 (N_14264,N_13997,N_13958);
nand U14265 (N_14265,N_13792,N_13864);
or U14266 (N_14266,N_13914,N_13994);
xnor U14267 (N_14267,N_13891,N_13882);
xnor U14268 (N_14268,N_13779,N_13938);
or U14269 (N_14269,N_13758,N_13838);
and U14270 (N_14270,N_13890,N_13668);
and U14271 (N_14271,N_13982,N_13854);
xor U14272 (N_14272,N_13986,N_13780);
or U14273 (N_14273,N_13801,N_13818);
nand U14274 (N_14274,N_13859,N_13842);
xor U14275 (N_14275,N_13641,N_13911);
or U14276 (N_14276,N_13882,N_13761);
and U14277 (N_14277,N_13726,N_13688);
or U14278 (N_14278,N_13867,N_13926);
nor U14279 (N_14279,N_13609,N_13629);
and U14280 (N_14280,N_13668,N_13674);
nand U14281 (N_14281,N_13769,N_13877);
nor U14282 (N_14282,N_13848,N_13639);
nor U14283 (N_14283,N_13669,N_13728);
or U14284 (N_14284,N_13638,N_13916);
xor U14285 (N_14285,N_13952,N_13961);
nor U14286 (N_14286,N_13673,N_13899);
xor U14287 (N_14287,N_13994,N_13835);
nor U14288 (N_14288,N_13781,N_13888);
nand U14289 (N_14289,N_13770,N_13996);
or U14290 (N_14290,N_13617,N_13897);
and U14291 (N_14291,N_13829,N_13619);
xnor U14292 (N_14292,N_13982,N_13632);
xor U14293 (N_14293,N_13751,N_13760);
and U14294 (N_14294,N_13986,N_13732);
nand U14295 (N_14295,N_13739,N_13923);
and U14296 (N_14296,N_13958,N_13784);
or U14297 (N_14297,N_13824,N_13946);
or U14298 (N_14298,N_13879,N_13603);
xor U14299 (N_14299,N_13923,N_13837);
and U14300 (N_14300,N_13711,N_13933);
and U14301 (N_14301,N_13954,N_13720);
or U14302 (N_14302,N_13603,N_13909);
and U14303 (N_14303,N_13966,N_13681);
or U14304 (N_14304,N_13700,N_13643);
or U14305 (N_14305,N_13853,N_13962);
and U14306 (N_14306,N_13672,N_13855);
nand U14307 (N_14307,N_13957,N_13776);
and U14308 (N_14308,N_13889,N_13991);
nor U14309 (N_14309,N_13704,N_13930);
xnor U14310 (N_14310,N_13978,N_13830);
and U14311 (N_14311,N_13732,N_13789);
and U14312 (N_14312,N_13623,N_13771);
xor U14313 (N_14313,N_13944,N_13966);
nor U14314 (N_14314,N_13862,N_13917);
nor U14315 (N_14315,N_13748,N_13620);
nand U14316 (N_14316,N_13937,N_13824);
nand U14317 (N_14317,N_13864,N_13992);
or U14318 (N_14318,N_13923,N_13878);
xnor U14319 (N_14319,N_13648,N_13841);
nand U14320 (N_14320,N_13666,N_13984);
and U14321 (N_14321,N_13994,N_13986);
nor U14322 (N_14322,N_13685,N_13784);
xor U14323 (N_14323,N_13630,N_13655);
nor U14324 (N_14324,N_13611,N_13928);
or U14325 (N_14325,N_13713,N_13734);
xor U14326 (N_14326,N_13733,N_13606);
xnor U14327 (N_14327,N_13878,N_13782);
xnor U14328 (N_14328,N_13715,N_13734);
nand U14329 (N_14329,N_13637,N_13802);
nand U14330 (N_14330,N_13844,N_13632);
nand U14331 (N_14331,N_13707,N_13910);
or U14332 (N_14332,N_13987,N_13741);
nor U14333 (N_14333,N_13855,N_13705);
xnor U14334 (N_14334,N_13914,N_13866);
and U14335 (N_14335,N_13600,N_13998);
and U14336 (N_14336,N_13792,N_13751);
and U14337 (N_14337,N_13692,N_13891);
xnor U14338 (N_14338,N_13922,N_13616);
and U14339 (N_14339,N_13756,N_13866);
and U14340 (N_14340,N_13930,N_13865);
and U14341 (N_14341,N_13634,N_13913);
and U14342 (N_14342,N_13959,N_13828);
and U14343 (N_14343,N_13756,N_13753);
nand U14344 (N_14344,N_13790,N_13614);
nor U14345 (N_14345,N_13841,N_13644);
or U14346 (N_14346,N_13670,N_13708);
nand U14347 (N_14347,N_13913,N_13777);
or U14348 (N_14348,N_13709,N_13955);
and U14349 (N_14349,N_13861,N_13697);
and U14350 (N_14350,N_13738,N_13948);
and U14351 (N_14351,N_13727,N_13623);
nand U14352 (N_14352,N_13705,N_13864);
nor U14353 (N_14353,N_13920,N_13803);
nand U14354 (N_14354,N_13848,N_13971);
nor U14355 (N_14355,N_13883,N_13950);
nor U14356 (N_14356,N_13610,N_13771);
or U14357 (N_14357,N_13956,N_13623);
and U14358 (N_14358,N_13994,N_13802);
nor U14359 (N_14359,N_13622,N_13905);
xor U14360 (N_14360,N_13975,N_13849);
nor U14361 (N_14361,N_13970,N_13843);
nor U14362 (N_14362,N_13673,N_13940);
or U14363 (N_14363,N_13688,N_13624);
or U14364 (N_14364,N_13818,N_13914);
xnor U14365 (N_14365,N_13617,N_13745);
and U14366 (N_14366,N_13875,N_13689);
and U14367 (N_14367,N_13732,N_13744);
nand U14368 (N_14368,N_13874,N_13633);
xor U14369 (N_14369,N_13762,N_13765);
nor U14370 (N_14370,N_13650,N_13721);
and U14371 (N_14371,N_13993,N_13820);
nand U14372 (N_14372,N_13923,N_13956);
and U14373 (N_14373,N_13865,N_13903);
nand U14374 (N_14374,N_13920,N_13804);
nor U14375 (N_14375,N_13899,N_13790);
nand U14376 (N_14376,N_13821,N_13797);
nand U14377 (N_14377,N_13996,N_13798);
and U14378 (N_14378,N_13823,N_13836);
and U14379 (N_14379,N_13827,N_13930);
nor U14380 (N_14380,N_13890,N_13664);
nor U14381 (N_14381,N_13854,N_13765);
nand U14382 (N_14382,N_13898,N_13682);
and U14383 (N_14383,N_13649,N_13823);
nand U14384 (N_14384,N_13791,N_13783);
xnor U14385 (N_14385,N_13605,N_13641);
nand U14386 (N_14386,N_13920,N_13887);
nor U14387 (N_14387,N_13772,N_13679);
and U14388 (N_14388,N_13762,N_13789);
or U14389 (N_14389,N_13723,N_13651);
nand U14390 (N_14390,N_13993,N_13718);
and U14391 (N_14391,N_13798,N_13987);
nor U14392 (N_14392,N_13873,N_13642);
and U14393 (N_14393,N_13935,N_13791);
nor U14394 (N_14394,N_13793,N_13691);
and U14395 (N_14395,N_13909,N_13766);
or U14396 (N_14396,N_13799,N_13935);
xnor U14397 (N_14397,N_13822,N_13716);
nor U14398 (N_14398,N_13670,N_13698);
nor U14399 (N_14399,N_13837,N_13944);
nand U14400 (N_14400,N_14094,N_14111);
or U14401 (N_14401,N_14205,N_14272);
or U14402 (N_14402,N_14026,N_14052);
xnor U14403 (N_14403,N_14070,N_14048);
or U14404 (N_14404,N_14043,N_14073);
nor U14405 (N_14405,N_14268,N_14109);
xnor U14406 (N_14406,N_14286,N_14361);
or U14407 (N_14407,N_14099,N_14334);
or U14408 (N_14408,N_14128,N_14105);
xnor U14409 (N_14409,N_14343,N_14092);
nand U14410 (N_14410,N_14011,N_14381);
or U14411 (N_14411,N_14395,N_14248);
xor U14412 (N_14412,N_14037,N_14013);
or U14413 (N_14413,N_14106,N_14084);
xnor U14414 (N_14414,N_14143,N_14309);
xnor U14415 (N_14415,N_14147,N_14333);
xnor U14416 (N_14416,N_14172,N_14022);
and U14417 (N_14417,N_14337,N_14151);
and U14418 (N_14418,N_14354,N_14207);
nand U14419 (N_14419,N_14368,N_14330);
nand U14420 (N_14420,N_14158,N_14173);
or U14421 (N_14421,N_14038,N_14371);
nand U14422 (N_14422,N_14169,N_14217);
nand U14423 (N_14423,N_14317,N_14004);
xor U14424 (N_14424,N_14076,N_14254);
nor U14425 (N_14425,N_14163,N_14285);
xnor U14426 (N_14426,N_14398,N_14122);
and U14427 (N_14427,N_14136,N_14377);
and U14428 (N_14428,N_14039,N_14003);
and U14429 (N_14429,N_14213,N_14081);
nand U14430 (N_14430,N_14063,N_14025);
and U14431 (N_14431,N_14168,N_14164);
nor U14432 (N_14432,N_14196,N_14127);
and U14433 (N_14433,N_14090,N_14244);
nor U14434 (N_14434,N_14262,N_14259);
and U14435 (N_14435,N_14057,N_14282);
nor U14436 (N_14436,N_14385,N_14249);
and U14437 (N_14437,N_14329,N_14382);
or U14438 (N_14438,N_14197,N_14340);
and U14439 (N_14439,N_14047,N_14346);
or U14440 (N_14440,N_14100,N_14365);
nor U14441 (N_14441,N_14328,N_14363);
and U14442 (N_14442,N_14206,N_14288);
xor U14443 (N_14443,N_14142,N_14133);
nand U14444 (N_14444,N_14120,N_14351);
nor U14445 (N_14445,N_14021,N_14201);
or U14446 (N_14446,N_14251,N_14059);
nor U14447 (N_14447,N_14289,N_14186);
and U14448 (N_14448,N_14373,N_14116);
and U14449 (N_14449,N_14091,N_14293);
nand U14450 (N_14450,N_14269,N_14126);
nor U14451 (N_14451,N_14235,N_14036);
and U14452 (N_14452,N_14029,N_14016);
nand U14453 (N_14453,N_14228,N_14352);
xor U14454 (N_14454,N_14291,N_14345);
xnor U14455 (N_14455,N_14212,N_14239);
or U14456 (N_14456,N_14087,N_14290);
or U14457 (N_14457,N_14135,N_14321);
xnor U14458 (N_14458,N_14181,N_14040);
nand U14459 (N_14459,N_14086,N_14359);
or U14460 (N_14460,N_14224,N_14166);
or U14461 (N_14461,N_14104,N_14215);
and U14462 (N_14462,N_14306,N_14374);
and U14463 (N_14463,N_14129,N_14171);
xor U14464 (N_14464,N_14218,N_14332);
xor U14465 (N_14465,N_14298,N_14231);
and U14466 (N_14466,N_14350,N_14032);
or U14467 (N_14467,N_14358,N_14055);
nand U14468 (N_14468,N_14221,N_14149);
nor U14469 (N_14469,N_14012,N_14256);
nor U14470 (N_14470,N_14216,N_14017);
and U14471 (N_14471,N_14214,N_14344);
xor U14472 (N_14472,N_14349,N_14211);
nor U14473 (N_14473,N_14240,N_14305);
xnor U14474 (N_14474,N_14390,N_14277);
or U14475 (N_14475,N_14190,N_14050);
nand U14476 (N_14476,N_14378,N_14131);
nor U14477 (N_14477,N_14083,N_14252);
or U14478 (N_14478,N_14322,N_14372);
and U14479 (N_14479,N_14366,N_14179);
nor U14480 (N_14480,N_14155,N_14316);
nor U14481 (N_14481,N_14257,N_14042);
nor U14482 (N_14482,N_14139,N_14118);
and U14483 (N_14483,N_14014,N_14130);
or U14484 (N_14484,N_14000,N_14194);
or U14485 (N_14485,N_14331,N_14255);
nor U14486 (N_14486,N_14008,N_14234);
nor U14487 (N_14487,N_14353,N_14189);
nand U14488 (N_14488,N_14261,N_14360);
xor U14489 (N_14489,N_14188,N_14125);
nor U14490 (N_14490,N_14225,N_14170);
xor U14491 (N_14491,N_14198,N_14101);
or U14492 (N_14492,N_14061,N_14020);
xor U14493 (N_14493,N_14204,N_14112);
xnor U14494 (N_14494,N_14064,N_14369);
nand U14495 (N_14495,N_14080,N_14270);
or U14496 (N_14496,N_14077,N_14274);
or U14497 (N_14497,N_14035,N_14028);
xnor U14498 (N_14498,N_14362,N_14200);
nand U14499 (N_14499,N_14024,N_14276);
nand U14500 (N_14500,N_14380,N_14030);
xor U14501 (N_14501,N_14138,N_14060);
nand U14502 (N_14502,N_14193,N_14156);
nand U14503 (N_14503,N_14237,N_14150);
and U14504 (N_14504,N_14312,N_14154);
xor U14505 (N_14505,N_14236,N_14279);
nor U14506 (N_14506,N_14260,N_14295);
nor U14507 (N_14507,N_14278,N_14089);
nor U14508 (N_14508,N_14157,N_14242);
nand U14509 (N_14509,N_14247,N_14132);
nor U14510 (N_14510,N_14069,N_14210);
or U14511 (N_14511,N_14273,N_14165);
and U14512 (N_14512,N_14324,N_14275);
or U14513 (N_14513,N_14308,N_14019);
xor U14514 (N_14514,N_14370,N_14307);
and U14515 (N_14515,N_14284,N_14113);
or U14516 (N_14516,N_14051,N_14005);
or U14517 (N_14517,N_14176,N_14271);
nor U14518 (N_14518,N_14015,N_14348);
nand U14519 (N_14519,N_14185,N_14357);
and U14520 (N_14520,N_14287,N_14031);
and U14521 (N_14521,N_14065,N_14085);
or U14522 (N_14522,N_14199,N_14192);
xor U14523 (N_14523,N_14148,N_14174);
and U14524 (N_14524,N_14023,N_14222);
nand U14525 (N_14525,N_14356,N_14182);
or U14526 (N_14526,N_14137,N_14297);
or U14527 (N_14527,N_14079,N_14146);
nor U14528 (N_14528,N_14396,N_14161);
nand U14529 (N_14529,N_14068,N_14313);
or U14530 (N_14530,N_14115,N_14376);
or U14531 (N_14531,N_14209,N_14009);
or U14532 (N_14532,N_14379,N_14219);
and U14533 (N_14533,N_14203,N_14062);
nand U14534 (N_14534,N_14058,N_14347);
or U14535 (N_14535,N_14241,N_14338);
xor U14536 (N_14536,N_14310,N_14007);
xor U14537 (N_14537,N_14053,N_14243);
and U14538 (N_14538,N_14299,N_14074);
nor U14539 (N_14539,N_14049,N_14121);
and U14540 (N_14540,N_14153,N_14180);
nor U14541 (N_14541,N_14386,N_14093);
and U14542 (N_14542,N_14342,N_14223);
and U14543 (N_14543,N_14304,N_14323);
and U14544 (N_14544,N_14245,N_14364);
nor U14545 (N_14545,N_14082,N_14018);
nor U14546 (N_14546,N_14162,N_14265);
nand U14547 (N_14547,N_14187,N_14391);
xor U14548 (N_14548,N_14384,N_14191);
and U14549 (N_14549,N_14263,N_14072);
and U14550 (N_14550,N_14341,N_14140);
and U14551 (N_14551,N_14102,N_14302);
or U14552 (N_14552,N_14208,N_14296);
and U14553 (N_14553,N_14399,N_14114);
nand U14554 (N_14554,N_14281,N_14107);
or U14555 (N_14555,N_14066,N_14110);
nand U14556 (N_14556,N_14144,N_14202);
xor U14557 (N_14557,N_14318,N_14336);
nand U14558 (N_14558,N_14388,N_14253);
nor U14559 (N_14559,N_14145,N_14183);
nand U14560 (N_14560,N_14033,N_14119);
or U14561 (N_14561,N_14264,N_14394);
and U14562 (N_14562,N_14292,N_14266);
nand U14563 (N_14563,N_14159,N_14027);
and U14564 (N_14564,N_14258,N_14319);
nand U14565 (N_14565,N_14001,N_14071);
nor U14566 (N_14566,N_14283,N_14046);
nand U14567 (N_14567,N_14355,N_14177);
xor U14568 (N_14568,N_14280,N_14389);
xor U14569 (N_14569,N_14045,N_14088);
and U14570 (N_14570,N_14375,N_14117);
nor U14571 (N_14571,N_14034,N_14230);
nand U14572 (N_14572,N_14175,N_14220);
and U14573 (N_14573,N_14238,N_14320);
xor U14574 (N_14574,N_14335,N_14097);
nor U14575 (N_14575,N_14054,N_14041);
nand U14576 (N_14576,N_14267,N_14103);
nor U14577 (N_14577,N_14315,N_14250);
and U14578 (N_14578,N_14096,N_14056);
nor U14579 (N_14579,N_14367,N_14108);
xor U14580 (N_14580,N_14006,N_14294);
or U14581 (N_14581,N_14160,N_14327);
or U14582 (N_14582,N_14393,N_14383);
and U14583 (N_14583,N_14226,N_14078);
xor U14584 (N_14584,N_14303,N_14232);
and U14585 (N_14585,N_14184,N_14195);
nand U14586 (N_14586,N_14326,N_14325);
nor U14587 (N_14587,N_14233,N_14387);
xor U14588 (N_14588,N_14010,N_14123);
xor U14589 (N_14589,N_14152,N_14314);
or U14590 (N_14590,N_14301,N_14124);
xnor U14591 (N_14591,N_14229,N_14095);
or U14592 (N_14592,N_14300,N_14098);
and U14593 (N_14593,N_14141,N_14067);
xnor U14594 (N_14594,N_14002,N_14246);
or U14595 (N_14595,N_14167,N_14134);
and U14596 (N_14596,N_14178,N_14397);
and U14597 (N_14597,N_14392,N_14075);
nor U14598 (N_14598,N_14227,N_14044);
nand U14599 (N_14599,N_14311,N_14339);
and U14600 (N_14600,N_14139,N_14302);
xor U14601 (N_14601,N_14002,N_14130);
or U14602 (N_14602,N_14229,N_14266);
or U14603 (N_14603,N_14367,N_14122);
nand U14604 (N_14604,N_14267,N_14391);
or U14605 (N_14605,N_14110,N_14219);
nand U14606 (N_14606,N_14356,N_14390);
xnor U14607 (N_14607,N_14098,N_14009);
nor U14608 (N_14608,N_14288,N_14289);
xnor U14609 (N_14609,N_14398,N_14204);
nor U14610 (N_14610,N_14101,N_14020);
nand U14611 (N_14611,N_14081,N_14289);
nor U14612 (N_14612,N_14129,N_14221);
xor U14613 (N_14613,N_14121,N_14024);
nand U14614 (N_14614,N_14315,N_14004);
xnor U14615 (N_14615,N_14015,N_14318);
or U14616 (N_14616,N_14281,N_14238);
xor U14617 (N_14617,N_14273,N_14212);
nor U14618 (N_14618,N_14052,N_14005);
nor U14619 (N_14619,N_14103,N_14348);
nand U14620 (N_14620,N_14332,N_14281);
and U14621 (N_14621,N_14355,N_14009);
xor U14622 (N_14622,N_14323,N_14226);
or U14623 (N_14623,N_14036,N_14030);
and U14624 (N_14624,N_14166,N_14085);
nand U14625 (N_14625,N_14165,N_14128);
nor U14626 (N_14626,N_14107,N_14292);
or U14627 (N_14627,N_14295,N_14269);
xor U14628 (N_14628,N_14184,N_14030);
nand U14629 (N_14629,N_14260,N_14240);
nand U14630 (N_14630,N_14005,N_14281);
nor U14631 (N_14631,N_14388,N_14002);
nand U14632 (N_14632,N_14294,N_14295);
xor U14633 (N_14633,N_14065,N_14206);
and U14634 (N_14634,N_14375,N_14188);
nand U14635 (N_14635,N_14378,N_14087);
xnor U14636 (N_14636,N_14364,N_14247);
and U14637 (N_14637,N_14070,N_14006);
nand U14638 (N_14638,N_14265,N_14100);
or U14639 (N_14639,N_14323,N_14105);
and U14640 (N_14640,N_14016,N_14206);
or U14641 (N_14641,N_14104,N_14048);
and U14642 (N_14642,N_14157,N_14360);
and U14643 (N_14643,N_14301,N_14063);
or U14644 (N_14644,N_14383,N_14257);
or U14645 (N_14645,N_14073,N_14028);
or U14646 (N_14646,N_14104,N_14067);
nand U14647 (N_14647,N_14399,N_14341);
nand U14648 (N_14648,N_14354,N_14318);
or U14649 (N_14649,N_14273,N_14113);
or U14650 (N_14650,N_14053,N_14075);
and U14651 (N_14651,N_14083,N_14008);
nor U14652 (N_14652,N_14279,N_14068);
nand U14653 (N_14653,N_14145,N_14196);
xor U14654 (N_14654,N_14296,N_14128);
or U14655 (N_14655,N_14290,N_14360);
nand U14656 (N_14656,N_14071,N_14198);
and U14657 (N_14657,N_14022,N_14227);
nand U14658 (N_14658,N_14141,N_14264);
nand U14659 (N_14659,N_14130,N_14108);
nor U14660 (N_14660,N_14029,N_14187);
nor U14661 (N_14661,N_14024,N_14058);
xnor U14662 (N_14662,N_14260,N_14355);
or U14663 (N_14663,N_14050,N_14241);
xor U14664 (N_14664,N_14197,N_14328);
xnor U14665 (N_14665,N_14007,N_14179);
nand U14666 (N_14666,N_14102,N_14390);
and U14667 (N_14667,N_14159,N_14060);
nor U14668 (N_14668,N_14349,N_14141);
and U14669 (N_14669,N_14051,N_14095);
or U14670 (N_14670,N_14235,N_14292);
nor U14671 (N_14671,N_14184,N_14319);
and U14672 (N_14672,N_14075,N_14046);
nor U14673 (N_14673,N_14239,N_14233);
xor U14674 (N_14674,N_14086,N_14207);
and U14675 (N_14675,N_14056,N_14218);
nor U14676 (N_14676,N_14242,N_14353);
xor U14677 (N_14677,N_14031,N_14008);
or U14678 (N_14678,N_14082,N_14028);
nor U14679 (N_14679,N_14236,N_14369);
or U14680 (N_14680,N_14134,N_14053);
and U14681 (N_14681,N_14264,N_14361);
xnor U14682 (N_14682,N_14354,N_14037);
nand U14683 (N_14683,N_14147,N_14384);
and U14684 (N_14684,N_14076,N_14109);
nor U14685 (N_14685,N_14002,N_14294);
nand U14686 (N_14686,N_14298,N_14058);
or U14687 (N_14687,N_14370,N_14131);
nand U14688 (N_14688,N_14076,N_14206);
and U14689 (N_14689,N_14020,N_14181);
nor U14690 (N_14690,N_14200,N_14186);
and U14691 (N_14691,N_14171,N_14219);
and U14692 (N_14692,N_14149,N_14390);
nand U14693 (N_14693,N_14126,N_14130);
xor U14694 (N_14694,N_14374,N_14090);
and U14695 (N_14695,N_14237,N_14238);
xnor U14696 (N_14696,N_14027,N_14145);
nand U14697 (N_14697,N_14080,N_14323);
xor U14698 (N_14698,N_14074,N_14081);
or U14699 (N_14699,N_14066,N_14086);
and U14700 (N_14700,N_14099,N_14386);
xnor U14701 (N_14701,N_14024,N_14348);
nor U14702 (N_14702,N_14028,N_14110);
or U14703 (N_14703,N_14027,N_14304);
xor U14704 (N_14704,N_14302,N_14369);
nor U14705 (N_14705,N_14115,N_14388);
nor U14706 (N_14706,N_14029,N_14353);
nand U14707 (N_14707,N_14068,N_14228);
or U14708 (N_14708,N_14144,N_14317);
xor U14709 (N_14709,N_14035,N_14327);
nor U14710 (N_14710,N_14168,N_14373);
or U14711 (N_14711,N_14239,N_14330);
nor U14712 (N_14712,N_14224,N_14376);
or U14713 (N_14713,N_14197,N_14205);
or U14714 (N_14714,N_14150,N_14257);
xor U14715 (N_14715,N_14378,N_14370);
or U14716 (N_14716,N_14348,N_14177);
nor U14717 (N_14717,N_14118,N_14067);
nand U14718 (N_14718,N_14213,N_14338);
and U14719 (N_14719,N_14101,N_14008);
and U14720 (N_14720,N_14111,N_14157);
nand U14721 (N_14721,N_14250,N_14296);
nor U14722 (N_14722,N_14111,N_14381);
or U14723 (N_14723,N_14128,N_14184);
nand U14724 (N_14724,N_14368,N_14191);
xor U14725 (N_14725,N_14237,N_14083);
xor U14726 (N_14726,N_14131,N_14148);
and U14727 (N_14727,N_14214,N_14270);
and U14728 (N_14728,N_14276,N_14085);
xor U14729 (N_14729,N_14142,N_14168);
and U14730 (N_14730,N_14129,N_14306);
and U14731 (N_14731,N_14052,N_14269);
and U14732 (N_14732,N_14179,N_14247);
and U14733 (N_14733,N_14394,N_14386);
or U14734 (N_14734,N_14117,N_14185);
and U14735 (N_14735,N_14176,N_14161);
nor U14736 (N_14736,N_14290,N_14342);
nand U14737 (N_14737,N_14270,N_14238);
xor U14738 (N_14738,N_14177,N_14253);
nand U14739 (N_14739,N_14140,N_14382);
and U14740 (N_14740,N_14098,N_14309);
or U14741 (N_14741,N_14162,N_14201);
nor U14742 (N_14742,N_14134,N_14119);
or U14743 (N_14743,N_14023,N_14057);
or U14744 (N_14744,N_14120,N_14070);
nor U14745 (N_14745,N_14270,N_14188);
xnor U14746 (N_14746,N_14115,N_14162);
nor U14747 (N_14747,N_14183,N_14205);
nor U14748 (N_14748,N_14121,N_14068);
xor U14749 (N_14749,N_14149,N_14173);
and U14750 (N_14750,N_14271,N_14340);
nand U14751 (N_14751,N_14002,N_14029);
or U14752 (N_14752,N_14355,N_14052);
xnor U14753 (N_14753,N_14399,N_14298);
and U14754 (N_14754,N_14344,N_14250);
and U14755 (N_14755,N_14129,N_14271);
and U14756 (N_14756,N_14061,N_14048);
nand U14757 (N_14757,N_14311,N_14010);
xnor U14758 (N_14758,N_14160,N_14185);
nand U14759 (N_14759,N_14296,N_14314);
nor U14760 (N_14760,N_14108,N_14052);
xnor U14761 (N_14761,N_14225,N_14085);
xnor U14762 (N_14762,N_14141,N_14008);
xnor U14763 (N_14763,N_14206,N_14382);
or U14764 (N_14764,N_14008,N_14231);
nor U14765 (N_14765,N_14146,N_14388);
and U14766 (N_14766,N_14268,N_14216);
xor U14767 (N_14767,N_14028,N_14264);
xor U14768 (N_14768,N_14120,N_14205);
xor U14769 (N_14769,N_14014,N_14140);
or U14770 (N_14770,N_14114,N_14276);
nand U14771 (N_14771,N_14227,N_14023);
and U14772 (N_14772,N_14096,N_14361);
xor U14773 (N_14773,N_14374,N_14219);
nor U14774 (N_14774,N_14198,N_14268);
and U14775 (N_14775,N_14264,N_14113);
nand U14776 (N_14776,N_14146,N_14298);
xnor U14777 (N_14777,N_14323,N_14111);
nand U14778 (N_14778,N_14282,N_14044);
and U14779 (N_14779,N_14079,N_14160);
or U14780 (N_14780,N_14147,N_14068);
or U14781 (N_14781,N_14384,N_14231);
nor U14782 (N_14782,N_14389,N_14047);
or U14783 (N_14783,N_14220,N_14006);
xor U14784 (N_14784,N_14077,N_14048);
and U14785 (N_14785,N_14157,N_14231);
or U14786 (N_14786,N_14394,N_14320);
nor U14787 (N_14787,N_14241,N_14270);
and U14788 (N_14788,N_14057,N_14140);
or U14789 (N_14789,N_14010,N_14006);
nor U14790 (N_14790,N_14341,N_14222);
xor U14791 (N_14791,N_14048,N_14188);
and U14792 (N_14792,N_14080,N_14299);
nand U14793 (N_14793,N_14316,N_14343);
xor U14794 (N_14794,N_14141,N_14217);
or U14795 (N_14795,N_14016,N_14266);
nor U14796 (N_14796,N_14096,N_14283);
xnor U14797 (N_14797,N_14226,N_14202);
nor U14798 (N_14798,N_14215,N_14154);
and U14799 (N_14799,N_14118,N_14095);
or U14800 (N_14800,N_14439,N_14520);
and U14801 (N_14801,N_14681,N_14786);
nand U14802 (N_14802,N_14459,N_14753);
nand U14803 (N_14803,N_14757,N_14725);
and U14804 (N_14804,N_14524,N_14656);
xnor U14805 (N_14805,N_14470,N_14473);
or U14806 (N_14806,N_14515,N_14564);
nor U14807 (N_14807,N_14488,N_14677);
nand U14808 (N_14808,N_14538,N_14478);
and U14809 (N_14809,N_14685,N_14576);
and U14810 (N_14810,N_14581,N_14794);
and U14811 (N_14811,N_14512,N_14412);
or U14812 (N_14812,N_14674,N_14710);
nand U14813 (N_14813,N_14768,N_14694);
xnor U14814 (N_14814,N_14454,N_14463);
nand U14815 (N_14815,N_14718,N_14483);
or U14816 (N_14816,N_14551,N_14643);
nor U14817 (N_14817,N_14622,N_14735);
xor U14818 (N_14818,N_14763,N_14627);
and U14819 (N_14819,N_14462,N_14783);
nor U14820 (N_14820,N_14562,N_14746);
xnor U14821 (N_14821,N_14587,N_14471);
nand U14822 (N_14822,N_14691,N_14772);
and U14823 (N_14823,N_14670,N_14719);
xnor U14824 (N_14824,N_14577,N_14608);
xor U14825 (N_14825,N_14417,N_14420);
and U14826 (N_14826,N_14578,N_14616);
or U14827 (N_14827,N_14623,N_14546);
xor U14828 (N_14828,N_14762,N_14765);
xor U14829 (N_14829,N_14791,N_14407);
or U14830 (N_14830,N_14662,N_14713);
nor U14831 (N_14831,N_14416,N_14641);
nand U14832 (N_14832,N_14590,N_14442);
nand U14833 (N_14833,N_14517,N_14777);
nor U14834 (N_14834,N_14775,N_14502);
or U14835 (N_14835,N_14599,N_14796);
nor U14836 (N_14836,N_14610,N_14501);
nand U14837 (N_14837,N_14704,N_14575);
nand U14838 (N_14838,N_14741,N_14711);
nor U14839 (N_14839,N_14460,N_14728);
and U14840 (N_14840,N_14537,N_14607);
nor U14841 (N_14841,N_14702,N_14489);
or U14842 (N_14842,N_14661,N_14697);
nand U14843 (N_14843,N_14550,N_14591);
nand U14844 (N_14844,N_14464,N_14522);
nor U14845 (N_14845,N_14596,N_14586);
or U14846 (N_14846,N_14499,N_14434);
xor U14847 (N_14847,N_14518,N_14679);
or U14848 (N_14848,N_14759,N_14745);
nand U14849 (N_14849,N_14769,N_14453);
and U14850 (N_14850,N_14655,N_14490);
or U14851 (N_14851,N_14668,N_14427);
nor U14852 (N_14852,N_14480,N_14498);
xnor U14853 (N_14853,N_14531,N_14560);
and U14854 (N_14854,N_14521,N_14536);
nand U14855 (N_14855,N_14738,N_14653);
xnor U14856 (N_14856,N_14636,N_14799);
nand U14857 (N_14857,N_14771,N_14760);
or U14858 (N_14858,N_14722,N_14472);
xor U14859 (N_14859,N_14751,N_14740);
nand U14860 (N_14860,N_14559,N_14708);
nor U14861 (N_14861,N_14781,N_14443);
nor U14862 (N_14862,N_14785,N_14500);
nand U14863 (N_14863,N_14479,N_14692);
and U14864 (N_14864,N_14743,N_14620);
nand U14865 (N_14865,N_14495,N_14458);
xnor U14866 (N_14866,N_14665,N_14695);
or U14867 (N_14867,N_14650,N_14657);
or U14868 (N_14868,N_14709,N_14510);
nor U14869 (N_14869,N_14592,N_14432);
and U14870 (N_14870,N_14739,N_14647);
nor U14871 (N_14871,N_14450,N_14602);
or U14872 (N_14872,N_14658,N_14606);
nor U14873 (N_14873,N_14487,N_14541);
nand U14874 (N_14874,N_14631,N_14526);
and U14875 (N_14875,N_14406,N_14570);
nand U14876 (N_14876,N_14424,N_14484);
xor U14877 (N_14877,N_14642,N_14689);
nor U14878 (N_14878,N_14737,N_14507);
nor U14879 (N_14879,N_14418,N_14566);
or U14880 (N_14880,N_14744,N_14544);
xor U14881 (N_14881,N_14761,N_14782);
xnor U14882 (N_14882,N_14696,N_14752);
xor U14883 (N_14883,N_14402,N_14456);
xnor U14884 (N_14884,N_14428,N_14633);
and U14885 (N_14885,N_14667,N_14605);
and U14886 (N_14886,N_14475,N_14648);
and U14887 (N_14887,N_14435,N_14686);
and U14888 (N_14888,N_14523,N_14496);
xor U14889 (N_14889,N_14569,N_14707);
or U14890 (N_14890,N_14654,N_14530);
and U14891 (N_14891,N_14614,N_14580);
and U14892 (N_14892,N_14469,N_14758);
xor U14893 (N_14893,N_14629,N_14535);
nor U14894 (N_14894,N_14584,N_14419);
xnor U14895 (N_14895,N_14409,N_14784);
or U14896 (N_14896,N_14663,N_14609);
and U14897 (N_14897,N_14764,N_14554);
xnor U14898 (N_14898,N_14730,N_14637);
nand U14899 (N_14899,N_14403,N_14563);
nor U14900 (N_14900,N_14508,N_14736);
and U14901 (N_14901,N_14579,N_14548);
or U14902 (N_14902,N_14749,N_14766);
xnor U14903 (N_14903,N_14513,N_14553);
nor U14904 (N_14904,N_14733,N_14767);
xor U14905 (N_14905,N_14613,N_14687);
xnor U14906 (N_14906,N_14747,N_14603);
or U14907 (N_14907,N_14600,N_14542);
nor U14908 (N_14908,N_14493,N_14754);
nor U14909 (N_14909,N_14703,N_14717);
and U14910 (N_14910,N_14669,N_14798);
and U14911 (N_14911,N_14452,N_14425);
nand U14912 (N_14912,N_14774,N_14660);
and U14913 (N_14913,N_14568,N_14492);
or U14914 (N_14914,N_14481,N_14755);
or U14915 (N_14915,N_14482,N_14683);
xnor U14916 (N_14916,N_14436,N_14748);
xor U14917 (N_14917,N_14601,N_14638);
nor U14918 (N_14918,N_14404,N_14441);
nor U14919 (N_14919,N_14506,N_14431);
xor U14920 (N_14920,N_14534,N_14491);
or U14921 (N_14921,N_14540,N_14672);
xnor U14922 (N_14922,N_14705,N_14438);
nor U14923 (N_14923,N_14617,N_14720);
or U14924 (N_14924,N_14726,N_14429);
xor U14925 (N_14925,N_14449,N_14455);
xor U14926 (N_14926,N_14573,N_14445);
or U14927 (N_14927,N_14497,N_14448);
nand U14928 (N_14928,N_14645,N_14780);
xnor U14929 (N_14929,N_14706,N_14734);
nand U14930 (N_14930,N_14572,N_14693);
or U14931 (N_14931,N_14666,N_14649);
or U14932 (N_14932,N_14451,N_14582);
nand U14933 (N_14933,N_14466,N_14675);
or U14934 (N_14934,N_14618,N_14626);
xnor U14935 (N_14935,N_14476,N_14595);
xnor U14936 (N_14936,N_14457,N_14678);
or U14937 (N_14937,N_14589,N_14615);
or U14938 (N_14938,N_14516,N_14400);
and U14939 (N_14939,N_14630,N_14509);
nor U14940 (N_14940,N_14405,N_14684);
nor U14941 (N_14941,N_14659,N_14423);
xor U14942 (N_14942,N_14477,N_14494);
nor U14943 (N_14943,N_14598,N_14621);
nand U14944 (N_14944,N_14715,N_14408);
nor U14945 (N_14945,N_14539,N_14440);
and U14946 (N_14946,N_14742,N_14532);
xor U14947 (N_14947,N_14511,N_14700);
nor U14948 (N_14948,N_14635,N_14619);
nand U14949 (N_14949,N_14699,N_14597);
nand U14950 (N_14950,N_14652,N_14413);
and U14951 (N_14951,N_14411,N_14433);
or U14952 (N_14952,N_14634,N_14611);
or U14953 (N_14953,N_14690,N_14793);
nor U14954 (N_14954,N_14547,N_14716);
nor U14955 (N_14955,N_14529,N_14625);
and U14956 (N_14956,N_14426,N_14731);
and U14957 (N_14957,N_14525,N_14410);
and U14958 (N_14958,N_14474,N_14787);
nand U14959 (N_14959,N_14555,N_14486);
xor U14960 (N_14960,N_14698,N_14792);
or U14961 (N_14961,N_14504,N_14519);
nand U14962 (N_14962,N_14797,N_14721);
xnor U14963 (N_14963,N_14505,N_14795);
or U14964 (N_14964,N_14401,N_14447);
and U14965 (N_14965,N_14682,N_14640);
or U14966 (N_14966,N_14461,N_14646);
nand U14967 (N_14967,N_14528,N_14485);
or U14968 (N_14968,N_14770,N_14514);
xor U14969 (N_14969,N_14556,N_14664);
xor U14970 (N_14970,N_14571,N_14465);
xnor U14971 (N_14971,N_14415,N_14789);
nor U14972 (N_14972,N_14727,N_14468);
or U14973 (N_14973,N_14594,N_14624);
xor U14974 (N_14974,N_14714,N_14676);
xnor U14975 (N_14975,N_14724,N_14779);
and U14976 (N_14976,N_14756,N_14437);
nor U14977 (N_14977,N_14444,N_14680);
nand U14978 (N_14978,N_14776,N_14567);
and U14979 (N_14979,N_14773,N_14604);
and U14980 (N_14980,N_14612,N_14723);
nor U14981 (N_14981,N_14588,N_14430);
or U14982 (N_14982,N_14673,N_14585);
xnor U14983 (N_14983,N_14545,N_14750);
or U14984 (N_14984,N_14788,N_14549);
xor U14985 (N_14985,N_14790,N_14778);
xnor U14986 (N_14986,N_14651,N_14527);
xor U14987 (N_14987,N_14552,N_14712);
nand U14988 (N_14988,N_14565,N_14543);
nand U14989 (N_14989,N_14628,N_14729);
nand U14990 (N_14990,N_14558,N_14671);
nand U14991 (N_14991,N_14503,N_14632);
or U14992 (N_14992,N_14732,N_14574);
nand U14993 (N_14993,N_14557,N_14421);
and U14994 (N_14994,N_14583,N_14467);
xor U14995 (N_14995,N_14422,N_14533);
nand U14996 (N_14996,N_14446,N_14561);
nor U14997 (N_14997,N_14639,N_14593);
or U14998 (N_14998,N_14701,N_14688);
nand U14999 (N_14999,N_14644,N_14414);
or U15000 (N_15000,N_14764,N_14522);
nor U15001 (N_15001,N_14464,N_14761);
xnor U15002 (N_15002,N_14795,N_14725);
nor U15003 (N_15003,N_14519,N_14791);
nand U15004 (N_15004,N_14543,N_14698);
nor U15005 (N_15005,N_14737,N_14746);
nand U15006 (N_15006,N_14645,N_14626);
or U15007 (N_15007,N_14406,N_14785);
xor U15008 (N_15008,N_14792,N_14720);
nor U15009 (N_15009,N_14622,N_14508);
and U15010 (N_15010,N_14638,N_14795);
nand U15011 (N_15011,N_14675,N_14728);
or U15012 (N_15012,N_14742,N_14466);
nor U15013 (N_15013,N_14694,N_14595);
or U15014 (N_15014,N_14713,N_14781);
and U15015 (N_15015,N_14673,N_14421);
or U15016 (N_15016,N_14683,N_14695);
nor U15017 (N_15017,N_14477,N_14577);
nand U15018 (N_15018,N_14482,N_14511);
or U15019 (N_15019,N_14784,N_14422);
nor U15020 (N_15020,N_14539,N_14558);
nand U15021 (N_15021,N_14605,N_14563);
nand U15022 (N_15022,N_14731,N_14719);
and U15023 (N_15023,N_14571,N_14569);
or U15024 (N_15024,N_14688,N_14541);
and U15025 (N_15025,N_14565,N_14522);
or U15026 (N_15026,N_14461,N_14651);
nor U15027 (N_15027,N_14642,N_14785);
nand U15028 (N_15028,N_14635,N_14641);
xor U15029 (N_15029,N_14719,N_14785);
and U15030 (N_15030,N_14592,N_14688);
nand U15031 (N_15031,N_14553,N_14767);
nor U15032 (N_15032,N_14651,N_14564);
or U15033 (N_15033,N_14434,N_14705);
or U15034 (N_15034,N_14506,N_14791);
nor U15035 (N_15035,N_14772,N_14790);
nor U15036 (N_15036,N_14453,N_14549);
xor U15037 (N_15037,N_14515,N_14421);
nand U15038 (N_15038,N_14423,N_14613);
and U15039 (N_15039,N_14475,N_14706);
or U15040 (N_15040,N_14608,N_14443);
xor U15041 (N_15041,N_14480,N_14579);
and U15042 (N_15042,N_14739,N_14620);
and U15043 (N_15043,N_14433,N_14783);
and U15044 (N_15044,N_14498,N_14430);
xor U15045 (N_15045,N_14651,N_14628);
xnor U15046 (N_15046,N_14684,N_14482);
or U15047 (N_15047,N_14721,N_14628);
and U15048 (N_15048,N_14623,N_14423);
and U15049 (N_15049,N_14476,N_14673);
xor U15050 (N_15050,N_14480,N_14587);
xnor U15051 (N_15051,N_14634,N_14669);
xnor U15052 (N_15052,N_14794,N_14683);
or U15053 (N_15053,N_14412,N_14571);
or U15054 (N_15054,N_14768,N_14654);
xor U15055 (N_15055,N_14659,N_14627);
nand U15056 (N_15056,N_14582,N_14721);
and U15057 (N_15057,N_14423,N_14528);
xor U15058 (N_15058,N_14523,N_14770);
or U15059 (N_15059,N_14501,N_14663);
nand U15060 (N_15060,N_14749,N_14503);
nand U15061 (N_15061,N_14651,N_14413);
and U15062 (N_15062,N_14749,N_14686);
xnor U15063 (N_15063,N_14574,N_14561);
xnor U15064 (N_15064,N_14632,N_14445);
and U15065 (N_15065,N_14797,N_14464);
and U15066 (N_15066,N_14584,N_14675);
nand U15067 (N_15067,N_14717,N_14406);
xnor U15068 (N_15068,N_14490,N_14713);
or U15069 (N_15069,N_14680,N_14774);
xor U15070 (N_15070,N_14770,N_14436);
nand U15071 (N_15071,N_14447,N_14755);
nand U15072 (N_15072,N_14515,N_14650);
xor U15073 (N_15073,N_14744,N_14590);
and U15074 (N_15074,N_14583,N_14515);
nand U15075 (N_15075,N_14658,N_14745);
or U15076 (N_15076,N_14535,N_14523);
and U15077 (N_15077,N_14544,N_14550);
xor U15078 (N_15078,N_14720,N_14475);
nor U15079 (N_15079,N_14695,N_14597);
xnor U15080 (N_15080,N_14597,N_14566);
and U15081 (N_15081,N_14660,N_14612);
and U15082 (N_15082,N_14711,N_14721);
nand U15083 (N_15083,N_14499,N_14680);
nor U15084 (N_15084,N_14660,N_14733);
and U15085 (N_15085,N_14440,N_14549);
or U15086 (N_15086,N_14551,N_14595);
and U15087 (N_15087,N_14535,N_14649);
or U15088 (N_15088,N_14566,N_14540);
nand U15089 (N_15089,N_14400,N_14584);
nand U15090 (N_15090,N_14434,N_14461);
or U15091 (N_15091,N_14716,N_14515);
nand U15092 (N_15092,N_14558,N_14732);
or U15093 (N_15093,N_14618,N_14487);
xor U15094 (N_15094,N_14587,N_14730);
xnor U15095 (N_15095,N_14596,N_14578);
xor U15096 (N_15096,N_14491,N_14641);
nor U15097 (N_15097,N_14639,N_14561);
or U15098 (N_15098,N_14557,N_14657);
nor U15099 (N_15099,N_14683,N_14511);
xnor U15100 (N_15100,N_14685,N_14682);
and U15101 (N_15101,N_14497,N_14600);
nand U15102 (N_15102,N_14554,N_14792);
and U15103 (N_15103,N_14527,N_14550);
nor U15104 (N_15104,N_14647,N_14797);
xor U15105 (N_15105,N_14577,N_14695);
nor U15106 (N_15106,N_14656,N_14433);
xnor U15107 (N_15107,N_14617,N_14746);
nand U15108 (N_15108,N_14421,N_14778);
and U15109 (N_15109,N_14727,N_14552);
nand U15110 (N_15110,N_14588,N_14778);
nor U15111 (N_15111,N_14607,N_14730);
nor U15112 (N_15112,N_14420,N_14446);
or U15113 (N_15113,N_14686,N_14503);
or U15114 (N_15114,N_14414,N_14527);
nand U15115 (N_15115,N_14752,N_14524);
xnor U15116 (N_15116,N_14772,N_14597);
nor U15117 (N_15117,N_14647,N_14679);
xor U15118 (N_15118,N_14613,N_14758);
xor U15119 (N_15119,N_14452,N_14640);
xor U15120 (N_15120,N_14791,N_14761);
nand U15121 (N_15121,N_14753,N_14623);
nor U15122 (N_15122,N_14709,N_14690);
nor U15123 (N_15123,N_14565,N_14616);
nor U15124 (N_15124,N_14738,N_14417);
nand U15125 (N_15125,N_14400,N_14767);
or U15126 (N_15126,N_14572,N_14716);
or U15127 (N_15127,N_14553,N_14679);
and U15128 (N_15128,N_14700,N_14638);
xor U15129 (N_15129,N_14647,N_14535);
or U15130 (N_15130,N_14572,N_14487);
and U15131 (N_15131,N_14406,N_14554);
nand U15132 (N_15132,N_14750,N_14743);
and U15133 (N_15133,N_14755,N_14683);
nor U15134 (N_15134,N_14584,N_14576);
xor U15135 (N_15135,N_14778,N_14661);
nor U15136 (N_15136,N_14533,N_14406);
xnor U15137 (N_15137,N_14430,N_14776);
xnor U15138 (N_15138,N_14682,N_14486);
xor U15139 (N_15139,N_14678,N_14674);
or U15140 (N_15140,N_14401,N_14663);
nand U15141 (N_15141,N_14634,N_14708);
xor U15142 (N_15142,N_14458,N_14506);
xor U15143 (N_15143,N_14590,N_14660);
and U15144 (N_15144,N_14418,N_14659);
and U15145 (N_15145,N_14618,N_14629);
xnor U15146 (N_15146,N_14513,N_14701);
nand U15147 (N_15147,N_14665,N_14751);
and U15148 (N_15148,N_14442,N_14517);
and U15149 (N_15149,N_14662,N_14710);
xor U15150 (N_15150,N_14481,N_14670);
nand U15151 (N_15151,N_14477,N_14401);
nand U15152 (N_15152,N_14686,N_14730);
and U15153 (N_15153,N_14444,N_14767);
nand U15154 (N_15154,N_14490,N_14648);
nand U15155 (N_15155,N_14522,N_14755);
xor U15156 (N_15156,N_14515,N_14633);
nor U15157 (N_15157,N_14480,N_14780);
and U15158 (N_15158,N_14685,N_14559);
xor U15159 (N_15159,N_14562,N_14573);
nor U15160 (N_15160,N_14480,N_14729);
or U15161 (N_15161,N_14784,N_14787);
nor U15162 (N_15162,N_14699,N_14525);
nor U15163 (N_15163,N_14431,N_14474);
and U15164 (N_15164,N_14498,N_14550);
or U15165 (N_15165,N_14706,N_14547);
nand U15166 (N_15166,N_14484,N_14562);
and U15167 (N_15167,N_14581,N_14590);
nor U15168 (N_15168,N_14545,N_14627);
and U15169 (N_15169,N_14614,N_14405);
nand U15170 (N_15170,N_14772,N_14743);
and U15171 (N_15171,N_14492,N_14460);
nor U15172 (N_15172,N_14566,N_14799);
nor U15173 (N_15173,N_14491,N_14580);
nand U15174 (N_15174,N_14724,N_14692);
or U15175 (N_15175,N_14600,N_14518);
nor U15176 (N_15176,N_14651,N_14705);
xnor U15177 (N_15177,N_14773,N_14463);
and U15178 (N_15178,N_14664,N_14792);
nor U15179 (N_15179,N_14755,N_14729);
or U15180 (N_15180,N_14627,N_14410);
and U15181 (N_15181,N_14571,N_14768);
nor U15182 (N_15182,N_14537,N_14446);
nand U15183 (N_15183,N_14617,N_14492);
and U15184 (N_15184,N_14572,N_14755);
nand U15185 (N_15185,N_14620,N_14708);
nor U15186 (N_15186,N_14646,N_14698);
nand U15187 (N_15187,N_14443,N_14580);
nor U15188 (N_15188,N_14780,N_14466);
and U15189 (N_15189,N_14657,N_14792);
nor U15190 (N_15190,N_14451,N_14611);
xnor U15191 (N_15191,N_14668,N_14633);
nand U15192 (N_15192,N_14523,N_14556);
xnor U15193 (N_15193,N_14400,N_14474);
xnor U15194 (N_15194,N_14718,N_14480);
nor U15195 (N_15195,N_14728,N_14647);
or U15196 (N_15196,N_14616,N_14519);
nand U15197 (N_15197,N_14730,N_14716);
nor U15198 (N_15198,N_14452,N_14575);
nand U15199 (N_15199,N_14657,N_14740);
or U15200 (N_15200,N_15197,N_14955);
nand U15201 (N_15201,N_14845,N_14988);
xor U15202 (N_15202,N_15065,N_14917);
or U15203 (N_15203,N_14931,N_14956);
xnor U15204 (N_15204,N_14913,N_15087);
and U15205 (N_15205,N_14916,N_15157);
or U15206 (N_15206,N_14823,N_14922);
xor U15207 (N_15207,N_15166,N_15152);
xor U15208 (N_15208,N_14850,N_15039);
or U15209 (N_15209,N_14882,N_15002);
nand U15210 (N_15210,N_15124,N_14972);
and U15211 (N_15211,N_15110,N_15162);
xor U15212 (N_15212,N_14885,N_15154);
and U15213 (N_15213,N_15114,N_15125);
and U15214 (N_15214,N_14883,N_14892);
and U15215 (N_15215,N_15075,N_15074);
nor U15216 (N_15216,N_14984,N_14944);
and U15217 (N_15217,N_15186,N_15155);
xnor U15218 (N_15218,N_14868,N_15103);
nand U15219 (N_15219,N_15137,N_14964);
and U15220 (N_15220,N_14992,N_15144);
nor U15221 (N_15221,N_15097,N_14876);
nand U15222 (N_15222,N_14981,N_14848);
xor U15223 (N_15223,N_15175,N_15031);
nor U15224 (N_15224,N_14865,N_14836);
nand U15225 (N_15225,N_14896,N_15193);
or U15226 (N_15226,N_14838,N_15133);
nor U15227 (N_15227,N_15094,N_14903);
xnor U15228 (N_15228,N_14982,N_15026);
xnor U15229 (N_15229,N_15120,N_15138);
nand U15230 (N_15230,N_14849,N_15135);
nand U15231 (N_15231,N_15093,N_15195);
nand U15232 (N_15232,N_15053,N_15073);
nor U15233 (N_15233,N_14936,N_15111);
and U15234 (N_15234,N_15156,N_14857);
and U15235 (N_15235,N_14867,N_14897);
and U15236 (N_15236,N_14859,N_15005);
and U15237 (N_15237,N_14828,N_14800);
or U15238 (N_15238,N_15022,N_15079);
or U15239 (N_15239,N_14934,N_14844);
xor U15240 (N_15240,N_15088,N_14959);
and U15241 (N_15241,N_15109,N_14863);
xnor U15242 (N_15242,N_15149,N_14938);
or U15243 (N_15243,N_15061,N_15054);
nand U15244 (N_15244,N_14921,N_15107);
and U15245 (N_15245,N_15178,N_15176);
and U15246 (N_15246,N_15052,N_14958);
nor U15247 (N_15247,N_15092,N_14855);
nor U15248 (N_15248,N_14949,N_15196);
and U15249 (N_15249,N_14852,N_15100);
nor U15250 (N_15250,N_14830,N_14995);
or U15251 (N_15251,N_15150,N_15055);
xnor U15252 (N_15252,N_14975,N_15012);
xnor U15253 (N_15253,N_15001,N_14813);
nand U15254 (N_15254,N_14856,N_15113);
nand U15255 (N_15255,N_15188,N_15173);
nand U15256 (N_15256,N_15187,N_14895);
xor U15257 (N_15257,N_15011,N_14909);
nand U15258 (N_15258,N_15102,N_14977);
nand U15259 (N_15259,N_14821,N_15014);
or U15260 (N_15260,N_14967,N_14884);
xor U15261 (N_15261,N_15036,N_15051);
nor U15262 (N_15262,N_15082,N_14819);
nor U15263 (N_15263,N_14901,N_14918);
or U15264 (N_15264,N_14814,N_14969);
nor U15265 (N_15265,N_15078,N_15008);
or U15266 (N_15266,N_14999,N_15108);
nor U15267 (N_15267,N_15115,N_15122);
and U15268 (N_15268,N_15081,N_15153);
nand U15269 (N_15269,N_14846,N_14954);
nand U15270 (N_15270,N_15063,N_15059);
nand U15271 (N_15271,N_15198,N_14872);
nand U15272 (N_15272,N_14888,N_14866);
or U15273 (N_15273,N_15170,N_14947);
xor U15274 (N_15274,N_14809,N_15179);
and U15275 (N_15275,N_15046,N_15016);
and U15276 (N_15276,N_14841,N_15140);
nand U15277 (N_15277,N_15148,N_15091);
xnor U15278 (N_15278,N_14923,N_15030);
nor U15279 (N_15279,N_15067,N_15032);
xor U15280 (N_15280,N_15168,N_14968);
and U15281 (N_15281,N_14948,N_14802);
and U15282 (N_15282,N_15123,N_14812);
and U15283 (N_15283,N_14805,N_14930);
or U15284 (N_15284,N_15143,N_14932);
nor U15285 (N_15285,N_14861,N_14827);
or U15286 (N_15286,N_15177,N_14891);
nand U15287 (N_15287,N_15021,N_15112);
and U15288 (N_15288,N_15080,N_14879);
nand U15289 (N_15289,N_14824,N_15043);
nor U15290 (N_15290,N_15020,N_15104);
and U15291 (N_15291,N_15129,N_15062);
and U15292 (N_15292,N_14979,N_14878);
xnor U15293 (N_15293,N_14914,N_15007);
nand U15294 (N_15294,N_14900,N_15139);
xor U15295 (N_15295,N_15130,N_15047);
xor U15296 (N_15296,N_14816,N_14801);
and U15297 (N_15297,N_14925,N_15025);
nand U15298 (N_15298,N_15167,N_15131);
xnor U15299 (N_15299,N_14858,N_14832);
and U15300 (N_15300,N_14899,N_14989);
nand U15301 (N_15301,N_15182,N_15040);
xnor U15302 (N_15302,N_14890,N_14950);
xnor U15303 (N_15303,N_15069,N_14919);
nor U15304 (N_15304,N_15145,N_15105);
nor U15305 (N_15305,N_14893,N_14862);
and U15306 (N_15306,N_14902,N_15165);
or U15307 (N_15307,N_15164,N_15057);
nor U15308 (N_15308,N_15098,N_15141);
or U15309 (N_15309,N_15000,N_14808);
nand U15310 (N_15310,N_15158,N_14843);
nand U15311 (N_15311,N_14842,N_15049);
nor U15312 (N_15312,N_15024,N_14965);
or U15313 (N_15313,N_14957,N_15127);
xor U15314 (N_15314,N_14831,N_15060);
and U15315 (N_15315,N_14839,N_15023);
nor U15316 (N_15316,N_14973,N_15086);
or U15317 (N_15317,N_14822,N_15018);
nor U15318 (N_15318,N_14974,N_14875);
or U15319 (N_15319,N_14905,N_14810);
or U15320 (N_15320,N_14997,N_15003);
and U15321 (N_15321,N_15095,N_14961);
and U15322 (N_15322,N_15096,N_15027);
nand U15323 (N_15323,N_15126,N_15034);
and U15324 (N_15324,N_14880,N_15045);
nand U15325 (N_15325,N_14978,N_14829);
or U15326 (N_15326,N_15085,N_14987);
nand U15327 (N_15327,N_14985,N_14898);
nor U15328 (N_15328,N_15072,N_14894);
xor U15329 (N_15329,N_15010,N_15071);
xor U15330 (N_15330,N_15189,N_15048);
and U15331 (N_15331,N_15044,N_15090);
xnor U15332 (N_15332,N_14906,N_14818);
and U15333 (N_15333,N_14970,N_15190);
xor U15334 (N_15334,N_15171,N_14806);
or U15335 (N_15335,N_15159,N_14869);
xor U15336 (N_15336,N_15089,N_15169);
xor U15337 (N_15337,N_14953,N_15161);
nand U15338 (N_15338,N_15151,N_14920);
and U15339 (N_15339,N_14837,N_15042);
nand U15340 (N_15340,N_14915,N_15035);
or U15341 (N_15341,N_15119,N_14889);
nand U15342 (N_15342,N_14966,N_14986);
or U15343 (N_15343,N_15056,N_15068);
nor U15344 (N_15344,N_15101,N_14952);
xnor U15345 (N_15345,N_15064,N_15033);
xnor U15346 (N_15346,N_15160,N_14825);
nor U15347 (N_15347,N_14935,N_14817);
and U15348 (N_15348,N_14983,N_14912);
or U15349 (N_15349,N_14803,N_15106);
or U15350 (N_15350,N_15185,N_14951);
nand U15351 (N_15351,N_14976,N_14908);
xnor U15352 (N_15352,N_14820,N_15077);
nor U15353 (N_15353,N_14811,N_15192);
nor U15354 (N_15354,N_15134,N_14933);
nor U15355 (N_15355,N_15028,N_15172);
xnor U15356 (N_15356,N_15019,N_14991);
nor U15357 (N_15357,N_14939,N_15183);
nand U15358 (N_15358,N_15142,N_14874);
nor U15359 (N_15359,N_15099,N_15136);
xnor U15360 (N_15360,N_14864,N_15084);
nand U15361 (N_15361,N_15118,N_14853);
and U15362 (N_15362,N_14873,N_14854);
and U15363 (N_15363,N_14804,N_14871);
and U15364 (N_15364,N_14960,N_14834);
xnor U15365 (N_15365,N_15117,N_14928);
nor U15366 (N_15366,N_14926,N_15076);
and U15367 (N_15367,N_14870,N_15037);
nor U15368 (N_15368,N_15184,N_14910);
and U15369 (N_15369,N_15038,N_14907);
and U15370 (N_15370,N_14937,N_15006);
nand U15371 (N_15371,N_15009,N_15013);
nand U15372 (N_15372,N_14833,N_14980);
xnor U15373 (N_15373,N_15132,N_14963);
or U15374 (N_15374,N_15146,N_15128);
or U15375 (N_15375,N_15121,N_15017);
and U15376 (N_15376,N_14929,N_14924);
or U15377 (N_15377,N_14971,N_15163);
or U15378 (N_15378,N_14962,N_14994);
xnor U15379 (N_15379,N_15194,N_15070);
nor U15380 (N_15380,N_14881,N_14860);
nand U15381 (N_15381,N_14886,N_15015);
xor U15382 (N_15382,N_14945,N_14941);
nor U15383 (N_15383,N_15191,N_14993);
xnor U15384 (N_15384,N_14877,N_14911);
or U15385 (N_15385,N_14942,N_14940);
nand U15386 (N_15386,N_14996,N_14815);
or U15387 (N_15387,N_15083,N_14847);
and U15388 (N_15388,N_14927,N_14835);
nand U15389 (N_15389,N_15050,N_15004);
and U15390 (N_15390,N_14887,N_14807);
nor U15391 (N_15391,N_14946,N_15199);
xor U15392 (N_15392,N_15181,N_14851);
nand U15393 (N_15393,N_14840,N_14998);
or U15394 (N_15394,N_14943,N_14904);
or U15395 (N_15395,N_15066,N_15116);
or U15396 (N_15396,N_15174,N_15041);
xnor U15397 (N_15397,N_15058,N_14826);
and U15398 (N_15398,N_15029,N_14990);
and U15399 (N_15399,N_15147,N_15180);
and U15400 (N_15400,N_15055,N_15148);
nor U15401 (N_15401,N_14905,N_15179);
xor U15402 (N_15402,N_14826,N_15017);
nor U15403 (N_15403,N_15021,N_14902);
or U15404 (N_15404,N_15148,N_15186);
nand U15405 (N_15405,N_15181,N_14931);
xor U15406 (N_15406,N_15103,N_15083);
and U15407 (N_15407,N_15130,N_15010);
nor U15408 (N_15408,N_14978,N_15025);
nor U15409 (N_15409,N_14889,N_15020);
and U15410 (N_15410,N_14934,N_14975);
nand U15411 (N_15411,N_14976,N_14981);
nand U15412 (N_15412,N_15160,N_15044);
nor U15413 (N_15413,N_15013,N_15183);
nand U15414 (N_15414,N_14938,N_15026);
or U15415 (N_15415,N_15165,N_15025);
xor U15416 (N_15416,N_14805,N_15028);
nor U15417 (N_15417,N_15082,N_14988);
and U15418 (N_15418,N_15159,N_15062);
nor U15419 (N_15419,N_14989,N_14806);
or U15420 (N_15420,N_15194,N_14819);
or U15421 (N_15421,N_15096,N_15032);
nor U15422 (N_15422,N_15098,N_15097);
nor U15423 (N_15423,N_15148,N_14878);
nand U15424 (N_15424,N_14816,N_14935);
or U15425 (N_15425,N_14823,N_15051);
nand U15426 (N_15426,N_15068,N_15173);
nand U15427 (N_15427,N_14946,N_15101);
or U15428 (N_15428,N_15159,N_14960);
xnor U15429 (N_15429,N_15117,N_14807);
nor U15430 (N_15430,N_14859,N_14963);
nor U15431 (N_15431,N_14874,N_14871);
xor U15432 (N_15432,N_14936,N_15074);
xnor U15433 (N_15433,N_14800,N_15174);
and U15434 (N_15434,N_15023,N_14971);
or U15435 (N_15435,N_14829,N_15016);
xor U15436 (N_15436,N_14908,N_15091);
or U15437 (N_15437,N_14900,N_14890);
xor U15438 (N_15438,N_14915,N_14858);
nand U15439 (N_15439,N_14980,N_14937);
xnor U15440 (N_15440,N_14843,N_14898);
or U15441 (N_15441,N_14991,N_15136);
or U15442 (N_15442,N_15187,N_15049);
xor U15443 (N_15443,N_14894,N_15187);
and U15444 (N_15444,N_14914,N_15123);
xor U15445 (N_15445,N_15027,N_15054);
or U15446 (N_15446,N_14991,N_14810);
and U15447 (N_15447,N_15015,N_15177);
nand U15448 (N_15448,N_14949,N_15189);
and U15449 (N_15449,N_14864,N_14978);
nor U15450 (N_15450,N_15084,N_14834);
xor U15451 (N_15451,N_14906,N_15003);
or U15452 (N_15452,N_14935,N_14812);
or U15453 (N_15453,N_15129,N_14926);
nor U15454 (N_15454,N_15133,N_14947);
and U15455 (N_15455,N_15165,N_15172);
and U15456 (N_15456,N_15110,N_14807);
xnor U15457 (N_15457,N_14929,N_14982);
xor U15458 (N_15458,N_14993,N_15160);
nand U15459 (N_15459,N_15147,N_14839);
nand U15460 (N_15460,N_15196,N_15097);
nand U15461 (N_15461,N_14819,N_15002);
xor U15462 (N_15462,N_14929,N_14947);
or U15463 (N_15463,N_14931,N_15112);
and U15464 (N_15464,N_15049,N_15167);
xor U15465 (N_15465,N_14898,N_15163);
and U15466 (N_15466,N_15062,N_14943);
xor U15467 (N_15467,N_15199,N_15193);
nor U15468 (N_15468,N_14874,N_15023);
nand U15469 (N_15469,N_14968,N_14975);
or U15470 (N_15470,N_14852,N_14842);
xnor U15471 (N_15471,N_15007,N_15141);
nor U15472 (N_15472,N_14920,N_15163);
nand U15473 (N_15473,N_15021,N_14895);
xor U15474 (N_15474,N_15027,N_14814);
xor U15475 (N_15475,N_15129,N_14960);
xor U15476 (N_15476,N_15021,N_14814);
xor U15477 (N_15477,N_14938,N_14805);
and U15478 (N_15478,N_15153,N_14832);
or U15479 (N_15479,N_14994,N_15090);
nor U15480 (N_15480,N_15075,N_15190);
nand U15481 (N_15481,N_15068,N_15067);
or U15482 (N_15482,N_15039,N_14848);
and U15483 (N_15483,N_14992,N_14881);
or U15484 (N_15484,N_14803,N_15123);
and U15485 (N_15485,N_14837,N_14988);
or U15486 (N_15486,N_15123,N_15003);
nor U15487 (N_15487,N_14841,N_14823);
nor U15488 (N_15488,N_14809,N_14905);
xnor U15489 (N_15489,N_14876,N_14835);
nor U15490 (N_15490,N_15017,N_14894);
and U15491 (N_15491,N_14930,N_14925);
nor U15492 (N_15492,N_14864,N_14883);
nand U15493 (N_15493,N_14952,N_14904);
nor U15494 (N_15494,N_14850,N_14960);
nor U15495 (N_15495,N_14981,N_15152);
nor U15496 (N_15496,N_14835,N_14971);
nand U15497 (N_15497,N_15020,N_14933);
xnor U15498 (N_15498,N_14878,N_15000);
nand U15499 (N_15499,N_14851,N_14861);
nand U15500 (N_15500,N_15123,N_15011);
and U15501 (N_15501,N_14979,N_14942);
nor U15502 (N_15502,N_14836,N_15000);
nor U15503 (N_15503,N_15111,N_14912);
or U15504 (N_15504,N_15054,N_14801);
or U15505 (N_15505,N_15167,N_14991);
and U15506 (N_15506,N_15144,N_14990);
and U15507 (N_15507,N_14829,N_14850);
nor U15508 (N_15508,N_14861,N_14806);
or U15509 (N_15509,N_14913,N_15102);
nor U15510 (N_15510,N_15111,N_14868);
nor U15511 (N_15511,N_15034,N_14941);
nand U15512 (N_15512,N_15087,N_14889);
nor U15513 (N_15513,N_14870,N_14967);
nor U15514 (N_15514,N_15004,N_15077);
or U15515 (N_15515,N_15187,N_14825);
or U15516 (N_15516,N_15164,N_14855);
and U15517 (N_15517,N_15157,N_15034);
or U15518 (N_15518,N_14956,N_14998);
xor U15519 (N_15519,N_14936,N_14802);
or U15520 (N_15520,N_15030,N_15139);
nand U15521 (N_15521,N_14819,N_15166);
nor U15522 (N_15522,N_15191,N_14807);
or U15523 (N_15523,N_15176,N_14821);
or U15524 (N_15524,N_14968,N_14907);
and U15525 (N_15525,N_14882,N_14862);
or U15526 (N_15526,N_14867,N_15033);
or U15527 (N_15527,N_14952,N_15184);
or U15528 (N_15528,N_14949,N_15100);
or U15529 (N_15529,N_15093,N_14932);
nor U15530 (N_15530,N_14943,N_15179);
nand U15531 (N_15531,N_15008,N_15053);
or U15532 (N_15532,N_14856,N_15155);
or U15533 (N_15533,N_15185,N_15114);
or U15534 (N_15534,N_14971,N_15028);
xnor U15535 (N_15535,N_14810,N_14926);
and U15536 (N_15536,N_14950,N_14859);
nor U15537 (N_15537,N_14894,N_14947);
nand U15538 (N_15538,N_15139,N_14825);
xor U15539 (N_15539,N_15117,N_14864);
nor U15540 (N_15540,N_14825,N_15154);
and U15541 (N_15541,N_14897,N_14955);
nor U15542 (N_15542,N_15150,N_14857);
nor U15543 (N_15543,N_15117,N_15006);
or U15544 (N_15544,N_14910,N_15032);
nor U15545 (N_15545,N_14943,N_15121);
nand U15546 (N_15546,N_15199,N_14953);
xor U15547 (N_15547,N_14825,N_15034);
nand U15548 (N_15548,N_14860,N_15118);
or U15549 (N_15549,N_14896,N_15008);
or U15550 (N_15550,N_15179,N_14858);
and U15551 (N_15551,N_14964,N_14931);
xor U15552 (N_15552,N_15194,N_15017);
and U15553 (N_15553,N_14906,N_14948);
nand U15554 (N_15554,N_14912,N_14807);
nor U15555 (N_15555,N_14907,N_14895);
xnor U15556 (N_15556,N_15168,N_15173);
or U15557 (N_15557,N_15020,N_14942);
and U15558 (N_15558,N_15026,N_14960);
or U15559 (N_15559,N_15127,N_15034);
and U15560 (N_15560,N_15146,N_15008);
nor U15561 (N_15561,N_15155,N_14826);
xnor U15562 (N_15562,N_14852,N_14907);
nand U15563 (N_15563,N_14991,N_15098);
and U15564 (N_15564,N_14982,N_15133);
nor U15565 (N_15565,N_14916,N_14909);
nor U15566 (N_15566,N_15031,N_15199);
xor U15567 (N_15567,N_15149,N_15180);
and U15568 (N_15568,N_14879,N_14834);
nand U15569 (N_15569,N_14916,N_15077);
and U15570 (N_15570,N_14874,N_15157);
and U15571 (N_15571,N_15187,N_14905);
or U15572 (N_15572,N_15026,N_15025);
or U15573 (N_15573,N_15005,N_15100);
nor U15574 (N_15574,N_15095,N_14880);
and U15575 (N_15575,N_15064,N_14986);
nand U15576 (N_15576,N_14849,N_14862);
nor U15577 (N_15577,N_15127,N_14935);
nor U15578 (N_15578,N_14967,N_14895);
or U15579 (N_15579,N_14933,N_15073);
and U15580 (N_15580,N_15124,N_15112);
and U15581 (N_15581,N_14898,N_15051);
or U15582 (N_15582,N_15147,N_15108);
and U15583 (N_15583,N_14924,N_15090);
nor U15584 (N_15584,N_15002,N_14885);
xnor U15585 (N_15585,N_15126,N_14978);
and U15586 (N_15586,N_15109,N_15012);
xor U15587 (N_15587,N_15131,N_15156);
nand U15588 (N_15588,N_14840,N_15143);
nor U15589 (N_15589,N_14976,N_14961);
xnor U15590 (N_15590,N_14868,N_15153);
nor U15591 (N_15591,N_15041,N_14811);
nand U15592 (N_15592,N_14875,N_15008);
nor U15593 (N_15593,N_14850,N_15057);
nor U15594 (N_15594,N_15103,N_14855);
or U15595 (N_15595,N_14809,N_15081);
or U15596 (N_15596,N_14848,N_14943);
or U15597 (N_15597,N_15051,N_15140);
nor U15598 (N_15598,N_15068,N_15149);
nor U15599 (N_15599,N_14971,N_14856);
or U15600 (N_15600,N_15231,N_15405);
and U15601 (N_15601,N_15222,N_15540);
xor U15602 (N_15602,N_15300,N_15253);
xor U15603 (N_15603,N_15455,N_15219);
nor U15604 (N_15604,N_15557,N_15331);
nor U15605 (N_15605,N_15578,N_15213);
xor U15606 (N_15606,N_15533,N_15262);
nand U15607 (N_15607,N_15296,N_15221);
nand U15608 (N_15608,N_15456,N_15391);
xor U15609 (N_15609,N_15348,N_15305);
nand U15610 (N_15610,N_15401,N_15563);
xnor U15611 (N_15611,N_15543,N_15410);
xnor U15612 (N_15612,N_15528,N_15488);
nand U15613 (N_15613,N_15395,N_15498);
xor U15614 (N_15614,N_15582,N_15465);
nand U15615 (N_15615,N_15323,N_15400);
nand U15616 (N_15616,N_15408,N_15306);
or U15617 (N_15617,N_15469,N_15333);
nand U15618 (N_15618,N_15482,N_15491);
xnor U15619 (N_15619,N_15251,N_15449);
and U15620 (N_15620,N_15367,N_15249);
and U15621 (N_15621,N_15413,N_15335);
xor U15622 (N_15622,N_15329,N_15307);
and U15623 (N_15623,N_15585,N_15421);
nand U15624 (N_15624,N_15514,N_15217);
nand U15625 (N_15625,N_15243,N_15384);
nor U15626 (N_15626,N_15264,N_15404);
and U15627 (N_15627,N_15471,N_15555);
or U15628 (N_15628,N_15229,N_15261);
xor U15629 (N_15629,N_15587,N_15492);
and U15630 (N_15630,N_15226,N_15537);
nor U15631 (N_15631,N_15411,N_15366);
nor U15632 (N_15632,N_15561,N_15422);
nand U15633 (N_15633,N_15551,N_15420);
xor U15634 (N_15634,N_15228,N_15448);
nand U15635 (N_15635,N_15525,N_15398);
nor U15636 (N_15636,N_15278,N_15495);
and U15637 (N_15637,N_15504,N_15403);
and U15638 (N_15638,N_15216,N_15480);
nor U15639 (N_15639,N_15241,N_15355);
and U15640 (N_15640,N_15426,N_15344);
or U15641 (N_15641,N_15215,N_15326);
and U15642 (N_15642,N_15233,N_15444);
nor U15643 (N_15643,N_15499,N_15571);
nand U15644 (N_15644,N_15373,N_15599);
and U15645 (N_15645,N_15507,N_15479);
xor U15646 (N_15646,N_15409,N_15521);
and U15647 (N_15647,N_15211,N_15201);
nand U15648 (N_15648,N_15535,N_15266);
xor U15649 (N_15649,N_15531,N_15227);
xnor U15650 (N_15650,N_15283,N_15375);
nor U15651 (N_15651,N_15462,N_15496);
nor U15652 (N_15652,N_15595,N_15493);
and U15653 (N_15653,N_15477,N_15316);
or U15654 (N_15654,N_15402,N_15284);
and U15655 (N_15655,N_15354,N_15321);
nor U15656 (N_15656,N_15206,N_15327);
xnor U15657 (N_15657,N_15271,N_15285);
and U15658 (N_15658,N_15447,N_15268);
xnor U15659 (N_15659,N_15299,N_15476);
nor U15660 (N_15660,N_15439,N_15387);
nand U15661 (N_15661,N_15519,N_15220);
or U15662 (N_15662,N_15510,N_15553);
or U15663 (N_15663,N_15598,N_15236);
and U15664 (N_15664,N_15362,N_15350);
nor U15665 (N_15665,N_15451,N_15437);
xnor U15666 (N_15666,N_15513,N_15511);
nor U15667 (N_15667,N_15383,N_15516);
nor U15668 (N_15668,N_15260,N_15341);
or U15669 (N_15669,N_15548,N_15256);
nand U15670 (N_15670,N_15474,N_15419);
nand U15671 (N_15671,N_15542,N_15520);
xor U15672 (N_15672,N_15346,N_15460);
nand U15673 (N_15673,N_15390,N_15472);
nand U15674 (N_15674,N_15435,N_15596);
or U15675 (N_15675,N_15224,N_15290);
xor U15676 (N_15676,N_15225,N_15489);
or U15677 (N_15677,N_15397,N_15374);
or U15678 (N_15678,N_15255,N_15239);
nor U15679 (N_15679,N_15454,N_15450);
and U15680 (N_15680,N_15440,N_15240);
nand U15681 (N_15681,N_15443,N_15467);
nand U15682 (N_15682,N_15281,N_15274);
nand U15683 (N_15683,N_15351,N_15509);
or U15684 (N_15684,N_15342,N_15369);
xnor U15685 (N_15685,N_15297,N_15556);
or U15686 (N_15686,N_15396,N_15487);
nor U15687 (N_15687,N_15330,N_15379);
and U15688 (N_15688,N_15502,N_15526);
nand U15689 (N_15689,N_15433,N_15218);
nor U15690 (N_15690,N_15317,N_15545);
nand U15691 (N_15691,N_15386,N_15282);
and U15692 (N_15692,N_15212,N_15572);
xnor U15693 (N_15693,N_15592,N_15416);
nand U15694 (N_15694,N_15376,N_15358);
nor U15695 (N_15695,N_15432,N_15564);
or U15696 (N_15696,N_15392,N_15473);
nor U15697 (N_15697,N_15552,N_15505);
xor U15698 (N_15698,N_15328,N_15209);
nor U15699 (N_15699,N_15320,N_15470);
or U15700 (N_15700,N_15332,N_15265);
or U15701 (N_15701,N_15272,N_15588);
nor U15702 (N_15702,N_15590,N_15234);
or U15703 (N_15703,N_15325,N_15324);
or U15704 (N_15704,N_15315,N_15550);
xnor U15705 (N_15705,N_15573,N_15593);
and U15706 (N_15706,N_15353,N_15377);
xor U15707 (N_15707,N_15304,N_15244);
nand U15708 (N_15708,N_15583,N_15512);
nand U15709 (N_15709,N_15584,N_15273);
nand U15710 (N_15710,N_15501,N_15457);
nor U15711 (N_15711,N_15562,N_15279);
nor U15712 (N_15712,N_15277,N_15577);
or U15713 (N_15713,N_15356,N_15500);
xnor U15714 (N_15714,N_15204,N_15539);
xor U15715 (N_15715,N_15475,N_15478);
or U15716 (N_15716,N_15291,N_15532);
nor U15717 (N_15717,N_15257,N_15567);
and U15718 (N_15718,N_15490,N_15360);
nand U15719 (N_15719,N_15597,N_15293);
or U15720 (N_15720,N_15363,N_15589);
nand U15721 (N_15721,N_15276,N_15442);
xor U15722 (N_15722,N_15549,N_15560);
xnor U15723 (N_15723,N_15267,N_15263);
nand U15724 (N_15724,N_15246,N_15202);
and U15725 (N_15725,N_15436,N_15463);
or U15726 (N_15726,N_15530,N_15295);
and U15727 (N_15727,N_15591,N_15481);
nor U15728 (N_15728,N_15406,N_15494);
and U15729 (N_15729,N_15428,N_15286);
xor U15730 (N_15730,N_15298,N_15389);
nand U15731 (N_15731,N_15459,N_15523);
and U15732 (N_15732,N_15486,N_15461);
or U15733 (N_15733,N_15289,N_15245);
nand U15734 (N_15734,N_15287,N_15214);
and U15735 (N_15735,N_15361,N_15203);
and U15736 (N_15736,N_15349,N_15388);
and U15737 (N_15737,N_15575,N_15334);
and U15738 (N_15738,N_15312,N_15441);
and U15739 (N_15739,N_15415,N_15453);
nor U15740 (N_15740,N_15232,N_15207);
or U15741 (N_15741,N_15452,N_15337);
xor U15742 (N_15742,N_15538,N_15424);
nand U15743 (N_15743,N_15301,N_15536);
and U15744 (N_15744,N_15497,N_15529);
nor U15745 (N_15745,N_15414,N_15258);
nand U15746 (N_15746,N_15508,N_15485);
and U15747 (N_15747,N_15541,N_15412);
and U15748 (N_15748,N_15208,N_15368);
or U15749 (N_15749,N_15322,N_15468);
nand U15750 (N_15750,N_15527,N_15235);
and U15751 (N_15751,N_15546,N_15434);
or U15752 (N_15752,N_15483,N_15319);
and U15753 (N_15753,N_15230,N_15394);
or U15754 (N_15754,N_15423,N_15242);
and U15755 (N_15755,N_15576,N_15431);
nor U15756 (N_15756,N_15568,N_15418);
nor U15757 (N_15757,N_15464,N_15574);
and U15758 (N_15758,N_15314,N_15382);
or U15759 (N_15759,N_15503,N_15364);
or U15760 (N_15760,N_15370,N_15238);
nand U15761 (N_15761,N_15318,N_15292);
and U15762 (N_15762,N_15407,N_15569);
or U15763 (N_15763,N_15294,N_15399);
xor U15764 (N_15764,N_15237,N_15357);
xor U15765 (N_15765,N_15484,N_15200);
and U15766 (N_15766,N_15248,N_15247);
xnor U15767 (N_15767,N_15347,N_15378);
and U15768 (N_15768,N_15269,N_15581);
nor U15769 (N_15769,N_15427,N_15380);
nor U15770 (N_15770,N_15417,N_15566);
or U15771 (N_15771,N_15446,N_15345);
and U15772 (N_15772,N_15438,N_15558);
xor U15773 (N_15773,N_15515,N_15565);
nand U15774 (N_15774,N_15302,N_15559);
nand U15775 (N_15775,N_15466,N_15544);
or U15776 (N_15776,N_15303,N_15343);
nand U15777 (N_15777,N_15458,N_15425);
or U15778 (N_15778,N_15259,N_15594);
nor U15779 (N_15779,N_15547,N_15522);
and U15780 (N_15780,N_15359,N_15311);
and U15781 (N_15781,N_15205,N_15430);
nor U15782 (N_15782,N_15365,N_15586);
nor U15783 (N_15783,N_15313,N_15309);
nand U15784 (N_15784,N_15308,N_15385);
xor U15785 (N_15785,N_15554,N_15579);
nand U15786 (N_15786,N_15570,N_15336);
nor U15787 (N_15787,N_15338,N_15445);
or U15788 (N_15788,N_15506,N_15352);
and U15789 (N_15789,N_15223,N_15250);
or U15790 (N_15790,N_15340,N_15254);
nor U15791 (N_15791,N_15288,N_15275);
or U15792 (N_15792,N_15339,N_15393);
or U15793 (N_15793,N_15517,N_15270);
and U15794 (N_15794,N_15580,N_15518);
nor U15795 (N_15795,N_15524,N_15252);
nor U15796 (N_15796,N_15210,N_15310);
xor U15797 (N_15797,N_15429,N_15372);
and U15798 (N_15798,N_15280,N_15371);
nand U15799 (N_15799,N_15381,N_15534);
and U15800 (N_15800,N_15423,N_15330);
xor U15801 (N_15801,N_15589,N_15249);
nor U15802 (N_15802,N_15344,N_15329);
and U15803 (N_15803,N_15409,N_15488);
nor U15804 (N_15804,N_15307,N_15368);
or U15805 (N_15805,N_15491,N_15516);
or U15806 (N_15806,N_15360,N_15429);
and U15807 (N_15807,N_15509,N_15304);
and U15808 (N_15808,N_15288,N_15415);
and U15809 (N_15809,N_15508,N_15350);
and U15810 (N_15810,N_15538,N_15430);
nor U15811 (N_15811,N_15243,N_15240);
xor U15812 (N_15812,N_15598,N_15461);
xnor U15813 (N_15813,N_15236,N_15244);
xnor U15814 (N_15814,N_15549,N_15521);
or U15815 (N_15815,N_15323,N_15575);
nor U15816 (N_15816,N_15293,N_15507);
nand U15817 (N_15817,N_15418,N_15348);
nand U15818 (N_15818,N_15250,N_15392);
nand U15819 (N_15819,N_15411,N_15248);
or U15820 (N_15820,N_15245,N_15569);
and U15821 (N_15821,N_15231,N_15589);
nor U15822 (N_15822,N_15261,N_15424);
nand U15823 (N_15823,N_15280,N_15401);
nand U15824 (N_15824,N_15384,N_15209);
xnor U15825 (N_15825,N_15565,N_15546);
or U15826 (N_15826,N_15337,N_15403);
or U15827 (N_15827,N_15497,N_15215);
and U15828 (N_15828,N_15444,N_15210);
and U15829 (N_15829,N_15581,N_15414);
nand U15830 (N_15830,N_15442,N_15595);
xor U15831 (N_15831,N_15480,N_15287);
or U15832 (N_15832,N_15231,N_15324);
nand U15833 (N_15833,N_15202,N_15413);
and U15834 (N_15834,N_15459,N_15302);
or U15835 (N_15835,N_15237,N_15244);
and U15836 (N_15836,N_15402,N_15285);
nor U15837 (N_15837,N_15362,N_15255);
xnor U15838 (N_15838,N_15386,N_15558);
nor U15839 (N_15839,N_15408,N_15293);
nand U15840 (N_15840,N_15248,N_15530);
nand U15841 (N_15841,N_15331,N_15366);
or U15842 (N_15842,N_15515,N_15491);
and U15843 (N_15843,N_15571,N_15258);
or U15844 (N_15844,N_15285,N_15338);
nor U15845 (N_15845,N_15250,N_15238);
nand U15846 (N_15846,N_15301,N_15397);
and U15847 (N_15847,N_15423,N_15542);
nor U15848 (N_15848,N_15257,N_15574);
xnor U15849 (N_15849,N_15248,N_15590);
nand U15850 (N_15850,N_15383,N_15441);
nor U15851 (N_15851,N_15515,N_15449);
xor U15852 (N_15852,N_15330,N_15550);
xor U15853 (N_15853,N_15256,N_15574);
xor U15854 (N_15854,N_15518,N_15506);
or U15855 (N_15855,N_15457,N_15347);
xor U15856 (N_15856,N_15481,N_15426);
or U15857 (N_15857,N_15245,N_15561);
xor U15858 (N_15858,N_15239,N_15267);
nor U15859 (N_15859,N_15307,N_15407);
nor U15860 (N_15860,N_15563,N_15375);
xor U15861 (N_15861,N_15376,N_15535);
or U15862 (N_15862,N_15267,N_15510);
nand U15863 (N_15863,N_15269,N_15332);
or U15864 (N_15864,N_15509,N_15581);
or U15865 (N_15865,N_15367,N_15421);
or U15866 (N_15866,N_15322,N_15260);
and U15867 (N_15867,N_15597,N_15580);
and U15868 (N_15868,N_15318,N_15505);
nand U15869 (N_15869,N_15324,N_15395);
nand U15870 (N_15870,N_15591,N_15435);
or U15871 (N_15871,N_15425,N_15238);
or U15872 (N_15872,N_15365,N_15585);
or U15873 (N_15873,N_15216,N_15295);
nand U15874 (N_15874,N_15451,N_15209);
nand U15875 (N_15875,N_15455,N_15241);
xor U15876 (N_15876,N_15534,N_15340);
nand U15877 (N_15877,N_15506,N_15241);
and U15878 (N_15878,N_15453,N_15253);
or U15879 (N_15879,N_15326,N_15236);
and U15880 (N_15880,N_15302,N_15417);
and U15881 (N_15881,N_15407,N_15286);
nor U15882 (N_15882,N_15491,N_15255);
nor U15883 (N_15883,N_15454,N_15377);
nor U15884 (N_15884,N_15368,N_15433);
xnor U15885 (N_15885,N_15310,N_15583);
nand U15886 (N_15886,N_15536,N_15226);
nand U15887 (N_15887,N_15579,N_15498);
xor U15888 (N_15888,N_15334,N_15306);
xor U15889 (N_15889,N_15347,N_15359);
or U15890 (N_15890,N_15261,N_15577);
xnor U15891 (N_15891,N_15357,N_15298);
nor U15892 (N_15892,N_15266,N_15482);
and U15893 (N_15893,N_15422,N_15433);
xor U15894 (N_15894,N_15537,N_15498);
nor U15895 (N_15895,N_15379,N_15243);
nand U15896 (N_15896,N_15357,N_15584);
nand U15897 (N_15897,N_15397,N_15261);
nor U15898 (N_15898,N_15527,N_15495);
and U15899 (N_15899,N_15475,N_15346);
nand U15900 (N_15900,N_15311,N_15375);
or U15901 (N_15901,N_15519,N_15347);
or U15902 (N_15902,N_15372,N_15318);
and U15903 (N_15903,N_15395,N_15237);
or U15904 (N_15904,N_15247,N_15356);
and U15905 (N_15905,N_15545,N_15511);
xor U15906 (N_15906,N_15532,N_15333);
and U15907 (N_15907,N_15574,N_15485);
nor U15908 (N_15908,N_15413,N_15423);
or U15909 (N_15909,N_15528,N_15489);
nand U15910 (N_15910,N_15338,N_15342);
and U15911 (N_15911,N_15529,N_15315);
and U15912 (N_15912,N_15440,N_15264);
or U15913 (N_15913,N_15441,N_15459);
or U15914 (N_15914,N_15456,N_15254);
and U15915 (N_15915,N_15545,N_15260);
and U15916 (N_15916,N_15490,N_15582);
and U15917 (N_15917,N_15320,N_15235);
nand U15918 (N_15918,N_15428,N_15274);
xor U15919 (N_15919,N_15282,N_15396);
and U15920 (N_15920,N_15251,N_15554);
and U15921 (N_15921,N_15380,N_15382);
xnor U15922 (N_15922,N_15478,N_15560);
or U15923 (N_15923,N_15328,N_15315);
nand U15924 (N_15924,N_15267,N_15250);
and U15925 (N_15925,N_15502,N_15385);
nand U15926 (N_15926,N_15359,N_15383);
nor U15927 (N_15927,N_15219,N_15257);
and U15928 (N_15928,N_15311,N_15259);
nand U15929 (N_15929,N_15262,N_15431);
nor U15930 (N_15930,N_15260,N_15334);
or U15931 (N_15931,N_15421,N_15547);
nand U15932 (N_15932,N_15324,N_15306);
or U15933 (N_15933,N_15249,N_15414);
xnor U15934 (N_15934,N_15529,N_15306);
nor U15935 (N_15935,N_15276,N_15304);
and U15936 (N_15936,N_15307,N_15281);
or U15937 (N_15937,N_15330,N_15254);
or U15938 (N_15938,N_15220,N_15474);
xnor U15939 (N_15939,N_15264,N_15546);
and U15940 (N_15940,N_15436,N_15385);
or U15941 (N_15941,N_15417,N_15540);
xnor U15942 (N_15942,N_15587,N_15444);
xnor U15943 (N_15943,N_15456,N_15353);
nand U15944 (N_15944,N_15203,N_15377);
nand U15945 (N_15945,N_15211,N_15484);
or U15946 (N_15946,N_15429,N_15402);
or U15947 (N_15947,N_15361,N_15267);
xnor U15948 (N_15948,N_15350,N_15511);
nand U15949 (N_15949,N_15335,N_15281);
nor U15950 (N_15950,N_15496,N_15399);
nand U15951 (N_15951,N_15363,N_15550);
nand U15952 (N_15952,N_15292,N_15547);
or U15953 (N_15953,N_15470,N_15474);
and U15954 (N_15954,N_15454,N_15228);
nor U15955 (N_15955,N_15399,N_15272);
and U15956 (N_15956,N_15599,N_15552);
or U15957 (N_15957,N_15210,N_15511);
nor U15958 (N_15958,N_15563,N_15570);
and U15959 (N_15959,N_15288,N_15530);
or U15960 (N_15960,N_15585,N_15271);
and U15961 (N_15961,N_15293,N_15480);
and U15962 (N_15962,N_15229,N_15561);
nor U15963 (N_15963,N_15322,N_15236);
xnor U15964 (N_15964,N_15532,N_15200);
or U15965 (N_15965,N_15341,N_15350);
nand U15966 (N_15966,N_15226,N_15248);
or U15967 (N_15967,N_15344,N_15285);
xnor U15968 (N_15968,N_15350,N_15578);
and U15969 (N_15969,N_15282,N_15556);
and U15970 (N_15970,N_15267,N_15310);
or U15971 (N_15971,N_15260,N_15517);
xnor U15972 (N_15972,N_15203,N_15535);
nand U15973 (N_15973,N_15386,N_15519);
xnor U15974 (N_15974,N_15372,N_15524);
nor U15975 (N_15975,N_15384,N_15473);
and U15976 (N_15976,N_15514,N_15376);
and U15977 (N_15977,N_15518,N_15468);
or U15978 (N_15978,N_15372,N_15573);
and U15979 (N_15979,N_15428,N_15589);
and U15980 (N_15980,N_15410,N_15289);
or U15981 (N_15981,N_15483,N_15508);
or U15982 (N_15982,N_15499,N_15532);
nand U15983 (N_15983,N_15264,N_15237);
nand U15984 (N_15984,N_15456,N_15321);
nor U15985 (N_15985,N_15517,N_15589);
or U15986 (N_15986,N_15419,N_15538);
nand U15987 (N_15987,N_15447,N_15207);
xnor U15988 (N_15988,N_15215,N_15280);
or U15989 (N_15989,N_15332,N_15369);
or U15990 (N_15990,N_15533,N_15201);
xor U15991 (N_15991,N_15537,N_15427);
or U15992 (N_15992,N_15392,N_15358);
and U15993 (N_15993,N_15262,N_15278);
xnor U15994 (N_15994,N_15522,N_15309);
xnor U15995 (N_15995,N_15532,N_15428);
xor U15996 (N_15996,N_15232,N_15383);
nand U15997 (N_15997,N_15309,N_15377);
xnor U15998 (N_15998,N_15242,N_15289);
and U15999 (N_15999,N_15395,N_15311);
xnor U16000 (N_16000,N_15808,N_15905);
or U16001 (N_16001,N_15797,N_15867);
and U16002 (N_16002,N_15823,N_15966);
xnor U16003 (N_16003,N_15718,N_15914);
nor U16004 (N_16004,N_15950,N_15902);
or U16005 (N_16005,N_15936,N_15999);
nand U16006 (N_16006,N_15657,N_15689);
nand U16007 (N_16007,N_15772,N_15921);
nand U16008 (N_16008,N_15782,N_15899);
or U16009 (N_16009,N_15670,N_15716);
xnor U16010 (N_16010,N_15763,N_15770);
xnor U16011 (N_16011,N_15774,N_15631);
or U16012 (N_16012,N_15813,N_15912);
and U16013 (N_16013,N_15788,N_15668);
or U16014 (N_16014,N_15874,N_15858);
and U16015 (N_16015,N_15927,N_15671);
xor U16016 (N_16016,N_15928,N_15614);
nand U16017 (N_16017,N_15913,N_15651);
nor U16018 (N_16018,N_15892,N_15962);
nor U16019 (N_16019,N_15849,N_15649);
nor U16020 (N_16020,N_15674,N_15945);
or U16021 (N_16021,N_15794,N_15617);
xnor U16022 (N_16022,N_15731,N_15854);
or U16023 (N_16023,N_15916,N_15604);
and U16024 (N_16024,N_15910,N_15785);
or U16025 (N_16025,N_15618,N_15876);
nor U16026 (N_16026,N_15663,N_15822);
nor U16027 (N_16027,N_15795,N_15694);
nor U16028 (N_16028,N_15812,N_15969);
nor U16029 (N_16029,N_15977,N_15690);
or U16030 (N_16030,N_15642,N_15881);
and U16031 (N_16031,N_15627,N_15875);
or U16032 (N_16032,N_15971,N_15850);
and U16033 (N_16033,N_15766,N_15641);
or U16034 (N_16034,N_15717,N_15890);
and U16035 (N_16035,N_15833,N_15681);
nor U16036 (N_16036,N_15883,N_15920);
or U16037 (N_16037,N_15778,N_15719);
nand U16038 (N_16038,N_15817,N_15853);
xnor U16039 (N_16039,N_15806,N_15838);
or U16040 (N_16040,N_15915,N_15987);
nand U16041 (N_16041,N_15677,N_15861);
xnor U16042 (N_16042,N_15897,N_15815);
nand U16043 (N_16043,N_15746,N_15870);
and U16044 (N_16044,N_15807,N_15738);
nor U16045 (N_16045,N_15675,N_15611);
and U16046 (N_16046,N_15843,N_15798);
or U16047 (N_16047,N_15931,N_15608);
nor U16048 (N_16048,N_15981,N_15992);
nor U16049 (N_16049,N_15852,N_15697);
xnor U16050 (N_16050,N_15740,N_15634);
or U16051 (N_16051,N_15877,N_15684);
and U16052 (N_16052,N_15848,N_15702);
or U16053 (N_16053,N_15695,N_15789);
or U16054 (N_16054,N_15868,N_15669);
xor U16055 (N_16055,N_15622,N_15722);
and U16056 (N_16056,N_15647,N_15776);
and U16057 (N_16057,N_15748,N_15872);
nor U16058 (N_16058,N_15687,N_15894);
or U16059 (N_16059,N_15990,N_15654);
nand U16060 (N_16060,N_15643,N_15715);
or U16061 (N_16061,N_15660,N_15781);
nor U16062 (N_16062,N_15942,N_15696);
xnor U16063 (N_16063,N_15636,N_15831);
xor U16064 (N_16064,N_15946,N_15811);
xnor U16065 (N_16065,N_15836,N_15683);
xor U16066 (N_16066,N_15994,N_15873);
xor U16067 (N_16067,N_15835,N_15821);
and U16068 (N_16068,N_15954,N_15984);
nand U16069 (N_16069,N_15713,N_15855);
nand U16070 (N_16070,N_15814,N_15603);
nand U16071 (N_16071,N_15924,N_15964);
xnor U16072 (N_16072,N_15919,N_15941);
nand U16073 (N_16073,N_15628,N_15693);
or U16074 (N_16074,N_15613,N_15819);
or U16075 (N_16075,N_15620,N_15757);
and U16076 (N_16076,N_15648,N_15727);
nor U16077 (N_16077,N_15704,N_15792);
nor U16078 (N_16078,N_15767,N_15830);
and U16079 (N_16079,N_15885,N_15764);
and U16080 (N_16080,N_15955,N_15856);
nand U16081 (N_16081,N_15989,N_15908);
nor U16082 (N_16082,N_15653,N_15923);
xor U16083 (N_16083,N_15975,N_15735);
and U16084 (N_16084,N_15956,N_15625);
and U16085 (N_16085,N_15898,N_15827);
nor U16086 (N_16086,N_15650,N_15786);
nor U16087 (N_16087,N_15859,N_15932);
and U16088 (N_16088,N_15829,N_15646);
and U16089 (N_16089,N_15633,N_15739);
xnor U16090 (N_16090,N_15879,N_15880);
nand U16091 (N_16091,N_15726,N_15865);
nand U16092 (N_16092,N_15601,N_15723);
and U16093 (N_16093,N_15972,N_15685);
or U16094 (N_16094,N_15623,N_15733);
xnor U16095 (N_16095,N_15711,N_15841);
and U16096 (N_16096,N_15790,N_15667);
or U16097 (N_16097,N_15791,N_15729);
and U16098 (N_16098,N_15743,N_15688);
and U16099 (N_16099,N_15960,N_15679);
xnor U16100 (N_16100,N_15871,N_15991);
or U16101 (N_16101,N_15672,N_15754);
and U16102 (N_16102,N_15953,N_15707);
and U16103 (N_16103,N_15665,N_15607);
xnor U16104 (N_16104,N_15918,N_15673);
or U16105 (N_16105,N_15706,N_15606);
xor U16106 (N_16106,N_15804,N_15737);
nor U16107 (N_16107,N_15692,N_15760);
xnor U16108 (N_16108,N_15957,N_15976);
xnor U16109 (N_16109,N_15952,N_15970);
xnor U16110 (N_16110,N_15997,N_15878);
nor U16111 (N_16111,N_15619,N_15869);
xor U16112 (N_16112,N_15917,N_15762);
and U16113 (N_16113,N_15904,N_15832);
and U16114 (N_16114,N_15745,N_15780);
xnor U16115 (N_16115,N_15837,N_15980);
and U16116 (N_16116,N_15828,N_15886);
nor U16117 (N_16117,N_15610,N_15996);
and U16118 (N_16118,N_15775,N_15901);
nor U16119 (N_16119,N_15751,N_15771);
nor U16120 (N_16120,N_15985,N_15664);
nor U16121 (N_16121,N_15777,N_15720);
and U16122 (N_16122,N_15699,N_15632);
and U16123 (N_16123,N_15965,N_15640);
and U16124 (N_16124,N_15686,N_15948);
nand U16125 (N_16125,N_15802,N_15982);
and U16126 (N_16126,N_15721,N_15995);
nor U16127 (N_16127,N_15734,N_15656);
nor U16128 (N_16128,N_15609,N_15926);
nand U16129 (N_16129,N_15978,N_15658);
and U16130 (N_16130,N_15624,N_15967);
xnor U16131 (N_16131,N_15616,N_15661);
or U16132 (N_16132,N_15801,N_15736);
xor U16133 (N_16133,N_15810,N_15612);
and U16134 (N_16134,N_15968,N_15889);
nor U16135 (N_16135,N_15973,N_15700);
and U16136 (N_16136,N_15787,N_15783);
nand U16137 (N_16137,N_15993,N_15750);
xnor U16138 (N_16138,N_15756,N_15834);
nor U16139 (N_16139,N_15799,N_15851);
nor U16140 (N_16140,N_15710,N_15714);
xnor U16141 (N_16141,N_15698,N_15730);
xnor U16142 (N_16142,N_15949,N_15638);
or U16143 (N_16143,N_15680,N_15888);
and U16144 (N_16144,N_15796,N_15988);
nor U16145 (N_16145,N_15842,N_15630);
nand U16146 (N_16146,N_15891,N_15826);
or U16147 (N_16147,N_15896,N_15705);
nor U16148 (N_16148,N_15906,N_15963);
nor U16149 (N_16149,N_15629,N_15742);
and U16150 (N_16150,N_15758,N_15895);
xnor U16151 (N_16151,N_15882,N_15749);
nor U16152 (N_16152,N_15933,N_15784);
or U16153 (N_16153,N_15864,N_15947);
nand U16154 (N_16154,N_15943,N_15925);
nand U16155 (N_16155,N_15983,N_15708);
nand U16156 (N_16156,N_15844,N_15659);
or U16157 (N_16157,N_15986,N_15884);
xnor U16158 (N_16158,N_15602,N_15959);
or U16159 (N_16159,N_15635,N_15958);
and U16160 (N_16160,N_15605,N_15655);
and U16161 (N_16161,N_15860,N_15809);
nand U16162 (N_16162,N_15759,N_15761);
nor U16163 (N_16163,N_15682,N_15845);
and U16164 (N_16164,N_15839,N_15626);
or U16165 (N_16165,N_15863,N_15678);
nor U16166 (N_16166,N_15752,N_15816);
nor U16167 (N_16167,N_15937,N_15951);
nand U16168 (N_16168,N_15747,N_15600);
xnor U16169 (N_16169,N_15857,N_15847);
xnor U16170 (N_16170,N_15911,N_15922);
nand U16171 (N_16171,N_15753,N_15769);
nor U16172 (N_16172,N_15755,N_15765);
nand U16173 (N_16173,N_15930,N_15741);
nor U16174 (N_16174,N_15793,N_15666);
xnor U16175 (N_16175,N_15805,N_15862);
xor U16176 (N_16176,N_15724,N_15998);
nand U16177 (N_16177,N_15637,N_15800);
nand U16178 (N_16178,N_15979,N_15615);
nand U16179 (N_16179,N_15961,N_15909);
or U16180 (N_16180,N_15929,N_15691);
xnor U16181 (N_16181,N_15676,N_15974);
or U16182 (N_16182,N_15840,N_15744);
nor U16183 (N_16183,N_15732,N_15621);
or U16184 (N_16184,N_15935,N_15645);
and U16185 (N_16185,N_15820,N_15803);
nor U16186 (N_16186,N_15725,N_15779);
and U16187 (N_16187,N_15703,N_15887);
or U16188 (N_16188,N_15846,N_15825);
xor U16189 (N_16189,N_15639,N_15818);
nand U16190 (N_16190,N_15934,N_15644);
or U16191 (N_16191,N_15939,N_15903);
and U16192 (N_16192,N_15940,N_15944);
or U16193 (N_16193,N_15907,N_15866);
xnor U16194 (N_16194,N_15662,N_15701);
nor U16195 (N_16195,N_15773,N_15728);
or U16196 (N_16196,N_15938,N_15709);
nor U16197 (N_16197,N_15900,N_15893);
or U16198 (N_16198,N_15652,N_15824);
xnor U16199 (N_16199,N_15768,N_15712);
and U16200 (N_16200,N_15834,N_15825);
nor U16201 (N_16201,N_15915,N_15855);
and U16202 (N_16202,N_15627,N_15920);
nand U16203 (N_16203,N_15763,N_15653);
or U16204 (N_16204,N_15756,N_15844);
xor U16205 (N_16205,N_15654,N_15635);
nand U16206 (N_16206,N_15915,N_15752);
and U16207 (N_16207,N_15645,N_15910);
and U16208 (N_16208,N_15843,N_15670);
xor U16209 (N_16209,N_15730,N_15896);
nor U16210 (N_16210,N_15913,N_15992);
nand U16211 (N_16211,N_15651,N_15719);
and U16212 (N_16212,N_15636,N_15791);
nand U16213 (N_16213,N_15995,N_15630);
nand U16214 (N_16214,N_15764,N_15744);
xnor U16215 (N_16215,N_15943,N_15968);
nand U16216 (N_16216,N_15888,N_15654);
nor U16217 (N_16217,N_15937,N_15835);
nand U16218 (N_16218,N_15659,N_15709);
nor U16219 (N_16219,N_15615,N_15934);
or U16220 (N_16220,N_15698,N_15823);
nor U16221 (N_16221,N_15948,N_15840);
or U16222 (N_16222,N_15652,N_15624);
xnor U16223 (N_16223,N_15835,N_15890);
or U16224 (N_16224,N_15937,N_15898);
or U16225 (N_16225,N_15991,N_15934);
nor U16226 (N_16226,N_15721,N_15909);
nor U16227 (N_16227,N_15667,N_15873);
nand U16228 (N_16228,N_15747,N_15973);
nor U16229 (N_16229,N_15726,N_15975);
nor U16230 (N_16230,N_15836,N_15997);
nand U16231 (N_16231,N_15824,N_15712);
or U16232 (N_16232,N_15809,N_15741);
and U16233 (N_16233,N_15757,N_15774);
and U16234 (N_16234,N_15974,N_15935);
and U16235 (N_16235,N_15818,N_15620);
and U16236 (N_16236,N_15924,N_15847);
xnor U16237 (N_16237,N_15674,N_15608);
and U16238 (N_16238,N_15653,N_15767);
and U16239 (N_16239,N_15646,N_15756);
and U16240 (N_16240,N_15865,N_15844);
nand U16241 (N_16241,N_15756,N_15960);
nor U16242 (N_16242,N_15893,N_15928);
and U16243 (N_16243,N_15740,N_15905);
and U16244 (N_16244,N_15935,N_15916);
xor U16245 (N_16245,N_15690,N_15660);
and U16246 (N_16246,N_15602,N_15807);
and U16247 (N_16247,N_15934,N_15865);
and U16248 (N_16248,N_15668,N_15980);
and U16249 (N_16249,N_15685,N_15637);
nor U16250 (N_16250,N_15812,N_15903);
xnor U16251 (N_16251,N_15647,N_15635);
or U16252 (N_16252,N_15821,N_15625);
xor U16253 (N_16253,N_15817,N_15618);
xor U16254 (N_16254,N_15789,N_15946);
or U16255 (N_16255,N_15974,N_15809);
or U16256 (N_16256,N_15809,N_15779);
nor U16257 (N_16257,N_15686,N_15970);
nand U16258 (N_16258,N_15878,N_15673);
nand U16259 (N_16259,N_15743,N_15677);
nor U16260 (N_16260,N_15875,N_15993);
and U16261 (N_16261,N_15634,N_15659);
nor U16262 (N_16262,N_15739,N_15889);
and U16263 (N_16263,N_15685,N_15665);
nand U16264 (N_16264,N_15935,N_15902);
xnor U16265 (N_16265,N_15943,N_15838);
or U16266 (N_16266,N_15899,N_15840);
nor U16267 (N_16267,N_15860,N_15776);
nor U16268 (N_16268,N_15815,N_15842);
nand U16269 (N_16269,N_15863,N_15707);
xor U16270 (N_16270,N_15631,N_15636);
nor U16271 (N_16271,N_15793,N_15795);
and U16272 (N_16272,N_15780,N_15849);
xnor U16273 (N_16273,N_15752,N_15948);
or U16274 (N_16274,N_15876,N_15833);
or U16275 (N_16275,N_15724,N_15849);
and U16276 (N_16276,N_15880,N_15903);
and U16277 (N_16277,N_15624,N_15948);
nor U16278 (N_16278,N_15689,N_15889);
nand U16279 (N_16279,N_15789,N_15896);
nor U16280 (N_16280,N_15984,N_15685);
nor U16281 (N_16281,N_15856,N_15754);
nor U16282 (N_16282,N_15604,N_15924);
or U16283 (N_16283,N_15904,N_15980);
or U16284 (N_16284,N_15867,N_15837);
nor U16285 (N_16285,N_15855,N_15925);
nand U16286 (N_16286,N_15667,N_15794);
or U16287 (N_16287,N_15992,N_15845);
and U16288 (N_16288,N_15633,N_15614);
and U16289 (N_16289,N_15927,N_15901);
or U16290 (N_16290,N_15892,N_15715);
or U16291 (N_16291,N_15768,N_15726);
nand U16292 (N_16292,N_15998,N_15973);
xnor U16293 (N_16293,N_15644,N_15627);
nor U16294 (N_16294,N_15818,N_15740);
nor U16295 (N_16295,N_15857,N_15959);
and U16296 (N_16296,N_15873,N_15746);
xnor U16297 (N_16297,N_15799,N_15903);
nor U16298 (N_16298,N_15670,N_15896);
and U16299 (N_16299,N_15651,N_15756);
and U16300 (N_16300,N_15786,N_15729);
or U16301 (N_16301,N_15786,N_15941);
xnor U16302 (N_16302,N_15631,N_15632);
xnor U16303 (N_16303,N_15616,N_15707);
nand U16304 (N_16304,N_15628,N_15918);
and U16305 (N_16305,N_15836,N_15633);
nand U16306 (N_16306,N_15677,N_15835);
and U16307 (N_16307,N_15691,N_15940);
nor U16308 (N_16308,N_15712,N_15757);
or U16309 (N_16309,N_15854,N_15696);
or U16310 (N_16310,N_15869,N_15692);
nand U16311 (N_16311,N_15784,N_15859);
nand U16312 (N_16312,N_15618,N_15873);
nor U16313 (N_16313,N_15785,N_15740);
xor U16314 (N_16314,N_15952,N_15754);
nor U16315 (N_16315,N_15726,N_15738);
xnor U16316 (N_16316,N_15830,N_15746);
nand U16317 (N_16317,N_15766,N_15915);
nand U16318 (N_16318,N_15932,N_15783);
or U16319 (N_16319,N_15884,N_15605);
or U16320 (N_16320,N_15673,N_15616);
and U16321 (N_16321,N_15626,N_15870);
nor U16322 (N_16322,N_15767,N_15724);
nand U16323 (N_16323,N_15982,N_15959);
or U16324 (N_16324,N_15628,N_15812);
and U16325 (N_16325,N_15602,N_15847);
nand U16326 (N_16326,N_15676,N_15953);
xor U16327 (N_16327,N_15790,N_15718);
or U16328 (N_16328,N_15822,N_15610);
nor U16329 (N_16329,N_15842,N_15910);
nand U16330 (N_16330,N_15856,N_15882);
or U16331 (N_16331,N_15805,N_15747);
nor U16332 (N_16332,N_15815,N_15693);
nand U16333 (N_16333,N_15609,N_15616);
and U16334 (N_16334,N_15636,N_15931);
or U16335 (N_16335,N_15667,N_15622);
or U16336 (N_16336,N_15946,N_15686);
nor U16337 (N_16337,N_15935,N_15789);
nand U16338 (N_16338,N_15897,N_15856);
xnor U16339 (N_16339,N_15635,N_15874);
nand U16340 (N_16340,N_15623,N_15709);
xnor U16341 (N_16341,N_15991,N_15989);
xnor U16342 (N_16342,N_15722,N_15737);
nand U16343 (N_16343,N_15915,N_15763);
and U16344 (N_16344,N_15619,N_15747);
and U16345 (N_16345,N_15642,N_15804);
xor U16346 (N_16346,N_15782,N_15670);
nand U16347 (N_16347,N_15967,N_15628);
nand U16348 (N_16348,N_15882,N_15744);
xnor U16349 (N_16349,N_15871,N_15646);
nor U16350 (N_16350,N_15907,N_15876);
nand U16351 (N_16351,N_15799,N_15647);
xor U16352 (N_16352,N_15617,N_15765);
or U16353 (N_16353,N_15947,N_15700);
nand U16354 (N_16354,N_15641,N_15803);
nor U16355 (N_16355,N_15859,N_15973);
nand U16356 (N_16356,N_15656,N_15708);
or U16357 (N_16357,N_15874,N_15728);
or U16358 (N_16358,N_15627,N_15642);
nor U16359 (N_16359,N_15861,N_15784);
xor U16360 (N_16360,N_15619,N_15971);
or U16361 (N_16361,N_15840,N_15943);
or U16362 (N_16362,N_15986,N_15905);
nor U16363 (N_16363,N_15880,N_15799);
and U16364 (N_16364,N_15838,N_15680);
nor U16365 (N_16365,N_15672,N_15940);
nor U16366 (N_16366,N_15870,N_15952);
nand U16367 (N_16367,N_15984,N_15838);
or U16368 (N_16368,N_15944,N_15686);
nand U16369 (N_16369,N_15909,N_15859);
and U16370 (N_16370,N_15985,N_15912);
nand U16371 (N_16371,N_15882,N_15769);
and U16372 (N_16372,N_15867,N_15738);
nor U16373 (N_16373,N_15961,N_15824);
nand U16374 (N_16374,N_15654,N_15752);
nor U16375 (N_16375,N_15907,N_15622);
xor U16376 (N_16376,N_15805,N_15790);
nand U16377 (N_16377,N_15680,N_15602);
xnor U16378 (N_16378,N_15997,N_15722);
xnor U16379 (N_16379,N_15947,N_15910);
xor U16380 (N_16380,N_15690,N_15956);
and U16381 (N_16381,N_15860,N_15917);
and U16382 (N_16382,N_15833,N_15809);
nand U16383 (N_16383,N_15617,N_15841);
nor U16384 (N_16384,N_15888,N_15762);
or U16385 (N_16385,N_15731,N_15806);
or U16386 (N_16386,N_15956,N_15993);
nor U16387 (N_16387,N_15642,N_15728);
xor U16388 (N_16388,N_15828,N_15618);
or U16389 (N_16389,N_15975,N_15716);
xnor U16390 (N_16390,N_15627,N_15746);
nand U16391 (N_16391,N_15906,N_15665);
nand U16392 (N_16392,N_15956,N_15759);
nand U16393 (N_16393,N_15930,N_15605);
and U16394 (N_16394,N_15696,N_15674);
xnor U16395 (N_16395,N_15941,N_15669);
and U16396 (N_16396,N_15705,N_15819);
nand U16397 (N_16397,N_15993,N_15613);
or U16398 (N_16398,N_15708,N_15864);
nor U16399 (N_16399,N_15800,N_15846);
xnor U16400 (N_16400,N_16109,N_16100);
xor U16401 (N_16401,N_16260,N_16286);
and U16402 (N_16402,N_16268,N_16381);
or U16403 (N_16403,N_16153,N_16399);
nor U16404 (N_16404,N_16246,N_16394);
nor U16405 (N_16405,N_16355,N_16353);
and U16406 (N_16406,N_16083,N_16138);
and U16407 (N_16407,N_16148,N_16347);
nand U16408 (N_16408,N_16054,N_16003);
and U16409 (N_16409,N_16267,N_16393);
xnor U16410 (N_16410,N_16330,N_16363);
or U16411 (N_16411,N_16318,N_16365);
and U16412 (N_16412,N_16266,N_16183);
nand U16413 (N_16413,N_16132,N_16019);
nand U16414 (N_16414,N_16004,N_16129);
nor U16415 (N_16415,N_16102,N_16050);
xnor U16416 (N_16416,N_16130,N_16325);
nor U16417 (N_16417,N_16263,N_16043);
xnor U16418 (N_16418,N_16396,N_16152);
xor U16419 (N_16419,N_16157,N_16141);
or U16420 (N_16420,N_16044,N_16150);
nor U16421 (N_16421,N_16240,N_16233);
and U16422 (N_16422,N_16234,N_16010);
xnor U16423 (N_16423,N_16339,N_16310);
nor U16424 (N_16424,N_16116,N_16271);
and U16425 (N_16425,N_16176,N_16344);
nor U16426 (N_16426,N_16211,N_16122);
nor U16427 (N_16427,N_16181,N_16162);
xnor U16428 (N_16428,N_16382,N_16217);
nor U16429 (N_16429,N_16345,N_16346);
xnor U16430 (N_16430,N_16289,N_16095);
nor U16431 (N_16431,N_16031,N_16232);
nand U16432 (N_16432,N_16080,N_16064);
and U16433 (N_16433,N_16287,N_16007);
and U16434 (N_16434,N_16320,N_16096);
nand U16435 (N_16435,N_16146,N_16250);
xor U16436 (N_16436,N_16302,N_16139);
xor U16437 (N_16437,N_16062,N_16072);
or U16438 (N_16438,N_16067,N_16155);
nor U16439 (N_16439,N_16312,N_16392);
or U16440 (N_16440,N_16262,N_16364);
and U16441 (N_16441,N_16055,N_16354);
xor U16442 (N_16442,N_16338,N_16305);
xor U16443 (N_16443,N_16342,N_16030);
nor U16444 (N_16444,N_16200,N_16202);
nand U16445 (N_16445,N_16060,N_16329);
and U16446 (N_16446,N_16280,N_16040);
or U16447 (N_16447,N_16229,N_16341);
xnor U16448 (N_16448,N_16015,N_16039);
nand U16449 (N_16449,N_16073,N_16105);
nand U16450 (N_16450,N_16035,N_16270);
nand U16451 (N_16451,N_16395,N_16056);
nand U16452 (N_16452,N_16236,N_16169);
nand U16453 (N_16453,N_16016,N_16121);
and U16454 (N_16454,N_16136,N_16158);
nor U16455 (N_16455,N_16391,N_16203);
nand U16456 (N_16456,N_16373,N_16154);
nand U16457 (N_16457,N_16235,N_16212);
xor U16458 (N_16458,N_16379,N_16282);
and U16459 (N_16459,N_16256,N_16206);
and U16460 (N_16460,N_16113,N_16265);
nand U16461 (N_16461,N_16065,N_16110);
nand U16462 (N_16462,N_16386,N_16023);
xor U16463 (N_16463,N_16241,N_16384);
nor U16464 (N_16464,N_16315,N_16316);
nand U16465 (N_16465,N_16002,N_16195);
nand U16466 (N_16466,N_16297,N_16193);
or U16467 (N_16467,N_16224,N_16168);
xor U16468 (N_16468,N_16245,N_16291);
and U16469 (N_16469,N_16127,N_16037);
xor U16470 (N_16470,N_16362,N_16008);
nor U16471 (N_16471,N_16009,N_16182);
nor U16472 (N_16472,N_16295,N_16149);
or U16473 (N_16473,N_16253,N_16128);
nand U16474 (N_16474,N_16348,N_16006);
nand U16475 (N_16475,N_16159,N_16198);
nor U16476 (N_16476,N_16140,N_16201);
nor U16477 (N_16477,N_16092,N_16349);
nor U16478 (N_16478,N_16078,N_16231);
xor U16479 (N_16479,N_16225,N_16052);
nand U16480 (N_16480,N_16205,N_16179);
or U16481 (N_16481,N_16356,N_16051);
and U16482 (N_16482,N_16022,N_16307);
xnor U16483 (N_16483,N_16228,N_16021);
xnor U16484 (N_16484,N_16081,N_16252);
xor U16485 (N_16485,N_16048,N_16388);
nand U16486 (N_16486,N_16374,N_16324);
and U16487 (N_16487,N_16368,N_16336);
nor U16488 (N_16488,N_16046,N_16099);
or U16489 (N_16489,N_16226,N_16276);
or U16490 (N_16490,N_16375,N_16389);
nand U16491 (N_16491,N_16207,N_16313);
xor U16492 (N_16492,N_16190,N_16020);
or U16493 (N_16493,N_16156,N_16126);
nor U16494 (N_16494,N_16334,N_16075);
or U16495 (N_16495,N_16086,N_16071);
and U16496 (N_16496,N_16213,N_16170);
and U16497 (N_16497,N_16074,N_16053);
or U16498 (N_16498,N_16028,N_16251);
or U16499 (N_16499,N_16208,N_16185);
nor U16500 (N_16500,N_16036,N_16358);
nor U16501 (N_16501,N_16269,N_16311);
nor U16502 (N_16502,N_16077,N_16088);
nor U16503 (N_16503,N_16013,N_16104);
and U16504 (N_16504,N_16283,N_16264);
xnor U16505 (N_16505,N_16167,N_16027);
xnor U16506 (N_16506,N_16084,N_16292);
and U16507 (N_16507,N_16000,N_16322);
nand U16508 (N_16508,N_16274,N_16131);
nand U16509 (N_16509,N_16238,N_16145);
xnor U16510 (N_16510,N_16390,N_16108);
or U16511 (N_16511,N_16220,N_16103);
nand U16512 (N_16512,N_16045,N_16335);
nor U16513 (N_16513,N_16175,N_16372);
or U16514 (N_16514,N_16079,N_16314);
and U16515 (N_16515,N_16112,N_16242);
nor U16516 (N_16516,N_16161,N_16069);
or U16517 (N_16517,N_16387,N_16106);
or U16518 (N_16518,N_16279,N_16143);
or U16519 (N_16519,N_16180,N_16214);
or U16520 (N_16520,N_16369,N_16142);
nor U16521 (N_16521,N_16293,N_16360);
and U16522 (N_16522,N_16350,N_16172);
or U16523 (N_16523,N_16398,N_16397);
xnor U16524 (N_16524,N_16239,N_16210);
or U16525 (N_16525,N_16063,N_16118);
xor U16526 (N_16526,N_16284,N_16194);
nor U16527 (N_16527,N_16093,N_16378);
nand U16528 (N_16528,N_16340,N_16101);
nor U16529 (N_16529,N_16133,N_16012);
xor U16530 (N_16530,N_16290,N_16371);
xor U16531 (N_16531,N_16370,N_16321);
and U16532 (N_16532,N_16304,N_16144);
or U16533 (N_16533,N_16090,N_16191);
nor U16534 (N_16534,N_16041,N_16296);
or U16535 (N_16535,N_16018,N_16385);
or U16536 (N_16536,N_16223,N_16085);
nand U16537 (N_16537,N_16024,N_16189);
nor U16538 (N_16538,N_16107,N_16124);
or U16539 (N_16539,N_16357,N_16165);
xnor U16540 (N_16540,N_16332,N_16288);
or U16541 (N_16541,N_16337,N_16058);
and U16542 (N_16542,N_16380,N_16306);
nand U16543 (N_16543,N_16331,N_16204);
xnor U16544 (N_16544,N_16299,N_16328);
xor U16545 (N_16545,N_16237,N_16171);
and U16546 (N_16546,N_16301,N_16326);
and U16547 (N_16547,N_16076,N_16070);
nand U16548 (N_16548,N_16091,N_16367);
or U16549 (N_16549,N_16351,N_16285);
nor U16550 (N_16550,N_16017,N_16177);
and U16551 (N_16551,N_16068,N_16300);
or U16552 (N_16552,N_16359,N_16029);
xor U16553 (N_16553,N_16082,N_16273);
and U16554 (N_16554,N_16218,N_16151);
nand U16555 (N_16555,N_16192,N_16244);
and U16556 (N_16556,N_16343,N_16255);
xnor U16557 (N_16557,N_16281,N_16174);
or U16558 (N_16558,N_16294,N_16137);
nand U16559 (N_16559,N_16303,N_16057);
nor U16560 (N_16560,N_16033,N_16261);
and U16561 (N_16561,N_16366,N_16376);
and U16562 (N_16562,N_16038,N_16049);
xor U16563 (N_16563,N_16184,N_16014);
xnor U16564 (N_16564,N_16361,N_16219);
xnor U16565 (N_16565,N_16216,N_16319);
or U16566 (N_16566,N_16333,N_16249);
nand U16567 (N_16567,N_16115,N_16209);
nor U16568 (N_16568,N_16034,N_16125);
and U16569 (N_16569,N_16199,N_16123);
nand U16570 (N_16570,N_16259,N_16222);
and U16571 (N_16571,N_16188,N_16026);
or U16572 (N_16572,N_16248,N_16173);
xnor U16573 (N_16573,N_16327,N_16377);
nand U16574 (N_16574,N_16215,N_16098);
or U16575 (N_16575,N_16196,N_16011);
nand U16576 (N_16576,N_16061,N_16277);
xor U16577 (N_16577,N_16097,N_16001);
nand U16578 (N_16578,N_16164,N_16230);
or U16579 (N_16579,N_16042,N_16186);
nor U16580 (N_16580,N_16254,N_16120);
xnor U16581 (N_16581,N_16114,N_16094);
nand U16582 (N_16582,N_16272,N_16160);
xnor U16583 (N_16583,N_16166,N_16089);
nand U16584 (N_16584,N_16323,N_16117);
xnor U16585 (N_16585,N_16147,N_16317);
nand U16586 (N_16586,N_16352,N_16298);
and U16587 (N_16587,N_16163,N_16221);
xor U16588 (N_16588,N_16257,N_16111);
xor U16589 (N_16589,N_16025,N_16178);
and U16590 (N_16590,N_16275,N_16308);
and U16591 (N_16591,N_16087,N_16243);
and U16592 (N_16592,N_16135,N_16066);
nand U16593 (N_16593,N_16119,N_16032);
or U16594 (N_16594,N_16383,N_16258);
nand U16595 (N_16595,N_16309,N_16059);
nand U16596 (N_16596,N_16187,N_16197);
and U16597 (N_16597,N_16247,N_16134);
xor U16598 (N_16598,N_16227,N_16047);
nor U16599 (N_16599,N_16278,N_16005);
xor U16600 (N_16600,N_16240,N_16172);
and U16601 (N_16601,N_16162,N_16019);
xor U16602 (N_16602,N_16076,N_16025);
or U16603 (N_16603,N_16340,N_16162);
nand U16604 (N_16604,N_16289,N_16363);
and U16605 (N_16605,N_16235,N_16154);
and U16606 (N_16606,N_16022,N_16321);
nand U16607 (N_16607,N_16264,N_16164);
and U16608 (N_16608,N_16261,N_16250);
xnor U16609 (N_16609,N_16390,N_16260);
or U16610 (N_16610,N_16379,N_16303);
and U16611 (N_16611,N_16159,N_16067);
nand U16612 (N_16612,N_16395,N_16274);
or U16613 (N_16613,N_16003,N_16205);
nand U16614 (N_16614,N_16351,N_16030);
or U16615 (N_16615,N_16357,N_16317);
and U16616 (N_16616,N_16062,N_16342);
or U16617 (N_16617,N_16338,N_16201);
nand U16618 (N_16618,N_16068,N_16327);
nor U16619 (N_16619,N_16199,N_16313);
xor U16620 (N_16620,N_16101,N_16099);
xnor U16621 (N_16621,N_16099,N_16189);
nand U16622 (N_16622,N_16139,N_16056);
and U16623 (N_16623,N_16325,N_16213);
nand U16624 (N_16624,N_16081,N_16362);
nor U16625 (N_16625,N_16353,N_16028);
xnor U16626 (N_16626,N_16022,N_16194);
xor U16627 (N_16627,N_16186,N_16313);
or U16628 (N_16628,N_16338,N_16053);
nand U16629 (N_16629,N_16081,N_16157);
nand U16630 (N_16630,N_16322,N_16097);
or U16631 (N_16631,N_16381,N_16009);
xnor U16632 (N_16632,N_16286,N_16284);
xor U16633 (N_16633,N_16270,N_16241);
and U16634 (N_16634,N_16175,N_16387);
xnor U16635 (N_16635,N_16322,N_16234);
nor U16636 (N_16636,N_16190,N_16104);
and U16637 (N_16637,N_16050,N_16145);
nor U16638 (N_16638,N_16350,N_16217);
or U16639 (N_16639,N_16133,N_16109);
nand U16640 (N_16640,N_16006,N_16101);
nand U16641 (N_16641,N_16036,N_16325);
or U16642 (N_16642,N_16351,N_16271);
nor U16643 (N_16643,N_16380,N_16368);
nand U16644 (N_16644,N_16151,N_16233);
nor U16645 (N_16645,N_16350,N_16046);
nand U16646 (N_16646,N_16118,N_16201);
nor U16647 (N_16647,N_16358,N_16360);
and U16648 (N_16648,N_16317,N_16383);
nor U16649 (N_16649,N_16127,N_16206);
xor U16650 (N_16650,N_16022,N_16191);
nand U16651 (N_16651,N_16306,N_16299);
and U16652 (N_16652,N_16342,N_16160);
and U16653 (N_16653,N_16374,N_16210);
xor U16654 (N_16654,N_16044,N_16002);
xnor U16655 (N_16655,N_16239,N_16174);
or U16656 (N_16656,N_16237,N_16072);
nor U16657 (N_16657,N_16368,N_16334);
nand U16658 (N_16658,N_16369,N_16389);
nor U16659 (N_16659,N_16212,N_16322);
or U16660 (N_16660,N_16321,N_16123);
or U16661 (N_16661,N_16027,N_16377);
or U16662 (N_16662,N_16136,N_16038);
and U16663 (N_16663,N_16257,N_16201);
xor U16664 (N_16664,N_16199,N_16336);
or U16665 (N_16665,N_16231,N_16378);
or U16666 (N_16666,N_16123,N_16105);
nor U16667 (N_16667,N_16157,N_16125);
nand U16668 (N_16668,N_16114,N_16386);
or U16669 (N_16669,N_16126,N_16200);
nand U16670 (N_16670,N_16195,N_16153);
xnor U16671 (N_16671,N_16250,N_16218);
nor U16672 (N_16672,N_16209,N_16350);
or U16673 (N_16673,N_16284,N_16361);
xor U16674 (N_16674,N_16030,N_16015);
nor U16675 (N_16675,N_16348,N_16242);
nand U16676 (N_16676,N_16205,N_16001);
xnor U16677 (N_16677,N_16117,N_16009);
and U16678 (N_16678,N_16209,N_16280);
nand U16679 (N_16679,N_16330,N_16276);
xnor U16680 (N_16680,N_16207,N_16389);
or U16681 (N_16681,N_16098,N_16219);
xnor U16682 (N_16682,N_16223,N_16371);
nand U16683 (N_16683,N_16197,N_16337);
or U16684 (N_16684,N_16334,N_16190);
xnor U16685 (N_16685,N_16039,N_16140);
nor U16686 (N_16686,N_16320,N_16281);
and U16687 (N_16687,N_16361,N_16029);
xor U16688 (N_16688,N_16201,N_16048);
and U16689 (N_16689,N_16001,N_16389);
or U16690 (N_16690,N_16343,N_16120);
nor U16691 (N_16691,N_16244,N_16124);
and U16692 (N_16692,N_16237,N_16061);
and U16693 (N_16693,N_16149,N_16128);
nor U16694 (N_16694,N_16281,N_16289);
or U16695 (N_16695,N_16109,N_16210);
and U16696 (N_16696,N_16003,N_16178);
nor U16697 (N_16697,N_16026,N_16123);
nand U16698 (N_16698,N_16341,N_16328);
and U16699 (N_16699,N_16041,N_16317);
and U16700 (N_16700,N_16182,N_16343);
or U16701 (N_16701,N_16102,N_16318);
xnor U16702 (N_16702,N_16260,N_16220);
or U16703 (N_16703,N_16377,N_16114);
nand U16704 (N_16704,N_16030,N_16098);
and U16705 (N_16705,N_16319,N_16181);
nand U16706 (N_16706,N_16215,N_16141);
and U16707 (N_16707,N_16143,N_16310);
nor U16708 (N_16708,N_16050,N_16185);
xor U16709 (N_16709,N_16215,N_16132);
nor U16710 (N_16710,N_16297,N_16359);
and U16711 (N_16711,N_16390,N_16224);
and U16712 (N_16712,N_16066,N_16027);
or U16713 (N_16713,N_16272,N_16195);
xor U16714 (N_16714,N_16182,N_16006);
nand U16715 (N_16715,N_16195,N_16030);
nand U16716 (N_16716,N_16272,N_16371);
and U16717 (N_16717,N_16286,N_16230);
or U16718 (N_16718,N_16278,N_16048);
nor U16719 (N_16719,N_16294,N_16277);
xor U16720 (N_16720,N_16219,N_16008);
and U16721 (N_16721,N_16260,N_16098);
xor U16722 (N_16722,N_16032,N_16285);
nor U16723 (N_16723,N_16172,N_16131);
nor U16724 (N_16724,N_16030,N_16211);
nand U16725 (N_16725,N_16069,N_16212);
and U16726 (N_16726,N_16136,N_16140);
or U16727 (N_16727,N_16273,N_16336);
and U16728 (N_16728,N_16299,N_16359);
xor U16729 (N_16729,N_16064,N_16249);
nand U16730 (N_16730,N_16179,N_16165);
and U16731 (N_16731,N_16282,N_16081);
nand U16732 (N_16732,N_16110,N_16211);
and U16733 (N_16733,N_16348,N_16249);
or U16734 (N_16734,N_16329,N_16068);
nand U16735 (N_16735,N_16245,N_16238);
and U16736 (N_16736,N_16132,N_16082);
and U16737 (N_16737,N_16155,N_16236);
nand U16738 (N_16738,N_16218,N_16280);
or U16739 (N_16739,N_16079,N_16075);
and U16740 (N_16740,N_16023,N_16223);
and U16741 (N_16741,N_16024,N_16265);
or U16742 (N_16742,N_16315,N_16243);
nand U16743 (N_16743,N_16137,N_16141);
nor U16744 (N_16744,N_16056,N_16264);
nand U16745 (N_16745,N_16083,N_16359);
xnor U16746 (N_16746,N_16123,N_16084);
nor U16747 (N_16747,N_16047,N_16201);
nand U16748 (N_16748,N_16327,N_16390);
and U16749 (N_16749,N_16294,N_16319);
nor U16750 (N_16750,N_16360,N_16357);
xnor U16751 (N_16751,N_16222,N_16369);
xnor U16752 (N_16752,N_16233,N_16131);
xor U16753 (N_16753,N_16398,N_16063);
or U16754 (N_16754,N_16114,N_16005);
nand U16755 (N_16755,N_16348,N_16191);
nor U16756 (N_16756,N_16181,N_16254);
nor U16757 (N_16757,N_16128,N_16115);
nor U16758 (N_16758,N_16291,N_16167);
or U16759 (N_16759,N_16251,N_16310);
nor U16760 (N_16760,N_16078,N_16375);
nand U16761 (N_16761,N_16185,N_16212);
xor U16762 (N_16762,N_16284,N_16002);
xor U16763 (N_16763,N_16329,N_16067);
nand U16764 (N_16764,N_16246,N_16181);
nor U16765 (N_16765,N_16103,N_16379);
nor U16766 (N_16766,N_16387,N_16261);
and U16767 (N_16767,N_16134,N_16024);
nand U16768 (N_16768,N_16118,N_16130);
nor U16769 (N_16769,N_16344,N_16234);
or U16770 (N_16770,N_16172,N_16305);
nor U16771 (N_16771,N_16251,N_16299);
nor U16772 (N_16772,N_16237,N_16295);
or U16773 (N_16773,N_16299,N_16090);
nor U16774 (N_16774,N_16102,N_16042);
nand U16775 (N_16775,N_16275,N_16361);
and U16776 (N_16776,N_16045,N_16155);
nor U16777 (N_16777,N_16029,N_16286);
and U16778 (N_16778,N_16333,N_16279);
and U16779 (N_16779,N_16061,N_16111);
xnor U16780 (N_16780,N_16208,N_16023);
and U16781 (N_16781,N_16351,N_16031);
or U16782 (N_16782,N_16267,N_16273);
xnor U16783 (N_16783,N_16092,N_16318);
nand U16784 (N_16784,N_16193,N_16095);
nand U16785 (N_16785,N_16389,N_16152);
and U16786 (N_16786,N_16039,N_16001);
and U16787 (N_16787,N_16191,N_16197);
nand U16788 (N_16788,N_16258,N_16032);
and U16789 (N_16789,N_16297,N_16264);
nor U16790 (N_16790,N_16385,N_16245);
xnor U16791 (N_16791,N_16074,N_16066);
nand U16792 (N_16792,N_16150,N_16298);
xor U16793 (N_16793,N_16311,N_16342);
or U16794 (N_16794,N_16202,N_16353);
nor U16795 (N_16795,N_16207,N_16325);
or U16796 (N_16796,N_16054,N_16181);
and U16797 (N_16797,N_16196,N_16164);
nor U16798 (N_16798,N_16029,N_16291);
xor U16799 (N_16799,N_16197,N_16032);
and U16800 (N_16800,N_16736,N_16633);
and U16801 (N_16801,N_16550,N_16554);
or U16802 (N_16802,N_16426,N_16651);
or U16803 (N_16803,N_16653,N_16737);
nand U16804 (N_16804,N_16549,N_16535);
xor U16805 (N_16805,N_16476,N_16412);
xor U16806 (N_16806,N_16501,N_16788);
nand U16807 (N_16807,N_16747,N_16526);
xnor U16808 (N_16808,N_16656,N_16486);
nand U16809 (N_16809,N_16527,N_16536);
or U16810 (N_16810,N_16512,N_16415);
and U16811 (N_16811,N_16459,N_16607);
xnor U16812 (N_16812,N_16752,N_16548);
nor U16813 (N_16813,N_16566,N_16629);
or U16814 (N_16814,N_16445,N_16614);
xor U16815 (N_16815,N_16406,N_16465);
xor U16816 (N_16816,N_16402,N_16751);
nand U16817 (N_16817,N_16538,N_16487);
or U16818 (N_16818,N_16668,N_16516);
nand U16819 (N_16819,N_16420,N_16617);
nand U16820 (N_16820,N_16759,N_16652);
nand U16821 (N_16821,N_16506,N_16715);
or U16822 (N_16822,N_16645,N_16589);
and U16823 (N_16823,N_16562,N_16563);
xor U16824 (N_16824,N_16489,N_16432);
or U16825 (N_16825,N_16770,N_16636);
xor U16826 (N_16826,N_16711,N_16613);
nor U16827 (N_16827,N_16655,N_16494);
and U16828 (N_16828,N_16525,N_16577);
nor U16829 (N_16829,N_16482,N_16514);
xor U16830 (N_16830,N_16599,N_16769);
xnor U16831 (N_16831,N_16582,N_16587);
nor U16832 (N_16832,N_16673,N_16541);
nor U16833 (N_16833,N_16513,N_16734);
xnor U16834 (N_16834,N_16620,N_16574);
nand U16835 (N_16835,N_16739,N_16778);
nand U16836 (N_16836,N_16744,N_16775);
nor U16837 (N_16837,N_16517,N_16542);
nand U16838 (N_16838,N_16404,N_16484);
nand U16839 (N_16839,N_16703,N_16621);
nand U16840 (N_16840,N_16416,N_16661);
nand U16841 (N_16841,N_16546,N_16596);
or U16842 (N_16842,N_16576,N_16697);
and U16843 (N_16843,N_16746,N_16608);
or U16844 (N_16844,N_16706,N_16594);
nor U16845 (N_16845,N_16559,N_16735);
xnor U16846 (N_16846,N_16713,N_16444);
or U16847 (N_16847,N_16678,N_16748);
or U16848 (N_16848,N_16741,N_16648);
nor U16849 (N_16849,N_16558,N_16709);
xnor U16850 (N_16850,N_16463,N_16449);
or U16851 (N_16851,N_16570,N_16635);
and U16852 (N_16852,N_16509,N_16529);
xnor U16853 (N_16853,N_16792,N_16772);
and U16854 (N_16854,N_16485,N_16531);
nand U16855 (N_16855,N_16627,N_16555);
nand U16856 (N_16856,N_16469,N_16436);
nor U16857 (N_16857,N_16685,N_16413);
and U16858 (N_16858,N_16600,N_16545);
nand U16859 (N_16859,N_16493,N_16647);
nor U16860 (N_16860,N_16722,N_16676);
nor U16861 (N_16861,N_16428,N_16716);
nand U16862 (N_16862,N_16616,N_16575);
xnor U16863 (N_16863,N_16679,N_16409);
and U16864 (N_16864,N_16433,N_16776);
xor U16865 (N_16865,N_16714,N_16528);
xor U16866 (N_16866,N_16782,N_16691);
nand U16867 (N_16867,N_16755,N_16461);
or U16868 (N_16868,N_16464,N_16448);
nand U16869 (N_16869,N_16625,N_16523);
nor U16870 (N_16870,N_16583,N_16641);
and U16871 (N_16871,N_16460,N_16794);
and U16872 (N_16872,N_16768,N_16662);
nand U16873 (N_16873,N_16692,N_16701);
xnor U16874 (N_16874,N_16508,N_16667);
and U16875 (N_16875,N_16753,N_16597);
or U16876 (N_16876,N_16586,N_16507);
nand U16877 (N_16877,N_16441,N_16694);
and U16878 (N_16878,N_16533,N_16591);
xnor U16879 (N_16879,N_16684,N_16455);
or U16880 (N_16880,N_16786,N_16474);
or U16881 (N_16881,N_16552,N_16442);
xnor U16882 (N_16882,N_16756,N_16758);
nand U16883 (N_16883,N_16793,N_16400);
nand U16884 (N_16884,N_16723,N_16665);
and U16885 (N_16885,N_16717,N_16405);
or U16886 (N_16886,N_16689,N_16708);
and U16887 (N_16887,N_16403,N_16573);
nand U16888 (N_16888,N_16423,N_16468);
xnor U16889 (N_16889,N_16624,N_16521);
nor U16890 (N_16890,N_16543,N_16443);
and U16891 (N_16891,N_16547,N_16557);
and U16892 (N_16892,N_16646,N_16712);
or U16893 (N_16893,N_16785,N_16481);
nor U16894 (N_16894,N_16478,N_16659);
xor U16895 (N_16895,N_16677,N_16431);
or U16896 (N_16896,N_16740,N_16610);
nand U16897 (N_16897,N_16532,N_16503);
nand U16898 (N_16898,N_16790,N_16687);
nor U16899 (N_16899,N_16688,N_16495);
nand U16900 (N_16900,N_16649,N_16754);
xnor U16901 (N_16901,N_16773,N_16681);
or U16902 (N_16902,N_16675,N_16450);
and U16903 (N_16903,N_16553,N_16766);
xor U16904 (N_16904,N_16795,N_16686);
nor U16905 (N_16905,N_16654,N_16605);
xnor U16906 (N_16906,N_16779,N_16764);
nand U16907 (N_16907,N_16519,N_16467);
xnor U16908 (N_16908,N_16567,N_16473);
xor U16909 (N_16909,N_16721,N_16693);
or U16910 (N_16910,N_16470,N_16727);
nor U16911 (N_16911,N_16435,N_16500);
or U16912 (N_16912,N_16551,N_16699);
xnor U16913 (N_16913,N_16743,N_16799);
nor U16914 (N_16914,N_16569,N_16611);
nor U16915 (N_16915,N_16437,N_16781);
or U16916 (N_16916,N_16411,N_16628);
nand U16917 (N_16917,N_16774,N_16477);
or U16918 (N_16918,N_16571,N_16642);
xnor U16919 (N_16919,N_16650,N_16408);
and U16920 (N_16920,N_16479,N_16632);
and U16921 (N_16921,N_16578,N_16522);
nand U16922 (N_16922,N_16490,N_16660);
and U16923 (N_16923,N_16695,N_16592);
xnor U16924 (N_16924,N_16762,N_16466);
xor U16925 (N_16925,N_16726,N_16622);
xnor U16926 (N_16926,N_16612,N_16540);
and U16927 (N_16927,N_16705,N_16637);
nor U16928 (N_16928,N_16704,N_16520);
and U16929 (N_16929,N_16707,N_16417);
or U16930 (N_16930,N_16742,N_16492);
and U16931 (N_16931,N_16798,N_16498);
or U16932 (N_16932,N_16789,N_16418);
nand U16933 (N_16933,N_16601,N_16718);
or U16934 (N_16934,N_16784,N_16603);
nor U16935 (N_16935,N_16407,N_16457);
nor U16936 (N_16936,N_16446,N_16401);
xnor U16937 (N_16937,N_16453,N_16452);
or U16938 (N_16938,N_16634,N_16499);
and U16939 (N_16939,N_16488,N_16422);
xor U16940 (N_16940,N_16439,N_16657);
nand U16941 (N_16941,N_16618,N_16585);
xor U16942 (N_16942,N_16698,N_16419);
nor U16943 (N_16943,N_16414,N_16638);
or U16944 (N_16944,N_16623,N_16609);
nor U16945 (N_16945,N_16757,N_16644);
nand U16946 (N_16946,N_16447,N_16593);
nand U16947 (N_16947,N_16424,N_16524);
nor U16948 (N_16948,N_16619,N_16510);
xor U16949 (N_16949,N_16544,N_16456);
nand U16950 (N_16950,N_16777,N_16666);
nand U16951 (N_16951,N_16561,N_16696);
and U16952 (N_16952,N_16710,N_16458);
and U16953 (N_16953,N_16750,N_16738);
xor U16954 (N_16954,N_16434,N_16671);
nand U16955 (N_16955,N_16680,N_16511);
xor U16956 (N_16956,N_16670,N_16530);
nand U16957 (N_16957,N_16471,N_16475);
and U16958 (N_16958,N_16763,N_16630);
or U16959 (N_16959,N_16472,N_16663);
or U16960 (N_16960,N_16796,N_16643);
and U16961 (N_16961,N_16640,N_16783);
nand U16962 (N_16962,N_16658,N_16719);
and U16963 (N_16963,N_16579,N_16539);
xor U16964 (N_16964,N_16556,N_16568);
xor U16965 (N_16965,N_16745,N_16462);
nor U16966 (N_16966,N_16502,N_16560);
nand U16967 (N_16967,N_16765,N_16421);
nor U16968 (N_16968,N_16787,N_16732);
or U16969 (N_16969,N_16606,N_16454);
nor U16970 (N_16970,N_16631,N_16505);
xnor U16971 (N_16971,N_16410,N_16598);
nand U16972 (N_16972,N_16565,N_16491);
nand U16973 (N_16973,N_16504,N_16590);
nor U16974 (N_16974,N_16728,N_16720);
nor U16975 (N_16975,N_16581,N_16672);
or U16976 (N_16976,N_16564,N_16690);
nand U16977 (N_16977,N_16664,N_16572);
and U16978 (N_16978,N_16749,N_16682);
nor U16979 (N_16979,N_16430,N_16761);
and U16980 (N_16980,N_16604,N_16440);
or U16981 (N_16981,N_16674,N_16669);
and U16982 (N_16982,N_16427,N_16760);
and U16983 (N_16983,N_16683,N_16700);
and U16984 (N_16984,N_16730,N_16731);
xnor U16985 (N_16985,N_16725,N_16639);
and U16986 (N_16986,N_16534,N_16580);
nand U16987 (N_16987,N_16429,N_16724);
nor U16988 (N_16988,N_16797,N_16425);
and U16989 (N_16989,N_16588,N_16496);
xnor U16990 (N_16990,N_16497,N_16780);
or U16991 (N_16991,N_16702,N_16733);
and U16992 (N_16992,N_16438,N_16451);
xnor U16993 (N_16993,N_16602,N_16626);
nor U16994 (N_16994,N_16480,N_16595);
or U16995 (N_16995,N_16615,N_16483);
xnor U16996 (N_16996,N_16767,N_16515);
nor U16997 (N_16997,N_16771,N_16729);
and U16998 (N_16998,N_16537,N_16584);
or U16999 (N_16999,N_16518,N_16791);
or U17000 (N_17000,N_16618,N_16608);
or U17001 (N_17001,N_16522,N_16773);
and U17002 (N_17002,N_16580,N_16740);
xnor U17003 (N_17003,N_16737,N_16703);
xor U17004 (N_17004,N_16649,N_16436);
xnor U17005 (N_17005,N_16527,N_16443);
or U17006 (N_17006,N_16427,N_16661);
nand U17007 (N_17007,N_16515,N_16544);
or U17008 (N_17008,N_16572,N_16508);
nand U17009 (N_17009,N_16456,N_16701);
and U17010 (N_17010,N_16713,N_16597);
nor U17011 (N_17011,N_16507,N_16727);
or U17012 (N_17012,N_16668,N_16666);
and U17013 (N_17013,N_16519,N_16708);
xnor U17014 (N_17014,N_16454,N_16661);
nand U17015 (N_17015,N_16619,N_16463);
and U17016 (N_17016,N_16443,N_16693);
xor U17017 (N_17017,N_16722,N_16493);
nand U17018 (N_17018,N_16789,N_16700);
and U17019 (N_17019,N_16450,N_16589);
nor U17020 (N_17020,N_16572,N_16703);
and U17021 (N_17021,N_16678,N_16636);
nand U17022 (N_17022,N_16781,N_16796);
and U17023 (N_17023,N_16473,N_16667);
xor U17024 (N_17024,N_16474,N_16484);
nand U17025 (N_17025,N_16621,N_16541);
or U17026 (N_17026,N_16589,N_16551);
nor U17027 (N_17027,N_16789,N_16571);
nor U17028 (N_17028,N_16797,N_16729);
nand U17029 (N_17029,N_16684,N_16538);
and U17030 (N_17030,N_16510,N_16677);
or U17031 (N_17031,N_16779,N_16780);
xor U17032 (N_17032,N_16760,N_16498);
xor U17033 (N_17033,N_16571,N_16667);
xor U17034 (N_17034,N_16694,N_16635);
nor U17035 (N_17035,N_16710,N_16688);
nor U17036 (N_17036,N_16535,N_16702);
nor U17037 (N_17037,N_16605,N_16425);
and U17038 (N_17038,N_16739,N_16761);
and U17039 (N_17039,N_16412,N_16614);
or U17040 (N_17040,N_16746,N_16497);
xnor U17041 (N_17041,N_16554,N_16504);
nor U17042 (N_17042,N_16774,N_16666);
nand U17043 (N_17043,N_16670,N_16710);
nor U17044 (N_17044,N_16551,N_16417);
or U17045 (N_17045,N_16695,N_16529);
and U17046 (N_17046,N_16621,N_16432);
or U17047 (N_17047,N_16514,N_16555);
nand U17048 (N_17048,N_16522,N_16609);
and U17049 (N_17049,N_16400,N_16531);
nand U17050 (N_17050,N_16666,N_16677);
or U17051 (N_17051,N_16669,N_16730);
and U17052 (N_17052,N_16769,N_16406);
xnor U17053 (N_17053,N_16765,N_16506);
and U17054 (N_17054,N_16506,N_16787);
nor U17055 (N_17055,N_16684,N_16667);
and U17056 (N_17056,N_16767,N_16783);
and U17057 (N_17057,N_16619,N_16492);
nand U17058 (N_17058,N_16769,N_16647);
or U17059 (N_17059,N_16491,N_16618);
nand U17060 (N_17060,N_16721,N_16491);
or U17061 (N_17061,N_16704,N_16535);
or U17062 (N_17062,N_16408,N_16506);
or U17063 (N_17063,N_16438,N_16409);
nor U17064 (N_17064,N_16518,N_16618);
nand U17065 (N_17065,N_16508,N_16540);
or U17066 (N_17066,N_16725,N_16470);
xor U17067 (N_17067,N_16579,N_16543);
nor U17068 (N_17068,N_16778,N_16538);
and U17069 (N_17069,N_16431,N_16620);
nand U17070 (N_17070,N_16769,N_16680);
xor U17071 (N_17071,N_16720,N_16571);
or U17072 (N_17072,N_16632,N_16414);
nor U17073 (N_17073,N_16409,N_16510);
xnor U17074 (N_17074,N_16635,N_16783);
nand U17075 (N_17075,N_16791,N_16431);
or U17076 (N_17076,N_16710,N_16778);
xor U17077 (N_17077,N_16711,N_16703);
xor U17078 (N_17078,N_16724,N_16646);
or U17079 (N_17079,N_16763,N_16619);
or U17080 (N_17080,N_16455,N_16490);
and U17081 (N_17081,N_16566,N_16725);
xor U17082 (N_17082,N_16579,N_16701);
or U17083 (N_17083,N_16532,N_16633);
nand U17084 (N_17084,N_16639,N_16719);
or U17085 (N_17085,N_16606,N_16735);
and U17086 (N_17086,N_16660,N_16514);
nand U17087 (N_17087,N_16612,N_16692);
or U17088 (N_17088,N_16546,N_16482);
xor U17089 (N_17089,N_16504,N_16719);
or U17090 (N_17090,N_16603,N_16477);
xnor U17091 (N_17091,N_16646,N_16615);
nand U17092 (N_17092,N_16444,N_16403);
and U17093 (N_17093,N_16710,N_16457);
nand U17094 (N_17094,N_16792,N_16746);
and U17095 (N_17095,N_16772,N_16497);
nand U17096 (N_17096,N_16790,N_16780);
or U17097 (N_17097,N_16520,N_16504);
and U17098 (N_17098,N_16567,N_16759);
xor U17099 (N_17099,N_16496,N_16614);
nand U17100 (N_17100,N_16663,N_16708);
and U17101 (N_17101,N_16563,N_16632);
xnor U17102 (N_17102,N_16704,N_16506);
nor U17103 (N_17103,N_16433,N_16520);
nor U17104 (N_17104,N_16441,N_16703);
xor U17105 (N_17105,N_16676,N_16423);
nor U17106 (N_17106,N_16423,N_16437);
xnor U17107 (N_17107,N_16677,N_16683);
xor U17108 (N_17108,N_16467,N_16472);
or U17109 (N_17109,N_16462,N_16568);
xnor U17110 (N_17110,N_16635,N_16437);
or U17111 (N_17111,N_16663,N_16478);
and U17112 (N_17112,N_16417,N_16592);
xnor U17113 (N_17113,N_16653,N_16721);
nor U17114 (N_17114,N_16562,N_16576);
or U17115 (N_17115,N_16431,N_16511);
or U17116 (N_17116,N_16698,N_16771);
xnor U17117 (N_17117,N_16778,N_16760);
xor U17118 (N_17118,N_16587,N_16444);
nor U17119 (N_17119,N_16431,N_16764);
nor U17120 (N_17120,N_16637,N_16426);
nand U17121 (N_17121,N_16750,N_16780);
xnor U17122 (N_17122,N_16663,N_16491);
or U17123 (N_17123,N_16479,N_16721);
or U17124 (N_17124,N_16460,N_16547);
nor U17125 (N_17125,N_16551,N_16630);
xor U17126 (N_17126,N_16750,N_16402);
xnor U17127 (N_17127,N_16519,N_16673);
and U17128 (N_17128,N_16552,N_16657);
or U17129 (N_17129,N_16457,N_16617);
xnor U17130 (N_17130,N_16427,N_16630);
or U17131 (N_17131,N_16570,N_16474);
nor U17132 (N_17132,N_16494,N_16732);
and U17133 (N_17133,N_16757,N_16503);
nor U17134 (N_17134,N_16658,N_16757);
xnor U17135 (N_17135,N_16557,N_16459);
or U17136 (N_17136,N_16517,N_16699);
xnor U17137 (N_17137,N_16673,N_16626);
and U17138 (N_17138,N_16771,N_16476);
or U17139 (N_17139,N_16777,N_16450);
or U17140 (N_17140,N_16768,N_16640);
nor U17141 (N_17141,N_16653,N_16644);
and U17142 (N_17142,N_16416,N_16766);
or U17143 (N_17143,N_16421,N_16472);
and U17144 (N_17144,N_16786,N_16581);
and U17145 (N_17145,N_16714,N_16558);
nor U17146 (N_17146,N_16781,N_16692);
and U17147 (N_17147,N_16749,N_16407);
and U17148 (N_17148,N_16449,N_16466);
nor U17149 (N_17149,N_16741,N_16454);
and U17150 (N_17150,N_16427,N_16446);
nor U17151 (N_17151,N_16648,N_16690);
nor U17152 (N_17152,N_16498,N_16744);
and U17153 (N_17153,N_16593,N_16432);
nand U17154 (N_17154,N_16756,N_16474);
or U17155 (N_17155,N_16621,N_16504);
nor U17156 (N_17156,N_16574,N_16731);
nor U17157 (N_17157,N_16424,N_16647);
or U17158 (N_17158,N_16476,N_16656);
xor U17159 (N_17159,N_16604,N_16692);
or U17160 (N_17160,N_16794,N_16432);
nand U17161 (N_17161,N_16585,N_16656);
xor U17162 (N_17162,N_16503,N_16590);
xor U17163 (N_17163,N_16720,N_16451);
or U17164 (N_17164,N_16428,N_16433);
and U17165 (N_17165,N_16637,N_16679);
and U17166 (N_17166,N_16506,N_16627);
nand U17167 (N_17167,N_16450,N_16503);
or U17168 (N_17168,N_16461,N_16770);
nand U17169 (N_17169,N_16419,N_16649);
and U17170 (N_17170,N_16507,N_16500);
xnor U17171 (N_17171,N_16519,N_16579);
nand U17172 (N_17172,N_16465,N_16463);
or U17173 (N_17173,N_16733,N_16639);
or U17174 (N_17174,N_16786,N_16754);
nand U17175 (N_17175,N_16584,N_16710);
nor U17176 (N_17176,N_16769,N_16717);
nand U17177 (N_17177,N_16517,N_16613);
nor U17178 (N_17178,N_16617,N_16552);
or U17179 (N_17179,N_16520,N_16623);
or U17180 (N_17180,N_16754,N_16777);
nor U17181 (N_17181,N_16616,N_16573);
nor U17182 (N_17182,N_16522,N_16513);
nor U17183 (N_17183,N_16575,N_16747);
xor U17184 (N_17184,N_16456,N_16523);
nand U17185 (N_17185,N_16483,N_16604);
nand U17186 (N_17186,N_16491,N_16735);
xor U17187 (N_17187,N_16485,N_16680);
and U17188 (N_17188,N_16471,N_16485);
nand U17189 (N_17189,N_16607,N_16660);
xor U17190 (N_17190,N_16677,N_16594);
xor U17191 (N_17191,N_16432,N_16545);
and U17192 (N_17192,N_16779,N_16685);
or U17193 (N_17193,N_16722,N_16450);
xnor U17194 (N_17194,N_16444,N_16685);
or U17195 (N_17195,N_16644,N_16451);
xor U17196 (N_17196,N_16633,N_16589);
xor U17197 (N_17197,N_16472,N_16600);
xnor U17198 (N_17198,N_16407,N_16644);
nor U17199 (N_17199,N_16522,N_16438);
nor U17200 (N_17200,N_17068,N_17126);
nand U17201 (N_17201,N_17178,N_16846);
nand U17202 (N_17202,N_17116,N_16881);
xnor U17203 (N_17203,N_16888,N_16828);
and U17204 (N_17204,N_16989,N_16963);
nor U17205 (N_17205,N_17015,N_17179);
or U17206 (N_17206,N_16841,N_17092);
nand U17207 (N_17207,N_17001,N_16968);
nand U17208 (N_17208,N_16877,N_17098);
and U17209 (N_17209,N_16848,N_17081);
or U17210 (N_17210,N_16894,N_16920);
xor U17211 (N_17211,N_16842,N_16991);
and U17212 (N_17212,N_17004,N_17132);
xor U17213 (N_17213,N_16984,N_17194);
nor U17214 (N_17214,N_17187,N_16999);
nand U17215 (N_17215,N_16830,N_17054);
xnor U17216 (N_17216,N_17086,N_16837);
xor U17217 (N_17217,N_16823,N_17186);
nor U17218 (N_17218,N_17005,N_16982);
nand U17219 (N_17219,N_17046,N_16878);
xor U17220 (N_17220,N_17029,N_16880);
or U17221 (N_17221,N_17141,N_17119);
xnor U17222 (N_17222,N_16988,N_16806);
or U17223 (N_17223,N_17078,N_17157);
xor U17224 (N_17224,N_16914,N_17095);
nor U17225 (N_17225,N_16922,N_17090);
or U17226 (N_17226,N_17168,N_17025);
nor U17227 (N_17227,N_17175,N_17166);
nor U17228 (N_17228,N_17070,N_17173);
nand U17229 (N_17229,N_16923,N_17097);
xnor U17230 (N_17230,N_17129,N_16975);
nand U17231 (N_17231,N_16800,N_16857);
and U17232 (N_17232,N_17082,N_16936);
nor U17233 (N_17233,N_16942,N_16972);
nand U17234 (N_17234,N_16986,N_16882);
nand U17235 (N_17235,N_17016,N_17118);
xnor U17236 (N_17236,N_16898,N_17061);
and U17237 (N_17237,N_17076,N_16971);
xnor U17238 (N_17238,N_16805,N_16930);
and U17239 (N_17239,N_17146,N_17162);
xor U17240 (N_17240,N_16820,N_17109);
and U17241 (N_17241,N_16812,N_17130);
or U17242 (N_17242,N_16918,N_17043);
and U17243 (N_17243,N_16978,N_17160);
and U17244 (N_17244,N_17135,N_17096);
and U17245 (N_17245,N_17040,N_17042);
and U17246 (N_17246,N_16943,N_17142);
or U17247 (N_17247,N_17191,N_16960);
nand U17248 (N_17248,N_17094,N_16887);
or U17249 (N_17249,N_17053,N_16939);
and U17250 (N_17250,N_16948,N_16906);
or U17251 (N_17251,N_17003,N_16973);
or U17252 (N_17252,N_17190,N_17120);
or U17253 (N_17253,N_17169,N_16854);
xor U17254 (N_17254,N_16919,N_17152);
xnor U17255 (N_17255,N_16916,N_17007);
or U17256 (N_17256,N_16938,N_17019);
xor U17257 (N_17257,N_17083,N_17136);
and U17258 (N_17258,N_17006,N_17115);
or U17259 (N_17259,N_17080,N_16904);
and U17260 (N_17260,N_17000,N_16941);
nand U17261 (N_17261,N_16905,N_16970);
xnor U17262 (N_17262,N_17125,N_17075);
and U17263 (N_17263,N_17101,N_16847);
nor U17264 (N_17264,N_17189,N_16872);
nand U17265 (N_17265,N_16876,N_17147);
nand U17266 (N_17266,N_16947,N_16909);
nor U17267 (N_17267,N_17170,N_17032);
xor U17268 (N_17268,N_17071,N_17059);
nor U17269 (N_17269,N_16911,N_17117);
xor U17270 (N_17270,N_17084,N_17184);
or U17271 (N_17271,N_17056,N_16816);
nor U17272 (N_17272,N_17140,N_16833);
nor U17273 (N_17273,N_17150,N_17148);
xnor U17274 (N_17274,N_16871,N_16944);
xor U17275 (N_17275,N_17023,N_17085);
xor U17276 (N_17276,N_16822,N_17038);
nor U17277 (N_17277,N_17156,N_16875);
nand U17278 (N_17278,N_17195,N_17108);
nand U17279 (N_17279,N_17065,N_17182);
nor U17280 (N_17280,N_16890,N_16891);
nor U17281 (N_17281,N_16856,N_17072);
or U17282 (N_17282,N_17067,N_17105);
xor U17283 (N_17283,N_17088,N_17091);
xnor U17284 (N_17284,N_17181,N_17111);
xnor U17285 (N_17285,N_16958,N_16921);
nor U17286 (N_17286,N_17133,N_16860);
xor U17287 (N_17287,N_17051,N_17018);
or U17288 (N_17288,N_16865,N_16874);
xor U17289 (N_17289,N_16900,N_16996);
and U17290 (N_17290,N_16831,N_17196);
nor U17291 (N_17291,N_16992,N_17177);
nand U17292 (N_17292,N_16907,N_17013);
or U17293 (N_17293,N_16803,N_16953);
nor U17294 (N_17294,N_17161,N_17030);
nor U17295 (N_17295,N_17134,N_17055);
or U17296 (N_17296,N_17192,N_17028);
or U17297 (N_17297,N_17089,N_16836);
xor U17298 (N_17298,N_16926,N_17188);
xor U17299 (N_17299,N_17021,N_16834);
xnor U17300 (N_17300,N_16811,N_16908);
nand U17301 (N_17301,N_16807,N_17121);
and U17302 (N_17302,N_16813,N_16951);
and U17303 (N_17303,N_17048,N_16902);
nand U17304 (N_17304,N_16917,N_17110);
or U17305 (N_17305,N_16845,N_16949);
nor U17306 (N_17306,N_17014,N_17041);
xor U17307 (N_17307,N_16934,N_16819);
and U17308 (N_17308,N_16851,N_16966);
and U17309 (N_17309,N_17167,N_17149);
nor U17310 (N_17310,N_16852,N_17022);
nor U17311 (N_17311,N_17012,N_17128);
and U17312 (N_17312,N_16903,N_16873);
and U17313 (N_17313,N_17138,N_16897);
nand U17314 (N_17314,N_17011,N_17087);
and U17315 (N_17315,N_17064,N_17180);
and U17316 (N_17316,N_16885,N_16866);
nand U17317 (N_17317,N_16915,N_17139);
nand U17318 (N_17318,N_17060,N_17113);
nand U17319 (N_17319,N_16843,N_17020);
nor U17320 (N_17320,N_17073,N_16884);
xnor U17321 (N_17321,N_16962,N_16853);
or U17322 (N_17322,N_16801,N_16952);
or U17323 (N_17323,N_17102,N_16964);
nand U17324 (N_17324,N_17106,N_16835);
nand U17325 (N_17325,N_16855,N_17069);
or U17326 (N_17326,N_17010,N_17031);
nor U17327 (N_17327,N_16869,N_17045);
and U17328 (N_17328,N_16932,N_17062);
or U17329 (N_17329,N_16827,N_17198);
nand U17330 (N_17330,N_17079,N_16849);
or U17331 (N_17331,N_17144,N_17009);
nand U17332 (N_17332,N_16980,N_16928);
nor U17333 (N_17333,N_16867,N_16979);
and U17334 (N_17334,N_16955,N_17112);
xnor U17335 (N_17335,N_16965,N_17026);
nand U17336 (N_17336,N_17027,N_16879);
nor U17337 (N_17337,N_17104,N_17037);
or U17338 (N_17338,N_16861,N_17151);
or U17339 (N_17339,N_16998,N_16954);
xor U17340 (N_17340,N_16957,N_16981);
nor U17341 (N_17341,N_16976,N_17124);
xor U17342 (N_17342,N_16839,N_16995);
xnor U17343 (N_17343,N_16946,N_17172);
xnor U17344 (N_17344,N_16924,N_17131);
or U17345 (N_17345,N_16945,N_17039);
nand U17346 (N_17346,N_16912,N_17050);
or U17347 (N_17347,N_16832,N_16892);
nand U17348 (N_17348,N_16899,N_16913);
nand U17349 (N_17349,N_16977,N_16961);
xnor U17350 (N_17350,N_16937,N_16838);
xnor U17351 (N_17351,N_16883,N_17171);
and U17352 (N_17352,N_16993,N_16985);
and U17353 (N_17353,N_17047,N_16818);
nor U17354 (N_17354,N_16983,N_16829);
nand U17355 (N_17355,N_16844,N_16959);
or U17356 (N_17356,N_16933,N_16814);
and U17357 (N_17357,N_16901,N_17143);
or U17358 (N_17358,N_16858,N_17008);
xnor U17359 (N_17359,N_17099,N_17154);
nor U17360 (N_17360,N_17137,N_17057);
nand U17361 (N_17361,N_16910,N_17193);
nor U17362 (N_17362,N_16817,N_17024);
nor U17363 (N_17363,N_16927,N_16967);
nand U17364 (N_17364,N_16826,N_16956);
xor U17365 (N_17365,N_17034,N_17122);
nand U17366 (N_17366,N_16940,N_16950);
nor U17367 (N_17367,N_16895,N_16931);
and U17368 (N_17368,N_16815,N_17058);
or U17369 (N_17369,N_17077,N_16974);
xnor U17370 (N_17370,N_17159,N_17114);
xor U17371 (N_17371,N_17017,N_17183);
nor U17372 (N_17372,N_17127,N_17158);
xor U17373 (N_17373,N_17052,N_16859);
nor U17374 (N_17374,N_16886,N_17123);
nor U17375 (N_17375,N_17074,N_17036);
nor U17376 (N_17376,N_16997,N_16821);
or U17377 (N_17377,N_17155,N_16990);
and U17378 (N_17378,N_17049,N_17174);
xor U17379 (N_17379,N_17093,N_17153);
xor U17380 (N_17380,N_16868,N_17185);
nor U17381 (N_17381,N_16850,N_16863);
xnor U17382 (N_17382,N_16862,N_16825);
nor U17383 (N_17383,N_17199,N_16925);
and U17384 (N_17384,N_17165,N_17100);
and U17385 (N_17385,N_16804,N_17044);
and U17386 (N_17386,N_16896,N_17002);
and U17387 (N_17387,N_17066,N_16935);
nor U17388 (N_17388,N_16929,N_16808);
xnor U17389 (N_17389,N_16969,N_16824);
xor U17390 (N_17390,N_17103,N_17164);
xor U17391 (N_17391,N_17063,N_17035);
xnor U17392 (N_17392,N_16893,N_17197);
and U17393 (N_17393,N_16810,N_17107);
and U17394 (N_17394,N_16987,N_17163);
xnor U17395 (N_17395,N_16870,N_17176);
or U17396 (N_17396,N_16809,N_17145);
nand U17397 (N_17397,N_16994,N_16802);
nor U17398 (N_17398,N_16864,N_16889);
nor U17399 (N_17399,N_16840,N_17033);
xor U17400 (N_17400,N_16883,N_16994);
nor U17401 (N_17401,N_16898,N_16851);
nand U17402 (N_17402,N_17018,N_16968);
nand U17403 (N_17403,N_16897,N_16995);
and U17404 (N_17404,N_16959,N_17027);
nor U17405 (N_17405,N_16936,N_16988);
and U17406 (N_17406,N_16834,N_17139);
xor U17407 (N_17407,N_17109,N_17160);
and U17408 (N_17408,N_17047,N_16902);
or U17409 (N_17409,N_16849,N_17191);
nor U17410 (N_17410,N_16861,N_16843);
nor U17411 (N_17411,N_16942,N_17182);
xor U17412 (N_17412,N_17033,N_17091);
nor U17413 (N_17413,N_17161,N_17023);
or U17414 (N_17414,N_17147,N_17007);
and U17415 (N_17415,N_16862,N_17118);
nor U17416 (N_17416,N_17163,N_16830);
xor U17417 (N_17417,N_16809,N_16910);
or U17418 (N_17418,N_17094,N_16826);
and U17419 (N_17419,N_16997,N_16854);
nand U17420 (N_17420,N_16930,N_16899);
nand U17421 (N_17421,N_17056,N_16933);
nor U17422 (N_17422,N_16836,N_16800);
nor U17423 (N_17423,N_16818,N_17027);
and U17424 (N_17424,N_17031,N_17190);
nand U17425 (N_17425,N_17024,N_16926);
xnor U17426 (N_17426,N_16851,N_16847);
nor U17427 (N_17427,N_16891,N_16883);
nor U17428 (N_17428,N_17093,N_17161);
nor U17429 (N_17429,N_16882,N_17192);
nor U17430 (N_17430,N_16806,N_17128);
or U17431 (N_17431,N_16944,N_17114);
nand U17432 (N_17432,N_16879,N_16840);
xor U17433 (N_17433,N_16989,N_17094);
and U17434 (N_17434,N_16986,N_17086);
and U17435 (N_17435,N_17018,N_17107);
and U17436 (N_17436,N_16960,N_17022);
xnor U17437 (N_17437,N_17184,N_16996);
xor U17438 (N_17438,N_17186,N_16903);
or U17439 (N_17439,N_16839,N_16971);
nor U17440 (N_17440,N_16898,N_17060);
nor U17441 (N_17441,N_16982,N_17064);
xnor U17442 (N_17442,N_16809,N_17022);
nor U17443 (N_17443,N_16837,N_16862);
and U17444 (N_17444,N_16962,N_16809);
or U17445 (N_17445,N_17128,N_17161);
nor U17446 (N_17446,N_17163,N_17030);
and U17447 (N_17447,N_17014,N_16925);
nand U17448 (N_17448,N_16897,N_16941);
xor U17449 (N_17449,N_17032,N_16840);
and U17450 (N_17450,N_17078,N_16833);
or U17451 (N_17451,N_17153,N_16980);
or U17452 (N_17452,N_16878,N_16834);
nand U17453 (N_17453,N_16835,N_17072);
nand U17454 (N_17454,N_16892,N_17174);
xor U17455 (N_17455,N_17136,N_16839);
nor U17456 (N_17456,N_17041,N_17005);
or U17457 (N_17457,N_16853,N_17035);
nor U17458 (N_17458,N_16961,N_17184);
xnor U17459 (N_17459,N_17049,N_16844);
or U17460 (N_17460,N_16925,N_16842);
xor U17461 (N_17461,N_16873,N_16973);
nand U17462 (N_17462,N_17084,N_16912);
nand U17463 (N_17463,N_16849,N_17161);
nor U17464 (N_17464,N_17055,N_16923);
xnor U17465 (N_17465,N_17021,N_17120);
nand U17466 (N_17466,N_17163,N_16935);
nor U17467 (N_17467,N_16914,N_17138);
xor U17468 (N_17468,N_17117,N_16992);
nor U17469 (N_17469,N_17076,N_17188);
or U17470 (N_17470,N_17160,N_16910);
xor U17471 (N_17471,N_16815,N_17123);
nor U17472 (N_17472,N_16939,N_17082);
xor U17473 (N_17473,N_17130,N_17163);
xnor U17474 (N_17474,N_16976,N_17012);
nand U17475 (N_17475,N_16955,N_17180);
nor U17476 (N_17476,N_16851,N_16843);
and U17477 (N_17477,N_17068,N_17041);
nand U17478 (N_17478,N_16871,N_16817);
xnor U17479 (N_17479,N_16918,N_17080);
and U17480 (N_17480,N_16974,N_16841);
xnor U17481 (N_17481,N_17091,N_16870);
nor U17482 (N_17482,N_16985,N_16862);
or U17483 (N_17483,N_16957,N_16905);
and U17484 (N_17484,N_17040,N_17041);
and U17485 (N_17485,N_17061,N_17095);
xor U17486 (N_17486,N_17106,N_16851);
nor U17487 (N_17487,N_16963,N_17001);
nand U17488 (N_17488,N_16902,N_16836);
xor U17489 (N_17489,N_17026,N_16868);
and U17490 (N_17490,N_17065,N_17020);
nand U17491 (N_17491,N_16847,N_16965);
nor U17492 (N_17492,N_16979,N_16880);
and U17493 (N_17493,N_17066,N_17044);
xor U17494 (N_17494,N_17175,N_16914);
nor U17495 (N_17495,N_16944,N_17100);
nand U17496 (N_17496,N_17087,N_16887);
xor U17497 (N_17497,N_16886,N_16879);
xor U17498 (N_17498,N_17035,N_17131);
and U17499 (N_17499,N_16889,N_16825);
and U17500 (N_17500,N_16897,N_17121);
xnor U17501 (N_17501,N_16998,N_16923);
nor U17502 (N_17502,N_16954,N_16991);
nand U17503 (N_17503,N_16882,N_17148);
nand U17504 (N_17504,N_16981,N_16984);
and U17505 (N_17505,N_17028,N_16826);
nor U17506 (N_17506,N_16844,N_17004);
nor U17507 (N_17507,N_17124,N_17109);
xor U17508 (N_17508,N_16972,N_17104);
and U17509 (N_17509,N_16960,N_16948);
and U17510 (N_17510,N_16925,N_16998);
nor U17511 (N_17511,N_16937,N_17090);
nor U17512 (N_17512,N_16886,N_16943);
and U17513 (N_17513,N_16857,N_16817);
nand U17514 (N_17514,N_17142,N_17146);
xnor U17515 (N_17515,N_16851,N_16875);
nand U17516 (N_17516,N_16920,N_17083);
nor U17517 (N_17517,N_16855,N_16955);
xor U17518 (N_17518,N_17085,N_16868);
or U17519 (N_17519,N_17029,N_16901);
xor U17520 (N_17520,N_16959,N_17016);
and U17521 (N_17521,N_16969,N_17021);
xnor U17522 (N_17522,N_16898,N_16849);
xor U17523 (N_17523,N_17138,N_17013);
and U17524 (N_17524,N_17147,N_16960);
and U17525 (N_17525,N_16961,N_16971);
and U17526 (N_17526,N_17162,N_16919);
and U17527 (N_17527,N_17103,N_17010);
or U17528 (N_17528,N_16845,N_16953);
nand U17529 (N_17529,N_17129,N_17077);
and U17530 (N_17530,N_16885,N_17155);
or U17531 (N_17531,N_17007,N_16826);
and U17532 (N_17532,N_17185,N_17009);
nor U17533 (N_17533,N_17173,N_16940);
and U17534 (N_17534,N_16875,N_16961);
or U17535 (N_17535,N_16966,N_17182);
or U17536 (N_17536,N_16960,N_17189);
xor U17537 (N_17537,N_16992,N_16981);
nor U17538 (N_17538,N_17031,N_17138);
nor U17539 (N_17539,N_17126,N_17030);
xnor U17540 (N_17540,N_17154,N_16972);
nand U17541 (N_17541,N_16960,N_16890);
and U17542 (N_17542,N_17116,N_17195);
and U17543 (N_17543,N_16813,N_16843);
nor U17544 (N_17544,N_17193,N_16960);
and U17545 (N_17545,N_17163,N_16906);
xor U17546 (N_17546,N_16916,N_17141);
or U17547 (N_17547,N_16803,N_17064);
and U17548 (N_17548,N_17120,N_17111);
nand U17549 (N_17549,N_16854,N_16898);
nor U17550 (N_17550,N_16802,N_16974);
or U17551 (N_17551,N_16958,N_16951);
nor U17552 (N_17552,N_17181,N_17120);
nor U17553 (N_17553,N_17042,N_16810);
or U17554 (N_17554,N_17162,N_16999);
xor U17555 (N_17555,N_17048,N_16903);
nor U17556 (N_17556,N_17068,N_16990);
xnor U17557 (N_17557,N_16802,N_17044);
xor U17558 (N_17558,N_17040,N_16902);
xor U17559 (N_17559,N_16913,N_16803);
and U17560 (N_17560,N_17075,N_16840);
nor U17561 (N_17561,N_16800,N_17195);
nor U17562 (N_17562,N_17055,N_16887);
and U17563 (N_17563,N_17083,N_16968);
nor U17564 (N_17564,N_16900,N_17198);
xnor U17565 (N_17565,N_16962,N_16944);
xnor U17566 (N_17566,N_17035,N_17028);
and U17567 (N_17567,N_17170,N_17003);
nor U17568 (N_17568,N_17185,N_16835);
nor U17569 (N_17569,N_16909,N_17179);
nand U17570 (N_17570,N_16869,N_17039);
or U17571 (N_17571,N_17100,N_17080);
and U17572 (N_17572,N_16888,N_17181);
and U17573 (N_17573,N_16976,N_16881);
nor U17574 (N_17574,N_17053,N_17107);
nand U17575 (N_17575,N_17160,N_17108);
nand U17576 (N_17576,N_16904,N_17083);
xor U17577 (N_17577,N_17161,N_16987);
or U17578 (N_17578,N_16867,N_17118);
nand U17579 (N_17579,N_17111,N_16861);
nor U17580 (N_17580,N_16881,N_17117);
nand U17581 (N_17581,N_16935,N_17070);
nand U17582 (N_17582,N_16805,N_17079);
xor U17583 (N_17583,N_17038,N_16902);
nand U17584 (N_17584,N_17079,N_17185);
xor U17585 (N_17585,N_17052,N_17113);
or U17586 (N_17586,N_17151,N_16884);
nor U17587 (N_17587,N_17145,N_17127);
or U17588 (N_17588,N_17023,N_17117);
nand U17589 (N_17589,N_17001,N_16983);
nor U17590 (N_17590,N_16820,N_16862);
nand U17591 (N_17591,N_17178,N_17097);
nand U17592 (N_17592,N_16867,N_17005);
nor U17593 (N_17593,N_16919,N_17133);
xor U17594 (N_17594,N_17014,N_17094);
nand U17595 (N_17595,N_17094,N_16853);
or U17596 (N_17596,N_16824,N_17167);
nor U17597 (N_17597,N_17122,N_17089);
or U17598 (N_17598,N_17097,N_17089);
nor U17599 (N_17599,N_16943,N_17067);
or U17600 (N_17600,N_17486,N_17257);
or U17601 (N_17601,N_17392,N_17246);
nand U17602 (N_17602,N_17493,N_17573);
nor U17603 (N_17603,N_17429,N_17581);
or U17604 (N_17604,N_17218,N_17456);
nor U17605 (N_17605,N_17331,N_17527);
xnor U17606 (N_17606,N_17343,N_17589);
or U17607 (N_17607,N_17567,N_17446);
or U17608 (N_17608,N_17220,N_17510);
or U17609 (N_17609,N_17405,N_17263);
nand U17610 (N_17610,N_17404,N_17275);
nor U17611 (N_17611,N_17340,N_17396);
nand U17612 (N_17612,N_17289,N_17598);
xor U17613 (N_17613,N_17465,N_17251);
and U17614 (N_17614,N_17454,N_17500);
nand U17615 (N_17615,N_17406,N_17517);
nand U17616 (N_17616,N_17415,N_17212);
nand U17617 (N_17617,N_17496,N_17498);
nor U17618 (N_17618,N_17325,N_17278);
and U17619 (N_17619,N_17252,N_17552);
nor U17620 (N_17620,N_17323,N_17580);
and U17621 (N_17621,N_17308,N_17485);
nor U17622 (N_17622,N_17386,N_17240);
nor U17623 (N_17623,N_17480,N_17588);
nand U17624 (N_17624,N_17563,N_17221);
xnor U17625 (N_17625,N_17298,N_17487);
nor U17626 (N_17626,N_17582,N_17248);
xor U17627 (N_17627,N_17381,N_17261);
xor U17628 (N_17628,N_17238,N_17526);
or U17629 (N_17629,N_17349,N_17488);
nand U17630 (N_17630,N_17472,N_17231);
xor U17631 (N_17631,N_17314,N_17514);
or U17632 (N_17632,N_17471,N_17372);
and U17633 (N_17633,N_17499,N_17360);
or U17634 (N_17634,N_17539,N_17395);
or U17635 (N_17635,N_17342,N_17365);
xor U17636 (N_17636,N_17225,N_17470);
or U17637 (N_17637,N_17203,N_17548);
and U17638 (N_17638,N_17215,N_17451);
xor U17639 (N_17639,N_17511,N_17286);
and U17640 (N_17640,N_17371,N_17434);
nor U17641 (N_17641,N_17358,N_17455);
nand U17642 (N_17642,N_17482,N_17583);
or U17643 (N_17643,N_17244,N_17418);
nor U17644 (N_17644,N_17576,N_17353);
xor U17645 (N_17645,N_17394,N_17422);
xnor U17646 (N_17646,N_17276,N_17309);
or U17647 (N_17647,N_17448,N_17361);
xnor U17648 (N_17648,N_17250,N_17544);
xnor U17649 (N_17649,N_17345,N_17299);
nor U17650 (N_17650,N_17237,N_17282);
or U17651 (N_17651,N_17380,N_17436);
nor U17652 (N_17652,N_17437,N_17214);
or U17653 (N_17653,N_17202,N_17297);
or U17654 (N_17654,N_17443,N_17397);
or U17655 (N_17655,N_17574,N_17586);
nor U17656 (N_17656,N_17599,N_17206);
and U17657 (N_17657,N_17277,N_17211);
and U17658 (N_17658,N_17462,N_17389);
or U17659 (N_17659,N_17233,N_17440);
nor U17660 (N_17660,N_17374,N_17337);
xnor U17661 (N_17661,N_17288,N_17505);
or U17662 (N_17662,N_17216,N_17270);
xor U17663 (N_17663,N_17529,N_17327);
or U17664 (N_17664,N_17584,N_17302);
and U17665 (N_17665,N_17333,N_17311);
xnor U17666 (N_17666,N_17304,N_17306);
and U17667 (N_17667,N_17312,N_17507);
xnor U17668 (N_17668,N_17439,N_17279);
and U17669 (N_17669,N_17255,N_17457);
and U17670 (N_17670,N_17525,N_17541);
nor U17671 (N_17671,N_17356,N_17452);
nand U17672 (N_17672,N_17408,N_17483);
or U17673 (N_17673,N_17272,N_17481);
xnor U17674 (N_17674,N_17398,N_17477);
or U17675 (N_17675,N_17503,N_17591);
xor U17676 (N_17676,N_17375,N_17569);
nand U17677 (N_17677,N_17593,N_17370);
or U17678 (N_17678,N_17217,N_17219);
xnor U17679 (N_17679,N_17550,N_17254);
or U17680 (N_17680,N_17473,N_17322);
nand U17681 (N_17681,N_17549,N_17538);
xnor U17682 (N_17682,N_17502,N_17540);
xnor U17683 (N_17683,N_17401,N_17319);
nor U17684 (N_17684,N_17543,N_17449);
or U17685 (N_17685,N_17256,N_17243);
xnor U17686 (N_17686,N_17478,N_17287);
nor U17687 (N_17687,N_17445,N_17284);
or U17688 (N_17688,N_17504,N_17561);
or U17689 (N_17689,N_17587,N_17423);
nor U17690 (N_17690,N_17283,N_17435);
or U17691 (N_17691,N_17348,N_17267);
or U17692 (N_17692,N_17513,N_17534);
or U17693 (N_17693,N_17391,N_17224);
nand U17694 (N_17694,N_17229,N_17508);
and U17695 (N_17695,N_17400,N_17377);
xnor U17696 (N_17696,N_17411,N_17533);
nor U17697 (N_17697,N_17274,N_17317);
nand U17698 (N_17698,N_17223,N_17491);
xor U17699 (N_17699,N_17557,N_17512);
and U17700 (N_17700,N_17303,N_17575);
or U17701 (N_17701,N_17554,N_17245);
nand U17702 (N_17702,N_17442,N_17560);
or U17703 (N_17703,N_17556,N_17373);
nand U17704 (N_17704,N_17438,N_17447);
xor U17705 (N_17705,N_17547,N_17518);
xnor U17706 (N_17706,N_17444,N_17249);
or U17707 (N_17707,N_17268,N_17357);
nor U17708 (N_17708,N_17232,N_17459);
nand U17709 (N_17709,N_17264,N_17516);
or U17710 (N_17710,N_17201,N_17200);
xnor U17711 (N_17711,N_17528,N_17281);
nand U17712 (N_17712,N_17355,N_17464);
xor U17713 (N_17713,N_17585,N_17292);
nand U17714 (N_17714,N_17553,N_17568);
nand U17715 (N_17715,N_17432,N_17463);
nor U17716 (N_17716,N_17242,N_17354);
nor U17717 (N_17717,N_17524,N_17426);
or U17718 (N_17718,N_17594,N_17383);
or U17719 (N_17719,N_17506,N_17326);
or U17720 (N_17720,N_17546,N_17388);
xor U17721 (N_17721,N_17376,N_17566);
and U17722 (N_17722,N_17346,N_17402);
or U17723 (N_17723,N_17328,N_17310);
nor U17724 (N_17724,N_17424,N_17522);
or U17725 (N_17725,N_17570,N_17536);
or U17726 (N_17726,N_17403,N_17597);
xnor U17727 (N_17727,N_17466,N_17321);
or U17728 (N_17728,N_17571,N_17519);
nand U17729 (N_17729,N_17207,N_17461);
nor U17730 (N_17730,N_17351,N_17595);
or U17731 (N_17731,N_17523,N_17565);
nor U17732 (N_17732,N_17430,N_17531);
nand U17733 (N_17733,N_17421,N_17542);
nor U17734 (N_17734,N_17271,N_17338);
nor U17735 (N_17735,N_17367,N_17259);
xor U17736 (N_17736,N_17280,N_17262);
nor U17737 (N_17737,N_17362,N_17460);
nor U17738 (N_17738,N_17562,N_17416);
or U17739 (N_17739,N_17399,N_17222);
nor U17740 (N_17740,N_17551,N_17545);
or U17741 (N_17741,N_17420,N_17204);
xor U17742 (N_17742,N_17450,N_17307);
nor U17743 (N_17743,N_17468,N_17425);
nor U17744 (N_17744,N_17407,N_17427);
or U17745 (N_17745,N_17414,N_17269);
and U17746 (N_17746,N_17295,N_17369);
and U17747 (N_17747,N_17318,N_17316);
or U17748 (N_17748,N_17339,N_17273);
xnor U17749 (N_17749,N_17209,N_17558);
nand U17750 (N_17750,N_17341,N_17347);
xor U17751 (N_17751,N_17555,N_17489);
nor U17752 (N_17752,N_17363,N_17492);
nor U17753 (N_17753,N_17332,N_17228);
nor U17754 (N_17754,N_17320,N_17359);
or U17755 (N_17755,N_17532,N_17296);
nor U17756 (N_17756,N_17413,N_17335);
or U17757 (N_17757,N_17501,N_17479);
nor U17758 (N_17758,N_17564,N_17592);
or U17759 (N_17759,N_17409,N_17227);
nor U17760 (N_17760,N_17329,N_17330);
nor U17761 (N_17761,N_17521,N_17324);
nor U17762 (N_17762,N_17520,N_17241);
or U17763 (N_17763,N_17537,N_17490);
nand U17764 (N_17764,N_17412,N_17260);
xor U17765 (N_17765,N_17266,N_17453);
xor U17766 (N_17766,N_17265,N_17382);
nor U17767 (N_17767,N_17535,N_17213);
or U17768 (N_17768,N_17475,N_17234);
nor U17769 (N_17769,N_17578,N_17334);
or U17770 (N_17770,N_17226,N_17344);
xnor U17771 (N_17771,N_17305,N_17253);
xor U17772 (N_17772,N_17431,N_17419);
nand U17773 (N_17773,N_17497,N_17293);
xor U17774 (N_17774,N_17495,N_17291);
nand U17775 (N_17775,N_17258,N_17384);
or U17776 (N_17776,N_17559,N_17290);
nor U17777 (N_17777,N_17469,N_17205);
xnor U17778 (N_17778,N_17247,N_17350);
xor U17779 (N_17779,N_17300,N_17210);
xnor U17780 (N_17780,N_17458,N_17467);
or U17781 (N_17781,N_17315,N_17410);
nand U17782 (N_17782,N_17208,N_17590);
nand U17783 (N_17783,N_17494,N_17379);
nand U17784 (N_17784,N_17572,N_17484);
xor U17785 (N_17785,N_17294,N_17366);
nand U17786 (N_17786,N_17378,N_17441);
xor U17787 (N_17787,N_17530,N_17239);
xnor U17788 (N_17788,N_17393,N_17236);
xor U17789 (N_17789,N_17474,N_17235);
or U17790 (N_17790,N_17417,N_17509);
nor U17791 (N_17791,N_17336,N_17301);
or U17792 (N_17792,N_17352,N_17368);
or U17793 (N_17793,N_17387,N_17390);
and U17794 (N_17794,N_17433,N_17596);
nand U17795 (N_17795,N_17579,N_17577);
or U17796 (N_17796,N_17230,N_17285);
nor U17797 (N_17797,N_17385,N_17313);
and U17798 (N_17798,N_17364,N_17428);
and U17799 (N_17799,N_17515,N_17476);
nand U17800 (N_17800,N_17376,N_17401);
nor U17801 (N_17801,N_17275,N_17579);
nand U17802 (N_17802,N_17546,N_17558);
and U17803 (N_17803,N_17511,N_17205);
xor U17804 (N_17804,N_17477,N_17377);
nor U17805 (N_17805,N_17400,N_17518);
nor U17806 (N_17806,N_17310,N_17206);
or U17807 (N_17807,N_17228,N_17493);
and U17808 (N_17808,N_17499,N_17555);
nor U17809 (N_17809,N_17472,N_17409);
nand U17810 (N_17810,N_17389,N_17486);
or U17811 (N_17811,N_17514,N_17387);
nor U17812 (N_17812,N_17407,N_17547);
or U17813 (N_17813,N_17534,N_17236);
nand U17814 (N_17814,N_17492,N_17426);
and U17815 (N_17815,N_17386,N_17532);
nand U17816 (N_17816,N_17415,N_17315);
nand U17817 (N_17817,N_17499,N_17551);
nand U17818 (N_17818,N_17210,N_17460);
nor U17819 (N_17819,N_17359,N_17318);
xnor U17820 (N_17820,N_17357,N_17465);
and U17821 (N_17821,N_17340,N_17272);
and U17822 (N_17822,N_17541,N_17348);
xnor U17823 (N_17823,N_17231,N_17538);
nand U17824 (N_17824,N_17456,N_17465);
or U17825 (N_17825,N_17470,N_17584);
xnor U17826 (N_17826,N_17581,N_17272);
nor U17827 (N_17827,N_17269,N_17561);
and U17828 (N_17828,N_17569,N_17541);
xor U17829 (N_17829,N_17549,N_17443);
and U17830 (N_17830,N_17517,N_17325);
or U17831 (N_17831,N_17520,N_17563);
or U17832 (N_17832,N_17473,N_17317);
xor U17833 (N_17833,N_17554,N_17385);
nand U17834 (N_17834,N_17337,N_17250);
or U17835 (N_17835,N_17561,N_17526);
and U17836 (N_17836,N_17454,N_17427);
and U17837 (N_17837,N_17532,N_17445);
and U17838 (N_17838,N_17217,N_17469);
xor U17839 (N_17839,N_17377,N_17443);
and U17840 (N_17840,N_17326,N_17373);
and U17841 (N_17841,N_17532,N_17535);
xor U17842 (N_17842,N_17210,N_17257);
nor U17843 (N_17843,N_17517,N_17476);
nor U17844 (N_17844,N_17491,N_17455);
and U17845 (N_17845,N_17432,N_17375);
nor U17846 (N_17846,N_17240,N_17441);
xor U17847 (N_17847,N_17377,N_17319);
xor U17848 (N_17848,N_17563,N_17476);
nand U17849 (N_17849,N_17521,N_17322);
or U17850 (N_17850,N_17549,N_17399);
or U17851 (N_17851,N_17365,N_17230);
or U17852 (N_17852,N_17347,N_17470);
nand U17853 (N_17853,N_17259,N_17487);
and U17854 (N_17854,N_17286,N_17229);
or U17855 (N_17855,N_17501,N_17200);
xor U17856 (N_17856,N_17389,N_17273);
nor U17857 (N_17857,N_17430,N_17307);
nor U17858 (N_17858,N_17582,N_17595);
nor U17859 (N_17859,N_17280,N_17225);
and U17860 (N_17860,N_17383,N_17476);
xor U17861 (N_17861,N_17486,N_17252);
and U17862 (N_17862,N_17274,N_17453);
xor U17863 (N_17863,N_17446,N_17447);
xor U17864 (N_17864,N_17446,N_17538);
or U17865 (N_17865,N_17450,N_17242);
or U17866 (N_17866,N_17445,N_17215);
and U17867 (N_17867,N_17565,N_17459);
or U17868 (N_17868,N_17507,N_17581);
nor U17869 (N_17869,N_17480,N_17393);
and U17870 (N_17870,N_17373,N_17421);
or U17871 (N_17871,N_17527,N_17498);
nor U17872 (N_17872,N_17542,N_17505);
and U17873 (N_17873,N_17266,N_17496);
nor U17874 (N_17874,N_17435,N_17388);
or U17875 (N_17875,N_17442,N_17507);
nand U17876 (N_17876,N_17456,N_17533);
nor U17877 (N_17877,N_17488,N_17213);
or U17878 (N_17878,N_17523,N_17414);
nand U17879 (N_17879,N_17231,N_17463);
or U17880 (N_17880,N_17498,N_17487);
nand U17881 (N_17881,N_17243,N_17437);
and U17882 (N_17882,N_17389,N_17342);
nand U17883 (N_17883,N_17588,N_17352);
xor U17884 (N_17884,N_17593,N_17468);
nor U17885 (N_17885,N_17220,N_17334);
nor U17886 (N_17886,N_17473,N_17480);
nand U17887 (N_17887,N_17582,N_17520);
xor U17888 (N_17888,N_17519,N_17490);
and U17889 (N_17889,N_17395,N_17565);
nand U17890 (N_17890,N_17524,N_17423);
or U17891 (N_17891,N_17525,N_17262);
nand U17892 (N_17892,N_17228,N_17550);
or U17893 (N_17893,N_17380,N_17470);
or U17894 (N_17894,N_17488,N_17230);
nand U17895 (N_17895,N_17297,N_17349);
or U17896 (N_17896,N_17228,N_17465);
or U17897 (N_17897,N_17533,N_17331);
xnor U17898 (N_17898,N_17453,N_17340);
and U17899 (N_17899,N_17353,N_17366);
xnor U17900 (N_17900,N_17522,N_17402);
and U17901 (N_17901,N_17446,N_17312);
nand U17902 (N_17902,N_17488,N_17212);
nor U17903 (N_17903,N_17575,N_17267);
and U17904 (N_17904,N_17510,N_17563);
or U17905 (N_17905,N_17285,N_17236);
nor U17906 (N_17906,N_17479,N_17255);
xor U17907 (N_17907,N_17595,N_17469);
nor U17908 (N_17908,N_17275,N_17412);
or U17909 (N_17909,N_17335,N_17362);
or U17910 (N_17910,N_17541,N_17212);
or U17911 (N_17911,N_17258,N_17420);
nand U17912 (N_17912,N_17579,N_17235);
or U17913 (N_17913,N_17411,N_17527);
nor U17914 (N_17914,N_17549,N_17555);
or U17915 (N_17915,N_17372,N_17499);
and U17916 (N_17916,N_17457,N_17287);
nand U17917 (N_17917,N_17314,N_17583);
and U17918 (N_17918,N_17211,N_17460);
nor U17919 (N_17919,N_17406,N_17259);
or U17920 (N_17920,N_17548,N_17457);
nor U17921 (N_17921,N_17241,N_17287);
nor U17922 (N_17922,N_17499,N_17525);
xor U17923 (N_17923,N_17275,N_17324);
nor U17924 (N_17924,N_17377,N_17426);
nor U17925 (N_17925,N_17249,N_17465);
nor U17926 (N_17926,N_17597,N_17336);
nor U17927 (N_17927,N_17390,N_17338);
nand U17928 (N_17928,N_17424,N_17441);
or U17929 (N_17929,N_17555,N_17302);
and U17930 (N_17930,N_17256,N_17342);
nor U17931 (N_17931,N_17440,N_17475);
xor U17932 (N_17932,N_17283,N_17523);
or U17933 (N_17933,N_17352,N_17284);
or U17934 (N_17934,N_17286,N_17441);
or U17935 (N_17935,N_17459,N_17213);
nor U17936 (N_17936,N_17540,N_17222);
xor U17937 (N_17937,N_17558,N_17525);
and U17938 (N_17938,N_17541,N_17495);
xor U17939 (N_17939,N_17496,N_17577);
nor U17940 (N_17940,N_17467,N_17247);
nor U17941 (N_17941,N_17306,N_17483);
or U17942 (N_17942,N_17213,N_17396);
nand U17943 (N_17943,N_17225,N_17446);
nand U17944 (N_17944,N_17265,N_17364);
or U17945 (N_17945,N_17387,N_17506);
nand U17946 (N_17946,N_17426,N_17261);
and U17947 (N_17947,N_17420,N_17440);
nand U17948 (N_17948,N_17442,N_17246);
and U17949 (N_17949,N_17526,N_17322);
nor U17950 (N_17950,N_17299,N_17342);
nor U17951 (N_17951,N_17536,N_17561);
nor U17952 (N_17952,N_17338,N_17205);
xor U17953 (N_17953,N_17364,N_17459);
nand U17954 (N_17954,N_17411,N_17484);
and U17955 (N_17955,N_17465,N_17308);
xnor U17956 (N_17956,N_17415,N_17259);
nor U17957 (N_17957,N_17298,N_17297);
and U17958 (N_17958,N_17240,N_17242);
nor U17959 (N_17959,N_17207,N_17554);
nor U17960 (N_17960,N_17420,N_17597);
and U17961 (N_17961,N_17297,N_17350);
and U17962 (N_17962,N_17420,N_17493);
nor U17963 (N_17963,N_17293,N_17530);
or U17964 (N_17964,N_17262,N_17306);
or U17965 (N_17965,N_17401,N_17444);
or U17966 (N_17966,N_17248,N_17221);
xor U17967 (N_17967,N_17550,N_17449);
nand U17968 (N_17968,N_17266,N_17590);
and U17969 (N_17969,N_17542,N_17585);
or U17970 (N_17970,N_17233,N_17378);
nor U17971 (N_17971,N_17519,N_17564);
nor U17972 (N_17972,N_17385,N_17228);
nor U17973 (N_17973,N_17488,N_17485);
nand U17974 (N_17974,N_17317,N_17351);
xnor U17975 (N_17975,N_17450,N_17346);
xor U17976 (N_17976,N_17448,N_17410);
and U17977 (N_17977,N_17232,N_17581);
nand U17978 (N_17978,N_17589,N_17595);
nand U17979 (N_17979,N_17467,N_17489);
nor U17980 (N_17980,N_17312,N_17465);
nor U17981 (N_17981,N_17530,N_17248);
or U17982 (N_17982,N_17375,N_17559);
xnor U17983 (N_17983,N_17473,N_17554);
nand U17984 (N_17984,N_17253,N_17510);
nor U17985 (N_17985,N_17430,N_17372);
xor U17986 (N_17986,N_17307,N_17475);
nor U17987 (N_17987,N_17422,N_17563);
or U17988 (N_17988,N_17306,N_17418);
or U17989 (N_17989,N_17446,N_17425);
nor U17990 (N_17990,N_17275,N_17486);
and U17991 (N_17991,N_17435,N_17359);
and U17992 (N_17992,N_17513,N_17486);
xor U17993 (N_17993,N_17350,N_17349);
or U17994 (N_17994,N_17589,N_17261);
and U17995 (N_17995,N_17370,N_17315);
xnor U17996 (N_17996,N_17529,N_17378);
xor U17997 (N_17997,N_17557,N_17515);
nor U17998 (N_17998,N_17471,N_17523);
or U17999 (N_17999,N_17326,N_17422);
nor U18000 (N_18000,N_17654,N_17770);
xor U18001 (N_18001,N_17860,N_17635);
xor U18002 (N_18002,N_17804,N_17851);
xnor U18003 (N_18003,N_17863,N_17815);
xnor U18004 (N_18004,N_17631,N_17980);
nor U18005 (N_18005,N_17945,N_17961);
xnor U18006 (N_18006,N_17866,N_17652);
nand U18007 (N_18007,N_17659,N_17898);
xor U18008 (N_18008,N_17943,N_17732);
and U18009 (N_18009,N_17979,N_17810);
nor U18010 (N_18010,N_17977,N_17890);
or U18011 (N_18011,N_17701,N_17621);
xnor U18012 (N_18012,N_17957,N_17773);
nand U18013 (N_18013,N_17953,N_17829);
or U18014 (N_18014,N_17681,N_17988);
nor U18015 (N_18015,N_17787,N_17775);
or U18016 (N_18016,N_17833,N_17784);
nand U18017 (N_18017,N_17794,N_17625);
nand U18018 (N_18018,N_17765,N_17856);
or U18019 (N_18019,N_17616,N_17710);
or U18020 (N_18020,N_17627,N_17912);
xnor U18021 (N_18021,N_17926,N_17666);
or U18022 (N_18022,N_17924,N_17682);
or U18023 (N_18023,N_17981,N_17747);
xor U18024 (N_18024,N_17764,N_17956);
or U18025 (N_18025,N_17954,N_17964);
or U18026 (N_18026,N_17626,N_17995);
xnor U18027 (N_18027,N_17600,N_17936);
and U18028 (N_18028,N_17842,N_17855);
or U18029 (N_18029,N_17861,N_17673);
xor U18030 (N_18030,N_17858,N_17947);
nor U18031 (N_18031,N_17997,N_17668);
and U18032 (N_18032,N_17606,N_17677);
nor U18033 (N_18033,N_17788,N_17660);
and U18034 (N_18034,N_17613,N_17727);
xor U18035 (N_18035,N_17739,N_17743);
nor U18036 (N_18036,N_17604,N_17644);
or U18037 (N_18037,N_17874,N_17744);
xor U18038 (N_18038,N_17708,N_17768);
and U18039 (N_18039,N_17657,N_17946);
nand U18040 (N_18040,N_17756,N_17812);
nor U18041 (N_18041,N_17748,N_17901);
and U18042 (N_18042,N_17751,N_17884);
or U18043 (N_18043,N_17862,N_17904);
nand U18044 (N_18044,N_17753,N_17822);
xor U18045 (N_18045,N_17647,N_17892);
nor U18046 (N_18046,N_17746,N_17993);
nand U18047 (N_18047,N_17785,N_17929);
xor U18048 (N_18048,N_17909,N_17941);
nor U18049 (N_18049,N_17820,N_17645);
nor U18050 (N_18050,N_17602,N_17601);
or U18051 (N_18051,N_17903,N_17694);
or U18052 (N_18052,N_17932,N_17796);
nor U18053 (N_18053,N_17769,N_17617);
nand U18054 (N_18054,N_17871,N_17832);
and U18055 (N_18055,N_17888,N_17913);
xor U18056 (N_18056,N_17891,N_17907);
xor U18057 (N_18057,N_17974,N_17758);
nor U18058 (N_18058,N_17779,N_17830);
or U18059 (N_18059,N_17911,N_17763);
nor U18060 (N_18060,N_17948,N_17847);
xnor U18061 (N_18061,N_17735,N_17843);
or U18062 (N_18062,N_17693,N_17823);
xnor U18063 (N_18063,N_17648,N_17699);
xnor U18064 (N_18064,N_17797,N_17879);
or U18065 (N_18065,N_17703,N_17940);
nand U18066 (N_18066,N_17618,N_17813);
or U18067 (N_18067,N_17986,N_17987);
xnor U18068 (N_18068,N_17878,N_17915);
and U18069 (N_18069,N_17725,N_17730);
or U18070 (N_18070,N_17609,N_17615);
or U18071 (N_18071,N_17837,N_17684);
nand U18072 (N_18072,N_17854,N_17695);
or U18073 (N_18073,N_17786,N_17723);
nor U18074 (N_18074,N_17908,N_17774);
xor U18075 (N_18075,N_17887,N_17629);
nor U18076 (N_18076,N_17937,N_17930);
nor U18077 (N_18077,N_17722,N_17881);
and U18078 (N_18078,N_17653,N_17916);
nand U18079 (N_18079,N_17959,N_17679);
or U18080 (N_18080,N_17641,N_17781);
xnor U18081 (N_18081,N_17938,N_17783);
xnor U18082 (N_18082,N_17857,N_17935);
xnor U18083 (N_18083,N_17726,N_17814);
and U18084 (N_18084,N_17894,N_17720);
xor U18085 (N_18085,N_17712,N_17738);
or U18086 (N_18086,N_17750,N_17840);
xnor U18087 (N_18087,N_17873,N_17877);
xnor U18088 (N_18088,N_17686,N_17754);
and U18089 (N_18089,N_17683,N_17972);
xor U18090 (N_18090,N_17605,N_17757);
nor U18091 (N_18091,N_17838,N_17885);
nor U18092 (N_18092,N_17949,N_17711);
and U18093 (N_18093,N_17841,N_17706);
nand U18094 (N_18094,N_17688,N_17990);
and U18095 (N_18095,N_17762,N_17975);
nor U18096 (N_18096,N_17705,N_17638);
xnor U18097 (N_18097,N_17870,N_17921);
nor U18098 (N_18098,N_17968,N_17655);
and U18099 (N_18099,N_17928,N_17782);
nor U18100 (N_18100,N_17734,N_17971);
nand U18101 (N_18101,N_17978,N_17767);
nand U18102 (N_18102,N_17772,N_17960);
xor U18103 (N_18103,N_17994,N_17914);
nor U18104 (N_18104,N_17792,N_17636);
nor U18105 (N_18105,N_17886,N_17640);
and U18106 (N_18106,N_17958,N_17882);
and U18107 (N_18107,N_17778,N_17620);
and U18108 (N_18108,N_17817,N_17728);
or U18109 (N_18109,N_17671,N_17713);
nand U18110 (N_18110,N_17608,N_17680);
xnor U18111 (N_18111,N_17985,N_17771);
or U18112 (N_18112,N_17759,N_17818);
nor U18113 (N_18113,N_17839,N_17632);
xnor U18114 (N_18114,N_17852,N_17678);
or U18115 (N_18115,N_17731,N_17630);
and U18116 (N_18116,N_17610,N_17718);
xnor U18117 (N_18117,N_17998,N_17761);
or U18118 (N_18118,N_17689,N_17777);
or U18119 (N_18119,N_17658,N_17969);
xor U18120 (N_18120,N_17844,N_17875);
nand U18121 (N_18121,N_17649,N_17868);
or U18122 (N_18122,N_17900,N_17633);
xor U18123 (N_18123,N_17973,N_17745);
and U18124 (N_18124,N_17933,N_17824);
and U18125 (N_18125,N_17790,N_17899);
nor U18126 (N_18126,N_17664,N_17809);
nor U18127 (N_18127,N_17611,N_17865);
and U18128 (N_18128,N_17724,N_17880);
and U18129 (N_18129,N_17793,N_17766);
xnor U18130 (N_18130,N_17674,N_17922);
nand U18131 (N_18131,N_17670,N_17942);
and U18132 (N_18132,N_17805,N_17827);
nand U18133 (N_18133,N_17834,N_17692);
xor U18134 (N_18134,N_17672,N_17826);
and U18135 (N_18135,N_17996,N_17895);
or U18136 (N_18136,N_17910,N_17850);
xor U18137 (N_18137,N_17691,N_17799);
and U18138 (N_18138,N_17696,N_17931);
nand U18139 (N_18139,N_17967,N_17853);
nand U18140 (N_18140,N_17897,N_17667);
xnor U18141 (N_18141,N_17889,N_17951);
nor U18142 (N_18142,N_17955,N_17637);
xor U18143 (N_18143,N_17729,N_17848);
nand U18144 (N_18144,N_17883,N_17776);
and U18145 (N_18145,N_17867,N_17800);
nand U18146 (N_18146,N_17685,N_17828);
nor U18147 (N_18147,N_17628,N_17736);
nor U18148 (N_18148,N_17803,N_17992);
nor U18149 (N_18149,N_17733,N_17950);
and U18150 (N_18150,N_17755,N_17927);
or U18151 (N_18151,N_17923,N_17917);
or U18152 (N_18152,N_17737,N_17920);
and U18153 (N_18153,N_17704,N_17749);
nand U18154 (N_18154,N_17965,N_17944);
nand U18155 (N_18155,N_17864,N_17811);
nor U18156 (N_18156,N_17687,N_17634);
nor U18157 (N_18157,N_17663,N_17845);
nand U18158 (N_18158,N_17623,N_17719);
and U18159 (N_18159,N_17825,N_17821);
and U18160 (N_18160,N_17607,N_17717);
nor U18161 (N_18161,N_17831,N_17721);
xnor U18162 (N_18162,N_17716,N_17795);
and U18163 (N_18163,N_17808,N_17983);
and U18164 (N_18164,N_17650,N_17614);
nor U18165 (N_18165,N_17819,N_17849);
or U18166 (N_18166,N_17690,N_17715);
xor U18167 (N_18167,N_17801,N_17806);
nor U18168 (N_18168,N_17962,N_17906);
xnor U18169 (N_18169,N_17697,N_17970);
xnor U18170 (N_18170,N_17791,N_17741);
nand U18171 (N_18171,N_17902,N_17982);
xnor U18172 (N_18172,N_17707,N_17918);
nand U18173 (N_18173,N_17622,N_17846);
xnor U18174 (N_18174,N_17642,N_17976);
nand U18175 (N_18175,N_17752,N_17963);
xnor U18176 (N_18176,N_17646,N_17893);
nor U18177 (N_18177,N_17662,N_17934);
xnor U18178 (N_18178,N_17702,N_17669);
xnor U18179 (N_18179,N_17859,N_17740);
nand U18180 (N_18180,N_17939,N_17639);
xor U18181 (N_18181,N_17919,N_17876);
or U18182 (N_18182,N_17661,N_17984);
and U18183 (N_18183,N_17742,N_17780);
xor U18184 (N_18184,N_17816,N_17714);
or U18185 (N_18185,N_17807,N_17905);
and U18186 (N_18186,N_17999,N_17675);
xnor U18187 (N_18187,N_17665,N_17966);
xor U18188 (N_18188,N_17991,N_17656);
nor U18189 (N_18189,N_17651,N_17925);
and U18190 (N_18190,N_17676,N_17952);
nor U18191 (N_18191,N_17896,N_17989);
nand U18192 (N_18192,N_17836,N_17624);
or U18193 (N_18193,N_17872,N_17835);
nand U18194 (N_18194,N_17760,N_17802);
or U18195 (N_18195,N_17869,N_17698);
nor U18196 (N_18196,N_17612,N_17603);
nand U18197 (N_18197,N_17789,N_17643);
nor U18198 (N_18198,N_17700,N_17619);
xnor U18199 (N_18199,N_17798,N_17709);
or U18200 (N_18200,N_17718,N_17946);
and U18201 (N_18201,N_17630,N_17766);
nor U18202 (N_18202,N_17738,N_17880);
and U18203 (N_18203,N_17771,N_17961);
nor U18204 (N_18204,N_17920,N_17672);
or U18205 (N_18205,N_17775,N_17949);
and U18206 (N_18206,N_17954,N_17641);
xnor U18207 (N_18207,N_17684,N_17716);
nor U18208 (N_18208,N_17745,N_17721);
xnor U18209 (N_18209,N_17921,N_17992);
xnor U18210 (N_18210,N_17715,N_17883);
nor U18211 (N_18211,N_17726,N_17926);
nor U18212 (N_18212,N_17872,N_17787);
xor U18213 (N_18213,N_17746,N_17843);
nor U18214 (N_18214,N_17701,N_17870);
and U18215 (N_18215,N_17854,N_17793);
or U18216 (N_18216,N_17769,N_17699);
nand U18217 (N_18217,N_17716,N_17780);
and U18218 (N_18218,N_17726,N_17864);
xnor U18219 (N_18219,N_17874,N_17649);
nor U18220 (N_18220,N_17777,N_17917);
xor U18221 (N_18221,N_17963,N_17785);
and U18222 (N_18222,N_17970,N_17926);
nor U18223 (N_18223,N_17749,N_17674);
xnor U18224 (N_18224,N_17898,N_17719);
nor U18225 (N_18225,N_17649,N_17728);
and U18226 (N_18226,N_17864,N_17898);
or U18227 (N_18227,N_17970,N_17640);
or U18228 (N_18228,N_17796,N_17963);
xor U18229 (N_18229,N_17689,N_17679);
nand U18230 (N_18230,N_17931,N_17800);
nor U18231 (N_18231,N_17878,N_17977);
xor U18232 (N_18232,N_17874,N_17745);
xnor U18233 (N_18233,N_17986,N_17616);
or U18234 (N_18234,N_17602,N_17905);
nor U18235 (N_18235,N_17639,N_17716);
or U18236 (N_18236,N_17880,N_17772);
nor U18237 (N_18237,N_17793,N_17749);
nor U18238 (N_18238,N_17678,N_17707);
nor U18239 (N_18239,N_17801,N_17615);
nand U18240 (N_18240,N_17955,N_17880);
or U18241 (N_18241,N_17618,N_17922);
nor U18242 (N_18242,N_17987,N_17779);
nand U18243 (N_18243,N_17744,N_17904);
nor U18244 (N_18244,N_17864,N_17660);
and U18245 (N_18245,N_17605,N_17820);
xnor U18246 (N_18246,N_17646,N_17672);
and U18247 (N_18247,N_17919,N_17851);
xor U18248 (N_18248,N_17608,N_17908);
nand U18249 (N_18249,N_17780,N_17705);
nand U18250 (N_18250,N_17699,N_17806);
nor U18251 (N_18251,N_17929,N_17630);
xnor U18252 (N_18252,N_17726,N_17737);
and U18253 (N_18253,N_17685,N_17839);
or U18254 (N_18254,N_17838,N_17977);
xor U18255 (N_18255,N_17619,N_17817);
xor U18256 (N_18256,N_17951,N_17804);
nand U18257 (N_18257,N_17971,N_17697);
and U18258 (N_18258,N_17920,N_17680);
and U18259 (N_18259,N_17991,N_17877);
and U18260 (N_18260,N_17750,N_17863);
or U18261 (N_18261,N_17618,N_17839);
and U18262 (N_18262,N_17670,N_17812);
and U18263 (N_18263,N_17786,N_17720);
nor U18264 (N_18264,N_17631,N_17790);
and U18265 (N_18265,N_17743,N_17614);
nand U18266 (N_18266,N_17842,N_17703);
and U18267 (N_18267,N_17979,N_17755);
nor U18268 (N_18268,N_17697,N_17796);
nor U18269 (N_18269,N_17816,N_17851);
xnor U18270 (N_18270,N_17920,N_17994);
nand U18271 (N_18271,N_17716,N_17872);
xor U18272 (N_18272,N_17729,N_17885);
xor U18273 (N_18273,N_17626,N_17845);
nand U18274 (N_18274,N_17963,N_17670);
and U18275 (N_18275,N_17885,N_17795);
or U18276 (N_18276,N_17967,N_17893);
or U18277 (N_18277,N_17788,N_17850);
or U18278 (N_18278,N_17745,N_17848);
xor U18279 (N_18279,N_17749,N_17611);
nand U18280 (N_18280,N_17790,N_17874);
nand U18281 (N_18281,N_17985,N_17742);
xor U18282 (N_18282,N_17770,N_17910);
nor U18283 (N_18283,N_17640,N_17767);
and U18284 (N_18284,N_17606,N_17876);
nor U18285 (N_18285,N_17661,N_17794);
xor U18286 (N_18286,N_17862,N_17839);
nand U18287 (N_18287,N_17908,N_17764);
nand U18288 (N_18288,N_17621,N_17812);
nor U18289 (N_18289,N_17764,N_17821);
or U18290 (N_18290,N_17840,N_17742);
nor U18291 (N_18291,N_17744,N_17676);
nor U18292 (N_18292,N_17998,N_17695);
nand U18293 (N_18293,N_17628,N_17884);
or U18294 (N_18294,N_17744,N_17662);
nand U18295 (N_18295,N_17663,N_17696);
nand U18296 (N_18296,N_17653,N_17792);
or U18297 (N_18297,N_17880,N_17982);
nor U18298 (N_18298,N_17978,N_17891);
xor U18299 (N_18299,N_17990,N_17671);
or U18300 (N_18300,N_17703,N_17911);
xor U18301 (N_18301,N_17877,N_17829);
and U18302 (N_18302,N_17726,N_17654);
xor U18303 (N_18303,N_17932,N_17641);
nand U18304 (N_18304,N_17729,N_17793);
and U18305 (N_18305,N_17739,N_17986);
xnor U18306 (N_18306,N_17860,N_17931);
nand U18307 (N_18307,N_17722,N_17764);
nand U18308 (N_18308,N_17720,N_17953);
and U18309 (N_18309,N_17798,N_17879);
or U18310 (N_18310,N_17940,N_17928);
xnor U18311 (N_18311,N_17664,N_17703);
xnor U18312 (N_18312,N_17914,N_17806);
nand U18313 (N_18313,N_17984,N_17605);
or U18314 (N_18314,N_17726,N_17766);
nand U18315 (N_18315,N_17783,N_17818);
nor U18316 (N_18316,N_17653,N_17975);
and U18317 (N_18317,N_17984,N_17692);
or U18318 (N_18318,N_17600,N_17713);
or U18319 (N_18319,N_17703,N_17808);
xnor U18320 (N_18320,N_17862,N_17856);
nand U18321 (N_18321,N_17604,N_17792);
xnor U18322 (N_18322,N_17906,N_17689);
xor U18323 (N_18323,N_17611,N_17754);
nand U18324 (N_18324,N_17734,N_17988);
and U18325 (N_18325,N_17780,N_17609);
and U18326 (N_18326,N_17948,N_17605);
xor U18327 (N_18327,N_17819,N_17737);
and U18328 (N_18328,N_17699,N_17748);
nand U18329 (N_18329,N_17904,N_17959);
nand U18330 (N_18330,N_17783,N_17724);
nand U18331 (N_18331,N_17839,N_17962);
nand U18332 (N_18332,N_17796,N_17623);
and U18333 (N_18333,N_17906,N_17736);
nand U18334 (N_18334,N_17650,N_17920);
and U18335 (N_18335,N_17637,N_17919);
nand U18336 (N_18336,N_17767,N_17650);
and U18337 (N_18337,N_17900,N_17639);
and U18338 (N_18338,N_17985,N_17702);
nand U18339 (N_18339,N_17958,N_17982);
xnor U18340 (N_18340,N_17705,N_17987);
and U18341 (N_18341,N_17926,N_17958);
or U18342 (N_18342,N_17891,N_17811);
nand U18343 (N_18343,N_17705,N_17682);
nor U18344 (N_18344,N_17768,N_17969);
and U18345 (N_18345,N_17946,N_17831);
nand U18346 (N_18346,N_17911,N_17805);
nor U18347 (N_18347,N_17698,N_17769);
nand U18348 (N_18348,N_17996,N_17861);
nor U18349 (N_18349,N_17738,N_17864);
and U18350 (N_18350,N_17747,N_17969);
nand U18351 (N_18351,N_17769,N_17810);
nor U18352 (N_18352,N_17705,N_17918);
or U18353 (N_18353,N_17878,N_17624);
nand U18354 (N_18354,N_17784,N_17944);
nor U18355 (N_18355,N_17623,N_17978);
xnor U18356 (N_18356,N_17647,N_17629);
xnor U18357 (N_18357,N_17871,N_17696);
or U18358 (N_18358,N_17732,N_17966);
nor U18359 (N_18359,N_17672,N_17844);
or U18360 (N_18360,N_17876,N_17624);
xor U18361 (N_18361,N_17940,N_17753);
or U18362 (N_18362,N_17685,N_17631);
xnor U18363 (N_18363,N_17977,N_17656);
xor U18364 (N_18364,N_17825,N_17836);
nor U18365 (N_18365,N_17959,N_17793);
nand U18366 (N_18366,N_17690,N_17766);
or U18367 (N_18367,N_17878,N_17764);
xnor U18368 (N_18368,N_17733,N_17945);
nand U18369 (N_18369,N_17972,N_17923);
nor U18370 (N_18370,N_17741,N_17898);
nor U18371 (N_18371,N_17878,N_17718);
nor U18372 (N_18372,N_17926,N_17725);
or U18373 (N_18373,N_17911,N_17939);
or U18374 (N_18374,N_17759,N_17651);
xor U18375 (N_18375,N_17845,N_17816);
nor U18376 (N_18376,N_17797,N_17961);
and U18377 (N_18377,N_17958,N_17738);
nand U18378 (N_18378,N_17898,N_17809);
xnor U18379 (N_18379,N_17817,N_17870);
nor U18380 (N_18380,N_17754,N_17636);
and U18381 (N_18381,N_17601,N_17643);
nor U18382 (N_18382,N_17728,N_17915);
nor U18383 (N_18383,N_17847,N_17723);
or U18384 (N_18384,N_17767,N_17803);
xnor U18385 (N_18385,N_17713,N_17786);
or U18386 (N_18386,N_17717,N_17898);
nor U18387 (N_18387,N_17726,N_17881);
nor U18388 (N_18388,N_17964,N_17898);
nand U18389 (N_18389,N_17621,N_17869);
and U18390 (N_18390,N_17714,N_17970);
nand U18391 (N_18391,N_17728,N_17726);
nor U18392 (N_18392,N_17943,N_17650);
xor U18393 (N_18393,N_17801,N_17881);
xnor U18394 (N_18394,N_17707,N_17973);
or U18395 (N_18395,N_17892,N_17816);
or U18396 (N_18396,N_17858,N_17753);
xnor U18397 (N_18397,N_17672,N_17634);
nor U18398 (N_18398,N_17916,N_17878);
nor U18399 (N_18399,N_17907,N_17660);
or U18400 (N_18400,N_18184,N_18375);
nand U18401 (N_18401,N_18220,N_18359);
nand U18402 (N_18402,N_18307,N_18104);
nor U18403 (N_18403,N_18042,N_18009);
nor U18404 (N_18404,N_18033,N_18177);
nor U18405 (N_18405,N_18024,N_18109);
nand U18406 (N_18406,N_18214,N_18153);
and U18407 (N_18407,N_18320,N_18158);
nor U18408 (N_18408,N_18298,N_18193);
or U18409 (N_18409,N_18358,N_18037);
and U18410 (N_18410,N_18395,N_18074);
or U18411 (N_18411,N_18336,N_18078);
nand U18412 (N_18412,N_18278,N_18082);
or U18413 (N_18413,N_18092,N_18079);
nor U18414 (N_18414,N_18056,N_18303);
or U18415 (N_18415,N_18094,N_18151);
and U18416 (N_18416,N_18199,N_18321);
nor U18417 (N_18417,N_18051,N_18241);
and U18418 (N_18418,N_18156,N_18299);
nand U18419 (N_18419,N_18260,N_18367);
nor U18420 (N_18420,N_18398,N_18050);
and U18421 (N_18421,N_18185,N_18253);
nor U18422 (N_18422,N_18231,N_18378);
nor U18423 (N_18423,N_18100,N_18120);
or U18424 (N_18424,N_18314,N_18179);
and U18425 (N_18425,N_18144,N_18101);
xnor U18426 (N_18426,N_18300,N_18129);
or U18427 (N_18427,N_18136,N_18066);
or U18428 (N_18428,N_18102,N_18125);
nand U18429 (N_18429,N_18067,N_18005);
xnor U18430 (N_18430,N_18335,N_18275);
and U18431 (N_18431,N_18325,N_18372);
or U18432 (N_18432,N_18259,N_18175);
xnor U18433 (N_18433,N_18306,N_18244);
nand U18434 (N_18434,N_18392,N_18202);
xor U18435 (N_18435,N_18097,N_18386);
xor U18436 (N_18436,N_18270,N_18046);
nor U18437 (N_18437,N_18208,N_18366);
nor U18438 (N_18438,N_18238,N_18133);
xnor U18439 (N_18439,N_18237,N_18107);
and U18440 (N_18440,N_18119,N_18317);
and U18441 (N_18441,N_18030,N_18025);
or U18442 (N_18442,N_18217,N_18164);
nor U18443 (N_18443,N_18354,N_18131);
nand U18444 (N_18444,N_18155,N_18069);
or U18445 (N_18445,N_18391,N_18165);
nor U18446 (N_18446,N_18178,N_18085);
xor U18447 (N_18447,N_18224,N_18264);
or U18448 (N_18448,N_18341,N_18140);
xor U18449 (N_18449,N_18271,N_18022);
nor U18450 (N_18450,N_18377,N_18373);
nand U18451 (N_18451,N_18138,N_18351);
nor U18452 (N_18452,N_18139,N_18044);
or U18453 (N_18453,N_18269,N_18363);
and U18454 (N_18454,N_18173,N_18329);
nor U18455 (N_18455,N_18200,N_18226);
xnor U18456 (N_18456,N_18334,N_18349);
nor U18457 (N_18457,N_18023,N_18362);
nand U18458 (N_18458,N_18324,N_18145);
nand U18459 (N_18459,N_18286,N_18028);
nor U18460 (N_18460,N_18014,N_18243);
or U18461 (N_18461,N_18262,N_18338);
nor U18462 (N_18462,N_18087,N_18390);
nand U18463 (N_18463,N_18147,N_18057);
xor U18464 (N_18464,N_18083,N_18365);
nand U18465 (N_18465,N_18121,N_18149);
nand U18466 (N_18466,N_18016,N_18148);
or U18467 (N_18467,N_18076,N_18397);
xnor U18468 (N_18468,N_18326,N_18291);
or U18469 (N_18469,N_18090,N_18382);
nor U18470 (N_18470,N_18011,N_18393);
or U18471 (N_18471,N_18127,N_18146);
and U18472 (N_18472,N_18080,N_18361);
and U18473 (N_18473,N_18331,N_18160);
and U18474 (N_18474,N_18305,N_18254);
or U18475 (N_18475,N_18252,N_18195);
nor U18476 (N_18476,N_18152,N_18013);
nand U18477 (N_18477,N_18181,N_18060);
nand U18478 (N_18478,N_18190,N_18111);
or U18479 (N_18479,N_18239,N_18012);
xnor U18480 (N_18480,N_18255,N_18123);
xnor U18481 (N_18481,N_18360,N_18137);
xor U18482 (N_18482,N_18285,N_18348);
nand U18483 (N_18483,N_18293,N_18374);
xnor U18484 (N_18484,N_18273,N_18343);
and U18485 (N_18485,N_18188,N_18384);
and U18486 (N_18486,N_18059,N_18337);
and U18487 (N_18487,N_18205,N_18388);
nor U18488 (N_18488,N_18265,N_18112);
or U18489 (N_18489,N_18268,N_18313);
nand U18490 (N_18490,N_18276,N_18197);
nand U18491 (N_18491,N_18026,N_18055);
xor U18492 (N_18492,N_18126,N_18210);
nor U18493 (N_18493,N_18062,N_18061);
xnor U18494 (N_18494,N_18345,N_18170);
nor U18495 (N_18495,N_18150,N_18098);
xnor U18496 (N_18496,N_18143,N_18093);
nand U18497 (N_18497,N_18027,N_18342);
and U18498 (N_18498,N_18357,N_18333);
nor U18499 (N_18499,N_18376,N_18000);
nor U18500 (N_18500,N_18118,N_18004);
and U18501 (N_18501,N_18394,N_18047);
nand U18502 (N_18502,N_18221,N_18154);
nand U18503 (N_18503,N_18058,N_18369);
and U18504 (N_18504,N_18176,N_18304);
nand U18505 (N_18505,N_18236,N_18251);
xnor U18506 (N_18506,N_18261,N_18172);
or U18507 (N_18507,N_18308,N_18171);
nor U18508 (N_18508,N_18387,N_18385);
and U18509 (N_18509,N_18319,N_18396);
xnor U18510 (N_18510,N_18364,N_18018);
nor U18511 (N_18511,N_18032,N_18266);
and U18512 (N_18512,N_18350,N_18234);
and U18513 (N_18513,N_18168,N_18029);
and U18514 (N_18514,N_18006,N_18064);
nor U18515 (N_18515,N_18211,N_18379);
nor U18516 (N_18516,N_18043,N_18277);
nor U18517 (N_18517,N_18183,N_18368);
or U18518 (N_18518,N_18225,N_18174);
and U18519 (N_18519,N_18216,N_18212);
nor U18520 (N_18520,N_18115,N_18247);
or U18521 (N_18521,N_18040,N_18162);
nor U18522 (N_18522,N_18302,N_18035);
xor U18523 (N_18523,N_18089,N_18399);
nor U18524 (N_18524,N_18157,N_18292);
xnor U18525 (N_18525,N_18381,N_18203);
and U18526 (N_18526,N_18034,N_18322);
and U18527 (N_18527,N_18191,N_18290);
and U18528 (N_18528,N_18287,N_18383);
and U18529 (N_18529,N_18167,N_18103);
nand U18530 (N_18530,N_18257,N_18219);
and U18531 (N_18531,N_18134,N_18207);
and U18532 (N_18532,N_18105,N_18249);
nor U18533 (N_18533,N_18288,N_18015);
nand U18534 (N_18534,N_18370,N_18189);
and U18535 (N_18535,N_18311,N_18073);
xnor U18536 (N_18536,N_18021,N_18213);
or U18537 (N_18537,N_18130,N_18049);
xor U18538 (N_18538,N_18201,N_18279);
and U18539 (N_18539,N_18301,N_18113);
nand U18540 (N_18540,N_18267,N_18256);
or U18541 (N_18541,N_18008,N_18124);
nor U18542 (N_18542,N_18346,N_18235);
or U18543 (N_18543,N_18328,N_18096);
and U18544 (N_18544,N_18116,N_18280);
or U18545 (N_18545,N_18187,N_18371);
nand U18546 (N_18546,N_18084,N_18297);
or U18547 (N_18547,N_18215,N_18258);
nand U18548 (N_18548,N_18229,N_18233);
nand U18549 (N_18549,N_18063,N_18209);
and U18550 (N_18550,N_18091,N_18281);
or U18551 (N_18551,N_18099,N_18355);
or U18552 (N_18552,N_18196,N_18204);
or U18553 (N_18553,N_18128,N_18206);
and U18554 (N_18554,N_18135,N_18077);
nand U18555 (N_18555,N_18053,N_18114);
or U18556 (N_18556,N_18352,N_18347);
and U18557 (N_18557,N_18036,N_18070);
or U18558 (N_18558,N_18192,N_18296);
nand U18559 (N_18559,N_18295,N_18380);
xor U18560 (N_18560,N_18072,N_18327);
nand U18561 (N_18561,N_18356,N_18010);
and U18562 (N_18562,N_18065,N_18017);
or U18563 (N_18563,N_18240,N_18106);
nor U18564 (N_18564,N_18223,N_18054);
xnor U18565 (N_18565,N_18052,N_18310);
or U18566 (N_18566,N_18117,N_18242);
nand U18567 (N_18567,N_18272,N_18071);
nand U18568 (N_18568,N_18284,N_18274);
nand U18569 (N_18569,N_18330,N_18194);
nor U18570 (N_18570,N_18166,N_18228);
nor U18571 (N_18571,N_18163,N_18161);
and U18572 (N_18572,N_18389,N_18002);
or U18573 (N_18573,N_18289,N_18186);
xnor U18574 (N_18574,N_18283,N_18250);
or U18575 (N_18575,N_18282,N_18068);
xor U18576 (N_18576,N_18142,N_18182);
nor U18577 (N_18577,N_18020,N_18230);
nor U18578 (N_18578,N_18110,N_18003);
nor U18579 (N_18579,N_18169,N_18086);
xor U18580 (N_18580,N_18232,N_18218);
nor U18581 (N_18581,N_18316,N_18344);
and U18582 (N_18582,N_18007,N_18227);
nor U18583 (N_18583,N_18180,N_18039);
nor U18584 (N_18584,N_18001,N_18108);
and U18585 (N_18585,N_18248,N_18353);
nor U18586 (N_18586,N_18088,N_18081);
nand U18587 (N_18587,N_18245,N_18141);
nand U18588 (N_18588,N_18323,N_18019);
xnor U18589 (N_18589,N_18095,N_18122);
or U18590 (N_18590,N_18309,N_18315);
and U18591 (N_18591,N_18045,N_18159);
and U18592 (N_18592,N_18198,N_18075);
xor U18593 (N_18593,N_18041,N_18294);
or U18594 (N_18594,N_18312,N_18031);
nand U18595 (N_18595,N_18038,N_18246);
xor U18596 (N_18596,N_18263,N_18318);
or U18597 (N_18597,N_18222,N_18332);
or U18598 (N_18598,N_18339,N_18048);
xor U18599 (N_18599,N_18340,N_18132);
or U18600 (N_18600,N_18134,N_18016);
and U18601 (N_18601,N_18054,N_18253);
xnor U18602 (N_18602,N_18234,N_18099);
and U18603 (N_18603,N_18256,N_18166);
xor U18604 (N_18604,N_18292,N_18372);
xor U18605 (N_18605,N_18074,N_18082);
nand U18606 (N_18606,N_18200,N_18359);
or U18607 (N_18607,N_18335,N_18273);
xnor U18608 (N_18608,N_18034,N_18002);
xor U18609 (N_18609,N_18158,N_18133);
nand U18610 (N_18610,N_18372,N_18262);
xnor U18611 (N_18611,N_18283,N_18047);
and U18612 (N_18612,N_18274,N_18082);
nand U18613 (N_18613,N_18094,N_18239);
or U18614 (N_18614,N_18059,N_18069);
xor U18615 (N_18615,N_18032,N_18279);
nor U18616 (N_18616,N_18372,N_18094);
nand U18617 (N_18617,N_18302,N_18358);
nor U18618 (N_18618,N_18390,N_18242);
and U18619 (N_18619,N_18190,N_18142);
and U18620 (N_18620,N_18146,N_18016);
nor U18621 (N_18621,N_18323,N_18037);
nor U18622 (N_18622,N_18123,N_18376);
nand U18623 (N_18623,N_18009,N_18386);
nor U18624 (N_18624,N_18377,N_18136);
or U18625 (N_18625,N_18035,N_18059);
nand U18626 (N_18626,N_18303,N_18354);
or U18627 (N_18627,N_18118,N_18148);
xnor U18628 (N_18628,N_18027,N_18090);
or U18629 (N_18629,N_18154,N_18348);
nor U18630 (N_18630,N_18116,N_18137);
nand U18631 (N_18631,N_18384,N_18054);
and U18632 (N_18632,N_18299,N_18142);
or U18633 (N_18633,N_18297,N_18382);
nor U18634 (N_18634,N_18071,N_18138);
or U18635 (N_18635,N_18045,N_18239);
and U18636 (N_18636,N_18312,N_18134);
nand U18637 (N_18637,N_18259,N_18295);
and U18638 (N_18638,N_18072,N_18344);
nand U18639 (N_18639,N_18134,N_18372);
nand U18640 (N_18640,N_18249,N_18357);
or U18641 (N_18641,N_18299,N_18090);
and U18642 (N_18642,N_18268,N_18393);
xor U18643 (N_18643,N_18338,N_18165);
xor U18644 (N_18644,N_18116,N_18237);
or U18645 (N_18645,N_18200,N_18125);
nor U18646 (N_18646,N_18251,N_18152);
nand U18647 (N_18647,N_18178,N_18144);
and U18648 (N_18648,N_18151,N_18380);
nor U18649 (N_18649,N_18203,N_18362);
and U18650 (N_18650,N_18381,N_18083);
or U18651 (N_18651,N_18384,N_18022);
xor U18652 (N_18652,N_18040,N_18353);
xnor U18653 (N_18653,N_18171,N_18367);
and U18654 (N_18654,N_18203,N_18245);
nand U18655 (N_18655,N_18337,N_18068);
xnor U18656 (N_18656,N_18112,N_18175);
and U18657 (N_18657,N_18061,N_18231);
nor U18658 (N_18658,N_18132,N_18026);
nor U18659 (N_18659,N_18367,N_18293);
or U18660 (N_18660,N_18133,N_18295);
nor U18661 (N_18661,N_18271,N_18097);
and U18662 (N_18662,N_18053,N_18090);
and U18663 (N_18663,N_18053,N_18139);
nor U18664 (N_18664,N_18162,N_18114);
nand U18665 (N_18665,N_18372,N_18070);
nor U18666 (N_18666,N_18207,N_18176);
and U18667 (N_18667,N_18346,N_18270);
or U18668 (N_18668,N_18342,N_18286);
or U18669 (N_18669,N_18376,N_18228);
nand U18670 (N_18670,N_18113,N_18256);
xor U18671 (N_18671,N_18172,N_18292);
nor U18672 (N_18672,N_18237,N_18177);
nand U18673 (N_18673,N_18129,N_18042);
nand U18674 (N_18674,N_18145,N_18029);
xor U18675 (N_18675,N_18000,N_18132);
or U18676 (N_18676,N_18297,N_18187);
and U18677 (N_18677,N_18319,N_18118);
nand U18678 (N_18678,N_18332,N_18093);
xor U18679 (N_18679,N_18270,N_18014);
nor U18680 (N_18680,N_18024,N_18190);
nand U18681 (N_18681,N_18310,N_18323);
and U18682 (N_18682,N_18031,N_18275);
xnor U18683 (N_18683,N_18205,N_18370);
xnor U18684 (N_18684,N_18339,N_18085);
nor U18685 (N_18685,N_18256,N_18058);
nor U18686 (N_18686,N_18170,N_18236);
nor U18687 (N_18687,N_18049,N_18031);
xor U18688 (N_18688,N_18127,N_18112);
xor U18689 (N_18689,N_18174,N_18364);
and U18690 (N_18690,N_18317,N_18273);
or U18691 (N_18691,N_18368,N_18042);
or U18692 (N_18692,N_18016,N_18093);
nor U18693 (N_18693,N_18153,N_18155);
nand U18694 (N_18694,N_18306,N_18233);
nor U18695 (N_18695,N_18185,N_18056);
and U18696 (N_18696,N_18319,N_18111);
and U18697 (N_18697,N_18209,N_18179);
or U18698 (N_18698,N_18221,N_18366);
xnor U18699 (N_18699,N_18267,N_18140);
nand U18700 (N_18700,N_18186,N_18359);
and U18701 (N_18701,N_18196,N_18361);
and U18702 (N_18702,N_18259,N_18138);
and U18703 (N_18703,N_18024,N_18194);
and U18704 (N_18704,N_18062,N_18385);
nand U18705 (N_18705,N_18017,N_18136);
nor U18706 (N_18706,N_18042,N_18394);
nor U18707 (N_18707,N_18215,N_18028);
nand U18708 (N_18708,N_18003,N_18001);
and U18709 (N_18709,N_18013,N_18003);
xor U18710 (N_18710,N_18152,N_18239);
nand U18711 (N_18711,N_18197,N_18220);
or U18712 (N_18712,N_18026,N_18282);
nor U18713 (N_18713,N_18323,N_18314);
or U18714 (N_18714,N_18079,N_18322);
and U18715 (N_18715,N_18360,N_18014);
xnor U18716 (N_18716,N_18004,N_18198);
nor U18717 (N_18717,N_18238,N_18139);
nor U18718 (N_18718,N_18357,N_18116);
nand U18719 (N_18719,N_18290,N_18382);
xor U18720 (N_18720,N_18124,N_18355);
or U18721 (N_18721,N_18040,N_18227);
and U18722 (N_18722,N_18019,N_18398);
or U18723 (N_18723,N_18219,N_18084);
nor U18724 (N_18724,N_18236,N_18341);
nand U18725 (N_18725,N_18042,N_18281);
nor U18726 (N_18726,N_18225,N_18346);
and U18727 (N_18727,N_18248,N_18314);
nor U18728 (N_18728,N_18257,N_18084);
nor U18729 (N_18729,N_18293,N_18112);
or U18730 (N_18730,N_18372,N_18137);
and U18731 (N_18731,N_18381,N_18073);
nor U18732 (N_18732,N_18086,N_18336);
nor U18733 (N_18733,N_18095,N_18323);
and U18734 (N_18734,N_18026,N_18081);
xor U18735 (N_18735,N_18194,N_18160);
nor U18736 (N_18736,N_18359,N_18052);
or U18737 (N_18737,N_18173,N_18197);
nor U18738 (N_18738,N_18080,N_18297);
or U18739 (N_18739,N_18319,N_18185);
xor U18740 (N_18740,N_18183,N_18152);
and U18741 (N_18741,N_18330,N_18181);
nand U18742 (N_18742,N_18351,N_18344);
xnor U18743 (N_18743,N_18218,N_18159);
or U18744 (N_18744,N_18116,N_18213);
or U18745 (N_18745,N_18324,N_18327);
or U18746 (N_18746,N_18117,N_18058);
xnor U18747 (N_18747,N_18114,N_18313);
nor U18748 (N_18748,N_18038,N_18021);
or U18749 (N_18749,N_18200,N_18091);
nand U18750 (N_18750,N_18228,N_18052);
xnor U18751 (N_18751,N_18117,N_18264);
xor U18752 (N_18752,N_18382,N_18362);
nor U18753 (N_18753,N_18007,N_18087);
xor U18754 (N_18754,N_18375,N_18349);
nor U18755 (N_18755,N_18052,N_18098);
or U18756 (N_18756,N_18065,N_18292);
nor U18757 (N_18757,N_18205,N_18082);
nand U18758 (N_18758,N_18004,N_18054);
and U18759 (N_18759,N_18188,N_18360);
nand U18760 (N_18760,N_18051,N_18068);
nor U18761 (N_18761,N_18268,N_18300);
and U18762 (N_18762,N_18169,N_18273);
or U18763 (N_18763,N_18206,N_18378);
nand U18764 (N_18764,N_18288,N_18002);
nand U18765 (N_18765,N_18204,N_18261);
and U18766 (N_18766,N_18301,N_18184);
nand U18767 (N_18767,N_18016,N_18264);
nor U18768 (N_18768,N_18142,N_18121);
nor U18769 (N_18769,N_18172,N_18397);
xnor U18770 (N_18770,N_18154,N_18303);
and U18771 (N_18771,N_18159,N_18022);
or U18772 (N_18772,N_18100,N_18385);
nor U18773 (N_18773,N_18218,N_18001);
or U18774 (N_18774,N_18189,N_18056);
xor U18775 (N_18775,N_18282,N_18120);
xnor U18776 (N_18776,N_18182,N_18289);
nand U18777 (N_18777,N_18176,N_18166);
nor U18778 (N_18778,N_18127,N_18084);
or U18779 (N_18779,N_18022,N_18305);
or U18780 (N_18780,N_18254,N_18045);
xnor U18781 (N_18781,N_18393,N_18343);
nor U18782 (N_18782,N_18127,N_18175);
nand U18783 (N_18783,N_18243,N_18078);
and U18784 (N_18784,N_18288,N_18378);
nor U18785 (N_18785,N_18250,N_18062);
and U18786 (N_18786,N_18019,N_18064);
xor U18787 (N_18787,N_18061,N_18282);
nand U18788 (N_18788,N_18399,N_18397);
or U18789 (N_18789,N_18121,N_18283);
and U18790 (N_18790,N_18340,N_18311);
or U18791 (N_18791,N_18357,N_18301);
or U18792 (N_18792,N_18057,N_18302);
nor U18793 (N_18793,N_18260,N_18188);
xor U18794 (N_18794,N_18230,N_18340);
nand U18795 (N_18795,N_18123,N_18303);
nor U18796 (N_18796,N_18198,N_18162);
nor U18797 (N_18797,N_18389,N_18127);
xor U18798 (N_18798,N_18150,N_18115);
nand U18799 (N_18799,N_18096,N_18132);
nand U18800 (N_18800,N_18413,N_18496);
nand U18801 (N_18801,N_18552,N_18776);
nand U18802 (N_18802,N_18597,N_18420);
xor U18803 (N_18803,N_18604,N_18679);
and U18804 (N_18804,N_18547,N_18755);
and U18805 (N_18805,N_18654,N_18521);
nor U18806 (N_18806,N_18467,N_18444);
xnor U18807 (N_18807,N_18516,N_18763);
nor U18808 (N_18808,N_18665,N_18466);
and U18809 (N_18809,N_18610,N_18422);
nand U18810 (N_18810,N_18515,N_18438);
nor U18811 (N_18811,N_18403,N_18781);
xnor U18812 (N_18812,N_18704,N_18684);
nor U18813 (N_18813,N_18450,N_18421);
or U18814 (N_18814,N_18626,N_18648);
and U18815 (N_18815,N_18465,N_18722);
nor U18816 (N_18816,N_18447,N_18631);
and U18817 (N_18817,N_18750,N_18771);
or U18818 (N_18818,N_18622,N_18678);
xor U18819 (N_18819,N_18479,N_18492);
nor U18820 (N_18820,N_18671,N_18502);
or U18821 (N_18821,N_18457,N_18688);
nand U18822 (N_18822,N_18498,N_18629);
xor U18823 (N_18823,N_18708,N_18746);
or U18824 (N_18824,N_18573,N_18605);
and U18825 (N_18825,N_18768,N_18402);
xor U18826 (N_18826,N_18484,N_18409);
nor U18827 (N_18827,N_18511,N_18675);
nor U18828 (N_18828,N_18408,N_18773);
or U18829 (N_18829,N_18764,N_18749);
or U18830 (N_18830,N_18545,N_18464);
and U18831 (N_18831,N_18461,N_18766);
xnor U18832 (N_18832,N_18485,N_18673);
nor U18833 (N_18833,N_18418,N_18714);
xnor U18834 (N_18834,N_18510,N_18655);
and U18835 (N_18835,N_18674,N_18400);
or U18836 (N_18836,N_18572,N_18682);
xnor U18837 (N_18837,N_18535,N_18579);
and U18838 (N_18838,N_18551,N_18434);
or U18839 (N_18839,N_18412,N_18627);
or U18840 (N_18840,N_18460,N_18612);
xor U18841 (N_18841,N_18554,N_18630);
and U18842 (N_18842,N_18735,N_18480);
or U18843 (N_18843,N_18454,N_18725);
and U18844 (N_18844,N_18401,N_18651);
nor U18845 (N_18845,N_18528,N_18715);
and U18846 (N_18846,N_18556,N_18497);
nor U18847 (N_18847,N_18690,N_18449);
xor U18848 (N_18848,N_18677,N_18570);
or U18849 (N_18849,N_18779,N_18659);
and U18850 (N_18850,N_18729,N_18649);
and U18851 (N_18851,N_18425,N_18482);
and U18852 (N_18852,N_18744,N_18531);
nor U18853 (N_18853,N_18711,N_18578);
and U18854 (N_18854,N_18529,N_18658);
nand U18855 (N_18855,N_18595,N_18685);
xnor U18856 (N_18856,N_18761,N_18488);
nor U18857 (N_18857,N_18797,N_18426);
xor U18858 (N_18858,N_18542,N_18562);
nor U18859 (N_18859,N_18698,N_18733);
nor U18860 (N_18860,N_18666,N_18693);
and U18861 (N_18861,N_18762,N_18724);
nand U18862 (N_18862,N_18726,N_18751);
nand U18863 (N_18863,N_18789,N_18441);
and U18864 (N_18864,N_18507,N_18536);
nand U18865 (N_18865,N_18534,N_18638);
and U18866 (N_18866,N_18526,N_18697);
nor U18867 (N_18867,N_18778,N_18608);
or U18868 (N_18868,N_18470,N_18676);
and U18869 (N_18869,N_18490,N_18427);
or U18870 (N_18870,N_18653,N_18472);
xnor U18871 (N_18871,N_18667,N_18481);
xor U18872 (N_18872,N_18474,N_18769);
xnor U18873 (N_18873,N_18601,N_18737);
xor U18874 (N_18874,N_18513,N_18491);
nor U18875 (N_18875,N_18709,N_18652);
xnor U18876 (N_18876,N_18719,N_18772);
nor U18877 (N_18877,N_18432,N_18512);
or U18878 (N_18878,N_18517,N_18743);
nor U18879 (N_18879,N_18431,N_18782);
xor U18880 (N_18880,N_18594,N_18723);
and U18881 (N_18881,N_18748,N_18456);
xor U18882 (N_18882,N_18643,N_18628);
xnor U18883 (N_18883,N_18641,N_18784);
or U18884 (N_18884,N_18646,N_18439);
and U18885 (N_18885,N_18523,N_18732);
or U18886 (N_18886,N_18742,N_18509);
or U18887 (N_18887,N_18462,N_18495);
or U18888 (N_18888,N_18463,N_18717);
xor U18889 (N_18889,N_18788,N_18741);
and U18890 (N_18890,N_18775,N_18691);
or U18891 (N_18891,N_18700,N_18642);
nand U18892 (N_18892,N_18696,N_18423);
nor U18893 (N_18893,N_18500,N_18670);
or U18894 (N_18894,N_18794,N_18455);
nand U18895 (N_18895,N_18720,N_18525);
xor U18896 (N_18896,N_18656,N_18428);
nand U18897 (N_18897,N_18745,N_18565);
xor U18898 (N_18898,N_18718,N_18406);
or U18899 (N_18899,N_18707,N_18616);
xor U18900 (N_18900,N_18633,N_18686);
xor U18901 (N_18901,N_18569,N_18543);
and U18902 (N_18902,N_18561,N_18581);
nand U18903 (N_18903,N_18692,N_18503);
nor U18904 (N_18904,N_18539,N_18681);
and U18905 (N_18905,N_18596,N_18792);
and U18906 (N_18906,N_18650,N_18560);
nand U18907 (N_18907,N_18548,N_18712);
or U18908 (N_18908,N_18527,N_18501);
and U18909 (N_18909,N_18756,N_18433);
xor U18910 (N_18910,N_18770,N_18524);
xor U18911 (N_18911,N_18533,N_18713);
nand U18912 (N_18912,N_18506,N_18430);
nor U18913 (N_18913,N_18519,N_18663);
and U18914 (N_18914,N_18760,N_18786);
xnor U18915 (N_18915,N_18669,N_18632);
nand U18916 (N_18916,N_18615,N_18623);
and U18917 (N_18917,N_18798,N_18473);
xor U18918 (N_18918,N_18793,N_18668);
xnor U18919 (N_18919,N_18494,N_18787);
nor U18920 (N_18920,N_18624,N_18514);
or U18921 (N_18921,N_18598,N_18419);
and U18922 (N_18922,N_18747,N_18574);
nor U18923 (N_18923,N_18404,N_18619);
or U18924 (N_18924,N_18532,N_18791);
or U18925 (N_18925,N_18695,N_18568);
nor U18926 (N_18926,N_18680,N_18589);
and U18927 (N_18927,N_18736,N_18607);
or U18928 (N_18928,N_18541,N_18540);
xnor U18929 (N_18929,N_18504,N_18505);
nand U18930 (N_18930,N_18443,N_18405);
and U18931 (N_18931,N_18731,N_18705);
nand U18932 (N_18932,N_18469,N_18647);
xor U18933 (N_18933,N_18437,N_18557);
nor U18934 (N_18934,N_18580,N_18618);
xor U18935 (N_18935,N_18739,N_18706);
or U18936 (N_18936,N_18699,N_18435);
and U18937 (N_18937,N_18458,N_18734);
and U18938 (N_18938,N_18774,N_18660);
and U18939 (N_18939,N_18687,N_18703);
nand U18940 (N_18940,N_18577,N_18661);
and U18941 (N_18941,N_18752,N_18783);
and U18942 (N_18942,N_18415,N_18520);
or U18943 (N_18943,N_18603,N_18702);
or U18944 (N_18944,N_18417,N_18489);
and U18945 (N_18945,N_18590,N_18446);
nand U18946 (N_18946,N_18440,N_18620);
or U18947 (N_18947,N_18617,N_18530);
or U18948 (N_18948,N_18586,N_18538);
nor U18949 (N_18949,N_18758,N_18799);
nor U18950 (N_18950,N_18411,N_18567);
or U18951 (N_18951,N_18635,N_18410);
or U18952 (N_18952,N_18710,N_18468);
or U18953 (N_18953,N_18478,N_18575);
or U18954 (N_18954,N_18727,N_18407);
or U18955 (N_18955,N_18716,N_18559);
or U18956 (N_18956,N_18599,N_18664);
nor U18957 (N_18957,N_18459,N_18765);
nor U18958 (N_18958,N_18471,N_18796);
nand U18959 (N_18959,N_18442,N_18644);
xor U18960 (N_18960,N_18721,N_18730);
xnor U18961 (N_18961,N_18592,N_18600);
or U18962 (N_18962,N_18740,N_18475);
nor U18963 (N_18963,N_18537,N_18553);
xor U18964 (N_18964,N_18753,N_18451);
or U18965 (N_18965,N_18564,N_18518);
or U18966 (N_18966,N_18728,N_18571);
nand U18967 (N_18967,N_18416,N_18445);
nor U18968 (N_18968,N_18499,N_18602);
or U18969 (N_18969,N_18453,N_18477);
nor U18970 (N_18970,N_18583,N_18587);
nand U18971 (N_18971,N_18544,N_18448);
xnor U18972 (N_18972,N_18585,N_18550);
or U18973 (N_18973,N_18672,N_18476);
and U18974 (N_18974,N_18613,N_18785);
xor U18975 (N_18975,N_18522,N_18645);
xor U18976 (N_18976,N_18609,N_18483);
or U18977 (N_18977,N_18639,N_18767);
and U18978 (N_18978,N_18584,N_18436);
or U18979 (N_18979,N_18689,N_18606);
xnor U18980 (N_18980,N_18625,N_18637);
or U18981 (N_18981,N_18738,N_18452);
xor U18982 (N_18982,N_18591,N_18780);
or U18983 (N_18983,N_18614,N_18757);
or U18984 (N_18984,N_18576,N_18508);
and U18985 (N_18985,N_18563,N_18662);
xnor U18986 (N_18986,N_18636,N_18754);
nand U18987 (N_18987,N_18640,N_18487);
and U18988 (N_18988,N_18566,N_18694);
xor U18989 (N_18989,N_18621,N_18414);
nor U18990 (N_18990,N_18493,N_18424);
nor U18991 (N_18991,N_18777,N_18795);
nor U18992 (N_18992,N_18759,N_18593);
or U18993 (N_18993,N_18588,N_18683);
nor U18994 (N_18994,N_18634,N_18657);
or U18995 (N_18995,N_18546,N_18549);
nand U18996 (N_18996,N_18611,N_18558);
or U18997 (N_18997,N_18582,N_18701);
nand U18998 (N_18998,N_18486,N_18429);
nand U18999 (N_18999,N_18790,N_18555);
nand U19000 (N_19000,N_18787,N_18757);
or U19001 (N_19001,N_18719,N_18591);
xor U19002 (N_19002,N_18408,N_18774);
nor U19003 (N_19003,N_18772,N_18587);
and U19004 (N_19004,N_18663,N_18736);
nand U19005 (N_19005,N_18589,N_18682);
and U19006 (N_19006,N_18575,N_18612);
or U19007 (N_19007,N_18626,N_18605);
or U19008 (N_19008,N_18453,N_18468);
xor U19009 (N_19009,N_18557,N_18461);
xnor U19010 (N_19010,N_18672,N_18634);
nand U19011 (N_19011,N_18403,N_18427);
nand U19012 (N_19012,N_18618,N_18441);
and U19013 (N_19013,N_18557,N_18645);
nor U19014 (N_19014,N_18490,N_18686);
xnor U19015 (N_19015,N_18698,N_18504);
xnor U19016 (N_19016,N_18570,N_18708);
nand U19017 (N_19017,N_18630,N_18616);
nor U19018 (N_19018,N_18495,N_18787);
nand U19019 (N_19019,N_18608,N_18702);
nand U19020 (N_19020,N_18564,N_18421);
nand U19021 (N_19021,N_18538,N_18400);
xor U19022 (N_19022,N_18591,N_18671);
or U19023 (N_19023,N_18737,N_18428);
xnor U19024 (N_19024,N_18673,N_18494);
xnor U19025 (N_19025,N_18449,N_18571);
xor U19026 (N_19026,N_18414,N_18570);
xnor U19027 (N_19027,N_18741,N_18508);
nor U19028 (N_19028,N_18481,N_18405);
or U19029 (N_19029,N_18546,N_18514);
xor U19030 (N_19030,N_18440,N_18436);
or U19031 (N_19031,N_18746,N_18713);
xor U19032 (N_19032,N_18521,N_18516);
nand U19033 (N_19033,N_18762,N_18630);
and U19034 (N_19034,N_18664,N_18532);
nand U19035 (N_19035,N_18651,N_18649);
xor U19036 (N_19036,N_18679,N_18509);
nor U19037 (N_19037,N_18514,N_18436);
nor U19038 (N_19038,N_18435,N_18701);
and U19039 (N_19039,N_18734,N_18402);
xor U19040 (N_19040,N_18654,N_18579);
and U19041 (N_19041,N_18714,N_18706);
or U19042 (N_19042,N_18573,N_18586);
xor U19043 (N_19043,N_18416,N_18517);
and U19044 (N_19044,N_18772,N_18631);
or U19045 (N_19045,N_18561,N_18754);
and U19046 (N_19046,N_18762,N_18436);
and U19047 (N_19047,N_18450,N_18759);
or U19048 (N_19048,N_18424,N_18658);
nand U19049 (N_19049,N_18666,N_18428);
nor U19050 (N_19050,N_18788,N_18784);
and U19051 (N_19051,N_18781,N_18720);
and U19052 (N_19052,N_18772,N_18449);
nand U19053 (N_19053,N_18764,N_18593);
or U19054 (N_19054,N_18624,N_18501);
nor U19055 (N_19055,N_18516,N_18444);
nand U19056 (N_19056,N_18772,N_18784);
xor U19057 (N_19057,N_18480,N_18628);
nand U19058 (N_19058,N_18623,N_18616);
xnor U19059 (N_19059,N_18451,N_18731);
nand U19060 (N_19060,N_18480,N_18525);
nor U19061 (N_19061,N_18648,N_18506);
nand U19062 (N_19062,N_18482,N_18616);
nor U19063 (N_19063,N_18464,N_18566);
xnor U19064 (N_19064,N_18530,N_18598);
nor U19065 (N_19065,N_18531,N_18517);
xor U19066 (N_19066,N_18668,N_18538);
nor U19067 (N_19067,N_18710,N_18550);
or U19068 (N_19068,N_18408,N_18592);
nand U19069 (N_19069,N_18504,N_18792);
xnor U19070 (N_19070,N_18755,N_18514);
and U19071 (N_19071,N_18707,N_18485);
xnor U19072 (N_19072,N_18422,N_18737);
or U19073 (N_19073,N_18489,N_18479);
or U19074 (N_19074,N_18461,N_18697);
xnor U19075 (N_19075,N_18746,N_18531);
xnor U19076 (N_19076,N_18700,N_18411);
or U19077 (N_19077,N_18562,N_18731);
and U19078 (N_19078,N_18407,N_18678);
nor U19079 (N_19079,N_18729,N_18430);
or U19080 (N_19080,N_18704,N_18481);
xnor U19081 (N_19081,N_18530,N_18799);
or U19082 (N_19082,N_18660,N_18513);
xnor U19083 (N_19083,N_18734,N_18723);
and U19084 (N_19084,N_18521,N_18599);
nand U19085 (N_19085,N_18413,N_18668);
nor U19086 (N_19086,N_18711,N_18531);
nand U19087 (N_19087,N_18529,N_18646);
xor U19088 (N_19088,N_18724,N_18662);
and U19089 (N_19089,N_18510,N_18762);
or U19090 (N_19090,N_18669,N_18411);
nor U19091 (N_19091,N_18518,N_18530);
and U19092 (N_19092,N_18631,N_18407);
nor U19093 (N_19093,N_18706,N_18598);
nor U19094 (N_19094,N_18500,N_18463);
and U19095 (N_19095,N_18715,N_18652);
or U19096 (N_19096,N_18662,N_18687);
or U19097 (N_19097,N_18765,N_18432);
or U19098 (N_19098,N_18607,N_18587);
or U19099 (N_19099,N_18511,N_18692);
and U19100 (N_19100,N_18696,N_18685);
nor U19101 (N_19101,N_18508,N_18561);
and U19102 (N_19102,N_18779,N_18658);
xor U19103 (N_19103,N_18694,N_18633);
and U19104 (N_19104,N_18616,N_18563);
and U19105 (N_19105,N_18723,N_18418);
nor U19106 (N_19106,N_18601,N_18784);
nor U19107 (N_19107,N_18665,N_18469);
and U19108 (N_19108,N_18542,N_18770);
and U19109 (N_19109,N_18588,N_18548);
xnor U19110 (N_19110,N_18617,N_18668);
nor U19111 (N_19111,N_18540,N_18744);
nand U19112 (N_19112,N_18598,N_18770);
nor U19113 (N_19113,N_18742,N_18630);
nor U19114 (N_19114,N_18694,N_18443);
and U19115 (N_19115,N_18756,N_18492);
xor U19116 (N_19116,N_18519,N_18724);
nand U19117 (N_19117,N_18403,N_18659);
and U19118 (N_19118,N_18592,N_18587);
or U19119 (N_19119,N_18560,N_18763);
nand U19120 (N_19120,N_18522,N_18523);
or U19121 (N_19121,N_18724,N_18736);
nand U19122 (N_19122,N_18673,N_18423);
and U19123 (N_19123,N_18648,N_18402);
nor U19124 (N_19124,N_18652,N_18663);
xnor U19125 (N_19125,N_18409,N_18734);
nand U19126 (N_19126,N_18572,N_18590);
and U19127 (N_19127,N_18549,N_18621);
or U19128 (N_19128,N_18404,N_18545);
and U19129 (N_19129,N_18787,N_18753);
nor U19130 (N_19130,N_18731,N_18737);
and U19131 (N_19131,N_18664,N_18441);
xnor U19132 (N_19132,N_18617,N_18551);
and U19133 (N_19133,N_18640,N_18518);
nand U19134 (N_19134,N_18455,N_18729);
nor U19135 (N_19135,N_18796,N_18470);
nand U19136 (N_19136,N_18525,N_18669);
nand U19137 (N_19137,N_18442,N_18596);
and U19138 (N_19138,N_18641,N_18723);
xor U19139 (N_19139,N_18651,N_18661);
nor U19140 (N_19140,N_18519,N_18612);
nand U19141 (N_19141,N_18417,N_18601);
nor U19142 (N_19142,N_18407,N_18795);
xnor U19143 (N_19143,N_18429,N_18703);
xnor U19144 (N_19144,N_18453,N_18504);
and U19145 (N_19145,N_18742,N_18651);
nor U19146 (N_19146,N_18452,N_18598);
nand U19147 (N_19147,N_18471,N_18423);
xnor U19148 (N_19148,N_18569,N_18635);
nor U19149 (N_19149,N_18457,N_18511);
xnor U19150 (N_19150,N_18775,N_18551);
or U19151 (N_19151,N_18626,N_18474);
or U19152 (N_19152,N_18481,N_18665);
or U19153 (N_19153,N_18528,N_18594);
and U19154 (N_19154,N_18659,N_18795);
nor U19155 (N_19155,N_18574,N_18748);
or U19156 (N_19156,N_18756,N_18459);
and U19157 (N_19157,N_18465,N_18577);
nand U19158 (N_19158,N_18665,N_18764);
or U19159 (N_19159,N_18709,N_18496);
nor U19160 (N_19160,N_18559,N_18456);
and U19161 (N_19161,N_18550,N_18447);
nand U19162 (N_19162,N_18402,N_18660);
or U19163 (N_19163,N_18428,N_18633);
nand U19164 (N_19164,N_18542,N_18549);
nand U19165 (N_19165,N_18658,N_18575);
nand U19166 (N_19166,N_18604,N_18493);
and U19167 (N_19167,N_18422,N_18616);
or U19168 (N_19168,N_18692,N_18571);
nor U19169 (N_19169,N_18709,N_18639);
and U19170 (N_19170,N_18466,N_18457);
xor U19171 (N_19171,N_18768,N_18474);
xor U19172 (N_19172,N_18415,N_18411);
xor U19173 (N_19173,N_18510,N_18506);
or U19174 (N_19174,N_18575,N_18713);
xor U19175 (N_19175,N_18715,N_18402);
xor U19176 (N_19176,N_18709,N_18731);
or U19177 (N_19177,N_18533,N_18689);
nor U19178 (N_19178,N_18702,N_18799);
and U19179 (N_19179,N_18455,N_18707);
xor U19180 (N_19180,N_18449,N_18410);
nand U19181 (N_19181,N_18517,N_18780);
nand U19182 (N_19182,N_18720,N_18404);
and U19183 (N_19183,N_18542,N_18495);
or U19184 (N_19184,N_18609,N_18462);
or U19185 (N_19185,N_18544,N_18716);
and U19186 (N_19186,N_18513,N_18612);
nand U19187 (N_19187,N_18510,N_18422);
and U19188 (N_19188,N_18563,N_18605);
nand U19189 (N_19189,N_18607,N_18718);
nand U19190 (N_19190,N_18593,N_18520);
xnor U19191 (N_19191,N_18479,N_18465);
or U19192 (N_19192,N_18551,N_18444);
nand U19193 (N_19193,N_18735,N_18424);
xor U19194 (N_19194,N_18722,N_18554);
nor U19195 (N_19195,N_18759,N_18599);
nand U19196 (N_19196,N_18719,N_18564);
xnor U19197 (N_19197,N_18608,N_18509);
xnor U19198 (N_19198,N_18586,N_18417);
xnor U19199 (N_19199,N_18787,N_18411);
and U19200 (N_19200,N_19160,N_18847);
xor U19201 (N_19201,N_18963,N_19130);
nor U19202 (N_19202,N_18973,N_18991);
xnor U19203 (N_19203,N_19137,N_19150);
xnor U19204 (N_19204,N_18879,N_19133);
nor U19205 (N_19205,N_19079,N_19178);
or U19206 (N_19206,N_18861,N_19011);
xnor U19207 (N_19207,N_18851,N_19076);
or U19208 (N_19208,N_19067,N_19113);
nand U19209 (N_19209,N_19016,N_18871);
and U19210 (N_19210,N_18969,N_19152);
or U19211 (N_19211,N_18918,N_18950);
nand U19212 (N_19212,N_19126,N_18986);
or U19213 (N_19213,N_19027,N_18814);
nand U19214 (N_19214,N_19001,N_18877);
xnor U19215 (N_19215,N_19115,N_18942);
and U19216 (N_19216,N_19087,N_18857);
nand U19217 (N_19217,N_18937,N_18941);
nand U19218 (N_19218,N_19002,N_18804);
nor U19219 (N_19219,N_18901,N_18919);
nand U19220 (N_19220,N_19052,N_19191);
or U19221 (N_19221,N_19118,N_18834);
nor U19222 (N_19222,N_18954,N_18939);
nor U19223 (N_19223,N_18890,N_18912);
nand U19224 (N_19224,N_19154,N_18846);
nand U19225 (N_19225,N_19101,N_18813);
and U19226 (N_19226,N_19054,N_18835);
and U19227 (N_19227,N_18805,N_18800);
xnor U19228 (N_19228,N_19182,N_18887);
nor U19229 (N_19229,N_19066,N_19139);
and U19230 (N_19230,N_19042,N_18981);
nor U19231 (N_19231,N_18898,N_19058);
nand U19232 (N_19232,N_19084,N_19043);
nand U19233 (N_19233,N_18976,N_19111);
or U19234 (N_19234,N_18970,N_18966);
and U19235 (N_19235,N_18867,N_18817);
xor U19236 (N_19236,N_18998,N_19104);
nand U19237 (N_19237,N_18825,N_19037);
or U19238 (N_19238,N_19125,N_18803);
and U19239 (N_19239,N_19049,N_18811);
or U19240 (N_19240,N_19140,N_18931);
and U19241 (N_19241,N_18995,N_18917);
or U19242 (N_19242,N_18810,N_18878);
nor U19243 (N_19243,N_18845,N_19156);
and U19244 (N_19244,N_19063,N_19145);
nand U19245 (N_19245,N_19081,N_19075);
xnor U19246 (N_19246,N_19183,N_19185);
xor U19247 (N_19247,N_18959,N_19094);
or U19248 (N_19248,N_19004,N_18983);
nand U19249 (N_19249,N_19162,N_19022);
or U19250 (N_19250,N_19007,N_18920);
nor U19251 (N_19251,N_19034,N_18909);
xnor U19252 (N_19252,N_19061,N_19073);
nand U19253 (N_19253,N_19192,N_19196);
nor U19254 (N_19254,N_18921,N_19151);
nand U19255 (N_19255,N_18911,N_19032);
or U19256 (N_19256,N_19129,N_19167);
nand U19257 (N_19257,N_19189,N_19047);
and U19258 (N_19258,N_18967,N_19065);
nor U19259 (N_19259,N_18815,N_18885);
xor U19260 (N_19260,N_19174,N_18893);
nor U19261 (N_19261,N_19109,N_18996);
nor U19262 (N_19262,N_19127,N_18923);
nor U19263 (N_19263,N_18906,N_19142);
and U19264 (N_19264,N_19048,N_19062);
nand U19265 (N_19265,N_18971,N_18934);
or U19266 (N_19266,N_18974,N_18808);
and U19267 (N_19267,N_19082,N_18872);
xor U19268 (N_19268,N_19057,N_18860);
and U19269 (N_19269,N_19106,N_19138);
and U19270 (N_19270,N_19021,N_18819);
nand U19271 (N_19271,N_19036,N_19060);
xor U19272 (N_19272,N_19128,N_18826);
xor U19273 (N_19273,N_18806,N_19055);
and U19274 (N_19274,N_18838,N_18985);
xor U19275 (N_19275,N_19013,N_18840);
or U19276 (N_19276,N_19157,N_19143);
and U19277 (N_19277,N_18952,N_19199);
xnor U19278 (N_19278,N_18975,N_19198);
and U19279 (N_19279,N_18957,N_18848);
xor U19280 (N_19280,N_18930,N_19144);
nand U19281 (N_19281,N_19184,N_19035);
or U19282 (N_19282,N_18895,N_18888);
nand U19283 (N_19283,N_19026,N_18854);
or U19284 (N_19284,N_18843,N_19018);
and U19285 (N_19285,N_18829,N_18870);
or U19286 (N_19286,N_19008,N_19141);
and U19287 (N_19287,N_19040,N_18948);
nand U19288 (N_19288,N_19175,N_18982);
nor U19289 (N_19289,N_19170,N_18896);
xnor U19290 (N_19290,N_18936,N_18944);
and U19291 (N_19291,N_18913,N_18801);
and U19292 (N_19292,N_19131,N_18947);
nor U19293 (N_19293,N_19046,N_19017);
and U19294 (N_19294,N_19136,N_18842);
and U19295 (N_19295,N_18924,N_19166);
nand U19296 (N_19296,N_18822,N_19187);
nand U19297 (N_19297,N_18999,N_19091);
nand U19298 (N_19298,N_18965,N_19064);
nor U19299 (N_19299,N_19014,N_18886);
nor U19300 (N_19300,N_18849,N_19159);
or U19301 (N_19301,N_18916,N_18943);
nand U19302 (N_19302,N_19181,N_19146);
nand U19303 (N_19303,N_18859,N_18892);
nand U19304 (N_19304,N_18980,N_19120);
and U19305 (N_19305,N_18858,N_18933);
and U19306 (N_19306,N_18964,N_18960);
and U19307 (N_19307,N_18821,N_18988);
nor U19308 (N_19308,N_19155,N_18836);
and U19309 (N_19309,N_19100,N_18908);
nand U19310 (N_19310,N_18946,N_19093);
or U19311 (N_19311,N_18928,N_19193);
and U19312 (N_19312,N_19161,N_18951);
or U19313 (N_19313,N_18956,N_19180);
nor U19314 (N_19314,N_18831,N_19194);
nand U19315 (N_19315,N_18997,N_19164);
nor U19316 (N_19316,N_19041,N_18863);
and U19317 (N_19317,N_19020,N_18961);
or U19318 (N_19318,N_19165,N_18881);
xor U19319 (N_19319,N_19090,N_19050);
xor U19320 (N_19320,N_18868,N_18977);
xnor U19321 (N_19321,N_19124,N_19158);
nor U19322 (N_19322,N_19024,N_19078);
and U19323 (N_19323,N_19039,N_19077);
and U19324 (N_19324,N_19147,N_19045);
nor U19325 (N_19325,N_19172,N_19068);
xor U19326 (N_19326,N_18828,N_19169);
nor U19327 (N_19327,N_19108,N_19117);
or U19328 (N_19328,N_18874,N_18992);
and U19329 (N_19329,N_18802,N_19059);
or U19330 (N_19330,N_19033,N_18899);
xnor U19331 (N_19331,N_19122,N_18869);
and U19332 (N_19332,N_19070,N_18962);
nand U19333 (N_19333,N_18866,N_18894);
nor U19334 (N_19334,N_18816,N_18862);
and U19335 (N_19335,N_18827,N_18987);
xor U19336 (N_19336,N_18875,N_18865);
and U19337 (N_19337,N_19163,N_18873);
nand U19338 (N_19338,N_19103,N_19171);
or U19339 (N_19339,N_18853,N_19051);
or U19340 (N_19340,N_19179,N_19168);
or U19341 (N_19341,N_19088,N_19096);
or U19342 (N_19342,N_18940,N_18905);
xnor U19343 (N_19343,N_18990,N_18891);
nor U19344 (N_19344,N_19099,N_19005);
nor U19345 (N_19345,N_19009,N_18958);
nand U19346 (N_19346,N_19085,N_19083);
nand U19347 (N_19347,N_19044,N_19038);
xnor U19348 (N_19348,N_19071,N_18949);
xor U19349 (N_19349,N_18935,N_19123);
xor U19350 (N_19350,N_18841,N_18830);
and U19351 (N_19351,N_18955,N_18903);
or U19352 (N_19352,N_19019,N_18889);
and U19353 (N_19353,N_19114,N_19148);
nand U19354 (N_19354,N_18883,N_18809);
nor U19355 (N_19355,N_18812,N_19010);
and U19356 (N_19356,N_19197,N_18922);
nor U19357 (N_19357,N_19098,N_19000);
or U19358 (N_19358,N_19153,N_19030);
nand U19359 (N_19359,N_19095,N_18907);
and U19360 (N_19360,N_19072,N_18910);
nor U19361 (N_19361,N_18914,N_19177);
or U19362 (N_19362,N_19105,N_18850);
xor U19363 (N_19363,N_18818,N_18945);
and U19364 (N_19364,N_18837,N_18979);
or U19365 (N_19365,N_18932,N_19186);
nor U19366 (N_19366,N_18833,N_19025);
nor U19367 (N_19367,N_19195,N_18993);
and U19368 (N_19368,N_18925,N_19190);
nor U19369 (N_19369,N_18807,N_18882);
or U19370 (N_19370,N_19015,N_18978);
nand U19371 (N_19371,N_19089,N_19031);
or U19372 (N_19372,N_19080,N_18994);
nand U19373 (N_19373,N_18902,N_19006);
nand U19374 (N_19374,N_18852,N_19074);
or U19375 (N_19375,N_18832,N_19173);
or U19376 (N_19376,N_18927,N_19012);
nand U19377 (N_19377,N_19112,N_18972);
xnor U19378 (N_19378,N_19029,N_19135);
nor U19379 (N_19379,N_19028,N_18844);
xor U19380 (N_19380,N_19069,N_18929);
nand U19381 (N_19381,N_18824,N_18855);
or U19382 (N_19382,N_19107,N_18876);
nor U19383 (N_19383,N_18864,N_19102);
nor U19384 (N_19384,N_18823,N_18820);
or U19385 (N_19385,N_19110,N_18900);
xnor U19386 (N_19386,N_19176,N_19053);
nand U19387 (N_19387,N_18953,N_19188);
or U19388 (N_19388,N_19097,N_19119);
nor U19389 (N_19389,N_18904,N_19056);
and U19390 (N_19390,N_19132,N_19116);
nor U19391 (N_19391,N_18938,N_19134);
xnor U19392 (N_19392,N_19121,N_18984);
and U19393 (N_19393,N_19086,N_19003);
nand U19394 (N_19394,N_18915,N_18839);
nor U19395 (N_19395,N_18968,N_18897);
xor U19396 (N_19396,N_18926,N_18884);
xor U19397 (N_19397,N_19149,N_18880);
xor U19398 (N_19398,N_18856,N_19092);
nor U19399 (N_19399,N_19023,N_18989);
and U19400 (N_19400,N_19072,N_18972);
and U19401 (N_19401,N_19157,N_19095);
and U19402 (N_19402,N_19059,N_18902);
nand U19403 (N_19403,N_19064,N_19126);
nand U19404 (N_19404,N_19133,N_19008);
nand U19405 (N_19405,N_19001,N_19105);
xnor U19406 (N_19406,N_18826,N_19060);
xnor U19407 (N_19407,N_18920,N_19030);
xor U19408 (N_19408,N_18959,N_18836);
and U19409 (N_19409,N_19045,N_19116);
xnor U19410 (N_19410,N_18999,N_19168);
and U19411 (N_19411,N_18820,N_19119);
nor U19412 (N_19412,N_18956,N_18966);
or U19413 (N_19413,N_18892,N_19071);
and U19414 (N_19414,N_18935,N_19143);
or U19415 (N_19415,N_18982,N_18951);
or U19416 (N_19416,N_19117,N_19072);
and U19417 (N_19417,N_19136,N_19031);
nand U19418 (N_19418,N_19100,N_19027);
xnor U19419 (N_19419,N_19120,N_18916);
nor U19420 (N_19420,N_18810,N_19044);
nand U19421 (N_19421,N_18884,N_18981);
and U19422 (N_19422,N_18826,N_18955);
xor U19423 (N_19423,N_19106,N_18970);
or U19424 (N_19424,N_18987,N_19075);
nor U19425 (N_19425,N_19141,N_19028);
xor U19426 (N_19426,N_19078,N_18938);
and U19427 (N_19427,N_19023,N_19057);
and U19428 (N_19428,N_18801,N_18920);
nand U19429 (N_19429,N_19032,N_18840);
or U19430 (N_19430,N_19129,N_19043);
nor U19431 (N_19431,N_18952,N_19150);
nand U19432 (N_19432,N_19023,N_18926);
and U19433 (N_19433,N_18884,N_18831);
or U19434 (N_19434,N_19094,N_19195);
nand U19435 (N_19435,N_18928,N_19142);
nand U19436 (N_19436,N_19046,N_19076);
or U19437 (N_19437,N_19083,N_18861);
or U19438 (N_19438,N_19095,N_19169);
nand U19439 (N_19439,N_19194,N_18852);
xnor U19440 (N_19440,N_19182,N_18954);
or U19441 (N_19441,N_19156,N_18880);
xnor U19442 (N_19442,N_19035,N_18923);
or U19443 (N_19443,N_18813,N_19092);
or U19444 (N_19444,N_19067,N_19187);
and U19445 (N_19445,N_18928,N_19075);
or U19446 (N_19446,N_18878,N_19053);
and U19447 (N_19447,N_18995,N_18989);
nor U19448 (N_19448,N_18897,N_19050);
nor U19449 (N_19449,N_19077,N_19078);
xor U19450 (N_19450,N_19188,N_18886);
xor U19451 (N_19451,N_19182,N_18827);
nor U19452 (N_19452,N_18869,N_19176);
or U19453 (N_19453,N_18811,N_18958);
nor U19454 (N_19454,N_18821,N_18945);
and U19455 (N_19455,N_19178,N_19023);
nor U19456 (N_19456,N_18858,N_18867);
nand U19457 (N_19457,N_18954,N_19026);
and U19458 (N_19458,N_18976,N_18808);
nor U19459 (N_19459,N_18805,N_18907);
nor U19460 (N_19460,N_18943,N_18847);
xor U19461 (N_19461,N_19155,N_18840);
or U19462 (N_19462,N_19118,N_18938);
or U19463 (N_19463,N_19196,N_18991);
or U19464 (N_19464,N_18991,N_18819);
nor U19465 (N_19465,N_18910,N_19086);
and U19466 (N_19466,N_18955,N_18983);
xnor U19467 (N_19467,N_18868,N_18965);
nand U19468 (N_19468,N_18835,N_18855);
or U19469 (N_19469,N_18873,N_19195);
or U19470 (N_19470,N_19039,N_18917);
or U19471 (N_19471,N_18846,N_18966);
xor U19472 (N_19472,N_18939,N_19153);
nand U19473 (N_19473,N_18808,N_18937);
and U19474 (N_19474,N_19198,N_18845);
and U19475 (N_19475,N_18839,N_19046);
nand U19476 (N_19476,N_19177,N_19048);
nand U19477 (N_19477,N_19174,N_18887);
or U19478 (N_19478,N_18882,N_18946);
nor U19479 (N_19479,N_18982,N_18916);
and U19480 (N_19480,N_19188,N_18972);
or U19481 (N_19481,N_19129,N_19162);
nand U19482 (N_19482,N_18975,N_19147);
xnor U19483 (N_19483,N_18881,N_18862);
nor U19484 (N_19484,N_18960,N_19072);
nand U19485 (N_19485,N_19102,N_19122);
nor U19486 (N_19486,N_18871,N_18925);
nor U19487 (N_19487,N_19000,N_19106);
nor U19488 (N_19488,N_19010,N_19129);
nand U19489 (N_19489,N_19039,N_18876);
or U19490 (N_19490,N_18850,N_19192);
or U19491 (N_19491,N_18864,N_18810);
xor U19492 (N_19492,N_18970,N_18864);
or U19493 (N_19493,N_19016,N_18942);
nand U19494 (N_19494,N_18961,N_18935);
xnor U19495 (N_19495,N_19147,N_19077);
nand U19496 (N_19496,N_18870,N_18998);
xnor U19497 (N_19497,N_18880,N_18894);
nor U19498 (N_19498,N_19060,N_18925);
or U19499 (N_19499,N_18899,N_18877);
nor U19500 (N_19500,N_19032,N_19059);
or U19501 (N_19501,N_19164,N_18839);
or U19502 (N_19502,N_19123,N_19142);
nor U19503 (N_19503,N_18898,N_19163);
and U19504 (N_19504,N_19067,N_18909);
nor U19505 (N_19505,N_18881,N_19101);
nor U19506 (N_19506,N_19081,N_19127);
xor U19507 (N_19507,N_18843,N_19037);
xor U19508 (N_19508,N_18843,N_18983);
or U19509 (N_19509,N_18938,N_18950);
nand U19510 (N_19510,N_18828,N_19117);
or U19511 (N_19511,N_18996,N_18945);
nor U19512 (N_19512,N_19103,N_18915);
nor U19513 (N_19513,N_19103,N_18864);
or U19514 (N_19514,N_18809,N_19143);
or U19515 (N_19515,N_18980,N_19176);
nor U19516 (N_19516,N_18972,N_19049);
or U19517 (N_19517,N_19151,N_18862);
xnor U19518 (N_19518,N_19173,N_18867);
nor U19519 (N_19519,N_19123,N_19016);
nor U19520 (N_19520,N_18920,N_18885);
nand U19521 (N_19521,N_18810,N_19163);
nand U19522 (N_19522,N_19086,N_18834);
or U19523 (N_19523,N_18839,N_19089);
nand U19524 (N_19524,N_19163,N_19050);
and U19525 (N_19525,N_19000,N_19092);
nand U19526 (N_19526,N_18951,N_19013);
nor U19527 (N_19527,N_19075,N_19199);
xor U19528 (N_19528,N_18901,N_19061);
xnor U19529 (N_19529,N_19134,N_19075);
and U19530 (N_19530,N_18851,N_19097);
xor U19531 (N_19531,N_19150,N_19162);
nor U19532 (N_19532,N_19070,N_18968);
xnor U19533 (N_19533,N_19093,N_18996);
or U19534 (N_19534,N_19173,N_18830);
or U19535 (N_19535,N_18954,N_19034);
and U19536 (N_19536,N_18824,N_19041);
nand U19537 (N_19537,N_19006,N_19149);
nand U19538 (N_19538,N_19010,N_18948);
nor U19539 (N_19539,N_19100,N_19061);
or U19540 (N_19540,N_18954,N_18816);
or U19541 (N_19541,N_18941,N_18901);
and U19542 (N_19542,N_18869,N_19038);
nor U19543 (N_19543,N_19145,N_18815);
nor U19544 (N_19544,N_19174,N_19165);
nor U19545 (N_19545,N_18918,N_19064);
and U19546 (N_19546,N_19141,N_19187);
and U19547 (N_19547,N_19026,N_18992);
nor U19548 (N_19548,N_19185,N_18952);
and U19549 (N_19549,N_19117,N_18886);
and U19550 (N_19550,N_18868,N_19198);
nand U19551 (N_19551,N_18925,N_18881);
and U19552 (N_19552,N_19061,N_19165);
or U19553 (N_19553,N_19052,N_19087);
or U19554 (N_19554,N_19064,N_19125);
xor U19555 (N_19555,N_18942,N_18882);
or U19556 (N_19556,N_18988,N_19134);
nand U19557 (N_19557,N_19031,N_18883);
or U19558 (N_19558,N_18952,N_19039);
nor U19559 (N_19559,N_19034,N_18894);
or U19560 (N_19560,N_19185,N_19179);
and U19561 (N_19561,N_19014,N_19172);
xnor U19562 (N_19562,N_18954,N_18897);
and U19563 (N_19563,N_19174,N_19105);
xor U19564 (N_19564,N_18853,N_18983);
or U19565 (N_19565,N_19017,N_19126);
nor U19566 (N_19566,N_18923,N_18932);
nand U19567 (N_19567,N_19103,N_18990);
nor U19568 (N_19568,N_19007,N_19120);
and U19569 (N_19569,N_18838,N_18902);
nor U19570 (N_19570,N_19171,N_18951);
nand U19571 (N_19571,N_19041,N_18988);
xor U19572 (N_19572,N_19190,N_19100);
and U19573 (N_19573,N_18859,N_19199);
or U19574 (N_19574,N_19000,N_19091);
or U19575 (N_19575,N_18837,N_18828);
xnor U19576 (N_19576,N_18857,N_18883);
and U19577 (N_19577,N_19140,N_18875);
or U19578 (N_19578,N_19030,N_18942);
nor U19579 (N_19579,N_19116,N_19181);
and U19580 (N_19580,N_18912,N_19030);
nand U19581 (N_19581,N_18899,N_18873);
nand U19582 (N_19582,N_18849,N_19125);
nor U19583 (N_19583,N_19178,N_19153);
or U19584 (N_19584,N_19065,N_19018);
nor U19585 (N_19585,N_18809,N_18926);
xor U19586 (N_19586,N_19063,N_18804);
or U19587 (N_19587,N_19149,N_18935);
xnor U19588 (N_19588,N_19173,N_18974);
nand U19589 (N_19589,N_18843,N_18973);
and U19590 (N_19590,N_18812,N_18820);
nor U19591 (N_19591,N_18870,N_18980);
and U19592 (N_19592,N_19119,N_18938);
nand U19593 (N_19593,N_19192,N_19117);
or U19594 (N_19594,N_18939,N_19084);
or U19595 (N_19595,N_19193,N_19084);
xnor U19596 (N_19596,N_18880,N_19127);
and U19597 (N_19597,N_19071,N_19016);
or U19598 (N_19598,N_18895,N_19140);
and U19599 (N_19599,N_19047,N_18996);
and U19600 (N_19600,N_19549,N_19498);
nand U19601 (N_19601,N_19358,N_19292);
nand U19602 (N_19602,N_19279,N_19266);
or U19603 (N_19603,N_19380,N_19249);
and U19604 (N_19604,N_19426,N_19512);
or U19605 (N_19605,N_19458,N_19444);
nand U19606 (N_19606,N_19390,N_19242);
nor U19607 (N_19607,N_19431,N_19471);
xnor U19608 (N_19608,N_19570,N_19245);
nor U19609 (N_19609,N_19463,N_19499);
and U19610 (N_19610,N_19328,N_19262);
or U19611 (N_19611,N_19568,N_19542);
nor U19612 (N_19612,N_19467,N_19539);
xor U19613 (N_19613,N_19434,N_19235);
xnor U19614 (N_19614,N_19450,N_19581);
or U19615 (N_19615,N_19415,N_19312);
nand U19616 (N_19616,N_19562,N_19445);
nor U19617 (N_19617,N_19550,N_19521);
or U19618 (N_19618,N_19525,N_19258);
and U19619 (N_19619,N_19409,N_19482);
nor U19620 (N_19620,N_19511,N_19345);
and U19621 (N_19621,N_19487,N_19578);
nand U19622 (N_19622,N_19425,N_19538);
or U19623 (N_19623,N_19288,N_19408);
nand U19624 (N_19624,N_19595,N_19532);
or U19625 (N_19625,N_19220,N_19502);
nand U19626 (N_19626,N_19490,N_19218);
nand U19627 (N_19627,N_19324,N_19453);
or U19628 (N_19628,N_19353,N_19384);
xnor U19629 (N_19629,N_19485,N_19295);
or U19630 (N_19630,N_19333,N_19572);
or U19631 (N_19631,N_19335,N_19286);
nor U19632 (N_19632,N_19522,N_19251);
xnor U19633 (N_19633,N_19418,N_19206);
and U19634 (N_19634,N_19347,N_19494);
nand U19635 (N_19635,N_19492,N_19533);
and U19636 (N_19636,N_19559,N_19460);
nand U19637 (N_19637,N_19212,N_19497);
or U19638 (N_19638,N_19513,N_19537);
xnor U19639 (N_19639,N_19464,N_19405);
and U19640 (N_19640,N_19489,N_19438);
or U19641 (N_19641,N_19457,N_19342);
and U19642 (N_19642,N_19493,N_19354);
or U19643 (N_19643,N_19466,N_19571);
or U19644 (N_19644,N_19423,N_19404);
nand U19645 (N_19645,N_19203,N_19569);
and U19646 (N_19646,N_19211,N_19310);
xnor U19647 (N_19647,N_19486,N_19383);
nor U19648 (N_19648,N_19302,N_19516);
or U19649 (N_19649,N_19228,N_19585);
nor U19650 (N_19650,N_19406,N_19505);
nor U19651 (N_19651,N_19282,N_19455);
and U19652 (N_19652,N_19399,N_19340);
and U19653 (N_19653,N_19337,N_19545);
or U19654 (N_19654,N_19241,N_19352);
xor U19655 (N_19655,N_19305,N_19285);
nand U19656 (N_19656,N_19276,N_19366);
nand U19657 (N_19657,N_19370,N_19309);
xnor U19658 (N_19658,N_19403,N_19429);
xnor U19659 (N_19659,N_19555,N_19209);
nand U19660 (N_19660,N_19402,N_19346);
and U19661 (N_19661,N_19243,N_19386);
xnor U19662 (N_19662,N_19433,N_19330);
nor U19663 (N_19663,N_19393,N_19259);
xor U19664 (N_19664,N_19520,N_19591);
and U19665 (N_19665,N_19563,N_19316);
xor U19666 (N_19666,N_19319,N_19435);
xor U19667 (N_19667,N_19514,N_19510);
or U19668 (N_19668,N_19400,N_19517);
nor U19669 (N_19669,N_19411,N_19265);
nor U19670 (N_19670,N_19558,N_19491);
or U19671 (N_19671,N_19326,N_19267);
and U19672 (N_19672,N_19541,N_19543);
nor U19673 (N_19673,N_19320,N_19246);
or U19674 (N_19674,N_19227,N_19307);
nor U19675 (N_19675,N_19391,N_19238);
xor U19676 (N_19676,N_19219,N_19588);
and U19677 (N_19677,N_19526,N_19233);
and U19678 (N_19678,N_19379,N_19407);
or U19679 (N_19679,N_19436,N_19261);
nor U19680 (N_19680,N_19461,N_19336);
and U19681 (N_19681,N_19350,N_19597);
or U19682 (N_19682,N_19318,N_19214);
nand U19683 (N_19683,N_19313,N_19546);
nand U19684 (N_19684,N_19274,N_19303);
and U19685 (N_19685,N_19557,N_19361);
xnor U19686 (N_19686,N_19574,N_19480);
or U19687 (N_19687,N_19293,N_19278);
nand U19688 (N_19688,N_19323,N_19584);
or U19689 (N_19689,N_19504,N_19417);
nand U19690 (N_19690,N_19495,N_19226);
nor U19691 (N_19691,N_19341,N_19388);
xor U19692 (N_19692,N_19580,N_19509);
and U19693 (N_19693,N_19441,N_19397);
nor U19694 (N_19694,N_19264,N_19410);
nor U19695 (N_19695,N_19240,N_19527);
and U19696 (N_19696,N_19465,N_19476);
or U19697 (N_19697,N_19396,N_19456);
and U19698 (N_19698,N_19506,N_19232);
and U19699 (N_19699,N_19225,N_19430);
and U19700 (N_19700,N_19277,N_19373);
and U19701 (N_19701,N_19413,N_19420);
nand U19702 (N_19702,N_19356,N_19582);
nor U19703 (N_19703,N_19377,N_19385);
or U19704 (N_19704,N_19298,N_19587);
xnor U19705 (N_19705,N_19416,N_19473);
and U19706 (N_19706,N_19357,N_19564);
xor U19707 (N_19707,N_19579,N_19381);
xnor U19708 (N_19708,N_19204,N_19221);
nor U19709 (N_19709,N_19394,N_19412);
or U19710 (N_19710,N_19334,N_19213);
and U19711 (N_19711,N_19311,N_19208);
or U19712 (N_19712,N_19589,N_19401);
and U19713 (N_19713,N_19553,N_19556);
or U19714 (N_19714,N_19577,N_19291);
nor U19715 (N_19715,N_19483,N_19325);
nand U19716 (N_19716,N_19314,N_19343);
and U19717 (N_19717,N_19253,N_19427);
or U19718 (N_19718,N_19359,N_19474);
nor U19719 (N_19719,N_19317,N_19573);
xor U19720 (N_19720,N_19338,N_19528);
or U19721 (N_19721,N_19363,N_19301);
or U19722 (N_19722,N_19560,N_19369);
nor U19723 (N_19723,N_19440,N_19280);
and U19724 (N_19724,N_19216,N_19501);
nand U19725 (N_19725,N_19566,N_19344);
nor U19726 (N_19726,N_19478,N_19231);
nor U19727 (N_19727,N_19367,N_19257);
or U19728 (N_19728,N_19376,N_19548);
xnor U19729 (N_19729,N_19364,N_19229);
or U19730 (N_19730,N_19244,N_19547);
and U19731 (N_19731,N_19500,N_19375);
and U19732 (N_19732,N_19387,N_19565);
and U19733 (N_19733,N_19224,N_19419);
xor U19734 (N_19734,N_19331,N_19348);
nor U19735 (N_19735,N_19552,N_19382);
or U19736 (N_19736,N_19508,N_19596);
nor U19737 (N_19737,N_19439,N_19551);
xor U19738 (N_19738,N_19462,N_19308);
and U19739 (N_19739,N_19446,N_19593);
nand U19740 (N_19740,N_19294,N_19247);
nor U19741 (N_19741,N_19398,N_19332);
or U19742 (N_19742,N_19534,N_19531);
nand U19743 (N_19743,N_19371,N_19583);
xor U19744 (N_19744,N_19300,N_19268);
xor U19745 (N_19745,N_19270,N_19496);
nor U19746 (N_19746,N_19222,N_19575);
and U19747 (N_19747,N_19205,N_19428);
nor U19748 (N_19748,N_19215,N_19524);
xor U19749 (N_19749,N_19479,N_19250);
and U19750 (N_19750,N_19468,N_19374);
nand U19751 (N_19751,N_19477,N_19260);
nand U19752 (N_19752,N_19217,N_19443);
and U19753 (N_19753,N_19594,N_19201);
xnor U19754 (N_19754,N_19207,N_19372);
nand U19755 (N_19755,N_19421,N_19432);
nand U19756 (N_19756,N_19561,N_19523);
nand U19757 (N_19757,N_19289,N_19378);
nor U19758 (N_19758,N_19287,N_19459);
and U19759 (N_19759,N_19297,N_19540);
and U19760 (N_19760,N_19454,N_19424);
nand U19761 (N_19761,N_19223,N_19484);
xor U19762 (N_19762,N_19451,N_19488);
or U19763 (N_19763,N_19481,N_19392);
nor U19764 (N_19764,N_19447,N_19470);
nor U19765 (N_19765,N_19237,N_19475);
or U19766 (N_19766,N_19503,N_19234);
and U19767 (N_19767,N_19269,N_19230);
xnor U19768 (N_19768,N_19329,N_19256);
or U19769 (N_19769,N_19327,N_19281);
and U19770 (N_19770,N_19284,N_19200);
nor U19771 (N_19771,N_19339,N_19322);
nor U19772 (N_19772,N_19263,N_19236);
or U19773 (N_19773,N_19254,N_19507);
nor U19774 (N_19774,N_19519,N_19598);
xnor U19775 (N_19775,N_19529,N_19275);
nor U19776 (N_19776,N_19365,N_19290);
nand U19777 (N_19777,N_19255,N_19202);
nor U19778 (N_19778,N_19349,N_19414);
and U19779 (N_19779,N_19306,N_19252);
nand U19780 (N_19780,N_19535,N_19395);
nand U19781 (N_19781,N_19360,N_19355);
nand U19782 (N_19782,N_19437,N_19248);
nand U19783 (N_19783,N_19304,N_19592);
and U19784 (N_19784,N_19299,N_19362);
xnor U19785 (N_19785,N_19389,N_19530);
or U19786 (N_19786,N_19554,N_19351);
nand U19787 (N_19787,N_19272,N_19368);
xnor U19788 (N_19788,N_19210,N_19271);
and U19789 (N_19789,N_19283,N_19576);
nor U19790 (N_19790,N_19518,N_19544);
xnor U19791 (N_19791,N_19449,N_19586);
or U19792 (N_19792,N_19469,N_19442);
and U19793 (N_19793,N_19296,N_19536);
nor U19794 (N_19794,N_19472,N_19321);
xor U19795 (N_19795,N_19315,N_19515);
or U19796 (N_19796,N_19448,N_19422);
nand U19797 (N_19797,N_19452,N_19567);
and U19798 (N_19798,N_19239,N_19599);
or U19799 (N_19799,N_19273,N_19590);
or U19800 (N_19800,N_19446,N_19213);
xnor U19801 (N_19801,N_19409,N_19353);
xnor U19802 (N_19802,N_19575,N_19569);
and U19803 (N_19803,N_19223,N_19381);
xnor U19804 (N_19804,N_19599,N_19361);
nand U19805 (N_19805,N_19289,N_19537);
nand U19806 (N_19806,N_19520,N_19572);
and U19807 (N_19807,N_19288,N_19359);
xnor U19808 (N_19808,N_19384,N_19465);
nand U19809 (N_19809,N_19480,N_19362);
and U19810 (N_19810,N_19440,N_19498);
nand U19811 (N_19811,N_19492,N_19439);
and U19812 (N_19812,N_19211,N_19439);
and U19813 (N_19813,N_19206,N_19201);
nor U19814 (N_19814,N_19540,N_19396);
xor U19815 (N_19815,N_19461,N_19314);
xnor U19816 (N_19816,N_19285,N_19366);
xnor U19817 (N_19817,N_19519,N_19389);
xnor U19818 (N_19818,N_19457,N_19405);
and U19819 (N_19819,N_19583,N_19448);
or U19820 (N_19820,N_19297,N_19332);
nand U19821 (N_19821,N_19251,N_19238);
nor U19822 (N_19822,N_19240,N_19391);
and U19823 (N_19823,N_19205,N_19389);
and U19824 (N_19824,N_19572,N_19551);
xor U19825 (N_19825,N_19553,N_19255);
nor U19826 (N_19826,N_19459,N_19360);
nand U19827 (N_19827,N_19508,N_19372);
and U19828 (N_19828,N_19408,N_19268);
or U19829 (N_19829,N_19388,N_19383);
nor U19830 (N_19830,N_19323,N_19526);
or U19831 (N_19831,N_19593,N_19548);
nand U19832 (N_19832,N_19533,N_19299);
and U19833 (N_19833,N_19499,N_19577);
xor U19834 (N_19834,N_19575,N_19567);
xor U19835 (N_19835,N_19267,N_19336);
nand U19836 (N_19836,N_19575,N_19409);
and U19837 (N_19837,N_19567,N_19313);
nor U19838 (N_19838,N_19416,N_19296);
nand U19839 (N_19839,N_19349,N_19422);
nand U19840 (N_19840,N_19260,N_19306);
nand U19841 (N_19841,N_19582,N_19391);
nand U19842 (N_19842,N_19401,N_19391);
nor U19843 (N_19843,N_19559,N_19429);
xor U19844 (N_19844,N_19522,N_19201);
nor U19845 (N_19845,N_19461,N_19258);
and U19846 (N_19846,N_19214,N_19570);
nand U19847 (N_19847,N_19591,N_19510);
nand U19848 (N_19848,N_19537,N_19558);
xor U19849 (N_19849,N_19281,N_19471);
nand U19850 (N_19850,N_19427,N_19419);
nor U19851 (N_19851,N_19562,N_19351);
nor U19852 (N_19852,N_19560,N_19530);
nand U19853 (N_19853,N_19462,N_19598);
and U19854 (N_19854,N_19523,N_19396);
nor U19855 (N_19855,N_19260,N_19421);
nand U19856 (N_19856,N_19241,N_19492);
nand U19857 (N_19857,N_19205,N_19378);
xnor U19858 (N_19858,N_19319,N_19317);
or U19859 (N_19859,N_19414,N_19578);
xnor U19860 (N_19860,N_19232,N_19329);
nand U19861 (N_19861,N_19452,N_19559);
nor U19862 (N_19862,N_19256,N_19471);
nand U19863 (N_19863,N_19216,N_19556);
or U19864 (N_19864,N_19343,N_19463);
or U19865 (N_19865,N_19537,N_19457);
or U19866 (N_19866,N_19479,N_19341);
nor U19867 (N_19867,N_19479,N_19598);
and U19868 (N_19868,N_19325,N_19535);
nand U19869 (N_19869,N_19439,N_19355);
and U19870 (N_19870,N_19552,N_19462);
nor U19871 (N_19871,N_19434,N_19414);
nor U19872 (N_19872,N_19290,N_19460);
and U19873 (N_19873,N_19435,N_19406);
and U19874 (N_19874,N_19500,N_19376);
and U19875 (N_19875,N_19430,N_19293);
and U19876 (N_19876,N_19478,N_19378);
and U19877 (N_19877,N_19295,N_19257);
or U19878 (N_19878,N_19297,N_19560);
and U19879 (N_19879,N_19243,N_19233);
or U19880 (N_19880,N_19352,N_19416);
nor U19881 (N_19881,N_19529,N_19350);
nor U19882 (N_19882,N_19463,N_19472);
and U19883 (N_19883,N_19333,N_19534);
or U19884 (N_19884,N_19273,N_19310);
or U19885 (N_19885,N_19247,N_19297);
and U19886 (N_19886,N_19263,N_19448);
or U19887 (N_19887,N_19267,N_19261);
nand U19888 (N_19888,N_19414,N_19229);
xnor U19889 (N_19889,N_19358,N_19278);
nor U19890 (N_19890,N_19487,N_19549);
and U19891 (N_19891,N_19384,N_19211);
nand U19892 (N_19892,N_19416,N_19210);
nand U19893 (N_19893,N_19279,N_19504);
xnor U19894 (N_19894,N_19443,N_19339);
nor U19895 (N_19895,N_19556,N_19482);
nand U19896 (N_19896,N_19401,N_19425);
nor U19897 (N_19897,N_19538,N_19525);
xnor U19898 (N_19898,N_19456,N_19595);
nand U19899 (N_19899,N_19311,N_19515);
nand U19900 (N_19900,N_19251,N_19398);
or U19901 (N_19901,N_19547,N_19276);
and U19902 (N_19902,N_19276,N_19543);
or U19903 (N_19903,N_19224,N_19333);
nand U19904 (N_19904,N_19323,N_19567);
nor U19905 (N_19905,N_19287,N_19490);
xor U19906 (N_19906,N_19215,N_19309);
nand U19907 (N_19907,N_19514,N_19555);
or U19908 (N_19908,N_19488,N_19454);
nor U19909 (N_19909,N_19208,N_19444);
xnor U19910 (N_19910,N_19551,N_19595);
nand U19911 (N_19911,N_19288,N_19263);
nand U19912 (N_19912,N_19452,N_19412);
nor U19913 (N_19913,N_19293,N_19279);
nand U19914 (N_19914,N_19519,N_19236);
and U19915 (N_19915,N_19240,N_19388);
or U19916 (N_19916,N_19413,N_19353);
xor U19917 (N_19917,N_19304,N_19558);
and U19918 (N_19918,N_19284,N_19352);
nand U19919 (N_19919,N_19260,N_19203);
or U19920 (N_19920,N_19213,N_19211);
nor U19921 (N_19921,N_19511,N_19528);
nor U19922 (N_19922,N_19457,N_19580);
xor U19923 (N_19923,N_19270,N_19454);
and U19924 (N_19924,N_19470,N_19230);
nor U19925 (N_19925,N_19578,N_19207);
xnor U19926 (N_19926,N_19390,N_19402);
xnor U19927 (N_19927,N_19549,N_19524);
nor U19928 (N_19928,N_19510,N_19548);
nand U19929 (N_19929,N_19362,N_19330);
and U19930 (N_19930,N_19261,N_19379);
nor U19931 (N_19931,N_19434,N_19550);
nor U19932 (N_19932,N_19226,N_19331);
nor U19933 (N_19933,N_19344,N_19208);
or U19934 (N_19934,N_19320,N_19509);
nand U19935 (N_19935,N_19227,N_19410);
or U19936 (N_19936,N_19400,N_19523);
nor U19937 (N_19937,N_19421,N_19337);
or U19938 (N_19938,N_19270,N_19425);
nand U19939 (N_19939,N_19333,N_19329);
xnor U19940 (N_19940,N_19291,N_19313);
or U19941 (N_19941,N_19569,N_19391);
or U19942 (N_19942,N_19572,N_19343);
nand U19943 (N_19943,N_19429,N_19523);
nand U19944 (N_19944,N_19549,N_19303);
nand U19945 (N_19945,N_19379,N_19334);
xor U19946 (N_19946,N_19275,N_19212);
nand U19947 (N_19947,N_19477,N_19221);
or U19948 (N_19948,N_19305,N_19240);
and U19949 (N_19949,N_19539,N_19431);
nor U19950 (N_19950,N_19474,N_19568);
nor U19951 (N_19951,N_19431,N_19385);
nand U19952 (N_19952,N_19393,N_19366);
nand U19953 (N_19953,N_19516,N_19305);
or U19954 (N_19954,N_19439,N_19330);
and U19955 (N_19955,N_19336,N_19441);
nand U19956 (N_19956,N_19549,N_19461);
xnor U19957 (N_19957,N_19422,N_19533);
xnor U19958 (N_19958,N_19579,N_19439);
and U19959 (N_19959,N_19430,N_19229);
or U19960 (N_19960,N_19292,N_19277);
xor U19961 (N_19961,N_19416,N_19440);
xnor U19962 (N_19962,N_19385,N_19263);
or U19963 (N_19963,N_19450,N_19346);
and U19964 (N_19964,N_19452,N_19277);
or U19965 (N_19965,N_19582,N_19550);
nand U19966 (N_19966,N_19372,N_19374);
nand U19967 (N_19967,N_19572,N_19415);
nand U19968 (N_19968,N_19254,N_19461);
and U19969 (N_19969,N_19377,N_19527);
or U19970 (N_19970,N_19582,N_19491);
or U19971 (N_19971,N_19518,N_19528);
or U19972 (N_19972,N_19354,N_19443);
nand U19973 (N_19973,N_19344,N_19246);
or U19974 (N_19974,N_19408,N_19330);
nand U19975 (N_19975,N_19263,N_19443);
nand U19976 (N_19976,N_19422,N_19275);
and U19977 (N_19977,N_19301,N_19267);
and U19978 (N_19978,N_19385,N_19332);
and U19979 (N_19979,N_19460,N_19425);
nor U19980 (N_19980,N_19383,N_19442);
nand U19981 (N_19981,N_19465,N_19487);
or U19982 (N_19982,N_19300,N_19594);
and U19983 (N_19983,N_19221,N_19389);
and U19984 (N_19984,N_19323,N_19370);
nand U19985 (N_19985,N_19503,N_19468);
or U19986 (N_19986,N_19400,N_19288);
and U19987 (N_19987,N_19461,N_19299);
and U19988 (N_19988,N_19324,N_19375);
and U19989 (N_19989,N_19366,N_19251);
nor U19990 (N_19990,N_19474,N_19579);
and U19991 (N_19991,N_19335,N_19381);
nor U19992 (N_19992,N_19389,N_19447);
nor U19993 (N_19993,N_19206,N_19252);
nand U19994 (N_19994,N_19486,N_19453);
and U19995 (N_19995,N_19537,N_19464);
nor U19996 (N_19996,N_19290,N_19390);
or U19997 (N_19997,N_19322,N_19529);
xnor U19998 (N_19998,N_19373,N_19420);
or U19999 (N_19999,N_19241,N_19366);
xnor UO_0 (O_0,N_19966,N_19840);
and UO_1 (O_1,N_19617,N_19727);
or UO_2 (O_2,N_19983,N_19600);
and UO_3 (O_3,N_19950,N_19639);
and UO_4 (O_4,N_19919,N_19706);
xor UO_5 (O_5,N_19795,N_19914);
and UO_6 (O_6,N_19916,N_19888);
nor UO_7 (O_7,N_19680,N_19673);
or UO_8 (O_8,N_19656,N_19887);
xnor UO_9 (O_9,N_19972,N_19738);
and UO_10 (O_10,N_19743,N_19976);
and UO_11 (O_11,N_19758,N_19883);
or UO_12 (O_12,N_19717,N_19659);
xor UO_13 (O_13,N_19688,N_19954);
and UO_14 (O_14,N_19642,N_19754);
xor UO_15 (O_15,N_19925,N_19830);
xnor UO_16 (O_16,N_19864,N_19943);
and UO_17 (O_17,N_19889,N_19924);
and UO_18 (O_18,N_19683,N_19613);
and UO_19 (O_19,N_19753,N_19751);
or UO_20 (O_20,N_19736,N_19968);
nand UO_21 (O_21,N_19681,N_19603);
nor UO_22 (O_22,N_19990,N_19759);
xnor UO_23 (O_23,N_19971,N_19749);
and UO_24 (O_24,N_19773,N_19674);
nor UO_25 (O_25,N_19652,N_19898);
xnor UO_26 (O_26,N_19609,N_19973);
or UO_27 (O_27,N_19788,N_19905);
nor UO_28 (O_28,N_19756,N_19839);
or UO_29 (O_29,N_19776,N_19655);
xor UO_30 (O_30,N_19610,N_19942);
and UO_31 (O_31,N_19821,N_19808);
and UO_32 (O_32,N_19775,N_19678);
and UO_33 (O_33,N_19915,N_19701);
nand UO_34 (O_34,N_19713,N_19904);
xor UO_35 (O_35,N_19782,N_19725);
nand UO_36 (O_36,N_19661,N_19800);
nand UO_37 (O_37,N_19822,N_19760);
or UO_38 (O_38,N_19764,N_19739);
and UO_39 (O_39,N_19921,N_19791);
xor UO_40 (O_40,N_19938,N_19970);
or UO_41 (O_41,N_19619,N_19869);
and UO_42 (O_42,N_19920,N_19832);
xnor UO_43 (O_43,N_19649,N_19944);
nand UO_44 (O_44,N_19768,N_19997);
nor UO_45 (O_45,N_19996,N_19923);
or UO_46 (O_46,N_19994,N_19828);
nor UO_47 (O_47,N_19690,N_19978);
nand UO_48 (O_48,N_19826,N_19867);
nor UO_49 (O_49,N_19992,N_19695);
and UO_50 (O_50,N_19730,N_19875);
or UO_51 (O_51,N_19824,N_19785);
or UO_52 (O_52,N_19606,N_19786);
and UO_53 (O_53,N_19857,N_19620);
nand UO_54 (O_54,N_19890,N_19918);
xor UO_55 (O_55,N_19902,N_19616);
xnor UO_56 (O_56,N_19658,N_19939);
and UO_57 (O_57,N_19692,N_19926);
or UO_58 (O_58,N_19952,N_19912);
and UO_59 (O_59,N_19720,N_19724);
nor UO_60 (O_60,N_19903,N_19940);
nand UO_61 (O_61,N_19820,N_19657);
nand UO_62 (O_62,N_19772,N_19982);
and UO_63 (O_63,N_19718,N_19856);
nand UO_64 (O_64,N_19851,N_19740);
xor UO_65 (O_65,N_19860,N_19941);
and UO_66 (O_66,N_19910,N_19817);
and UO_67 (O_67,N_19933,N_19750);
or UO_68 (O_68,N_19669,N_19605);
and UO_69 (O_69,N_19638,N_19899);
or UO_70 (O_70,N_19805,N_19797);
nand UO_71 (O_71,N_19614,N_19648);
or UO_72 (O_72,N_19841,N_19909);
xnor UO_73 (O_73,N_19861,N_19960);
nor UO_74 (O_74,N_19927,N_19951);
xor UO_75 (O_75,N_19858,N_19862);
or UO_76 (O_76,N_19794,N_19676);
and UO_77 (O_77,N_19715,N_19825);
nand UO_78 (O_78,N_19789,N_19716);
or UO_79 (O_79,N_19687,N_19908);
xnor UO_80 (O_80,N_19814,N_19991);
or UO_81 (O_81,N_19932,N_19769);
nand UO_82 (O_82,N_19654,N_19777);
or UO_83 (O_83,N_19917,N_19846);
nand UO_84 (O_84,N_19765,N_19700);
nand UO_85 (O_85,N_19728,N_19627);
or UO_86 (O_86,N_19913,N_19670);
or UO_87 (O_87,N_19980,N_19963);
nor UO_88 (O_88,N_19636,N_19757);
nand UO_89 (O_89,N_19866,N_19635);
or UO_90 (O_90,N_19693,N_19849);
nor UO_91 (O_91,N_19865,N_19957);
xnor UO_92 (O_92,N_19696,N_19843);
and UO_93 (O_93,N_19998,N_19784);
and UO_94 (O_94,N_19622,N_19819);
nand UO_95 (O_95,N_19704,N_19884);
or UO_96 (O_96,N_19880,N_19611);
or UO_97 (O_97,N_19995,N_19677);
nand UO_98 (O_98,N_19747,N_19623);
xor UO_99 (O_99,N_19896,N_19831);
nor UO_100 (O_100,N_19956,N_19945);
and UO_101 (O_101,N_19816,N_19807);
and UO_102 (O_102,N_19874,N_19999);
and UO_103 (O_103,N_19781,N_19930);
nand UO_104 (O_104,N_19767,N_19709);
nand UO_105 (O_105,N_19705,N_19762);
and UO_106 (O_106,N_19792,N_19868);
nor UO_107 (O_107,N_19981,N_19891);
nand UO_108 (O_108,N_19612,N_19958);
and UO_109 (O_109,N_19664,N_19936);
and UO_110 (O_110,N_19697,N_19802);
xor UO_111 (O_111,N_19987,N_19876);
xnor UO_112 (O_112,N_19601,N_19702);
nand UO_113 (O_113,N_19947,N_19922);
and UO_114 (O_114,N_19872,N_19878);
xnor UO_115 (O_115,N_19722,N_19885);
xor UO_116 (O_116,N_19827,N_19796);
nor UO_117 (O_117,N_19721,N_19985);
or UO_118 (O_118,N_19892,N_19615);
nand UO_119 (O_119,N_19929,N_19684);
nand UO_120 (O_120,N_19602,N_19848);
xnor UO_121 (O_121,N_19964,N_19886);
and UO_122 (O_122,N_19685,N_19748);
nor UO_123 (O_123,N_19879,N_19967);
or UO_124 (O_124,N_19948,N_19607);
xor UO_125 (O_125,N_19937,N_19618);
nand UO_126 (O_126,N_19818,N_19621);
or UO_127 (O_127,N_19842,N_19726);
and UO_128 (O_128,N_19911,N_19699);
xnor UO_129 (O_129,N_19900,N_19640);
xor UO_130 (O_130,N_19986,N_19643);
nor UO_131 (O_131,N_19719,N_19853);
xnor UO_132 (O_132,N_19928,N_19668);
nand UO_133 (O_133,N_19604,N_19835);
or UO_134 (O_134,N_19955,N_19984);
nand UO_135 (O_135,N_19812,N_19894);
nand UO_136 (O_136,N_19710,N_19780);
or UO_137 (O_137,N_19946,N_19895);
nor UO_138 (O_138,N_19778,N_19810);
or UO_139 (O_139,N_19979,N_19901);
nor UO_140 (O_140,N_19799,N_19637);
nor UO_141 (O_141,N_19608,N_19694);
and UO_142 (O_142,N_19679,N_19633);
nand UO_143 (O_143,N_19752,N_19703);
nand UO_144 (O_144,N_19771,N_19766);
and UO_145 (O_145,N_19714,N_19823);
or UO_146 (O_146,N_19790,N_19949);
nand UO_147 (O_147,N_19634,N_19737);
nand UO_148 (O_148,N_19708,N_19698);
nor UO_149 (O_149,N_19993,N_19733);
and UO_150 (O_150,N_19855,N_19965);
or UO_151 (O_151,N_19630,N_19646);
nand UO_152 (O_152,N_19893,N_19744);
xnor UO_153 (O_153,N_19844,N_19953);
nor UO_154 (O_154,N_19871,N_19763);
xnor UO_155 (O_155,N_19829,N_19734);
or UO_156 (O_156,N_19645,N_19897);
nand UO_157 (O_157,N_19707,N_19755);
and UO_158 (O_158,N_19854,N_19974);
and UO_159 (O_159,N_19870,N_19761);
xnor UO_160 (O_160,N_19837,N_19809);
xnor UO_161 (O_161,N_19806,N_19798);
nand UO_162 (O_162,N_19977,N_19961);
nor UO_163 (O_163,N_19732,N_19804);
xor UO_164 (O_164,N_19813,N_19735);
nand UO_165 (O_165,N_19989,N_19779);
xor UO_166 (O_166,N_19975,N_19850);
nor UO_167 (O_167,N_19731,N_19774);
or UO_168 (O_168,N_19691,N_19833);
or UO_169 (O_169,N_19624,N_19742);
nand UO_170 (O_170,N_19847,N_19834);
or UO_171 (O_171,N_19815,N_19882);
xor UO_172 (O_172,N_19988,N_19859);
nand UO_173 (O_173,N_19845,N_19959);
or UO_174 (O_174,N_19644,N_19663);
and UO_175 (O_175,N_19675,N_19934);
or UO_176 (O_176,N_19723,N_19852);
and UO_177 (O_177,N_19907,N_19682);
or UO_178 (O_178,N_19962,N_19651);
and UO_179 (O_179,N_19628,N_19793);
xor UO_180 (O_180,N_19650,N_19665);
nand UO_181 (O_181,N_19741,N_19801);
nor UO_182 (O_182,N_19671,N_19881);
or UO_183 (O_183,N_19631,N_19787);
xor UO_184 (O_184,N_19729,N_19745);
and UO_185 (O_185,N_19660,N_19647);
nand UO_186 (O_186,N_19626,N_19653);
and UO_187 (O_187,N_19969,N_19931);
or UO_188 (O_188,N_19803,N_19877);
xor UO_189 (O_189,N_19712,N_19783);
or UO_190 (O_190,N_19873,N_19632);
and UO_191 (O_191,N_19746,N_19770);
nand UO_192 (O_192,N_19641,N_19625);
xnor UO_193 (O_193,N_19629,N_19711);
and UO_194 (O_194,N_19666,N_19811);
and UO_195 (O_195,N_19662,N_19906);
nand UO_196 (O_196,N_19863,N_19838);
nand UO_197 (O_197,N_19667,N_19836);
and UO_198 (O_198,N_19672,N_19689);
and UO_199 (O_199,N_19935,N_19686);
and UO_200 (O_200,N_19956,N_19756);
nor UO_201 (O_201,N_19954,N_19710);
and UO_202 (O_202,N_19872,N_19860);
nor UO_203 (O_203,N_19892,N_19851);
nor UO_204 (O_204,N_19992,N_19924);
nand UO_205 (O_205,N_19875,N_19987);
nand UO_206 (O_206,N_19897,N_19611);
and UO_207 (O_207,N_19671,N_19767);
nand UO_208 (O_208,N_19825,N_19815);
and UO_209 (O_209,N_19633,N_19677);
nor UO_210 (O_210,N_19644,N_19697);
and UO_211 (O_211,N_19676,N_19647);
or UO_212 (O_212,N_19966,N_19970);
and UO_213 (O_213,N_19882,N_19627);
nor UO_214 (O_214,N_19918,N_19823);
and UO_215 (O_215,N_19681,N_19853);
or UO_216 (O_216,N_19907,N_19961);
and UO_217 (O_217,N_19816,N_19997);
and UO_218 (O_218,N_19719,N_19870);
xnor UO_219 (O_219,N_19770,N_19787);
and UO_220 (O_220,N_19861,N_19655);
xor UO_221 (O_221,N_19698,N_19693);
or UO_222 (O_222,N_19819,N_19715);
and UO_223 (O_223,N_19638,N_19904);
nor UO_224 (O_224,N_19857,N_19686);
nand UO_225 (O_225,N_19976,N_19616);
nand UO_226 (O_226,N_19606,N_19805);
nand UO_227 (O_227,N_19840,N_19717);
nand UO_228 (O_228,N_19777,N_19951);
and UO_229 (O_229,N_19874,N_19957);
or UO_230 (O_230,N_19969,N_19788);
or UO_231 (O_231,N_19632,N_19779);
nor UO_232 (O_232,N_19851,N_19958);
or UO_233 (O_233,N_19734,N_19789);
nand UO_234 (O_234,N_19824,N_19812);
or UO_235 (O_235,N_19656,N_19783);
nand UO_236 (O_236,N_19893,N_19731);
and UO_237 (O_237,N_19750,N_19711);
nor UO_238 (O_238,N_19759,N_19652);
xor UO_239 (O_239,N_19828,N_19767);
and UO_240 (O_240,N_19938,N_19777);
or UO_241 (O_241,N_19842,N_19724);
nor UO_242 (O_242,N_19618,N_19919);
and UO_243 (O_243,N_19645,N_19957);
nor UO_244 (O_244,N_19851,N_19628);
nor UO_245 (O_245,N_19659,N_19629);
and UO_246 (O_246,N_19981,N_19637);
xor UO_247 (O_247,N_19711,N_19894);
nand UO_248 (O_248,N_19814,N_19820);
and UO_249 (O_249,N_19856,N_19794);
nand UO_250 (O_250,N_19885,N_19730);
and UO_251 (O_251,N_19843,N_19764);
and UO_252 (O_252,N_19669,N_19639);
or UO_253 (O_253,N_19812,N_19809);
or UO_254 (O_254,N_19962,N_19638);
nor UO_255 (O_255,N_19891,N_19733);
xor UO_256 (O_256,N_19807,N_19679);
nand UO_257 (O_257,N_19862,N_19850);
and UO_258 (O_258,N_19986,N_19926);
xnor UO_259 (O_259,N_19866,N_19996);
nor UO_260 (O_260,N_19770,N_19696);
nand UO_261 (O_261,N_19893,N_19718);
xnor UO_262 (O_262,N_19627,N_19644);
nand UO_263 (O_263,N_19863,N_19796);
xor UO_264 (O_264,N_19975,N_19844);
nor UO_265 (O_265,N_19879,N_19686);
and UO_266 (O_266,N_19979,N_19843);
or UO_267 (O_267,N_19914,N_19950);
nand UO_268 (O_268,N_19979,N_19788);
or UO_269 (O_269,N_19632,N_19851);
or UO_270 (O_270,N_19979,N_19705);
nor UO_271 (O_271,N_19748,N_19893);
and UO_272 (O_272,N_19932,N_19720);
nand UO_273 (O_273,N_19895,N_19634);
and UO_274 (O_274,N_19899,N_19963);
nor UO_275 (O_275,N_19630,N_19634);
xor UO_276 (O_276,N_19929,N_19609);
nand UO_277 (O_277,N_19688,N_19715);
nand UO_278 (O_278,N_19848,N_19941);
and UO_279 (O_279,N_19843,N_19678);
and UO_280 (O_280,N_19621,N_19764);
nand UO_281 (O_281,N_19989,N_19637);
and UO_282 (O_282,N_19926,N_19838);
and UO_283 (O_283,N_19779,N_19918);
and UO_284 (O_284,N_19814,N_19615);
and UO_285 (O_285,N_19847,N_19977);
nor UO_286 (O_286,N_19800,N_19654);
nand UO_287 (O_287,N_19953,N_19778);
or UO_288 (O_288,N_19985,N_19739);
nor UO_289 (O_289,N_19993,N_19944);
or UO_290 (O_290,N_19834,N_19792);
or UO_291 (O_291,N_19911,N_19867);
and UO_292 (O_292,N_19818,N_19833);
and UO_293 (O_293,N_19778,N_19606);
nand UO_294 (O_294,N_19648,N_19967);
nand UO_295 (O_295,N_19917,N_19883);
or UO_296 (O_296,N_19788,N_19962);
nor UO_297 (O_297,N_19874,N_19905);
nand UO_298 (O_298,N_19740,N_19653);
xnor UO_299 (O_299,N_19960,N_19985);
nor UO_300 (O_300,N_19906,N_19750);
or UO_301 (O_301,N_19788,N_19674);
nand UO_302 (O_302,N_19664,N_19722);
nand UO_303 (O_303,N_19752,N_19614);
and UO_304 (O_304,N_19789,N_19781);
nand UO_305 (O_305,N_19771,N_19852);
or UO_306 (O_306,N_19923,N_19933);
or UO_307 (O_307,N_19618,N_19911);
nor UO_308 (O_308,N_19698,N_19606);
xnor UO_309 (O_309,N_19956,N_19645);
and UO_310 (O_310,N_19795,N_19891);
or UO_311 (O_311,N_19645,N_19654);
nor UO_312 (O_312,N_19681,N_19665);
xor UO_313 (O_313,N_19746,N_19991);
or UO_314 (O_314,N_19857,N_19993);
or UO_315 (O_315,N_19996,N_19857);
xnor UO_316 (O_316,N_19739,N_19929);
xnor UO_317 (O_317,N_19995,N_19793);
and UO_318 (O_318,N_19600,N_19631);
and UO_319 (O_319,N_19653,N_19900);
nand UO_320 (O_320,N_19814,N_19773);
or UO_321 (O_321,N_19672,N_19606);
and UO_322 (O_322,N_19654,N_19880);
and UO_323 (O_323,N_19694,N_19617);
and UO_324 (O_324,N_19846,N_19750);
nor UO_325 (O_325,N_19769,N_19695);
xor UO_326 (O_326,N_19909,N_19721);
xor UO_327 (O_327,N_19976,N_19862);
or UO_328 (O_328,N_19971,N_19989);
xnor UO_329 (O_329,N_19828,N_19974);
nor UO_330 (O_330,N_19878,N_19602);
nand UO_331 (O_331,N_19747,N_19820);
nor UO_332 (O_332,N_19912,N_19721);
or UO_333 (O_333,N_19711,N_19899);
nor UO_334 (O_334,N_19956,N_19636);
or UO_335 (O_335,N_19932,N_19684);
xnor UO_336 (O_336,N_19991,N_19797);
or UO_337 (O_337,N_19941,N_19874);
xor UO_338 (O_338,N_19993,N_19653);
or UO_339 (O_339,N_19642,N_19963);
and UO_340 (O_340,N_19928,N_19770);
or UO_341 (O_341,N_19969,N_19790);
xor UO_342 (O_342,N_19834,N_19842);
and UO_343 (O_343,N_19948,N_19786);
nor UO_344 (O_344,N_19885,N_19696);
nor UO_345 (O_345,N_19602,N_19774);
or UO_346 (O_346,N_19972,N_19856);
nand UO_347 (O_347,N_19990,N_19781);
and UO_348 (O_348,N_19740,N_19713);
and UO_349 (O_349,N_19810,N_19871);
xor UO_350 (O_350,N_19858,N_19850);
xor UO_351 (O_351,N_19874,N_19923);
or UO_352 (O_352,N_19857,N_19998);
or UO_353 (O_353,N_19952,N_19665);
nor UO_354 (O_354,N_19682,N_19819);
nand UO_355 (O_355,N_19972,N_19622);
and UO_356 (O_356,N_19646,N_19623);
or UO_357 (O_357,N_19727,N_19774);
nand UO_358 (O_358,N_19792,N_19623);
and UO_359 (O_359,N_19605,N_19949);
nand UO_360 (O_360,N_19961,N_19746);
or UO_361 (O_361,N_19999,N_19871);
or UO_362 (O_362,N_19639,N_19954);
nand UO_363 (O_363,N_19998,N_19850);
nand UO_364 (O_364,N_19674,N_19754);
xnor UO_365 (O_365,N_19683,N_19635);
xor UO_366 (O_366,N_19936,N_19883);
nand UO_367 (O_367,N_19749,N_19841);
xnor UO_368 (O_368,N_19972,N_19651);
nand UO_369 (O_369,N_19652,N_19614);
or UO_370 (O_370,N_19687,N_19826);
xnor UO_371 (O_371,N_19748,N_19935);
or UO_372 (O_372,N_19953,N_19703);
xnor UO_373 (O_373,N_19803,N_19917);
or UO_374 (O_374,N_19818,N_19682);
nor UO_375 (O_375,N_19703,N_19851);
or UO_376 (O_376,N_19663,N_19792);
xor UO_377 (O_377,N_19713,N_19774);
or UO_378 (O_378,N_19879,N_19902);
xor UO_379 (O_379,N_19936,N_19738);
and UO_380 (O_380,N_19787,N_19663);
and UO_381 (O_381,N_19747,N_19825);
or UO_382 (O_382,N_19983,N_19680);
xor UO_383 (O_383,N_19764,N_19836);
nand UO_384 (O_384,N_19726,N_19616);
nand UO_385 (O_385,N_19754,N_19870);
or UO_386 (O_386,N_19997,N_19664);
and UO_387 (O_387,N_19603,N_19781);
nor UO_388 (O_388,N_19600,N_19632);
nand UO_389 (O_389,N_19886,N_19790);
nand UO_390 (O_390,N_19891,N_19945);
and UO_391 (O_391,N_19762,N_19722);
or UO_392 (O_392,N_19628,N_19941);
xor UO_393 (O_393,N_19726,N_19640);
or UO_394 (O_394,N_19726,N_19864);
xnor UO_395 (O_395,N_19823,N_19778);
or UO_396 (O_396,N_19703,N_19714);
and UO_397 (O_397,N_19607,N_19879);
nor UO_398 (O_398,N_19734,N_19759);
nand UO_399 (O_399,N_19653,N_19749);
nand UO_400 (O_400,N_19649,N_19647);
nand UO_401 (O_401,N_19775,N_19927);
nor UO_402 (O_402,N_19755,N_19692);
nand UO_403 (O_403,N_19846,N_19627);
and UO_404 (O_404,N_19827,N_19653);
and UO_405 (O_405,N_19735,N_19855);
and UO_406 (O_406,N_19657,N_19751);
and UO_407 (O_407,N_19796,N_19902);
and UO_408 (O_408,N_19921,N_19879);
nand UO_409 (O_409,N_19668,N_19727);
nand UO_410 (O_410,N_19818,N_19907);
nand UO_411 (O_411,N_19800,N_19820);
or UO_412 (O_412,N_19910,N_19833);
and UO_413 (O_413,N_19710,N_19977);
and UO_414 (O_414,N_19716,N_19995);
nand UO_415 (O_415,N_19807,N_19676);
nor UO_416 (O_416,N_19622,N_19713);
xor UO_417 (O_417,N_19761,N_19784);
nand UO_418 (O_418,N_19814,N_19999);
nor UO_419 (O_419,N_19625,N_19882);
nand UO_420 (O_420,N_19890,N_19861);
xnor UO_421 (O_421,N_19997,N_19929);
nand UO_422 (O_422,N_19927,N_19992);
or UO_423 (O_423,N_19724,N_19791);
nand UO_424 (O_424,N_19645,N_19952);
xnor UO_425 (O_425,N_19708,N_19830);
xor UO_426 (O_426,N_19663,N_19688);
nand UO_427 (O_427,N_19956,N_19646);
nor UO_428 (O_428,N_19869,N_19649);
xnor UO_429 (O_429,N_19617,N_19890);
nand UO_430 (O_430,N_19693,N_19956);
and UO_431 (O_431,N_19995,N_19883);
nor UO_432 (O_432,N_19992,N_19943);
nand UO_433 (O_433,N_19783,N_19923);
or UO_434 (O_434,N_19954,N_19727);
nand UO_435 (O_435,N_19612,N_19981);
nor UO_436 (O_436,N_19717,N_19603);
xnor UO_437 (O_437,N_19895,N_19741);
and UO_438 (O_438,N_19979,N_19690);
or UO_439 (O_439,N_19894,N_19863);
nor UO_440 (O_440,N_19835,N_19996);
and UO_441 (O_441,N_19983,N_19659);
nand UO_442 (O_442,N_19695,N_19716);
nand UO_443 (O_443,N_19975,N_19882);
xor UO_444 (O_444,N_19992,N_19881);
xor UO_445 (O_445,N_19687,N_19696);
and UO_446 (O_446,N_19831,N_19904);
nor UO_447 (O_447,N_19627,N_19912);
nor UO_448 (O_448,N_19973,N_19978);
and UO_449 (O_449,N_19799,N_19945);
nand UO_450 (O_450,N_19741,N_19900);
and UO_451 (O_451,N_19648,N_19633);
nor UO_452 (O_452,N_19906,N_19635);
xnor UO_453 (O_453,N_19895,N_19612);
nand UO_454 (O_454,N_19761,N_19960);
nor UO_455 (O_455,N_19640,N_19919);
and UO_456 (O_456,N_19691,N_19912);
and UO_457 (O_457,N_19856,N_19873);
or UO_458 (O_458,N_19803,N_19980);
and UO_459 (O_459,N_19706,N_19731);
nor UO_460 (O_460,N_19921,N_19631);
nor UO_461 (O_461,N_19617,N_19704);
xor UO_462 (O_462,N_19762,N_19977);
or UO_463 (O_463,N_19805,N_19770);
nand UO_464 (O_464,N_19958,N_19856);
or UO_465 (O_465,N_19607,N_19795);
or UO_466 (O_466,N_19811,N_19737);
and UO_467 (O_467,N_19847,N_19733);
or UO_468 (O_468,N_19713,N_19953);
nand UO_469 (O_469,N_19936,N_19787);
or UO_470 (O_470,N_19703,N_19914);
xnor UO_471 (O_471,N_19707,N_19959);
nand UO_472 (O_472,N_19743,N_19643);
xnor UO_473 (O_473,N_19725,N_19798);
nor UO_474 (O_474,N_19826,N_19794);
nand UO_475 (O_475,N_19779,N_19926);
xor UO_476 (O_476,N_19983,N_19619);
nand UO_477 (O_477,N_19727,N_19918);
xor UO_478 (O_478,N_19658,N_19999);
nor UO_479 (O_479,N_19688,N_19839);
and UO_480 (O_480,N_19780,N_19834);
or UO_481 (O_481,N_19858,N_19728);
nand UO_482 (O_482,N_19947,N_19806);
nand UO_483 (O_483,N_19907,N_19672);
or UO_484 (O_484,N_19876,N_19685);
and UO_485 (O_485,N_19695,N_19623);
and UO_486 (O_486,N_19796,N_19995);
nor UO_487 (O_487,N_19931,N_19740);
nor UO_488 (O_488,N_19942,N_19697);
or UO_489 (O_489,N_19764,N_19671);
or UO_490 (O_490,N_19671,N_19860);
nand UO_491 (O_491,N_19913,N_19928);
and UO_492 (O_492,N_19717,N_19903);
xor UO_493 (O_493,N_19973,N_19619);
xor UO_494 (O_494,N_19934,N_19801);
nor UO_495 (O_495,N_19796,N_19872);
or UO_496 (O_496,N_19651,N_19945);
and UO_497 (O_497,N_19909,N_19783);
or UO_498 (O_498,N_19831,N_19618);
and UO_499 (O_499,N_19688,N_19995);
nand UO_500 (O_500,N_19710,N_19873);
nor UO_501 (O_501,N_19867,N_19831);
nor UO_502 (O_502,N_19699,N_19761);
nand UO_503 (O_503,N_19691,N_19904);
nand UO_504 (O_504,N_19977,N_19821);
or UO_505 (O_505,N_19657,N_19759);
and UO_506 (O_506,N_19821,N_19686);
nor UO_507 (O_507,N_19918,N_19913);
or UO_508 (O_508,N_19869,N_19822);
nand UO_509 (O_509,N_19973,N_19952);
nand UO_510 (O_510,N_19617,N_19832);
nand UO_511 (O_511,N_19675,N_19611);
or UO_512 (O_512,N_19923,N_19850);
or UO_513 (O_513,N_19958,N_19766);
nand UO_514 (O_514,N_19817,N_19987);
or UO_515 (O_515,N_19973,N_19927);
or UO_516 (O_516,N_19818,N_19754);
and UO_517 (O_517,N_19853,N_19795);
xnor UO_518 (O_518,N_19968,N_19919);
nand UO_519 (O_519,N_19874,N_19830);
or UO_520 (O_520,N_19661,N_19827);
nor UO_521 (O_521,N_19849,N_19819);
xnor UO_522 (O_522,N_19669,N_19609);
and UO_523 (O_523,N_19776,N_19718);
or UO_524 (O_524,N_19714,N_19729);
and UO_525 (O_525,N_19686,N_19865);
xor UO_526 (O_526,N_19926,N_19652);
and UO_527 (O_527,N_19979,N_19767);
or UO_528 (O_528,N_19617,N_19786);
xor UO_529 (O_529,N_19654,N_19900);
and UO_530 (O_530,N_19711,N_19957);
or UO_531 (O_531,N_19692,N_19824);
nor UO_532 (O_532,N_19758,N_19775);
nand UO_533 (O_533,N_19779,N_19897);
nor UO_534 (O_534,N_19858,N_19719);
nor UO_535 (O_535,N_19804,N_19707);
and UO_536 (O_536,N_19913,N_19948);
nor UO_537 (O_537,N_19987,N_19776);
or UO_538 (O_538,N_19722,N_19977);
and UO_539 (O_539,N_19869,N_19798);
nor UO_540 (O_540,N_19810,N_19965);
nor UO_541 (O_541,N_19854,N_19698);
nor UO_542 (O_542,N_19680,N_19753);
and UO_543 (O_543,N_19767,N_19650);
nor UO_544 (O_544,N_19835,N_19603);
nand UO_545 (O_545,N_19645,N_19709);
xnor UO_546 (O_546,N_19752,N_19974);
and UO_547 (O_547,N_19697,N_19810);
nand UO_548 (O_548,N_19930,N_19643);
nor UO_549 (O_549,N_19694,N_19982);
xnor UO_550 (O_550,N_19797,N_19834);
or UO_551 (O_551,N_19671,N_19692);
or UO_552 (O_552,N_19819,N_19921);
nor UO_553 (O_553,N_19801,N_19682);
or UO_554 (O_554,N_19847,N_19868);
or UO_555 (O_555,N_19795,N_19965);
xor UO_556 (O_556,N_19686,N_19676);
or UO_557 (O_557,N_19771,N_19649);
and UO_558 (O_558,N_19629,N_19830);
and UO_559 (O_559,N_19950,N_19628);
xnor UO_560 (O_560,N_19784,N_19887);
nand UO_561 (O_561,N_19729,N_19942);
nor UO_562 (O_562,N_19893,N_19863);
or UO_563 (O_563,N_19965,N_19908);
xnor UO_564 (O_564,N_19985,N_19975);
and UO_565 (O_565,N_19724,N_19779);
or UO_566 (O_566,N_19835,N_19656);
nand UO_567 (O_567,N_19707,N_19908);
xnor UO_568 (O_568,N_19967,N_19899);
nand UO_569 (O_569,N_19688,N_19755);
nor UO_570 (O_570,N_19816,N_19682);
nor UO_571 (O_571,N_19980,N_19641);
nand UO_572 (O_572,N_19855,N_19682);
nor UO_573 (O_573,N_19608,N_19710);
or UO_574 (O_574,N_19815,N_19716);
xor UO_575 (O_575,N_19826,N_19725);
or UO_576 (O_576,N_19906,N_19961);
xor UO_577 (O_577,N_19678,N_19784);
and UO_578 (O_578,N_19638,N_19881);
nor UO_579 (O_579,N_19712,N_19751);
and UO_580 (O_580,N_19705,N_19754);
and UO_581 (O_581,N_19908,N_19914);
and UO_582 (O_582,N_19900,N_19601);
and UO_583 (O_583,N_19781,N_19821);
nand UO_584 (O_584,N_19834,N_19632);
nand UO_585 (O_585,N_19654,N_19980);
nand UO_586 (O_586,N_19802,N_19744);
or UO_587 (O_587,N_19855,N_19769);
nor UO_588 (O_588,N_19922,N_19679);
nand UO_589 (O_589,N_19701,N_19725);
and UO_590 (O_590,N_19767,N_19693);
nor UO_591 (O_591,N_19853,N_19934);
xnor UO_592 (O_592,N_19963,N_19792);
nor UO_593 (O_593,N_19772,N_19972);
and UO_594 (O_594,N_19692,N_19892);
nor UO_595 (O_595,N_19848,N_19637);
xor UO_596 (O_596,N_19755,N_19608);
or UO_597 (O_597,N_19731,N_19734);
and UO_598 (O_598,N_19624,N_19999);
nand UO_599 (O_599,N_19806,N_19799);
and UO_600 (O_600,N_19670,N_19816);
and UO_601 (O_601,N_19709,N_19730);
and UO_602 (O_602,N_19916,N_19849);
nor UO_603 (O_603,N_19846,N_19723);
or UO_604 (O_604,N_19904,N_19644);
or UO_605 (O_605,N_19716,N_19840);
xor UO_606 (O_606,N_19987,N_19834);
or UO_607 (O_607,N_19815,N_19945);
and UO_608 (O_608,N_19673,N_19613);
and UO_609 (O_609,N_19959,N_19690);
nor UO_610 (O_610,N_19785,N_19685);
nand UO_611 (O_611,N_19777,N_19836);
xor UO_612 (O_612,N_19810,N_19933);
xor UO_613 (O_613,N_19642,N_19996);
or UO_614 (O_614,N_19880,N_19839);
nor UO_615 (O_615,N_19845,N_19615);
nor UO_616 (O_616,N_19915,N_19634);
nor UO_617 (O_617,N_19862,N_19601);
nor UO_618 (O_618,N_19914,N_19618);
nor UO_619 (O_619,N_19744,N_19674);
and UO_620 (O_620,N_19728,N_19937);
xnor UO_621 (O_621,N_19644,N_19958);
nand UO_622 (O_622,N_19789,N_19607);
xor UO_623 (O_623,N_19689,N_19764);
nor UO_624 (O_624,N_19797,N_19705);
or UO_625 (O_625,N_19743,N_19899);
nor UO_626 (O_626,N_19861,N_19941);
nand UO_627 (O_627,N_19817,N_19898);
or UO_628 (O_628,N_19756,N_19872);
nand UO_629 (O_629,N_19839,N_19647);
nand UO_630 (O_630,N_19884,N_19749);
nor UO_631 (O_631,N_19666,N_19662);
or UO_632 (O_632,N_19692,N_19658);
xnor UO_633 (O_633,N_19967,N_19870);
or UO_634 (O_634,N_19704,N_19804);
xnor UO_635 (O_635,N_19795,N_19929);
and UO_636 (O_636,N_19988,N_19781);
nor UO_637 (O_637,N_19867,N_19728);
nor UO_638 (O_638,N_19858,N_19996);
or UO_639 (O_639,N_19855,N_19979);
xor UO_640 (O_640,N_19823,N_19928);
nand UO_641 (O_641,N_19641,N_19777);
or UO_642 (O_642,N_19879,N_19945);
nand UO_643 (O_643,N_19959,N_19970);
nor UO_644 (O_644,N_19671,N_19870);
and UO_645 (O_645,N_19874,N_19837);
nor UO_646 (O_646,N_19644,N_19613);
xnor UO_647 (O_647,N_19990,N_19848);
xor UO_648 (O_648,N_19975,N_19648);
or UO_649 (O_649,N_19754,N_19790);
or UO_650 (O_650,N_19805,N_19736);
nor UO_651 (O_651,N_19859,N_19642);
nand UO_652 (O_652,N_19834,N_19859);
and UO_653 (O_653,N_19619,N_19884);
xnor UO_654 (O_654,N_19601,N_19921);
or UO_655 (O_655,N_19638,N_19954);
and UO_656 (O_656,N_19909,N_19620);
nand UO_657 (O_657,N_19779,N_19879);
and UO_658 (O_658,N_19681,N_19866);
nand UO_659 (O_659,N_19962,N_19908);
or UO_660 (O_660,N_19609,N_19855);
xnor UO_661 (O_661,N_19714,N_19607);
xnor UO_662 (O_662,N_19888,N_19880);
and UO_663 (O_663,N_19679,N_19719);
or UO_664 (O_664,N_19950,N_19826);
nor UO_665 (O_665,N_19820,N_19965);
and UO_666 (O_666,N_19677,N_19673);
xor UO_667 (O_667,N_19842,N_19636);
or UO_668 (O_668,N_19787,N_19923);
or UO_669 (O_669,N_19976,N_19733);
or UO_670 (O_670,N_19890,N_19741);
nand UO_671 (O_671,N_19774,N_19666);
and UO_672 (O_672,N_19996,N_19892);
or UO_673 (O_673,N_19918,N_19915);
or UO_674 (O_674,N_19624,N_19813);
nor UO_675 (O_675,N_19850,N_19941);
xor UO_676 (O_676,N_19792,N_19790);
nand UO_677 (O_677,N_19831,N_19783);
and UO_678 (O_678,N_19943,N_19890);
or UO_679 (O_679,N_19863,N_19690);
nand UO_680 (O_680,N_19782,N_19870);
nor UO_681 (O_681,N_19682,N_19735);
nand UO_682 (O_682,N_19659,N_19721);
nand UO_683 (O_683,N_19801,N_19609);
and UO_684 (O_684,N_19877,N_19942);
xor UO_685 (O_685,N_19952,N_19979);
nand UO_686 (O_686,N_19986,N_19858);
nor UO_687 (O_687,N_19898,N_19637);
nor UO_688 (O_688,N_19811,N_19977);
nor UO_689 (O_689,N_19775,N_19810);
and UO_690 (O_690,N_19867,N_19991);
or UO_691 (O_691,N_19888,N_19994);
and UO_692 (O_692,N_19805,N_19661);
or UO_693 (O_693,N_19830,N_19709);
xor UO_694 (O_694,N_19717,N_19790);
nor UO_695 (O_695,N_19779,N_19923);
or UO_696 (O_696,N_19685,N_19914);
nor UO_697 (O_697,N_19815,N_19640);
nor UO_698 (O_698,N_19733,N_19640);
and UO_699 (O_699,N_19982,N_19799);
and UO_700 (O_700,N_19962,N_19794);
nand UO_701 (O_701,N_19730,N_19889);
nand UO_702 (O_702,N_19777,N_19944);
xor UO_703 (O_703,N_19611,N_19761);
nand UO_704 (O_704,N_19739,N_19632);
nand UO_705 (O_705,N_19928,N_19937);
and UO_706 (O_706,N_19933,N_19749);
nor UO_707 (O_707,N_19748,N_19830);
and UO_708 (O_708,N_19794,N_19745);
nor UO_709 (O_709,N_19606,N_19868);
nor UO_710 (O_710,N_19878,N_19773);
nand UO_711 (O_711,N_19787,N_19916);
nor UO_712 (O_712,N_19944,N_19880);
or UO_713 (O_713,N_19833,N_19665);
and UO_714 (O_714,N_19610,N_19666);
xnor UO_715 (O_715,N_19971,N_19747);
and UO_716 (O_716,N_19764,N_19740);
xor UO_717 (O_717,N_19921,N_19804);
nand UO_718 (O_718,N_19642,N_19774);
xnor UO_719 (O_719,N_19733,N_19791);
nor UO_720 (O_720,N_19940,N_19980);
nand UO_721 (O_721,N_19917,N_19637);
nor UO_722 (O_722,N_19839,N_19803);
xnor UO_723 (O_723,N_19871,N_19863);
and UO_724 (O_724,N_19829,N_19657);
or UO_725 (O_725,N_19704,N_19602);
and UO_726 (O_726,N_19647,N_19973);
nor UO_727 (O_727,N_19940,N_19918);
nor UO_728 (O_728,N_19918,N_19987);
or UO_729 (O_729,N_19731,N_19777);
xnor UO_730 (O_730,N_19795,N_19650);
or UO_731 (O_731,N_19615,N_19702);
or UO_732 (O_732,N_19909,N_19675);
or UO_733 (O_733,N_19964,N_19922);
or UO_734 (O_734,N_19878,N_19886);
nand UO_735 (O_735,N_19888,N_19853);
xor UO_736 (O_736,N_19648,N_19900);
and UO_737 (O_737,N_19655,N_19976);
or UO_738 (O_738,N_19702,N_19935);
xor UO_739 (O_739,N_19796,N_19903);
nand UO_740 (O_740,N_19617,N_19764);
or UO_741 (O_741,N_19704,N_19957);
nor UO_742 (O_742,N_19954,N_19882);
nand UO_743 (O_743,N_19607,N_19797);
nand UO_744 (O_744,N_19796,N_19880);
nor UO_745 (O_745,N_19928,N_19737);
nor UO_746 (O_746,N_19836,N_19956);
xor UO_747 (O_747,N_19655,N_19944);
nand UO_748 (O_748,N_19871,N_19984);
nand UO_749 (O_749,N_19990,N_19742);
or UO_750 (O_750,N_19898,N_19857);
nor UO_751 (O_751,N_19998,N_19728);
or UO_752 (O_752,N_19870,N_19657);
or UO_753 (O_753,N_19638,N_19652);
and UO_754 (O_754,N_19620,N_19759);
xnor UO_755 (O_755,N_19850,N_19765);
and UO_756 (O_756,N_19607,N_19822);
and UO_757 (O_757,N_19686,N_19944);
and UO_758 (O_758,N_19600,N_19757);
nor UO_759 (O_759,N_19997,N_19901);
nor UO_760 (O_760,N_19705,N_19670);
nand UO_761 (O_761,N_19694,N_19734);
nand UO_762 (O_762,N_19966,N_19900);
xor UO_763 (O_763,N_19617,N_19607);
nor UO_764 (O_764,N_19776,N_19703);
and UO_765 (O_765,N_19667,N_19963);
or UO_766 (O_766,N_19669,N_19972);
and UO_767 (O_767,N_19780,N_19736);
nand UO_768 (O_768,N_19792,N_19610);
nand UO_769 (O_769,N_19999,N_19873);
nand UO_770 (O_770,N_19972,N_19842);
and UO_771 (O_771,N_19771,N_19867);
or UO_772 (O_772,N_19814,N_19975);
or UO_773 (O_773,N_19765,N_19913);
or UO_774 (O_774,N_19763,N_19952);
nand UO_775 (O_775,N_19975,N_19970);
xnor UO_776 (O_776,N_19995,N_19939);
nor UO_777 (O_777,N_19678,N_19605);
and UO_778 (O_778,N_19730,N_19959);
or UO_779 (O_779,N_19817,N_19976);
nand UO_780 (O_780,N_19611,N_19926);
nand UO_781 (O_781,N_19757,N_19789);
nor UO_782 (O_782,N_19895,N_19832);
or UO_783 (O_783,N_19925,N_19996);
or UO_784 (O_784,N_19630,N_19739);
xor UO_785 (O_785,N_19634,N_19809);
or UO_786 (O_786,N_19954,N_19866);
nor UO_787 (O_787,N_19617,N_19870);
nand UO_788 (O_788,N_19922,N_19689);
nand UO_789 (O_789,N_19773,N_19684);
xor UO_790 (O_790,N_19663,N_19818);
xor UO_791 (O_791,N_19644,N_19893);
nor UO_792 (O_792,N_19605,N_19909);
nand UO_793 (O_793,N_19939,N_19800);
or UO_794 (O_794,N_19704,N_19885);
xnor UO_795 (O_795,N_19765,N_19862);
nor UO_796 (O_796,N_19739,N_19884);
or UO_797 (O_797,N_19802,N_19719);
or UO_798 (O_798,N_19998,N_19922);
and UO_799 (O_799,N_19855,N_19821);
and UO_800 (O_800,N_19678,N_19857);
xor UO_801 (O_801,N_19640,N_19686);
nand UO_802 (O_802,N_19832,N_19911);
or UO_803 (O_803,N_19814,N_19691);
or UO_804 (O_804,N_19827,N_19928);
xnor UO_805 (O_805,N_19787,N_19963);
or UO_806 (O_806,N_19963,N_19628);
nor UO_807 (O_807,N_19949,N_19800);
or UO_808 (O_808,N_19910,N_19955);
nor UO_809 (O_809,N_19626,N_19666);
or UO_810 (O_810,N_19957,N_19756);
and UO_811 (O_811,N_19951,N_19616);
nand UO_812 (O_812,N_19705,N_19896);
or UO_813 (O_813,N_19726,N_19830);
or UO_814 (O_814,N_19702,N_19963);
nand UO_815 (O_815,N_19965,N_19982);
nor UO_816 (O_816,N_19605,N_19830);
nand UO_817 (O_817,N_19798,N_19827);
and UO_818 (O_818,N_19723,N_19789);
nor UO_819 (O_819,N_19703,N_19609);
xnor UO_820 (O_820,N_19607,N_19738);
nor UO_821 (O_821,N_19846,N_19978);
nand UO_822 (O_822,N_19829,N_19636);
or UO_823 (O_823,N_19689,N_19645);
or UO_824 (O_824,N_19989,N_19655);
nand UO_825 (O_825,N_19868,N_19796);
nand UO_826 (O_826,N_19709,N_19996);
xnor UO_827 (O_827,N_19742,N_19715);
xor UO_828 (O_828,N_19821,N_19983);
nand UO_829 (O_829,N_19698,N_19957);
nand UO_830 (O_830,N_19973,N_19753);
nand UO_831 (O_831,N_19808,N_19663);
and UO_832 (O_832,N_19942,N_19926);
and UO_833 (O_833,N_19687,N_19804);
xnor UO_834 (O_834,N_19977,N_19708);
nand UO_835 (O_835,N_19839,N_19958);
xor UO_836 (O_836,N_19610,N_19841);
and UO_837 (O_837,N_19997,N_19854);
and UO_838 (O_838,N_19882,N_19859);
and UO_839 (O_839,N_19690,N_19825);
nand UO_840 (O_840,N_19820,N_19895);
nand UO_841 (O_841,N_19920,N_19891);
nor UO_842 (O_842,N_19904,N_19945);
nor UO_843 (O_843,N_19885,N_19978);
and UO_844 (O_844,N_19614,N_19832);
nor UO_845 (O_845,N_19943,N_19610);
nand UO_846 (O_846,N_19757,N_19623);
xnor UO_847 (O_847,N_19744,N_19675);
or UO_848 (O_848,N_19855,N_19919);
and UO_849 (O_849,N_19639,N_19658);
nand UO_850 (O_850,N_19987,N_19944);
nor UO_851 (O_851,N_19655,N_19630);
xnor UO_852 (O_852,N_19604,N_19779);
and UO_853 (O_853,N_19974,N_19977);
nor UO_854 (O_854,N_19642,N_19626);
nor UO_855 (O_855,N_19741,N_19775);
and UO_856 (O_856,N_19812,N_19750);
and UO_857 (O_857,N_19981,N_19939);
and UO_858 (O_858,N_19923,N_19668);
xor UO_859 (O_859,N_19620,N_19847);
and UO_860 (O_860,N_19786,N_19613);
and UO_861 (O_861,N_19706,N_19878);
xor UO_862 (O_862,N_19601,N_19788);
and UO_863 (O_863,N_19746,N_19839);
or UO_864 (O_864,N_19728,N_19859);
xor UO_865 (O_865,N_19845,N_19758);
nor UO_866 (O_866,N_19752,N_19715);
xnor UO_867 (O_867,N_19889,N_19822);
nand UO_868 (O_868,N_19692,N_19915);
xor UO_869 (O_869,N_19969,N_19669);
or UO_870 (O_870,N_19849,N_19782);
nor UO_871 (O_871,N_19752,N_19724);
and UO_872 (O_872,N_19828,N_19935);
and UO_873 (O_873,N_19889,N_19833);
and UO_874 (O_874,N_19755,N_19876);
or UO_875 (O_875,N_19883,N_19781);
or UO_876 (O_876,N_19903,N_19712);
nor UO_877 (O_877,N_19657,N_19925);
or UO_878 (O_878,N_19665,N_19927);
nand UO_879 (O_879,N_19660,N_19853);
and UO_880 (O_880,N_19951,N_19996);
or UO_881 (O_881,N_19622,N_19893);
or UO_882 (O_882,N_19974,N_19779);
or UO_883 (O_883,N_19895,N_19748);
xnor UO_884 (O_884,N_19636,N_19805);
nor UO_885 (O_885,N_19934,N_19870);
nor UO_886 (O_886,N_19866,N_19811);
xnor UO_887 (O_887,N_19645,N_19767);
xnor UO_888 (O_888,N_19627,N_19877);
nand UO_889 (O_889,N_19898,N_19946);
nor UO_890 (O_890,N_19889,N_19613);
xor UO_891 (O_891,N_19682,N_19664);
or UO_892 (O_892,N_19893,N_19945);
xor UO_893 (O_893,N_19667,N_19680);
xnor UO_894 (O_894,N_19741,N_19837);
or UO_895 (O_895,N_19776,N_19723);
nand UO_896 (O_896,N_19725,N_19755);
xor UO_897 (O_897,N_19747,N_19636);
nor UO_898 (O_898,N_19838,N_19866);
or UO_899 (O_899,N_19995,N_19659);
and UO_900 (O_900,N_19893,N_19719);
nand UO_901 (O_901,N_19728,N_19838);
and UO_902 (O_902,N_19662,N_19904);
or UO_903 (O_903,N_19818,N_19771);
or UO_904 (O_904,N_19603,N_19648);
xor UO_905 (O_905,N_19760,N_19774);
nor UO_906 (O_906,N_19705,N_19736);
xor UO_907 (O_907,N_19967,N_19812);
nor UO_908 (O_908,N_19799,N_19913);
and UO_909 (O_909,N_19931,N_19697);
nor UO_910 (O_910,N_19622,N_19804);
xor UO_911 (O_911,N_19747,N_19607);
nand UO_912 (O_912,N_19800,N_19906);
or UO_913 (O_913,N_19671,N_19965);
nor UO_914 (O_914,N_19936,N_19754);
nor UO_915 (O_915,N_19841,N_19634);
xnor UO_916 (O_916,N_19918,N_19909);
nand UO_917 (O_917,N_19983,N_19882);
or UO_918 (O_918,N_19627,N_19958);
xnor UO_919 (O_919,N_19693,N_19862);
nand UO_920 (O_920,N_19835,N_19999);
nor UO_921 (O_921,N_19786,N_19873);
and UO_922 (O_922,N_19681,N_19754);
or UO_923 (O_923,N_19626,N_19913);
nand UO_924 (O_924,N_19764,N_19687);
nor UO_925 (O_925,N_19928,N_19701);
xor UO_926 (O_926,N_19691,N_19649);
nand UO_927 (O_927,N_19785,N_19877);
nor UO_928 (O_928,N_19666,N_19851);
nand UO_929 (O_929,N_19809,N_19603);
and UO_930 (O_930,N_19864,N_19821);
or UO_931 (O_931,N_19806,N_19751);
and UO_932 (O_932,N_19624,N_19857);
xnor UO_933 (O_933,N_19875,N_19751);
or UO_934 (O_934,N_19698,N_19650);
nor UO_935 (O_935,N_19672,N_19736);
and UO_936 (O_936,N_19672,N_19819);
and UO_937 (O_937,N_19980,N_19668);
xor UO_938 (O_938,N_19611,N_19835);
nor UO_939 (O_939,N_19661,N_19747);
or UO_940 (O_940,N_19853,N_19931);
xnor UO_941 (O_941,N_19641,N_19811);
and UO_942 (O_942,N_19872,N_19699);
and UO_943 (O_943,N_19709,N_19706);
and UO_944 (O_944,N_19915,N_19816);
xnor UO_945 (O_945,N_19722,N_19696);
nand UO_946 (O_946,N_19917,N_19726);
nor UO_947 (O_947,N_19991,N_19872);
and UO_948 (O_948,N_19851,N_19805);
xor UO_949 (O_949,N_19912,N_19724);
nor UO_950 (O_950,N_19704,N_19768);
or UO_951 (O_951,N_19877,N_19920);
nand UO_952 (O_952,N_19910,N_19871);
nand UO_953 (O_953,N_19874,N_19919);
nor UO_954 (O_954,N_19952,N_19641);
nor UO_955 (O_955,N_19966,N_19995);
or UO_956 (O_956,N_19946,N_19888);
nand UO_957 (O_957,N_19619,N_19936);
xnor UO_958 (O_958,N_19963,N_19882);
or UO_959 (O_959,N_19768,N_19736);
xor UO_960 (O_960,N_19723,N_19839);
and UO_961 (O_961,N_19734,N_19785);
and UO_962 (O_962,N_19933,N_19708);
nand UO_963 (O_963,N_19655,N_19678);
nor UO_964 (O_964,N_19804,N_19815);
or UO_965 (O_965,N_19697,N_19772);
nor UO_966 (O_966,N_19626,N_19994);
nand UO_967 (O_967,N_19946,N_19803);
nor UO_968 (O_968,N_19807,N_19765);
xor UO_969 (O_969,N_19931,N_19714);
xor UO_970 (O_970,N_19675,N_19736);
nand UO_971 (O_971,N_19921,N_19613);
nand UO_972 (O_972,N_19729,N_19783);
nand UO_973 (O_973,N_19767,N_19757);
nand UO_974 (O_974,N_19609,N_19870);
nor UO_975 (O_975,N_19682,N_19692);
nor UO_976 (O_976,N_19859,N_19856);
or UO_977 (O_977,N_19671,N_19719);
nand UO_978 (O_978,N_19890,N_19678);
nand UO_979 (O_979,N_19764,N_19802);
nor UO_980 (O_980,N_19872,N_19636);
nor UO_981 (O_981,N_19667,N_19687);
or UO_982 (O_982,N_19828,N_19963);
nor UO_983 (O_983,N_19841,N_19778);
nand UO_984 (O_984,N_19614,N_19954);
nor UO_985 (O_985,N_19903,N_19735);
xor UO_986 (O_986,N_19931,N_19707);
xnor UO_987 (O_987,N_19971,N_19895);
and UO_988 (O_988,N_19984,N_19674);
and UO_989 (O_989,N_19735,N_19624);
nor UO_990 (O_990,N_19868,N_19913);
nand UO_991 (O_991,N_19875,N_19864);
xnor UO_992 (O_992,N_19765,N_19968);
nand UO_993 (O_993,N_19839,N_19760);
nor UO_994 (O_994,N_19919,N_19864);
xor UO_995 (O_995,N_19900,N_19883);
xor UO_996 (O_996,N_19799,N_19702);
xnor UO_997 (O_997,N_19838,N_19620);
xnor UO_998 (O_998,N_19918,N_19944);
nor UO_999 (O_999,N_19922,N_19741);
xnor UO_1000 (O_1000,N_19799,N_19881);
nand UO_1001 (O_1001,N_19787,N_19732);
and UO_1002 (O_1002,N_19803,N_19617);
and UO_1003 (O_1003,N_19674,N_19909);
or UO_1004 (O_1004,N_19906,N_19720);
nor UO_1005 (O_1005,N_19723,N_19637);
nor UO_1006 (O_1006,N_19764,N_19652);
nand UO_1007 (O_1007,N_19891,N_19939);
xor UO_1008 (O_1008,N_19627,N_19778);
or UO_1009 (O_1009,N_19950,N_19716);
nor UO_1010 (O_1010,N_19737,N_19671);
or UO_1011 (O_1011,N_19659,N_19851);
xor UO_1012 (O_1012,N_19609,N_19808);
and UO_1013 (O_1013,N_19946,N_19960);
nor UO_1014 (O_1014,N_19839,N_19854);
or UO_1015 (O_1015,N_19957,N_19822);
nand UO_1016 (O_1016,N_19649,N_19959);
or UO_1017 (O_1017,N_19603,N_19871);
nand UO_1018 (O_1018,N_19678,N_19834);
and UO_1019 (O_1019,N_19836,N_19940);
or UO_1020 (O_1020,N_19781,N_19658);
nor UO_1021 (O_1021,N_19667,N_19632);
nand UO_1022 (O_1022,N_19710,N_19793);
and UO_1023 (O_1023,N_19652,N_19706);
or UO_1024 (O_1024,N_19895,N_19969);
nor UO_1025 (O_1025,N_19994,N_19965);
or UO_1026 (O_1026,N_19920,N_19655);
and UO_1027 (O_1027,N_19721,N_19934);
xor UO_1028 (O_1028,N_19876,N_19723);
xor UO_1029 (O_1029,N_19813,N_19879);
nor UO_1030 (O_1030,N_19732,N_19854);
or UO_1031 (O_1031,N_19831,N_19979);
xnor UO_1032 (O_1032,N_19603,N_19908);
nand UO_1033 (O_1033,N_19776,N_19726);
and UO_1034 (O_1034,N_19703,N_19725);
xnor UO_1035 (O_1035,N_19756,N_19616);
nand UO_1036 (O_1036,N_19654,N_19875);
nor UO_1037 (O_1037,N_19654,N_19901);
and UO_1038 (O_1038,N_19754,N_19676);
or UO_1039 (O_1039,N_19699,N_19836);
or UO_1040 (O_1040,N_19679,N_19704);
nor UO_1041 (O_1041,N_19662,N_19807);
nand UO_1042 (O_1042,N_19741,N_19762);
and UO_1043 (O_1043,N_19854,N_19878);
nor UO_1044 (O_1044,N_19876,N_19671);
nor UO_1045 (O_1045,N_19673,N_19745);
and UO_1046 (O_1046,N_19941,N_19665);
and UO_1047 (O_1047,N_19699,N_19624);
xnor UO_1048 (O_1048,N_19971,N_19922);
nand UO_1049 (O_1049,N_19903,N_19944);
nand UO_1050 (O_1050,N_19658,N_19976);
and UO_1051 (O_1051,N_19641,N_19971);
nor UO_1052 (O_1052,N_19713,N_19667);
and UO_1053 (O_1053,N_19679,N_19945);
and UO_1054 (O_1054,N_19606,N_19654);
nor UO_1055 (O_1055,N_19913,N_19941);
nor UO_1056 (O_1056,N_19970,N_19868);
and UO_1057 (O_1057,N_19798,N_19876);
or UO_1058 (O_1058,N_19739,N_19754);
xor UO_1059 (O_1059,N_19835,N_19859);
nor UO_1060 (O_1060,N_19643,N_19690);
xnor UO_1061 (O_1061,N_19764,N_19829);
and UO_1062 (O_1062,N_19924,N_19843);
nor UO_1063 (O_1063,N_19818,N_19936);
nor UO_1064 (O_1064,N_19946,N_19750);
and UO_1065 (O_1065,N_19616,N_19978);
xor UO_1066 (O_1066,N_19653,N_19747);
nand UO_1067 (O_1067,N_19841,N_19601);
or UO_1068 (O_1068,N_19989,N_19852);
nor UO_1069 (O_1069,N_19717,N_19894);
nand UO_1070 (O_1070,N_19657,N_19907);
nand UO_1071 (O_1071,N_19979,N_19771);
or UO_1072 (O_1072,N_19785,N_19724);
nor UO_1073 (O_1073,N_19853,N_19993);
or UO_1074 (O_1074,N_19885,N_19710);
or UO_1075 (O_1075,N_19847,N_19732);
nand UO_1076 (O_1076,N_19640,N_19737);
and UO_1077 (O_1077,N_19717,N_19699);
and UO_1078 (O_1078,N_19727,N_19634);
nand UO_1079 (O_1079,N_19977,N_19655);
nand UO_1080 (O_1080,N_19902,N_19794);
and UO_1081 (O_1081,N_19980,N_19782);
or UO_1082 (O_1082,N_19882,N_19614);
xnor UO_1083 (O_1083,N_19825,N_19742);
and UO_1084 (O_1084,N_19991,N_19848);
nand UO_1085 (O_1085,N_19721,N_19798);
and UO_1086 (O_1086,N_19798,N_19803);
nand UO_1087 (O_1087,N_19649,N_19667);
nand UO_1088 (O_1088,N_19636,N_19646);
nand UO_1089 (O_1089,N_19781,N_19753);
or UO_1090 (O_1090,N_19837,N_19716);
xnor UO_1091 (O_1091,N_19884,N_19692);
nand UO_1092 (O_1092,N_19687,N_19928);
and UO_1093 (O_1093,N_19941,N_19718);
nor UO_1094 (O_1094,N_19817,N_19671);
or UO_1095 (O_1095,N_19795,N_19733);
or UO_1096 (O_1096,N_19825,N_19693);
nand UO_1097 (O_1097,N_19887,N_19814);
xnor UO_1098 (O_1098,N_19810,N_19796);
or UO_1099 (O_1099,N_19646,N_19801);
nand UO_1100 (O_1100,N_19963,N_19837);
xor UO_1101 (O_1101,N_19671,N_19659);
nor UO_1102 (O_1102,N_19653,N_19944);
nor UO_1103 (O_1103,N_19819,N_19762);
or UO_1104 (O_1104,N_19686,N_19985);
xnor UO_1105 (O_1105,N_19713,N_19710);
and UO_1106 (O_1106,N_19666,N_19806);
xnor UO_1107 (O_1107,N_19825,N_19967);
and UO_1108 (O_1108,N_19643,N_19797);
and UO_1109 (O_1109,N_19901,N_19608);
nand UO_1110 (O_1110,N_19888,N_19808);
and UO_1111 (O_1111,N_19949,N_19884);
xnor UO_1112 (O_1112,N_19833,N_19637);
nand UO_1113 (O_1113,N_19741,N_19924);
nand UO_1114 (O_1114,N_19908,N_19616);
nand UO_1115 (O_1115,N_19852,N_19802);
or UO_1116 (O_1116,N_19960,N_19619);
and UO_1117 (O_1117,N_19868,N_19703);
xor UO_1118 (O_1118,N_19706,N_19781);
or UO_1119 (O_1119,N_19726,N_19827);
or UO_1120 (O_1120,N_19751,N_19771);
nand UO_1121 (O_1121,N_19740,N_19981);
nand UO_1122 (O_1122,N_19800,N_19994);
or UO_1123 (O_1123,N_19702,N_19755);
or UO_1124 (O_1124,N_19906,N_19930);
nor UO_1125 (O_1125,N_19892,N_19897);
nand UO_1126 (O_1126,N_19772,N_19950);
nand UO_1127 (O_1127,N_19613,N_19955);
xor UO_1128 (O_1128,N_19682,N_19944);
nor UO_1129 (O_1129,N_19776,N_19877);
or UO_1130 (O_1130,N_19951,N_19781);
xor UO_1131 (O_1131,N_19940,N_19745);
or UO_1132 (O_1132,N_19620,N_19659);
nor UO_1133 (O_1133,N_19938,N_19825);
nand UO_1134 (O_1134,N_19760,N_19814);
nand UO_1135 (O_1135,N_19917,N_19727);
nor UO_1136 (O_1136,N_19959,N_19617);
or UO_1137 (O_1137,N_19682,N_19600);
nor UO_1138 (O_1138,N_19779,N_19686);
nand UO_1139 (O_1139,N_19954,N_19619);
xor UO_1140 (O_1140,N_19839,N_19670);
or UO_1141 (O_1141,N_19618,N_19753);
nand UO_1142 (O_1142,N_19712,N_19607);
or UO_1143 (O_1143,N_19998,N_19877);
nand UO_1144 (O_1144,N_19868,N_19699);
nand UO_1145 (O_1145,N_19768,N_19771);
nand UO_1146 (O_1146,N_19638,N_19837);
nor UO_1147 (O_1147,N_19801,N_19908);
and UO_1148 (O_1148,N_19670,N_19975);
or UO_1149 (O_1149,N_19717,N_19608);
nor UO_1150 (O_1150,N_19658,N_19843);
and UO_1151 (O_1151,N_19888,N_19814);
xor UO_1152 (O_1152,N_19646,N_19656);
and UO_1153 (O_1153,N_19692,N_19999);
nor UO_1154 (O_1154,N_19950,N_19889);
nand UO_1155 (O_1155,N_19665,N_19988);
xnor UO_1156 (O_1156,N_19831,N_19739);
and UO_1157 (O_1157,N_19718,N_19618);
nand UO_1158 (O_1158,N_19615,N_19719);
or UO_1159 (O_1159,N_19824,N_19815);
nand UO_1160 (O_1160,N_19652,N_19757);
or UO_1161 (O_1161,N_19796,N_19876);
and UO_1162 (O_1162,N_19765,N_19881);
xor UO_1163 (O_1163,N_19838,N_19670);
or UO_1164 (O_1164,N_19852,N_19687);
and UO_1165 (O_1165,N_19734,N_19797);
nand UO_1166 (O_1166,N_19870,N_19653);
nand UO_1167 (O_1167,N_19712,N_19678);
nor UO_1168 (O_1168,N_19648,N_19925);
nor UO_1169 (O_1169,N_19867,N_19822);
and UO_1170 (O_1170,N_19692,N_19921);
nor UO_1171 (O_1171,N_19668,N_19710);
and UO_1172 (O_1172,N_19717,N_19973);
nand UO_1173 (O_1173,N_19709,N_19849);
or UO_1174 (O_1174,N_19862,N_19958);
or UO_1175 (O_1175,N_19797,N_19713);
and UO_1176 (O_1176,N_19735,N_19656);
nand UO_1177 (O_1177,N_19813,N_19912);
nor UO_1178 (O_1178,N_19835,N_19953);
xnor UO_1179 (O_1179,N_19690,N_19775);
or UO_1180 (O_1180,N_19800,N_19987);
xor UO_1181 (O_1181,N_19802,N_19781);
nand UO_1182 (O_1182,N_19701,N_19958);
or UO_1183 (O_1183,N_19665,N_19618);
and UO_1184 (O_1184,N_19689,N_19917);
nor UO_1185 (O_1185,N_19800,N_19928);
or UO_1186 (O_1186,N_19996,N_19635);
and UO_1187 (O_1187,N_19841,N_19743);
nand UO_1188 (O_1188,N_19979,N_19808);
or UO_1189 (O_1189,N_19913,N_19980);
nand UO_1190 (O_1190,N_19751,N_19717);
or UO_1191 (O_1191,N_19756,N_19733);
and UO_1192 (O_1192,N_19964,N_19981);
or UO_1193 (O_1193,N_19846,N_19633);
nand UO_1194 (O_1194,N_19907,N_19977);
nand UO_1195 (O_1195,N_19990,N_19992);
nor UO_1196 (O_1196,N_19905,N_19681);
or UO_1197 (O_1197,N_19983,N_19995);
nand UO_1198 (O_1198,N_19976,N_19859);
and UO_1199 (O_1199,N_19908,N_19618);
or UO_1200 (O_1200,N_19877,N_19777);
and UO_1201 (O_1201,N_19984,N_19823);
xor UO_1202 (O_1202,N_19859,N_19645);
and UO_1203 (O_1203,N_19740,N_19886);
nor UO_1204 (O_1204,N_19619,N_19986);
nor UO_1205 (O_1205,N_19914,N_19878);
xnor UO_1206 (O_1206,N_19786,N_19876);
nor UO_1207 (O_1207,N_19826,N_19956);
nand UO_1208 (O_1208,N_19953,N_19666);
nand UO_1209 (O_1209,N_19614,N_19933);
xnor UO_1210 (O_1210,N_19681,N_19982);
nand UO_1211 (O_1211,N_19787,N_19685);
or UO_1212 (O_1212,N_19733,N_19886);
and UO_1213 (O_1213,N_19697,N_19639);
nor UO_1214 (O_1214,N_19977,N_19804);
nand UO_1215 (O_1215,N_19963,N_19861);
xnor UO_1216 (O_1216,N_19718,N_19831);
and UO_1217 (O_1217,N_19835,N_19807);
and UO_1218 (O_1218,N_19977,N_19999);
nor UO_1219 (O_1219,N_19632,N_19924);
and UO_1220 (O_1220,N_19750,N_19855);
or UO_1221 (O_1221,N_19984,N_19694);
nand UO_1222 (O_1222,N_19968,N_19904);
nand UO_1223 (O_1223,N_19915,N_19845);
or UO_1224 (O_1224,N_19992,N_19802);
nand UO_1225 (O_1225,N_19893,N_19875);
nand UO_1226 (O_1226,N_19869,N_19703);
or UO_1227 (O_1227,N_19868,N_19975);
xor UO_1228 (O_1228,N_19669,N_19674);
nand UO_1229 (O_1229,N_19722,N_19786);
and UO_1230 (O_1230,N_19802,N_19972);
xnor UO_1231 (O_1231,N_19973,N_19671);
or UO_1232 (O_1232,N_19707,N_19729);
nor UO_1233 (O_1233,N_19827,N_19622);
nand UO_1234 (O_1234,N_19684,N_19849);
xor UO_1235 (O_1235,N_19749,N_19739);
and UO_1236 (O_1236,N_19609,N_19651);
nor UO_1237 (O_1237,N_19791,N_19697);
and UO_1238 (O_1238,N_19904,N_19989);
and UO_1239 (O_1239,N_19926,N_19856);
nand UO_1240 (O_1240,N_19754,N_19694);
xor UO_1241 (O_1241,N_19980,N_19742);
or UO_1242 (O_1242,N_19700,N_19679);
nor UO_1243 (O_1243,N_19662,N_19603);
nor UO_1244 (O_1244,N_19648,N_19688);
and UO_1245 (O_1245,N_19677,N_19916);
and UO_1246 (O_1246,N_19742,N_19683);
and UO_1247 (O_1247,N_19822,N_19752);
nand UO_1248 (O_1248,N_19945,N_19957);
xnor UO_1249 (O_1249,N_19984,N_19966);
xnor UO_1250 (O_1250,N_19648,N_19935);
or UO_1251 (O_1251,N_19823,N_19872);
xnor UO_1252 (O_1252,N_19920,N_19986);
nor UO_1253 (O_1253,N_19782,N_19641);
xnor UO_1254 (O_1254,N_19698,N_19804);
nor UO_1255 (O_1255,N_19929,N_19675);
xor UO_1256 (O_1256,N_19996,N_19924);
or UO_1257 (O_1257,N_19810,N_19841);
or UO_1258 (O_1258,N_19630,N_19636);
nor UO_1259 (O_1259,N_19947,N_19686);
nand UO_1260 (O_1260,N_19642,N_19939);
xor UO_1261 (O_1261,N_19686,N_19777);
nor UO_1262 (O_1262,N_19928,N_19796);
and UO_1263 (O_1263,N_19694,N_19757);
nand UO_1264 (O_1264,N_19695,N_19776);
and UO_1265 (O_1265,N_19954,N_19894);
nor UO_1266 (O_1266,N_19962,N_19622);
or UO_1267 (O_1267,N_19778,N_19819);
nor UO_1268 (O_1268,N_19637,N_19772);
and UO_1269 (O_1269,N_19736,N_19657);
nand UO_1270 (O_1270,N_19825,N_19726);
nor UO_1271 (O_1271,N_19771,N_19976);
or UO_1272 (O_1272,N_19720,N_19940);
nand UO_1273 (O_1273,N_19612,N_19877);
or UO_1274 (O_1274,N_19655,N_19657);
or UO_1275 (O_1275,N_19744,N_19635);
nand UO_1276 (O_1276,N_19871,N_19604);
or UO_1277 (O_1277,N_19696,N_19731);
nor UO_1278 (O_1278,N_19972,N_19746);
nor UO_1279 (O_1279,N_19837,N_19723);
or UO_1280 (O_1280,N_19685,N_19797);
xor UO_1281 (O_1281,N_19718,N_19678);
and UO_1282 (O_1282,N_19992,N_19772);
nor UO_1283 (O_1283,N_19634,N_19726);
nor UO_1284 (O_1284,N_19978,N_19922);
xnor UO_1285 (O_1285,N_19876,N_19928);
nand UO_1286 (O_1286,N_19643,N_19967);
or UO_1287 (O_1287,N_19988,N_19972);
nand UO_1288 (O_1288,N_19918,N_19981);
xor UO_1289 (O_1289,N_19866,N_19931);
xor UO_1290 (O_1290,N_19902,N_19621);
nor UO_1291 (O_1291,N_19709,N_19665);
nand UO_1292 (O_1292,N_19756,N_19794);
nor UO_1293 (O_1293,N_19663,N_19615);
nand UO_1294 (O_1294,N_19641,N_19710);
xnor UO_1295 (O_1295,N_19695,N_19928);
or UO_1296 (O_1296,N_19616,N_19615);
or UO_1297 (O_1297,N_19848,N_19841);
nor UO_1298 (O_1298,N_19613,N_19934);
and UO_1299 (O_1299,N_19674,N_19857);
nor UO_1300 (O_1300,N_19646,N_19916);
nor UO_1301 (O_1301,N_19974,N_19843);
xor UO_1302 (O_1302,N_19925,N_19948);
and UO_1303 (O_1303,N_19891,N_19698);
nor UO_1304 (O_1304,N_19829,N_19791);
nand UO_1305 (O_1305,N_19968,N_19963);
nand UO_1306 (O_1306,N_19951,N_19656);
or UO_1307 (O_1307,N_19706,N_19678);
nand UO_1308 (O_1308,N_19968,N_19693);
nand UO_1309 (O_1309,N_19889,N_19986);
xor UO_1310 (O_1310,N_19887,N_19644);
and UO_1311 (O_1311,N_19768,N_19641);
or UO_1312 (O_1312,N_19887,N_19783);
or UO_1313 (O_1313,N_19732,N_19860);
nand UO_1314 (O_1314,N_19966,N_19948);
xor UO_1315 (O_1315,N_19837,N_19737);
or UO_1316 (O_1316,N_19631,N_19722);
nand UO_1317 (O_1317,N_19626,N_19661);
and UO_1318 (O_1318,N_19880,N_19668);
xor UO_1319 (O_1319,N_19796,N_19973);
and UO_1320 (O_1320,N_19649,N_19759);
nand UO_1321 (O_1321,N_19988,N_19839);
nor UO_1322 (O_1322,N_19970,N_19879);
nand UO_1323 (O_1323,N_19638,N_19857);
nand UO_1324 (O_1324,N_19663,N_19636);
or UO_1325 (O_1325,N_19744,N_19837);
or UO_1326 (O_1326,N_19731,N_19902);
nor UO_1327 (O_1327,N_19642,N_19621);
nor UO_1328 (O_1328,N_19889,N_19732);
nand UO_1329 (O_1329,N_19711,N_19760);
and UO_1330 (O_1330,N_19794,N_19600);
or UO_1331 (O_1331,N_19865,N_19776);
nand UO_1332 (O_1332,N_19604,N_19783);
nand UO_1333 (O_1333,N_19912,N_19967);
and UO_1334 (O_1334,N_19746,N_19883);
nor UO_1335 (O_1335,N_19798,N_19749);
and UO_1336 (O_1336,N_19932,N_19738);
or UO_1337 (O_1337,N_19952,N_19898);
nor UO_1338 (O_1338,N_19757,N_19980);
and UO_1339 (O_1339,N_19768,N_19748);
nand UO_1340 (O_1340,N_19891,N_19710);
or UO_1341 (O_1341,N_19667,N_19719);
nor UO_1342 (O_1342,N_19841,N_19974);
nor UO_1343 (O_1343,N_19621,N_19734);
or UO_1344 (O_1344,N_19751,N_19621);
xnor UO_1345 (O_1345,N_19666,N_19956);
nand UO_1346 (O_1346,N_19973,N_19980);
or UO_1347 (O_1347,N_19979,N_19629);
or UO_1348 (O_1348,N_19887,N_19714);
xor UO_1349 (O_1349,N_19920,N_19728);
and UO_1350 (O_1350,N_19725,N_19882);
xnor UO_1351 (O_1351,N_19789,N_19795);
and UO_1352 (O_1352,N_19684,N_19672);
or UO_1353 (O_1353,N_19852,N_19965);
nand UO_1354 (O_1354,N_19838,N_19939);
nor UO_1355 (O_1355,N_19644,N_19698);
nand UO_1356 (O_1356,N_19983,N_19805);
nor UO_1357 (O_1357,N_19650,N_19662);
nand UO_1358 (O_1358,N_19723,N_19773);
or UO_1359 (O_1359,N_19705,N_19848);
and UO_1360 (O_1360,N_19677,N_19940);
nand UO_1361 (O_1361,N_19867,N_19937);
or UO_1362 (O_1362,N_19698,N_19942);
nor UO_1363 (O_1363,N_19769,N_19925);
or UO_1364 (O_1364,N_19942,N_19870);
xnor UO_1365 (O_1365,N_19638,N_19763);
nor UO_1366 (O_1366,N_19982,N_19809);
and UO_1367 (O_1367,N_19942,N_19700);
nand UO_1368 (O_1368,N_19714,N_19648);
nand UO_1369 (O_1369,N_19998,N_19602);
and UO_1370 (O_1370,N_19675,N_19729);
and UO_1371 (O_1371,N_19834,N_19613);
or UO_1372 (O_1372,N_19689,N_19868);
nor UO_1373 (O_1373,N_19786,N_19671);
or UO_1374 (O_1374,N_19665,N_19976);
and UO_1375 (O_1375,N_19701,N_19932);
and UO_1376 (O_1376,N_19880,N_19747);
nand UO_1377 (O_1377,N_19963,N_19948);
and UO_1378 (O_1378,N_19994,N_19854);
or UO_1379 (O_1379,N_19613,N_19782);
or UO_1380 (O_1380,N_19745,N_19738);
nand UO_1381 (O_1381,N_19806,N_19883);
nor UO_1382 (O_1382,N_19947,N_19851);
nand UO_1383 (O_1383,N_19806,N_19880);
xor UO_1384 (O_1384,N_19842,N_19970);
nor UO_1385 (O_1385,N_19661,N_19940);
nor UO_1386 (O_1386,N_19904,N_19776);
or UO_1387 (O_1387,N_19967,N_19782);
nand UO_1388 (O_1388,N_19908,N_19852);
xnor UO_1389 (O_1389,N_19979,N_19848);
xor UO_1390 (O_1390,N_19710,N_19671);
nand UO_1391 (O_1391,N_19958,N_19771);
nor UO_1392 (O_1392,N_19906,N_19956);
nand UO_1393 (O_1393,N_19812,N_19966);
and UO_1394 (O_1394,N_19682,N_19696);
and UO_1395 (O_1395,N_19903,N_19696);
nor UO_1396 (O_1396,N_19933,N_19900);
or UO_1397 (O_1397,N_19760,N_19804);
and UO_1398 (O_1398,N_19625,N_19971);
xor UO_1399 (O_1399,N_19825,N_19785);
and UO_1400 (O_1400,N_19789,N_19673);
and UO_1401 (O_1401,N_19816,N_19687);
xor UO_1402 (O_1402,N_19966,N_19615);
xor UO_1403 (O_1403,N_19660,N_19829);
nand UO_1404 (O_1404,N_19885,N_19810);
nor UO_1405 (O_1405,N_19846,N_19900);
or UO_1406 (O_1406,N_19930,N_19908);
nand UO_1407 (O_1407,N_19787,N_19775);
nor UO_1408 (O_1408,N_19633,N_19686);
nor UO_1409 (O_1409,N_19770,N_19732);
or UO_1410 (O_1410,N_19695,N_19691);
nor UO_1411 (O_1411,N_19613,N_19734);
nand UO_1412 (O_1412,N_19631,N_19996);
and UO_1413 (O_1413,N_19735,N_19628);
nor UO_1414 (O_1414,N_19970,N_19704);
xor UO_1415 (O_1415,N_19659,N_19783);
nor UO_1416 (O_1416,N_19888,N_19953);
nand UO_1417 (O_1417,N_19896,N_19640);
xor UO_1418 (O_1418,N_19770,N_19634);
nor UO_1419 (O_1419,N_19933,N_19828);
and UO_1420 (O_1420,N_19638,N_19660);
or UO_1421 (O_1421,N_19977,N_19840);
nand UO_1422 (O_1422,N_19763,N_19828);
nor UO_1423 (O_1423,N_19780,N_19643);
nor UO_1424 (O_1424,N_19657,N_19624);
or UO_1425 (O_1425,N_19767,N_19724);
nand UO_1426 (O_1426,N_19962,N_19857);
nand UO_1427 (O_1427,N_19982,N_19790);
or UO_1428 (O_1428,N_19799,N_19661);
and UO_1429 (O_1429,N_19809,N_19983);
nand UO_1430 (O_1430,N_19953,N_19738);
or UO_1431 (O_1431,N_19618,N_19874);
nor UO_1432 (O_1432,N_19916,N_19650);
or UO_1433 (O_1433,N_19650,N_19611);
xnor UO_1434 (O_1434,N_19717,N_19812);
or UO_1435 (O_1435,N_19783,N_19934);
or UO_1436 (O_1436,N_19742,N_19866);
and UO_1437 (O_1437,N_19867,N_19935);
or UO_1438 (O_1438,N_19695,N_19829);
nand UO_1439 (O_1439,N_19784,N_19798);
and UO_1440 (O_1440,N_19842,N_19964);
nor UO_1441 (O_1441,N_19715,N_19602);
nor UO_1442 (O_1442,N_19674,N_19986);
or UO_1443 (O_1443,N_19916,N_19614);
or UO_1444 (O_1444,N_19913,N_19752);
and UO_1445 (O_1445,N_19784,N_19903);
and UO_1446 (O_1446,N_19719,N_19828);
xnor UO_1447 (O_1447,N_19864,N_19707);
xnor UO_1448 (O_1448,N_19941,N_19762);
nor UO_1449 (O_1449,N_19717,N_19692);
and UO_1450 (O_1450,N_19867,N_19844);
nor UO_1451 (O_1451,N_19672,N_19709);
nor UO_1452 (O_1452,N_19976,N_19984);
and UO_1453 (O_1453,N_19630,N_19760);
and UO_1454 (O_1454,N_19721,N_19759);
nand UO_1455 (O_1455,N_19871,N_19779);
nor UO_1456 (O_1456,N_19648,N_19658);
nor UO_1457 (O_1457,N_19734,N_19997);
and UO_1458 (O_1458,N_19613,N_19841);
nor UO_1459 (O_1459,N_19745,N_19943);
and UO_1460 (O_1460,N_19928,N_19601);
nand UO_1461 (O_1461,N_19629,N_19666);
or UO_1462 (O_1462,N_19952,N_19964);
and UO_1463 (O_1463,N_19926,N_19602);
nor UO_1464 (O_1464,N_19867,N_19906);
or UO_1465 (O_1465,N_19728,N_19827);
nor UO_1466 (O_1466,N_19910,N_19778);
nor UO_1467 (O_1467,N_19601,N_19867);
or UO_1468 (O_1468,N_19795,N_19886);
or UO_1469 (O_1469,N_19711,N_19850);
nand UO_1470 (O_1470,N_19854,N_19992);
or UO_1471 (O_1471,N_19767,N_19706);
nor UO_1472 (O_1472,N_19632,N_19876);
nor UO_1473 (O_1473,N_19957,N_19969);
or UO_1474 (O_1474,N_19901,N_19681);
and UO_1475 (O_1475,N_19997,N_19873);
or UO_1476 (O_1476,N_19907,N_19713);
nor UO_1477 (O_1477,N_19617,N_19650);
and UO_1478 (O_1478,N_19609,N_19829);
nor UO_1479 (O_1479,N_19752,N_19647);
nor UO_1480 (O_1480,N_19927,N_19685);
xor UO_1481 (O_1481,N_19883,N_19875);
or UO_1482 (O_1482,N_19806,N_19915);
nor UO_1483 (O_1483,N_19646,N_19999);
and UO_1484 (O_1484,N_19991,N_19902);
and UO_1485 (O_1485,N_19926,N_19792);
or UO_1486 (O_1486,N_19887,N_19623);
xor UO_1487 (O_1487,N_19662,N_19920);
and UO_1488 (O_1488,N_19786,N_19825);
xnor UO_1489 (O_1489,N_19613,N_19614);
or UO_1490 (O_1490,N_19723,N_19656);
or UO_1491 (O_1491,N_19632,N_19882);
xor UO_1492 (O_1492,N_19842,N_19870);
or UO_1493 (O_1493,N_19952,N_19815);
nor UO_1494 (O_1494,N_19827,N_19696);
xor UO_1495 (O_1495,N_19607,N_19690);
nand UO_1496 (O_1496,N_19883,N_19838);
and UO_1497 (O_1497,N_19603,N_19755);
nor UO_1498 (O_1498,N_19792,N_19976);
nand UO_1499 (O_1499,N_19612,N_19804);
xnor UO_1500 (O_1500,N_19962,N_19671);
or UO_1501 (O_1501,N_19990,N_19916);
and UO_1502 (O_1502,N_19941,N_19700);
nand UO_1503 (O_1503,N_19922,N_19614);
and UO_1504 (O_1504,N_19911,N_19771);
xnor UO_1505 (O_1505,N_19697,N_19986);
or UO_1506 (O_1506,N_19809,N_19919);
nor UO_1507 (O_1507,N_19867,N_19618);
nor UO_1508 (O_1508,N_19898,N_19838);
or UO_1509 (O_1509,N_19726,N_19690);
nand UO_1510 (O_1510,N_19884,N_19801);
and UO_1511 (O_1511,N_19812,N_19746);
or UO_1512 (O_1512,N_19686,N_19663);
xnor UO_1513 (O_1513,N_19713,N_19882);
nor UO_1514 (O_1514,N_19871,N_19711);
nor UO_1515 (O_1515,N_19731,N_19750);
nor UO_1516 (O_1516,N_19847,N_19674);
nand UO_1517 (O_1517,N_19998,N_19646);
nor UO_1518 (O_1518,N_19792,N_19871);
or UO_1519 (O_1519,N_19785,N_19869);
nand UO_1520 (O_1520,N_19980,N_19785);
and UO_1521 (O_1521,N_19765,N_19630);
and UO_1522 (O_1522,N_19668,N_19982);
or UO_1523 (O_1523,N_19734,N_19777);
xnor UO_1524 (O_1524,N_19771,N_19895);
or UO_1525 (O_1525,N_19729,N_19846);
nand UO_1526 (O_1526,N_19852,N_19974);
or UO_1527 (O_1527,N_19955,N_19921);
nor UO_1528 (O_1528,N_19715,N_19764);
nand UO_1529 (O_1529,N_19636,N_19946);
xnor UO_1530 (O_1530,N_19704,N_19949);
and UO_1531 (O_1531,N_19852,N_19998);
or UO_1532 (O_1532,N_19729,N_19693);
and UO_1533 (O_1533,N_19723,N_19739);
nand UO_1534 (O_1534,N_19625,N_19947);
xor UO_1535 (O_1535,N_19716,N_19843);
nor UO_1536 (O_1536,N_19748,N_19756);
nand UO_1537 (O_1537,N_19994,N_19636);
nand UO_1538 (O_1538,N_19701,N_19989);
and UO_1539 (O_1539,N_19776,N_19977);
or UO_1540 (O_1540,N_19759,N_19724);
nor UO_1541 (O_1541,N_19606,N_19655);
nor UO_1542 (O_1542,N_19703,N_19698);
nor UO_1543 (O_1543,N_19823,N_19916);
nand UO_1544 (O_1544,N_19975,N_19962);
and UO_1545 (O_1545,N_19704,N_19658);
xnor UO_1546 (O_1546,N_19708,N_19866);
nor UO_1547 (O_1547,N_19818,N_19678);
nand UO_1548 (O_1548,N_19613,N_19883);
and UO_1549 (O_1549,N_19840,N_19721);
and UO_1550 (O_1550,N_19745,N_19633);
nor UO_1551 (O_1551,N_19881,N_19751);
nor UO_1552 (O_1552,N_19737,N_19876);
or UO_1553 (O_1553,N_19888,N_19983);
or UO_1554 (O_1554,N_19886,N_19623);
xnor UO_1555 (O_1555,N_19952,N_19659);
and UO_1556 (O_1556,N_19817,N_19977);
and UO_1557 (O_1557,N_19793,N_19925);
nand UO_1558 (O_1558,N_19934,N_19664);
and UO_1559 (O_1559,N_19629,N_19658);
nand UO_1560 (O_1560,N_19931,N_19636);
nor UO_1561 (O_1561,N_19761,N_19990);
and UO_1562 (O_1562,N_19956,N_19996);
or UO_1563 (O_1563,N_19797,N_19842);
xnor UO_1564 (O_1564,N_19857,N_19839);
nor UO_1565 (O_1565,N_19745,N_19879);
or UO_1566 (O_1566,N_19913,N_19696);
and UO_1567 (O_1567,N_19670,N_19674);
or UO_1568 (O_1568,N_19732,N_19749);
xor UO_1569 (O_1569,N_19894,N_19822);
or UO_1570 (O_1570,N_19964,N_19726);
nor UO_1571 (O_1571,N_19789,N_19837);
or UO_1572 (O_1572,N_19929,N_19723);
or UO_1573 (O_1573,N_19918,N_19613);
xnor UO_1574 (O_1574,N_19628,N_19994);
nor UO_1575 (O_1575,N_19728,N_19846);
nor UO_1576 (O_1576,N_19952,N_19721);
xor UO_1577 (O_1577,N_19942,N_19927);
xnor UO_1578 (O_1578,N_19689,N_19988);
nor UO_1579 (O_1579,N_19950,N_19718);
xor UO_1580 (O_1580,N_19835,N_19895);
and UO_1581 (O_1581,N_19945,N_19662);
nor UO_1582 (O_1582,N_19893,N_19986);
xnor UO_1583 (O_1583,N_19738,N_19638);
nor UO_1584 (O_1584,N_19723,N_19626);
nor UO_1585 (O_1585,N_19869,N_19941);
nor UO_1586 (O_1586,N_19822,N_19974);
nor UO_1587 (O_1587,N_19982,N_19997);
and UO_1588 (O_1588,N_19724,N_19749);
or UO_1589 (O_1589,N_19745,N_19973);
or UO_1590 (O_1590,N_19942,N_19791);
nand UO_1591 (O_1591,N_19797,N_19751);
nor UO_1592 (O_1592,N_19988,N_19906);
xor UO_1593 (O_1593,N_19664,N_19842);
nand UO_1594 (O_1594,N_19811,N_19659);
nand UO_1595 (O_1595,N_19617,N_19876);
nand UO_1596 (O_1596,N_19811,N_19961);
or UO_1597 (O_1597,N_19759,N_19600);
nor UO_1598 (O_1598,N_19728,N_19981);
xnor UO_1599 (O_1599,N_19684,N_19717);
nor UO_1600 (O_1600,N_19943,N_19939);
nand UO_1601 (O_1601,N_19652,N_19849);
or UO_1602 (O_1602,N_19606,N_19927);
xor UO_1603 (O_1603,N_19618,N_19666);
and UO_1604 (O_1604,N_19839,N_19917);
and UO_1605 (O_1605,N_19789,N_19814);
or UO_1606 (O_1606,N_19873,N_19964);
or UO_1607 (O_1607,N_19656,N_19857);
and UO_1608 (O_1608,N_19769,N_19727);
nor UO_1609 (O_1609,N_19824,N_19765);
xor UO_1610 (O_1610,N_19638,N_19780);
or UO_1611 (O_1611,N_19842,N_19656);
nor UO_1612 (O_1612,N_19840,N_19764);
xnor UO_1613 (O_1613,N_19875,N_19638);
and UO_1614 (O_1614,N_19626,N_19926);
nand UO_1615 (O_1615,N_19600,N_19943);
xor UO_1616 (O_1616,N_19731,N_19905);
nor UO_1617 (O_1617,N_19845,N_19746);
nand UO_1618 (O_1618,N_19859,N_19966);
and UO_1619 (O_1619,N_19941,N_19837);
nor UO_1620 (O_1620,N_19963,N_19833);
nand UO_1621 (O_1621,N_19718,N_19702);
xnor UO_1622 (O_1622,N_19668,N_19687);
and UO_1623 (O_1623,N_19943,N_19825);
nor UO_1624 (O_1624,N_19694,N_19862);
or UO_1625 (O_1625,N_19966,N_19988);
xnor UO_1626 (O_1626,N_19749,N_19990);
nand UO_1627 (O_1627,N_19898,N_19682);
nand UO_1628 (O_1628,N_19860,N_19655);
nand UO_1629 (O_1629,N_19608,N_19604);
and UO_1630 (O_1630,N_19869,N_19642);
or UO_1631 (O_1631,N_19672,N_19933);
nand UO_1632 (O_1632,N_19659,N_19736);
nor UO_1633 (O_1633,N_19944,N_19860);
xnor UO_1634 (O_1634,N_19774,N_19683);
nor UO_1635 (O_1635,N_19806,N_19817);
and UO_1636 (O_1636,N_19949,N_19823);
and UO_1637 (O_1637,N_19976,N_19952);
or UO_1638 (O_1638,N_19686,N_19856);
xor UO_1639 (O_1639,N_19970,N_19865);
xnor UO_1640 (O_1640,N_19836,N_19852);
nor UO_1641 (O_1641,N_19863,N_19932);
nor UO_1642 (O_1642,N_19840,N_19871);
nor UO_1643 (O_1643,N_19641,N_19986);
xnor UO_1644 (O_1644,N_19975,N_19624);
nand UO_1645 (O_1645,N_19847,N_19915);
or UO_1646 (O_1646,N_19761,N_19777);
xnor UO_1647 (O_1647,N_19875,N_19718);
and UO_1648 (O_1648,N_19696,N_19730);
xor UO_1649 (O_1649,N_19619,N_19928);
xnor UO_1650 (O_1650,N_19851,N_19669);
nand UO_1651 (O_1651,N_19713,N_19777);
xnor UO_1652 (O_1652,N_19843,N_19685);
nand UO_1653 (O_1653,N_19686,N_19735);
or UO_1654 (O_1654,N_19677,N_19828);
and UO_1655 (O_1655,N_19810,N_19850);
and UO_1656 (O_1656,N_19643,N_19928);
nand UO_1657 (O_1657,N_19617,N_19761);
nor UO_1658 (O_1658,N_19606,N_19766);
and UO_1659 (O_1659,N_19882,N_19685);
and UO_1660 (O_1660,N_19874,N_19829);
or UO_1661 (O_1661,N_19813,N_19995);
nor UO_1662 (O_1662,N_19905,N_19945);
and UO_1663 (O_1663,N_19885,N_19793);
or UO_1664 (O_1664,N_19757,N_19893);
and UO_1665 (O_1665,N_19990,N_19841);
nor UO_1666 (O_1666,N_19960,N_19959);
or UO_1667 (O_1667,N_19844,N_19826);
and UO_1668 (O_1668,N_19899,N_19851);
xor UO_1669 (O_1669,N_19946,N_19841);
nor UO_1670 (O_1670,N_19940,N_19788);
nor UO_1671 (O_1671,N_19711,N_19778);
nand UO_1672 (O_1672,N_19683,N_19695);
xor UO_1673 (O_1673,N_19750,N_19877);
and UO_1674 (O_1674,N_19924,N_19891);
nand UO_1675 (O_1675,N_19977,N_19768);
or UO_1676 (O_1676,N_19813,N_19970);
nor UO_1677 (O_1677,N_19778,N_19642);
nor UO_1678 (O_1678,N_19851,N_19800);
and UO_1679 (O_1679,N_19905,N_19817);
and UO_1680 (O_1680,N_19679,N_19709);
xnor UO_1681 (O_1681,N_19812,N_19628);
nor UO_1682 (O_1682,N_19955,N_19818);
and UO_1683 (O_1683,N_19904,N_19939);
nor UO_1684 (O_1684,N_19663,N_19605);
nand UO_1685 (O_1685,N_19626,N_19863);
nor UO_1686 (O_1686,N_19859,N_19971);
nand UO_1687 (O_1687,N_19887,N_19830);
nand UO_1688 (O_1688,N_19927,N_19978);
or UO_1689 (O_1689,N_19902,N_19661);
nand UO_1690 (O_1690,N_19933,N_19848);
and UO_1691 (O_1691,N_19905,N_19721);
and UO_1692 (O_1692,N_19806,N_19651);
nor UO_1693 (O_1693,N_19901,N_19645);
or UO_1694 (O_1694,N_19601,N_19600);
or UO_1695 (O_1695,N_19881,N_19879);
xnor UO_1696 (O_1696,N_19739,N_19923);
nand UO_1697 (O_1697,N_19861,N_19729);
xor UO_1698 (O_1698,N_19896,N_19863);
or UO_1699 (O_1699,N_19909,N_19851);
and UO_1700 (O_1700,N_19867,N_19625);
xnor UO_1701 (O_1701,N_19829,N_19901);
and UO_1702 (O_1702,N_19735,N_19955);
xnor UO_1703 (O_1703,N_19601,N_19796);
xor UO_1704 (O_1704,N_19765,N_19866);
xor UO_1705 (O_1705,N_19690,N_19950);
or UO_1706 (O_1706,N_19677,N_19618);
nor UO_1707 (O_1707,N_19939,N_19738);
nor UO_1708 (O_1708,N_19653,N_19804);
and UO_1709 (O_1709,N_19757,N_19604);
nor UO_1710 (O_1710,N_19763,N_19780);
nand UO_1711 (O_1711,N_19922,N_19707);
nor UO_1712 (O_1712,N_19893,N_19970);
xnor UO_1713 (O_1713,N_19789,N_19719);
nand UO_1714 (O_1714,N_19902,N_19924);
xor UO_1715 (O_1715,N_19666,N_19620);
or UO_1716 (O_1716,N_19835,N_19908);
xnor UO_1717 (O_1717,N_19841,N_19994);
and UO_1718 (O_1718,N_19640,N_19769);
nor UO_1719 (O_1719,N_19686,N_19766);
xnor UO_1720 (O_1720,N_19827,N_19618);
nor UO_1721 (O_1721,N_19872,N_19687);
and UO_1722 (O_1722,N_19986,N_19895);
or UO_1723 (O_1723,N_19993,N_19633);
xor UO_1724 (O_1724,N_19965,N_19897);
xor UO_1725 (O_1725,N_19926,N_19801);
nand UO_1726 (O_1726,N_19750,N_19968);
nor UO_1727 (O_1727,N_19925,N_19759);
nor UO_1728 (O_1728,N_19889,N_19681);
nand UO_1729 (O_1729,N_19837,N_19640);
and UO_1730 (O_1730,N_19623,N_19965);
and UO_1731 (O_1731,N_19824,N_19686);
or UO_1732 (O_1732,N_19657,N_19740);
xor UO_1733 (O_1733,N_19891,N_19986);
xnor UO_1734 (O_1734,N_19943,N_19616);
or UO_1735 (O_1735,N_19674,N_19929);
xnor UO_1736 (O_1736,N_19854,N_19951);
xor UO_1737 (O_1737,N_19662,N_19816);
and UO_1738 (O_1738,N_19958,N_19991);
nand UO_1739 (O_1739,N_19803,N_19697);
xor UO_1740 (O_1740,N_19698,N_19692);
xor UO_1741 (O_1741,N_19615,N_19629);
or UO_1742 (O_1742,N_19740,N_19829);
xnor UO_1743 (O_1743,N_19869,N_19759);
nand UO_1744 (O_1744,N_19794,N_19648);
nand UO_1745 (O_1745,N_19729,N_19802);
nor UO_1746 (O_1746,N_19912,N_19910);
nand UO_1747 (O_1747,N_19934,N_19943);
and UO_1748 (O_1748,N_19737,N_19867);
xnor UO_1749 (O_1749,N_19937,N_19991);
nor UO_1750 (O_1750,N_19675,N_19898);
xor UO_1751 (O_1751,N_19735,N_19731);
xor UO_1752 (O_1752,N_19743,N_19883);
and UO_1753 (O_1753,N_19759,N_19952);
xnor UO_1754 (O_1754,N_19925,N_19637);
nor UO_1755 (O_1755,N_19897,N_19948);
nand UO_1756 (O_1756,N_19979,N_19648);
nor UO_1757 (O_1757,N_19899,N_19973);
nor UO_1758 (O_1758,N_19789,N_19653);
nor UO_1759 (O_1759,N_19907,N_19952);
xnor UO_1760 (O_1760,N_19863,N_19779);
and UO_1761 (O_1761,N_19730,N_19925);
or UO_1762 (O_1762,N_19900,N_19961);
or UO_1763 (O_1763,N_19954,N_19783);
xor UO_1764 (O_1764,N_19774,N_19971);
and UO_1765 (O_1765,N_19771,N_19691);
nor UO_1766 (O_1766,N_19970,N_19734);
nand UO_1767 (O_1767,N_19746,N_19955);
xor UO_1768 (O_1768,N_19711,N_19696);
nand UO_1769 (O_1769,N_19899,N_19664);
nor UO_1770 (O_1770,N_19771,N_19748);
and UO_1771 (O_1771,N_19613,N_19850);
and UO_1772 (O_1772,N_19774,N_19905);
or UO_1773 (O_1773,N_19704,N_19836);
and UO_1774 (O_1774,N_19992,N_19880);
nand UO_1775 (O_1775,N_19861,N_19965);
nor UO_1776 (O_1776,N_19729,N_19602);
and UO_1777 (O_1777,N_19681,N_19847);
nor UO_1778 (O_1778,N_19775,N_19849);
xor UO_1779 (O_1779,N_19631,N_19903);
and UO_1780 (O_1780,N_19718,N_19795);
or UO_1781 (O_1781,N_19608,N_19636);
and UO_1782 (O_1782,N_19805,N_19946);
nand UO_1783 (O_1783,N_19892,N_19952);
and UO_1784 (O_1784,N_19813,N_19825);
nand UO_1785 (O_1785,N_19628,N_19786);
nor UO_1786 (O_1786,N_19898,N_19924);
xor UO_1787 (O_1787,N_19680,N_19981);
nand UO_1788 (O_1788,N_19850,N_19748);
and UO_1789 (O_1789,N_19981,N_19707);
or UO_1790 (O_1790,N_19638,N_19729);
xor UO_1791 (O_1791,N_19944,N_19667);
nor UO_1792 (O_1792,N_19789,N_19992);
or UO_1793 (O_1793,N_19857,N_19852);
or UO_1794 (O_1794,N_19785,N_19911);
xnor UO_1795 (O_1795,N_19779,N_19852);
nand UO_1796 (O_1796,N_19913,N_19835);
nor UO_1797 (O_1797,N_19832,N_19877);
xnor UO_1798 (O_1798,N_19701,N_19604);
nor UO_1799 (O_1799,N_19624,N_19943);
and UO_1800 (O_1800,N_19622,N_19824);
nand UO_1801 (O_1801,N_19938,N_19873);
or UO_1802 (O_1802,N_19972,N_19957);
and UO_1803 (O_1803,N_19966,N_19703);
xnor UO_1804 (O_1804,N_19623,N_19626);
or UO_1805 (O_1805,N_19773,N_19652);
nor UO_1806 (O_1806,N_19681,N_19981);
nor UO_1807 (O_1807,N_19936,N_19746);
nor UO_1808 (O_1808,N_19619,N_19887);
nor UO_1809 (O_1809,N_19873,N_19987);
and UO_1810 (O_1810,N_19803,N_19918);
and UO_1811 (O_1811,N_19624,N_19737);
nor UO_1812 (O_1812,N_19822,N_19930);
nand UO_1813 (O_1813,N_19746,N_19865);
and UO_1814 (O_1814,N_19701,N_19695);
nor UO_1815 (O_1815,N_19979,N_19819);
or UO_1816 (O_1816,N_19762,N_19933);
nor UO_1817 (O_1817,N_19819,N_19739);
or UO_1818 (O_1818,N_19633,N_19909);
xnor UO_1819 (O_1819,N_19912,N_19659);
nand UO_1820 (O_1820,N_19766,N_19678);
nand UO_1821 (O_1821,N_19782,N_19777);
nor UO_1822 (O_1822,N_19776,N_19795);
and UO_1823 (O_1823,N_19914,N_19892);
or UO_1824 (O_1824,N_19985,N_19823);
and UO_1825 (O_1825,N_19723,N_19681);
xnor UO_1826 (O_1826,N_19715,N_19725);
and UO_1827 (O_1827,N_19617,N_19651);
and UO_1828 (O_1828,N_19988,N_19734);
xor UO_1829 (O_1829,N_19993,N_19906);
or UO_1830 (O_1830,N_19884,N_19885);
xnor UO_1831 (O_1831,N_19790,N_19741);
nand UO_1832 (O_1832,N_19972,N_19761);
nor UO_1833 (O_1833,N_19636,N_19917);
nor UO_1834 (O_1834,N_19931,N_19782);
and UO_1835 (O_1835,N_19766,N_19786);
xnor UO_1836 (O_1836,N_19778,N_19637);
nand UO_1837 (O_1837,N_19630,N_19958);
and UO_1838 (O_1838,N_19941,N_19644);
nand UO_1839 (O_1839,N_19955,N_19665);
and UO_1840 (O_1840,N_19893,N_19704);
nand UO_1841 (O_1841,N_19924,N_19773);
nor UO_1842 (O_1842,N_19803,N_19880);
or UO_1843 (O_1843,N_19757,N_19626);
or UO_1844 (O_1844,N_19767,N_19761);
or UO_1845 (O_1845,N_19942,N_19797);
and UO_1846 (O_1846,N_19680,N_19704);
nor UO_1847 (O_1847,N_19833,N_19952);
and UO_1848 (O_1848,N_19925,N_19797);
nor UO_1849 (O_1849,N_19785,N_19752);
nand UO_1850 (O_1850,N_19923,N_19915);
xor UO_1851 (O_1851,N_19852,N_19657);
nand UO_1852 (O_1852,N_19913,N_19726);
or UO_1853 (O_1853,N_19790,N_19814);
xnor UO_1854 (O_1854,N_19825,N_19602);
nand UO_1855 (O_1855,N_19828,N_19693);
and UO_1856 (O_1856,N_19837,N_19818);
nor UO_1857 (O_1857,N_19979,N_19934);
nand UO_1858 (O_1858,N_19926,N_19788);
nand UO_1859 (O_1859,N_19717,N_19851);
nand UO_1860 (O_1860,N_19775,N_19826);
nand UO_1861 (O_1861,N_19646,N_19901);
xor UO_1862 (O_1862,N_19907,N_19730);
nand UO_1863 (O_1863,N_19698,N_19728);
and UO_1864 (O_1864,N_19681,N_19610);
or UO_1865 (O_1865,N_19944,N_19938);
nor UO_1866 (O_1866,N_19603,N_19673);
or UO_1867 (O_1867,N_19611,N_19621);
nor UO_1868 (O_1868,N_19839,N_19690);
and UO_1869 (O_1869,N_19841,N_19779);
nor UO_1870 (O_1870,N_19980,N_19658);
or UO_1871 (O_1871,N_19680,N_19890);
and UO_1872 (O_1872,N_19718,N_19842);
or UO_1873 (O_1873,N_19782,N_19963);
nand UO_1874 (O_1874,N_19740,N_19778);
nor UO_1875 (O_1875,N_19749,N_19673);
or UO_1876 (O_1876,N_19873,N_19747);
or UO_1877 (O_1877,N_19832,N_19787);
nor UO_1878 (O_1878,N_19668,N_19633);
and UO_1879 (O_1879,N_19620,N_19986);
nor UO_1880 (O_1880,N_19879,N_19946);
and UO_1881 (O_1881,N_19607,N_19694);
nor UO_1882 (O_1882,N_19978,N_19941);
nand UO_1883 (O_1883,N_19740,N_19946);
nor UO_1884 (O_1884,N_19985,N_19924);
or UO_1885 (O_1885,N_19974,N_19842);
nor UO_1886 (O_1886,N_19856,N_19937);
nor UO_1887 (O_1887,N_19615,N_19624);
nor UO_1888 (O_1888,N_19894,N_19932);
and UO_1889 (O_1889,N_19806,N_19945);
xnor UO_1890 (O_1890,N_19824,N_19848);
xnor UO_1891 (O_1891,N_19738,N_19641);
and UO_1892 (O_1892,N_19746,N_19940);
or UO_1893 (O_1893,N_19860,N_19926);
and UO_1894 (O_1894,N_19623,N_19798);
or UO_1895 (O_1895,N_19741,N_19699);
and UO_1896 (O_1896,N_19860,N_19618);
and UO_1897 (O_1897,N_19990,N_19778);
xor UO_1898 (O_1898,N_19667,N_19768);
nor UO_1899 (O_1899,N_19908,N_19752);
nor UO_1900 (O_1900,N_19762,N_19925);
xnor UO_1901 (O_1901,N_19668,N_19616);
xnor UO_1902 (O_1902,N_19977,N_19635);
xnor UO_1903 (O_1903,N_19906,N_19798);
nor UO_1904 (O_1904,N_19607,N_19792);
or UO_1905 (O_1905,N_19638,N_19607);
or UO_1906 (O_1906,N_19638,N_19849);
nor UO_1907 (O_1907,N_19734,N_19888);
xnor UO_1908 (O_1908,N_19663,N_19950);
or UO_1909 (O_1909,N_19764,N_19623);
nor UO_1910 (O_1910,N_19656,N_19934);
nand UO_1911 (O_1911,N_19720,N_19936);
or UO_1912 (O_1912,N_19874,N_19762);
xor UO_1913 (O_1913,N_19946,N_19632);
xnor UO_1914 (O_1914,N_19812,N_19686);
nand UO_1915 (O_1915,N_19829,N_19931);
nor UO_1916 (O_1916,N_19648,N_19827);
nor UO_1917 (O_1917,N_19633,N_19712);
nor UO_1918 (O_1918,N_19954,N_19844);
or UO_1919 (O_1919,N_19770,N_19752);
nand UO_1920 (O_1920,N_19881,N_19861);
or UO_1921 (O_1921,N_19717,N_19758);
and UO_1922 (O_1922,N_19832,N_19912);
and UO_1923 (O_1923,N_19810,N_19700);
and UO_1924 (O_1924,N_19950,N_19778);
nand UO_1925 (O_1925,N_19851,N_19694);
nand UO_1926 (O_1926,N_19803,N_19957);
or UO_1927 (O_1927,N_19819,N_19808);
and UO_1928 (O_1928,N_19634,N_19769);
or UO_1929 (O_1929,N_19945,N_19619);
and UO_1930 (O_1930,N_19641,N_19867);
nand UO_1931 (O_1931,N_19814,N_19963);
nor UO_1932 (O_1932,N_19727,N_19793);
or UO_1933 (O_1933,N_19887,N_19711);
or UO_1934 (O_1934,N_19849,N_19930);
nand UO_1935 (O_1935,N_19849,N_19862);
and UO_1936 (O_1936,N_19713,N_19876);
and UO_1937 (O_1937,N_19824,N_19620);
and UO_1938 (O_1938,N_19775,N_19908);
nor UO_1939 (O_1939,N_19856,N_19762);
and UO_1940 (O_1940,N_19830,N_19698);
xnor UO_1941 (O_1941,N_19603,N_19604);
xor UO_1942 (O_1942,N_19672,N_19856);
nor UO_1943 (O_1943,N_19744,N_19642);
xnor UO_1944 (O_1944,N_19935,N_19836);
and UO_1945 (O_1945,N_19892,N_19733);
or UO_1946 (O_1946,N_19760,N_19930);
xnor UO_1947 (O_1947,N_19805,N_19935);
xnor UO_1948 (O_1948,N_19943,N_19783);
nand UO_1949 (O_1949,N_19980,N_19737);
nor UO_1950 (O_1950,N_19609,N_19934);
xnor UO_1951 (O_1951,N_19813,N_19846);
nor UO_1952 (O_1952,N_19960,N_19905);
nor UO_1953 (O_1953,N_19666,N_19955);
and UO_1954 (O_1954,N_19632,N_19828);
or UO_1955 (O_1955,N_19773,N_19847);
nand UO_1956 (O_1956,N_19817,N_19871);
nand UO_1957 (O_1957,N_19809,N_19922);
nand UO_1958 (O_1958,N_19777,N_19711);
nand UO_1959 (O_1959,N_19643,N_19669);
nand UO_1960 (O_1960,N_19692,N_19899);
or UO_1961 (O_1961,N_19915,N_19602);
or UO_1962 (O_1962,N_19620,N_19854);
nand UO_1963 (O_1963,N_19630,N_19827);
or UO_1964 (O_1964,N_19928,N_19748);
nand UO_1965 (O_1965,N_19953,N_19704);
nand UO_1966 (O_1966,N_19933,N_19608);
nand UO_1967 (O_1967,N_19624,N_19876);
or UO_1968 (O_1968,N_19769,N_19613);
xor UO_1969 (O_1969,N_19860,N_19875);
nand UO_1970 (O_1970,N_19884,N_19781);
and UO_1971 (O_1971,N_19767,N_19637);
nor UO_1972 (O_1972,N_19725,N_19671);
nand UO_1973 (O_1973,N_19873,N_19641);
nor UO_1974 (O_1974,N_19934,N_19685);
nand UO_1975 (O_1975,N_19664,N_19662);
nor UO_1976 (O_1976,N_19793,N_19743);
nor UO_1977 (O_1977,N_19752,N_19944);
nand UO_1978 (O_1978,N_19787,N_19951);
nor UO_1979 (O_1979,N_19766,N_19644);
and UO_1980 (O_1980,N_19712,N_19806);
nor UO_1981 (O_1981,N_19878,N_19678);
nor UO_1982 (O_1982,N_19908,N_19727);
and UO_1983 (O_1983,N_19945,N_19729);
nor UO_1984 (O_1984,N_19762,N_19735);
xnor UO_1985 (O_1985,N_19657,N_19776);
xnor UO_1986 (O_1986,N_19997,N_19804);
or UO_1987 (O_1987,N_19833,N_19944);
and UO_1988 (O_1988,N_19747,N_19739);
or UO_1989 (O_1989,N_19951,N_19883);
nand UO_1990 (O_1990,N_19614,N_19955);
nand UO_1991 (O_1991,N_19885,N_19777);
or UO_1992 (O_1992,N_19699,N_19975);
and UO_1993 (O_1993,N_19605,N_19818);
or UO_1994 (O_1994,N_19691,N_19650);
or UO_1995 (O_1995,N_19762,N_19613);
nor UO_1996 (O_1996,N_19984,N_19989);
nand UO_1997 (O_1997,N_19944,N_19755);
nand UO_1998 (O_1998,N_19856,N_19881);
nand UO_1999 (O_1999,N_19746,N_19669);
nor UO_2000 (O_2000,N_19620,N_19849);
nand UO_2001 (O_2001,N_19793,N_19970);
or UO_2002 (O_2002,N_19653,N_19686);
nor UO_2003 (O_2003,N_19710,N_19968);
nand UO_2004 (O_2004,N_19823,N_19977);
nor UO_2005 (O_2005,N_19634,N_19702);
nor UO_2006 (O_2006,N_19989,N_19813);
or UO_2007 (O_2007,N_19751,N_19827);
nand UO_2008 (O_2008,N_19707,N_19764);
xnor UO_2009 (O_2009,N_19889,N_19963);
or UO_2010 (O_2010,N_19627,N_19987);
nor UO_2011 (O_2011,N_19800,N_19881);
nand UO_2012 (O_2012,N_19754,N_19872);
and UO_2013 (O_2013,N_19660,N_19765);
or UO_2014 (O_2014,N_19968,N_19858);
xor UO_2015 (O_2015,N_19692,N_19777);
and UO_2016 (O_2016,N_19977,N_19949);
and UO_2017 (O_2017,N_19612,N_19632);
nand UO_2018 (O_2018,N_19724,N_19707);
nor UO_2019 (O_2019,N_19951,N_19613);
xor UO_2020 (O_2020,N_19941,N_19808);
and UO_2021 (O_2021,N_19619,N_19971);
nand UO_2022 (O_2022,N_19694,N_19663);
nand UO_2023 (O_2023,N_19928,N_19815);
nor UO_2024 (O_2024,N_19666,N_19923);
nor UO_2025 (O_2025,N_19714,N_19854);
and UO_2026 (O_2026,N_19642,N_19785);
and UO_2027 (O_2027,N_19823,N_19937);
or UO_2028 (O_2028,N_19897,N_19635);
nor UO_2029 (O_2029,N_19863,N_19995);
xnor UO_2030 (O_2030,N_19661,N_19769);
or UO_2031 (O_2031,N_19601,N_19614);
or UO_2032 (O_2032,N_19956,N_19703);
nand UO_2033 (O_2033,N_19861,N_19610);
xnor UO_2034 (O_2034,N_19861,N_19797);
nand UO_2035 (O_2035,N_19627,N_19810);
and UO_2036 (O_2036,N_19651,N_19804);
nor UO_2037 (O_2037,N_19675,N_19988);
or UO_2038 (O_2038,N_19720,N_19909);
nand UO_2039 (O_2039,N_19604,N_19849);
and UO_2040 (O_2040,N_19659,N_19746);
and UO_2041 (O_2041,N_19815,N_19855);
nor UO_2042 (O_2042,N_19986,N_19882);
and UO_2043 (O_2043,N_19801,N_19750);
or UO_2044 (O_2044,N_19840,N_19766);
nand UO_2045 (O_2045,N_19831,N_19627);
nor UO_2046 (O_2046,N_19799,N_19986);
xor UO_2047 (O_2047,N_19649,N_19924);
or UO_2048 (O_2048,N_19834,N_19818);
or UO_2049 (O_2049,N_19913,N_19766);
nand UO_2050 (O_2050,N_19608,N_19855);
nor UO_2051 (O_2051,N_19977,N_19852);
and UO_2052 (O_2052,N_19895,N_19736);
and UO_2053 (O_2053,N_19626,N_19791);
nor UO_2054 (O_2054,N_19918,N_19899);
and UO_2055 (O_2055,N_19874,N_19852);
nor UO_2056 (O_2056,N_19782,N_19672);
and UO_2057 (O_2057,N_19961,N_19692);
nor UO_2058 (O_2058,N_19882,N_19633);
nor UO_2059 (O_2059,N_19618,N_19635);
and UO_2060 (O_2060,N_19718,N_19746);
xnor UO_2061 (O_2061,N_19801,N_19689);
or UO_2062 (O_2062,N_19746,N_19899);
or UO_2063 (O_2063,N_19720,N_19783);
or UO_2064 (O_2064,N_19754,N_19922);
nor UO_2065 (O_2065,N_19700,N_19980);
or UO_2066 (O_2066,N_19814,N_19636);
or UO_2067 (O_2067,N_19891,N_19958);
or UO_2068 (O_2068,N_19864,N_19891);
nand UO_2069 (O_2069,N_19907,N_19688);
or UO_2070 (O_2070,N_19954,N_19825);
or UO_2071 (O_2071,N_19908,N_19974);
nand UO_2072 (O_2072,N_19907,N_19850);
and UO_2073 (O_2073,N_19847,N_19781);
xor UO_2074 (O_2074,N_19958,N_19801);
or UO_2075 (O_2075,N_19933,N_19820);
nand UO_2076 (O_2076,N_19841,N_19707);
xor UO_2077 (O_2077,N_19977,N_19800);
xnor UO_2078 (O_2078,N_19646,N_19653);
nor UO_2079 (O_2079,N_19906,N_19888);
nand UO_2080 (O_2080,N_19802,N_19753);
or UO_2081 (O_2081,N_19856,N_19633);
nand UO_2082 (O_2082,N_19788,N_19790);
or UO_2083 (O_2083,N_19872,N_19778);
or UO_2084 (O_2084,N_19882,N_19608);
and UO_2085 (O_2085,N_19813,N_19819);
and UO_2086 (O_2086,N_19828,N_19903);
or UO_2087 (O_2087,N_19841,N_19888);
xor UO_2088 (O_2088,N_19637,N_19818);
xnor UO_2089 (O_2089,N_19693,N_19801);
xor UO_2090 (O_2090,N_19969,N_19851);
nor UO_2091 (O_2091,N_19751,N_19880);
xnor UO_2092 (O_2092,N_19636,N_19738);
nand UO_2093 (O_2093,N_19965,N_19605);
nor UO_2094 (O_2094,N_19709,N_19677);
nor UO_2095 (O_2095,N_19638,N_19805);
or UO_2096 (O_2096,N_19683,N_19897);
or UO_2097 (O_2097,N_19850,N_19826);
or UO_2098 (O_2098,N_19985,N_19842);
nor UO_2099 (O_2099,N_19817,N_19788);
and UO_2100 (O_2100,N_19680,N_19606);
nor UO_2101 (O_2101,N_19694,N_19760);
or UO_2102 (O_2102,N_19996,N_19617);
and UO_2103 (O_2103,N_19924,N_19758);
xor UO_2104 (O_2104,N_19956,N_19902);
nand UO_2105 (O_2105,N_19806,N_19619);
and UO_2106 (O_2106,N_19840,N_19842);
nand UO_2107 (O_2107,N_19741,N_19755);
and UO_2108 (O_2108,N_19883,N_19926);
nand UO_2109 (O_2109,N_19890,N_19716);
or UO_2110 (O_2110,N_19738,N_19631);
nor UO_2111 (O_2111,N_19625,N_19997);
nor UO_2112 (O_2112,N_19680,N_19881);
and UO_2113 (O_2113,N_19848,N_19726);
nor UO_2114 (O_2114,N_19999,N_19799);
nand UO_2115 (O_2115,N_19963,N_19942);
xor UO_2116 (O_2116,N_19612,N_19783);
nor UO_2117 (O_2117,N_19987,N_19622);
and UO_2118 (O_2118,N_19986,N_19991);
nand UO_2119 (O_2119,N_19949,N_19992);
xnor UO_2120 (O_2120,N_19915,N_19799);
and UO_2121 (O_2121,N_19898,N_19758);
xor UO_2122 (O_2122,N_19655,N_19684);
nand UO_2123 (O_2123,N_19845,N_19902);
nor UO_2124 (O_2124,N_19951,N_19871);
nor UO_2125 (O_2125,N_19910,N_19710);
nand UO_2126 (O_2126,N_19608,N_19702);
nor UO_2127 (O_2127,N_19999,N_19843);
and UO_2128 (O_2128,N_19617,N_19866);
and UO_2129 (O_2129,N_19758,N_19669);
and UO_2130 (O_2130,N_19793,N_19651);
and UO_2131 (O_2131,N_19609,N_19671);
nand UO_2132 (O_2132,N_19689,N_19752);
and UO_2133 (O_2133,N_19680,N_19829);
nand UO_2134 (O_2134,N_19604,N_19760);
nand UO_2135 (O_2135,N_19680,N_19810);
and UO_2136 (O_2136,N_19758,N_19958);
nor UO_2137 (O_2137,N_19917,N_19879);
nor UO_2138 (O_2138,N_19827,N_19886);
or UO_2139 (O_2139,N_19624,N_19835);
or UO_2140 (O_2140,N_19787,N_19984);
and UO_2141 (O_2141,N_19879,N_19808);
nor UO_2142 (O_2142,N_19682,N_19697);
xor UO_2143 (O_2143,N_19827,N_19643);
or UO_2144 (O_2144,N_19652,N_19639);
nor UO_2145 (O_2145,N_19978,N_19721);
or UO_2146 (O_2146,N_19659,N_19777);
xnor UO_2147 (O_2147,N_19654,N_19667);
and UO_2148 (O_2148,N_19772,N_19874);
nand UO_2149 (O_2149,N_19744,N_19792);
nor UO_2150 (O_2150,N_19883,N_19954);
nand UO_2151 (O_2151,N_19708,N_19650);
nand UO_2152 (O_2152,N_19983,N_19964);
and UO_2153 (O_2153,N_19619,N_19665);
nand UO_2154 (O_2154,N_19805,N_19993);
or UO_2155 (O_2155,N_19833,N_19964);
and UO_2156 (O_2156,N_19758,N_19763);
nand UO_2157 (O_2157,N_19918,N_19759);
and UO_2158 (O_2158,N_19767,N_19711);
nand UO_2159 (O_2159,N_19872,N_19906);
nand UO_2160 (O_2160,N_19683,N_19812);
and UO_2161 (O_2161,N_19665,N_19792);
nor UO_2162 (O_2162,N_19840,N_19837);
nand UO_2163 (O_2163,N_19903,N_19930);
and UO_2164 (O_2164,N_19602,N_19677);
xnor UO_2165 (O_2165,N_19930,N_19821);
xnor UO_2166 (O_2166,N_19706,N_19655);
and UO_2167 (O_2167,N_19703,N_19848);
and UO_2168 (O_2168,N_19962,N_19602);
and UO_2169 (O_2169,N_19789,N_19664);
nor UO_2170 (O_2170,N_19804,N_19602);
and UO_2171 (O_2171,N_19946,N_19612);
nor UO_2172 (O_2172,N_19773,N_19981);
or UO_2173 (O_2173,N_19812,N_19840);
and UO_2174 (O_2174,N_19647,N_19884);
nor UO_2175 (O_2175,N_19947,N_19637);
nand UO_2176 (O_2176,N_19958,N_19671);
nand UO_2177 (O_2177,N_19905,N_19684);
nand UO_2178 (O_2178,N_19606,N_19709);
and UO_2179 (O_2179,N_19685,N_19765);
nor UO_2180 (O_2180,N_19951,N_19671);
nor UO_2181 (O_2181,N_19749,N_19846);
nor UO_2182 (O_2182,N_19983,N_19912);
or UO_2183 (O_2183,N_19697,N_19853);
and UO_2184 (O_2184,N_19729,N_19918);
nand UO_2185 (O_2185,N_19788,N_19638);
nand UO_2186 (O_2186,N_19999,N_19797);
nor UO_2187 (O_2187,N_19895,N_19823);
nor UO_2188 (O_2188,N_19642,N_19923);
xnor UO_2189 (O_2189,N_19730,N_19630);
nor UO_2190 (O_2190,N_19616,N_19975);
and UO_2191 (O_2191,N_19707,N_19999);
nor UO_2192 (O_2192,N_19767,N_19787);
and UO_2193 (O_2193,N_19883,N_19851);
or UO_2194 (O_2194,N_19992,N_19748);
xor UO_2195 (O_2195,N_19660,N_19623);
and UO_2196 (O_2196,N_19617,N_19730);
or UO_2197 (O_2197,N_19835,N_19615);
xnor UO_2198 (O_2198,N_19743,N_19979);
and UO_2199 (O_2199,N_19627,N_19739);
nand UO_2200 (O_2200,N_19793,N_19677);
nand UO_2201 (O_2201,N_19721,N_19767);
nor UO_2202 (O_2202,N_19827,N_19950);
nand UO_2203 (O_2203,N_19870,N_19700);
and UO_2204 (O_2204,N_19723,N_19934);
xnor UO_2205 (O_2205,N_19973,N_19859);
nor UO_2206 (O_2206,N_19836,N_19927);
nand UO_2207 (O_2207,N_19851,N_19636);
and UO_2208 (O_2208,N_19935,N_19633);
xnor UO_2209 (O_2209,N_19791,N_19624);
or UO_2210 (O_2210,N_19796,N_19629);
and UO_2211 (O_2211,N_19870,N_19993);
and UO_2212 (O_2212,N_19716,N_19799);
nand UO_2213 (O_2213,N_19759,N_19881);
nand UO_2214 (O_2214,N_19744,N_19886);
xor UO_2215 (O_2215,N_19806,N_19932);
nor UO_2216 (O_2216,N_19632,N_19729);
nand UO_2217 (O_2217,N_19811,N_19859);
and UO_2218 (O_2218,N_19963,N_19789);
xor UO_2219 (O_2219,N_19946,N_19976);
nor UO_2220 (O_2220,N_19731,N_19818);
or UO_2221 (O_2221,N_19620,N_19795);
or UO_2222 (O_2222,N_19977,N_19944);
nor UO_2223 (O_2223,N_19889,N_19972);
nor UO_2224 (O_2224,N_19881,N_19963);
and UO_2225 (O_2225,N_19658,N_19928);
nor UO_2226 (O_2226,N_19707,N_19614);
or UO_2227 (O_2227,N_19858,N_19775);
nand UO_2228 (O_2228,N_19901,N_19859);
nand UO_2229 (O_2229,N_19822,N_19785);
xnor UO_2230 (O_2230,N_19899,N_19926);
or UO_2231 (O_2231,N_19720,N_19612);
nand UO_2232 (O_2232,N_19832,N_19719);
and UO_2233 (O_2233,N_19943,N_19654);
and UO_2234 (O_2234,N_19804,N_19665);
xor UO_2235 (O_2235,N_19990,N_19812);
and UO_2236 (O_2236,N_19817,N_19861);
nor UO_2237 (O_2237,N_19713,N_19870);
xnor UO_2238 (O_2238,N_19959,N_19663);
nor UO_2239 (O_2239,N_19683,N_19906);
nor UO_2240 (O_2240,N_19625,N_19973);
xor UO_2241 (O_2241,N_19611,N_19929);
nand UO_2242 (O_2242,N_19618,N_19602);
nor UO_2243 (O_2243,N_19839,N_19699);
nor UO_2244 (O_2244,N_19630,N_19862);
xor UO_2245 (O_2245,N_19982,N_19976);
nor UO_2246 (O_2246,N_19986,N_19997);
and UO_2247 (O_2247,N_19866,N_19660);
nand UO_2248 (O_2248,N_19808,N_19873);
or UO_2249 (O_2249,N_19620,N_19773);
nand UO_2250 (O_2250,N_19968,N_19745);
and UO_2251 (O_2251,N_19630,N_19988);
nor UO_2252 (O_2252,N_19827,N_19978);
nand UO_2253 (O_2253,N_19799,N_19865);
nand UO_2254 (O_2254,N_19670,N_19959);
or UO_2255 (O_2255,N_19625,N_19900);
and UO_2256 (O_2256,N_19942,N_19674);
nand UO_2257 (O_2257,N_19767,N_19685);
nand UO_2258 (O_2258,N_19672,N_19926);
and UO_2259 (O_2259,N_19924,N_19960);
or UO_2260 (O_2260,N_19652,N_19798);
xor UO_2261 (O_2261,N_19767,N_19804);
and UO_2262 (O_2262,N_19826,N_19711);
and UO_2263 (O_2263,N_19726,N_19881);
or UO_2264 (O_2264,N_19637,N_19978);
xnor UO_2265 (O_2265,N_19896,N_19748);
nor UO_2266 (O_2266,N_19895,N_19838);
or UO_2267 (O_2267,N_19794,N_19687);
xor UO_2268 (O_2268,N_19749,N_19776);
nor UO_2269 (O_2269,N_19989,N_19916);
xor UO_2270 (O_2270,N_19607,N_19618);
nand UO_2271 (O_2271,N_19675,N_19691);
nor UO_2272 (O_2272,N_19765,N_19886);
or UO_2273 (O_2273,N_19887,N_19974);
xor UO_2274 (O_2274,N_19810,N_19910);
nor UO_2275 (O_2275,N_19652,N_19988);
and UO_2276 (O_2276,N_19950,N_19818);
nand UO_2277 (O_2277,N_19994,N_19913);
nor UO_2278 (O_2278,N_19613,N_19649);
nand UO_2279 (O_2279,N_19721,N_19705);
xor UO_2280 (O_2280,N_19851,N_19971);
xor UO_2281 (O_2281,N_19866,N_19988);
nor UO_2282 (O_2282,N_19655,N_19965);
nor UO_2283 (O_2283,N_19891,N_19919);
xor UO_2284 (O_2284,N_19937,N_19948);
xor UO_2285 (O_2285,N_19913,N_19784);
xor UO_2286 (O_2286,N_19892,N_19955);
xor UO_2287 (O_2287,N_19902,N_19890);
xnor UO_2288 (O_2288,N_19760,N_19657);
or UO_2289 (O_2289,N_19618,N_19922);
or UO_2290 (O_2290,N_19723,N_19648);
and UO_2291 (O_2291,N_19816,N_19786);
and UO_2292 (O_2292,N_19894,N_19937);
nand UO_2293 (O_2293,N_19652,N_19826);
or UO_2294 (O_2294,N_19958,N_19802);
nand UO_2295 (O_2295,N_19640,N_19988);
nand UO_2296 (O_2296,N_19981,N_19878);
xor UO_2297 (O_2297,N_19977,N_19644);
and UO_2298 (O_2298,N_19846,N_19675);
and UO_2299 (O_2299,N_19865,N_19755);
or UO_2300 (O_2300,N_19753,N_19823);
nand UO_2301 (O_2301,N_19980,N_19943);
nor UO_2302 (O_2302,N_19964,N_19815);
nor UO_2303 (O_2303,N_19873,N_19735);
or UO_2304 (O_2304,N_19650,N_19868);
or UO_2305 (O_2305,N_19927,N_19910);
and UO_2306 (O_2306,N_19870,N_19794);
nand UO_2307 (O_2307,N_19806,N_19741);
nand UO_2308 (O_2308,N_19837,N_19714);
nor UO_2309 (O_2309,N_19658,N_19735);
and UO_2310 (O_2310,N_19902,N_19803);
nor UO_2311 (O_2311,N_19893,N_19913);
or UO_2312 (O_2312,N_19821,N_19753);
and UO_2313 (O_2313,N_19651,N_19977);
nor UO_2314 (O_2314,N_19631,N_19893);
nand UO_2315 (O_2315,N_19633,N_19973);
or UO_2316 (O_2316,N_19849,N_19881);
xor UO_2317 (O_2317,N_19891,N_19645);
nand UO_2318 (O_2318,N_19967,N_19985);
and UO_2319 (O_2319,N_19655,N_19909);
nor UO_2320 (O_2320,N_19965,N_19919);
nand UO_2321 (O_2321,N_19810,N_19669);
xor UO_2322 (O_2322,N_19754,N_19947);
xor UO_2323 (O_2323,N_19702,N_19897);
and UO_2324 (O_2324,N_19713,N_19686);
nor UO_2325 (O_2325,N_19686,N_19946);
and UO_2326 (O_2326,N_19742,N_19716);
or UO_2327 (O_2327,N_19973,N_19866);
xnor UO_2328 (O_2328,N_19920,N_19863);
and UO_2329 (O_2329,N_19632,N_19721);
nand UO_2330 (O_2330,N_19893,N_19801);
and UO_2331 (O_2331,N_19676,N_19944);
xor UO_2332 (O_2332,N_19946,N_19831);
nand UO_2333 (O_2333,N_19898,N_19997);
xor UO_2334 (O_2334,N_19760,N_19949);
or UO_2335 (O_2335,N_19665,N_19746);
nand UO_2336 (O_2336,N_19987,N_19977);
nand UO_2337 (O_2337,N_19916,N_19944);
nand UO_2338 (O_2338,N_19899,N_19694);
and UO_2339 (O_2339,N_19709,N_19814);
or UO_2340 (O_2340,N_19877,N_19674);
and UO_2341 (O_2341,N_19839,N_19649);
xor UO_2342 (O_2342,N_19824,N_19910);
or UO_2343 (O_2343,N_19874,N_19608);
and UO_2344 (O_2344,N_19753,N_19873);
nand UO_2345 (O_2345,N_19962,N_19973);
nor UO_2346 (O_2346,N_19910,N_19838);
xor UO_2347 (O_2347,N_19645,N_19984);
or UO_2348 (O_2348,N_19931,N_19922);
or UO_2349 (O_2349,N_19916,N_19752);
or UO_2350 (O_2350,N_19932,N_19925);
nor UO_2351 (O_2351,N_19995,N_19666);
nor UO_2352 (O_2352,N_19749,N_19876);
nor UO_2353 (O_2353,N_19836,N_19614);
nor UO_2354 (O_2354,N_19910,N_19609);
and UO_2355 (O_2355,N_19984,N_19677);
nand UO_2356 (O_2356,N_19637,N_19906);
xor UO_2357 (O_2357,N_19963,N_19887);
and UO_2358 (O_2358,N_19951,N_19905);
xnor UO_2359 (O_2359,N_19886,N_19818);
nor UO_2360 (O_2360,N_19670,N_19830);
and UO_2361 (O_2361,N_19841,N_19877);
or UO_2362 (O_2362,N_19708,N_19641);
and UO_2363 (O_2363,N_19776,N_19952);
and UO_2364 (O_2364,N_19660,N_19607);
xor UO_2365 (O_2365,N_19843,N_19921);
nor UO_2366 (O_2366,N_19628,N_19659);
xor UO_2367 (O_2367,N_19606,N_19789);
or UO_2368 (O_2368,N_19810,N_19772);
and UO_2369 (O_2369,N_19698,N_19952);
nand UO_2370 (O_2370,N_19882,N_19629);
xor UO_2371 (O_2371,N_19842,N_19788);
and UO_2372 (O_2372,N_19800,N_19915);
and UO_2373 (O_2373,N_19605,N_19664);
nor UO_2374 (O_2374,N_19621,N_19898);
xnor UO_2375 (O_2375,N_19646,N_19765);
and UO_2376 (O_2376,N_19621,N_19720);
nor UO_2377 (O_2377,N_19631,N_19739);
and UO_2378 (O_2378,N_19722,N_19943);
and UO_2379 (O_2379,N_19624,N_19916);
xor UO_2380 (O_2380,N_19881,N_19985);
xor UO_2381 (O_2381,N_19739,N_19635);
nand UO_2382 (O_2382,N_19956,N_19960);
nand UO_2383 (O_2383,N_19738,N_19752);
xnor UO_2384 (O_2384,N_19720,N_19802);
xor UO_2385 (O_2385,N_19730,N_19869);
and UO_2386 (O_2386,N_19750,N_19723);
nor UO_2387 (O_2387,N_19779,N_19968);
xnor UO_2388 (O_2388,N_19887,N_19617);
nand UO_2389 (O_2389,N_19932,N_19904);
nand UO_2390 (O_2390,N_19843,N_19808);
nand UO_2391 (O_2391,N_19943,N_19998);
nor UO_2392 (O_2392,N_19750,N_19897);
or UO_2393 (O_2393,N_19885,N_19642);
xnor UO_2394 (O_2394,N_19951,N_19670);
and UO_2395 (O_2395,N_19803,N_19778);
nand UO_2396 (O_2396,N_19996,N_19788);
xnor UO_2397 (O_2397,N_19628,N_19779);
nor UO_2398 (O_2398,N_19721,N_19662);
or UO_2399 (O_2399,N_19835,N_19625);
xnor UO_2400 (O_2400,N_19802,N_19953);
nand UO_2401 (O_2401,N_19829,N_19932);
nand UO_2402 (O_2402,N_19660,N_19816);
nor UO_2403 (O_2403,N_19923,N_19979);
and UO_2404 (O_2404,N_19963,N_19815);
nor UO_2405 (O_2405,N_19731,N_19875);
nor UO_2406 (O_2406,N_19980,N_19902);
xor UO_2407 (O_2407,N_19903,N_19833);
and UO_2408 (O_2408,N_19896,N_19627);
nand UO_2409 (O_2409,N_19837,N_19937);
xnor UO_2410 (O_2410,N_19776,N_19624);
or UO_2411 (O_2411,N_19894,N_19874);
or UO_2412 (O_2412,N_19760,N_19744);
nand UO_2413 (O_2413,N_19704,N_19969);
or UO_2414 (O_2414,N_19979,N_19844);
and UO_2415 (O_2415,N_19891,N_19870);
xor UO_2416 (O_2416,N_19605,N_19929);
nand UO_2417 (O_2417,N_19623,N_19611);
nor UO_2418 (O_2418,N_19982,N_19841);
and UO_2419 (O_2419,N_19860,N_19798);
and UO_2420 (O_2420,N_19631,N_19815);
nor UO_2421 (O_2421,N_19659,N_19848);
nand UO_2422 (O_2422,N_19692,N_19911);
nor UO_2423 (O_2423,N_19898,N_19766);
nor UO_2424 (O_2424,N_19801,N_19938);
and UO_2425 (O_2425,N_19678,N_19879);
nor UO_2426 (O_2426,N_19910,N_19870);
and UO_2427 (O_2427,N_19628,N_19866);
nand UO_2428 (O_2428,N_19830,N_19783);
and UO_2429 (O_2429,N_19898,N_19820);
xor UO_2430 (O_2430,N_19936,N_19991);
nand UO_2431 (O_2431,N_19619,N_19788);
xor UO_2432 (O_2432,N_19976,N_19920);
and UO_2433 (O_2433,N_19812,N_19834);
nand UO_2434 (O_2434,N_19665,N_19736);
nand UO_2435 (O_2435,N_19729,N_19917);
and UO_2436 (O_2436,N_19910,N_19894);
and UO_2437 (O_2437,N_19996,N_19931);
nor UO_2438 (O_2438,N_19722,N_19763);
nand UO_2439 (O_2439,N_19836,N_19695);
nand UO_2440 (O_2440,N_19907,N_19988);
nor UO_2441 (O_2441,N_19606,N_19746);
and UO_2442 (O_2442,N_19608,N_19979);
xnor UO_2443 (O_2443,N_19814,N_19721);
nor UO_2444 (O_2444,N_19996,N_19911);
and UO_2445 (O_2445,N_19867,N_19930);
xor UO_2446 (O_2446,N_19793,N_19942);
and UO_2447 (O_2447,N_19803,N_19925);
nor UO_2448 (O_2448,N_19649,N_19787);
xor UO_2449 (O_2449,N_19968,N_19607);
xnor UO_2450 (O_2450,N_19746,N_19794);
nand UO_2451 (O_2451,N_19711,N_19725);
and UO_2452 (O_2452,N_19934,N_19883);
nand UO_2453 (O_2453,N_19715,N_19604);
or UO_2454 (O_2454,N_19865,N_19761);
and UO_2455 (O_2455,N_19703,N_19726);
or UO_2456 (O_2456,N_19764,N_19702);
and UO_2457 (O_2457,N_19759,N_19941);
xor UO_2458 (O_2458,N_19631,N_19618);
nor UO_2459 (O_2459,N_19803,N_19718);
and UO_2460 (O_2460,N_19691,N_19916);
nor UO_2461 (O_2461,N_19928,N_19671);
and UO_2462 (O_2462,N_19646,N_19857);
xnor UO_2463 (O_2463,N_19848,N_19851);
xnor UO_2464 (O_2464,N_19666,N_19637);
or UO_2465 (O_2465,N_19879,N_19769);
or UO_2466 (O_2466,N_19619,N_19990);
xnor UO_2467 (O_2467,N_19790,N_19858);
xnor UO_2468 (O_2468,N_19958,N_19887);
nor UO_2469 (O_2469,N_19959,N_19681);
nand UO_2470 (O_2470,N_19709,N_19965);
nor UO_2471 (O_2471,N_19902,N_19769);
nor UO_2472 (O_2472,N_19889,N_19840);
xor UO_2473 (O_2473,N_19749,N_19703);
nor UO_2474 (O_2474,N_19950,N_19780);
or UO_2475 (O_2475,N_19871,N_19879);
xor UO_2476 (O_2476,N_19951,N_19826);
or UO_2477 (O_2477,N_19969,N_19967);
nor UO_2478 (O_2478,N_19750,N_19770);
xor UO_2479 (O_2479,N_19809,N_19658);
nor UO_2480 (O_2480,N_19852,N_19624);
and UO_2481 (O_2481,N_19821,N_19694);
nor UO_2482 (O_2482,N_19889,N_19821);
xor UO_2483 (O_2483,N_19801,N_19891);
or UO_2484 (O_2484,N_19941,N_19647);
nand UO_2485 (O_2485,N_19848,N_19863);
xnor UO_2486 (O_2486,N_19893,N_19968);
and UO_2487 (O_2487,N_19751,N_19910);
nand UO_2488 (O_2488,N_19758,N_19609);
xor UO_2489 (O_2489,N_19898,N_19964);
nand UO_2490 (O_2490,N_19732,N_19796);
nor UO_2491 (O_2491,N_19680,N_19634);
nor UO_2492 (O_2492,N_19685,N_19802);
or UO_2493 (O_2493,N_19706,N_19938);
nor UO_2494 (O_2494,N_19991,N_19695);
xnor UO_2495 (O_2495,N_19778,N_19971);
nor UO_2496 (O_2496,N_19751,N_19838);
xnor UO_2497 (O_2497,N_19603,N_19898);
xnor UO_2498 (O_2498,N_19995,N_19763);
or UO_2499 (O_2499,N_19750,N_19952);
endmodule