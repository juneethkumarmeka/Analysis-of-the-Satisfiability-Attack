module basic_2500_25000_3000_8_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_1083,In_560);
nand U1 (N_1,In_849,In_1949);
xnor U2 (N_2,In_2411,In_2014);
nor U3 (N_3,In_304,In_639);
nor U4 (N_4,In_2025,In_1796);
xnor U5 (N_5,In_1917,In_767);
and U6 (N_6,In_1702,In_884);
nand U7 (N_7,In_2365,In_585);
or U8 (N_8,In_563,In_1946);
or U9 (N_9,In_1303,In_1831);
nand U10 (N_10,In_2312,In_1575);
nor U11 (N_11,In_728,In_1270);
and U12 (N_12,In_1935,In_1271);
or U13 (N_13,In_256,In_2325);
or U14 (N_14,In_1669,In_1834);
nor U15 (N_15,In_996,In_743);
and U16 (N_16,In_647,In_2206);
and U17 (N_17,In_1724,In_1485);
or U18 (N_18,In_1297,In_257);
or U19 (N_19,In_1244,In_1247);
nor U20 (N_20,In_2301,In_1838);
nand U21 (N_21,In_1887,In_1585);
xnor U22 (N_22,In_58,In_1554);
nor U23 (N_23,In_537,In_139);
or U24 (N_24,In_1673,In_581);
and U25 (N_25,In_548,In_1489);
and U26 (N_26,In_510,In_2335);
and U27 (N_27,In_1505,In_681);
nor U28 (N_28,In_662,In_673);
or U29 (N_29,In_1202,In_117);
or U30 (N_30,In_1191,In_1320);
nor U31 (N_31,In_221,In_1392);
nand U32 (N_32,In_1009,In_684);
or U33 (N_33,In_2475,In_2017);
or U34 (N_34,In_1389,In_1963);
or U35 (N_35,In_1626,In_1900);
nor U36 (N_36,In_1678,In_1890);
and U37 (N_37,In_817,In_1049);
xor U38 (N_38,In_392,In_176);
nand U39 (N_39,In_710,In_1893);
nand U40 (N_40,In_2306,In_1472);
or U41 (N_41,In_164,In_80);
xor U42 (N_42,In_920,In_306);
or U43 (N_43,In_1291,In_580);
nand U44 (N_44,In_2094,In_1707);
and U45 (N_45,In_1265,In_2121);
nand U46 (N_46,In_282,In_1363);
nor U47 (N_47,In_2370,In_2103);
nor U48 (N_48,In_1823,In_215);
or U49 (N_49,In_1637,In_2087);
nor U50 (N_50,In_2456,In_289);
xnor U51 (N_51,In_940,In_1751);
and U52 (N_52,In_790,In_2490);
nor U53 (N_53,In_2059,In_1753);
or U54 (N_54,In_1734,In_1667);
nor U55 (N_55,In_1569,In_1118);
and U56 (N_56,In_1361,In_1953);
nand U57 (N_57,In_1690,In_1179);
or U58 (N_58,In_2351,In_2040);
or U59 (N_59,In_520,In_2406);
nor U60 (N_60,In_183,In_49);
or U61 (N_61,In_2491,In_1916);
nor U62 (N_62,In_52,In_1155);
xnor U63 (N_63,In_1616,In_1051);
nor U64 (N_64,In_345,In_1222);
nor U65 (N_65,In_909,In_1475);
nand U66 (N_66,In_532,In_424);
nand U67 (N_67,In_1706,In_1653);
nand U68 (N_68,In_124,In_1962);
nor U69 (N_69,In_1108,In_1292);
nor U70 (N_70,In_629,In_2086);
nor U71 (N_71,In_1205,In_2063);
nor U72 (N_72,In_848,In_2056);
or U73 (N_73,In_2319,In_177);
and U74 (N_74,In_1967,In_1038);
or U75 (N_75,In_2262,In_154);
nor U76 (N_76,In_396,In_1728);
and U77 (N_77,In_1506,In_989);
nor U78 (N_78,In_951,In_357);
and U79 (N_79,In_957,In_1522);
nor U80 (N_80,In_1033,In_2323);
and U81 (N_81,In_2116,In_811);
and U82 (N_82,In_1134,In_1801);
nand U83 (N_83,In_212,In_336);
nor U84 (N_84,In_2449,In_889);
and U85 (N_85,In_825,In_543);
or U86 (N_86,In_1130,In_1727);
nor U87 (N_87,In_1842,In_1725);
nand U88 (N_88,In_490,In_934);
or U89 (N_89,In_1857,In_2190);
and U90 (N_90,In_1476,In_1880);
nand U91 (N_91,In_1206,In_1456);
xor U92 (N_92,In_171,In_2037);
xor U93 (N_93,In_2023,In_1666);
and U94 (N_94,In_1220,In_1581);
nand U95 (N_95,In_1611,In_1825);
nand U96 (N_96,In_2254,In_1198);
nand U97 (N_97,In_261,In_1470);
nor U98 (N_98,In_1371,In_668);
and U99 (N_99,In_343,In_1789);
nor U100 (N_100,In_1419,In_970);
or U101 (N_101,In_919,In_732);
or U102 (N_102,In_2144,In_819);
nand U103 (N_103,In_202,In_2194);
or U104 (N_104,In_92,In_635);
or U105 (N_105,In_739,In_2229);
nand U106 (N_106,In_44,In_2071);
or U107 (N_107,In_2459,In_1888);
xor U108 (N_108,In_2452,In_1113);
nor U109 (N_109,In_2293,In_1210);
or U110 (N_110,In_2230,In_2280);
nand U111 (N_111,In_795,In_584);
nor U112 (N_112,In_1047,In_1922);
or U113 (N_113,In_1605,In_1040);
nand U114 (N_114,In_809,In_1336);
or U115 (N_115,In_249,In_2150);
nand U116 (N_116,In_1741,In_1462);
xnor U117 (N_117,In_738,In_1993);
or U118 (N_118,In_1995,In_1004);
or U119 (N_119,In_2467,In_199);
or U120 (N_120,In_897,In_1037);
nand U121 (N_121,In_218,In_1186);
or U122 (N_122,In_279,In_1024);
or U123 (N_123,In_1345,In_245);
nand U124 (N_124,In_1212,In_29);
nor U125 (N_125,In_858,In_313);
nand U126 (N_126,In_1433,In_677);
or U127 (N_127,In_979,In_1633);
or U128 (N_128,In_954,In_1593);
nor U129 (N_129,In_2118,In_1532);
nand U130 (N_130,In_2385,In_1832);
nor U131 (N_131,In_1194,In_496);
nand U132 (N_132,In_1393,In_1928);
xor U133 (N_133,In_655,In_488);
nor U134 (N_134,In_975,In_481);
and U135 (N_135,In_450,In_337);
nand U136 (N_136,In_415,In_1164);
and U137 (N_137,In_1290,In_658);
nor U138 (N_138,In_562,In_2033);
nand U139 (N_139,In_615,In_1580);
nand U140 (N_140,In_1570,In_700);
nand U141 (N_141,In_1641,In_1800);
and U142 (N_142,In_2122,In_2314);
or U143 (N_143,In_59,In_526);
and U144 (N_144,In_1481,In_485);
or U145 (N_145,In_851,In_2376);
nor U146 (N_146,In_54,In_2353);
and U147 (N_147,In_796,In_38);
or U148 (N_148,In_2439,In_2266);
and U149 (N_149,In_427,In_2251);
xor U150 (N_150,In_1793,In_570);
or U151 (N_151,In_1597,In_822);
and U152 (N_152,In_947,In_77);
xnor U153 (N_153,In_404,In_149);
or U154 (N_154,In_1338,In_731);
and U155 (N_155,In_948,In_187);
nor U156 (N_156,In_1237,In_255);
xnor U157 (N_157,In_1714,In_987);
or U158 (N_158,In_805,In_1994);
xor U159 (N_159,In_1471,In_32);
nor U160 (N_160,In_2123,In_39);
or U161 (N_161,In_2067,In_1460);
or U162 (N_162,In_778,In_1968);
and U163 (N_163,In_1548,In_1883);
or U164 (N_164,In_2447,In_96);
nor U165 (N_165,In_482,In_2480);
and U166 (N_166,In_228,In_2349);
and U167 (N_167,In_985,In_1116);
or U168 (N_168,In_239,In_763);
xor U169 (N_169,In_899,In_327);
or U170 (N_170,In_2455,In_1982);
xnor U171 (N_171,In_1816,In_373);
or U172 (N_172,In_1552,In_911);
or U173 (N_173,In_56,In_2303);
and U174 (N_174,In_564,In_1703);
nand U175 (N_175,In_1933,In_2494);
nor U176 (N_176,In_33,In_921);
nand U177 (N_177,In_235,In_1936);
xor U178 (N_178,In_425,In_25);
nor U179 (N_179,In_1156,In_1814);
nand U180 (N_180,In_1971,In_2361);
and U181 (N_181,In_358,In_1892);
or U182 (N_182,In_2112,In_2205);
nor U183 (N_183,In_271,In_1467);
xnor U184 (N_184,In_1781,In_650);
and U185 (N_185,In_412,In_2287);
nor U186 (N_186,In_968,In_2263);
nand U187 (N_187,In_544,In_572);
nand U188 (N_188,In_1366,In_259);
nand U189 (N_189,In_785,In_1160);
or U190 (N_190,In_2394,In_1414);
or U191 (N_191,In_1868,In_1687);
nor U192 (N_192,In_836,In_2126);
nand U193 (N_193,In_2000,In_950);
xnor U194 (N_194,In_589,In_445);
and U195 (N_195,In_1642,In_2080);
nor U196 (N_196,In_2364,In_1573);
and U197 (N_197,In_123,In_144);
nand U198 (N_198,In_1073,In_1434);
nor U199 (N_199,In_733,In_620);
and U200 (N_200,In_2155,In_2345);
nand U201 (N_201,In_361,In_1520);
and U202 (N_202,In_1269,In_1177);
and U203 (N_203,In_1097,In_1306);
nand U204 (N_204,In_16,In_439);
and U205 (N_205,In_1263,In_293);
nand U206 (N_206,In_258,In_764);
xor U207 (N_207,In_2259,In_2318);
and U208 (N_208,In_1420,In_1693);
and U209 (N_209,In_19,In_857);
nor U210 (N_210,In_76,In_319);
xnor U211 (N_211,In_147,In_2214);
or U212 (N_212,In_2195,In_1343);
nor U213 (N_213,In_2288,In_1466);
nor U214 (N_214,In_2138,In_1030);
or U215 (N_215,In_15,In_1899);
and U216 (N_216,In_1443,In_850);
nor U217 (N_217,In_596,In_2409);
or U218 (N_218,In_833,In_156);
or U219 (N_219,In_1509,In_1511);
or U220 (N_220,In_573,In_2337);
and U221 (N_221,In_1864,In_974);
and U222 (N_222,In_1283,In_777);
or U223 (N_223,In_1952,In_971);
and U224 (N_224,In_1856,In_555);
nand U225 (N_225,In_1382,In_941);
nand U226 (N_226,In_112,In_414);
or U227 (N_227,In_2240,In_2030);
nor U228 (N_228,In_2149,In_2437);
and U229 (N_229,In_372,In_2381);
nor U230 (N_230,In_341,In_2342);
or U231 (N_231,In_1977,In_2196);
nor U232 (N_232,In_384,In_1068);
nor U233 (N_233,In_515,In_1188);
nor U234 (N_234,In_1135,In_2410);
and U235 (N_235,In_1440,In_1874);
nor U236 (N_236,In_2108,In_1930);
nand U237 (N_237,In_627,In_748);
nand U238 (N_238,In_806,In_522);
and U239 (N_239,In_945,In_2078);
nand U240 (N_240,In_839,In_2493);
and U241 (N_241,In_533,In_191);
xnor U242 (N_242,In_2111,In_1256);
nand U243 (N_243,In_2168,In_1299);
or U244 (N_244,In_108,In_1154);
or U245 (N_245,In_2284,In_682);
or U246 (N_246,In_538,In_346);
and U247 (N_247,In_686,In_633);
or U248 (N_248,In_351,In_1512);
and U249 (N_249,In_2137,In_1293);
and U250 (N_250,In_2373,In_442);
nand U251 (N_251,In_1077,In_1426);
nor U252 (N_252,In_408,In_1048);
xor U253 (N_253,In_2298,In_1317);
xor U254 (N_254,In_1430,In_625);
and U255 (N_255,In_1418,In_1975);
nand U256 (N_256,In_550,In_1891);
nor U257 (N_257,In_2484,In_248);
xor U258 (N_258,In_1733,In_617);
nor U259 (N_259,In_2226,In_2401);
nor U260 (N_260,In_2243,In_541);
nand U261 (N_261,In_1468,In_172);
nand U262 (N_262,In_1984,In_1139);
xor U263 (N_263,In_2244,In_469);
and U264 (N_264,In_2273,In_877);
and U265 (N_265,In_669,In_1799);
xor U266 (N_266,In_2400,In_251);
nand U267 (N_267,In_1412,In_547);
and U268 (N_268,In_2065,In_509);
or U269 (N_269,In_1101,In_1736);
or U270 (N_270,In_2089,In_1078);
and U271 (N_271,In_493,In_1233);
and U272 (N_272,In_2344,In_1207);
or U273 (N_273,In_1007,In_666);
or U274 (N_274,In_896,In_1192);
nand U275 (N_275,In_582,In_2486);
nand U276 (N_276,In_2479,In_826);
nor U277 (N_277,In_71,In_2258);
nand U278 (N_278,In_1855,In_861);
nand U279 (N_279,In_1094,In_2020);
or U280 (N_280,In_1529,In_1251);
nor U281 (N_281,In_269,In_2236);
xnor U282 (N_282,In_745,In_73);
nor U283 (N_283,In_207,In_1127);
or U284 (N_284,In_1375,In_1045);
nor U285 (N_285,In_1332,In_1881);
xor U286 (N_286,In_1016,In_1172);
nand U287 (N_287,In_2180,In_2470);
or U288 (N_288,In_579,In_479);
and U289 (N_289,In_905,In_2022);
nand U290 (N_290,In_1395,In_267);
nor U291 (N_291,In_2327,In_2350);
nand U292 (N_292,In_231,In_2153);
nand U293 (N_293,In_1232,In_1308);
or U294 (N_294,In_13,In_1408);
nor U295 (N_295,In_881,In_1587);
nor U296 (N_296,In_605,In_967);
nor U297 (N_297,In_1711,In_693);
nand U298 (N_298,In_1621,In_998);
nand U299 (N_299,In_1992,In_1589);
or U300 (N_300,In_1015,In_1833);
nor U301 (N_301,In_477,In_1630);
and U302 (N_302,In_2378,In_136);
and U303 (N_303,In_1301,In_339);
or U304 (N_304,In_1316,In_2464);
nor U305 (N_305,In_1309,In_2179);
or U306 (N_306,In_638,In_2292);
nand U307 (N_307,In_283,In_460);
or U308 (N_308,In_2395,In_1131);
nand U309 (N_309,In_914,In_298);
or U310 (N_310,In_2264,In_497);
and U311 (N_311,In_632,In_2203);
and U312 (N_312,In_1786,In_1594);
nand U313 (N_313,In_1406,In_1093);
nor U314 (N_314,In_1720,In_1954);
and U315 (N_315,In_350,In_137);
and U316 (N_316,In_518,In_2139);
nand U317 (N_317,In_2483,In_1404);
nand U318 (N_318,In_2471,In_1488);
or U319 (N_319,In_290,In_1439);
xor U320 (N_320,In_505,In_1879);
xor U321 (N_321,In_990,In_2165);
nand U322 (N_322,In_1791,In_1431);
nand U323 (N_323,In_935,In_1662);
or U324 (N_324,In_1717,In_872);
or U325 (N_325,In_976,In_208);
nor U326 (N_326,In_276,In_1624);
xor U327 (N_327,In_2274,In_774);
nand U328 (N_328,In_1973,In_1780);
and U329 (N_329,In_1726,In_2296);
and U330 (N_330,In_1835,In_2261);
and U331 (N_331,In_1173,In_723);
nand U332 (N_332,In_2221,In_1377);
nand U333 (N_333,In_2047,In_1959);
or U334 (N_334,In_2387,In_800);
and U335 (N_335,In_753,In_265);
and U336 (N_336,In_1010,In_2291);
or U337 (N_337,In_2382,In_2418);
nand U338 (N_338,In_318,In_1153);
and U339 (N_339,In_1671,In_2430);
nand U340 (N_340,In_353,In_1072);
nand U341 (N_341,In_2004,In_1795);
and U342 (N_342,In_1159,In_646);
xor U343 (N_343,In_1017,In_366);
or U344 (N_344,In_328,In_871);
or U345 (N_345,In_195,In_1769);
nand U346 (N_346,In_1111,In_691);
nor U347 (N_347,In_1854,In_1120);
nor U348 (N_348,In_1884,In_40);
and U349 (N_349,In_772,In_2106);
or U350 (N_350,In_1960,In_882);
and U351 (N_351,In_491,In_1810);
or U352 (N_352,In_51,In_1782);
or U353 (N_353,In_527,In_813);
nor U354 (N_354,In_2006,In_1474);
and U355 (N_355,In_679,In_344);
or U356 (N_356,In_1204,In_34);
or U357 (N_357,In_1729,In_2013);
nand U358 (N_358,In_608,In_2039);
nand U359 (N_359,In_364,In_820);
xnor U360 (N_360,In_938,In_793);
nor U361 (N_361,In_1340,In_1503);
nor U362 (N_362,In_609,In_1806);
or U363 (N_363,In_818,In_201);
nand U364 (N_364,In_1105,In_1924);
nor U365 (N_365,In_1402,In_250);
and U366 (N_366,In_1110,In_624);
nand U367 (N_367,In_1321,In_2201);
or U368 (N_368,In_665,In_588);
nor U369 (N_369,In_428,In_703);
or U370 (N_370,In_1465,In_2212);
nand U371 (N_371,In_1115,In_473);
and U372 (N_372,In_2241,In_1571);
and U373 (N_373,In_446,In_1525);
nor U374 (N_374,In_883,In_1421);
nor U375 (N_375,In_1266,In_12);
nor U376 (N_376,In_837,In_854);
nand U377 (N_377,In_1167,In_2249);
nor U378 (N_378,In_1812,In_1683);
nor U379 (N_379,In_1904,In_2222);
xnor U380 (N_380,In_2285,In_844);
and U381 (N_381,In_1639,In_284);
nand U382 (N_382,In_335,In_2247);
and U383 (N_383,In_1502,In_2101);
nand U384 (N_384,In_1788,In_1372);
and U385 (N_385,In_233,In_46);
nor U386 (N_386,In_1850,In_678);
xnor U387 (N_387,In_1107,In_9);
or U388 (N_388,In_797,In_2482);
nor U389 (N_389,In_461,In_842);
nand U390 (N_390,In_1578,In_1150);
and U391 (N_391,In_1761,In_2461);
xor U392 (N_392,In_2311,In_1557);
nor U393 (N_393,In_1853,In_1352);
nor U394 (N_394,In_1356,In_119);
nand U395 (N_395,In_1945,In_988);
or U396 (N_396,In_730,In_2443);
nor U397 (N_397,In_1902,In_574);
nor U398 (N_398,In_1568,In_159);
and U399 (N_399,In_1651,In_2310);
nor U400 (N_400,In_1305,In_26);
or U401 (N_401,In_696,In_1413);
and U402 (N_402,In_459,In_1636);
nor U403 (N_403,In_799,In_88);
and U404 (N_404,In_1985,In_1988);
nor U405 (N_405,In_1288,In_1384);
or U406 (N_406,In_903,In_565);
xnor U407 (N_407,In_557,In_1223);
or U408 (N_408,In_1640,In_1817);
xor U409 (N_409,In_158,In_1063);
or U410 (N_410,In_1184,In_663);
or U411 (N_411,In_213,In_2446);
nor U412 (N_412,In_592,In_1871);
nor U413 (N_413,In_782,In_628);
nor U414 (N_414,In_641,In_1808);
or U415 (N_415,In_152,In_1410);
nand U416 (N_416,In_242,In_1849);
or U417 (N_417,In_642,In_1248);
nor U418 (N_418,In_1185,In_2386);
or U419 (N_419,In_1219,In_155);
or U420 (N_420,In_53,In_688);
xor U421 (N_421,In_1543,In_1608);
nor U422 (N_422,In_910,In_2469);
and U423 (N_423,In_1089,In_913);
nor U424 (N_424,In_1286,In_1003);
nand U425 (N_425,In_294,In_246);
and U426 (N_426,In_334,In_2355);
nor U427 (N_427,In_1043,In_2423);
xnor U428 (N_428,In_901,In_873);
and U429 (N_429,In_1969,In_1919);
nor U430 (N_430,In_2322,In_2330);
nor U431 (N_431,In_1121,In_2073);
and U432 (N_432,In_569,In_2340);
nand U433 (N_433,In_1674,In_2474);
nand U434 (N_434,In_953,In_1367);
and U435 (N_435,In_1261,In_2135);
or U436 (N_436,In_1061,In_959);
or U437 (N_437,In_1490,In_1365);
or U438 (N_438,In_463,In_253);
xnor U439 (N_439,In_260,In_1405);
or U440 (N_440,In_1335,In_1203);
and U441 (N_441,In_1712,In_1182);
nand U442 (N_442,In_1328,In_45);
and U443 (N_443,In_734,In_1664);
nor U444 (N_444,In_89,In_1401);
nor U445 (N_445,In_701,In_2267);
nand U446 (N_446,In_499,In_1540);
or U447 (N_447,In_2079,In_1311);
and U448 (N_448,In_1620,In_1227);
xnor U449 (N_449,In_904,In_21);
or U450 (N_450,In_2202,In_273);
or U451 (N_451,In_129,In_1106);
or U452 (N_452,In_352,In_1768);
and U453 (N_453,In_1912,In_1889);
nor U454 (N_454,In_2231,In_441);
nor U455 (N_455,In_2057,In_300);
nand U456 (N_456,In_431,In_132);
and U457 (N_457,In_2356,In_1199);
and U458 (N_458,In_2268,In_2487);
and U459 (N_459,In_769,In_101);
nand U460 (N_460,In_394,In_1705);
and U461 (N_461,In_1586,In_1294);
nand U462 (N_462,In_1021,In_1224);
or U463 (N_463,In_1565,In_1530);
and U464 (N_464,In_1022,In_2277);
xnor U465 (N_465,In_148,In_438);
nand U466 (N_466,In_278,In_1028);
and U467 (N_467,In_1828,In_410);
nor U468 (N_468,In_2127,In_621);
and U469 (N_469,In_558,In_1486);
or U470 (N_470,In_167,In_236);
nor U471 (N_471,In_1964,In_1147);
and U472 (N_472,In_2095,In_2207);
nand U473 (N_473,In_740,In_1508);
and U474 (N_474,In_786,In_692);
xnor U475 (N_475,In_2304,In_2043);
or U476 (N_476,In_175,In_2140);
and U477 (N_477,In_190,In_1926);
nor U478 (N_478,In_649,In_2166);
nor U479 (N_479,In_1046,In_2415);
nor U480 (N_480,In_1353,In_832);
nand U481 (N_481,In_867,In_241);
nand U482 (N_482,In_2425,In_1001);
and U483 (N_483,In_530,In_163);
and U484 (N_484,In_2465,In_890);
nand U485 (N_485,In_2115,In_1746);
nand U486 (N_486,In_2290,In_776);
or U487 (N_487,In_590,In_2429);
and U488 (N_488,In_531,In_1941);
and U489 (N_489,In_784,In_1461);
xor U490 (N_490,In_676,In_2399);
nand U491 (N_491,In_2388,In_1104);
or U492 (N_492,In_468,In_1379);
nand U493 (N_493,In_1555,In_2100);
nor U494 (N_494,In_1445,In_1193);
or U495 (N_495,In_741,In_2245);
nand U496 (N_496,In_2018,In_1655);
nor U497 (N_497,In_23,In_1749);
nor U498 (N_498,In_234,In_1627);
nor U499 (N_499,In_787,In_138);
or U500 (N_500,In_1974,In_180);
nor U501 (N_501,In_1663,In_69);
nor U502 (N_502,In_1645,In_694);
and U503 (N_503,In_1095,In_247);
nor U504 (N_504,In_2334,In_1);
and U505 (N_505,In_1322,In_2283);
nor U506 (N_506,In_845,In_1142);
or U507 (N_507,In_2427,In_1437);
nand U508 (N_508,In_157,In_2129);
or U509 (N_509,In_2199,In_430);
and U510 (N_510,In_2237,In_729);
and U511 (N_511,In_41,In_1754);
or U512 (N_512,In_2072,In_1381);
xor U513 (N_513,In_1370,In_952);
and U514 (N_514,In_1787,In_330);
or U515 (N_515,In_1258,In_893);
xor U516 (N_516,In_1403,In_79);
nand U517 (N_517,In_1700,In_467);
xor U518 (N_518,In_1562,In_1329);
nand U519 (N_519,In_1064,In_603);
and U520 (N_520,In_874,In_436);
nand U521 (N_521,In_939,In_1019);
or U522 (N_522,In_2054,In_545);
and U523 (N_523,In_1757,In_888);
xor U524 (N_524,In_1012,In_1138);
and U525 (N_525,In_1837,In_2160);
and U526 (N_526,In_1628,In_390);
nor U527 (N_527,In_317,In_2270);
xnor U528 (N_528,In_664,In_852);
nand U529 (N_529,In_1915,In_517);
nor U530 (N_530,In_203,In_1027);
nand U531 (N_531,In_2050,In_1556);
nor U532 (N_532,In_583,In_1006);
nor U533 (N_533,In_2156,In_393);
and U534 (N_534,In_266,In_705);
or U535 (N_535,In_1619,In_1152);
or U536 (N_536,In_1696,In_1133);
nor U537 (N_537,In_853,In_168);
nor U538 (N_538,In_2407,In_2492);
nor U539 (N_539,In_2031,In_1128);
or U540 (N_540,In_2404,In_1615);
nand U541 (N_541,In_2462,In_1685);
and U542 (N_542,In_2223,In_523);
nand U543 (N_543,In_360,In_122);
nand U544 (N_544,In_2498,In_1400);
nor U545 (N_545,In_752,In_105);
nor U546 (N_546,In_2148,In_656);
nand U547 (N_547,In_2473,In_1980);
nor U548 (N_548,In_756,In_2213);
xor U549 (N_549,In_440,In_2016);
nand U550 (N_550,In_2120,In_416);
nand U551 (N_551,In_296,In_93);
and U552 (N_552,In_553,In_1877);
or U553 (N_553,In_1518,In_2300);
and U554 (N_554,In_1528,In_1387);
or U555 (N_555,In_1901,In_72);
or U556 (N_556,In_761,In_2170);
nand U557 (N_557,In_2051,In_192);
or U558 (N_558,In_2389,In_2143);
and U559 (N_559,In_2392,In_1920);
nand U560 (N_560,In_81,In_338);
or U561 (N_561,In_977,In_1348);
or U562 (N_562,In_966,In_85);
or U563 (N_563,In_1598,In_2426);
and U564 (N_564,In_98,In_2088);
nor U565 (N_565,In_918,In_2281);
nor U566 (N_566,In_48,In_2279);
xor U567 (N_567,In_1416,In_814);
nor U568 (N_568,In_1228,In_1238);
nand U569 (N_569,In_1344,In_1876);
nand U570 (N_570,In_1357,In_483);
nor U571 (N_571,In_1307,In_2015);
or U572 (N_572,In_323,In_17);
and U573 (N_573,In_1302,In_2360);
or U574 (N_574,In_452,In_402);
nand U575 (N_575,In_456,In_1783);
nand U576 (N_576,In_1454,In_1638);
and U577 (N_577,In_1961,In_1146);
nand U578 (N_578,In_2052,In_1459);
nand U579 (N_579,In_6,In_2489);
and U580 (N_580,In_2107,In_1070);
or U581 (N_581,In_1148,In_1295);
nand U582 (N_582,In_1745,In_2081);
or U583 (N_583,In_2257,In_808);
nor U584 (N_584,In_2227,In_419);
nand U585 (N_585,In_1298,In_2162);
nor U586 (N_586,In_1802,In_549);
nor U587 (N_587,In_2357,In_2110);
nor U588 (N_588,In_798,In_2154);
and U589 (N_589,In_403,In_1602);
nand U590 (N_590,In_1275,In_385);
or U591 (N_591,In_1574,In_1660);
and U592 (N_592,In_1976,In_1748);
nand U593 (N_593,In_1981,In_447);
or U594 (N_594,In_1723,In_1591);
nor U595 (N_595,In_232,In_880);
nor U596 (N_596,In_65,In_311);
nor U597 (N_597,In_860,In_1273);
or U598 (N_598,In_471,In_1042);
nand U599 (N_599,In_1829,In_1304);
nor U600 (N_600,In_254,In_2152);
and U601 (N_601,In_2299,In_348);
or U602 (N_602,In_619,In_125);
or U603 (N_603,In_1692,In_908);
nor U604 (N_604,In_1008,In_1385);
and U605 (N_605,In_1358,In_1947);
or U606 (N_606,In_1035,In_1181);
nand U607 (N_607,In_1840,In_1774);
nor U608 (N_608,In_2495,In_1607);
nand U609 (N_609,In_1386,In_474);
and U610 (N_610,In_2458,In_121);
nand U611 (N_611,In_1325,In_1399);
nor U612 (N_612,In_1075,In_1259);
or U613 (N_613,In_369,In_773);
nor U614 (N_614,In_1526,In_434);
or U615 (N_615,In_1494,In_587);
nor U616 (N_616,In_1618,In_2472);
and U617 (N_617,In_575,In_1939);
nand U618 (N_618,In_1438,In_1533);
or U619 (N_619,In_2055,In_342);
xnor U620 (N_620,In_104,In_329);
xnor U621 (N_621,In_1583,In_946);
nor U622 (N_622,In_2019,In_868);
and U623 (N_623,In_521,In_288);
nand U624 (N_624,In_524,In_1300);
nand U625 (N_625,In_2232,In_1735);
or U626 (N_626,In_1938,In_1521);
or U627 (N_627,In_916,In_1821);
and U628 (N_628,In_82,In_552);
nand U629 (N_629,In_2233,In_1350);
or U630 (N_630,In_862,In_1514);
nor U631 (N_631,In_973,In_1276);
nand U632 (N_632,In_1435,In_18);
nand U633 (N_633,In_2225,In_405);
or U634 (N_634,In_610,In_2041);
and U635 (N_635,In_771,In_494);
nor U636 (N_636,In_1601,In_162);
or U637 (N_637,In_8,In_224);
nand U638 (N_638,In_68,In_1242);
nand U639 (N_639,In_1560,In_965);
or U640 (N_640,In_2420,In_810);
nand U641 (N_641,In_2219,In_1029);
nand U642 (N_642,In_1260,In_297);
nand U643 (N_643,In_2048,In_2085);
or U644 (N_644,In_2218,In_2324);
nor U645 (N_645,In_1098,In_2302);
and U646 (N_646,In_2275,In_687);
nand U647 (N_647,In_1174,In_5);
nor U648 (N_648,In_1847,In_775);
or U649 (N_649,In_511,In_602);
and U650 (N_650,In_454,In_1145);
xnor U651 (N_651,In_528,In_1798);
and U652 (N_652,In_2009,In_870);
or U653 (N_653,In_924,In_243);
or U654 (N_654,In_3,In_1240);
nor U655 (N_655,In_1044,In_316);
and U656 (N_656,In_707,In_1955);
or U657 (N_657,In_237,In_1844);
nand U658 (N_658,In_783,In_2159);
nor U659 (N_659,In_1897,In_1661);
and U660 (N_660,In_539,In_1176);
nor U661 (N_661,In_2074,In_380);
or U662 (N_662,In_1178,In_2397);
and U663 (N_663,In_1549,In_2070);
xor U664 (N_664,In_27,In_1695);
nand U665 (N_665,In_1872,In_1241);
nand U666 (N_666,In_1417,In_2362);
or U667 (N_667,In_1069,In_1542);
nor U668 (N_668,In_1125,In_1141);
nand U669 (N_669,In_131,In_932);
nor U670 (N_670,In_1285,In_1682);
and U671 (N_671,In_1065,In_1126);
and U672 (N_672,In_1144,In_1990);
xnor U673 (N_673,In_2188,In_2255);
xor U674 (N_674,In_2133,In_1341);
nor U675 (N_675,In_1934,In_1544);
xnor U676 (N_676,In_895,In_1970);
nor U677 (N_677,In_697,In_1906);
or U678 (N_678,In_78,In_1183);
and U679 (N_679,In_2192,In_1081);
nand U680 (N_680,In_2408,In_2248);
and U681 (N_681,In_1436,In_2238);
nand U682 (N_682,In_1841,In_1866);
and U683 (N_683,In_885,In_226);
and U684 (N_684,In_1209,In_1091);
and U685 (N_685,In_2032,In_604);
nand U686 (N_686,In_1617,In_1958);
xor U687 (N_687,In_2035,In_2380);
and U688 (N_688,In_1606,In_331);
or U689 (N_689,In_936,In_2313);
and U690 (N_690,In_299,In_1584);
nand U691 (N_691,In_751,In_1052);
nor U692 (N_692,In_1650,In_193);
nor U693 (N_693,In_1805,In_766);
and U694 (N_694,In_1564,In_1545);
nand U695 (N_695,In_1878,In_1267);
nor U696 (N_696,In_1572,In_1858);
and U697 (N_697,In_94,In_1453);
nand U698 (N_698,In_2338,In_1524);
nand U699 (N_699,In_2282,In_2099);
nor U700 (N_700,In_2189,In_1681);
and U701 (N_701,In_188,In_770);
xor U702 (N_702,In_2228,In_923);
and U703 (N_703,In_371,In_718);
nand U704 (N_704,In_1342,In_644);
nor U705 (N_705,In_1020,In_1764);
xor U706 (N_706,In_823,In_1862);
or U707 (N_707,In_675,In_2347);
nor U708 (N_708,In_958,In_1360);
or U709 (N_709,In_519,In_1213);
or U710 (N_710,In_1998,In_865);
nand U711 (N_711,In_185,In_1279);
or U712 (N_712,In_2440,In_1596);
nand U713 (N_713,In_1446,In_906);
nand U714 (N_714,In_922,In_846);
xnor U715 (N_715,In_2242,In_1163);
nand U716 (N_716,In_325,In_140);
or U717 (N_717,In_97,In_1676);
nand U718 (N_718,In_654,In_153);
and U719 (N_719,In_2371,In_2090);
or U720 (N_720,In_302,In_1337);
nor U721 (N_721,In_1765,In_466);
and U722 (N_722,In_2053,In_712);
and U723 (N_723,In_1092,In_1200);
nor U724 (N_724,In_2007,In_1407);
xnor U725 (N_725,In_614,In_500);
and U726 (N_726,In_1351,In_2390);
xor U727 (N_727,In_2253,In_2366);
nand U728 (N_728,In_1217,In_1349);
and U729 (N_729,In_1716,In_1333);
or U730 (N_730,In_367,In_999);
or U731 (N_731,In_111,In_829);
xor U732 (N_732,In_126,In_64);
xor U733 (N_733,In_1277,In_2384);
or U734 (N_734,In_2182,In_1775);
nand U735 (N_735,In_991,In_1250);
and U736 (N_736,In_960,In_2476);
xnor U737 (N_737,In_781,In_525);
xor U738 (N_738,In_435,In_1648);
or U739 (N_739,In_2286,In_220);
nand U740 (N_740,In_1313,In_135);
and U741 (N_741,In_312,In_95);
nand U742 (N_742,In_828,In_1635);
nor U743 (N_743,In_1576,In_616);
nand U744 (N_744,In_225,In_437);
nor U745 (N_745,In_1253,In_115);
or U746 (N_746,In_409,In_110);
nor U747 (N_747,In_0,In_1054);
and U748 (N_748,In_516,In_1684);
xnor U749 (N_749,In_280,In_643);
and U750 (N_750,In_14,In_1561);
nand U751 (N_751,In_1894,In_362);
or U752 (N_752,In_1701,In_270);
or U753 (N_753,In_375,In_512);
or U754 (N_754,In_30,In_1603);
or U755 (N_755,In_2308,In_2091);
or U756 (N_756,In_1658,In_2215);
xnor U757 (N_757,In_1709,In_305);
and U758 (N_758,In_2130,In_2058);
or U759 (N_759,In_1908,In_1918);
nor U760 (N_760,In_1473,In_1315);
nand U761 (N_761,In_1031,In_622);
and U762 (N_762,In_1262,In_2068);
and U763 (N_763,In_2066,In_1268);
nand U764 (N_764,In_2481,In_840);
and U765 (N_765,In_894,In_413);
or U766 (N_766,In_540,In_1944);
nand U767 (N_767,In_926,In_2003);
xor U768 (N_768,In_1815,In_421);
nor U769 (N_769,In_1444,In_735);
or U770 (N_770,In_2485,In_2331);
nand U771 (N_771,In_1394,In_1869);
and U772 (N_772,In_1216,In_640);
nor U773 (N_773,In_2172,In_2069);
nor U774 (N_774,In_381,In_1708);
and U775 (N_775,In_489,In_1280);
nor U776 (N_776,In_1513,In_1794);
nor U777 (N_777,In_1195,In_1625);
nand U778 (N_778,In_1978,In_554);
or U779 (N_779,In_1809,In_70);
nand U780 (N_780,In_716,In_2317);
nand U781 (N_781,In_303,In_891);
xnor U782 (N_782,In_1956,In_824);
and U783 (N_783,In_2042,In_2477);
nor U784 (N_784,In_2082,In_1369);
nor U785 (N_785,In_630,In_2169);
and U786 (N_786,In_1623,In_1510);
nor U787 (N_787,In_1050,In_2422);
or U788 (N_788,In_2200,In_1318);
nand U789 (N_789,In_1234,In_788);
or U790 (N_790,In_1937,In_636);
nor U791 (N_791,In_310,In_102);
and U792 (N_792,In_2432,In_1538);
nand U793 (N_793,In_1374,In_1319);
or U794 (N_794,In_462,In_863);
nand U795 (N_795,In_964,In_103);
or U796 (N_796,In_1517,In_2332);
and U797 (N_797,In_22,In_750);
and U798 (N_798,In_2119,In_1744);
or U799 (N_799,In_1066,In_1721);
or U800 (N_800,In_1927,In_736);
nor U801 (N_801,In_376,In_354);
nand U802 (N_802,In_2008,In_2369);
nor U803 (N_803,In_1675,In_10);
and U804 (N_804,In_1644,In_551);
nor U805 (N_805,In_422,In_320);
xor U806 (N_806,In_801,In_42);
nand U807 (N_807,In_206,In_2488);
or U808 (N_808,In_314,In_1824);
or U809 (N_809,In_209,In_2451);
nand U810 (N_810,In_2177,In_765);
xor U811 (N_811,In_1088,In_618);
nand U812 (N_812,In_984,In_830);
nor U813 (N_813,In_892,In_1117);
nor U814 (N_814,In_1477,In_1913);
nor U815 (N_815,In_2186,In_281);
nand U816 (N_816,In_2125,In_1225);
nor U817 (N_817,In_426,In_1931);
and U818 (N_818,In_1762,In_986);
nor U819 (N_819,In_1274,In_2348);
and U820 (N_820,In_2083,In_695);
nand U821 (N_821,In_982,In_2367);
and U822 (N_822,In_2002,In_146);
nor U823 (N_823,In_1704,In_690);
and U824 (N_824,In_62,In_704);
and U825 (N_825,In_2497,In_648);
or U826 (N_826,In_535,In_301);
nand U827 (N_827,In_368,In_1826);
and U828 (N_828,In_1599,In_2448);
nand U829 (N_829,In_1229,In_1999);
and U830 (N_830,In_931,In_1496);
nor U831 (N_831,In_90,In_347);
nand U832 (N_832,In_2184,In_114);
or U833 (N_833,In_1519,In_2076);
or U834 (N_834,In_1208,In_709);
or U835 (N_835,In_2209,In_698);
and U836 (N_836,In_1491,In_2478);
nand U837 (N_837,In_1634,In_1929);
nand U838 (N_838,In_1013,In_1151);
and U839 (N_839,In_1827,In_1114);
nor U840 (N_840,In_1284,In_2109);
xor U841 (N_841,In_1861,In_900);
or U842 (N_842,In_1631,In_1822);
or U843 (N_843,In_130,In_1767);
xnor U844 (N_844,In_141,In_1469);
and U845 (N_845,In_2010,In_1739);
xnor U846 (N_846,In_1424,In_1296);
nand U847 (N_847,In_599,In_1423);
and U848 (N_848,In_268,In_210);
nand U849 (N_849,In_1507,In_1679);
nand U850 (N_850,In_2151,In_128);
or U851 (N_851,In_1622,In_1710);
and U852 (N_852,In_972,In_1686);
nor U853 (N_853,In_383,In_61);
nor U854 (N_854,In_1190,In_2321);
or U855 (N_855,In_1820,In_613);
and U856 (N_856,In_1415,In_1694);
nand U857 (N_857,In_444,In_1478);
nor U858 (N_858,In_708,In_2114);
and U859 (N_859,In_432,In_838);
nand U860 (N_860,In_1873,In_907);
nand U861 (N_861,In_1482,In_591);
and U862 (N_862,In_2157,In_1071);
and U863 (N_863,In_1447,In_275);
xor U864 (N_864,In_264,In_1197);
nor U865 (N_865,In_324,In_626);
xor U866 (N_866,In_295,In_1497);
xor U867 (N_867,In_2176,In_2217);
nor U868 (N_868,In_1737,In_1039);
nand U869 (N_869,In_746,In_1032);
or U870 (N_870,In_387,In_2341);
nor U871 (N_871,In_2431,In_2174);
nand U872 (N_872,In_1082,In_184);
or U873 (N_873,In_11,In_377);
nand U874 (N_874,In_1553,In_943);
xor U875 (N_875,In_768,In_2289);
and U876 (N_876,In_1175,In_1378);
or U877 (N_877,In_2045,In_386);
nor U878 (N_878,In_925,In_683);
xnor U879 (N_879,In_949,In_802);
and U880 (N_880,In_2128,In_1536);
nor U881 (N_881,In_600,In_634);
nor U882 (N_882,In_2358,In_400);
nor U883 (N_883,In_2193,In_407);
nor U884 (N_884,In_898,In_2269);
or U885 (N_885,In_758,In_2104);
and U886 (N_886,In_755,In_1323);
xnor U887 (N_887,In_1688,In_855);
or U888 (N_888,In_2134,In_1790);
nor U889 (N_889,In_1909,In_113);
nor U890 (N_890,In_1778,In_1699);
or U891 (N_891,In_1652,In_1773);
nor U892 (N_892,In_847,In_1187);
and U893 (N_893,In_1018,In_831);
nor U894 (N_894,In_1632,In_2027);
xnor U895 (N_895,In_2036,In_389);
nand U896 (N_896,In_457,In_1314);
nor U897 (N_897,In_2442,In_1196);
nand U898 (N_898,In_1698,In_50);
xor U899 (N_899,In_886,In_1484);
nand U900 (N_900,In_1983,In_1487);
and U901 (N_901,In_2499,In_107);
nand U902 (N_902,In_1846,In_2428);
nor U903 (N_903,In_2320,In_35);
and U904 (N_904,In_2234,In_1149);
nand U905 (N_905,In_1914,In_2265);
nand U906 (N_906,In_1763,In_1215);
nand U907 (N_907,In_1921,In_754);
or U908 (N_908,In_611,In_1498);
and U909 (N_909,In_1797,In_214);
nor U910 (N_910,In_1388,In_1910);
xnor U911 (N_911,In_170,In_1818);
nand U912 (N_912,In_127,In_2145);
or U913 (N_913,In_930,In_1002);
nand U914 (N_914,In_60,In_1932);
or U915 (N_915,In_762,In_2272);
and U916 (N_916,In_992,In_1074);
nand U917 (N_917,In_2175,In_37);
nand U918 (N_918,In_2496,In_759);
or U919 (N_919,In_2185,In_1221);
or U920 (N_920,In_1731,In_2105);
and U921 (N_921,In_2438,In_1776);
nand U922 (N_922,In_36,In_1236);
xnor U923 (N_923,In_169,In_1339);
nor U924 (N_924,In_1537,In_1550);
and U925 (N_925,In_1715,In_1755);
nand U926 (N_926,In_1680,In_561);
nor U927 (N_927,In_504,In_1766);
nand U928 (N_928,In_1249,In_689);
nand U929 (N_929,In_1257,In_876);
and U930 (N_930,In_2113,In_1500);
or U931 (N_931,In_1950,In_1732);
nand U932 (N_932,In_1122,In_651);
or U933 (N_933,In_835,In_715);
and U934 (N_934,In_1836,In_2256);
or U935 (N_935,In_556,In_1090);
nand U936 (N_936,In_382,In_1011);
xor U937 (N_937,In_57,In_2309);
xor U938 (N_938,In_1541,In_2424);
nand U939 (N_939,In_1547,In_1951);
nor U940 (N_940,In_571,In_227);
nor U941 (N_941,In_2271,In_721);
xor U942 (N_942,In_1231,In_487);
nand U943 (N_943,In_1364,In_915);
and U944 (N_944,In_197,In_67);
and U945 (N_945,In_2163,In_464);
xor U946 (N_946,In_1158,In_812);
xnor U947 (N_947,In_878,In_216);
nand U948 (N_948,In_744,In_2316);
nand U949 (N_949,In_1034,In_1025);
and U950 (N_950,In_1409,In_74);
nand U951 (N_951,In_1136,In_2276);
and U952 (N_952,In_2391,In_2450);
or U953 (N_953,In_196,In_1480);
nand U954 (N_954,In_1898,In_1396);
and U955 (N_955,In_1023,In_815);
and U956 (N_956,In_1281,In_2178);
nor U957 (N_957,In_2328,In_470);
nor U958 (N_958,In_1255,In_399);
and U959 (N_959,In_1539,In_1807);
and U960 (N_960,In_204,In_443);
nand U961 (N_961,In_711,In_1427);
and U962 (N_962,In_1719,In_321);
or U963 (N_963,In_1312,In_174);
nand U964 (N_964,In_1112,In_2024);
nor U965 (N_965,In_827,In_980);
or U966 (N_966,In_2239,In_1180);
xnor U967 (N_967,In_2460,In_2167);
nor U968 (N_968,In_631,In_1230);
nand U969 (N_969,In_856,In_165);
xor U970 (N_970,In_1422,In_1600);
and U971 (N_971,In_1852,In_285);
and U972 (N_972,In_2092,In_423);
and U973 (N_973,In_962,In_2379);
and U974 (N_974,In_637,In_1863);
nand U975 (N_975,In_1428,In_2096);
nor U976 (N_976,In_230,In_142);
nand U977 (N_977,In_2377,In_722);
xor U978 (N_978,In_2398,In_1535);
nor U979 (N_979,In_821,In_356);
and U980 (N_980,In_2278,In_1330);
and U981 (N_981,In_1103,In_912);
nand U982 (N_982,In_2333,In_1646);
and U983 (N_983,In_577,In_727);
and U984 (N_984,In_1123,In_2363);
and U985 (N_985,In_2005,In_674);
and U986 (N_986,In_2433,In_1851);
nor U987 (N_987,In_374,In_1129);
nand U988 (N_988,In_1779,In_143);
and U989 (N_989,In_713,In_2235);
and U990 (N_990,In_2026,In_1086);
nand U991 (N_991,In_794,In_2315);
xor U992 (N_992,In_1079,In_804);
nand U993 (N_993,In_395,In_2417);
nor U994 (N_994,In_484,In_2061);
nand U995 (N_995,In_1373,In_2396);
nand U996 (N_996,In_1359,In_63);
or U997 (N_997,In_2158,In_1668);
nor U998 (N_998,In_1245,In_2142);
and U999 (N_999,In_455,In_1579);
and U1000 (N_1000,In_333,In_1758);
and U1001 (N_1001,In_1563,In_659);
and U1002 (N_1002,In_1750,In_2060);
nand U1003 (N_1003,In_507,In_1398);
and U1004 (N_1004,In_1582,In_2183);
nand U1005 (N_1005,In_2028,In_1432);
nor U1006 (N_1006,In_1559,In_1346);
or U1007 (N_1007,In_465,In_2210);
xnor U1008 (N_1008,In_286,In_84);
nand U1009 (N_1009,In_513,In_2064);
nor U1010 (N_1010,In_2368,In_1875);
nor U1011 (N_1011,In_340,In_1614);
nand U1012 (N_1012,In_2124,In_28);
and U1013 (N_1013,In_2435,In_1493);
xor U1014 (N_1014,In_2359,In_917);
nand U1015 (N_1015,In_542,In_1354);
or U1016 (N_1016,In_1479,In_1590);
and U1017 (N_1017,In_1463,In_1102);
and U1018 (N_1018,In_398,In_2383);
or U1019 (N_1019,In_1997,In_1986);
nand U1020 (N_1020,In_702,In_1534);
nand U1021 (N_1021,In_1448,In_724);
nor U1022 (N_1022,In_244,In_291);
and U1023 (N_1023,In_1331,In_1609);
nand U1024 (N_1024,In_757,In_1551);
or U1025 (N_1025,In_1450,In_1738);
nand U1026 (N_1026,In_1492,In_1132);
and U1027 (N_1027,In_476,In_379);
nor U1028 (N_1028,In_150,In_315);
nor U1029 (N_1029,In_397,In_106);
or U1030 (N_1030,In_277,In_869);
and U1031 (N_1031,In_671,In_503);
nand U1032 (N_1032,In_238,In_370);
and U1033 (N_1033,In_685,In_606);
or U1034 (N_1034,In_1740,In_1925);
and U1035 (N_1035,In_969,In_2305);
nor U1036 (N_1036,In_2414,In_566);
nand U1037 (N_1037,In_287,In_1979);
nand U1038 (N_1038,In_182,In_1109);
nand U1039 (N_1039,In_2029,In_502);
and U1040 (N_1040,In_1803,In_1722);
and U1041 (N_1041,In_1647,In_349);
and U1042 (N_1042,In_994,In_1326);
nor U1043 (N_1043,In_2034,In_725);
or U1044 (N_1044,In_2187,In_363);
and U1045 (N_1045,In_1495,In_2);
nor U1046 (N_1046,In_546,In_807);
nor U1047 (N_1047,In_1771,In_448);
nand U1048 (N_1048,In_1804,In_2466);
xor U1049 (N_1049,In_593,In_472);
nor U1050 (N_1050,In_714,In_453);
and U1051 (N_1051,In_1566,In_749);
or U1052 (N_1052,In_20,In_1060);
nand U1053 (N_1053,In_2339,In_607);
xor U1054 (N_1054,In_1243,In_2146);
and U1055 (N_1055,In_274,In_2001);
nor U1056 (N_1056,In_928,In_109);
nor U1057 (N_1057,In_1239,In_534);
and U1058 (N_1058,In_2403,In_1165);
nand U1059 (N_1059,In_160,In_780);
nor U1060 (N_1060,In_887,In_2164);
or U1061 (N_1061,In_1966,In_2375);
nand U1062 (N_1062,In_1991,In_2093);
or U1063 (N_1063,In_2436,In_1546);
nand U1064 (N_1064,In_1211,In_816);
nand U1065 (N_1065,In_492,In_929);
and U1066 (N_1066,In_1940,In_726);
nand U1067 (N_1067,In_2098,In_529);
nand U1068 (N_1068,In_2294,In_1752);
nor U1069 (N_1069,In_879,In_1713);
xor U1070 (N_1070,In_401,In_2374);
nor U1071 (N_1071,In_161,In_2136);
or U1072 (N_1072,In_1201,In_568);
and U1073 (N_1073,In_332,In_219);
nor U1074 (N_1074,In_1441,In_937);
nor U1075 (N_1075,In_1604,In_902);
or U1076 (N_1076,In_1000,In_576);
or U1077 (N_1077,In_1143,In_2224);
xor U1078 (N_1078,In_378,In_1041);
and U1079 (N_1079,In_418,In_1499);
and U1080 (N_1080,In_1665,In_1278);
and U1081 (N_1081,In_1397,In_2454);
nand U1082 (N_1082,In_1140,In_2131);
nand U1083 (N_1083,In_1189,In_717);
xnor U1084 (N_1084,In_263,In_1458);
or U1085 (N_1085,In_449,In_961);
and U1086 (N_1086,In_2445,In_1629);
nor U1087 (N_1087,In_1886,In_1996);
nand U1088 (N_1088,In_657,In_145);
nor U1089 (N_1089,In_1659,In_1455);
nor U1090 (N_1090,In_1811,In_198);
or U1091 (N_1091,In_1895,In_2141);
and U1092 (N_1092,In_1324,In_1697);
xnor U1093 (N_1093,In_1657,In_1390);
or U1094 (N_1094,In_1062,In_151);
nor U1095 (N_1095,In_652,In_1756);
and U1096 (N_1096,In_406,In_417);
xnor U1097 (N_1097,In_2021,In_1848);
nor U1098 (N_1098,In_223,In_1264);
or U1099 (N_1099,In_670,In_2453);
and U1100 (N_1100,In_1080,In_2208);
and U1101 (N_1101,In_211,In_2173);
xor U1102 (N_1102,In_742,In_1943);
and U1103 (N_1103,In_66,In_1896);
nand U1104 (N_1104,In_120,In_309);
nand U1105 (N_1105,In_2038,In_536);
and U1106 (N_1106,In_252,In_292);
nor U1107 (N_1107,In_116,In_1376);
nor U1108 (N_1108,In_1613,In_1656);
and U1109 (N_1109,In_2250,In_1612);
nand U1110 (N_1110,In_189,In_420);
nor U1111 (N_1111,In_2326,In_433);
nor U1112 (N_1112,In_1056,In_2468);
nor U1113 (N_1113,In_598,In_2413);
or U1114 (N_1114,In_789,In_791);
nand U1115 (N_1115,In_981,In_2204);
or U1116 (N_1116,In_1772,In_1170);
nor U1117 (N_1117,In_1246,In_173);
and U1118 (N_1118,In_2405,In_326);
and U1119 (N_1119,In_480,In_1885);
xnor U1120 (N_1120,In_1558,In_1567);
nor U1121 (N_1121,In_1691,In_720);
or U1122 (N_1122,In_194,In_623);
xor U1123 (N_1123,In_1310,In_944);
and U1124 (N_1124,In_1903,In_1577);
nand U1125 (N_1125,In_4,In_1026);
nor U1126 (N_1126,In_1449,In_1036);
or U1127 (N_1127,In_1882,In_559);
nor U1128 (N_1128,In_2132,In_978);
xnor U1129 (N_1129,In_1162,In_1588);
xnor U1130 (N_1130,In_2421,In_2402);
nand U1131 (N_1131,In_1067,In_7);
nand U1132 (N_1132,In_1654,In_365);
nand U1133 (N_1133,In_514,In_843);
nand U1134 (N_1134,In_87,In_1451);
nor U1135 (N_1135,In_2295,In_1865);
nand U1136 (N_1136,In_567,In_942);
nor U1137 (N_1137,In_2077,In_1643);
xnor U1138 (N_1138,In_506,In_2343);
or U1139 (N_1139,In_355,In_1058);
and U1140 (N_1140,In_1957,In_645);
nand U1141 (N_1141,In_2372,In_75);
nor U1142 (N_1142,In_1911,In_205);
and U1143 (N_1143,In_1334,In_272);
nand U1144 (N_1144,In_1527,In_2393);
and U1145 (N_1145,In_1287,In_501);
nand U1146 (N_1146,In_927,In_834);
nand U1147 (N_1147,In_933,In_1515);
nand U1148 (N_1148,In_1327,In_2044);
xnor U1149 (N_1149,In_2329,In_24);
nor U1150 (N_1150,In_1157,In_2412);
or U1151 (N_1151,In_1839,In_2012);
nor U1152 (N_1152,In_864,In_359);
nand U1153 (N_1153,In_2062,In_2197);
nor U1154 (N_1154,In_2161,In_1531);
or U1155 (N_1155,In_178,In_1923);
and U1156 (N_1156,In_1464,In_1948);
or U1157 (N_1157,In_1411,In_200);
and U1158 (N_1158,In_1516,In_2434);
nor U1159 (N_1159,In_2307,In_1235);
and U1160 (N_1160,In_2457,In_1905);
and U1161 (N_1161,In_100,In_1595);
nor U1162 (N_1162,In_779,In_2444);
nand U1163 (N_1163,In_1096,In_1226);
nand U1164 (N_1164,In_262,In_1845);
xnor U1165 (N_1165,In_1784,In_1689);
nand U1166 (N_1166,In_1014,In_2297);
nor U1167 (N_1167,In_2181,In_1457);
or U1168 (N_1168,In_2346,In_1483);
and U1169 (N_1169,In_1649,In_86);
nor U1170 (N_1170,In_2216,In_429);
nor U1171 (N_1171,In_660,In_1759);
and U1172 (N_1172,In_322,In_699);
nor U1173 (N_1173,In_2354,In_1907);
and U1174 (N_1174,In_1362,In_2352);
nor U1175 (N_1175,In_1452,In_388);
or U1176 (N_1176,In_1137,In_737);
xnor U1177 (N_1177,In_43,In_1087);
and U1178 (N_1178,In_963,In_747);
or U1179 (N_1179,In_2191,In_875);
nand U1180 (N_1180,In_1870,In_586);
or U1181 (N_1181,In_1942,In_661);
nor U1182 (N_1182,In_498,In_803);
nor U1183 (N_1183,In_2084,In_1171);
nand U1184 (N_1184,In_55,In_1368);
and U1185 (N_1185,In_2419,In_1843);
and U1186 (N_1186,In_983,In_1677);
and U1187 (N_1187,In_2097,In_2075);
or U1188 (N_1188,In_133,In_308);
xor U1189 (N_1189,In_1355,In_1053);
nor U1190 (N_1190,In_91,In_229);
and U1191 (N_1191,In_1076,In_2102);
or U1192 (N_1192,In_222,In_1972);
nand U1193 (N_1193,In_451,In_1218);
nand U1194 (N_1194,In_166,In_1830);
xor U1195 (N_1195,In_1289,In_1747);
and U1196 (N_1196,In_601,In_1859);
nor U1197 (N_1197,In_1523,In_83);
nand U1198 (N_1198,In_993,In_2416);
nor U1199 (N_1199,In_1383,In_458);
and U1200 (N_1200,In_1504,In_1168);
nor U1201 (N_1201,In_1085,In_2198);
and U1202 (N_1202,In_672,In_1670);
nand U1203 (N_1203,In_578,In_859);
xor U1204 (N_1204,In_1254,In_2171);
nor U1205 (N_1205,In_1166,In_1282);
or U1206 (N_1206,In_1425,In_181);
and U1207 (N_1207,In_1057,In_1989);
xor U1208 (N_1208,In_680,In_997);
or U1209 (N_1209,In_2336,In_995);
nor U1210 (N_1210,In_1084,In_475);
or U1211 (N_1211,In_1819,In_31);
and U1212 (N_1212,In_1672,In_134);
or U1213 (N_1213,In_1743,In_47);
nand U1214 (N_1214,In_1442,In_2246);
nor U1215 (N_1215,In_1987,In_1099);
nand U1216 (N_1216,In_495,In_2220);
and U1217 (N_1217,In_508,In_1760);
or U1218 (N_1218,In_1777,In_2260);
nor U1219 (N_1219,In_1100,In_1718);
nand U1220 (N_1220,In_179,In_1501);
and U1221 (N_1221,In_1610,In_955);
nor U1222 (N_1222,In_1965,In_2147);
and U1223 (N_1223,In_2011,In_1380);
nor U1224 (N_1224,In_391,In_1169);
and U1225 (N_1225,In_2049,In_760);
or U1226 (N_1226,In_1785,In_1860);
nor U1227 (N_1227,In_1391,In_1055);
and U1228 (N_1228,In_2211,In_2463);
nand U1229 (N_1229,In_719,In_1124);
and U1230 (N_1230,In_1742,In_667);
nor U1231 (N_1231,In_1730,In_706);
nor U1232 (N_1232,In_956,In_186);
nor U1233 (N_1233,In_307,In_486);
xnor U1234 (N_1234,In_99,In_240);
nand U1235 (N_1235,In_411,In_217);
nor U1236 (N_1236,In_594,In_1813);
and U1237 (N_1237,In_2441,In_1272);
and U1238 (N_1238,In_1592,In_1429);
and U1239 (N_1239,In_792,In_597);
or U1240 (N_1240,In_1059,In_2117);
or U1241 (N_1241,In_2046,In_478);
xor U1242 (N_1242,In_1214,In_866);
nand U1243 (N_1243,In_841,In_1867);
nor U1244 (N_1244,In_1161,In_1792);
nor U1245 (N_1245,In_1252,In_1770);
or U1246 (N_1246,In_653,In_1005);
or U1247 (N_1247,In_1119,In_118);
xor U1248 (N_1248,In_595,In_1347);
nand U1249 (N_1249,In_2252,In_612);
nand U1250 (N_1250,In_2182,In_1036);
and U1251 (N_1251,In_1840,In_825);
and U1252 (N_1252,In_927,In_583);
or U1253 (N_1253,In_2112,In_2176);
nor U1254 (N_1254,In_1958,In_227);
nor U1255 (N_1255,In_1769,In_1661);
and U1256 (N_1256,In_1310,In_1391);
nor U1257 (N_1257,In_1973,In_603);
and U1258 (N_1258,In_1418,In_1017);
nor U1259 (N_1259,In_2355,In_446);
or U1260 (N_1260,In_546,In_140);
and U1261 (N_1261,In_2309,In_1918);
nand U1262 (N_1262,In_2470,In_567);
or U1263 (N_1263,In_521,In_2171);
nor U1264 (N_1264,In_663,In_2360);
and U1265 (N_1265,In_101,In_1419);
and U1266 (N_1266,In_2064,In_208);
or U1267 (N_1267,In_2414,In_1277);
nor U1268 (N_1268,In_503,In_1834);
nor U1269 (N_1269,In_718,In_574);
xnor U1270 (N_1270,In_2155,In_2111);
and U1271 (N_1271,In_288,In_1293);
nor U1272 (N_1272,In_746,In_2118);
and U1273 (N_1273,In_823,In_2085);
nand U1274 (N_1274,In_55,In_151);
and U1275 (N_1275,In_799,In_2363);
and U1276 (N_1276,In_48,In_305);
and U1277 (N_1277,In_1517,In_2350);
and U1278 (N_1278,In_1177,In_2097);
nor U1279 (N_1279,In_405,In_2009);
nand U1280 (N_1280,In_1139,In_2448);
and U1281 (N_1281,In_1840,In_2108);
nor U1282 (N_1282,In_1566,In_2348);
xor U1283 (N_1283,In_708,In_2201);
xor U1284 (N_1284,In_991,In_1151);
and U1285 (N_1285,In_2313,In_605);
nand U1286 (N_1286,In_1613,In_253);
or U1287 (N_1287,In_199,In_313);
and U1288 (N_1288,In_1461,In_152);
nor U1289 (N_1289,In_446,In_1234);
or U1290 (N_1290,In_1905,In_303);
nand U1291 (N_1291,In_1616,In_2398);
or U1292 (N_1292,In_901,In_277);
xor U1293 (N_1293,In_2179,In_1064);
and U1294 (N_1294,In_428,In_2380);
and U1295 (N_1295,In_563,In_252);
xor U1296 (N_1296,In_2009,In_1625);
nand U1297 (N_1297,In_694,In_2481);
nand U1298 (N_1298,In_1062,In_1391);
xor U1299 (N_1299,In_332,In_589);
xor U1300 (N_1300,In_1734,In_200);
or U1301 (N_1301,In_864,In_29);
nand U1302 (N_1302,In_755,In_310);
or U1303 (N_1303,In_1970,In_2134);
nand U1304 (N_1304,In_2186,In_2441);
or U1305 (N_1305,In_2355,In_1218);
and U1306 (N_1306,In_1443,In_60);
xnor U1307 (N_1307,In_1836,In_635);
or U1308 (N_1308,In_533,In_1854);
and U1309 (N_1309,In_791,In_426);
nand U1310 (N_1310,In_1842,In_1371);
nand U1311 (N_1311,In_927,In_1219);
xor U1312 (N_1312,In_1543,In_960);
or U1313 (N_1313,In_169,In_640);
or U1314 (N_1314,In_1013,In_1949);
and U1315 (N_1315,In_2049,In_1005);
or U1316 (N_1316,In_399,In_889);
or U1317 (N_1317,In_1566,In_1929);
or U1318 (N_1318,In_2254,In_620);
nor U1319 (N_1319,In_1431,In_555);
and U1320 (N_1320,In_144,In_817);
nor U1321 (N_1321,In_1792,In_1696);
xnor U1322 (N_1322,In_963,In_501);
or U1323 (N_1323,In_1081,In_1935);
nand U1324 (N_1324,In_2413,In_1475);
nand U1325 (N_1325,In_1212,In_395);
xnor U1326 (N_1326,In_774,In_379);
or U1327 (N_1327,In_729,In_1281);
and U1328 (N_1328,In_237,In_1441);
nand U1329 (N_1329,In_2233,In_2483);
xor U1330 (N_1330,In_744,In_2219);
nor U1331 (N_1331,In_708,In_841);
nand U1332 (N_1332,In_713,In_1400);
and U1333 (N_1333,In_1205,In_1689);
or U1334 (N_1334,In_1631,In_1493);
nand U1335 (N_1335,In_259,In_454);
and U1336 (N_1336,In_618,In_1721);
and U1337 (N_1337,In_1877,In_1247);
and U1338 (N_1338,In_2002,In_969);
nor U1339 (N_1339,In_320,In_1750);
nand U1340 (N_1340,In_2159,In_1330);
nand U1341 (N_1341,In_1732,In_1536);
and U1342 (N_1342,In_723,In_1392);
or U1343 (N_1343,In_1340,In_1224);
nand U1344 (N_1344,In_2074,In_1121);
or U1345 (N_1345,In_2372,In_1809);
and U1346 (N_1346,In_2106,In_2360);
or U1347 (N_1347,In_2327,In_480);
nor U1348 (N_1348,In_1069,In_2172);
nand U1349 (N_1349,In_2472,In_1131);
nor U1350 (N_1350,In_456,In_1750);
xor U1351 (N_1351,In_2270,In_2039);
and U1352 (N_1352,In_780,In_874);
xor U1353 (N_1353,In_2401,In_893);
nor U1354 (N_1354,In_2181,In_1670);
nor U1355 (N_1355,In_1215,In_2023);
and U1356 (N_1356,In_1005,In_2343);
xor U1357 (N_1357,In_638,In_221);
or U1358 (N_1358,In_599,In_1914);
nand U1359 (N_1359,In_1577,In_1557);
or U1360 (N_1360,In_1571,In_2301);
nor U1361 (N_1361,In_2192,In_63);
xor U1362 (N_1362,In_755,In_1491);
nand U1363 (N_1363,In_1890,In_398);
nor U1364 (N_1364,In_1477,In_56);
nand U1365 (N_1365,In_1935,In_2124);
and U1366 (N_1366,In_1575,In_1954);
or U1367 (N_1367,In_1041,In_1206);
and U1368 (N_1368,In_180,In_2005);
and U1369 (N_1369,In_1686,In_1269);
nor U1370 (N_1370,In_222,In_1316);
nand U1371 (N_1371,In_62,In_939);
nand U1372 (N_1372,In_328,In_2221);
or U1373 (N_1373,In_2329,In_1877);
nand U1374 (N_1374,In_1670,In_2042);
nor U1375 (N_1375,In_1222,In_1506);
and U1376 (N_1376,In_822,In_1538);
or U1377 (N_1377,In_567,In_962);
xor U1378 (N_1378,In_1646,In_1258);
nor U1379 (N_1379,In_101,In_1404);
or U1380 (N_1380,In_2068,In_1635);
nor U1381 (N_1381,In_24,In_248);
or U1382 (N_1382,In_306,In_2287);
xnor U1383 (N_1383,In_2021,In_875);
xor U1384 (N_1384,In_587,In_2491);
or U1385 (N_1385,In_1223,In_1815);
or U1386 (N_1386,In_1444,In_907);
and U1387 (N_1387,In_736,In_1946);
and U1388 (N_1388,In_348,In_279);
or U1389 (N_1389,In_1960,In_1399);
nor U1390 (N_1390,In_563,In_1139);
nand U1391 (N_1391,In_602,In_1467);
or U1392 (N_1392,In_1997,In_1715);
and U1393 (N_1393,In_2029,In_1676);
xor U1394 (N_1394,In_700,In_835);
and U1395 (N_1395,In_2028,In_1014);
nor U1396 (N_1396,In_2412,In_932);
or U1397 (N_1397,In_1326,In_720);
and U1398 (N_1398,In_650,In_979);
and U1399 (N_1399,In_110,In_1562);
or U1400 (N_1400,In_962,In_1706);
nand U1401 (N_1401,In_981,In_1809);
or U1402 (N_1402,In_1080,In_1581);
nor U1403 (N_1403,In_1095,In_2218);
nand U1404 (N_1404,In_655,In_1209);
or U1405 (N_1405,In_47,In_1127);
nand U1406 (N_1406,In_868,In_2263);
or U1407 (N_1407,In_1694,In_2262);
xor U1408 (N_1408,In_2467,In_723);
or U1409 (N_1409,In_916,In_1158);
or U1410 (N_1410,In_52,In_1371);
nand U1411 (N_1411,In_1826,In_2056);
xnor U1412 (N_1412,In_2283,In_414);
and U1413 (N_1413,In_1815,In_609);
and U1414 (N_1414,In_1600,In_1929);
nor U1415 (N_1415,In_1608,In_1192);
nor U1416 (N_1416,In_1912,In_119);
xnor U1417 (N_1417,In_1964,In_1357);
or U1418 (N_1418,In_2002,In_96);
and U1419 (N_1419,In_2086,In_877);
nand U1420 (N_1420,In_912,In_2208);
and U1421 (N_1421,In_784,In_1602);
and U1422 (N_1422,In_1841,In_911);
nand U1423 (N_1423,In_443,In_723);
nand U1424 (N_1424,In_1981,In_492);
nand U1425 (N_1425,In_1022,In_868);
nand U1426 (N_1426,In_1173,In_691);
or U1427 (N_1427,In_2102,In_2172);
nand U1428 (N_1428,In_1602,In_1390);
nor U1429 (N_1429,In_1896,In_2428);
and U1430 (N_1430,In_967,In_793);
or U1431 (N_1431,In_1888,In_201);
nor U1432 (N_1432,In_467,In_1763);
xor U1433 (N_1433,In_1412,In_1907);
xor U1434 (N_1434,In_2147,In_1499);
and U1435 (N_1435,In_2497,In_227);
nor U1436 (N_1436,In_58,In_1153);
and U1437 (N_1437,In_770,In_1608);
or U1438 (N_1438,In_836,In_1360);
and U1439 (N_1439,In_1168,In_1428);
or U1440 (N_1440,In_1234,In_180);
nand U1441 (N_1441,In_546,In_2194);
and U1442 (N_1442,In_1108,In_545);
and U1443 (N_1443,In_1569,In_1148);
and U1444 (N_1444,In_494,In_1883);
nor U1445 (N_1445,In_2307,In_40);
or U1446 (N_1446,In_1433,In_571);
nand U1447 (N_1447,In_1198,In_1595);
or U1448 (N_1448,In_244,In_572);
or U1449 (N_1449,In_334,In_1228);
nand U1450 (N_1450,In_2451,In_2351);
and U1451 (N_1451,In_1185,In_915);
nor U1452 (N_1452,In_1264,In_776);
or U1453 (N_1453,In_2300,In_2205);
and U1454 (N_1454,In_1312,In_244);
xor U1455 (N_1455,In_331,In_226);
nor U1456 (N_1456,In_1325,In_509);
nand U1457 (N_1457,In_21,In_2495);
or U1458 (N_1458,In_217,In_35);
nor U1459 (N_1459,In_342,In_730);
nand U1460 (N_1460,In_1280,In_272);
and U1461 (N_1461,In_618,In_1824);
xor U1462 (N_1462,In_865,In_671);
nor U1463 (N_1463,In_1189,In_166);
nor U1464 (N_1464,In_460,In_2211);
nor U1465 (N_1465,In_1900,In_944);
xnor U1466 (N_1466,In_1278,In_1731);
or U1467 (N_1467,In_1420,In_283);
xnor U1468 (N_1468,In_1790,In_2277);
nor U1469 (N_1469,In_452,In_1970);
and U1470 (N_1470,In_1168,In_1575);
nand U1471 (N_1471,In_490,In_2499);
nand U1472 (N_1472,In_358,In_737);
and U1473 (N_1473,In_497,In_2211);
or U1474 (N_1474,In_2063,In_2120);
or U1475 (N_1475,In_1982,In_1317);
nor U1476 (N_1476,In_70,In_1523);
and U1477 (N_1477,In_362,In_735);
nand U1478 (N_1478,In_1919,In_963);
or U1479 (N_1479,In_1152,In_1359);
or U1480 (N_1480,In_7,In_2442);
and U1481 (N_1481,In_329,In_506);
xor U1482 (N_1482,In_813,In_1899);
or U1483 (N_1483,In_115,In_1535);
or U1484 (N_1484,In_1112,In_1636);
nor U1485 (N_1485,In_2138,In_1533);
xnor U1486 (N_1486,In_203,In_1295);
or U1487 (N_1487,In_2326,In_1835);
nor U1488 (N_1488,In_1968,In_384);
and U1489 (N_1489,In_2166,In_1489);
xnor U1490 (N_1490,In_2158,In_2440);
and U1491 (N_1491,In_241,In_385);
nand U1492 (N_1492,In_2421,In_691);
and U1493 (N_1493,In_1283,In_1906);
nand U1494 (N_1494,In_813,In_1408);
xor U1495 (N_1495,In_1531,In_219);
xor U1496 (N_1496,In_2350,In_90);
nor U1497 (N_1497,In_1669,In_535);
xnor U1498 (N_1498,In_1377,In_245);
and U1499 (N_1499,In_1804,In_1032);
nand U1500 (N_1500,In_1122,In_363);
and U1501 (N_1501,In_1752,In_1615);
nor U1502 (N_1502,In_1843,In_2133);
and U1503 (N_1503,In_93,In_705);
nand U1504 (N_1504,In_1452,In_1991);
nand U1505 (N_1505,In_2,In_1923);
nand U1506 (N_1506,In_309,In_217);
nand U1507 (N_1507,In_1660,In_1250);
or U1508 (N_1508,In_197,In_2222);
nand U1509 (N_1509,In_17,In_788);
nor U1510 (N_1510,In_2025,In_1446);
nand U1511 (N_1511,In_2172,In_677);
and U1512 (N_1512,In_1730,In_419);
or U1513 (N_1513,In_621,In_632);
nand U1514 (N_1514,In_548,In_1414);
and U1515 (N_1515,In_146,In_33);
and U1516 (N_1516,In_2264,In_2181);
or U1517 (N_1517,In_2075,In_1987);
nor U1518 (N_1518,In_638,In_1779);
or U1519 (N_1519,In_881,In_688);
and U1520 (N_1520,In_118,In_269);
nor U1521 (N_1521,In_793,In_451);
and U1522 (N_1522,In_814,In_820);
and U1523 (N_1523,In_2363,In_2413);
nor U1524 (N_1524,In_254,In_2201);
and U1525 (N_1525,In_1910,In_2010);
or U1526 (N_1526,In_1273,In_53);
or U1527 (N_1527,In_1318,In_2417);
nand U1528 (N_1528,In_1068,In_484);
nor U1529 (N_1529,In_80,In_1819);
or U1530 (N_1530,In_1911,In_54);
nand U1531 (N_1531,In_1887,In_676);
and U1532 (N_1532,In_2191,In_1647);
or U1533 (N_1533,In_0,In_1165);
and U1534 (N_1534,In_336,In_1482);
nand U1535 (N_1535,In_2007,In_2337);
or U1536 (N_1536,In_932,In_2075);
nand U1537 (N_1537,In_464,In_511);
nor U1538 (N_1538,In_1657,In_1687);
nor U1539 (N_1539,In_1609,In_322);
nor U1540 (N_1540,In_917,In_1987);
and U1541 (N_1541,In_1067,In_1580);
nor U1542 (N_1542,In_1774,In_928);
and U1543 (N_1543,In_336,In_1963);
and U1544 (N_1544,In_1120,In_1705);
nor U1545 (N_1545,In_692,In_2351);
or U1546 (N_1546,In_1337,In_544);
or U1547 (N_1547,In_1176,In_511);
and U1548 (N_1548,In_1632,In_912);
or U1549 (N_1549,In_1539,In_266);
xor U1550 (N_1550,In_1496,In_1800);
nand U1551 (N_1551,In_267,In_1193);
xnor U1552 (N_1552,In_1286,In_403);
or U1553 (N_1553,In_1210,In_94);
xnor U1554 (N_1554,In_1270,In_384);
and U1555 (N_1555,In_2316,In_989);
nor U1556 (N_1556,In_272,In_1683);
or U1557 (N_1557,In_1592,In_1108);
nand U1558 (N_1558,In_2081,In_880);
nor U1559 (N_1559,In_2446,In_987);
xnor U1560 (N_1560,In_1627,In_2007);
or U1561 (N_1561,In_2347,In_204);
nand U1562 (N_1562,In_2474,In_2193);
and U1563 (N_1563,In_1696,In_2342);
nand U1564 (N_1564,In_430,In_823);
nand U1565 (N_1565,In_555,In_1148);
nand U1566 (N_1566,In_2118,In_480);
and U1567 (N_1567,In_2116,In_923);
nand U1568 (N_1568,In_737,In_339);
and U1569 (N_1569,In_2247,In_1559);
nand U1570 (N_1570,In_1701,In_574);
or U1571 (N_1571,In_104,In_1033);
nand U1572 (N_1572,In_1621,In_6);
nand U1573 (N_1573,In_1326,In_2073);
nor U1574 (N_1574,In_1926,In_1840);
and U1575 (N_1575,In_1035,In_1535);
nor U1576 (N_1576,In_2060,In_1562);
nor U1577 (N_1577,In_18,In_1547);
or U1578 (N_1578,In_252,In_1550);
or U1579 (N_1579,In_1945,In_64);
xnor U1580 (N_1580,In_78,In_1752);
or U1581 (N_1581,In_1894,In_1757);
xor U1582 (N_1582,In_1837,In_1057);
xnor U1583 (N_1583,In_646,In_1369);
nand U1584 (N_1584,In_1111,In_7);
and U1585 (N_1585,In_693,In_624);
and U1586 (N_1586,In_757,In_2323);
nand U1587 (N_1587,In_1374,In_1038);
or U1588 (N_1588,In_1278,In_877);
nor U1589 (N_1589,In_1718,In_2081);
and U1590 (N_1590,In_1344,In_329);
nand U1591 (N_1591,In_578,In_1724);
or U1592 (N_1592,In_930,In_438);
or U1593 (N_1593,In_672,In_1943);
nand U1594 (N_1594,In_2011,In_46);
xnor U1595 (N_1595,In_1464,In_1949);
nand U1596 (N_1596,In_239,In_1376);
xor U1597 (N_1597,In_192,In_2208);
and U1598 (N_1598,In_644,In_125);
or U1599 (N_1599,In_57,In_580);
and U1600 (N_1600,In_2451,In_294);
or U1601 (N_1601,In_1835,In_2244);
and U1602 (N_1602,In_377,In_2130);
nand U1603 (N_1603,In_1665,In_2108);
or U1604 (N_1604,In_610,In_863);
and U1605 (N_1605,In_844,In_778);
or U1606 (N_1606,In_2235,In_1776);
and U1607 (N_1607,In_1346,In_981);
nor U1608 (N_1608,In_2007,In_88);
or U1609 (N_1609,In_982,In_1440);
and U1610 (N_1610,In_2430,In_2187);
or U1611 (N_1611,In_538,In_953);
nor U1612 (N_1612,In_272,In_1525);
xor U1613 (N_1613,In_2128,In_1537);
nand U1614 (N_1614,In_1025,In_489);
or U1615 (N_1615,In_0,In_225);
nor U1616 (N_1616,In_642,In_438);
and U1617 (N_1617,In_2127,In_1499);
or U1618 (N_1618,In_2424,In_360);
nand U1619 (N_1619,In_849,In_1315);
or U1620 (N_1620,In_1426,In_80);
nor U1621 (N_1621,In_413,In_1692);
or U1622 (N_1622,In_246,In_20);
nand U1623 (N_1623,In_387,In_2105);
or U1624 (N_1624,In_1596,In_1330);
xnor U1625 (N_1625,In_386,In_163);
nor U1626 (N_1626,In_806,In_1295);
xnor U1627 (N_1627,In_2220,In_1680);
nand U1628 (N_1628,In_943,In_748);
nor U1629 (N_1629,In_2188,In_680);
xnor U1630 (N_1630,In_987,In_2182);
or U1631 (N_1631,In_748,In_335);
and U1632 (N_1632,In_262,In_14);
or U1633 (N_1633,In_1740,In_239);
or U1634 (N_1634,In_643,In_2418);
nor U1635 (N_1635,In_462,In_70);
xnor U1636 (N_1636,In_409,In_293);
xnor U1637 (N_1637,In_301,In_1141);
and U1638 (N_1638,In_85,In_124);
nor U1639 (N_1639,In_1114,In_32);
nand U1640 (N_1640,In_1303,In_1040);
or U1641 (N_1641,In_1938,In_648);
nor U1642 (N_1642,In_2265,In_853);
nor U1643 (N_1643,In_486,In_390);
or U1644 (N_1644,In_2345,In_978);
and U1645 (N_1645,In_1807,In_2269);
or U1646 (N_1646,In_121,In_2489);
and U1647 (N_1647,In_2110,In_824);
or U1648 (N_1648,In_2126,In_2440);
xnor U1649 (N_1649,In_647,In_2304);
xnor U1650 (N_1650,In_989,In_36);
nor U1651 (N_1651,In_180,In_114);
or U1652 (N_1652,In_2371,In_666);
or U1653 (N_1653,In_1116,In_720);
nand U1654 (N_1654,In_802,In_1874);
nand U1655 (N_1655,In_2097,In_411);
nand U1656 (N_1656,In_1965,In_1515);
and U1657 (N_1657,In_1731,In_863);
nand U1658 (N_1658,In_866,In_709);
and U1659 (N_1659,In_2269,In_2212);
nand U1660 (N_1660,In_1975,In_474);
or U1661 (N_1661,In_657,In_2159);
nand U1662 (N_1662,In_385,In_2128);
nand U1663 (N_1663,In_1979,In_490);
and U1664 (N_1664,In_152,In_2343);
or U1665 (N_1665,In_1335,In_713);
and U1666 (N_1666,In_996,In_138);
nor U1667 (N_1667,In_2152,In_1072);
or U1668 (N_1668,In_1752,In_1966);
or U1669 (N_1669,In_1038,In_1785);
or U1670 (N_1670,In_1181,In_427);
nor U1671 (N_1671,In_2047,In_1534);
and U1672 (N_1672,In_1546,In_227);
or U1673 (N_1673,In_1169,In_685);
xnor U1674 (N_1674,In_1417,In_1033);
xor U1675 (N_1675,In_394,In_369);
nand U1676 (N_1676,In_1261,In_154);
nand U1677 (N_1677,In_738,In_695);
or U1678 (N_1678,In_516,In_2454);
and U1679 (N_1679,In_1532,In_1197);
and U1680 (N_1680,In_2187,In_583);
or U1681 (N_1681,In_561,In_588);
or U1682 (N_1682,In_97,In_1728);
and U1683 (N_1683,In_1729,In_2388);
or U1684 (N_1684,In_919,In_2279);
and U1685 (N_1685,In_264,In_435);
and U1686 (N_1686,In_566,In_2013);
nor U1687 (N_1687,In_2183,In_2263);
nor U1688 (N_1688,In_613,In_600);
nand U1689 (N_1689,In_426,In_1017);
nor U1690 (N_1690,In_768,In_1577);
nor U1691 (N_1691,In_455,In_876);
nand U1692 (N_1692,In_967,In_156);
and U1693 (N_1693,In_2317,In_1757);
xor U1694 (N_1694,In_2303,In_158);
xnor U1695 (N_1695,In_1640,In_2414);
and U1696 (N_1696,In_2193,In_2426);
and U1697 (N_1697,In_2434,In_1969);
and U1698 (N_1698,In_113,In_1773);
and U1699 (N_1699,In_917,In_2030);
xnor U1700 (N_1700,In_2335,In_2118);
or U1701 (N_1701,In_325,In_630);
nand U1702 (N_1702,In_1810,In_1023);
nor U1703 (N_1703,In_1602,In_530);
and U1704 (N_1704,In_2183,In_543);
nor U1705 (N_1705,In_232,In_2405);
or U1706 (N_1706,In_2135,In_1511);
and U1707 (N_1707,In_1016,In_176);
and U1708 (N_1708,In_1802,In_1975);
or U1709 (N_1709,In_1640,In_1456);
or U1710 (N_1710,In_1072,In_1390);
nand U1711 (N_1711,In_1017,In_1995);
and U1712 (N_1712,In_2401,In_2051);
xnor U1713 (N_1713,In_1926,In_1986);
nand U1714 (N_1714,In_207,In_2451);
nor U1715 (N_1715,In_881,In_1258);
nand U1716 (N_1716,In_1714,In_2297);
and U1717 (N_1717,In_314,In_1716);
and U1718 (N_1718,In_2178,In_654);
nor U1719 (N_1719,In_2177,In_1683);
nand U1720 (N_1720,In_1497,In_806);
or U1721 (N_1721,In_1837,In_1595);
nor U1722 (N_1722,In_295,In_137);
or U1723 (N_1723,In_441,In_924);
nand U1724 (N_1724,In_1512,In_363);
and U1725 (N_1725,In_1701,In_133);
xor U1726 (N_1726,In_886,In_1511);
nand U1727 (N_1727,In_664,In_277);
nor U1728 (N_1728,In_175,In_2232);
nand U1729 (N_1729,In_1677,In_2116);
and U1730 (N_1730,In_326,In_16);
and U1731 (N_1731,In_2311,In_733);
nand U1732 (N_1732,In_639,In_1021);
nor U1733 (N_1733,In_422,In_1847);
nand U1734 (N_1734,In_1742,In_2162);
nor U1735 (N_1735,In_1859,In_862);
nor U1736 (N_1736,In_2471,In_415);
or U1737 (N_1737,In_1094,In_1420);
and U1738 (N_1738,In_146,In_1572);
nand U1739 (N_1739,In_18,In_270);
or U1740 (N_1740,In_330,In_2336);
and U1741 (N_1741,In_1316,In_2282);
or U1742 (N_1742,In_1518,In_1126);
nor U1743 (N_1743,In_1474,In_1748);
or U1744 (N_1744,In_962,In_1139);
nor U1745 (N_1745,In_1662,In_1850);
xor U1746 (N_1746,In_2040,In_858);
nor U1747 (N_1747,In_937,In_2232);
xor U1748 (N_1748,In_2362,In_360);
xor U1749 (N_1749,In_2117,In_1499);
or U1750 (N_1750,In_141,In_2062);
and U1751 (N_1751,In_1756,In_887);
and U1752 (N_1752,In_1950,In_1525);
nand U1753 (N_1753,In_201,In_1666);
or U1754 (N_1754,In_716,In_1448);
nand U1755 (N_1755,In_90,In_719);
nor U1756 (N_1756,In_1747,In_799);
or U1757 (N_1757,In_999,In_1611);
nand U1758 (N_1758,In_1528,In_1464);
and U1759 (N_1759,In_1826,In_502);
nand U1760 (N_1760,In_1445,In_1379);
nor U1761 (N_1761,In_2287,In_2459);
nand U1762 (N_1762,In_1174,In_1018);
xnor U1763 (N_1763,In_2272,In_832);
nand U1764 (N_1764,In_391,In_921);
nand U1765 (N_1765,In_626,In_586);
xnor U1766 (N_1766,In_357,In_2197);
nor U1767 (N_1767,In_994,In_843);
nor U1768 (N_1768,In_1049,In_1289);
xor U1769 (N_1769,In_1408,In_385);
nor U1770 (N_1770,In_428,In_1034);
nor U1771 (N_1771,In_2381,In_2297);
nor U1772 (N_1772,In_7,In_532);
nor U1773 (N_1773,In_863,In_2309);
or U1774 (N_1774,In_1545,In_1703);
or U1775 (N_1775,In_2432,In_140);
or U1776 (N_1776,In_1608,In_1147);
nor U1777 (N_1777,In_744,In_2341);
and U1778 (N_1778,In_2354,In_1889);
nand U1779 (N_1779,In_2360,In_73);
nand U1780 (N_1780,In_1951,In_2382);
and U1781 (N_1781,In_1793,In_2029);
and U1782 (N_1782,In_1248,In_1303);
or U1783 (N_1783,In_670,In_1623);
and U1784 (N_1784,In_1712,In_84);
and U1785 (N_1785,In_364,In_518);
xor U1786 (N_1786,In_550,In_543);
nand U1787 (N_1787,In_1430,In_1619);
nand U1788 (N_1788,In_1131,In_1017);
and U1789 (N_1789,In_2206,In_202);
or U1790 (N_1790,In_1570,In_1121);
or U1791 (N_1791,In_1209,In_826);
nor U1792 (N_1792,In_695,In_1880);
or U1793 (N_1793,In_1526,In_1706);
nand U1794 (N_1794,In_711,In_1404);
or U1795 (N_1795,In_2396,In_499);
or U1796 (N_1796,In_1087,In_469);
nand U1797 (N_1797,In_504,In_650);
and U1798 (N_1798,In_443,In_2345);
and U1799 (N_1799,In_810,In_723);
nand U1800 (N_1800,In_1702,In_571);
nand U1801 (N_1801,In_1798,In_2085);
and U1802 (N_1802,In_1839,In_2251);
xnor U1803 (N_1803,In_1979,In_971);
and U1804 (N_1804,In_1263,In_1599);
or U1805 (N_1805,In_1815,In_70);
nand U1806 (N_1806,In_1124,In_1990);
xnor U1807 (N_1807,In_2301,In_1459);
nand U1808 (N_1808,In_244,In_2299);
nor U1809 (N_1809,In_1961,In_1911);
xor U1810 (N_1810,In_567,In_263);
nor U1811 (N_1811,In_814,In_2477);
or U1812 (N_1812,In_1722,In_1898);
or U1813 (N_1813,In_1272,In_1021);
or U1814 (N_1814,In_1295,In_1345);
nor U1815 (N_1815,In_1326,In_1805);
nand U1816 (N_1816,In_94,In_2250);
nand U1817 (N_1817,In_2116,In_1477);
and U1818 (N_1818,In_1295,In_1545);
and U1819 (N_1819,In_392,In_2233);
nor U1820 (N_1820,In_1971,In_1927);
nand U1821 (N_1821,In_1795,In_2356);
or U1822 (N_1822,In_2143,In_2208);
and U1823 (N_1823,In_1792,In_1407);
nor U1824 (N_1824,In_2234,In_185);
or U1825 (N_1825,In_119,In_1766);
nor U1826 (N_1826,In_1983,In_981);
or U1827 (N_1827,In_82,In_507);
nand U1828 (N_1828,In_658,In_1599);
nor U1829 (N_1829,In_902,In_202);
and U1830 (N_1830,In_448,In_632);
or U1831 (N_1831,In_2497,In_2164);
nand U1832 (N_1832,In_521,In_585);
nand U1833 (N_1833,In_1951,In_634);
and U1834 (N_1834,In_1914,In_1101);
nand U1835 (N_1835,In_2393,In_784);
and U1836 (N_1836,In_2383,In_9);
and U1837 (N_1837,In_2177,In_674);
or U1838 (N_1838,In_345,In_1943);
or U1839 (N_1839,In_434,In_1317);
nand U1840 (N_1840,In_2422,In_2430);
nand U1841 (N_1841,In_1626,In_38);
nor U1842 (N_1842,In_577,In_2243);
or U1843 (N_1843,In_64,In_1490);
and U1844 (N_1844,In_215,In_1816);
and U1845 (N_1845,In_1643,In_1072);
and U1846 (N_1846,In_1408,In_418);
and U1847 (N_1847,In_149,In_1137);
nand U1848 (N_1848,In_1661,In_2283);
and U1849 (N_1849,In_1576,In_1640);
nor U1850 (N_1850,In_1920,In_2091);
nor U1851 (N_1851,In_1315,In_2212);
and U1852 (N_1852,In_301,In_1167);
or U1853 (N_1853,In_1655,In_1032);
or U1854 (N_1854,In_633,In_2378);
and U1855 (N_1855,In_1986,In_2174);
and U1856 (N_1856,In_2039,In_2375);
xnor U1857 (N_1857,In_226,In_525);
nor U1858 (N_1858,In_1351,In_2192);
xnor U1859 (N_1859,In_1353,In_1328);
or U1860 (N_1860,In_682,In_1882);
and U1861 (N_1861,In_2330,In_1487);
or U1862 (N_1862,In_780,In_1525);
nand U1863 (N_1863,In_1900,In_1251);
or U1864 (N_1864,In_1556,In_1279);
nor U1865 (N_1865,In_1804,In_2071);
and U1866 (N_1866,In_216,In_436);
nand U1867 (N_1867,In_1154,In_1774);
xor U1868 (N_1868,In_557,In_1163);
and U1869 (N_1869,In_480,In_183);
xor U1870 (N_1870,In_1453,In_1593);
and U1871 (N_1871,In_165,In_1656);
or U1872 (N_1872,In_1530,In_2261);
nand U1873 (N_1873,In_223,In_1178);
or U1874 (N_1874,In_919,In_168);
or U1875 (N_1875,In_2252,In_1664);
nand U1876 (N_1876,In_943,In_399);
nand U1877 (N_1877,In_2171,In_576);
nand U1878 (N_1878,In_1255,In_1827);
nor U1879 (N_1879,In_1593,In_2425);
nand U1880 (N_1880,In_1600,In_2272);
nor U1881 (N_1881,In_1038,In_1280);
nand U1882 (N_1882,In_895,In_347);
or U1883 (N_1883,In_1902,In_1750);
and U1884 (N_1884,In_350,In_2331);
nor U1885 (N_1885,In_2453,In_1045);
nand U1886 (N_1886,In_1221,In_1961);
and U1887 (N_1887,In_88,In_807);
nor U1888 (N_1888,In_1972,In_1769);
nor U1889 (N_1889,In_2440,In_910);
or U1890 (N_1890,In_950,In_717);
nor U1891 (N_1891,In_2013,In_1075);
xnor U1892 (N_1892,In_2365,In_801);
or U1893 (N_1893,In_57,In_239);
and U1894 (N_1894,In_109,In_1780);
or U1895 (N_1895,In_1931,In_2032);
or U1896 (N_1896,In_1041,In_115);
or U1897 (N_1897,In_1311,In_820);
or U1898 (N_1898,In_2241,In_1623);
or U1899 (N_1899,In_1986,In_1471);
or U1900 (N_1900,In_1934,In_225);
nor U1901 (N_1901,In_2254,In_146);
nor U1902 (N_1902,In_251,In_1269);
or U1903 (N_1903,In_1108,In_857);
nor U1904 (N_1904,In_1369,In_457);
nor U1905 (N_1905,In_1944,In_1448);
and U1906 (N_1906,In_1954,In_1866);
nand U1907 (N_1907,In_1028,In_345);
or U1908 (N_1908,In_1355,In_792);
nand U1909 (N_1909,In_992,In_921);
and U1910 (N_1910,In_71,In_645);
nand U1911 (N_1911,In_1878,In_1432);
and U1912 (N_1912,In_1066,In_2083);
and U1913 (N_1913,In_2000,In_2498);
and U1914 (N_1914,In_1084,In_1021);
or U1915 (N_1915,In_566,In_790);
or U1916 (N_1916,In_335,In_435);
or U1917 (N_1917,In_1271,In_2470);
xor U1918 (N_1918,In_1718,In_1484);
or U1919 (N_1919,In_1520,In_1031);
nand U1920 (N_1920,In_71,In_1826);
nor U1921 (N_1921,In_942,In_1738);
nand U1922 (N_1922,In_519,In_928);
or U1923 (N_1923,In_1406,In_767);
or U1924 (N_1924,In_1177,In_2109);
or U1925 (N_1925,In_1348,In_1478);
and U1926 (N_1926,In_207,In_1554);
or U1927 (N_1927,In_623,In_1192);
nand U1928 (N_1928,In_766,In_455);
or U1929 (N_1929,In_669,In_2447);
nand U1930 (N_1930,In_1591,In_580);
nand U1931 (N_1931,In_2450,In_2439);
nor U1932 (N_1932,In_894,In_656);
xnor U1933 (N_1933,In_20,In_672);
and U1934 (N_1934,In_782,In_787);
and U1935 (N_1935,In_111,In_1052);
nand U1936 (N_1936,In_1592,In_704);
and U1937 (N_1937,In_343,In_2171);
nor U1938 (N_1938,In_1533,In_2032);
or U1939 (N_1939,In_1304,In_940);
nor U1940 (N_1940,In_1406,In_726);
and U1941 (N_1941,In_186,In_572);
and U1942 (N_1942,In_2130,In_554);
nor U1943 (N_1943,In_1383,In_747);
nor U1944 (N_1944,In_2161,In_2430);
and U1945 (N_1945,In_1542,In_2024);
nand U1946 (N_1946,In_2119,In_1506);
nand U1947 (N_1947,In_1487,In_880);
nand U1948 (N_1948,In_2181,In_2419);
and U1949 (N_1949,In_1884,In_1333);
and U1950 (N_1950,In_2498,In_1123);
nor U1951 (N_1951,In_1342,In_1336);
or U1952 (N_1952,In_338,In_125);
and U1953 (N_1953,In_529,In_1522);
nand U1954 (N_1954,In_1009,In_1416);
or U1955 (N_1955,In_344,In_988);
xnor U1956 (N_1956,In_612,In_847);
or U1957 (N_1957,In_1323,In_1919);
and U1958 (N_1958,In_1549,In_1741);
nand U1959 (N_1959,In_1254,In_953);
nand U1960 (N_1960,In_950,In_1143);
and U1961 (N_1961,In_864,In_1079);
nand U1962 (N_1962,In_877,In_2425);
nand U1963 (N_1963,In_2371,In_960);
nor U1964 (N_1964,In_2192,In_1124);
and U1965 (N_1965,In_2254,In_116);
or U1966 (N_1966,In_2108,In_1228);
and U1967 (N_1967,In_1526,In_1222);
and U1968 (N_1968,In_785,In_1367);
or U1969 (N_1969,In_587,In_1991);
and U1970 (N_1970,In_332,In_2061);
and U1971 (N_1971,In_1009,In_848);
and U1972 (N_1972,In_209,In_1686);
or U1973 (N_1973,In_1660,In_1504);
and U1974 (N_1974,In_451,In_2249);
nor U1975 (N_1975,In_750,In_1166);
nand U1976 (N_1976,In_605,In_1419);
xnor U1977 (N_1977,In_334,In_1469);
nor U1978 (N_1978,In_1592,In_728);
nand U1979 (N_1979,In_53,In_363);
and U1980 (N_1980,In_198,In_2388);
nand U1981 (N_1981,In_1271,In_872);
and U1982 (N_1982,In_87,In_922);
nor U1983 (N_1983,In_2285,In_2112);
nand U1984 (N_1984,In_2196,In_2337);
nor U1985 (N_1985,In_2344,In_1368);
or U1986 (N_1986,In_69,In_2494);
nor U1987 (N_1987,In_2117,In_2015);
and U1988 (N_1988,In_2196,In_528);
nor U1989 (N_1989,In_2034,In_1638);
and U1990 (N_1990,In_2444,In_454);
nor U1991 (N_1991,In_707,In_1203);
or U1992 (N_1992,In_885,In_856);
xor U1993 (N_1993,In_845,In_1463);
or U1994 (N_1994,In_721,In_1840);
nor U1995 (N_1995,In_1456,In_1510);
or U1996 (N_1996,In_1304,In_822);
nor U1997 (N_1997,In_1674,In_1987);
nand U1998 (N_1998,In_1062,In_2290);
nand U1999 (N_1999,In_1909,In_183);
or U2000 (N_2000,In_1281,In_2357);
or U2001 (N_2001,In_2143,In_1546);
nor U2002 (N_2002,In_1934,In_2222);
nor U2003 (N_2003,In_1812,In_384);
nor U2004 (N_2004,In_1017,In_1529);
and U2005 (N_2005,In_256,In_583);
xor U2006 (N_2006,In_2266,In_1177);
and U2007 (N_2007,In_214,In_1881);
or U2008 (N_2008,In_1548,In_1901);
xnor U2009 (N_2009,In_1105,In_798);
nand U2010 (N_2010,In_358,In_1662);
xnor U2011 (N_2011,In_254,In_540);
nor U2012 (N_2012,In_1689,In_792);
xor U2013 (N_2013,In_130,In_1185);
and U2014 (N_2014,In_2353,In_522);
nor U2015 (N_2015,In_1772,In_583);
or U2016 (N_2016,In_440,In_1819);
and U2017 (N_2017,In_1570,In_54);
xnor U2018 (N_2018,In_1805,In_1672);
or U2019 (N_2019,In_1995,In_1892);
nand U2020 (N_2020,In_479,In_432);
nand U2021 (N_2021,In_41,In_1372);
and U2022 (N_2022,In_1553,In_639);
xor U2023 (N_2023,In_2267,In_837);
and U2024 (N_2024,In_530,In_828);
nand U2025 (N_2025,In_807,In_399);
nand U2026 (N_2026,In_1597,In_1366);
nand U2027 (N_2027,In_2201,In_205);
nor U2028 (N_2028,In_1852,In_1986);
nor U2029 (N_2029,In_35,In_337);
and U2030 (N_2030,In_1440,In_774);
or U2031 (N_2031,In_1341,In_782);
nand U2032 (N_2032,In_1064,In_524);
xor U2033 (N_2033,In_581,In_1404);
and U2034 (N_2034,In_424,In_1151);
nor U2035 (N_2035,In_877,In_1352);
and U2036 (N_2036,In_261,In_1480);
or U2037 (N_2037,In_494,In_631);
or U2038 (N_2038,In_2456,In_2346);
xnor U2039 (N_2039,In_161,In_619);
nand U2040 (N_2040,In_1141,In_2485);
nor U2041 (N_2041,In_1154,In_1189);
nand U2042 (N_2042,In_1982,In_1540);
nor U2043 (N_2043,In_99,In_491);
xnor U2044 (N_2044,In_947,In_1531);
and U2045 (N_2045,In_137,In_1046);
xor U2046 (N_2046,In_1076,In_1035);
or U2047 (N_2047,In_972,In_2241);
and U2048 (N_2048,In_1334,In_1911);
or U2049 (N_2049,In_153,In_851);
nand U2050 (N_2050,In_2440,In_2315);
and U2051 (N_2051,In_804,In_294);
nor U2052 (N_2052,In_466,In_1833);
or U2053 (N_2053,In_183,In_744);
or U2054 (N_2054,In_2193,In_1024);
nand U2055 (N_2055,In_903,In_456);
nand U2056 (N_2056,In_351,In_2493);
xor U2057 (N_2057,In_605,In_2345);
nor U2058 (N_2058,In_1017,In_321);
or U2059 (N_2059,In_1427,In_1550);
nor U2060 (N_2060,In_443,In_115);
nor U2061 (N_2061,In_1209,In_609);
or U2062 (N_2062,In_1681,In_176);
nand U2063 (N_2063,In_270,In_379);
nor U2064 (N_2064,In_103,In_1146);
nand U2065 (N_2065,In_2389,In_726);
nor U2066 (N_2066,In_966,In_1909);
nand U2067 (N_2067,In_2109,In_492);
or U2068 (N_2068,In_691,In_187);
and U2069 (N_2069,In_1565,In_11);
nor U2070 (N_2070,In_2439,In_1458);
and U2071 (N_2071,In_1804,In_95);
xnor U2072 (N_2072,In_1376,In_1107);
nor U2073 (N_2073,In_248,In_1984);
and U2074 (N_2074,In_1304,In_1958);
nor U2075 (N_2075,In_1573,In_1044);
nor U2076 (N_2076,In_663,In_287);
xor U2077 (N_2077,In_1105,In_2223);
and U2078 (N_2078,In_1961,In_1340);
or U2079 (N_2079,In_804,In_1963);
nand U2080 (N_2080,In_1922,In_1309);
or U2081 (N_2081,In_1433,In_592);
xor U2082 (N_2082,In_677,In_992);
and U2083 (N_2083,In_932,In_1386);
nor U2084 (N_2084,In_2457,In_958);
and U2085 (N_2085,In_2059,In_2035);
and U2086 (N_2086,In_2278,In_216);
or U2087 (N_2087,In_694,In_788);
and U2088 (N_2088,In_1589,In_1662);
and U2089 (N_2089,In_2187,In_2418);
nand U2090 (N_2090,In_513,In_1731);
xor U2091 (N_2091,In_1651,In_1298);
nand U2092 (N_2092,In_685,In_544);
and U2093 (N_2093,In_1336,In_2156);
nor U2094 (N_2094,In_559,In_1751);
or U2095 (N_2095,In_686,In_2096);
nor U2096 (N_2096,In_831,In_809);
nand U2097 (N_2097,In_110,In_265);
nand U2098 (N_2098,In_158,In_2333);
or U2099 (N_2099,In_1238,In_324);
xnor U2100 (N_2100,In_380,In_2489);
nor U2101 (N_2101,In_813,In_486);
nand U2102 (N_2102,In_185,In_153);
and U2103 (N_2103,In_1577,In_2157);
and U2104 (N_2104,In_895,In_1863);
xnor U2105 (N_2105,In_321,In_1430);
nor U2106 (N_2106,In_2109,In_1067);
nand U2107 (N_2107,In_2213,In_1589);
nor U2108 (N_2108,In_51,In_1387);
nor U2109 (N_2109,In_833,In_1099);
and U2110 (N_2110,In_1791,In_1725);
nor U2111 (N_2111,In_981,In_1583);
or U2112 (N_2112,In_1307,In_727);
and U2113 (N_2113,In_54,In_1049);
and U2114 (N_2114,In_35,In_1407);
nor U2115 (N_2115,In_12,In_1224);
or U2116 (N_2116,In_1731,In_982);
and U2117 (N_2117,In_1963,In_1010);
and U2118 (N_2118,In_1222,In_673);
or U2119 (N_2119,In_480,In_2070);
nor U2120 (N_2120,In_1879,In_1534);
nor U2121 (N_2121,In_2463,In_1465);
nand U2122 (N_2122,In_112,In_1771);
xnor U2123 (N_2123,In_639,In_1492);
and U2124 (N_2124,In_941,In_461);
nor U2125 (N_2125,In_563,In_915);
nor U2126 (N_2126,In_981,In_685);
and U2127 (N_2127,In_942,In_1519);
and U2128 (N_2128,In_277,In_1546);
xor U2129 (N_2129,In_1543,In_584);
nand U2130 (N_2130,In_2201,In_36);
xor U2131 (N_2131,In_1103,In_282);
and U2132 (N_2132,In_446,In_1408);
and U2133 (N_2133,In_616,In_1033);
or U2134 (N_2134,In_725,In_1617);
nand U2135 (N_2135,In_1038,In_2350);
xnor U2136 (N_2136,In_2362,In_651);
nand U2137 (N_2137,In_1925,In_558);
and U2138 (N_2138,In_1611,In_502);
nand U2139 (N_2139,In_1562,In_2418);
or U2140 (N_2140,In_1196,In_135);
xnor U2141 (N_2141,In_1848,In_792);
and U2142 (N_2142,In_108,In_1074);
or U2143 (N_2143,In_970,In_1089);
nor U2144 (N_2144,In_1959,In_2425);
nand U2145 (N_2145,In_1691,In_1887);
xnor U2146 (N_2146,In_582,In_1335);
or U2147 (N_2147,In_258,In_131);
and U2148 (N_2148,In_2296,In_2063);
or U2149 (N_2149,In_1795,In_559);
or U2150 (N_2150,In_2260,In_1694);
or U2151 (N_2151,In_678,In_2098);
xor U2152 (N_2152,In_1838,In_1463);
nor U2153 (N_2153,In_975,In_291);
or U2154 (N_2154,In_2452,In_378);
nand U2155 (N_2155,In_2435,In_621);
and U2156 (N_2156,In_2414,In_104);
xnor U2157 (N_2157,In_1113,In_1728);
nand U2158 (N_2158,In_405,In_1651);
nor U2159 (N_2159,In_1903,In_1291);
nor U2160 (N_2160,In_1322,In_1299);
and U2161 (N_2161,In_353,In_1096);
nor U2162 (N_2162,In_1049,In_1061);
nand U2163 (N_2163,In_1384,In_1047);
nor U2164 (N_2164,In_1751,In_391);
or U2165 (N_2165,In_318,In_1900);
nor U2166 (N_2166,In_956,In_685);
and U2167 (N_2167,In_1390,In_1243);
nand U2168 (N_2168,In_1187,In_2424);
or U2169 (N_2169,In_696,In_829);
nand U2170 (N_2170,In_214,In_2360);
and U2171 (N_2171,In_1606,In_1474);
or U2172 (N_2172,In_409,In_1629);
nor U2173 (N_2173,In_925,In_1344);
or U2174 (N_2174,In_1022,In_430);
nor U2175 (N_2175,In_1459,In_369);
nand U2176 (N_2176,In_705,In_780);
and U2177 (N_2177,In_1140,In_2450);
or U2178 (N_2178,In_2395,In_809);
nand U2179 (N_2179,In_1611,In_1356);
or U2180 (N_2180,In_565,In_1338);
nand U2181 (N_2181,In_1022,In_1895);
and U2182 (N_2182,In_1054,In_893);
nand U2183 (N_2183,In_421,In_975);
nor U2184 (N_2184,In_1333,In_19);
xnor U2185 (N_2185,In_266,In_413);
nand U2186 (N_2186,In_799,In_338);
nand U2187 (N_2187,In_600,In_119);
nor U2188 (N_2188,In_857,In_800);
nand U2189 (N_2189,In_1976,In_232);
xor U2190 (N_2190,In_906,In_1808);
and U2191 (N_2191,In_945,In_419);
or U2192 (N_2192,In_1002,In_2226);
and U2193 (N_2193,In_1250,In_616);
nand U2194 (N_2194,In_876,In_1364);
xnor U2195 (N_2195,In_767,In_506);
nor U2196 (N_2196,In_242,In_2372);
nor U2197 (N_2197,In_603,In_1351);
nand U2198 (N_2198,In_1050,In_2021);
or U2199 (N_2199,In_2486,In_1182);
or U2200 (N_2200,In_1116,In_151);
or U2201 (N_2201,In_41,In_2489);
nand U2202 (N_2202,In_1772,In_1340);
xor U2203 (N_2203,In_411,In_637);
or U2204 (N_2204,In_409,In_2264);
or U2205 (N_2205,In_1696,In_1712);
nand U2206 (N_2206,In_2189,In_1350);
nor U2207 (N_2207,In_1993,In_56);
nor U2208 (N_2208,In_1527,In_1378);
nor U2209 (N_2209,In_1401,In_1479);
or U2210 (N_2210,In_516,In_260);
and U2211 (N_2211,In_2385,In_642);
and U2212 (N_2212,In_1694,In_1661);
nor U2213 (N_2213,In_2072,In_412);
or U2214 (N_2214,In_2451,In_2266);
nand U2215 (N_2215,In_1478,In_2152);
nand U2216 (N_2216,In_1029,In_2331);
xor U2217 (N_2217,In_590,In_2453);
and U2218 (N_2218,In_463,In_1793);
nor U2219 (N_2219,In_480,In_518);
or U2220 (N_2220,In_286,In_2213);
nor U2221 (N_2221,In_510,In_2106);
and U2222 (N_2222,In_1345,In_1689);
and U2223 (N_2223,In_74,In_2005);
nand U2224 (N_2224,In_2335,In_1549);
and U2225 (N_2225,In_1883,In_980);
and U2226 (N_2226,In_2110,In_1625);
or U2227 (N_2227,In_284,In_324);
and U2228 (N_2228,In_412,In_1304);
and U2229 (N_2229,In_564,In_1621);
nand U2230 (N_2230,In_660,In_229);
nor U2231 (N_2231,In_1709,In_2150);
or U2232 (N_2232,In_1701,In_1790);
nand U2233 (N_2233,In_199,In_996);
nor U2234 (N_2234,In_2045,In_2138);
and U2235 (N_2235,In_1689,In_2122);
nand U2236 (N_2236,In_1053,In_2216);
nand U2237 (N_2237,In_215,In_621);
xnor U2238 (N_2238,In_2310,In_1780);
nor U2239 (N_2239,In_469,In_1855);
or U2240 (N_2240,In_309,In_1363);
and U2241 (N_2241,In_2193,In_218);
or U2242 (N_2242,In_933,In_2401);
nand U2243 (N_2243,In_257,In_2193);
xnor U2244 (N_2244,In_448,In_2145);
or U2245 (N_2245,In_2409,In_953);
nand U2246 (N_2246,In_1990,In_2020);
nand U2247 (N_2247,In_923,In_355);
and U2248 (N_2248,In_641,In_476);
nand U2249 (N_2249,In_2257,In_1340);
nand U2250 (N_2250,In_2403,In_2100);
nand U2251 (N_2251,In_1596,In_616);
nor U2252 (N_2252,In_1997,In_413);
or U2253 (N_2253,In_368,In_1987);
nor U2254 (N_2254,In_2360,In_1937);
nand U2255 (N_2255,In_934,In_2362);
nor U2256 (N_2256,In_810,In_866);
nand U2257 (N_2257,In_765,In_1965);
nand U2258 (N_2258,In_1350,In_2091);
or U2259 (N_2259,In_2130,In_2105);
nand U2260 (N_2260,In_1614,In_174);
nand U2261 (N_2261,In_2428,In_1941);
or U2262 (N_2262,In_137,In_206);
and U2263 (N_2263,In_389,In_499);
and U2264 (N_2264,In_1594,In_2051);
or U2265 (N_2265,In_2354,In_493);
or U2266 (N_2266,In_1241,In_409);
nor U2267 (N_2267,In_1294,In_838);
nor U2268 (N_2268,In_2133,In_2228);
nor U2269 (N_2269,In_2151,In_827);
and U2270 (N_2270,In_1440,In_903);
and U2271 (N_2271,In_1017,In_787);
and U2272 (N_2272,In_2464,In_2032);
nor U2273 (N_2273,In_990,In_521);
and U2274 (N_2274,In_2315,In_1956);
and U2275 (N_2275,In_959,In_1717);
nor U2276 (N_2276,In_2057,In_967);
or U2277 (N_2277,In_917,In_2338);
nor U2278 (N_2278,In_56,In_1446);
nor U2279 (N_2279,In_371,In_1739);
and U2280 (N_2280,In_261,In_520);
nor U2281 (N_2281,In_970,In_2285);
and U2282 (N_2282,In_1217,In_1901);
or U2283 (N_2283,In_1861,In_2350);
or U2284 (N_2284,In_1827,In_51);
nand U2285 (N_2285,In_629,In_2258);
and U2286 (N_2286,In_2122,In_2303);
or U2287 (N_2287,In_1035,In_601);
xor U2288 (N_2288,In_334,In_911);
or U2289 (N_2289,In_1731,In_2071);
or U2290 (N_2290,In_594,In_1753);
or U2291 (N_2291,In_2376,In_1819);
nor U2292 (N_2292,In_2368,In_260);
nor U2293 (N_2293,In_1905,In_1294);
or U2294 (N_2294,In_679,In_2319);
and U2295 (N_2295,In_1230,In_2254);
nand U2296 (N_2296,In_114,In_1742);
nand U2297 (N_2297,In_905,In_1990);
or U2298 (N_2298,In_559,In_2468);
and U2299 (N_2299,In_2419,In_2176);
nand U2300 (N_2300,In_1978,In_1968);
or U2301 (N_2301,In_1439,In_997);
and U2302 (N_2302,In_248,In_1081);
or U2303 (N_2303,In_958,In_1059);
or U2304 (N_2304,In_1981,In_479);
and U2305 (N_2305,In_1358,In_160);
nand U2306 (N_2306,In_2111,In_816);
nor U2307 (N_2307,In_2479,In_1787);
nand U2308 (N_2308,In_1430,In_881);
nor U2309 (N_2309,In_1502,In_93);
or U2310 (N_2310,In_1318,In_2410);
xor U2311 (N_2311,In_2087,In_587);
nor U2312 (N_2312,In_1728,In_1215);
xor U2313 (N_2313,In_1447,In_2326);
xor U2314 (N_2314,In_2329,In_1884);
or U2315 (N_2315,In_148,In_1244);
and U2316 (N_2316,In_1676,In_1754);
xor U2317 (N_2317,In_497,In_1870);
or U2318 (N_2318,In_96,In_1498);
nor U2319 (N_2319,In_342,In_1266);
or U2320 (N_2320,In_253,In_299);
nor U2321 (N_2321,In_1835,In_951);
or U2322 (N_2322,In_581,In_1276);
nor U2323 (N_2323,In_392,In_2372);
nor U2324 (N_2324,In_2063,In_318);
or U2325 (N_2325,In_666,In_1099);
and U2326 (N_2326,In_1339,In_813);
xor U2327 (N_2327,In_1431,In_1503);
and U2328 (N_2328,In_276,In_829);
or U2329 (N_2329,In_1263,In_2061);
and U2330 (N_2330,In_1166,In_2102);
nor U2331 (N_2331,In_546,In_56);
and U2332 (N_2332,In_1699,In_572);
and U2333 (N_2333,In_507,In_932);
and U2334 (N_2334,In_1513,In_865);
or U2335 (N_2335,In_87,In_1391);
nand U2336 (N_2336,In_1985,In_1417);
nor U2337 (N_2337,In_1095,In_940);
xnor U2338 (N_2338,In_1990,In_1696);
or U2339 (N_2339,In_1508,In_2057);
or U2340 (N_2340,In_1409,In_1160);
xnor U2341 (N_2341,In_213,In_2124);
and U2342 (N_2342,In_2332,In_1379);
nand U2343 (N_2343,In_627,In_2365);
xor U2344 (N_2344,In_550,In_567);
nor U2345 (N_2345,In_702,In_1446);
nand U2346 (N_2346,In_791,In_48);
xor U2347 (N_2347,In_65,In_33);
nand U2348 (N_2348,In_1344,In_2442);
nand U2349 (N_2349,In_1652,In_1407);
or U2350 (N_2350,In_974,In_2386);
nand U2351 (N_2351,In_540,In_1694);
nand U2352 (N_2352,In_1717,In_1931);
nand U2353 (N_2353,In_1348,In_1342);
nor U2354 (N_2354,In_478,In_1263);
xnor U2355 (N_2355,In_865,In_1063);
nor U2356 (N_2356,In_1151,In_830);
xor U2357 (N_2357,In_437,In_2335);
nand U2358 (N_2358,In_1761,In_580);
and U2359 (N_2359,In_1529,In_70);
or U2360 (N_2360,In_1912,In_1710);
or U2361 (N_2361,In_281,In_1793);
nand U2362 (N_2362,In_1244,In_2417);
nand U2363 (N_2363,In_1804,In_1132);
or U2364 (N_2364,In_2270,In_159);
xnor U2365 (N_2365,In_1357,In_1472);
nor U2366 (N_2366,In_2296,In_171);
xnor U2367 (N_2367,In_1260,In_1507);
nor U2368 (N_2368,In_443,In_436);
or U2369 (N_2369,In_879,In_1779);
nor U2370 (N_2370,In_1070,In_1055);
nand U2371 (N_2371,In_2491,In_540);
nand U2372 (N_2372,In_1385,In_288);
or U2373 (N_2373,In_2067,In_836);
xnor U2374 (N_2374,In_1326,In_1976);
and U2375 (N_2375,In_1904,In_99);
or U2376 (N_2376,In_1384,In_1521);
or U2377 (N_2377,In_193,In_1792);
nand U2378 (N_2378,In_1966,In_1701);
or U2379 (N_2379,In_1935,In_887);
nand U2380 (N_2380,In_1767,In_364);
nor U2381 (N_2381,In_938,In_1771);
and U2382 (N_2382,In_2100,In_2116);
xnor U2383 (N_2383,In_1880,In_1649);
xnor U2384 (N_2384,In_196,In_428);
and U2385 (N_2385,In_1231,In_1918);
nand U2386 (N_2386,In_1959,In_1201);
nand U2387 (N_2387,In_2286,In_1245);
nand U2388 (N_2388,In_1158,In_299);
and U2389 (N_2389,In_1178,In_2245);
and U2390 (N_2390,In_1288,In_2103);
and U2391 (N_2391,In_1425,In_514);
and U2392 (N_2392,In_1616,In_2277);
nor U2393 (N_2393,In_1581,In_2019);
xor U2394 (N_2394,In_996,In_651);
xor U2395 (N_2395,In_2297,In_856);
and U2396 (N_2396,In_1568,In_189);
and U2397 (N_2397,In_1452,In_425);
and U2398 (N_2398,In_1242,In_632);
nand U2399 (N_2399,In_2219,In_1721);
and U2400 (N_2400,In_1141,In_2121);
or U2401 (N_2401,In_131,In_898);
or U2402 (N_2402,In_1002,In_627);
and U2403 (N_2403,In_1097,In_1366);
nor U2404 (N_2404,In_461,In_841);
nand U2405 (N_2405,In_1070,In_246);
or U2406 (N_2406,In_535,In_794);
nand U2407 (N_2407,In_1379,In_1823);
and U2408 (N_2408,In_1794,In_876);
and U2409 (N_2409,In_1852,In_2150);
nand U2410 (N_2410,In_279,In_2188);
and U2411 (N_2411,In_2371,In_350);
and U2412 (N_2412,In_496,In_929);
nand U2413 (N_2413,In_983,In_1048);
nor U2414 (N_2414,In_707,In_1362);
or U2415 (N_2415,In_884,In_357);
nor U2416 (N_2416,In_2425,In_1829);
nand U2417 (N_2417,In_1230,In_2211);
nand U2418 (N_2418,In_1205,In_1161);
and U2419 (N_2419,In_1259,In_581);
nand U2420 (N_2420,In_2434,In_595);
nor U2421 (N_2421,In_1347,In_924);
and U2422 (N_2422,In_1615,In_152);
and U2423 (N_2423,In_944,In_1993);
or U2424 (N_2424,In_617,In_2406);
xor U2425 (N_2425,In_2148,In_2098);
or U2426 (N_2426,In_419,In_505);
or U2427 (N_2427,In_1402,In_1844);
or U2428 (N_2428,In_2057,In_424);
or U2429 (N_2429,In_1845,In_1853);
or U2430 (N_2430,In_2344,In_1881);
nand U2431 (N_2431,In_645,In_666);
nor U2432 (N_2432,In_1946,In_433);
or U2433 (N_2433,In_2479,In_994);
and U2434 (N_2434,In_2251,In_1005);
nand U2435 (N_2435,In_326,In_2427);
nand U2436 (N_2436,In_698,In_1717);
and U2437 (N_2437,In_1887,In_1298);
and U2438 (N_2438,In_1155,In_2393);
nor U2439 (N_2439,In_139,In_1475);
nor U2440 (N_2440,In_2364,In_1850);
nor U2441 (N_2441,In_2497,In_194);
and U2442 (N_2442,In_822,In_1378);
and U2443 (N_2443,In_1849,In_2497);
and U2444 (N_2444,In_1312,In_821);
nor U2445 (N_2445,In_1154,In_1538);
and U2446 (N_2446,In_1465,In_2461);
and U2447 (N_2447,In_2118,In_739);
and U2448 (N_2448,In_1896,In_1199);
and U2449 (N_2449,In_544,In_1468);
and U2450 (N_2450,In_1841,In_657);
nand U2451 (N_2451,In_270,In_2466);
nor U2452 (N_2452,In_1461,In_950);
nor U2453 (N_2453,In_961,In_1800);
nand U2454 (N_2454,In_926,In_1367);
nand U2455 (N_2455,In_1628,In_666);
nand U2456 (N_2456,In_978,In_523);
nor U2457 (N_2457,In_1263,In_724);
nor U2458 (N_2458,In_841,In_2125);
or U2459 (N_2459,In_2441,In_1209);
xor U2460 (N_2460,In_2451,In_2160);
or U2461 (N_2461,In_580,In_2036);
nor U2462 (N_2462,In_1550,In_1817);
or U2463 (N_2463,In_2441,In_2460);
nor U2464 (N_2464,In_755,In_478);
or U2465 (N_2465,In_963,In_599);
nand U2466 (N_2466,In_2303,In_224);
and U2467 (N_2467,In_1895,In_1502);
nor U2468 (N_2468,In_2389,In_1023);
and U2469 (N_2469,In_551,In_268);
nor U2470 (N_2470,In_179,In_512);
or U2471 (N_2471,In_1808,In_1683);
and U2472 (N_2472,In_373,In_1781);
nand U2473 (N_2473,In_408,In_1990);
or U2474 (N_2474,In_1186,In_1953);
and U2475 (N_2475,In_358,In_755);
nor U2476 (N_2476,In_1676,In_1892);
nor U2477 (N_2477,In_2045,In_2355);
or U2478 (N_2478,In_417,In_1677);
and U2479 (N_2479,In_1476,In_740);
or U2480 (N_2480,In_2224,In_831);
nor U2481 (N_2481,In_261,In_104);
nor U2482 (N_2482,In_1861,In_285);
nand U2483 (N_2483,In_1434,In_1400);
nand U2484 (N_2484,In_2226,In_2061);
and U2485 (N_2485,In_159,In_1917);
xor U2486 (N_2486,In_1333,In_2022);
or U2487 (N_2487,In_608,In_1580);
nand U2488 (N_2488,In_1470,In_1471);
and U2489 (N_2489,In_2121,In_1580);
nor U2490 (N_2490,In_1981,In_1294);
nand U2491 (N_2491,In_382,In_1655);
or U2492 (N_2492,In_2020,In_871);
and U2493 (N_2493,In_672,In_255);
and U2494 (N_2494,In_2463,In_1444);
nand U2495 (N_2495,In_104,In_1787);
nor U2496 (N_2496,In_577,In_2149);
or U2497 (N_2497,In_1306,In_1851);
nand U2498 (N_2498,In_2016,In_892);
xnor U2499 (N_2499,In_977,In_573);
nor U2500 (N_2500,In_1682,In_387);
nand U2501 (N_2501,In_823,In_983);
nand U2502 (N_2502,In_512,In_2039);
and U2503 (N_2503,In_1486,In_1656);
nor U2504 (N_2504,In_2043,In_907);
and U2505 (N_2505,In_100,In_226);
nor U2506 (N_2506,In_839,In_416);
or U2507 (N_2507,In_1467,In_2059);
and U2508 (N_2508,In_1746,In_273);
or U2509 (N_2509,In_1352,In_2422);
and U2510 (N_2510,In_1005,In_1576);
xor U2511 (N_2511,In_2363,In_1347);
or U2512 (N_2512,In_378,In_1679);
or U2513 (N_2513,In_103,In_1762);
nor U2514 (N_2514,In_1737,In_2163);
nand U2515 (N_2515,In_1704,In_269);
and U2516 (N_2516,In_837,In_90);
or U2517 (N_2517,In_2314,In_95);
and U2518 (N_2518,In_2463,In_65);
or U2519 (N_2519,In_1179,In_1648);
or U2520 (N_2520,In_1426,In_829);
nand U2521 (N_2521,In_111,In_1400);
nor U2522 (N_2522,In_652,In_1528);
nor U2523 (N_2523,In_2000,In_163);
nor U2524 (N_2524,In_981,In_980);
xor U2525 (N_2525,In_3,In_897);
or U2526 (N_2526,In_1808,In_1976);
or U2527 (N_2527,In_270,In_2233);
or U2528 (N_2528,In_1487,In_1009);
xnor U2529 (N_2529,In_385,In_1764);
nor U2530 (N_2530,In_643,In_554);
nand U2531 (N_2531,In_1194,In_1971);
or U2532 (N_2532,In_2289,In_2434);
nand U2533 (N_2533,In_90,In_1383);
or U2534 (N_2534,In_1831,In_1567);
or U2535 (N_2535,In_870,In_1034);
or U2536 (N_2536,In_1888,In_2252);
and U2537 (N_2537,In_124,In_941);
nand U2538 (N_2538,In_1399,In_404);
or U2539 (N_2539,In_2177,In_2154);
or U2540 (N_2540,In_2103,In_1054);
nand U2541 (N_2541,In_1073,In_578);
or U2542 (N_2542,In_1051,In_2259);
or U2543 (N_2543,In_454,In_968);
or U2544 (N_2544,In_609,In_971);
xnor U2545 (N_2545,In_1876,In_1096);
xor U2546 (N_2546,In_1859,In_1406);
nand U2547 (N_2547,In_1168,In_1736);
or U2548 (N_2548,In_131,In_272);
or U2549 (N_2549,In_2028,In_1999);
xnor U2550 (N_2550,In_819,In_804);
nor U2551 (N_2551,In_1277,In_403);
nor U2552 (N_2552,In_711,In_568);
nor U2553 (N_2553,In_784,In_535);
and U2554 (N_2554,In_1972,In_15);
nand U2555 (N_2555,In_2004,In_1558);
nor U2556 (N_2556,In_1461,In_1426);
xnor U2557 (N_2557,In_486,In_508);
nand U2558 (N_2558,In_1920,In_23);
nor U2559 (N_2559,In_1429,In_10);
and U2560 (N_2560,In_1945,In_1607);
nor U2561 (N_2561,In_2014,In_1573);
nand U2562 (N_2562,In_374,In_1100);
nand U2563 (N_2563,In_68,In_789);
and U2564 (N_2564,In_562,In_1488);
xor U2565 (N_2565,In_2070,In_1901);
xnor U2566 (N_2566,In_2316,In_222);
xor U2567 (N_2567,In_972,In_2178);
and U2568 (N_2568,In_2067,In_1022);
nor U2569 (N_2569,In_377,In_291);
xor U2570 (N_2570,In_850,In_1815);
and U2571 (N_2571,In_1028,In_41);
nor U2572 (N_2572,In_499,In_1198);
xor U2573 (N_2573,In_397,In_1893);
and U2574 (N_2574,In_663,In_1422);
nand U2575 (N_2575,In_2322,In_947);
nor U2576 (N_2576,In_435,In_952);
or U2577 (N_2577,In_1153,In_832);
or U2578 (N_2578,In_1249,In_2160);
nor U2579 (N_2579,In_380,In_148);
or U2580 (N_2580,In_1278,In_1231);
and U2581 (N_2581,In_70,In_2017);
nand U2582 (N_2582,In_1833,In_1032);
nor U2583 (N_2583,In_1955,In_2230);
or U2584 (N_2584,In_56,In_1928);
nand U2585 (N_2585,In_2234,In_1133);
and U2586 (N_2586,In_1217,In_217);
nand U2587 (N_2587,In_1281,In_2016);
nor U2588 (N_2588,In_1843,In_2003);
nor U2589 (N_2589,In_2067,In_1702);
or U2590 (N_2590,In_415,In_1617);
xnor U2591 (N_2591,In_1560,In_2156);
or U2592 (N_2592,In_148,In_2363);
and U2593 (N_2593,In_492,In_632);
or U2594 (N_2594,In_2031,In_2081);
and U2595 (N_2595,In_1886,In_2413);
nand U2596 (N_2596,In_1485,In_2294);
nand U2597 (N_2597,In_2328,In_478);
nand U2598 (N_2598,In_432,In_1509);
nor U2599 (N_2599,In_620,In_2002);
or U2600 (N_2600,In_2175,In_2288);
nand U2601 (N_2601,In_661,In_1820);
or U2602 (N_2602,In_621,In_2100);
nor U2603 (N_2603,In_133,In_995);
xor U2604 (N_2604,In_1807,In_349);
xnor U2605 (N_2605,In_439,In_275);
xnor U2606 (N_2606,In_1820,In_2083);
nand U2607 (N_2607,In_230,In_1757);
nor U2608 (N_2608,In_1969,In_253);
nor U2609 (N_2609,In_1823,In_1607);
and U2610 (N_2610,In_2021,In_1465);
or U2611 (N_2611,In_1942,In_2302);
nand U2612 (N_2612,In_1973,In_2106);
or U2613 (N_2613,In_1178,In_157);
and U2614 (N_2614,In_1217,In_1118);
nand U2615 (N_2615,In_1575,In_206);
or U2616 (N_2616,In_417,In_2348);
or U2617 (N_2617,In_1178,In_767);
nor U2618 (N_2618,In_947,In_409);
nor U2619 (N_2619,In_674,In_2161);
and U2620 (N_2620,In_2295,In_1691);
nand U2621 (N_2621,In_1254,In_697);
and U2622 (N_2622,In_947,In_1304);
nand U2623 (N_2623,In_1292,In_1440);
xor U2624 (N_2624,In_1105,In_114);
xnor U2625 (N_2625,In_756,In_173);
xnor U2626 (N_2626,In_2121,In_1341);
or U2627 (N_2627,In_422,In_421);
xor U2628 (N_2628,In_2354,In_736);
or U2629 (N_2629,In_1274,In_2214);
nand U2630 (N_2630,In_402,In_1406);
or U2631 (N_2631,In_389,In_526);
or U2632 (N_2632,In_366,In_1630);
and U2633 (N_2633,In_336,In_1554);
nor U2634 (N_2634,In_2223,In_253);
nand U2635 (N_2635,In_119,In_576);
or U2636 (N_2636,In_1971,In_667);
nor U2637 (N_2637,In_806,In_1168);
nand U2638 (N_2638,In_390,In_707);
nor U2639 (N_2639,In_1916,In_1827);
and U2640 (N_2640,In_2493,In_1335);
nand U2641 (N_2641,In_1923,In_910);
nand U2642 (N_2642,In_565,In_1579);
nand U2643 (N_2643,In_1628,In_1201);
nand U2644 (N_2644,In_1794,In_2496);
and U2645 (N_2645,In_783,In_370);
or U2646 (N_2646,In_1271,In_116);
nand U2647 (N_2647,In_1303,In_2154);
nor U2648 (N_2648,In_1701,In_2047);
or U2649 (N_2649,In_2187,In_1627);
and U2650 (N_2650,In_1573,In_2132);
nor U2651 (N_2651,In_2235,In_2142);
or U2652 (N_2652,In_1347,In_842);
xor U2653 (N_2653,In_21,In_961);
nor U2654 (N_2654,In_1705,In_1523);
nor U2655 (N_2655,In_84,In_1425);
or U2656 (N_2656,In_1116,In_405);
nor U2657 (N_2657,In_615,In_196);
and U2658 (N_2658,In_510,In_1595);
nand U2659 (N_2659,In_2394,In_2277);
nor U2660 (N_2660,In_202,In_1087);
nor U2661 (N_2661,In_1796,In_2002);
nand U2662 (N_2662,In_2489,In_1019);
nor U2663 (N_2663,In_766,In_1762);
nor U2664 (N_2664,In_404,In_883);
and U2665 (N_2665,In_2198,In_1936);
nor U2666 (N_2666,In_1446,In_71);
and U2667 (N_2667,In_886,In_149);
nor U2668 (N_2668,In_1785,In_2404);
and U2669 (N_2669,In_1152,In_398);
and U2670 (N_2670,In_2078,In_1920);
nor U2671 (N_2671,In_260,In_1703);
or U2672 (N_2672,In_643,In_1397);
nor U2673 (N_2673,In_267,In_395);
nor U2674 (N_2674,In_198,In_299);
nand U2675 (N_2675,In_1498,In_987);
or U2676 (N_2676,In_2452,In_1387);
or U2677 (N_2677,In_2109,In_1088);
and U2678 (N_2678,In_1786,In_2182);
or U2679 (N_2679,In_1389,In_1760);
nand U2680 (N_2680,In_156,In_2270);
or U2681 (N_2681,In_1850,In_1833);
nand U2682 (N_2682,In_1511,In_1127);
nand U2683 (N_2683,In_311,In_1690);
and U2684 (N_2684,In_222,In_2007);
nand U2685 (N_2685,In_2334,In_542);
xnor U2686 (N_2686,In_818,In_216);
and U2687 (N_2687,In_2200,In_187);
nand U2688 (N_2688,In_428,In_1888);
xor U2689 (N_2689,In_2294,In_2317);
or U2690 (N_2690,In_1332,In_1864);
or U2691 (N_2691,In_1766,In_470);
nand U2692 (N_2692,In_195,In_1314);
xnor U2693 (N_2693,In_1519,In_2398);
nor U2694 (N_2694,In_708,In_1451);
and U2695 (N_2695,In_1000,In_1049);
nand U2696 (N_2696,In_805,In_1490);
or U2697 (N_2697,In_548,In_2034);
nor U2698 (N_2698,In_1922,In_172);
nand U2699 (N_2699,In_1023,In_1319);
nand U2700 (N_2700,In_2405,In_1973);
nand U2701 (N_2701,In_2278,In_382);
and U2702 (N_2702,In_2369,In_1745);
nand U2703 (N_2703,In_1856,In_1718);
and U2704 (N_2704,In_1728,In_308);
and U2705 (N_2705,In_692,In_1801);
and U2706 (N_2706,In_685,In_2098);
nor U2707 (N_2707,In_1122,In_339);
nand U2708 (N_2708,In_561,In_564);
and U2709 (N_2709,In_2409,In_119);
and U2710 (N_2710,In_59,In_530);
xor U2711 (N_2711,In_863,In_199);
nand U2712 (N_2712,In_772,In_1564);
nand U2713 (N_2713,In_1013,In_1261);
nand U2714 (N_2714,In_1146,In_1017);
and U2715 (N_2715,In_432,In_2181);
and U2716 (N_2716,In_767,In_2149);
xnor U2717 (N_2717,In_1335,In_331);
and U2718 (N_2718,In_1465,In_1727);
or U2719 (N_2719,In_910,In_361);
nor U2720 (N_2720,In_1501,In_1880);
nand U2721 (N_2721,In_1612,In_943);
and U2722 (N_2722,In_1437,In_1244);
nor U2723 (N_2723,In_57,In_1488);
and U2724 (N_2724,In_635,In_1039);
nand U2725 (N_2725,In_939,In_779);
nand U2726 (N_2726,In_245,In_1182);
or U2727 (N_2727,In_2115,In_436);
or U2728 (N_2728,In_1467,In_214);
or U2729 (N_2729,In_185,In_149);
or U2730 (N_2730,In_1297,In_1886);
or U2731 (N_2731,In_713,In_1970);
or U2732 (N_2732,In_532,In_620);
nand U2733 (N_2733,In_1301,In_611);
or U2734 (N_2734,In_1378,In_1631);
nor U2735 (N_2735,In_1246,In_1861);
and U2736 (N_2736,In_1211,In_166);
nor U2737 (N_2737,In_2158,In_1044);
and U2738 (N_2738,In_552,In_1674);
or U2739 (N_2739,In_277,In_638);
and U2740 (N_2740,In_570,In_2335);
nand U2741 (N_2741,In_1447,In_287);
or U2742 (N_2742,In_1831,In_1276);
nor U2743 (N_2743,In_2116,In_1812);
xnor U2744 (N_2744,In_1237,In_488);
or U2745 (N_2745,In_2398,In_2017);
nand U2746 (N_2746,In_2225,In_1618);
nand U2747 (N_2747,In_13,In_803);
nand U2748 (N_2748,In_1846,In_113);
nand U2749 (N_2749,In_1223,In_1504);
and U2750 (N_2750,In_317,In_962);
or U2751 (N_2751,In_292,In_2461);
nor U2752 (N_2752,In_1850,In_168);
nor U2753 (N_2753,In_183,In_2034);
nor U2754 (N_2754,In_2435,In_1300);
or U2755 (N_2755,In_978,In_1160);
nor U2756 (N_2756,In_304,In_1877);
nand U2757 (N_2757,In_1427,In_953);
or U2758 (N_2758,In_2302,In_157);
nor U2759 (N_2759,In_1050,In_1546);
nor U2760 (N_2760,In_2282,In_292);
nor U2761 (N_2761,In_1163,In_197);
nor U2762 (N_2762,In_1136,In_913);
or U2763 (N_2763,In_2277,In_478);
or U2764 (N_2764,In_1812,In_1813);
and U2765 (N_2765,In_1992,In_2319);
or U2766 (N_2766,In_2063,In_2280);
or U2767 (N_2767,In_499,In_1918);
or U2768 (N_2768,In_2173,In_1610);
and U2769 (N_2769,In_2201,In_2219);
nand U2770 (N_2770,In_7,In_632);
nand U2771 (N_2771,In_750,In_2172);
and U2772 (N_2772,In_958,In_1549);
or U2773 (N_2773,In_2193,In_194);
and U2774 (N_2774,In_1847,In_61);
or U2775 (N_2775,In_420,In_1662);
nor U2776 (N_2776,In_1129,In_2079);
or U2777 (N_2777,In_344,In_1549);
xnor U2778 (N_2778,In_1532,In_1408);
nand U2779 (N_2779,In_2276,In_2151);
and U2780 (N_2780,In_1793,In_1603);
nand U2781 (N_2781,In_1196,In_145);
xnor U2782 (N_2782,In_78,In_2055);
or U2783 (N_2783,In_2246,In_401);
nand U2784 (N_2784,In_1323,In_1675);
and U2785 (N_2785,In_395,In_1417);
or U2786 (N_2786,In_529,In_911);
nor U2787 (N_2787,In_1670,In_2252);
nor U2788 (N_2788,In_894,In_710);
or U2789 (N_2789,In_1924,In_713);
and U2790 (N_2790,In_1454,In_160);
or U2791 (N_2791,In_451,In_2221);
and U2792 (N_2792,In_2351,In_2069);
or U2793 (N_2793,In_117,In_263);
nor U2794 (N_2794,In_1634,In_400);
and U2795 (N_2795,In_1558,In_197);
and U2796 (N_2796,In_2146,In_1921);
nand U2797 (N_2797,In_786,In_1068);
and U2798 (N_2798,In_824,In_2232);
nand U2799 (N_2799,In_1428,In_384);
nor U2800 (N_2800,In_2162,In_1472);
nand U2801 (N_2801,In_369,In_81);
nand U2802 (N_2802,In_2265,In_1755);
or U2803 (N_2803,In_1987,In_1981);
nor U2804 (N_2804,In_1807,In_2034);
nand U2805 (N_2805,In_41,In_1375);
nand U2806 (N_2806,In_549,In_597);
nand U2807 (N_2807,In_1660,In_1903);
nand U2808 (N_2808,In_1100,In_269);
or U2809 (N_2809,In_772,In_2072);
xor U2810 (N_2810,In_2252,In_2202);
or U2811 (N_2811,In_1935,In_131);
and U2812 (N_2812,In_342,In_632);
and U2813 (N_2813,In_68,In_0);
nor U2814 (N_2814,In_2489,In_1802);
and U2815 (N_2815,In_1719,In_1817);
nor U2816 (N_2816,In_1862,In_1334);
or U2817 (N_2817,In_1480,In_1206);
or U2818 (N_2818,In_1623,In_405);
nand U2819 (N_2819,In_1171,In_2433);
nand U2820 (N_2820,In_2225,In_2263);
xor U2821 (N_2821,In_272,In_338);
and U2822 (N_2822,In_388,In_829);
or U2823 (N_2823,In_1205,In_1576);
nor U2824 (N_2824,In_836,In_53);
or U2825 (N_2825,In_420,In_557);
nand U2826 (N_2826,In_1544,In_1552);
and U2827 (N_2827,In_679,In_2223);
or U2828 (N_2828,In_834,In_1129);
and U2829 (N_2829,In_2379,In_222);
xor U2830 (N_2830,In_1480,In_1715);
and U2831 (N_2831,In_1313,In_327);
nor U2832 (N_2832,In_2065,In_791);
nor U2833 (N_2833,In_1728,In_910);
or U2834 (N_2834,In_2475,In_1053);
or U2835 (N_2835,In_1854,In_934);
or U2836 (N_2836,In_1041,In_930);
nand U2837 (N_2837,In_1125,In_2111);
nand U2838 (N_2838,In_395,In_4);
nor U2839 (N_2839,In_2359,In_1804);
xor U2840 (N_2840,In_1685,In_1427);
nor U2841 (N_2841,In_699,In_1749);
xnor U2842 (N_2842,In_2366,In_905);
nand U2843 (N_2843,In_1110,In_277);
nor U2844 (N_2844,In_1604,In_172);
nor U2845 (N_2845,In_2401,In_1365);
and U2846 (N_2846,In_1480,In_317);
or U2847 (N_2847,In_1913,In_2133);
nor U2848 (N_2848,In_222,In_1597);
and U2849 (N_2849,In_1828,In_887);
or U2850 (N_2850,In_2315,In_134);
nor U2851 (N_2851,In_198,In_2297);
nand U2852 (N_2852,In_804,In_2458);
and U2853 (N_2853,In_121,In_308);
and U2854 (N_2854,In_502,In_362);
and U2855 (N_2855,In_40,In_188);
nand U2856 (N_2856,In_118,In_1478);
or U2857 (N_2857,In_1905,In_308);
or U2858 (N_2858,In_1863,In_2211);
and U2859 (N_2859,In_2075,In_2081);
and U2860 (N_2860,In_619,In_1684);
nor U2861 (N_2861,In_1480,In_1968);
nand U2862 (N_2862,In_885,In_7);
and U2863 (N_2863,In_2293,In_428);
nand U2864 (N_2864,In_2305,In_2498);
nor U2865 (N_2865,In_2203,In_2419);
nor U2866 (N_2866,In_742,In_1419);
nand U2867 (N_2867,In_1938,In_614);
nand U2868 (N_2868,In_319,In_823);
or U2869 (N_2869,In_578,In_2051);
or U2870 (N_2870,In_1491,In_246);
and U2871 (N_2871,In_501,In_408);
nand U2872 (N_2872,In_527,In_2303);
and U2873 (N_2873,In_613,In_1823);
nand U2874 (N_2874,In_24,In_1796);
and U2875 (N_2875,In_2183,In_1356);
xnor U2876 (N_2876,In_1909,In_2052);
or U2877 (N_2877,In_937,In_1003);
or U2878 (N_2878,In_113,In_1039);
and U2879 (N_2879,In_2400,In_2170);
nor U2880 (N_2880,In_1332,In_197);
and U2881 (N_2881,In_1869,In_1776);
or U2882 (N_2882,In_2443,In_1191);
nand U2883 (N_2883,In_1264,In_749);
and U2884 (N_2884,In_1663,In_986);
nand U2885 (N_2885,In_996,In_2408);
nand U2886 (N_2886,In_888,In_365);
or U2887 (N_2887,In_1942,In_2197);
or U2888 (N_2888,In_1714,In_1698);
nand U2889 (N_2889,In_655,In_882);
and U2890 (N_2890,In_1331,In_452);
nand U2891 (N_2891,In_432,In_2256);
nor U2892 (N_2892,In_1866,In_1776);
nand U2893 (N_2893,In_1552,In_1468);
or U2894 (N_2894,In_652,In_644);
nand U2895 (N_2895,In_27,In_725);
and U2896 (N_2896,In_1260,In_857);
nand U2897 (N_2897,In_1337,In_1757);
nor U2898 (N_2898,In_446,In_2419);
nand U2899 (N_2899,In_880,In_1907);
or U2900 (N_2900,In_637,In_353);
xor U2901 (N_2901,In_850,In_2371);
nor U2902 (N_2902,In_157,In_2270);
and U2903 (N_2903,In_166,In_2206);
or U2904 (N_2904,In_871,In_1462);
nor U2905 (N_2905,In_1347,In_99);
and U2906 (N_2906,In_482,In_1465);
nand U2907 (N_2907,In_1630,In_525);
or U2908 (N_2908,In_1075,In_442);
nand U2909 (N_2909,In_1830,In_1708);
nor U2910 (N_2910,In_249,In_1530);
nor U2911 (N_2911,In_2026,In_858);
xor U2912 (N_2912,In_1020,In_1119);
xnor U2913 (N_2913,In_1203,In_1835);
nand U2914 (N_2914,In_234,In_2134);
nand U2915 (N_2915,In_519,In_977);
and U2916 (N_2916,In_2030,In_710);
nor U2917 (N_2917,In_187,In_271);
nand U2918 (N_2918,In_1173,In_22);
and U2919 (N_2919,In_281,In_1057);
nor U2920 (N_2920,In_1146,In_111);
or U2921 (N_2921,In_806,In_414);
and U2922 (N_2922,In_2077,In_1124);
nand U2923 (N_2923,In_1673,In_34);
xor U2924 (N_2924,In_814,In_1502);
and U2925 (N_2925,In_1441,In_1940);
nand U2926 (N_2926,In_372,In_1914);
nor U2927 (N_2927,In_979,In_1739);
or U2928 (N_2928,In_682,In_1647);
nor U2929 (N_2929,In_797,In_1478);
nand U2930 (N_2930,In_2218,In_963);
xnor U2931 (N_2931,In_654,In_1453);
and U2932 (N_2932,In_1275,In_533);
and U2933 (N_2933,In_1765,In_676);
and U2934 (N_2934,In_1210,In_23);
and U2935 (N_2935,In_2029,In_771);
xor U2936 (N_2936,In_2251,In_1770);
or U2937 (N_2937,In_1886,In_1405);
xnor U2938 (N_2938,In_2066,In_108);
and U2939 (N_2939,In_327,In_674);
nor U2940 (N_2940,In_673,In_1379);
or U2941 (N_2941,In_208,In_315);
nor U2942 (N_2942,In_120,In_261);
or U2943 (N_2943,In_318,In_579);
nand U2944 (N_2944,In_1676,In_29);
or U2945 (N_2945,In_326,In_1726);
or U2946 (N_2946,In_1873,In_45);
or U2947 (N_2947,In_2059,In_1106);
nor U2948 (N_2948,In_737,In_1568);
nor U2949 (N_2949,In_2284,In_2055);
nor U2950 (N_2950,In_1887,In_600);
nor U2951 (N_2951,In_1288,In_1272);
and U2952 (N_2952,In_1243,In_2078);
nor U2953 (N_2953,In_2118,In_119);
or U2954 (N_2954,In_117,In_556);
or U2955 (N_2955,In_901,In_80);
xnor U2956 (N_2956,In_708,In_1560);
or U2957 (N_2957,In_874,In_999);
or U2958 (N_2958,In_406,In_1445);
and U2959 (N_2959,In_395,In_542);
nor U2960 (N_2960,In_2209,In_1873);
nor U2961 (N_2961,In_1725,In_162);
nand U2962 (N_2962,In_1982,In_1239);
nor U2963 (N_2963,In_1237,In_415);
or U2964 (N_2964,In_1137,In_473);
or U2965 (N_2965,In_1848,In_102);
nor U2966 (N_2966,In_622,In_868);
nand U2967 (N_2967,In_2377,In_2273);
and U2968 (N_2968,In_120,In_1951);
or U2969 (N_2969,In_379,In_2444);
or U2970 (N_2970,In_667,In_270);
or U2971 (N_2971,In_1193,In_1642);
or U2972 (N_2972,In_46,In_904);
nor U2973 (N_2973,In_2382,In_2366);
xnor U2974 (N_2974,In_1980,In_1518);
or U2975 (N_2975,In_2027,In_687);
and U2976 (N_2976,In_1261,In_249);
nand U2977 (N_2977,In_1864,In_1649);
or U2978 (N_2978,In_631,In_1070);
and U2979 (N_2979,In_541,In_1564);
nor U2980 (N_2980,In_2143,In_2274);
and U2981 (N_2981,In_539,In_736);
nor U2982 (N_2982,In_1605,In_1437);
and U2983 (N_2983,In_740,In_1421);
xnor U2984 (N_2984,In_1258,In_1652);
or U2985 (N_2985,In_431,In_1665);
nand U2986 (N_2986,In_202,In_1);
or U2987 (N_2987,In_2343,In_867);
or U2988 (N_2988,In_1559,In_921);
and U2989 (N_2989,In_1237,In_2349);
and U2990 (N_2990,In_1052,In_866);
nand U2991 (N_2991,In_630,In_749);
nor U2992 (N_2992,In_977,In_1653);
nand U2993 (N_2993,In_758,In_1945);
or U2994 (N_2994,In_1243,In_1178);
nand U2995 (N_2995,In_2366,In_1847);
nor U2996 (N_2996,In_1394,In_1680);
nand U2997 (N_2997,In_846,In_1890);
or U2998 (N_2998,In_328,In_1500);
nand U2999 (N_2999,In_533,In_1031);
nor U3000 (N_3000,In_398,In_1868);
or U3001 (N_3001,In_2017,In_339);
and U3002 (N_3002,In_1665,In_2263);
or U3003 (N_3003,In_295,In_1292);
or U3004 (N_3004,In_1540,In_2356);
nor U3005 (N_3005,In_348,In_1924);
and U3006 (N_3006,In_759,In_931);
or U3007 (N_3007,In_505,In_33);
and U3008 (N_3008,In_664,In_2350);
and U3009 (N_3009,In_2093,In_1885);
nand U3010 (N_3010,In_1218,In_774);
nand U3011 (N_3011,In_1734,In_1439);
nor U3012 (N_3012,In_49,In_1228);
nor U3013 (N_3013,In_1398,In_703);
xor U3014 (N_3014,In_2412,In_1924);
xor U3015 (N_3015,In_2099,In_1409);
nand U3016 (N_3016,In_475,In_1216);
nor U3017 (N_3017,In_201,In_2014);
nor U3018 (N_3018,In_396,In_1873);
and U3019 (N_3019,In_2124,In_451);
or U3020 (N_3020,In_1873,In_1127);
and U3021 (N_3021,In_1906,In_1875);
or U3022 (N_3022,In_824,In_330);
nand U3023 (N_3023,In_2292,In_1724);
and U3024 (N_3024,In_1310,In_1912);
or U3025 (N_3025,In_1968,In_815);
nor U3026 (N_3026,In_974,In_1865);
nand U3027 (N_3027,In_920,In_380);
and U3028 (N_3028,In_2178,In_1719);
nor U3029 (N_3029,In_1946,In_2378);
nand U3030 (N_3030,In_359,In_1881);
nor U3031 (N_3031,In_326,In_559);
nand U3032 (N_3032,In_1544,In_683);
and U3033 (N_3033,In_38,In_533);
nor U3034 (N_3034,In_462,In_2413);
and U3035 (N_3035,In_2103,In_2470);
or U3036 (N_3036,In_1910,In_1457);
and U3037 (N_3037,In_1680,In_524);
and U3038 (N_3038,In_878,In_357);
xnor U3039 (N_3039,In_325,In_1507);
and U3040 (N_3040,In_2132,In_1972);
and U3041 (N_3041,In_65,In_751);
xor U3042 (N_3042,In_2304,In_2420);
nand U3043 (N_3043,In_1926,In_2185);
and U3044 (N_3044,In_2239,In_1223);
xor U3045 (N_3045,In_351,In_1541);
and U3046 (N_3046,In_1530,In_1248);
xor U3047 (N_3047,In_625,In_2015);
nand U3048 (N_3048,In_1917,In_2136);
and U3049 (N_3049,In_1228,In_1178);
xor U3050 (N_3050,In_2285,In_1479);
nor U3051 (N_3051,In_1886,In_2344);
nand U3052 (N_3052,In_1078,In_788);
and U3053 (N_3053,In_2353,In_2458);
nor U3054 (N_3054,In_1032,In_1682);
nor U3055 (N_3055,In_1449,In_1880);
or U3056 (N_3056,In_78,In_35);
nor U3057 (N_3057,In_878,In_1834);
nand U3058 (N_3058,In_1147,In_790);
nand U3059 (N_3059,In_2147,In_2091);
or U3060 (N_3060,In_2042,In_74);
and U3061 (N_3061,In_2284,In_247);
xor U3062 (N_3062,In_507,In_139);
or U3063 (N_3063,In_2251,In_2231);
nor U3064 (N_3064,In_2075,In_239);
and U3065 (N_3065,In_1485,In_1364);
nand U3066 (N_3066,In_1350,In_2306);
or U3067 (N_3067,In_2016,In_396);
nand U3068 (N_3068,In_1325,In_1710);
or U3069 (N_3069,In_1021,In_2042);
or U3070 (N_3070,In_466,In_2378);
and U3071 (N_3071,In_2482,In_237);
or U3072 (N_3072,In_550,In_314);
and U3073 (N_3073,In_1219,In_1401);
nor U3074 (N_3074,In_707,In_1956);
nor U3075 (N_3075,In_1078,In_2458);
nor U3076 (N_3076,In_479,In_2475);
or U3077 (N_3077,In_1685,In_1036);
or U3078 (N_3078,In_673,In_547);
nand U3079 (N_3079,In_1144,In_918);
or U3080 (N_3080,In_248,In_2349);
and U3081 (N_3081,In_796,In_1577);
nand U3082 (N_3082,In_970,In_1045);
xor U3083 (N_3083,In_546,In_1111);
xnor U3084 (N_3084,In_1153,In_932);
and U3085 (N_3085,In_1938,In_186);
and U3086 (N_3086,In_447,In_224);
and U3087 (N_3087,In_2253,In_1268);
nor U3088 (N_3088,In_244,In_275);
and U3089 (N_3089,In_2308,In_430);
nand U3090 (N_3090,In_369,In_363);
nand U3091 (N_3091,In_2437,In_421);
or U3092 (N_3092,In_386,In_2388);
or U3093 (N_3093,In_2231,In_1494);
nand U3094 (N_3094,In_1140,In_835);
nand U3095 (N_3095,In_1091,In_2010);
nand U3096 (N_3096,In_1895,In_14);
nor U3097 (N_3097,In_1965,In_2472);
or U3098 (N_3098,In_1119,In_1801);
nor U3099 (N_3099,In_514,In_2407);
nand U3100 (N_3100,In_486,In_923);
and U3101 (N_3101,In_1137,In_1297);
and U3102 (N_3102,In_66,In_2004);
nor U3103 (N_3103,In_452,In_1699);
nand U3104 (N_3104,In_2228,In_720);
or U3105 (N_3105,In_2058,In_854);
nor U3106 (N_3106,In_2135,In_1739);
or U3107 (N_3107,In_1654,In_2392);
nand U3108 (N_3108,In_2105,In_597);
or U3109 (N_3109,In_1910,In_2152);
nand U3110 (N_3110,In_1835,In_1385);
and U3111 (N_3111,In_327,In_824);
or U3112 (N_3112,In_1078,In_1364);
nand U3113 (N_3113,In_2152,In_714);
or U3114 (N_3114,In_1877,In_1582);
and U3115 (N_3115,In_2448,In_424);
nand U3116 (N_3116,In_2433,In_2162);
nand U3117 (N_3117,In_419,In_862);
and U3118 (N_3118,In_1343,In_2435);
nand U3119 (N_3119,In_1688,In_1653);
and U3120 (N_3120,In_1304,In_732);
nor U3121 (N_3121,In_1867,In_1210);
or U3122 (N_3122,In_876,In_1989);
xor U3123 (N_3123,In_1218,In_619);
nand U3124 (N_3124,In_479,In_765);
nand U3125 (N_3125,N_2728,N_1678);
nor U3126 (N_3126,N_1412,N_3015);
xnor U3127 (N_3127,N_1582,N_1058);
and U3128 (N_3128,N_883,N_1866);
nor U3129 (N_3129,N_327,N_211);
nor U3130 (N_3130,N_1192,N_1804);
nand U3131 (N_3131,N_1629,N_2755);
nand U3132 (N_3132,N_2568,N_3098);
or U3133 (N_3133,N_1294,N_181);
nor U3134 (N_3134,N_1300,N_278);
nor U3135 (N_3135,N_1765,N_397);
and U3136 (N_3136,N_460,N_2454);
nor U3137 (N_3137,N_1504,N_1221);
or U3138 (N_3138,N_1716,N_368);
xor U3139 (N_3139,N_2994,N_1074);
nor U3140 (N_3140,N_781,N_3017);
nor U3141 (N_3141,N_1578,N_1186);
nor U3142 (N_3142,N_1906,N_1386);
or U3143 (N_3143,N_1503,N_1828);
xnor U3144 (N_3144,N_229,N_1704);
and U3145 (N_3145,N_2777,N_1585);
or U3146 (N_3146,N_1448,N_410);
nand U3147 (N_3147,N_2687,N_499);
nand U3148 (N_3148,N_1723,N_844);
xnor U3149 (N_3149,N_1075,N_651);
or U3150 (N_3150,N_2092,N_2027);
or U3151 (N_3151,N_816,N_1392);
or U3152 (N_3152,N_593,N_1326);
nor U3153 (N_3153,N_1683,N_1854);
and U3154 (N_3154,N_1462,N_2465);
and U3155 (N_3155,N_1897,N_1528);
and U3156 (N_3156,N_792,N_306);
nand U3157 (N_3157,N_2914,N_1441);
nor U3158 (N_3158,N_1818,N_1374);
and U3159 (N_3159,N_517,N_388);
nand U3160 (N_3160,N_2525,N_70);
xnor U3161 (N_3161,N_1369,N_1244);
or U3162 (N_3162,N_2952,N_148);
or U3163 (N_3163,N_1946,N_1117);
nand U3164 (N_3164,N_2129,N_2577);
or U3165 (N_3165,N_833,N_1486);
nor U3166 (N_3166,N_1699,N_1167);
nor U3167 (N_3167,N_1144,N_2721);
nor U3168 (N_3168,N_2285,N_1176);
nand U3169 (N_3169,N_1129,N_2245);
xor U3170 (N_3170,N_2183,N_2156);
nor U3171 (N_3171,N_2540,N_1912);
and U3172 (N_3172,N_2731,N_2303);
nand U3173 (N_3173,N_2034,N_117);
xor U3174 (N_3174,N_2225,N_2533);
or U3175 (N_3175,N_2956,N_17);
and U3176 (N_3176,N_2154,N_1188);
xnor U3177 (N_3177,N_1230,N_56);
and U3178 (N_3178,N_2595,N_1212);
nand U3179 (N_3179,N_2060,N_969);
or U3180 (N_3180,N_2635,N_3018);
nand U3181 (N_3181,N_2006,N_2432);
and U3182 (N_3182,N_2502,N_1204);
or U3183 (N_3183,N_94,N_2246);
or U3184 (N_3184,N_1352,N_1123);
and U3185 (N_3185,N_860,N_374);
nand U3186 (N_3186,N_1868,N_2624);
nand U3187 (N_3187,N_28,N_987);
nand U3188 (N_3188,N_756,N_1611);
nor U3189 (N_3189,N_878,N_2761);
and U3190 (N_3190,N_616,N_2269);
nand U3191 (N_3191,N_2516,N_438);
nand U3192 (N_3192,N_1207,N_2035);
or U3193 (N_3193,N_347,N_2209);
and U3194 (N_3194,N_2153,N_1345);
nand U3195 (N_3195,N_282,N_2016);
nor U3196 (N_3196,N_2140,N_2998);
nor U3197 (N_3197,N_632,N_275);
nand U3198 (N_3198,N_2809,N_2707);
nand U3199 (N_3199,N_526,N_149);
or U3200 (N_3200,N_1876,N_2197);
nand U3201 (N_3201,N_1776,N_3032);
or U3202 (N_3202,N_34,N_780);
nand U3203 (N_3203,N_2498,N_239);
nor U3204 (N_3204,N_1996,N_1577);
nand U3205 (N_3205,N_2822,N_1157);
or U3206 (N_3206,N_2037,N_900);
nor U3207 (N_3207,N_1251,N_185);
nor U3208 (N_3208,N_1465,N_2767);
xnor U3209 (N_3209,N_947,N_2446);
or U3210 (N_3210,N_596,N_2388);
xnor U3211 (N_3211,N_1275,N_2987);
nand U3212 (N_3212,N_2840,N_1116);
and U3213 (N_3213,N_2575,N_1012);
nand U3214 (N_3214,N_458,N_906);
and U3215 (N_3215,N_1241,N_1359);
or U3216 (N_3216,N_1601,N_233);
or U3217 (N_3217,N_289,N_1179);
and U3218 (N_3218,N_2397,N_1424);
or U3219 (N_3219,N_2963,N_2050);
and U3220 (N_3220,N_1226,N_2729);
and U3221 (N_3221,N_2422,N_1445);
nor U3222 (N_3222,N_779,N_3097);
nor U3223 (N_3223,N_662,N_1924);
or U3224 (N_3224,N_2002,N_49);
or U3225 (N_3225,N_288,N_1256);
and U3226 (N_3226,N_1978,N_2828);
and U3227 (N_3227,N_1511,N_1314);
nor U3228 (N_3228,N_3026,N_1926);
or U3229 (N_3229,N_2769,N_2574);
xnor U3230 (N_3230,N_2396,N_3052);
nor U3231 (N_3231,N_2940,N_144);
or U3232 (N_3232,N_3068,N_2166);
or U3233 (N_3233,N_715,N_1846);
or U3234 (N_3234,N_1457,N_535);
or U3235 (N_3235,N_1280,N_2055);
nand U3236 (N_3236,N_2988,N_2336);
and U3237 (N_3237,N_697,N_669);
or U3238 (N_3238,N_99,N_1108);
nand U3239 (N_3239,N_1677,N_107);
nor U3240 (N_3240,N_751,N_1217);
nand U3241 (N_3241,N_445,N_1834);
nand U3242 (N_3242,N_3027,N_2487);
or U3243 (N_3243,N_2556,N_796);
nor U3244 (N_3244,N_1891,N_655);
and U3245 (N_3245,N_2645,N_1824);
nand U3246 (N_3246,N_2636,N_3058);
nand U3247 (N_3247,N_2118,N_2802);
nor U3248 (N_3248,N_262,N_2283);
nand U3249 (N_3249,N_1443,N_300);
nand U3250 (N_3250,N_2992,N_1248);
nor U3251 (N_3251,N_970,N_1228);
nand U3252 (N_3252,N_2036,N_2149);
or U3253 (N_3253,N_162,N_2794);
nor U3254 (N_3254,N_2261,N_281);
and U3255 (N_3255,N_483,N_267);
xnor U3256 (N_3256,N_2929,N_2862);
nand U3257 (N_3257,N_894,N_90);
xor U3258 (N_3258,N_691,N_1184);
or U3259 (N_3259,N_2483,N_2365);
or U3260 (N_3260,N_1253,N_415);
nand U3261 (N_3261,N_319,N_2028);
and U3262 (N_3262,N_2442,N_2095);
and U3263 (N_3263,N_113,N_530);
xnor U3264 (N_3264,N_1757,N_2468);
nand U3265 (N_3265,N_826,N_63);
xnor U3266 (N_3266,N_2870,N_2739);
nand U3267 (N_3267,N_1049,N_2850);
nor U3268 (N_3268,N_961,N_1975);
xor U3269 (N_3269,N_1954,N_2589);
and U3270 (N_3270,N_2832,N_1728);
xnor U3271 (N_3271,N_854,N_2298);
or U3272 (N_3272,N_732,N_1466);
or U3273 (N_3273,N_150,N_1539);
or U3274 (N_3274,N_451,N_1567);
nor U3275 (N_3275,N_509,N_227);
nand U3276 (N_3276,N_2811,N_98);
nor U3277 (N_3277,N_750,N_1974);
nand U3278 (N_3278,N_1496,N_1853);
or U3279 (N_3279,N_856,N_1);
and U3280 (N_3280,N_396,N_1752);
nand U3281 (N_3281,N_882,N_1324);
nand U3282 (N_3282,N_1463,N_2404);
and U3283 (N_3283,N_2205,N_84);
nor U3284 (N_3284,N_159,N_543);
nor U3285 (N_3285,N_2433,N_1426);
nand U3286 (N_3286,N_2380,N_2594);
and U3287 (N_3287,N_2909,N_2390);
and U3288 (N_3288,N_515,N_681);
xor U3289 (N_3289,N_1003,N_488);
xnor U3290 (N_3290,N_177,N_2180);
and U3291 (N_3291,N_1987,N_644);
or U3292 (N_3292,N_2999,N_2689);
and U3293 (N_3293,N_168,N_1387);
or U3294 (N_3294,N_2893,N_119);
nand U3295 (N_3295,N_2626,N_1415);
nand U3296 (N_3296,N_114,N_2529);
or U3297 (N_3297,N_1737,N_1825);
or U3298 (N_3298,N_2743,N_680);
nor U3299 (N_3299,N_529,N_1024);
nand U3300 (N_3300,N_1316,N_2590);
and U3301 (N_3301,N_1779,N_3061);
xnor U3302 (N_3302,N_2795,N_283);
and U3303 (N_3303,N_1715,N_2207);
xnor U3304 (N_3304,N_65,N_2165);
nor U3305 (N_3305,N_716,N_1771);
or U3306 (N_3306,N_2376,N_1794);
nor U3307 (N_3307,N_2251,N_2668);
nor U3308 (N_3308,N_139,N_1812);
nand U3309 (N_3309,N_654,N_2872);
or U3310 (N_3310,N_258,N_138);
xnor U3311 (N_3311,N_1178,N_320);
nand U3312 (N_3312,N_2733,N_1410);
nand U3313 (N_3313,N_510,N_2902);
and U3314 (N_3314,N_2810,N_994);
and U3315 (N_3315,N_2409,N_171);
or U3316 (N_3316,N_2650,N_1747);
and U3317 (N_3317,N_1498,N_2630);
nor U3318 (N_3318,N_2351,N_2646);
or U3319 (N_3319,N_3116,N_2657);
nor U3320 (N_3320,N_1833,N_182);
nor U3321 (N_3321,N_3094,N_2905);
nand U3322 (N_3322,N_1686,N_2638);
nor U3323 (N_3323,N_2127,N_2497);
or U3324 (N_3324,N_904,N_3117);
nand U3325 (N_3325,N_2248,N_1624);
nand U3326 (N_3326,N_2232,N_124);
xor U3327 (N_3327,N_763,N_2263);
nand U3328 (N_3328,N_224,N_2470);
nor U3329 (N_3329,N_1468,N_1673);
nand U3330 (N_3330,N_131,N_271);
nor U3331 (N_3331,N_1175,N_1357);
xor U3332 (N_3332,N_2607,N_230);
nor U3333 (N_3333,N_785,N_197);
or U3334 (N_3334,N_1620,N_175);
nor U3335 (N_3335,N_2756,N_1181);
nor U3336 (N_3336,N_196,N_711);
nor U3337 (N_3337,N_1666,N_2026);
or U3338 (N_3338,N_2892,N_400);
nor U3339 (N_3339,N_2679,N_2184);
nor U3340 (N_3340,N_1682,N_853);
and U3341 (N_3341,N_2538,N_2262);
xor U3342 (N_3342,N_2210,N_2472);
and U3343 (N_3343,N_1231,N_3041);
nand U3344 (N_3344,N_2667,N_471);
nor U3345 (N_3345,N_161,N_3114);
nand U3346 (N_3346,N_427,N_414);
nand U3347 (N_3347,N_2356,N_2882);
nor U3348 (N_3348,N_1595,N_3118);
and U3349 (N_3349,N_85,N_2337);
or U3350 (N_3350,N_2951,N_1636);
nand U3351 (N_3351,N_494,N_2633);
and U3352 (N_3352,N_2628,N_292);
nor U3353 (N_3353,N_2461,N_2255);
or U3354 (N_3354,N_2946,N_3102);
nand U3355 (N_3355,N_1870,N_2596);
or U3356 (N_3356,N_670,N_495);
nand U3357 (N_3357,N_992,N_1836);
nor U3358 (N_3358,N_2553,N_1667);
nor U3359 (N_3359,N_787,N_633);
nor U3360 (N_3360,N_1336,N_46);
nor U3361 (N_3361,N_1398,N_805);
nand U3362 (N_3362,N_1235,N_1646);
nand U3363 (N_3363,N_837,N_1533);
and U3364 (N_3364,N_696,N_761);
nor U3365 (N_3365,N_1238,N_1898);
and U3366 (N_3366,N_2128,N_2250);
or U3367 (N_3367,N_2825,N_454);
nor U3368 (N_3368,N_2955,N_1239);
or U3369 (N_3369,N_1132,N_2355);
nor U3370 (N_3370,N_2482,N_1696);
nor U3371 (N_3371,N_1334,N_2344);
or U3372 (N_3372,N_2964,N_467);
nand U3373 (N_3373,N_1951,N_842);
or U3374 (N_3374,N_2239,N_1007);
or U3375 (N_3375,N_2204,N_1093);
or U3376 (N_3376,N_1698,N_1370);
nor U3377 (N_3377,N_2307,N_2325);
and U3378 (N_3378,N_2869,N_525);
and U3379 (N_3379,N_2928,N_429);
nor U3380 (N_3380,N_1397,N_1489);
nor U3381 (N_3381,N_3012,N_1593);
nor U3382 (N_3382,N_1384,N_2868);
xor U3383 (N_3383,N_1830,N_565);
nor U3384 (N_3384,N_3120,N_2618);
or U3385 (N_3385,N_1842,N_1546);
nand U3386 (N_3386,N_2823,N_1621);
xor U3387 (N_3387,N_1979,N_1071);
nor U3388 (N_3388,N_1261,N_2906);
and U3389 (N_3389,N_877,N_563);
nand U3390 (N_3390,N_2069,N_2780);
nand U3391 (N_3391,N_2517,N_305);
or U3392 (N_3392,N_567,N_1930);
or U3393 (N_3393,N_619,N_1714);
nor U3394 (N_3394,N_1029,N_2421);
or U3395 (N_3395,N_285,N_103);
nor U3396 (N_3396,N_1764,N_834);
nand U3397 (N_3397,N_442,N_2073);
nor U3398 (N_3398,N_2690,N_2723);
and U3399 (N_3399,N_949,N_1135);
and U3400 (N_3400,N_1363,N_800);
nor U3401 (N_3401,N_1148,N_2136);
or U3402 (N_3402,N_653,N_973);
and U3403 (N_3403,N_2550,N_3083);
nor U3404 (N_3404,N_2453,N_2025);
nand U3405 (N_3405,N_980,N_1480);
nand U3406 (N_3406,N_1614,N_3050);
or U3407 (N_3407,N_322,N_23);
nor U3408 (N_3408,N_2041,N_1695);
and U3409 (N_3409,N_1660,N_1894);
nand U3410 (N_3410,N_3010,N_1527);
and U3411 (N_3411,N_1201,N_1992);
and U3412 (N_3412,N_1915,N_2314);
nor U3413 (N_3413,N_2427,N_614);
and U3414 (N_3414,N_999,N_3100);
nand U3415 (N_3415,N_2061,N_1240);
or U3416 (N_3416,N_1933,N_2889);
or U3417 (N_3417,N_1113,N_922);
nand U3418 (N_3418,N_2477,N_3040);
or U3419 (N_3419,N_2576,N_2692);
and U3420 (N_3420,N_222,N_2324);
nand U3421 (N_3421,N_2853,N_2103);
or U3422 (N_3422,N_1160,N_20);
and U3423 (N_3423,N_2503,N_2284);
or U3424 (N_3424,N_504,N_2785);
or U3425 (N_3425,N_2078,N_588);
xnor U3426 (N_3426,N_830,N_1631);
or U3427 (N_3427,N_1538,N_2168);
nor U3428 (N_3428,N_1396,N_1705);
or U3429 (N_3429,N_1761,N_2102);
nor U3430 (N_3430,N_933,N_1997);
and U3431 (N_3431,N_1693,N_3104);
or U3432 (N_3432,N_424,N_1990);
and U3433 (N_3433,N_753,N_2022);
nand U3434 (N_3434,N_544,N_2004);
and U3435 (N_3435,N_1454,N_241);
nand U3436 (N_3436,N_2977,N_342);
nand U3437 (N_3437,N_1436,N_1409);
nand U3438 (N_3438,N_1786,N_1375);
nand U3439 (N_3439,N_38,N_2975);
nand U3440 (N_3440,N_967,N_1080);
nand U3441 (N_3441,N_1483,N_1420);
nor U3442 (N_3442,N_3006,N_343);
nor U3443 (N_3443,N_1896,N_885);
or U3444 (N_3444,N_2530,N_2105);
xnor U3445 (N_3445,N_13,N_1822);
nand U3446 (N_3446,N_353,N_2849);
nand U3447 (N_3447,N_2973,N_174);
and U3448 (N_3448,N_946,N_1164);
nor U3449 (N_3449,N_915,N_1152);
nand U3450 (N_3450,N_2684,N_804);
nand U3451 (N_3451,N_2212,N_940);
nand U3452 (N_3452,N_1471,N_1808);
or U3453 (N_3453,N_1576,N_1855);
or U3454 (N_3454,N_811,N_996);
nand U3455 (N_3455,N_236,N_2367);
or U3456 (N_3456,N_1917,N_694);
nor U3457 (N_3457,N_3,N_96);
nand U3458 (N_3458,N_2171,N_1858);
or U3459 (N_3459,N_2411,N_80);
nand U3460 (N_3460,N_752,N_2490);
nand U3461 (N_3461,N_1865,N_2867);
xnor U3462 (N_3462,N_2455,N_1684);
and U3463 (N_3463,N_2837,N_1881);
and U3464 (N_3464,N_1928,N_2895);
nand U3465 (N_3465,N_1028,N_741);
nor U3466 (N_3466,N_965,N_2845);
nor U3467 (N_3467,N_279,N_1574);
or U3468 (N_3468,N_255,N_1569);
xnor U3469 (N_3469,N_1205,N_2056);
or U3470 (N_3470,N_502,N_2301);
xor U3471 (N_3471,N_81,N_988);
or U3472 (N_3472,N_1563,N_2256);
xnor U3473 (N_3473,N_1467,N_1118);
or U3474 (N_3474,N_1430,N_2151);
or U3475 (N_3475,N_959,N_208);
and U3476 (N_3476,N_1340,N_2659);
and U3477 (N_3477,N_1701,N_789);
or U3478 (N_3478,N_2013,N_176);
and U3479 (N_3479,N_982,N_3124);
xor U3480 (N_3480,N_428,N_768);
nor U3481 (N_3481,N_2098,N_1022);
xor U3482 (N_3482,N_522,N_102);
or U3483 (N_3483,N_2749,N_1267);
and U3484 (N_3484,N_1146,N_2218);
and U3485 (N_3485,N_2855,N_3108);
nor U3486 (N_3486,N_1656,N_2741);
or U3487 (N_3487,N_2313,N_2548);
nand U3488 (N_3488,N_1615,N_2966);
and U3489 (N_3489,N_2185,N_1276);
or U3490 (N_3490,N_2641,N_634);
nand U3491 (N_3491,N_2759,N_1011);
nor U3492 (N_3492,N_1802,N_1216);
and U3493 (N_3493,N_1208,N_2651);
and U3494 (N_3494,N_2170,N_1242);
and U3495 (N_3495,N_2935,N_2216);
or U3496 (N_3496,N_2824,N_0);
or U3497 (N_3497,N_2143,N_589);
nor U3498 (N_3498,N_441,N_2228);
nand U3499 (N_3499,N_2656,N_250);
nand U3500 (N_3500,N_2713,N_448);
or U3501 (N_3501,N_1610,N_432);
or U3502 (N_3502,N_1137,N_160);
and U3503 (N_3503,N_1998,N_749);
or U3504 (N_3504,N_1461,N_1709);
nor U3505 (N_3505,N_1281,N_120);
or U3506 (N_3506,N_136,N_1637);
nand U3507 (N_3507,N_886,N_325);
xor U3508 (N_3508,N_1922,N_2562);
and U3509 (N_3509,N_2040,N_587);
xor U3510 (N_3510,N_635,N_1403);
nand U3511 (N_3511,N_1827,N_1639);
nor U3512 (N_3512,N_1872,N_650);
nor U3513 (N_3513,N_3080,N_1880);
nand U3514 (N_3514,N_2671,N_2718);
and U3515 (N_3515,N_1783,N_455);
or U3516 (N_3516,N_2787,N_31);
and U3517 (N_3517,N_1306,N_260);
or U3518 (N_3518,N_2392,N_1298);
xor U3519 (N_3519,N_387,N_599);
nand U3520 (N_3520,N_2965,N_2672);
xor U3521 (N_3521,N_453,N_1382);
xor U3522 (N_3522,N_872,N_3106);
and U3523 (N_3523,N_639,N_2495);
nand U3524 (N_3524,N_1391,N_101);
and U3525 (N_3525,N_1196,N_2160);
and U3526 (N_3526,N_1635,N_1961);
and U3527 (N_3527,N_3008,N_2799);
or U3528 (N_3528,N_1318,N_487);
nor U3529 (N_3529,N_1308,N_73);
nor U3530 (N_3530,N_2155,N_2711);
or U3531 (N_3531,N_1311,N_106);
and U3532 (N_3532,N_1407,N_825);
nand U3533 (N_3533,N_1588,N_829);
or U3534 (N_3534,N_2510,N_1084);
nor U3535 (N_3535,N_776,N_2830);
nor U3536 (N_3536,N_1659,N_2348);
or U3537 (N_3537,N_3092,N_401);
nand U3538 (N_3538,N_3033,N_2901);
nand U3539 (N_3539,N_465,N_2775);
nor U3540 (N_3540,N_1814,N_2046);
and U3541 (N_3541,N_1032,N_2831);
xor U3542 (N_3542,N_170,N_2735);
nand U3543 (N_3543,N_2587,N_489);
or U3544 (N_3544,N_2619,N_2076);
and U3545 (N_3545,N_130,N_112);
nor U3546 (N_3546,N_2790,N_1101);
and U3547 (N_3547,N_2876,N_188);
and U3548 (N_3548,N_2608,N_1114);
or U3549 (N_3549,N_2669,N_1428);
and U3550 (N_3550,N_2896,N_2750);
nor U3551 (N_3551,N_2859,N_1554);
xor U3552 (N_3552,N_273,N_491);
or U3553 (N_3553,N_2466,N_1692);
nand U3554 (N_3554,N_570,N_1969);
and U3555 (N_3555,N_1293,N_2015);
nor U3556 (N_3556,N_1879,N_1097);
nand U3557 (N_3557,N_2585,N_2700);
or U3558 (N_3558,N_3034,N_604);
xor U3559 (N_3559,N_1339,N_344);
and U3560 (N_3560,N_2358,N_2484);
nand U3561 (N_3561,N_318,N_665);
and U3562 (N_3562,N_1284,N_2760);
nor U3563 (N_3563,N_2989,N_1914);
nand U3564 (N_3564,N_1531,N_1929);
and U3565 (N_3565,N_2191,N_1634);
nand U3566 (N_3566,N_1519,N_2969);
nand U3567 (N_3567,N_901,N_2099);
or U3568 (N_3568,N_1122,N_1545);
or U3569 (N_3569,N_1406,N_2474);
and U3570 (N_3570,N_151,N_2138);
or U3571 (N_3571,N_2292,N_55);
and U3572 (N_3572,N_2379,N_62);
nand U3573 (N_3573,N_251,N_380);
nor U3574 (N_3574,N_2236,N_2227);
or U3575 (N_3575,N_1800,N_786);
nor U3576 (N_3576,N_2815,N_1838);
nand U3577 (N_3577,N_215,N_1939);
nand U3578 (N_3578,N_3076,N_2047);
nand U3579 (N_3579,N_1171,N_2215);
nor U3580 (N_3580,N_2531,N_134);
nor U3581 (N_3581,N_2082,N_2458);
and U3582 (N_3582,N_1020,N_389);
or U3583 (N_3583,N_314,N_1875);
or U3584 (N_3584,N_12,N_2984);
nand U3585 (N_3585,N_1680,N_147);
and U3586 (N_3586,N_2898,N_1512);
xnor U3587 (N_3587,N_33,N_2835);
nor U3588 (N_3588,N_1948,N_1000);
nand U3589 (N_3589,N_554,N_953);
and U3590 (N_3590,N_433,N_1050);
and U3591 (N_3591,N_1159,N_1245);
and U3592 (N_3592,N_573,N_3024);
nand U3593 (N_3593,N_1505,N_720);
nor U3594 (N_3594,N_1104,N_730);
nor U3595 (N_3595,N_2464,N_2592);
nand U3596 (N_3596,N_492,N_1850);
or U3597 (N_3597,N_2259,N_1076);
or U3598 (N_3598,N_1191,N_1087);
and U3599 (N_3599,N_474,N_937);
or U3600 (N_3600,N_2268,N_173);
and U3601 (N_3601,N_615,N_3057);
nor U3602 (N_3602,N_1154,N_1126);
and U3603 (N_3603,N_2788,N_807);
and U3604 (N_3604,N_2058,N_2967);
and U3605 (N_3605,N_1373,N_1568);
nand U3606 (N_3606,N_2983,N_2162);
and U3607 (N_3607,N_1031,N_524);
nand U3608 (N_3608,N_1524,N_2980);
and U3609 (N_3609,N_1556,N_1072);
xnor U3610 (N_3610,N_406,N_2808);
nand U3611 (N_3611,N_1991,N_1331);
xnor U3612 (N_3612,N_3063,N_2352);
nand U3613 (N_3613,N_274,N_2601);
and U3614 (N_3614,N_935,N_1143);
xnor U3615 (N_3615,N_821,N_2096);
nor U3616 (N_3616,N_1027,N_2569);
nor U3617 (N_3617,N_1973,N_2214);
nor U3618 (N_3618,N_2039,N_129);
or U3619 (N_3619,N_2528,N_3107);
or U3620 (N_3620,N_2784,N_774);
nand U3621 (N_3621,N_1453,N_1419);
nor U3622 (N_3622,N_2198,N_562);
and U3623 (N_3623,N_2920,N_1163);
xnor U3624 (N_3624,N_1984,N_2677);
nor U3625 (N_3625,N_2,N_675);
or U3626 (N_3626,N_1165,N_1422);
or U3627 (N_3627,N_143,N_2509);
nor U3628 (N_3628,N_2826,N_1711);
and U3629 (N_3629,N_2142,N_1197);
xor U3630 (N_3630,N_793,N_2834);
nand U3631 (N_3631,N_1425,N_2350);
and U3632 (N_3632,N_1156,N_1558);
nor U3633 (N_3633,N_2506,N_1001);
nand U3634 (N_3634,N_1056,N_699);
or U3635 (N_3635,N_672,N_1856);
nand U3636 (N_3636,N_2504,N_1439);
xor U3637 (N_3637,N_1520,N_1602);
nand U3638 (N_3638,N_810,N_1459);
nor U3639 (N_3639,N_1408,N_2402);
and U3640 (N_3640,N_2091,N_2158);
nor U3641 (N_3641,N_1218,N_1060);
nor U3642 (N_3642,N_2841,N_167);
xor U3643 (N_3643,N_1706,N_425);
or U3644 (N_3644,N_426,N_977);
or U3645 (N_3645,N_1110,N_199);
or U3646 (N_3646,N_1343,N_1727);
and U3647 (N_3647,N_640,N_2271);
nor U3648 (N_3648,N_10,N_423);
nand U3649 (N_3649,N_2018,N_2202);
and U3650 (N_3650,N_1623,N_1292);
nand U3651 (N_3651,N_303,N_1338);
or U3652 (N_3652,N_790,N_1405);
nand U3653 (N_3653,N_2836,N_264);
nor U3654 (N_3654,N_1313,N_2100);
nor U3655 (N_3655,N_1354,N_2195);
nor U3656 (N_3656,N_436,N_2240);
nand U3657 (N_3657,N_2449,N_299);
nor U3658 (N_3658,N_2972,N_405);
or U3659 (N_3659,N_2448,N_841);
xor U3660 (N_3660,N_1088,N_1254);
nor U3661 (N_3661,N_295,N_2148);
and U3662 (N_3662,N_2447,N_1742);
nor U3663 (N_3663,N_1795,N_2778);
or U3664 (N_3664,N_700,N_2133);
xor U3665 (N_3665,N_1793,N_439);
nand U3666 (N_3666,N_927,N_2068);
nor U3667 (N_3667,N_1642,N_201);
and U3668 (N_3668,N_2147,N_1940);
and U3669 (N_3669,N_68,N_466);
or U3670 (N_3670,N_61,N_1364);
or U3671 (N_3671,N_2792,N_1575);
and U3672 (N_3672,N_1166,N_861);
nand U3673 (N_3673,N_2126,N_1750);
and U3674 (N_3674,N_1630,N_952);
nand U3675 (N_3675,N_2706,N_1388);
nor U3676 (N_3676,N_2319,N_331);
or U3677 (N_3677,N_1931,N_658);
nand U3678 (N_3678,N_307,N_155);
or U3679 (N_3679,N_1499,N_1767);
xnor U3680 (N_3680,N_2104,N_3065);
and U3681 (N_3681,N_207,N_345);
and U3682 (N_3682,N_2593,N_1815);
nor U3683 (N_3683,N_2950,N_659);
or U3684 (N_3684,N_2776,N_2330);
nor U3685 (N_3685,N_1658,N_336);
or U3686 (N_3686,N_2237,N_2891);
nor U3687 (N_3687,N_2833,N_729);
xor U3688 (N_3688,N_2107,N_1353);
or U3689 (N_3689,N_2979,N_2182);
or U3690 (N_3690,N_115,N_895);
xor U3691 (N_3691,N_1982,N_2609);
or U3692 (N_3692,N_3036,N_2429);
and U3693 (N_3693,N_2927,N_2694);
and U3694 (N_3694,N_477,N_3009);
nand U3695 (N_3695,N_2316,N_2363);
and U3696 (N_3696,N_673,N_2384);
or U3697 (N_3697,N_740,N_583);
or U3698 (N_3698,N_2897,N_3087);
nand U3699 (N_3699,N_269,N_2632);
nand U3700 (N_3700,N_247,N_622);
nor U3701 (N_3701,N_1733,N_602);
and U3702 (N_3702,N_723,N_2771);
xor U3703 (N_3703,N_3022,N_909);
or U3704 (N_3704,N_717,N_1542);
nand U3705 (N_3705,N_668,N_1572);
nand U3706 (N_3706,N_1657,N_93);
or U3707 (N_3707,N_2648,N_2716);
nand U3708 (N_3708,N_880,N_1222);
xnor U3709 (N_3709,N_1932,N_1413);
nand U3710 (N_3710,N_3122,N_1895);
xnor U3711 (N_3711,N_983,N_1700);
nor U3712 (N_3712,N_2652,N_2812);
or U3713 (N_3713,N_1919,N_437);
nand U3714 (N_3714,N_2747,N_1307);
and U3715 (N_3715,N_799,N_2132);
or U3716 (N_3716,N_2054,N_2796);
or U3717 (N_3717,N_2059,N_773);
nor U3718 (N_3718,N_2885,N_795);
nor U3719 (N_3719,N_1317,N_1648);
and U3720 (N_3720,N_2740,N_2564);
nand U3721 (N_3721,N_788,N_1342);
nor U3722 (N_3722,N_2924,N_2244);
nand U3723 (N_3723,N_2431,N_1874);
nand U3724 (N_3724,N_1526,N_2134);
nor U3725 (N_3725,N_698,N_1018);
nor U3726 (N_3726,N_2177,N_352);
nor U3727 (N_3727,N_2274,N_1147);
and U3728 (N_3728,N_1911,N_764);
nand U3729 (N_3729,N_431,N_1530);
xor U3730 (N_3730,N_180,N_1916);
nor U3731 (N_3731,N_1893,N_2097);
nand U3732 (N_3732,N_190,N_2378);
and U3733 (N_3733,N_2478,N_1995);
and U3734 (N_3734,N_111,N_2121);
nor U3735 (N_3735,N_542,N_1100);
nand U3736 (N_3736,N_824,N_108);
nor U3737 (N_3737,N_1209,N_1679);
nor U3738 (N_3738,N_1083,N_858);
nand U3739 (N_3739,N_2217,N_1068);
nand U3740 (N_3740,N_1758,N_546);
or U3741 (N_3741,N_1044,N_2546);
or U3742 (N_3742,N_363,N_2640);
nor U3743 (N_3743,N_3045,N_2685);
and U3744 (N_3744,N_1172,N_1010);
or U3745 (N_3745,N_1045,N_71);
or U3746 (N_3746,N_1772,N_268);
nand U3747 (N_3747,N_1485,N_1959);
or U3748 (N_3748,N_1401,N_931);
nand U3749 (N_3749,N_3000,N_1805);
nor U3750 (N_3750,N_244,N_1320);
or U3751 (N_3751,N_985,N_459);
nand U3752 (N_3752,N_1039,N_721);
and U3753 (N_3753,N_1849,N_361);
nand U3754 (N_3754,N_1938,N_666);
xor U3755 (N_3755,N_2727,N_819);
and U3756 (N_3756,N_1607,N_884);
nor U3757 (N_3757,N_2071,N_2866);
and U3758 (N_3758,N_195,N_745);
nand U3759 (N_3759,N_402,N_2990);
nand U3760 (N_3760,N_1839,N_67);
or U3761 (N_3761,N_1790,N_2695);
and U3762 (N_3762,N_532,N_302);
nand U3763 (N_3763,N_1885,N_2604);
and U3764 (N_3764,N_690,N_2086);
and U3765 (N_3765,N_2175,N_2705);
and U3766 (N_3766,N_1474,N_1863);
xor U3767 (N_3767,N_1383,N_547);
nor U3768 (N_3768,N_118,N_1905);
nor U3769 (N_3769,N_777,N_942);
and U3770 (N_3770,N_2588,N_850);
nand U3771 (N_3771,N_3043,N_330);
nor U3772 (N_3772,N_2560,N_2108);
and U3773 (N_3773,N_30,N_1477);
and U3774 (N_3774,N_769,N_1350);
nor U3775 (N_3775,N_1549,N_1517);
nor U3776 (N_3776,N_1021,N_934);
nor U3777 (N_3777,N_1450,N_747);
xor U3778 (N_3778,N_912,N_1203);
nor U3779 (N_3779,N_1282,N_881);
nand U3780 (N_3780,N_815,N_1478);
nand U3781 (N_3781,N_500,N_2545);
or U3782 (N_3782,N_818,N_1968);
nand U3783 (N_3783,N_2910,N_1541);
nand U3784 (N_3784,N_1655,N_2664);
and U3785 (N_3785,N_47,N_2567);
xnor U3786 (N_3786,N_29,N_537);
nand U3787 (N_3787,N_2444,N_1584);
or U3788 (N_3788,N_2085,N_1768);
nand U3789 (N_3789,N_2493,N_686);
xor U3790 (N_3790,N_2030,N_2273);
and U3791 (N_3791,N_198,N_873);
nor U3792 (N_3792,N_920,N_24);
or U3793 (N_3793,N_2873,N_618);
xor U3794 (N_3794,N_1377,N_2272);
and U3795 (N_3795,N_2420,N_2070);
xnor U3796 (N_3796,N_2426,N_1941);
xnor U3797 (N_3797,N_2317,N_2361);
and U3798 (N_3798,N_862,N_876);
and U3799 (N_3799,N_214,N_2923);
nand U3800 (N_3800,N_1886,N_3030);
or U3801 (N_3801,N_528,N_1367);
or U3802 (N_3802,N_323,N_1440);
and U3803 (N_3803,N_1283,N_3099);
nand U3804 (N_3804,N_1883,N_1150);
nor U3805 (N_3805,N_919,N_1435);
nor U3806 (N_3806,N_1089,N_2513);
nand U3807 (N_3807,N_913,N_1232);
nand U3808 (N_3808,N_2770,N_1119);
nand U3809 (N_3809,N_1328,N_1797);
and U3810 (N_3810,N_1079,N_2491);
nor U3811 (N_3811,N_1491,N_91);
or U3812 (N_3812,N_1297,N_1550);
and U3813 (N_3813,N_1355,N_828);
nor U3814 (N_3814,N_298,N_1889);
nor U3815 (N_3815,N_1787,N_216);
or U3816 (N_3816,N_2364,N_461);
and U3817 (N_3817,N_265,N_978);
nand U3818 (N_3818,N_1500,N_1271);
or U3819 (N_3819,N_1438,N_2450);
xnor U3820 (N_3820,N_384,N_313);
or U3821 (N_3821,N_412,N_2456);
xor U3822 (N_3822,N_1404,N_1807);
nand U3823 (N_3823,N_1085,N_1092);
or U3824 (N_3824,N_2894,N_1273);
and U3825 (N_3825,N_2766,N_1059);
or U3826 (N_3826,N_2079,N_2598);
nor U3827 (N_3827,N_990,N_870);
nand U3828 (N_3828,N_468,N_2745);
nor U3829 (N_3829,N_2492,N_3004);
nand U3830 (N_3830,N_1162,N_2874);
nor U3831 (N_3831,N_240,N_333);
nand U3832 (N_3832,N_2900,N_3096);
nor U3833 (N_3833,N_1361,N_11);
xnor U3834 (N_3834,N_3105,N_359);
or U3835 (N_3835,N_2736,N_1739);
and U3836 (N_3836,N_613,N_2916);
nor U3837 (N_3837,N_2627,N_2253);
and U3838 (N_3838,N_2381,N_341);
nor U3839 (N_3839,N_2666,N_629);
nor U3840 (N_3840,N_2698,N_737);
nand U3841 (N_3841,N_2820,N_657);
nand U3842 (N_3842,N_261,N_1746);
xnor U3843 (N_3843,N_1262,N_2024);
and U3844 (N_3844,N_1037,N_1091);
and U3845 (N_3845,N_2331,N_2933);
nor U3846 (N_3846,N_2976,N_2334);
nand U3847 (N_3847,N_1920,N_294);
nor U3848 (N_3848,N_1323,N_1745);
and U3849 (N_3849,N_2786,N_286);
or U3850 (N_3850,N_2637,N_661);
nor U3851 (N_3851,N_2257,N_478);
or U3852 (N_3852,N_2798,N_899);
or U3853 (N_3853,N_1033,N_2954);
or U3854 (N_3854,N_116,N_2343);
nand U3855 (N_3855,N_1832,N_312);
or U3856 (N_3856,N_1259,N_1820);
or U3857 (N_3857,N_2179,N_293);
nand U3858 (N_3858,N_377,N_739);
nand U3859 (N_3859,N_3011,N_1892);
nor U3860 (N_3860,N_2305,N_1199);
nor U3861 (N_3861,N_1234,N_334);
or U3862 (N_3862,N_582,N_1233);
nand U3863 (N_3863,N_2926,N_2800);
nand U3864 (N_3864,N_340,N_1936);
or U3865 (N_3865,N_1884,N_2757);
and U3866 (N_3866,N_2581,N_1111);
nand U3867 (N_3867,N_2049,N_383);
nor U3868 (N_3868,N_1054,N_1016);
nand U3869 (N_3869,N_248,N_2720);
nand U3870 (N_3870,N_1730,N_2174);
and U3871 (N_3871,N_1432,N_464);
nand U3872 (N_3872,N_2416,N_2021);
xnor U3873 (N_3873,N_2925,N_1532);
or U3874 (N_3874,N_2557,N_2345);
nand U3875 (N_3875,N_2554,N_527);
or U3876 (N_3876,N_2008,N_3095);
or U3877 (N_3877,N_575,N_903);
and U3878 (N_3878,N_1702,N_597);
nand U3879 (N_3879,N_1744,N_92);
xor U3880 (N_3880,N_569,N_1304);
xnor U3881 (N_3881,N_3069,N_2114);
and U3882 (N_3882,N_1472,N_2401);
nand U3883 (N_3883,N_1460,N_391);
nor U3884 (N_3884,N_1098,N_1312);
nor U3885 (N_3885,N_802,N_2083);
and U3886 (N_3886,N_2489,N_1553);
nor U3887 (N_3887,N_2852,N_351);
nand U3888 (N_3888,N_871,N_798);
nand U3889 (N_3889,N_3082,N_760);
nand U3890 (N_3890,N_2340,N_2903);
or U3891 (N_3891,N_3016,N_2877);
nand U3892 (N_3892,N_1710,N_2200);
nor U3893 (N_3893,N_2681,N_971);
xor U3894 (N_3894,N_2821,N_280);
nor U3895 (N_3895,N_418,N_1942);
nor U3896 (N_3896,N_1057,N_791);
or U3897 (N_3897,N_2383,N_708);
and U3898 (N_3898,N_2135,N_2220);
xor U3899 (N_3899,N_2074,N_775);
nor U3900 (N_3900,N_186,N_2730);
or U3901 (N_3901,N_2277,N_419);
xor U3902 (N_3902,N_3090,N_1712);
or U3903 (N_3903,N_939,N_1633);
and U3904 (N_3904,N_2514,N_1697);
and U3905 (N_3905,N_1583,N_997);
nand U3906 (N_3906,N_39,N_2377);
and U3907 (N_3907,N_1268,N_783);
xnor U3908 (N_3908,N_2960,N_956);
or U3909 (N_3909,N_945,N_2369);
xor U3910 (N_3910,N_2643,N_2304);
nor U3911 (N_3911,N_1763,N_2782);
nand U3912 (N_3912,N_1581,N_914);
or U3913 (N_3913,N_3005,N_921);
nor U3914 (N_3914,N_2725,N_625);
and U3915 (N_3915,N_733,N_631);
xnor U3916 (N_3916,N_1606,N_2571);
nor U3917 (N_3917,N_2413,N_586);
nand U3918 (N_3918,N_2765,N_2373);
or U3919 (N_3919,N_158,N_1535);
or U3920 (N_3920,N_2322,N_2254);
or U3921 (N_3921,N_2899,N_2291);
or U3922 (N_3922,N_1481,N_1213);
nor U3923 (N_3923,N_172,N_2005);
nor U3924 (N_3924,N_2486,N_189);
nand U3925 (N_3925,N_1004,N_2682);
nor U3926 (N_3926,N_536,N_1703);
and U3927 (N_3927,N_2839,N_2505);
xnor U3928 (N_3928,N_2109,N_2696);
nor U3929 (N_3929,N_637,N_1743);
nand U3930 (N_3930,N_1887,N_1473);
and U3931 (N_3931,N_1983,N_1193);
or U3932 (N_3932,N_910,N_2995);
nand U3933 (N_3933,N_2480,N_566);
or U3934 (N_3934,N_2715,N_350);
nand U3935 (N_3935,N_297,N_1770);
or U3936 (N_3936,N_1841,N_77);
and U3937 (N_3937,N_449,N_2347);
and U3938 (N_3938,N_2410,N_671);
nor U3939 (N_3939,N_2558,N_1513);
nor U3940 (N_3940,N_1127,N_3044);
or U3941 (N_3941,N_123,N_2534);
and U3942 (N_3942,N_2201,N_1066);
and U3943 (N_3943,N_2359,N_2192);
xnor U3944 (N_3944,N_2961,N_1260);
and U3945 (N_3945,N_356,N_2805);
and U3946 (N_3946,N_2360,N_1337);
and U3947 (N_3947,N_1640,N_2710);
xnor U3948 (N_3948,N_2772,N_664);
and U3949 (N_3949,N_989,N_2403);
and U3950 (N_3950,N_1360,N_863);
nor U3951 (N_3951,N_1851,N_2675);
or U3952 (N_3952,N_2230,N_48);
or U3953 (N_3953,N_122,N_2057);
xnor U3954 (N_3954,N_59,N_16);
xor U3955 (N_3955,N_1970,N_1971);
and U3956 (N_3956,N_2958,N_1775);
nor U3957 (N_3957,N_2003,N_2971);
and U3958 (N_3958,N_1540,N_310);
and U3959 (N_3959,N_2508,N_1943);
and U3960 (N_3960,N_2613,N_3075);
or U3961 (N_3961,N_2907,N_1067);
nor U3962 (N_3962,N_812,N_2499);
nand U3963 (N_3963,N_1376,N_755);
xnor U3964 (N_3964,N_2843,N_1258);
and U3965 (N_3965,N_2663,N_879);
and U3966 (N_3966,N_1806,N_888);
xnor U3967 (N_3967,N_1766,N_918);
or U3968 (N_3968,N_1910,N_1810);
nand U3969 (N_3969,N_234,N_838);
nor U3970 (N_3970,N_25,N_1561);
and U3971 (N_3971,N_1507,N_875);
xnor U3972 (N_3972,N_2816,N_2243);
and U3973 (N_3973,N_1918,N_2573);
nor U3974 (N_3974,N_964,N_1303);
and U3975 (N_3975,N_1963,N_15);
and U3976 (N_3976,N_1823,N_1663);
or U3977 (N_3977,N_1741,N_767);
nand U3978 (N_3978,N_2642,N_125);
nor U3979 (N_3979,N_277,N_2931);
and U3980 (N_3980,N_963,N_142);
and U3981 (N_3981,N_398,N_1690);
or U3982 (N_3982,N_2748,N_864);
or U3983 (N_3983,N_152,N_2265);
nor U3984 (N_3984,N_328,N_572);
or U3985 (N_3985,N_1740,N_1206);
and U3986 (N_3986,N_2332,N_420);
nand U3987 (N_3987,N_1378,N_2346);
and U3988 (N_3988,N_378,N_135);
or U3989 (N_3989,N_1713,N_724);
nand U3990 (N_3990,N_1813,N_1608);
nand U3991 (N_3991,N_486,N_1335);
nand U3992 (N_3992,N_1506,N_1064);
nand U3993 (N_3993,N_905,N_591);
nand U3994 (N_3994,N_1236,N_2222);
and U3995 (N_3995,N_1626,N_1837);
and U3996 (N_3996,N_409,N_2851);
nand U3997 (N_3997,N_1096,N_2918);
or U3998 (N_3998,N_986,N_846);
nor U3999 (N_3999,N_1599,N_2023);
or U4000 (N_4000,N_757,N_291);
nor U4001 (N_4001,N_2282,N_2247);
xor U4002 (N_4002,N_2676,N_386);
nor U4003 (N_4003,N_1272,N_1346);
nand U4004 (N_4004,N_1774,N_2300);
nand U4005 (N_4005,N_902,N_1490);
and U4006 (N_4006,N_1960,N_3051);
nand U4007 (N_4007,N_1264,N_218);
and U4008 (N_4008,N_808,N_1564);
and U4009 (N_4009,N_2908,N_1400);
nor U4010 (N_4010,N_2275,N_954);
or U4011 (N_4011,N_1180,N_2959);
or U4012 (N_4012,N_434,N_1330);
or U4013 (N_4013,N_1627,N_620);
or U4014 (N_4014,N_373,N_966);
xor U4015 (N_4015,N_2603,N_9);
nand U4016 (N_4016,N_141,N_2398);
nand U4017 (N_4017,N_1131,N_187);
nand U4018 (N_4018,N_232,N_245);
and U4019 (N_4019,N_2144,N_1589);
nand U4020 (N_4020,N_1190,N_1112);
and U4021 (N_4021,N_476,N_2288);
or U4022 (N_4022,N_2986,N_1349);
nand U4023 (N_4023,N_689,N_2229);
or U4024 (N_4024,N_2141,N_4);
or U4025 (N_4025,N_2467,N_1651);
and U4026 (N_4026,N_2408,N_1452);
nor U4027 (N_4027,N_1475,N_581);
nand U4028 (N_4028,N_809,N_2693);
nand U4029 (N_4029,N_1344,N_1138);
nor U4030 (N_4030,N_335,N_121);
or U4031 (N_4031,N_1246,N_2789);
nand U4032 (N_4032,N_2445,N_2865);
nand U4033 (N_4033,N_1009,N_1945);
nand U4034 (N_4034,N_2169,N_649);
nor U4035 (N_4035,N_381,N_2625);
nand U4036 (N_4036,N_710,N_746);
nor U4037 (N_4037,N_1619,N_1579);
and U4038 (N_4038,N_1062,N_1736);
or U4039 (N_4039,N_1211,N_676);
nor U4040 (N_4040,N_2067,N_2342);
or U4041 (N_4041,N_538,N_719);
nor U4042 (N_4042,N_1831,N_422);
xnor U4043 (N_4043,N_1002,N_2075);
xor U4044 (N_4044,N_1130,N_628);
or U4045 (N_4045,N_457,N_519);
xor U4046 (N_4046,N_2053,N_1155);
nor U4047 (N_4047,N_309,N_332);
xor U4048 (N_4048,N_1537,N_1121);
nor U4049 (N_4049,N_1487,N_2532);
nor U4050 (N_4050,N_1981,N_1801);
nor U4051 (N_4051,N_2370,N_2527);
nor U4052 (N_4052,N_1061,N_1548);
or U4053 (N_4053,N_1479,N_1169);
nand U4054 (N_4054,N_2864,N_2081);
and U4055 (N_4055,N_944,N_209);
nand U4056 (N_4056,N_2249,N_1476);
or U4057 (N_4057,N_2551,N_2814);
nor U4058 (N_4058,N_3037,N_440);
and U4059 (N_4059,N_1124,N_709);
nor U4060 (N_4060,N_2312,N_2917);
nand U4061 (N_4061,N_1402,N_2258);
nand U4062 (N_4062,N_590,N_203);
nor U4063 (N_4063,N_2044,N_1470);
or U4064 (N_4064,N_2064,N_1161);
and U4065 (N_4065,N_2744,N_1099);
xor U4066 (N_4066,N_210,N_2267);
nor U4067 (N_4067,N_1458,N_1671);
nor U4068 (N_4068,N_1215,N_559);
nor U4069 (N_4069,N_2634,N_695);
xnor U4070 (N_4070,N_1200,N_2860);
nor U4071 (N_4071,N_2968,N_2719);
nor U4072 (N_4072,N_272,N_2512);
and U4073 (N_4073,N_1956,N_1962);
xor U4074 (N_4074,N_212,N_3023);
nor U4075 (N_4075,N_1006,N_2717);
xor U4076 (N_4076,N_60,N_1128);
or U4077 (N_4077,N_1724,N_1860);
and U4078 (N_4078,N_688,N_3019);
nand U4079 (N_4079,N_1691,N_627);
nor U4080 (N_4080,N_1444,N_1665);
and U4081 (N_4081,N_1518,N_762);
xor U4082 (N_4082,N_907,N_957);
and U4083 (N_4083,N_2911,N_2701);
nor U4084 (N_4084,N_770,N_2494);
nor U4085 (N_4085,N_2206,N_683);
and U4086 (N_4086,N_346,N_1909);
and U4087 (N_4087,N_472,N_2981);
and U4088 (N_4088,N_1675,N_2199);
nor U4089 (N_4089,N_2606,N_2544);
or U4090 (N_4090,N_1026,N_1322);
or U4091 (N_4091,N_348,N_2120);
nor U4092 (N_4092,N_771,N_97);
nand U4093 (N_4093,N_2691,N_3020);
nor U4094 (N_4094,N_1136,N_3042);
and U4095 (N_4095,N_2724,N_2339);
nor U4096 (N_4096,N_2187,N_2947);
nor U4097 (N_4097,N_2080,N_1015);
xnor U4098 (N_4098,N_1844,N_924);
and U4099 (N_4099,N_1210,N_1754);
or U4100 (N_4100,N_1177,N_551);
nor U4101 (N_4101,N_52,N_1685);
and U4102 (N_4102,N_1798,N_311);
and U4103 (N_4103,N_1255,N_679);
nor U4104 (N_4104,N_3003,N_1613);
nor U4105 (N_4105,N_2130,N_2622);
nand U4106 (N_4106,N_2605,N_6);
nor U4107 (N_4107,N_972,N_831);
and U4108 (N_4108,N_2939,N_610);
nor U4109 (N_4109,N_516,N_2435);
nor U4110 (N_4110,N_2818,N_2854);
or U4111 (N_4111,N_1081,N_2842);
or U4112 (N_4112,N_1013,N_1688);
and U4113 (N_4113,N_936,N_2653);
or U4114 (N_4114,N_1719,N_1955);
nand U4115 (N_4115,N_2597,N_2387);
and U4116 (N_4116,N_592,N_1817);
or U4117 (N_4117,N_479,N_202);
and U4118 (N_4118,N_827,N_2938);
and U4119 (N_4119,N_5,N_1571);
nor U4120 (N_4120,N_86,N_2323);
nand U4121 (N_4121,N_2172,N_213);
nand U4122 (N_4122,N_3119,N_714);
or U4123 (N_4123,N_2213,N_2357);
and U4124 (N_4124,N_928,N_2113);
nand U4125 (N_4125,N_534,N_2443);
or U4126 (N_4126,N_2211,N_1644);
nand U4127 (N_4127,N_2302,N_2507);
nor U4128 (N_4128,N_2112,N_2572);
nor U4129 (N_4129,N_399,N_521);
or U4130 (N_4130,N_1023,N_2286);
nor U4131 (N_4131,N_576,N_1878);
nor U4132 (N_4132,N_1289,N_1952);
nand U4133 (N_4133,N_707,N_1816);
or U4134 (N_4134,N_1647,N_2194);
and U4135 (N_4135,N_1341,N_1566);
or U4136 (N_4136,N_1557,N_2000);
nand U4137 (N_4137,N_430,N_2932);
and U4138 (N_4138,N_501,N_2221);
nor U4139 (N_4139,N_74,N_1762);
and U4140 (N_4140,N_1994,N_58);
or U4141 (N_4141,N_2394,N_560);
nand U4142 (N_4142,N_3013,N_2937);
nor U4143 (N_4143,N_110,N_1645);
nand U4144 (N_4144,N_183,N_843);
and U4145 (N_4145,N_1040,N_991);
nor U4146 (N_4146,N_1105,N_2459);
or U4147 (N_4147,N_713,N_2310);
nor U4148 (N_4148,N_2327,N_1829);
and U4149 (N_4149,N_2709,N_276);
or U4150 (N_4150,N_1356,N_1301);
and U4151 (N_4151,N_1622,N_2418);
or U4152 (N_4152,N_2803,N_371);
and U4153 (N_4153,N_911,N_246);
or U4154 (N_4154,N_482,N_2611);
nand U4155 (N_4155,N_2886,N_370);
nand U4156 (N_4156,N_1777,N_765);
or U4157 (N_4157,N_865,N_984);
and U4158 (N_4158,N_2620,N_2726);
or U4159 (N_4159,N_54,N_2065);
nand U4160 (N_4160,N_1985,N_2762);
nor U4161 (N_4161,N_981,N_2029);
nand U4162 (N_4162,N_1785,N_766);
nand U4163 (N_4163,N_1077,N_1748);
nor U4164 (N_4164,N_550,N_847);
or U4165 (N_4165,N_2742,N_1069);
and U4166 (N_4166,N_2583,N_1173);
or U4167 (N_4167,N_1133,N_1890);
nand U4168 (N_4168,N_2846,N_36);
and U4169 (N_4169,N_2294,N_1560);
xnor U4170 (N_4170,N_3088,N_2578);
nor U4171 (N_4171,N_2321,N_2235);
and U4172 (N_4172,N_568,N_889);
nor U4173 (N_4173,N_1725,N_254);
nand U4174 (N_4174,N_1923,N_1309);
xor U4175 (N_4175,N_1269,N_2537);
nand U4176 (N_4176,N_2173,N_1005);
or U4177 (N_4177,N_2318,N_1497);
xor U4178 (N_4178,N_2419,N_1195);
nor U4179 (N_4179,N_758,N_2045);
nand U4180 (N_4180,N_2231,N_2783);
nand U4181 (N_4181,N_1070,N_2565);
nor U4182 (N_4182,N_1869,N_520);
nand U4183 (N_4183,N_2522,N_1149);
and U4184 (N_4184,N_2779,N_2993);
nor U4185 (N_4185,N_1708,N_2801);
xor U4186 (N_4186,N_41,N_339);
nor U4187 (N_4187,N_82,N_2093);
or U4188 (N_4188,N_849,N_1362);
nand U4189 (N_4189,N_2829,N_2661);
and U4190 (N_4190,N_109,N_2425);
nor U4191 (N_4191,N_803,N_703);
nor U4192 (N_4192,N_2732,N_580);
nor U4193 (N_4193,N_3055,N_3007);
nor U4194 (N_4194,N_1502,N_3066);
or U4195 (N_4195,N_1266,N_2371);
and U4196 (N_4196,N_3014,N_1017);
xor U4197 (N_4197,N_2066,N_2806);
and U4198 (N_4198,N_513,N_867);
nand U4199 (N_4199,N_1446,N_1536);
nor U4200 (N_4200,N_3078,N_42);
nand U4201 (N_4201,N_1041,N_78);
nand U4202 (N_4202,N_1469,N_498);
or U4203 (N_4203,N_1654,N_678);
or U4204 (N_4204,N_1953,N_955);
nand U4205 (N_4205,N_545,N_79);
xor U4206 (N_4206,N_2878,N_355);
nand U4207 (N_4207,N_836,N_908);
nand U4208 (N_4208,N_1977,N_1421);
nor U4209 (N_4209,N_2471,N_228);
nand U4210 (N_4210,N_1902,N_18);
nand U4211 (N_4211,N_296,N_3071);
or U4212 (N_4212,N_485,N_778);
nor U4213 (N_4213,N_2704,N_390);
nor U4214 (N_4214,N_839,N_578);
or U4215 (N_4215,N_754,N_1508);
nand U4216 (N_4216,N_897,N_727);
or U4217 (N_4217,N_2469,N_366);
and U4218 (N_4218,N_354,N_1107);
or U4219 (N_4219,N_2945,N_2116);
nor U4220 (N_4220,N_2974,N_1257);
nor U4221 (N_4221,N_718,N_2299);
nand U4222 (N_4222,N_2407,N_1676);
nor U4223 (N_4223,N_701,N_1034);
nor U4224 (N_4224,N_1385,N_1738);
xor U4225 (N_4225,N_1274,N_404);
nor U4226 (N_4226,N_2880,N_595);
or U4227 (N_4227,N_165,N_1734);
nand U4228 (N_4228,N_2252,N_2629);
or U4229 (N_4229,N_2032,N_2038);
nor U4230 (N_4230,N_2734,N_553);
and U4231 (N_4231,N_2631,N_1456);
and U4232 (N_4232,N_2481,N_656);
or U4233 (N_4233,N_2460,N_1451);
or U4234 (N_4234,N_663,N_69);
xor U4235 (N_4235,N_2758,N_2020);
nor U4236 (N_4236,N_1437,N_259);
nand U4237 (N_4237,N_512,N_1986);
nand U4238 (N_4238,N_2296,N_2052);
or U4239 (N_4239,N_64,N_226);
xnor U4240 (N_4240,N_1603,N_925);
nand U4241 (N_4241,N_1555,N_137);
xor U4242 (N_4242,N_1036,N_1115);
and U4243 (N_4243,N_2354,N_2436);
nand U4244 (N_4244,N_2764,N_178);
nand U4245 (N_4245,N_2543,N_1449);
nor U4246 (N_4246,N_376,N_164);
and U4247 (N_4247,N_2012,N_2485);
nand U4248 (N_4248,N_416,N_1857);
and U4249 (N_4249,N_2496,N_2161);
nand U4250 (N_4250,N_1109,N_349);
nor U4251 (N_4251,N_242,N_362);
nor U4252 (N_4252,N_1811,N_1609);
or U4253 (N_4253,N_1501,N_2007);
nand U4254 (N_4254,N_2281,N_2752);
and U4255 (N_4255,N_1707,N_630);
and U4256 (N_4256,N_2680,N_1617);
nor U4257 (N_4257,N_1618,N_2017);
or U4258 (N_4258,N_2395,N_252);
xnor U4259 (N_4259,N_450,N_2043);
or U4260 (N_4260,N_2515,N_1957);
nand U4261 (N_4261,N_2586,N_308);
nor U4262 (N_4262,N_35,N_2655);
and U4263 (N_4263,N_3039,N_473);
nor U4264 (N_4264,N_1587,N_2295);
or U4265 (N_4265,N_1521,N_2382);
nand U4266 (N_4266,N_851,N_2488);
or U4267 (N_4267,N_2942,N_514);
nor U4268 (N_4268,N_1042,N_2982);
and U4269 (N_4269,N_1411,N_1168);
and U4270 (N_4270,N_243,N_2699);
and U4271 (N_4271,N_759,N_1514);
nand U4272 (N_4272,N_1174,N_1780);
and U4273 (N_4273,N_1753,N_2329);
xnor U4274 (N_4274,N_1299,N_1321);
xor U4275 (N_4275,N_667,N_206);
and U4276 (N_4276,N_1395,N_1721);
xor U4277 (N_4277,N_1224,N_205);
nand U4278 (N_4278,N_605,N_1901);
nand U4279 (N_4279,N_574,N_2122);
and U4280 (N_4280,N_3110,N_1731);
or U4281 (N_4281,N_1389,N_329);
nor U4282 (N_4282,N_315,N_1046);
or U4283 (N_4283,N_3085,N_2591);
or U4284 (N_4284,N_1843,N_470);
nand U4285 (N_4285,N_2670,N_890);
xor U4286 (N_4286,N_2838,N_1125);
nand U4287 (N_4287,N_166,N_284);
nor U4288 (N_4288,N_1625,N_2189);
nand U4289 (N_4289,N_2712,N_2362);
nand U4290 (N_4290,N_2871,N_2941);
or U4291 (N_4291,N_481,N_1759);
xnor U4292 (N_4292,N_1944,N_1263);
nand U4293 (N_4293,N_408,N_2523);
or U4294 (N_4294,N_2559,N_1225);
nor U4295 (N_4295,N_3072,N_2375);
nor U4296 (N_4296,N_2368,N_83);
or U4297 (N_4297,N_2341,N_2500);
and U4298 (N_4298,N_2890,N_1605);
and U4299 (N_4299,N_447,N_192);
and U4300 (N_4300,N_3035,N_2563);
xor U4301 (N_4301,N_742,N_577);
or U4302 (N_4302,N_2674,N_2479);
or U4303 (N_4303,N_1821,N_557);
xnor U4304 (N_4304,N_1019,N_2561);
nand U4305 (N_4305,N_2145,N_2031);
xnor U4306 (N_4306,N_1662,N_3079);
or U4307 (N_4307,N_2238,N_1735);
or U4308 (N_4308,N_813,N_411);
nor U4309 (N_4309,N_3021,N_2106);
nor U4310 (N_4310,N_1597,N_444);
or U4311 (N_4311,N_2428,N_1379);
nor U4312 (N_4312,N_2738,N_1120);
nand U4313 (N_4313,N_2163,N_2051);
nor U4314 (N_4314,N_1652,N_266);
xor U4315 (N_4315,N_235,N_1934);
nor U4316 (N_4316,N_801,N_2649);
xor U4317 (N_4317,N_194,N_140);
nor U4318 (N_4318,N_561,N_2414);
nor U4319 (N_4319,N_87,N_1882);
nor U4320 (N_4320,N_2524,N_1055);
nand U4321 (N_4321,N_1988,N_1145);
or U4322 (N_4322,N_2320,N_1523);
nor U4323 (N_4323,N_2440,N_2462);
nor U4324 (N_4324,N_2660,N_2048);
or U4325 (N_4325,N_2110,N_1366);
or U4326 (N_4326,N_2552,N_2297);
nand U4327 (N_4327,N_2270,N_1782);
nor U4328 (N_4328,N_929,N_2623);
nor U4329 (N_4329,N_3029,N_1789);
or U4330 (N_4330,N_1778,N_2856);
nand U4331 (N_4331,N_1516,N_1949);
or U4332 (N_4332,N_2164,N_652);
nor U4333 (N_4333,N_2930,N_2328);
nand U4334 (N_4334,N_645,N_2858);
and U4335 (N_4335,N_2196,N_817);
nor U4336 (N_4336,N_104,N_2881);
or U4337 (N_4337,N_2566,N_2226);
or U4338 (N_4338,N_1488,N_712);
and U4339 (N_4339,N_731,N_146);
and U4340 (N_4340,N_2152,N_2178);
nor U4341 (N_4341,N_1302,N_1103);
or U4342 (N_4342,N_2751,N_2599);
nand U4343 (N_4343,N_531,N_364);
xor U4344 (N_4344,N_1903,N_1967);
nand U4345 (N_4345,N_1431,N_2260);
or U4346 (N_4346,N_2117,N_1864);
and U4347 (N_4347,N_3111,N_249);
nor U4348 (N_4348,N_743,N_705);
nor U4349 (N_4349,N_2915,N_1214);
or U4350 (N_4350,N_1586,N_891);
and U4351 (N_4351,N_1534,N_736);
or U4352 (N_4352,N_797,N_3091);
nor U4353 (N_4353,N_1094,N_2266);
nand U4354 (N_4354,N_2405,N_3109);
nor U4355 (N_4355,N_2883,N_1202);
xor U4356 (N_4356,N_1873,N_1543);
and U4357 (N_4357,N_2600,N_617);
nor U4358 (N_4358,N_722,N_95);
and U4359 (N_4359,N_3046,N_1427);
nand U4360 (N_4360,N_1095,N_2962);
nand U4361 (N_4361,N_1351,N_2241);
xnor U4362 (N_4362,N_958,N_1935);
nor U4363 (N_4363,N_1220,N_784);
nor U4364 (N_4364,N_893,N_2612);
or U4365 (N_4365,N_1494,N_3053);
xnor U4366 (N_4366,N_270,N_3049);
and U4367 (N_4367,N_290,N_1198);
nand U4368 (N_4368,N_1862,N_1598);
nand U4369 (N_4369,N_2683,N_51);
xor U4370 (N_4370,N_2501,N_1799);
or U4371 (N_4371,N_2996,N_126);
or U4372 (N_4372,N_2219,N_1073);
nor U4373 (N_4373,N_1966,N_682);
nand U4374 (N_4374,N_3074,N_1249);
nand U4375 (N_4375,N_2223,N_1877);
nor U4376 (N_4376,N_1792,N_163);
and U4377 (N_4377,N_855,N_2234);
nor U4378 (N_4378,N_1399,N_2084);
or U4379 (N_4379,N_253,N_179);
nor U4380 (N_4380,N_1529,N_2279);
or U4381 (N_4381,N_507,N_132);
and U4382 (N_4382,N_3093,N_2584);
nand U4383 (N_4383,N_1773,N_1547);
and U4384 (N_4384,N_2547,N_1464);
or U4385 (N_4385,N_21,N_2697);
nor U4386 (N_4386,N_2521,N_1826);
nor U4387 (N_4387,N_2137,N_1223);
and U4388 (N_4388,N_1183,N_1591);
or U4389 (N_4389,N_2159,N_642);
and U4390 (N_4390,N_2437,N_2406);
xnor U4391 (N_4391,N_1078,N_869);
nand U4392 (N_4392,N_660,N_1937);
and U4393 (N_4393,N_539,N_598);
nor U4394 (N_4394,N_2804,N_2844);
nand U4395 (N_4395,N_3054,N_2819);
and U4396 (N_4396,N_263,N_1756);
xor U4397 (N_4397,N_1729,N_1393);
nor U4398 (N_4398,N_1958,N_1030);
or U4399 (N_4399,N_1980,N_579);
and U4400 (N_4400,N_1592,N_1653);
nor U4401 (N_4401,N_1888,N_998);
nor U4402 (N_4402,N_324,N_1845);
nor U4403 (N_4403,N_2457,N_2953);
or U4404 (N_4404,N_1749,N_2009);
nand U4405 (N_4405,N_1333,N_2861);
or U4406 (N_4406,N_375,N_962);
nand U4407 (N_4407,N_156,N_2579);
nor U4408 (N_4408,N_2644,N_2186);
and U4409 (N_4409,N_1788,N_1194);
xor U4410 (N_4410,N_72,N_1278);
and U4411 (N_4411,N_1852,N_191);
or U4412 (N_4412,N_1237,N_3070);
and U4413 (N_4413,N_2934,N_646);
xor U4414 (N_4414,N_2308,N_2306);
or U4415 (N_4415,N_2139,N_2813);
nand U4416 (N_4416,N_2922,N_2722);
xnor U4417 (N_4417,N_782,N_608);
xor U4418 (N_4418,N_1689,N_2985);
nand U4419 (N_4419,N_127,N_744);
xnor U4420 (N_4420,N_1722,N_2884);
nor U4421 (N_4421,N_316,N_1287);
nor U4422 (N_4422,N_2555,N_53);
and U4423 (N_4423,N_1769,N_1065);
nand U4424 (N_4424,N_393,N_1285);
xnor U4425 (N_4425,N_1142,N_968);
nor U4426 (N_4426,N_1052,N_1803);
xnor U4427 (N_4427,N_2439,N_1347);
or U4428 (N_4428,N_3060,N_806);
nand U4429 (N_4429,N_2658,N_2452);
nor U4430 (N_4430,N_2580,N_1859);
or U4431 (N_4431,N_413,N_2879);
or U4432 (N_4432,N_2264,N_2827);
nand U4433 (N_4433,N_452,N_2944);
or U4434 (N_4434,N_2333,N_2276);
or U4435 (N_4435,N_2602,N_2791);
or U4436 (N_4436,N_1904,N_2417);
or U4437 (N_4437,N_2774,N_564);
nor U4438 (N_4438,N_840,N_1515);
and U4439 (N_4439,N_558,N_814);
nand U4440 (N_4440,N_636,N_40);
and U4441 (N_4441,N_287,N_1669);
or U4442 (N_4442,N_518,N_748);
or U4443 (N_4443,N_2293,N_2746);
xnor U4444 (N_4444,N_1681,N_1947);
nand U4445 (N_4445,N_2678,N_1510);
and U4446 (N_4446,N_369,N_2539);
or U4447 (N_4447,N_2654,N_357);
nor U4448 (N_4448,N_200,N_857);
xnor U4449 (N_4449,N_571,N_365);
nor U4450 (N_4450,N_2451,N_916);
nor U4451 (N_4451,N_2203,N_1270);
and U4452 (N_4452,N_2549,N_105);
and U4453 (N_4453,N_540,N_2190);
or U4454 (N_4454,N_392,N_995);
and U4455 (N_4455,N_26,N_184);
and U4456 (N_4456,N_638,N_1509);
nor U4457 (N_4457,N_1551,N_1993);
and U4458 (N_4458,N_2438,N_1038);
or U4459 (N_4459,N_2101,N_1455);
and U4460 (N_4460,N_496,N_1008);
nor U4461 (N_4461,N_1048,N_624);
or U4462 (N_4462,N_974,N_2193);
nor U4463 (N_4463,N_1329,N_446);
or U4464 (N_4464,N_979,N_2476);
nand U4465 (N_4465,N_1327,N_1141);
nor U4466 (N_4466,N_2518,N_3025);
and U4467 (N_4467,N_1718,N_89);
or U4468 (N_4468,N_1182,N_417);
or U4469 (N_4469,N_75,N_2415);
and U4470 (N_4470,N_1380,N_2763);
or U4471 (N_4471,N_372,N_1247);
and U4472 (N_4472,N_2089,N_100);
or U4473 (N_4473,N_1310,N_1423);
xor U4474 (N_4474,N_898,N_217);
nor U4475 (N_4475,N_157,N_3081);
xor U4476 (N_4476,N_523,N_2290);
nor U4477 (N_4477,N_1965,N_1791);
nand U4478 (N_4478,N_859,N_1552);
or U4479 (N_4479,N_367,N_1429);
or U4480 (N_4480,N_951,N_611);
and U4481 (N_4481,N_1760,N_1484);
nand U4482 (N_4482,N_1755,N_1604);
nor U4483 (N_4483,N_1999,N_1720);
or U4484 (N_4484,N_3103,N_1390);
nor U4485 (N_4485,N_2019,N_641);
xnor U4486 (N_4486,N_50,N_726);
xnor U4487 (N_4487,N_2125,N_1381);
or U4488 (N_4488,N_772,N_3067);
xnor U4489 (N_4489,N_193,N_2123);
or U4490 (N_4490,N_14,N_2280);
nand U4491 (N_4491,N_1819,N_1106);
nand U4492 (N_4492,N_2781,N_1187);
nor U4493 (N_4493,N_704,N_1047);
nand U4494 (N_4494,N_76,N_2943);
or U4495 (N_4495,N_2913,N_926);
nand U4496 (N_4496,N_1672,N_1840);
nand U4497 (N_4497,N_1559,N_1632);
nand U4498 (N_4498,N_1908,N_2921);
or U4499 (N_4499,N_2366,N_976);
xnor U4500 (N_4500,N_1590,N_2146);
or U4501 (N_4501,N_2912,N_623);
nor U4502 (N_4502,N_1867,N_852);
nand U4503 (N_4503,N_2014,N_2315);
and U4504 (N_4504,N_848,N_1495);
nand U4505 (N_4505,N_1219,N_1976);
and U4506 (N_4506,N_2991,N_1641);
nor U4507 (N_4507,N_1522,N_674);
nand U4508 (N_4508,N_1972,N_621);
xor U4509 (N_4509,N_2997,N_1279);
or U4510 (N_4510,N_822,N_552);
or U4511 (N_4511,N_395,N_1348);
nor U4512 (N_4512,N_943,N_1305);
or U4513 (N_4513,N_556,N_2124);
or U4514 (N_4514,N_497,N_223);
xnor U4515 (N_4515,N_480,N_3101);
or U4516 (N_4516,N_917,N_1913);
nor U4517 (N_4517,N_1596,N_7);
nor U4518 (N_4518,N_1649,N_503);
and U4519 (N_4519,N_475,N_2807);
nor U4520 (N_4520,N_585,N_1927);
and U4521 (N_4521,N_43,N_154);
nor U4522 (N_4522,N_1043,N_2541);
or U4523 (N_4523,N_337,N_1687);
nand U4524 (N_4524,N_385,N_2400);
xor U4525 (N_4525,N_2242,N_1252);
nor U4526 (N_4526,N_594,N_2188);
xor U4527 (N_4527,N_493,N_3048);
xnor U4528 (N_4528,N_1185,N_27);
nor U4529 (N_4529,N_1809,N_2904);
or U4530 (N_4530,N_1417,N_794);
nand U4531 (N_4531,N_1871,N_1414);
nor U4532 (N_4532,N_1291,N_993);
xnor U4533 (N_4533,N_874,N_1796);
and U4534 (N_4534,N_2349,N_2434);
nand U4535 (N_4535,N_2374,N_220);
nor U4536 (N_4536,N_2150,N_647);
nand U4537 (N_4537,N_941,N_32);
nor U4538 (N_4538,N_1732,N_2737);
and U4539 (N_4539,N_1848,N_237);
nand U4540 (N_4540,N_1014,N_2978);
nand U4541 (N_4541,N_1861,N_866);
nor U4542 (N_4542,N_706,N_2688);
or U4543 (N_4543,N_2424,N_1670);
or U4544 (N_4544,N_1153,N_3031);
and U4545 (N_4545,N_301,N_1493);
nor U4546 (N_4546,N_2817,N_1139);
and U4547 (N_4547,N_2665,N_541);
or U4548 (N_4548,N_1492,N_2119);
nand U4549 (N_4549,N_1925,N_1053);
nand U4550 (N_4550,N_2001,N_169);
nor U4551 (N_4551,N_2326,N_1286);
nor U4552 (N_4552,N_2703,N_1442);
or U4553 (N_4553,N_1315,N_1628);
and U4554 (N_4554,N_600,N_462);
nor U4555 (N_4555,N_930,N_2463);
xnor U4556 (N_4556,N_1900,N_533);
and U4557 (N_4557,N_3112,N_221);
and U4558 (N_4558,N_2010,N_2848);
nor U4559 (N_4559,N_1102,N_463);
nor U4560 (N_4560,N_1565,N_2617);
or U4561 (N_4561,N_677,N_37);
or U4562 (N_4562,N_685,N_2793);
nor U4563 (N_4563,N_868,N_1229);
xor U4564 (N_4564,N_738,N_128);
nor U4565 (N_4565,N_950,N_609);
nor U4566 (N_4566,N_823,N_1170);
nand U4567 (N_4567,N_1950,N_2949);
nand U4568 (N_4568,N_2094,N_1227);
nand U4569 (N_4569,N_358,N_326);
nor U4570 (N_4570,N_2863,N_1573);
nor U4571 (N_4571,N_820,N_643);
nand U4572 (N_4572,N_225,N_3001);
and U4573 (N_4573,N_725,N_1525);
nor U4574 (N_4574,N_2033,N_1151);
or U4575 (N_4575,N_734,N_1580);
or U4576 (N_4576,N_2338,N_2335);
nor U4577 (N_4577,N_1140,N_256);
or U4578 (N_4578,N_505,N_626);
nand U4579 (N_4579,N_2919,N_57);
nor U4580 (N_4580,N_394,N_2639);
or U4581 (N_4581,N_1358,N_443);
and U4582 (N_4582,N_45,N_379);
nor U4583 (N_4583,N_456,N_3115);
and U4584 (N_4584,N_2615,N_1051);
nor U4585 (N_4585,N_133,N_2088);
nand U4586 (N_4586,N_2647,N_88);
nand U4587 (N_4587,N_2430,N_2768);
xnor U4588 (N_4588,N_2157,N_1447);
nand U4589 (N_4589,N_204,N_2423);
or U4590 (N_4590,N_2278,N_1332);
or U4591 (N_4591,N_2936,N_2393);
nand U4592 (N_4592,N_1570,N_3002);
nand U4593 (N_4593,N_360,N_469);
nor U4594 (N_4594,N_2614,N_1290);
nand U4595 (N_4595,N_2797,N_2686);
nor U4596 (N_4596,N_2412,N_1418);
nor U4597 (N_4597,N_1835,N_1243);
nand U4598 (N_4598,N_2391,N_1989);
or U4599 (N_4599,N_3047,N_1368);
or U4600 (N_4600,N_975,N_3086);
and U4601 (N_4601,N_511,N_484);
nand U4602 (N_4602,N_407,N_153);
nor U4603 (N_4603,N_321,N_1433);
nor U4604 (N_4604,N_2289,N_238);
nor U4605 (N_4605,N_1288,N_1296);
or U4606 (N_4606,N_735,N_2167);
and U4607 (N_4607,N_2536,N_1082);
xor U4608 (N_4608,N_1781,N_2063);
xor U4609 (N_4609,N_1265,N_2399);
nand U4610 (N_4610,N_1612,N_2176);
or U4611 (N_4611,N_3059,N_1594);
or U4612 (N_4612,N_3064,N_2714);
or U4613 (N_4613,N_257,N_2582);
or U4614 (N_4614,N_1717,N_2353);
and U4615 (N_4615,N_548,N_22);
and U4616 (N_4616,N_702,N_2090);
xor U4617 (N_4617,N_1674,N_2389);
and U4618 (N_4618,N_435,N_66);
nand U4619 (N_4619,N_403,N_2208);
or U4620 (N_4620,N_2773,N_2131);
nor U4621 (N_4621,N_231,N_606);
nor U4622 (N_4622,N_338,N_2888);
or U4623 (N_4623,N_3056,N_2519);
nand U4624 (N_4624,N_2224,N_687);
and U4625 (N_4625,N_2673,N_2441);
and U4626 (N_4626,N_2385,N_1158);
or U4627 (N_4627,N_584,N_2473);
nand U4628 (N_4628,N_1664,N_1371);
nor U4629 (N_4629,N_887,N_1694);
or U4630 (N_4630,N_692,N_1134);
nand U4631 (N_4631,N_2386,N_2511);
and U4632 (N_4632,N_1544,N_2072);
nand U4633 (N_4633,N_2887,N_3123);
or U4634 (N_4634,N_2311,N_1638);
and U4635 (N_4635,N_1025,N_1899);
xor U4636 (N_4636,N_948,N_1372);
and U4637 (N_4637,N_960,N_2535);
or U4638 (N_4638,N_648,N_3038);
nor U4639 (N_4639,N_2754,N_684);
nor U4640 (N_4640,N_1847,N_2616);
nand U4641 (N_4641,N_1434,N_2042);
nand U4642 (N_4642,N_2702,N_2181);
and U4643 (N_4643,N_1295,N_1751);
nor U4644 (N_4644,N_603,N_1325);
and U4645 (N_4645,N_382,N_3089);
and U4646 (N_4646,N_1319,N_1063);
xnor U4647 (N_4647,N_2287,N_2309);
nor U4648 (N_4648,N_892,N_1600);
and U4649 (N_4649,N_1482,N_2662);
nand U4650 (N_4650,N_2610,N_896);
or U4651 (N_4651,N_2520,N_3084);
or U4652 (N_4652,N_2111,N_1035);
and U4653 (N_4653,N_1661,N_607);
xnor U4654 (N_4654,N_304,N_1921);
nor U4655 (N_4655,N_421,N_1616);
nand U4656 (N_4656,N_832,N_549);
and U4657 (N_4657,N_1650,N_2847);
nand U4658 (N_4658,N_2857,N_2372);
nand U4659 (N_4659,N_2233,N_1250);
nor U4660 (N_4660,N_1964,N_3062);
nand U4661 (N_4661,N_317,N_932);
nor U4662 (N_4662,N_2708,N_1189);
nor U4663 (N_4663,N_1726,N_1907);
nor U4664 (N_4664,N_2475,N_2526);
nand U4665 (N_4665,N_2570,N_2087);
nor U4666 (N_4666,N_3073,N_2875);
and U4667 (N_4667,N_8,N_44);
nor U4668 (N_4668,N_219,N_3121);
nor U4669 (N_4669,N_728,N_601);
nor U4670 (N_4670,N_1668,N_923);
or U4671 (N_4671,N_2970,N_835);
and U4672 (N_4672,N_693,N_3113);
nand U4673 (N_4673,N_845,N_19);
or U4674 (N_4674,N_1416,N_2948);
nor U4675 (N_4675,N_1643,N_1365);
nor U4676 (N_4676,N_555,N_2957);
or U4677 (N_4677,N_1784,N_2062);
and U4678 (N_4678,N_3028,N_2542);
nor U4679 (N_4679,N_612,N_506);
xor U4680 (N_4680,N_1277,N_490);
and U4681 (N_4681,N_1090,N_1562);
nand U4682 (N_4682,N_3077,N_2621);
nand U4683 (N_4683,N_508,N_938);
xnor U4684 (N_4684,N_145,N_2753);
xnor U4685 (N_4685,N_2115,N_2011);
nor U4686 (N_4686,N_1394,N_2077);
nor U4687 (N_4687,N_1086,N_2319);
nand U4688 (N_4688,N_1032,N_1734);
nand U4689 (N_4689,N_1787,N_2648);
nor U4690 (N_4690,N_1720,N_394);
and U4691 (N_4691,N_481,N_1565);
nand U4692 (N_4692,N_2094,N_116);
or U4693 (N_4693,N_468,N_1570);
or U4694 (N_4694,N_415,N_1055);
nand U4695 (N_4695,N_2394,N_2430);
or U4696 (N_4696,N_1359,N_2623);
and U4697 (N_4697,N_300,N_40);
xnor U4698 (N_4698,N_2828,N_499);
and U4699 (N_4699,N_532,N_952);
and U4700 (N_4700,N_1630,N_382);
nor U4701 (N_4701,N_1315,N_2214);
nand U4702 (N_4702,N_2157,N_3042);
xor U4703 (N_4703,N_747,N_2706);
and U4704 (N_4704,N_1495,N_1474);
or U4705 (N_4705,N_547,N_505);
xnor U4706 (N_4706,N_1766,N_193);
or U4707 (N_4707,N_793,N_2360);
nand U4708 (N_4708,N_4,N_1923);
xor U4709 (N_4709,N_2900,N_1442);
nand U4710 (N_4710,N_1071,N_138);
nor U4711 (N_4711,N_1231,N_1374);
or U4712 (N_4712,N_2659,N_1529);
nor U4713 (N_4713,N_1917,N_10);
nor U4714 (N_4714,N_1722,N_1291);
nor U4715 (N_4715,N_557,N_3099);
or U4716 (N_4716,N_476,N_1794);
or U4717 (N_4717,N_208,N_2007);
nor U4718 (N_4718,N_1462,N_2814);
nor U4719 (N_4719,N_379,N_2876);
or U4720 (N_4720,N_1380,N_1069);
nor U4721 (N_4721,N_2348,N_1434);
and U4722 (N_4722,N_161,N_1710);
nor U4723 (N_4723,N_2536,N_2209);
and U4724 (N_4724,N_1199,N_896);
xnor U4725 (N_4725,N_2466,N_2820);
nand U4726 (N_4726,N_1363,N_304);
and U4727 (N_4727,N_653,N_1936);
and U4728 (N_4728,N_2042,N_1437);
or U4729 (N_4729,N_30,N_607);
nand U4730 (N_4730,N_1469,N_1775);
or U4731 (N_4731,N_874,N_2949);
nand U4732 (N_4732,N_1999,N_677);
nor U4733 (N_4733,N_700,N_2902);
and U4734 (N_4734,N_323,N_2983);
nand U4735 (N_4735,N_1980,N_2794);
and U4736 (N_4736,N_757,N_1071);
nand U4737 (N_4737,N_2409,N_2186);
or U4738 (N_4738,N_1034,N_823);
or U4739 (N_4739,N_2164,N_1135);
nor U4740 (N_4740,N_810,N_2574);
nor U4741 (N_4741,N_1069,N_2519);
and U4742 (N_4742,N_1034,N_1139);
nand U4743 (N_4743,N_698,N_2588);
nand U4744 (N_4744,N_0,N_106);
and U4745 (N_4745,N_1407,N_495);
or U4746 (N_4746,N_2720,N_2608);
nor U4747 (N_4747,N_597,N_466);
nand U4748 (N_4748,N_2323,N_2015);
or U4749 (N_4749,N_2436,N_1954);
nor U4750 (N_4750,N_1035,N_1728);
and U4751 (N_4751,N_2728,N_1836);
nor U4752 (N_4752,N_1555,N_668);
and U4753 (N_4753,N_984,N_1410);
or U4754 (N_4754,N_2876,N_0);
or U4755 (N_4755,N_2062,N_2369);
nor U4756 (N_4756,N_1909,N_2744);
and U4757 (N_4757,N_796,N_2939);
xor U4758 (N_4758,N_1784,N_2833);
or U4759 (N_4759,N_2669,N_972);
or U4760 (N_4760,N_2741,N_1882);
or U4761 (N_4761,N_2822,N_1932);
and U4762 (N_4762,N_573,N_2458);
xor U4763 (N_4763,N_2151,N_631);
nand U4764 (N_4764,N_2910,N_623);
nand U4765 (N_4765,N_2515,N_2102);
and U4766 (N_4766,N_373,N_1113);
and U4767 (N_4767,N_484,N_48);
nor U4768 (N_4768,N_1913,N_2379);
and U4769 (N_4769,N_1509,N_2675);
xor U4770 (N_4770,N_115,N_827);
nand U4771 (N_4771,N_1045,N_245);
xor U4772 (N_4772,N_2115,N_1468);
or U4773 (N_4773,N_1071,N_2629);
nor U4774 (N_4774,N_2605,N_2426);
and U4775 (N_4775,N_3057,N_1945);
or U4776 (N_4776,N_2658,N_366);
and U4777 (N_4777,N_2192,N_727);
or U4778 (N_4778,N_44,N_2241);
nand U4779 (N_4779,N_505,N_1502);
nand U4780 (N_4780,N_1672,N_1295);
or U4781 (N_4781,N_1921,N_211);
nor U4782 (N_4782,N_414,N_1449);
xnor U4783 (N_4783,N_3001,N_1369);
or U4784 (N_4784,N_2508,N_213);
nand U4785 (N_4785,N_1444,N_1528);
and U4786 (N_4786,N_1657,N_1478);
or U4787 (N_4787,N_2691,N_2855);
nand U4788 (N_4788,N_482,N_2604);
nor U4789 (N_4789,N_1948,N_3093);
nand U4790 (N_4790,N_2463,N_2138);
nor U4791 (N_4791,N_577,N_245);
nor U4792 (N_4792,N_515,N_2328);
or U4793 (N_4793,N_1121,N_2009);
xor U4794 (N_4794,N_2495,N_1868);
nand U4795 (N_4795,N_1644,N_329);
nor U4796 (N_4796,N_1698,N_434);
nand U4797 (N_4797,N_2990,N_1003);
nor U4798 (N_4798,N_23,N_249);
nor U4799 (N_4799,N_2912,N_1180);
nor U4800 (N_4800,N_387,N_26);
or U4801 (N_4801,N_717,N_2645);
nand U4802 (N_4802,N_2636,N_1855);
nand U4803 (N_4803,N_3005,N_2552);
or U4804 (N_4804,N_2474,N_425);
nand U4805 (N_4805,N_511,N_762);
nand U4806 (N_4806,N_900,N_645);
or U4807 (N_4807,N_502,N_1666);
nand U4808 (N_4808,N_749,N_312);
or U4809 (N_4809,N_738,N_2480);
nand U4810 (N_4810,N_1722,N_1033);
nand U4811 (N_4811,N_254,N_876);
or U4812 (N_4812,N_2129,N_2292);
or U4813 (N_4813,N_2022,N_1704);
or U4814 (N_4814,N_630,N_1950);
xor U4815 (N_4815,N_1605,N_2148);
or U4816 (N_4816,N_1781,N_519);
or U4817 (N_4817,N_1472,N_1597);
or U4818 (N_4818,N_1017,N_1042);
nand U4819 (N_4819,N_376,N_567);
nor U4820 (N_4820,N_1364,N_1000);
nor U4821 (N_4821,N_1297,N_1663);
or U4822 (N_4822,N_2310,N_561);
nand U4823 (N_4823,N_1026,N_919);
xor U4824 (N_4824,N_531,N_718);
nand U4825 (N_4825,N_138,N_1682);
xnor U4826 (N_4826,N_2091,N_451);
and U4827 (N_4827,N_920,N_2470);
or U4828 (N_4828,N_917,N_2995);
nand U4829 (N_4829,N_1485,N_920);
and U4830 (N_4830,N_2654,N_3056);
nor U4831 (N_4831,N_2689,N_1519);
or U4832 (N_4832,N_2735,N_627);
nor U4833 (N_4833,N_2256,N_689);
nor U4834 (N_4834,N_1323,N_1343);
nor U4835 (N_4835,N_2672,N_2147);
and U4836 (N_4836,N_2285,N_655);
nand U4837 (N_4837,N_2016,N_2841);
nor U4838 (N_4838,N_3033,N_2324);
or U4839 (N_4839,N_86,N_1477);
or U4840 (N_4840,N_1405,N_1240);
nand U4841 (N_4841,N_2682,N_2622);
or U4842 (N_4842,N_424,N_1368);
nor U4843 (N_4843,N_61,N_498);
or U4844 (N_4844,N_791,N_2033);
nor U4845 (N_4845,N_868,N_500);
or U4846 (N_4846,N_972,N_750);
nor U4847 (N_4847,N_874,N_2945);
and U4848 (N_4848,N_576,N_1857);
nand U4849 (N_4849,N_725,N_1247);
or U4850 (N_4850,N_75,N_2916);
or U4851 (N_4851,N_1858,N_919);
and U4852 (N_4852,N_367,N_747);
and U4853 (N_4853,N_517,N_603);
and U4854 (N_4854,N_94,N_2653);
xor U4855 (N_4855,N_1494,N_1237);
xnor U4856 (N_4856,N_376,N_1595);
or U4857 (N_4857,N_2605,N_1331);
or U4858 (N_4858,N_2509,N_1433);
nor U4859 (N_4859,N_750,N_952);
and U4860 (N_4860,N_225,N_1221);
nand U4861 (N_4861,N_595,N_599);
and U4862 (N_4862,N_2836,N_501);
xor U4863 (N_4863,N_1981,N_177);
nor U4864 (N_4864,N_2358,N_876);
and U4865 (N_4865,N_438,N_125);
or U4866 (N_4866,N_1723,N_186);
nand U4867 (N_4867,N_1137,N_2612);
nor U4868 (N_4868,N_1228,N_2425);
xnor U4869 (N_4869,N_257,N_369);
nand U4870 (N_4870,N_2823,N_688);
nand U4871 (N_4871,N_1674,N_1132);
or U4872 (N_4872,N_416,N_2074);
and U4873 (N_4873,N_2597,N_1661);
or U4874 (N_4874,N_2955,N_1136);
nor U4875 (N_4875,N_2520,N_2790);
and U4876 (N_4876,N_792,N_56);
or U4877 (N_4877,N_1147,N_2977);
nor U4878 (N_4878,N_552,N_1128);
xnor U4879 (N_4879,N_1582,N_417);
nor U4880 (N_4880,N_1116,N_2035);
nor U4881 (N_4881,N_2424,N_1978);
or U4882 (N_4882,N_2029,N_807);
and U4883 (N_4883,N_176,N_2211);
xor U4884 (N_4884,N_2261,N_1908);
nand U4885 (N_4885,N_726,N_1677);
nand U4886 (N_4886,N_2333,N_2988);
xnor U4887 (N_4887,N_1200,N_527);
and U4888 (N_4888,N_2821,N_1868);
nor U4889 (N_4889,N_1522,N_2138);
nand U4890 (N_4890,N_2299,N_698);
or U4891 (N_4891,N_980,N_1054);
nand U4892 (N_4892,N_1571,N_1793);
nor U4893 (N_4893,N_22,N_479);
nor U4894 (N_4894,N_101,N_504);
nor U4895 (N_4895,N_788,N_832);
or U4896 (N_4896,N_1931,N_381);
nor U4897 (N_4897,N_2619,N_107);
or U4898 (N_4898,N_2806,N_680);
and U4899 (N_4899,N_1755,N_2721);
xnor U4900 (N_4900,N_604,N_2276);
nand U4901 (N_4901,N_1990,N_1146);
nor U4902 (N_4902,N_1594,N_2288);
nand U4903 (N_4903,N_773,N_566);
nand U4904 (N_4904,N_802,N_2064);
or U4905 (N_4905,N_2239,N_419);
xnor U4906 (N_4906,N_1628,N_1696);
or U4907 (N_4907,N_1584,N_1900);
nor U4908 (N_4908,N_895,N_136);
xor U4909 (N_4909,N_391,N_156);
or U4910 (N_4910,N_2516,N_2631);
and U4911 (N_4911,N_2743,N_2954);
and U4912 (N_4912,N_1918,N_2393);
nor U4913 (N_4913,N_350,N_2386);
nor U4914 (N_4914,N_2449,N_755);
and U4915 (N_4915,N_1763,N_1950);
or U4916 (N_4916,N_38,N_1740);
nor U4917 (N_4917,N_1521,N_48);
and U4918 (N_4918,N_1520,N_810);
nor U4919 (N_4919,N_2136,N_921);
nor U4920 (N_4920,N_2883,N_1852);
nor U4921 (N_4921,N_1644,N_2585);
or U4922 (N_4922,N_1763,N_1729);
nor U4923 (N_4923,N_1789,N_1713);
nand U4924 (N_4924,N_747,N_2474);
nor U4925 (N_4925,N_1431,N_1563);
and U4926 (N_4926,N_2759,N_1147);
and U4927 (N_4927,N_1754,N_2804);
nand U4928 (N_4928,N_1245,N_2189);
and U4929 (N_4929,N_2100,N_1905);
or U4930 (N_4930,N_1778,N_2344);
nand U4931 (N_4931,N_2244,N_2615);
and U4932 (N_4932,N_2702,N_1153);
or U4933 (N_4933,N_2205,N_1389);
and U4934 (N_4934,N_957,N_79);
nor U4935 (N_4935,N_496,N_1554);
or U4936 (N_4936,N_78,N_2067);
or U4937 (N_4937,N_1852,N_1009);
and U4938 (N_4938,N_2753,N_2610);
nor U4939 (N_4939,N_2211,N_3115);
nor U4940 (N_4940,N_1626,N_2418);
xnor U4941 (N_4941,N_2569,N_1404);
or U4942 (N_4942,N_1313,N_1810);
and U4943 (N_4943,N_2241,N_1828);
xor U4944 (N_4944,N_2057,N_1238);
nor U4945 (N_4945,N_725,N_1900);
or U4946 (N_4946,N_703,N_3123);
nor U4947 (N_4947,N_2432,N_2339);
and U4948 (N_4948,N_574,N_580);
nor U4949 (N_4949,N_273,N_1507);
nand U4950 (N_4950,N_1895,N_1059);
and U4951 (N_4951,N_580,N_2133);
and U4952 (N_4952,N_1674,N_1294);
and U4953 (N_4953,N_554,N_2327);
nand U4954 (N_4954,N_89,N_949);
and U4955 (N_4955,N_2011,N_3);
or U4956 (N_4956,N_1421,N_1543);
and U4957 (N_4957,N_2733,N_1637);
and U4958 (N_4958,N_470,N_1174);
nor U4959 (N_4959,N_703,N_2777);
nor U4960 (N_4960,N_924,N_682);
nor U4961 (N_4961,N_1025,N_1877);
nor U4962 (N_4962,N_1601,N_2306);
or U4963 (N_4963,N_1341,N_215);
nand U4964 (N_4964,N_1368,N_1047);
and U4965 (N_4965,N_382,N_109);
nor U4966 (N_4966,N_59,N_1660);
and U4967 (N_4967,N_1258,N_1895);
nand U4968 (N_4968,N_2837,N_857);
nor U4969 (N_4969,N_2336,N_1001);
nor U4970 (N_4970,N_1433,N_92);
and U4971 (N_4971,N_1520,N_1019);
nor U4972 (N_4972,N_1550,N_1);
nor U4973 (N_4973,N_2161,N_2181);
nor U4974 (N_4974,N_1742,N_2679);
nand U4975 (N_4975,N_3,N_1667);
nand U4976 (N_4976,N_949,N_1067);
nor U4977 (N_4977,N_3092,N_2477);
or U4978 (N_4978,N_605,N_2901);
or U4979 (N_4979,N_876,N_2248);
nor U4980 (N_4980,N_1691,N_87);
and U4981 (N_4981,N_1793,N_138);
or U4982 (N_4982,N_301,N_2799);
nand U4983 (N_4983,N_2989,N_354);
nor U4984 (N_4984,N_1011,N_841);
and U4985 (N_4985,N_2220,N_794);
or U4986 (N_4986,N_1792,N_159);
nand U4987 (N_4987,N_267,N_2847);
nand U4988 (N_4988,N_767,N_1170);
nand U4989 (N_4989,N_1133,N_901);
or U4990 (N_4990,N_2620,N_2658);
and U4991 (N_4991,N_1095,N_2189);
and U4992 (N_4992,N_1011,N_3028);
and U4993 (N_4993,N_1043,N_718);
or U4994 (N_4994,N_1139,N_240);
nand U4995 (N_4995,N_2736,N_1020);
xnor U4996 (N_4996,N_893,N_90);
nand U4997 (N_4997,N_2621,N_178);
and U4998 (N_4998,N_1980,N_3111);
nand U4999 (N_4999,N_2152,N_2938);
nand U5000 (N_5000,N_1925,N_493);
nand U5001 (N_5001,N_847,N_250);
nor U5002 (N_5002,N_2097,N_1083);
and U5003 (N_5003,N_2161,N_1306);
or U5004 (N_5004,N_1548,N_444);
nand U5005 (N_5005,N_2134,N_2106);
or U5006 (N_5006,N_961,N_1306);
and U5007 (N_5007,N_901,N_2927);
xor U5008 (N_5008,N_1227,N_2699);
nor U5009 (N_5009,N_3044,N_1789);
nand U5010 (N_5010,N_2381,N_1596);
nor U5011 (N_5011,N_1118,N_1398);
or U5012 (N_5012,N_1441,N_627);
or U5013 (N_5013,N_781,N_809);
nand U5014 (N_5014,N_1591,N_2511);
or U5015 (N_5015,N_2310,N_347);
nor U5016 (N_5016,N_148,N_2877);
nand U5017 (N_5017,N_301,N_509);
nor U5018 (N_5018,N_3017,N_1302);
nor U5019 (N_5019,N_760,N_1005);
xnor U5020 (N_5020,N_1779,N_1848);
or U5021 (N_5021,N_2468,N_2677);
nand U5022 (N_5022,N_3069,N_1732);
and U5023 (N_5023,N_1463,N_1263);
and U5024 (N_5024,N_2000,N_618);
nor U5025 (N_5025,N_124,N_23);
nor U5026 (N_5026,N_1917,N_1173);
nor U5027 (N_5027,N_964,N_2814);
or U5028 (N_5028,N_1852,N_604);
nand U5029 (N_5029,N_1109,N_2144);
or U5030 (N_5030,N_1598,N_702);
and U5031 (N_5031,N_1162,N_1016);
xnor U5032 (N_5032,N_1076,N_157);
and U5033 (N_5033,N_1960,N_872);
nand U5034 (N_5034,N_1116,N_51);
xnor U5035 (N_5035,N_2699,N_685);
nand U5036 (N_5036,N_859,N_596);
nand U5037 (N_5037,N_1444,N_1989);
nand U5038 (N_5038,N_2213,N_1038);
xnor U5039 (N_5039,N_2071,N_1157);
and U5040 (N_5040,N_1791,N_395);
or U5041 (N_5041,N_784,N_1484);
and U5042 (N_5042,N_2638,N_1301);
xnor U5043 (N_5043,N_1719,N_1381);
and U5044 (N_5044,N_1801,N_2039);
or U5045 (N_5045,N_746,N_3031);
nor U5046 (N_5046,N_2060,N_2764);
nand U5047 (N_5047,N_1659,N_755);
or U5048 (N_5048,N_211,N_205);
or U5049 (N_5049,N_1845,N_2176);
xnor U5050 (N_5050,N_293,N_938);
nand U5051 (N_5051,N_2792,N_361);
nor U5052 (N_5052,N_2525,N_1737);
nand U5053 (N_5053,N_2590,N_2605);
or U5054 (N_5054,N_3011,N_2861);
nand U5055 (N_5055,N_64,N_2584);
and U5056 (N_5056,N_2084,N_917);
nor U5057 (N_5057,N_580,N_1878);
or U5058 (N_5058,N_2437,N_1549);
and U5059 (N_5059,N_988,N_645);
and U5060 (N_5060,N_2696,N_830);
and U5061 (N_5061,N_1967,N_956);
nand U5062 (N_5062,N_2064,N_2341);
nor U5063 (N_5063,N_800,N_1945);
nand U5064 (N_5064,N_643,N_2922);
nor U5065 (N_5065,N_1562,N_618);
or U5066 (N_5066,N_2641,N_1199);
and U5067 (N_5067,N_2949,N_977);
or U5068 (N_5068,N_787,N_324);
nor U5069 (N_5069,N_1238,N_822);
xnor U5070 (N_5070,N_2414,N_2025);
nand U5071 (N_5071,N_1080,N_1009);
xor U5072 (N_5072,N_2163,N_252);
nor U5073 (N_5073,N_524,N_2464);
and U5074 (N_5074,N_7,N_3007);
nor U5075 (N_5075,N_816,N_2823);
and U5076 (N_5076,N_1672,N_651);
xor U5077 (N_5077,N_2336,N_1612);
nor U5078 (N_5078,N_1676,N_442);
or U5079 (N_5079,N_2939,N_2640);
nor U5080 (N_5080,N_3108,N_1668);
and U5081 (N_5081,N_2654,N_2246);
or U5082 (N_5082,N_2403,N_63);
nand U5083 (N_5083,N_232,N_2708);
nand U5084 (N_5084,N_913,N_2043);
nand U5085 (N_5085,N_1048,N_2249);
or U5086 (N_5086,N_2644,N_1842);
xnor U5087 (N_5087,N_2629,N_2785);
nand U5088 (N_5088,N_977,N_2603);
nor U5089 (N_5089,N_1159,N_1840);
or U5090 (N_5090,N_1434,N_131);
and U5091 (N_5091,N_319,N_1244);
and U5092 (N_5092,N_307,N_358);
or U5093 (N_5093,N_895,N_1771);
and U5094 (N_5094,N_673,N_2490);
and U5095 (N_5095,N_274,N_2520);
and U5096 (N_5096,N_22,N_107);
or U5097 (N_5097,N_2668,N_3010);
nor U5098 (N_5098,N_945,N_2764);
or U5099 (N_5099,N_1714,N_2017);
or U5100 (N_5100,N_359,N_2171);
nand U5101 (N_5101,N_814,N_1738);
nand U5102 (N_5102,N_628,N_1426);
nand U5103 (N_5103,N_1076,N_950);
nand U5104 (N_5104,N_1945,N_826);
nor U5105 (N_5105,N_2419,N_424);
xor U5106 (N_5106,N_2440,N_878);
xor U5107 (N_5107,N_2838,N_418);
and U5108 (N_5108,N_1433,N_77);
nor U5109 (N_5109,N_2112,N_2873);
nand U5110 (N_5110,N_604,N_1912);
nor U5111 (N_5111,N_2360,N_2881);
and U5112 (N_5112,N_217,N_885);
and U5113 (N_5113,N_3047,N_3027);
or U5114 (N_5114,N_664,N_920);
nor U5115 (N_5115,N_528,N_922);
or U5116 (N_5116,N_352,N_1676);
xor U5117 (N_5117,N_1962,N_1007);
or U5118 (N_5118,N_428,N_2421);
or U5119 (N_5119,N_1929,N_2587);
or U5120 (N_5120,N_2762,N_2519);
nand U5121 (N_5121,N_2566,N_2637);
or U5122 (N_5122,N_2541,N_3075);
nor U5123 (N_5123,N_2308,N_911);
and U5124 (N_5124,N_2089,N_3086);
nand U5125 (N_5125,N_2574,N_1164);
or U5126 (N_5126,N_1657,N_2918);
or U5127 (N_5127,N_1474,N_1589);
nand U5128 (N_5128,N_2621,N_106);
nor U5129 (N_5129,N_2977,N_1767);
nor U5130 (N_5130,N_834,N_951);
or U5131 (N_5131,N_1560,N_2011);
or U5132 (N_5132,N_1048,N_109);
and U5133 (N_5133,N_1545,N_2428);
or U5134 (N_5134,N_2414,N_2703);
nor U5135 (N_5135,N_1241,N_1830);
xor U5136 (N_5136,N_2730,N_1436);
nand U5137 (N_5137,N_1246,N_2660);
nor U5138 (N_5138,N_960,N_1062);
and U5139 (N_5139,N_667,N_682);
and U5140 (N_5140,N_2873,N_631);
nor U5141 (N_5141,N_2172,N_1781);
nor U5142 (N_5142,N_186,N_1558);
and U5143 (N_5143,N_79,N_317);
xor U5144 (N_5144,N_695,N_1503);
xor U5145 (N_5145,N_1084,N_1596);
or U5146 (N_5146,N_751,N_2881);
nand U5147 (N_5147,N_1000,N_223);
xnor U5148 (N_5148,N_1767,N_1359);
nand U5149 (N_5149,N_978,N_2587);
and U5150 (N_5150,N_1982,N_2574);
nand U5151 (N_5151,N_1043,N_647);
nor U5152 (N_5152,N_2810,N_2979);
nor U5153 (N_5153,N_918,N_277);
and U5154 (N_5154,N_343,N_322);
nor U5155 (N_5155,N_544,N_1886);
nor U5156 (N_5156,N_2419,N_968);
or U5157 (N_5157,N_2970,N_1762);
xnor U5158 (N_5158,N_2365,N_39);
or U5159 (N_5159,N_2967,N_375);
or U5160 (N_5160,N_891,N_1479);
nand U5161 (N_5161,N_2071,N_585);
nand U5162 (N_5162,N_1816,N_1841);
and U5163 (N_5163,N_453,N_678);
nand U5164 (N_5164,N_2829,N_2786);
nor U5165 (N_5165,N_2893,N_2626);
or U5166 (N_5166,N_1130,N_2977);
or U5167 (N_5167,N_1044,N_596);
xnor U5168 (N_5168,N_258,N_240);
nor U5169 (N_5169,N_3027,N_1418);
nor U5170 (N_5170,N_2973,N_2122);
nor U5171 (N_5171,N_1355,N_2669);
nand U5172 (N_5172,N_2837,N_2909);
nor U5173 (N_5173,N_2230,N_76);
or U5174 (N_5174,N_2738,N_30);
nand U5175 (N_5175,N_2788,N_2696);
nand U5176 (N_5176,N_2634,N_2246);
nor U5177 (N_5177,N_1394,N_2168);
nor U5178 (N_5178,N_3026,N_1936);
and U5179 (N_5179,N_839,N_708);
and U5180 (N_5180,N_1564,N_2355);
nor U5181 (N_5181,N_2075,N_2092);
or U5182 (N_5182,N_2870,N_69);
nand U5183 (N_5183,N_3044,N_2772);
nand U5184 (N_5184,N_1632,N_571);
or U5185 (N_5185,N_3001,N_1900);
or U5186 (N_5186,N_1765,N_346);
nand U5187 (N_5187,N_585,N_1234);
nor U5188 (N_5188,N_978,N_1760);
nand U5189 (N_5189,N_2893,N_2941);
or U5190 (N_5190,N_2847,N_203);
nand U5191 (N_5191,N_1582,N_1649);
and U5192 (N_5192,N_1356,N_1957);
nand U5193 (N_5193,N_2604,N_2836);
nor U5194 (N_5194,N_432,N_2121);
or U5195 (N_5195,N_1198,N_1667);
nor U5196 (N_5196,N_2041,N_1975);
or U5197 (N_5197,N_2840,N_376);
nor U5198 (N_5198,N_138,N_2596);
nand U5199 (N_5199,N_2236,N_2067);
or U5200 (N_5200,N_67,N_2043);
xor U5201 (N_5201,N_217,N_1567);
nand U5202 (N_5202,N_2149,N_406);
nor U5203 (N_5203,N_1628,N_144);
nand U5204 (N_5204,N_2797,N_1896);
nand U5205 (N_5205,N_485,N_180);
nor U5206 (N_5206,N_561,N_270);
or U5207 (N_5207,N_846,N_395);
and U5208 (N_5208,N_2164,N_2217);
nor U5209 (N_5209,N_2883,N_575);
and U5210 (N_5210,N_2023,N_1888);
nor U5211 (N_5211,N_1812,N_1529);
or U5212 (N_5212,N_1055,N_1121);
and U5213 (N_5213,N_2114,N_1308);
nor U5214 (N_5214,N_580,N_117);
or U5215 (N_5215,N_682,N_1705);
nor U5216 (N_5216,N_1071,N_437);
or U5217 (N_5217,N_1628,N_223);
nor U5218 (N_5218,N_2779,N_1857);
nor U5219 (N_5219,N_2295,N_1808);
nor U5220 (N_5220,N_2737,N_1682);
and U5221 (N_5221,N_2453,N_3055);
and U5222 (N_5222,N_2805,N_2527);
nand U5223 (N_5223,N_1343,N_1855);
and U5224 (N_5224,N_2644,N_401);
nor U5225 (N_5225,N_1172,N_342);
xnor U5226 (N_5226,N_2190,N_2798);
nor U5227 (N_5227,N_1694,N_1945);
nor U5228 (N_5228,N_3032,N_2446);
nor U5229 (N_5229,N_1106,N_3036);
nand U5230 (N_5230,N_3016,N_1271);
nand U5231 (N_5231,N_17,N_1068);
or U5232 (N_5232,N_2481,N_2534);
and U5233 (N_5233,N_907,N_1966);
nand U5234 (N_5234,N_1191,N_2735);
nor U5235 (N_5235,N_306,N_1983);
or U5236 (N_5236,N_382,N_2589);
and U5237 (N_5237,N_2167,N_1028);
and U5238 (N_5238,N_1123,N_2855);
and U5239 (N_5239,N_2512,N_2534);
nand U5240 (N_5240,N_745,N_1425);
or U5241 (N_5241,N_2944,N_2749);
nor U5242 (N_5242,N_2562,N_1016);
or U5243 (N_5243,N_212,N_1174);
or U5244 (N_5244,N_1428,N_328);
or U5245 (N_5245,N_360,N_331);
nand U5246 (N_5246,N_767,N_1069);
xnor U5247 (N_5247,N_776,N_2691);
nand U5248 (N_5248,N_2667,N_2641);
or U5249 (N_5249,N_2229,N_2269);
nor U5250 (N_5250,N_1019,N_1169);
xor U5251 (N_5251,N_511,N_1694);
or U5252 (N_5252,N_322,N_772);
or U5253 (N_5253,N_178,N_257);
xnor U5254 (N_5254,N_3007,N_296);
or U5255 (N_5255,N_1909,N_1394);
and U5256 (N_5256,N_2451,N_1263);
nand U5257 (N_5257,N_2273,N_2987);
nor U5258 (N_5258,N_1041,N_1400);
nor U5259 (N_5259,N_2690,N_711);
or U5260 (N_5260,N_200,N_1181);
or U5261 (N_5261,N_1045,N_1465);
or U5262 (N_5262,N_1971,N_687);
and U5263 (N_5263,N_1527,N_2132);
nand U5264 (N_5264,N_294,N_1793);
nor U5265 (N_5265,N_1559,N_518);
and U5266 (N_5266,N_1223,N_171);
or U5267 (N_5267,N_17,N_2091);
nor U5268 (N_5268,N_577,N_255);
nand U5269 (N_5269,N_1700,N_2465);
nor U5270 (N_5270,N_2531,N_2324);
nand U5271 (N_5271,N_297,N_2143);
and U5272 (N_5272,N_509,N_1798);
and U5273 (N_5273,N_1748,N_1261);
nand U5274 (N_5274,N_653,N_2956);
nand U5275 (N_5275,N_305,N_74);
nor U5276 (N_5276,N_1724,N_272);
or U5277 (N_5277,N_1918,N_2655);
or U5278 (N_5278,N_3115,N_2545);
or U5279 (N_5279,N_1617,N_763);
xnor U5280 (N_5280,N_153,N_1694);
and U5281 (N_5281,N_1619,N_2302);
nand U5282 (N_5282,N_1562,N_284);
nand U5283 (N_5283,N_2738,N_2016);
and U5284 (N_5284,N_2359,N_410);
nor U5285 (N_5285,N_2333,N_2873);
nand U5286 (N_5286,N_520,N_983);
or U5287 (N_5287,N_664,N_691);
and U5288 (N_5288,N_1916,N_3110);
xor U5289 (N_5289,N_2533,N_991);
xor U5290 (N_5290,N_55,N_409);
nor U5291 (N_5291,N_223,N_137);
nor U5292 (N_5292,N_39,N_357);
xnor U5293 (N_5293,N_978,N_338);
and U5294 (N_5294,N_484,N_725);
nand U5295 (N_5295,N_1267,N_1274);
and U5296 (N_5296,N_1838,N_940);
nand U5297 (N_5297,N_1586,N_760);
and U5298 (N_5298,N_746,N_1684);
or U5299 (N_5299,N_2803,N_3019);
nand U5300 (N_5300,N_1240,N_1510);
and U5301 (N_5301,N_1171,N_1560);
xor U5302 (N_5302,N_229,N_1332);
nand U5303 (N_5303,N_2433,N_2567);
or U5304 (N_5304,N_3098,N_2474);
nor U5305 (N_5305,N_2609,N_682);
or U5306 (N_5306,N_1476,N_1250);
and U5307 (N_5307,N_1764,N_2440);
or U5308 (N_5308,N_60,N_1189);
nand U5309 (N_5309,N_2072,N_1757);
nand U5310 (N_5310,N_1666,N_2529);
nand U5311 (N_5311,N_2749,N_2016);
nor U5312 (N_5312,N_2729,N_723);
and U5313 (N_5313,N_2457,N_1444);
nand U5314 (N_5314,N_2584,N_1047);
or U5315 (N_5315,N_1543,N_2269);
or U5316 (N_5316,N_750,N_1664);
or U5317 (N_5317,N_2655,N_2002);
xor U5318 (N_5318,N_2122,N_1490);
and U5319 (N_5319,N_2820,N_208);
and U5320 (N_5320,N_2923,N_658);
or U5321 (N_5321,N_1996,N_3024);
and U5322 (N_5322,N_2434,N_2105);
and U5323 (N_5323,N_1733,N_817);
nor U5324 (N_5324,N_2549,N_2622);
and U5325 (N_5325,N_2975,N_28);
or U5326 (N_5326,N_475,N_3033);
nor U5327 (N_5327,N_1731,N_2859);
or U5328 (N_5328,N_2832,N_2248);
nor U5329 (N_5329,N_181,N_2976);
xnor U5330 (N_5330,N_2527,N_1963);
or U5331 (N_5331,N_1,N_1508);
nand U5332 (N_5332,N_1766,N_3002);
nor U5333 (N_5333,N_474,N_670);
or U5334 (N_5334,N_2183,N_89);
nor U5335 (N_5335,N_3103,N_81);
nor U5336 (N_5336,N_2563,N_1092);
nand U5337 (N_5337,N_1392,N_2547);
xor U5338 (N_5338,N_2723,N_2885);
nor U5339 (N_5339,N_3053,N_2234);
nor U5340 (N_5340,N_764,N_803);
or U5341 (N_5341,N_1311,N_1360);
or U5342 (N_5342,N_828,N_637);
nor U5343 (N_5343,N_993,N_1252);
nand U5344 (N_5344,N_2653,N_1292);
or U5345 (N_5345,N_1138,N_2297);
nor U5346 (N_5346,N_333,N_319);
xnor U5347 (N_5347,N_1106,N_900);
nand U5348 (N_5348,N_2179,N_269);
and U5349 (N_5349,N_2633,N_3032);
and U5350 (N_5350,N_827,N_19);
xor U5351 (N_5351,N_3037,N_2214);
or U5352 (N_5352,N_2190,N_2154);
nand U5353 (N_5353,N_600,N_828);
nand U5354 (N_5354,N_1366,N_2256);
xor U5355 (N_5355,N_490,N_1098);
nor U5356 (N_5356,N_763,N_1059);
and U5357 (N_5357,N_1308,N_456);
or U5358 (N_5358,N_2022,N_23);
or U5359 (N_5359,N_2167,N_1994);
nand U5360 (N_5360,N_448,N_2809);
and U5361 (N_5361,N_2044,N_203);
or U5362 (N_5362,N_396,N_2692);
or U5363 (N_5363,N_2858,N_1920);
nor U5364 (N_5364,N_1905,N_593);
nand U5365 (N_5365,N_1253,N_1100);
nor U5366 (N_5366,N_2935,N_2237);
or U5367 (N_5367,N_914,N_2257);
nand U5368 (N_5368,N_2366,N_1412);
or U5369 (N_5369,N_2279,N_2629);
or U5370 (N_5370,N_2730,N_1924);
or U5371 (N_5371,N_2642,N_1116);
nor U5372 (N_5372,N_2399,N_164);
nor U5373 (N_5373,N_1431,N_1907);
or U5374 (N_5374,N_1826,N_2629);
or U5375 (N_5375,N_2989,N_864);
nor U5376 (N_5376,N_1265,N_1349);
and U5377 (N_5377,N_979,N_2256);
nand U5378 (N_5378,N_1084,N_642);
or U5379 (N_5379,N_1616,N_947);
nand U5380 (N_5380,N_2439,N_1983);
and U5381 (N_5381,N_1608,N_519);
xnor U5382 (N_5382,N_1149,N_2921);
nand U5383 (N_5383,N_716,N_1308);
nor U5384 (N_5384,N_21,N_26);
nand U5385 (N_5385,N_2860,N_1256);
or U5386 (N_5386,N_1365,N_2548);
nand U5387 (N_5387,N_2170,N_1108);
nor U5388 (N_5388,N_309,N_190);
nand U5389 (N_5389,N_923,N_1131);
nand U5390 (N_5390,N_1241,N_416);
nand U5391 (N_5391,N_2190,N_2433);
nor U5392 (N_5392,N_983,N_1599);
and U5393 (N_5393,N_16,N_1795);
or U5394 (N_5394,N_245,N_2872);
nand U5395 (N_5395,N_2141,N_175);
or U5396 (N_5396,N_3027,N_1706);
nand U5397 (N_5397,N_594,N_3078);
nor U5398 (N_5398,N_309,N_843);
nor U5399 (N_5399,N_957,N_44);
or U5400 (N_5400,N_669,N_1622);
nor U5401 (N_5401,N_2721,N_146);
nor U5402 (N_5402,N_2764,N_2268);
and U5403 (N_5403,N_473,N_1616);
or U5404 (N_5404,N_1014,N_2997);
or U5405 (N_5405,N_2087,N_362);
nor U5406 (N_5406,N_2423,N_244);
nor U5407 (N_5407,N_2254,N_2800);
or U5408 (N_5408,N_2079,N_2469);
nand U5409 (N_5409,N_68,N_2586);
and U5410 (N_5410,N_1629,N_262);
nand U5411 (N_5411,N_135,N_1865);
xor U5412 (N_5412,N_264,N_228);
nand U5413 (N_5413,N_881,N_1898);
nor U5414 (N_5414,N_275,N_2506);
nand U5415 (N_5415,N_830,N_1573);
or U5416 (N_5416,N_737,N_2335);
or U5417 (N_5417,N_1827,N_1702);
and U5418 (N_5418,N_406,N_2141);
xor U5419 (N_5419,N_2763,N_538);
or U5420 (N_5420,N_367,N_815);
and U5421 (N_5421,N_1946,N_1351);
nand U5422 (N_5422,N_296,N_1058);
or U5423 (N_5423,N_2761,N_332);
and U5424 (N_5424,N_880,N_909);
nand U5425 (N_5425,N_2777,N_1016);
or U5426 (N_5426,N_2096,N_2564);
nor U5427 (N_5427,N_578,N_1823);
nand U5428 (N_5428,N_2793,N_2390);
and U5429 (N_5429,N_639,N_2581);
or U5430 (N_5430,N_2537,N_1061);
xnor U5431 (N_5431,N_2443,N_1141);
and U5432 (N_5432,N_1644,N_2049);
nand U5433 (N_5433,N_929,N_392);
or U5434 (N_5434,N_2210,N_1473);
nor U5435 (N_5435,N_2915,N_2165);
and U5436 (N_5436,N_82,N_24);
nor U5437 (N_5437,N_3116,N_509);
nor U5438 (N_5438,N_904,N_2839);
nor U5439 (N_5439,N_2711,N_2699);
nor U5440 (N_5440,N_1692,N_2755);
and U5441 (N_5441,N_2146,N_529);
nor U5442 (N_5442,N_261,N_2745);
and U5443 (N_5443,N_2277,N_2139);
or U5444 (N_5444,N_2425,N_343);
xor U5445 (N_5445,N_1235,N_2201);
nand U5446 (N_5446,N_2047,N_405);
and U5447 (N_5447,N_1943,N_344);
nor U5448 (N_5448,N_149,N_1183);
or U5449 (N_5449,N_448,N_1191);
nor U5450 (N_5450,N_2260,N_2354);
and U5451 (N_5451,N_2780,N_1749);
xnor U5452 (N_5452,N_2357,N_400);
nor U5453 (N_5453,N_2462,N_935);
nor U5454 (N_5454,N_1625,N_41);
xor U5455 (N_5455,N_2525,N_2321);
and U5456 (N_5456,N_2052,N_1389);
nor U5457 (N_5457,N_1032,N_2696);
nor U5458 (N_5458,N_2135,N_971);
or U5459 (N_5459,N_2572,N_2851);
nor U5460 (N_5460,N_953,N_1030);
or U5461 (N_5461,N_2096,N_3081);
nand U5462 (N_5462,N_929,N_682);
or U5463 (N_5463,N_1657,N_929);
nor U5464 (N_5464,N_2012,N_1937);
xor U5465 (N_5465,N_1412,N_3004);
nand U5466 (N_5466,N_3057,N_2867);
or U5467 (N_5467,N_923,N_479);
nor U5468 (N_5468,N_95,N_2625);
nor U5469 (N_5469,N_1964,N_1245);
and U5470 (N_5470,N_2050,N_2558);
or U5471 (N_5471,N_2438,N_666);
or U5472 (N_5472,N_567,N_1497);
nand U5473 (N_5473,N_2973,N_577);
and U5474 (N_5474,N_2568,N_208);
nor U5475 (N_5475,N_1242,N_2867);
nand U5476 (N_5476,N_3095,N_2026);
and U5477 (N_5477,N_945,N_2508);
nand U5478 (N_5478,N_2443,N_286);
nor U5479 (N_5479,N_739,N_46);
nand U5480 (N_5480,N_2231,N_726);
xor U5481 (N_5481,N_791,N_1270);
nand U5482 (N_5482,N_2209,N_722);
and U5483 (N_5483,N_184,N_2733);
nand U5484 (N_5484,N_1755,N_1464);
or U5485 (N_5485,N_1989,N_2231);
or U5486 (N_5486,N_3004,N_3045);
nand U5487 (N_5487,N_1032,N_476);
nand U5488 (N_5488,N_2338,N_852);
and U5489 (N_5489,N_311,N_2278);
or U5490 (N_5490,N_591,N_566);
xor U5491 (N_5491,N_2073,N_2082);
nor U5492 (N_5492,N_1687,N_747);
or U5493 (N_5493,N_3014,N_657);
or U5494 (N_5494,N_1776,N_3058);
nand U5495 (N_5495,N_666,N_1180);
nor U5496 (N_5496,N_773,N_1211);
and U5497 (N_5497,N_2978,N_1577);
and U5498 (N_5498,N_52,N_331);
nand U5499 (N_5499,N_2572,N_1284);
nor U5500 (N_5500,N_627,N_1678);
and U5501 (N_5501,N_535,N_629);
nand U5502 (N_5502,N_2561,N_663);
or U5503 (N_5503,N_207,N_2789);
and U5504 (N_5504,N_1223,N_1854);
or U5505 (N_5505,N_701,N_1140);
nand U5506 (N_5506,N_500,N_2392);
nand U5507 (N_5507,N_2133,N_198);
or U5508 (N_5508,N_2890,N_2660);
or U5509 (N_5509,N_2348,N_1444);
nor U5510 (N_5510,N_2478,N_313);
or U5511 (N_5511,N_2304,N_2494);
or U5512 (N_5512,N_1864,N_1438);
and U5513 (N_5513,N_1024,N_1702);
nor U5514 (N_5514,N_2572,N_1020);
or U5515 (N_5515,N_328,N_2249);
nor U5516 (N_5516,N_2431,N_2486);
and U5517 (N_5517,N_485,N_2103);
and U5518 (N_5518,N_2528,N_2744);
or U5519 (N_5519,N_1673,N_799);
or U5520 (N_5520,N_1692,N_1712);
nor U5521 (N_5521,N_1303,N_313);
nor U5522 (N_5522,N_640,N_2883);
or U5523 (N_5523,N_1160,N_1893);
or U5524 (N_5524,N_1582,N_1418);
nand U5525 (N_5525,N_341,N_2663);
nand U5526 (N_5526,N_2746,N_461);
nor U5527 (N_5527,N_361,N_2068);
nor U5528 (N_5528,N_368,N_2465);
or U5529 (N_5529,N_2942,N_2814);
nor U5530 (N_5530,N_1766,N_629);
nor U5531 (N_5531,N_2595,N_1683);
nor U5532 (N_5532,N_1901,N_75);
and U5533 (N_5533,N_232,N_83);
and U5534 (N_5534,N_1062,N_2033);
nor U5535 (N_5535,N_728,N_1121);
nor U5536 (N_5536,N_1539,N_2091);
nand U5537 (N_5537,N_2810,N_328);
nand U5538 (N_5538,N_1114,N_598);
xor U5539 (N_5539,N_1602,N_1572);
or U5540 (N_5540,N_393,N_57);
or U5541 (N_5541,N_2631,N_1548);
or U5542 (N_5542,N_593,N_2970);
or U5543 (N_5543,N_979,N_1424);
or U5544 (N_5544,N_2724,N_2196);
or U5545 (N_5545,N_36,N_1490);
nand U5546 (N_5546,N_2901,N_791);
nor U5547 (N_5547,N_3123,N_1532);
nor U5548 (N_5548,N_1358,N_824);
or U5549 (N_5549,N_780,N_1114);
nor U5550 (N_5550,N_911,N_2633);
nand U5551 (N_5551,N_2864,N_1736);
or U5552 (N_5552,N_2013,N_1620);
and U5553 (N_5553,N_184,N_2328);
or U5554 (N_5554,N_2195,N_614);
nor U5555 (N_5555,N_1920,N_2273);
nand U5556 (N_5556,N_418,N_2655);
nor U5557 (N_5557,N_2149,N_773);
nor U5558 (N_5558,N_794,N_401);
nand U5559 (N_5559,N_140,N_3107);
nor U5560 (N_5560,N_1369,N_1280);
nand U5561 (N_5561,N_2790,N_382);
or U5562 (N_5562,N_629,N_1142);
or U5563 (N_5563,N_1500,N_1776);
xor U5564 (N_5564,N_1064,N_304);
nand U5565 (N_5565,N_554,N_2763);
nand U5566 (N_5566,N_160,N_16);
or U5567 (N_5567,N_27,N_1682);
nand U5568 (N_5568,N_756,N_333);
and U5569 (N_5569,N_2066,N_2030);
and U5570 (N_5570,N_552,N_2893);
and U5571 (N_5571,N_2131,N_1152);
or U5572 (N_5572,N_1390,N_2896);
nor U5573 (N_5573,N_1890,N_3003);
and U5574 (N_5574,N_1044,N_1325);
nor U5575 (N_5575,N_266,N_2254);
nor U5576 (N_5576,N_402,N_496);
nor U5577 (N_5577,N_26,N_1264);
nor U5578 (N_5578,N_728,N_1774);
or U5579 (N_5579,N_1059,N_86);
nand U5580 (N_5580,N_26,N_672);
xnor U5581 (N_5581,N_2253,N_1990);
and U5582 (N_5582,N_1987,N_2565);
nor U5583 (N_5583,N_3085,N_309);
and U5584 (N_5584,N_2938,N_1815);
nand U5585 (N_5585,N_455,N_1059);
or U5586 (N_5586,N_1379,N_863);
and U5587 (N_5587,N_483,N_2271);
nor U5588 (N_5588,N_309,N_363);
nor U5589 (N_5589,N_1871,N_2835);
and U5590 (N_5590,N_2758,N_893);
and U5591 (N_5591,N_1658,N_263);
nand U5592 (N_5592,N_1847,N_1681);
and U5593 (N_5593,N_516,N_2981);
nor U5594 (N_5594,N_2853,N_271);
xnor U5595 (N_5595,N_1332,N_1675);
and U5596 (N_5596,N_1355,N_184);
and U5597 (N_5597,N_1605,N_1337);
nor U5598 (N_5598,N_2196,N_1888);
nand U5599 (N_5599,N_1744,N_1420);
nand U5600 (N_5600,N_1569,N_2246);
nor U5601 (N_5601,N_859,N_3104);
nor U5602 (N_5602,N_770,N_995);
nor U5603 (N_5603,N_161,N_208);
nor U5604 (N_5604,N_2546,N_1847);
nor U5605 (N_5605,N_1396,N_282);
or U5606 (N_5606,N_1604,N_1971);
nand U5607 (N_5607,N_2378,N_2745);
or U5608 (N_5608,N_1746,N_2751);
xnor U5609 (N_5609,N_2952,N_2306);
xor U5610 (N_5610,N_2058,N_1646);
xor U5611 (N_5611,N_2093,N_1632);
xor U5612 (N_5612,N_451,N_1257);
xor U5613 (N_5613,N_1718,N_91);
and U5614 (N_5614,N_1888,N_1204);
or U5615 (N_5615,N_2550,N_1725);
nand U5616 (N_5616,N_2489,N_2069);
xnor U5617 (N_5617,N_1588,N_1708);
nand U5618 (N_5618,N_2290,N_2733);
nor U5619 (N_5619,N_608,N_2532);
nor U5620 (N_5620,N_155,N_2916);
or U5621 (N_5621,N_1716,N_373);
xor U5622 (N_5622,N_1288,N_2644);
nor U5623 (N_5623,N_2208,N_934);
nor U5624 (N_5624,N_2470,N_2905);
or U5625 (N_5625,N_2581,N_1635);
nand U5626 (N_5626,N_1607,N_2614);
and U5627 (N_5627,N_166,N_1794);
xnor U5628 (N_5628,N_853,N_2252);
nand U5629 (N_5629,N_3031,N_121);
nand U5630 (N_5630,N_740,N_124);
nor U5631 (N_5631,N_820,N_868);
nand U5632 (N_5632,N_1756,N_1995);
nand U5633 (N_5633,N_364,N_1790);
xnor U5634 (N_5634,N_161,N_369);
xnor U5635 (N_5635,N_1435,N_1865);
nand U5636 (N_5636,N_1945,N_697);
xnor U5637 (N_5637,N_1028,N_594);
nor U5638 (N_5638,N_3095,N_2822);
or U5639 (N_5639,N_1991,N_2349);
nor U5640 (N_5640,N_2301,N_1452);
or U5641 (N_5641,N_2005,N_2421);
and U5642 (N_5642,N_658,N_2096);
nand U5643 (N_5643,N_1140,N_1653);
nand U5644 (N_5644,N_171,N_2156);
or U5645 (N_5645,N_759,N_1183);
or U5646 (N_5646,N_617,N_1068);
nor U5647 (N_5647,N_2772,N_216);
nor U5648 (N_5648,N_1083,N_491);
nor U5649 (N_5649,N_2107,N_960);
and U5650 (N_5650,N_682,N_2869);
and U5651 (N_5651,N_1053,N_744);
nand U5652 (N_5652,N_1788,N_2067);
and U5653 (N_5653,N_236,N_1141);
nand U5654 (N_5654,N_1667,N_2717);
or U5655 (N_5655,N_4,N_63);
and U5656 (N_5656,N_2251,N_960);
and U5657 (N_5657,N_152,N_162);
and U5658 (N_5658,N_1570,N_1242);
nand U5659 (N_5659,N_847,N_1030);
nor U5660 (N_5660,N_744,N_1160);
nand U5661 (N_5661,N_2481,N_1642);
nor U5662 (N_5662,N_688,N_2991);
nand U5663 (N_5663,N_2023,N_161);
nor U5664 (N_5664,N_3096,N_2173);
nor U5665 (N_5665,N_340,N_1110);
and U5666 (N_5666,N_611,N_1106);
and U5667 (N_5667,N_893,N_2292);
or U5668 (N_5668,N_407,N_2651);
nor U5669 (N_5669,N_712,N_983);
xnor U5670 (N_5670,N_2215,N_2324);
and U5671 (N_5671,N_372,N_706);
and U5672 (N_5672,N_192,N_1790);
nor U5673 (N_5673,N_268,N_1178);
nor U5674 (N_5674,N_466,N_1962);
nor U5675 (N_5675,N_2641,N_1476);
and U5676 (N_5676,N_977,N_1425);
nor U5677 (N_5677,N_2951,N_534);
and U5678 (N_5678,N_1658,N_1078);
and U5679 (N_5679,N_632,N_2342);
nor U5680 (N_5680,N_844,N_1423);
and U5681 (N_5681,N_1603,N_486);
or U5682 (N_5682,N_957,N_3009);
and U5683 (N_5683,N_2371,N_2548);
nor U5684 (N_5684,N_3079,N_2510);
xor U5685 (N_5685,N_2612,N_186);
and U5686 (N_5686,N_2838,N_237);
nor U5687 (N_5687,N_1742,N_2088);
or U5688 (N_5688,N_2178,N_1754);
and U5689 (N_5689,N_524,N_2502);
or U5690 (N_5690,N_2556,N_1128);
or U5691 (N_5691,N_2828,N_309);
xnor U5692 (N_5692,N_1080,N_613);
and U5693 (N_5693,N_2895,N_1097);
or U5694 (N_5694,N_1107,N_586);
and U5695 (N_5695,N_1254,N_2365);
and U5696 (N_5696,N_910,N_648);
nor U5697 (N_5697,N_1656,N_1731);
nand U5698 (N_5698,N_1329,N_2248);
nand U5699 (N_5699,N_1529,N_2065);
or U5700 (N_5700,N_1137,N_2411);
or U5701 (N_5701,N_1462,N_2105);
and U5702 (N_5702,N_1453,N_1209);
or U5703 (N_5703,N_1920,N_435);
nand U5704 (N_5704,N_1853,N_2456);
nand U5705 (N_5705,N_1219,N_1324);
or U5706 (N_5706,N_2357,N_1242);
or U5707 (N_5707,N_911,N_920);
nand U5708 (N_5708,N_2594,N_750);
nor U5709 (N_5709,N_2588,N_241);
and U5710 (N_5710,N_2932,N_1354);
nor U5711 (N_5711,N_1894,N_1694);
and U5712 (N_5712,N_660,N_818);
nand U5713 (N_5713,N_388,N_1690);
or U5714 (N_5714,N_2642,N_112);
nor U5715 (N_5715,N_774,N_762);
nor U5716 (N_5716,N_1587,N_2545);
or U5717 (N_5717,N_860,N_1918);
or U5718 (N_5718,N_575,N_694);
xor U5719 (N_5719,N_2282,N_1627);
and U5720 (N_5720,N_557,N_309);
xnor U5721 (N_5721,N_2947,N_1203);
nor U5722 (N_5722,N_2385,N_2927);
xor U5723 (N_5723,N_2028,N_2885);
and U5724 (N_5724,N_3109,N_1444);
and U5725 (N_5725,N_2316,N_1888);
xor U5726 (N_5726,N_1970,N_1972);
nand U5727 (N_5727,N_2403,N_1047);
nor U5728 (N_5728,N_2394,N_2084);
nor U5729 (N_5729,N_1116,N_2595);
or U5730 (N_5730,N_54,N_1585);
or U5731 (N_5731,N_1393,N_1609);
nor U5732 (N_5732,N_2882,N_2755);
nor U5733 (N_5733,N_2973,N_3006);
nor U5734 (N_5734,N_946,N_72);
xnor U5735 (N_5735,N_546,N_1319);
nand U5736 (N_5736,N_25,N_2795);
and U5737 (N_5737,N_1192,N_298);
xor U5738 (N_5738,N_185,N_2509);
and U5739 (N_5739,N_1105,N_2040);
nor U5740 (N_5740,N_923,N_900);
nand U5741 (N_5741,N_2328,N_113);
nor U5742 (N_5742,N_1533,N_250);
nor U5743 (N_5743,N_1829,N_1988);
or U5744 (N_5744,N_2526,N_1829);
or U5745 (N_5745,N_1549,N_2443);
nand U5746 (N_5746,N_686,N_1918);
and U5747 (N_5747,N_1362,N_1211);
or U5748 (N_5748,N_152,N_282);
and U5749 (N_5749,N_3025,N_467);
nand U5750 (N_5750,N_1972,N_2265);
and U5751 (N_5751,N_2386,N_867);
or U5752 (N_5752,N_208,N_2519);
nand U5753 (N_5753,N_2818,N_2995);
and U5754 (N_5754,N_409,N_1966);
nor U5755 (N_5755,N_1434,N_528);
nor U5756 (N_5756,N_725,N_2693);
nand U5757 (N_5757,N_2193,N_1034);
nand U5758 (N_5758,N_836,N_696);
or U5759 (N_5759,N_518,N_889);
nand U5760 (N_5760,N_941,N_1382);
and U5761 (N_5761,N_316,N_504);
or U5762 (N_5762,N_91,N_1327);
or U5763 (N_5763,N_1651,N_1344);
xnor U5764 (N_5764,N_3104,N_1060);
nand U5765 (N_5765,N_2685,N_352);
or U5766 (N_5766,N_417,N_2481);
xnor U5767 (N_5767,N_1928,N_1680);
nor U5768 (N_5768,N_2778,N_1546);
xnor U5769 (N_5769,N_11,N_2394);
nor U5770 (N_5770,N_1278,N_2407);
and U5771 (N_5771,N_815,N_1739);
nor U5772 (N_5772,N_1945,N_2937);
or U5773 (N_5773,N_393,N_2281);
nand U5774 (N_5774,N_1964,N_1110);
nor U5775 (N_5775,N_2597,N_76);
or U5776 (N_5776,N_2072,N_2964);
nor U5777 (N_5777,N_2568,N_171);
nand U5778 (N_5778,N_1123,N_2185);
nand U5779 (N_5779,N_2090,N_769);
and U5780 (N_5780,N_340,N_1108);
nand U5781 (N_5781,N_1069,N_2128);
or U5782 (N_5782,N_712,N_2889);
or U5783 (N_5783,N_864,N_1091);
nand U5784 (N_5784,N_553,N_2958);
nand U5785 (N_5785,N_368,N_199);
nand U5786 (N_5786,N_2365,N_2679);
or U5787 (N_5787,N_1186,N_1365);
nand U5788 (N_5788,N_2987,N_1276);
or U5789 (N_5789,N_2630,N_1236);
nand U5790 (N_5790,N_1548,N_2625);
and U5791 (N_5791,N_12,N_2080);
nor U5792 (N_5792,N_2022,N_2730);
or U5793 (N_5793,N_2906,N_1137);
nor U5794 (N_5794,N_1960,N_2818);
nand U5795 (N_5795,N_19,N_933);
or U5796 (N_5796,N_2524,N_606);
nand U5797 (N_5797,N_755,N_2802);
nand U5798 (N_5798,N_1716,N_1973);
nor U5799 (N_5799,N_627,N_1648);
nand U5800 (N_5800,N_3013,N_751);
or U5801 (N_5801,N_54,N_945);
or U5802 (N_5802,N_2569,N_2570);
or U5803 (N_5803,N_1263,N_3012);
and U5804 (N_5804,N_2764,N_2874);
xor U5805 (N_5805,N_205,N_447);
nand U5806 (N_5806,N_282,N_1294);
nand U5807 (N_5807,N_1010,N_791);
nand U5808 (N_5808,N_1649,N_2563);
and U5809 (N_5809,N_1919,N_2374);
nor U5810 (N_5810,N_817,N_2107);
and U5811 (N_5811,N_196,N_1977);
nand U5812 (N_5812,N_2703,N_300);
xor U5813 (N_5813,N_1817,N_2599);
or U5814 (N_5814,N_167,N_249);
or U5815 (N_5815,N_1580,N_1544);
and U5816 (N_5816,N_2315,N_3009);
nand U5817 (N_5817,N_3000,N_2633);
or U5818 (N_5818,N_464,N_1993);
and U5819 (N_5819,N_1547,N_407);
or U5820 (N_5820,N_931,N_230);
nand U5821 (N_5821,N_1564,N_3124);
or U5822 (N_5822,N_2300,N_960);
or U5823 (N_5823,N_2983,N_1556);
nand U5824 (N_5824,N_251,N_1292);
or U5825 (N_5825,N_580,N_1229);
and U5826 (N_5826,N_1840,N_1896);
xnor U5827 (N_5827,N_2979,N_984);
or U5828 (N_5828,N_975,N_2766);
or U5829 (N_5829,N_3048,N_973);
nor U5830 (N_5830,N_1267,N_651);
or U5831 (N_5831,N_100,N_663);
and U5832 (N_5832,N_386,N_98);
or U5833 (N_5833,N_703,N_2927);
xnor U5834 (N_5834,N_1908,N_363);
or U5835 (N_5835,N_2123,N_1569);
and U5836 (N_5836,N_320,N_123);
or U5837 (N_5837,N_1282,N_1537);
nand U5838 (N_5838,N_1310,N_383);
and U5839 (N_5839,N_2382,N_2596);
and U5840 (N_5840,N_789,N_2309);
nand U5841 (N_5841,N_1493,N_1291);
or U5842 (N_5842,N_1445,N_671);
or U5843 (N_5843,N_1159,N_2409);
xnor U5844 (N_5844,N_3098,N_632);
nand U5845 (N_5845,N_2887,N_3085);
nor U5846 (N_5846,N_1172,N_72);
and U5847 (N_5847,N_1494,N_1124);
nand U5848 (N_5848,N_1516,N_1275);
and U5849 (N_5849,N_1713,N_2784);
xor U5850 (N_5850,N_2423,N_2355);
and U5851 (N_5851,N_144,N_2587);
or U5852 (N_5852,N_1160,N_1459);
or U5853 (N_5853,N_2686,N_341);
nor U5854 (N_5854,N_1417,N_562);
or U5855 (N_5855,N_1536,N_1637);
nor U5856 (N_5856,N_334,N_686);
nand U5857 (N_5857,N_703,N_2583);
nor U5858 (N_5858,N_1983,N_1997);
or U5859 (N_5859,N_2429,N_1234);
or U5860 (N_5860,N_1737,N_2865);
and U5861 (N_5861,N_132,N_2330);
or U5862 (N_5862,N_497,N_2349);
or U5863 (N_5863,N_530,N_1738);
or U5864 (N_5864,N_1931,N_1963);
and U5865 (N_5865,N_2953,N_1876);
or U5866 (N_5866,N_344,N_698);
or U5867 (N_5867,N_648,N_1391);
or U5868 (N_5868,N_2415,N_1096);
and U5869 (N_5869,N_2511,N_2211);
nor U5870 (N_5870,N_956,N_2673);
and U5871 (N_5871,N_353,N_536);
xnor U5872 (N_5872,N_908,N_110);
nand U5873 (N_5873,N_1215,N_701);
or U5874 (N_5874,N_1270,N_1809);
nand U5875 (N_5875,N_1230,N_2769);
and U5876 (N_5876,N_1177,N_1616);
nor U5877 (N_5877,N_2539,N_976);
nor U5878 (N_5878,N_2954,N_2425);
or U5879 (N_5879,N_990,N_248);
and U5880 (N_5880,N_2055,N_2735);
and U5881 (N_5881,N_2032,N_154);
and U5882 (N_5882,N_2117,N_1218);
and U5883 (N_5883,N_2009,N_2539);
nor U5884 (N_5884,N_1051,N_1914);
xor U5885 (N_5885,N_327,N_1849);
nor U5886 (N_5886,N_1067,N_1340);
nand U5887 (N_5887,N_2380,N_2756);
or U5888 (N_5888,N_300,N_532);
or U5889 (N_5889,N_97,N_2854);
nand U5890 (N_5890,N_835,N_1541);
nor U5891 (N_5891,N_192,N_271);
xnor U5892 (N_5892,N_1066,N_2701);
and U5893 (N_5893,N_438,N_2664);
and U5894 (N_5894,N_1964,N_1813);
nand U5895 (N_5895,N_2617,N_2046);
nand U5896 (N_5896,N_552,N_598);
nor U5897 (N_5897,N_2653,N_2422);
nor U5898 (N_5898,N_2185,N_178);
or U5899 (N_5899,N_685,N_2451);
or U5900 (N_5900,N_2206,N_1204);
xnor U5901 (N_5901,N_791,N_2291);
or U5902 (N_5902,N_2173,N_2761);
or U5903 (N_5903,N_2152,N_2317);
or U5904 (N_5904,N_1554,N_1449);
or U5905 (N_5905,N_2748,N_971);
or U5906 (N_5906,N_2817,N_940);
or U5907 (N_5907,N_2080,N_739);
and U5908 (N_5908,N_939,N_2996);
nand U5909 (N_5909,N_1003,N_990);
nand U5910 (N_5910,N_340,N_1857);
nor U5911 (N_5911,N_2518,N_2492);
nor U5912 (N_5912,N_2460,N_801);
nand U5913 (N_5913,N_1851,N_1842);
and U5914 (N_5914,N_475,N_3011);
or U5915 (N_5915,N_158,N_1650);
nor U5916 (N_5916,N_1179,N_894);
and U5917 (N_5917,N_1490,N_172);
nand U5918 (N_5918,N_2372,N_2259);
or U5919 (N_5919,N_291,N_2375);
or U5920 (N_5920,N_167,N_2913);
nand U5921 (N_5921,N_452,N_900);
nor U5922 (N_5922,N_1514,N_1727);
nand U5923 (N_5923,N_1178,N_1418);
nand U5924 (N_5924,N_1593,N_209);
and U5925 (N_5925,N_462,N_3061);
nand U5926 (N_5926,N_1089,N_1607);
and U5927 (N_5927,N_2379,N_2228);
nand U5928 (N_5928,N_2569,N_2657);
nor U5929 (N_5929,N_555,N_1640);
nand U5930 (N_5930,N_798,N_813);
nand U5931 (N_5931,N_2369,N_3119);
nor U5932 (N_5932,N_2163,N_2283);
nor U5933 (N_5933,N_1451,N_1226);
xor U5934 (N_5934,N_882,N_248);
xnor U5935 (N_5935,N_2860,N_269);
nand U5936 (N_5936,N_3001,N_2168);
xnor U5937 (N_5937,N_2966,N_868);
or U5938 (N_5938,N_1477,N_88);
nor U5939 (N_5939,N_1074,N_2765);
nor U5940 (N_5940,N_1424,N_1982);
or U5941 (N_5941,N_1208,N_155);
nor U5942 (N_5942,N_21,N_2420);
or U5943 (N_5943,N_1372,N_1845);
xor U5944 (N_5944,N_1030,N_2481);
or U5945 (N_5945,N_1126,N_2746);
and U5946 (N_5946,N_2395,N_1016);
nor U5947 (N_5947,N_2014,N_887);
and U5948 (N_5948,N_1199,N_2269);
and U5949 (N_5949,N_2686,N_601);
nor U5950 (N_5950,N_2749,N_1222);
xnor U5951 (N_5951,N_206,N_2057);
or U5952 (N_5952,N_1261,N_2500);
nand U5953 (N_5953,N_320,N_2665);
and U5954 (N_5954,N_1770,N_546);
nand U5955 (N_5955,N_1252,N_2357);
nand U5956 (N_5956,N_2495,N_1014);
or U5957 (N_5957,N_2317,N_824);
or U5958 (N_5958,N_2378,N_1025);
and U5959 (N_5959,N_1019,N_1221);
or U5960 (N_5960,N_1753,N_1577);
nor U5961 (N_5961,N_1891,N_560);
and U5962 (N_5962,N_561,N_2502);
and U5963 (N_5963,N_2012,N_1690);
and U5964 (N_5964,N_2088,N_2717);
nand U5965 (N_5965,N_108,N_1742);
nand U5966 (N_5966,N_2752,N_2746);
or U5967 (N_5967,N_2278,N_1335);
or U5968 (N_5968,N_398,N_2819);
nor U5969 (N_5969,N_2874,N_2046);
and U5970 (N_5970,N_2558,N_2977);
nor U5971 (N_5971,N_496,N_3009);
xnor U5972 (N_5972,N_197,N_1682);
and U5973 (N_5973,N_393,N_2451);
and U5974 (N_5974,N_816,N_46);
nor U5975 (N_5975,N_2015,N_2490);
and U5976 (N_5976,N_1517,N_144);
nand U5977 (N_5977,N_2763,N_1821);
or U5978 (N_5978,N_2304,N_953);
or U5979 (N_5979,N_961,N_153);
nor U5980 (N_5980,N_2339,N_1553);
nand U5981 (N_5981,N_1117,N_1472);
nor U5982 (N_5982,N_656,N_3001);
or U5983 (N_5983,N_376,N_2685);
or U5984 (N_5984,N_984,N_1822);
and U5985 (N_5985,N_3041,N_819);
or U5986 (N_5986,N_1443,N_1655);
or U5987 (N_5987,N_1,N_430);
nand U5988 (N_5988,N_752,N_316);
or U5989 (N_5989,N_2323,N_2394);
nor U5990 (N_5990,N_2275,N_2050);
nand U5991 (N_5991,N_3108,N_2609);
or U5992 (N_5992,N_1498,N_839);
nand U5993 (N_5993,N_2742,N_1483);
and U5994 (N_5994,N_461,N_2697);
nor U5995 (N_5995,N_1933,N_2134);
and U5996 (N_5996,N_574,N_3107);
and U5997 (N_5997,N_2326,N_898);
nand U5998 (N_5998,N_2474,N_1587);
or U5999 (N_5999,N_335,N_2903);
nor U6000 (N_6000,N_2466,N_591);
nor U6001 (N_6001,N_2210,N_2735);
nor U6002 (N_6002,N_2571,N_58);
or U6003 (N_6003,N_2715,N_641);
nor U6004 (N_6004,N_633,N_1214);
nor U6005 (N_6005,N_192,N_1022);
or U6006 (N_6006,N_1118,N_2938);
and U6007 (N_6007,N_1127,N_2971);
and U6008 (N_6008,N_1648,N_173);
or U6009 (N_6009,N_2017,N_1332);
and U6010 (N_6010,N_1935,N_127);
xnor U6011 (N_6011,N_556,N_270);
nand U6012 (N_6012,N_2648,N_2536);
nor U6013 (N_6013,N_923,N_2361);
nand U6014 (N_6014,N_70,N_1880);
or U6015 (N_6015,N_1866,N_2797);
nand U6016 (N_6016,N_545,N_407);
nor U6017 (N_6017,N_1666,N_2940);
nand U6018 (N_6018,N_64,N_65);
or U6019 (N_6019,N_2983,N_2182);
and U6020 (N_6020,N_2335,N_2158);
or U6021 (N_6021,N_1868,N_1417);
nor U6022 (N_6022,N_578,N_1048);
and U6023 (N_6023,N_700,N_2705);
xnor U6024 (N_6024,N_2118,N_2698);
nor U6025 (N_6025,N_2682,N_2179);
nor U6026 (N_6026,N_170,N_1306);
or U6027 (N_6027,N_1707,N_3006);
nand U6028 (N_6028,N_131,N_2800);
xnor U6029 (N_6029,N_1563,N_2331);
nand U6030 (N_6030,N_1156,N_249);
nand U6031 (N_6031,N_2775,N_278);
nor U6032 (N_6032,N_1606,N_3028);
or U6033 (N_6033,N_3004,N_1858);
nor U6034 (N_6034,N_305,N_1658);
or U6035 (N_6035,N_1080,N_936);
or U6036 (N_6036,N_155,N_674);
nor U6037 (N_6037,N_984,N_2295);
or U6038 (N_6038,N_0,N_783);
or U6039 (N_6039,N_910,N_340);
or U6040 (N_6040,N_679,N_1632);
nor U6041 (N_6041,N_1132,N_1286);
nor U6042 (N_6042,N_677,N_297);
nand U6043 (N_6043,N_1814,N_2901);
or U6044 (N_6044,N_1040,N_1036);
xnor U6045 (N_6045,N_804,N_421);
or U6046 (N_6046,N_2858,N_257);
and U6047 (N_6047,N_1564,N_1089);
or U6048 (N_6048,N_450,N_2214);
nor U6049 (N_6049,N_1104,N_982);
nor U6050 (N_6050,N_413,N_2664);
and U6051 (N_6051,N_2085,N_758);
or U6052 (N_6052,N_729,N_3100);
and U6053 (N_6053,N_3036,N_2232);
and U6054 (N_6054,N_2980,N_2935);
nor U6055 (N_6055,N_1244,N_1210);
or U6056 (N_6056,N_872,N_487);
or U6057 (N_6057,N_219,N_1307);
or U6058 (N_6058,N_3064,N_1646);
or U6059 (N_6059,N_106,N_366);
nand U6060 (N_6060,N_1263,N_2643);
or U6061 (N_6061,N_142,N_930);
and U6062 (N_6062,N_1121,N_1150);
nand U6063 (N_6063,N_2095,N_2026);
or U6064 (N_6064,N_597,N_794);
nand U6065 (N_6065,N_2658,N_1069);
xnor U6066 (N_6066,N_2844,N_1531);
or U6067 (N_6067,N_1912,N_1692);
or U6068 (N_6068,N_1723,N_102);
nor U6069 (N_6069,N_340,N_1648);
nor U6070 (N_6070,N_1164,N_1101);
and U6071 (N_6071,N_436,N_918);
or U6072 (N_6072,N_63,N_2916);
nor U6073 (N_6073,N_2112,N_1222);
or U6074 (N_6074,N_1138,N_524);
and U6075 (N_6075,N_586,N_1807);
or U6076 (N_6076,N_1889,N_3100);
nor U6077 (N_6077,N_702,N_1218);
or U6078 (N_6078,N_2103,N_2368);
xnor U6079 (N_6079,N_2642,N_2747);
nand U6080 (N_6080,N_2140,N_2648);
and U6081 (N_6081,N_1,N_1317);
or U6082 (N_6082,N_2092,N_1636);
nor U6083 (N_6083,N_3017,N_546);
and U6084 (N_6084,N_2162,N_1850);
and U6085 (N_6085,N_2633,N_2293);
nand U6086 (N_6086,N_556,N_888);
and U6087 (N_6087,N_1607,N_2239);
or U6088 (N_6088,N_2199,N_1204);
nand U6089 (N_6089,N_775,N_923);
or U6090 (N_6090,N_174,N_1151);
nand U6091 (N_6091,N_612,N_2624);
or U6092 (N_6092,N_1052,N_2482);
or U6093 (N_6093,N_1017,N_1459);
xnor U6094 (N_6094,N_2812,N_1528);
nor U6095 (N_6095,N_1447,N_2919);
xor U6096 (N_6096,N_1294,N_2231);
and U6097 (N_6097,N_1455,N_2175);
nor U6098 (N_6098,N_926,N_2670);
and U6099 (N_6099,N_837,N_1217);
nand U6100 (N_6100,N_20,N_2717);
nor U6101 (N_6101,N_875,N_3122);
nor U6102 (N_6102,N_1000,N_1275);
and U6103 (N_6103,N_1729,N_2906);
or U6104 (N_6104,N_1811,N_1245);
or U6105 (N_6105,N_1008,N_1024);
xnor U6106 (N_6106,N_292,N_602);
nor U6107 (N_6107,N_59,N_2918);
nor U6108 (N_6108,N_854,N_853);
nand U6109 (N_6109,N_132,N_1370);
or U6110 (N_6110,N_2109,N_1361);
nor U6111 (N_6111,N_2727,N_886);
nand U6112 (N_6112,N_2753,N_420);
nor U6113 (N_6113,N_2299,N_1255);
nor U6114 (N_6114,N_40,N_984);
xnor U6115 (N_6115,N_2807,N_3034);
nand U6116 (N_6116,N_3056,N_628);
or U6117 (N_6117,N_282,N_1387);
nor U6118 (N_6118,N_2719,N_2733);
nand U6119 (N_6119,N_1313,N_492);
nand U6120 (N_6120,N_1127,N_1146);
xnor U6121 (N_6121,N_2517,N_591);
or U6122 (N_6122,N_2289,N_338);
nor U6123 (N_6123,N_2801,N_1399);
nor U6124 (N_6124,N_2029,N_1089);
or U6125 (N_6125,N_1630,N_2037);
and U6126 (N_6126,N_483,N_841);
nand U6127 (N_6127,N_2025,N_1079);
and U6128 (N_6128,N_1278,N_1954);
or U6129 (N_6129,N_1876,N_627);
nor U6130 (N_6130,N_9,N_2215);
xnor U6131 (N_6131,N_136,N_1396);
and U6132 (N_6132,N_2793,N_1625);
nor U6133 (N_6133,N_1244,N_559);
or U6134 (N_6134,N_1935,N_3056);
or U6135 (N_6135,N_1830,N_2538);
nor U6136 (N_6136,N_2265,N_441);
or U6137 (N_6137,N_2481,N_258);
nor U6138 (N_6138,N_1323,N_2357);
and U6139 (N_6139,N_3013,N_1367);
nand U6140 (N_6140,N_1827,N_1275);
and U6141 (N_6141,N_347,N_2915);
nor U6142 (N_6142,N_1809,N_2422);
and U6143 (N_6143,N_3032,N_1801);
nand U6144 (N_6144,N_1496,N_719);
or U6145 (N_6145,N_458,N_2714);
nand U6146 (N_6146,N_1508,N_1095);
nor U6147 (N_6147,N_416,N_2279);
nand U6148 (N_6148,N_617,N_1747);
and U6149 (N_6149,N_1963,N_2307);
and U6150 (N_6150,N_398,N_1744);
nand U6151 (N_6151,N_251,N_1316);
nand U6152 (N_6152,N_2363,N_1940);
nand U6153 (N_6153,N_1775,N_2251);
and U6154 (N_6154,N_1923,N_470);
or U6155 (N_6155,N_340,N_2661);
or U6156 (N_6156,N_22,N_591);
nand U6157 (N_6157,N_745,N_116);
and U6158 (N_6158,N_2986,N_1703);
nand U6159 (N_6159,N_575,N_2004);
or U6160 (N_6160,N_830,N_393);
nand U6161 (N_6161,N_1310,N_2188);
and U6162 (N_6162,N_275,N_1234);
and U6163 (N_6163,N_824,N_1585);
and U6164 (N_6164,N_2257,N_619);
nand U6165 (N_6165,N_3047,N_2832);
xor U6166 (N_6166,N_211,N_1554);
and U6167 (N_6167,N_1570,N_1916);
nand U6168 (N_6168,N_1608,N_2629);
and U6169 (N_6169,N_1408,N_1313);
xor U6170 (N_6170,N_2735,N_391);
or U6171 (N_6171,N_2688,N_1913);
nor U6172 (N_6172,N_139,N_501);
nor U6173 (N_6173,N_292,N_2750);
or U6174 (N_6174,N_1130,N_309);
xor U6175 (N_6175,N_1718,N_1964);
nor U6176 (N_6176,N_1865,N_506);
nand U6177 (N_6177,N_2290,N_2408);
nand U6178 (N_6178,N_512,N_1747);
nand U6179 (N_6179,N_1749,N_1288);
nor U6180 (N_6180,N_2702,N_2687);
or U6181 (N_6181,N_1351,N_3021);
and U6182 (N_6182,N_2502,N_2280);
and U6183 (N_6183,N_226,N_804);
or U6184 (N_6184,N_2603,N_2863);
and U6185 (N_6185,N_1325,N_1384);
or U6186 (N_6186,N_967,N_2565);
xnor U6187 (N_6187,N_2496,N_2835);
nor U6188 (N_6188,N_223,N_1989);
and U6189 (N_6189,N_1686,N_86);
nor U6190 (N_6190,N_1330,N_2073);
nand U6191 (N_6191,N_2280,N_404);
xor U6192 (N_6192,N_713,N_1714);
and U6193 (N_6193,N_964,N_2959);
xnor U6194 (N_6194,N_701,N_1515);
nor U6195 (N_6195,N_2404,N_1618);
xor U6196 (N_6196,N_1319,N_364);
and U6197 (N_6197,N_1370,N_722);
xor U6198 (N_6198,N_1228,N_600);
nand U6199 (N_6199,N_271,N_767);
nand U6200 (N_6200,N_1183,N_459);
nor U6201 (N_6201,N_240,N_1249);
nand U6202 (N_6202,N_0,N_1341);
or U6203 (N_6203,N_1825,N_2107);
nor U6204 (N_6204,N_1887,N_1792);
and U6205 (N_6205,N_37,N_2789);
or U6206 (N_6206,N_2478,N_84);
nand U6207 (N_6207,N_874,N_2868);
nand U6208 (N_6208,N_2403,N_587);
nor U6209 (N_6209,N_3034,N_945);
xor U6210 (N_6210,N_395,N_1218);
nor U6211 (N_6211,N_379,N_558);
and U6212 (N_6212,N_1078,N_1236);
and U6213 (N_6213,N_2192,N_1984);
and U6214 (N_6214,N_1196,N_2279);
or U6215 (N_6215,N_2061,N_65);
nand U6216 (N_6216,N_2159,N_145);
nor U6217 (N_6217,N_1663,N_2152);
nor U6218 (N_6218,N_2734,N_740);
nand U6219 (N_6219,N_2210,N_1184);
nor U6220 (N_6220,N_2662,N_385);
or U6221 (N_6221,N_228,N_1152);
nand U6222 (N_6222,N_785,N_1016);
and U6223 (N_6223,N_1242,N_2469);
and U6224 (N_6224,N_108,N_2773);
xor U6225 (N_6225,N_2919,N_2077);
or U6226 (N_6226,N_908,N_3118);
nand U6227 (N_6227,N_599,N_781);
nor U6228 (N_6228,N_883,N_2235);
nor U6229 (N_6229,N_539,N_940);
and U6230 (N_6230,N_2339,N_2570);
nor U6231 (N_6231,N_981,N_2328);
xor U6232 (N_6232,N_531,N_1982);
and U6233 (N_6233,N_61,N_1185);
nand U6234 (N_6234,N_2183,N_1080);
nand U6235 (N_6235,N_3097,N_1947);
and U6236 (N_6236,N_1362,N_2498);
and U6237 (N_6237,N_2746,N_1633);
xnor U6238 (N_6238,N_2231,N_2274);
nor U6239 (N_6239,N_891,N_660);
nand U6240 (N_6240,N_1998,N_1287);
and U6241 (N_6241,N_1543,N_1519);
and U6242 (N_6242,N_2700,N_1874);
or U6243 (N_6243,N_1394,N_2293);
and U6244 (N_6244,N_1506,N_442);
xor U6245 (N_6245,N_788,N_557);
nor U6246 (N_6246,N_2434,N_1693);
nor U6247 (N_6247,N_549,N_2326);
nand U6248 (N_6248,N_1302,N_660);
nor U6249 (N_6249,N_582,N_1748);
nor U6250 (N_6250,N_4121,N_4505);
nand U6251 (N_6251,N_4177,N_5374);
or U6252 (N_6252,N_3208,N_3670);
nor U6253 (N_6253,N_4440,N_3937);
nor U6254 (N_6254,N_3494,N_4904);
or U6255 (N_6255,N_3555,N_5398);
and U6256 (N_6256,N_4903,N_6013);
nor U6257 (N_6257,N_4523,N_3802);
nor U6258 (N_6258,N_5224,N_4267);
nand U6259 (N_6259,N_6134,N_4047);
nor U6260 (N_6260,N_6052,N_5114);
or U6261 (N_6261,N_4392,N_6037);
and U6262 (N_6262,N_5811,N_5622);
nand U6263 (N_6263,N_5864,N_3828);
nand U6264 (N_6264,N_4421,N_4941);
nor U6265 (N_6265,N_3462,N_3948);
nor U6266 (N_6266,N_5530,N_3360);
nand U6267 (N_6267,N_4023,N_5677);
or U6268 (N_6268,N_5316,N_4947);
or U6269 (N_6269,N_5230,N_4720);
nor U6270 (N_6270,N_4160,N_3709);
or U6271 (N_6271,N_3553,N_3356);
nor U6272 (N_6272,N_5023,N_3759);
nor U6273 (N_6273,N_3599,N_3924);
xnor U6274 (N_6274,N_4622,N_3724);
and U6275 (N_6275,N_5275,N_5024);
and U6276 (N_6276,N_6071,N_3886);
and U6277 (N_6277,N_4724,N_4530);
or U6278 (N_6278,N_3812,N_5472);
and U6279 (N_6279,N_3605,N_5640);
and U6280 (N_6280,N_5556,N_5404);
and U6281 (N_6281,N_5710,N_5691);
and U6282 (N_6282,N_6166,N_4165);
nand U6283 (N_6283,N_3327,N_5800);
and U6284 (N_6284,N_4119,N_3297);
or U6285 (N_6285,N_4925,N_4367);
or U6286 (N_6286,N_5718,N_5132);
nand U6287 (N_6287,N_5507,N_5003);
xor U6288 (N_6288,N_3939,N_5694);
xor U6289 (N_6289,N_5151,N_4113);
or U6290 (N_6290,N_5304,N_4384);
or U6291 (N_6291,N_3324,N_4747);
nor U6292 (N_6292,N_3193,N_4923);
and U6293 (N_6293,N_4460,N_5381);
and U6294 (N_6294,N_5774,N_4285);
and U6295 (N_6295,N_5908,N_3721);
nand U6296 (N_6296,N_3662,N_4757);
xor U6297 (N_6297,N_5070,N_4551);
nor U6298 (N_6298,N_4883,N_5687);
or U6299 (N_6299,N_5169,N_3281);
or U6300 (N_6300,N_6109,N_5413);
nor U6301 (N_6301,N_5784,N_3813);
or U6302 (N_6302,N_3716,N_3596);
or U6303 (N_6303,N_5568,N_3621);
nor U6304 (N_6304,N_4279,N_3769);
nor U6305 (N_6305,N_4965,N_5515);
nand U6306 (N_6306,N_5342,N_4576);
nor U6307 (N_6307,N_3756,N_5550);
and U6308 (N_6308,N_3291,N_6048);
xnor U6309 (N_6309,N_5088,N_3307);
nor U6310 (N_6310,N_3166,N_3567);
or U6311 (N_6311,N_5836,N_3400);
nand U6312 (N_6312,N_5803,N_4933);
or U6313 (N_6313,N_4985,N_3664);
xor U6314 (N_6314,N_4344,N_5223);
and U6315 (N_6315,N_6099,N_4178);
nor U6316 (N_6316,N_4703,N_5337);
nor U6317 (N_6317,N_5134,N_5427);
nand U6318 (N_6318,N_3995,N_4887);
or U6319 (N_6319,N_5684,N_3699);
nor U6320 (N_6320,N_4281,N_3614);
nand U6321 (N_6321,N_6075,N_3339);
xor U6322 (N_6322,N_3783,N_5778);
and U6323 (N_6323,N_3870,N_3689);
and U6324 (N_6324,N_5650,N_3710);
and U6325 (N_6325,N_6015,N_4426);
nor U6326 (N_6326,N_4345,N_5872);
and U6327 (N_6327,N_3698,N_4553);
nor U6328 (N_6328,N_3365,N_4256);
nand U6329 (N_6329,N_6120,N_5212);
xnor U6330 (N_6330,N_4782,N_4522);
nor U6331 (N_6331,N_4362,N_6116);
and U6332 (N_6332,N_5179,N_4766);
or U6333 (N_6333,N_3965,N_5729);
xnor U6334 (N_6334,N_3545,N_3781);
nor U6335 (N_6335,N_5032,N_4577);
xor U6336 (N_6336,N_6202,N_4041);
nand U6337 (N_6337,N_4272,N_5081);
nor U6338 (N_6338,N_3369,N_4462);
or U6339 (N_6339,N_5076,N_6069);
or U6340 (N_6340,N_3142,N_5971);
nor U6341 (N_6341,N_3498,N_5228);
nand U6342 (N_6342,N_3550,N_6242);
or U6343 (N_6343,N_5518,N_5166);
or U6344 (N_6344,N_5731,N_3469);
xor U6345 (N_6345,N_4400,N_4060);
xnor U6346 (N_6346,N_4005,N_3129);
nor U6347 (N_6347,N_5601,N_3925);
or U6348 (N_6348,N_3933,N_3635);
and U6349 (N_6349,N_3987,N_4250);
or U6350 (N_6350,N_5757,N_4994);
nor U6351 (N_6351,N_6246,N_3714);
nor U6352 (N_6352,N_5943,N_3482);
nor U6353 (N_6353,N_4222,N_3554);
or U6354 (N_6354,N_5322,N_5524);
nor U6355 (N_6355,N_3632,N_4917);
xnor U6356 (N_6356,N_4278,N_5865);
nand U6357 (N_6357,N_4702,N_3520);
or U6358 (N_6358,N_3736,N_5012);
and U6359 (N_6359,N_3475,N_5192);
and U6360 (N_6360,N_5537,N_4475);
and U6361 (N_6361,N_6045,N_5558);
xnor U6362 (N_6362,N_5257,N_4737);
nor U6363 (N_6363,N_4940,N_5593);
nand U6364 (N_6364,N_3273,N_3201);
and U6365 (N_6365,N_3474,N_3859);
nor U6366 (N_6366,N_6035,N_5418);
and U6367 (N_6367,N_4111,N_4274);
nand U6368 (N_6368,N_5309,N_3223);
or U6369 (N_6369,N_4218,N_5915);
and U6370 (N_6370,N_5749,N_4856);
nand U6371 (N_6371,N_4340,N_4488);
or U6372 (N_6372,N_4775,N_6153);
and U6373 (N_6373,N_3808,N_3486);
nor U6374 (N_6374,N_3209,N_5875);
nor U6375 (N_6375,N_3126,N_5352);
xor U6376 (N_6376,N_4434,N_5891);
nor U6377 (N_6377,N_4152,N_5609);
nor U6378 (N_6378,N_3231,N_6235);
or U6379 (N_6379,N_5119,N_3835);
and U6380 (N_6380,N_5849,N_5141);
nor U6381 (N_6381,N_5520,N_4351);
or U6382 (N_6382,N_4070,N_4337);
nand U6383 (N_6383,N_4103,N_3165);
and U6384 (N_6384,N_5676,N_3881);
nand U6385 (N_6385,N_3815,N_4497);
or U6386 (N_6386,N_5722,N_3125);
nand U6387 (N_6387,N_3315,N_5137);
xor U6388 (N_6388,N_4495,N_5978);
and U6389 (N_6389,N_3237,N_6210);
nand U6390 (N_6390,N_3861,N_5871);
nand U6391 (N_6391,N_5690,N_5017);
xor U6392 (N_6392,N_4466,N_5576);
nand U6393 (N_6393,N_4543,N_4777);
nand U6394 (N_6394,N_6151,N_6174);
nor U6395 (N_6395,N_3233,N_3323);
nor U6396 (N_6396,N_3580,N_6133);
nor U6397 (N_6397,N_4311,N_3500);
or U6398 (N_6398,N_4208,N_4455);
nand U6399 (N_6399,N_4671,N_4874);
or U6400 (N_6400,N_3650,N_5913);
and U6401 (N_6401,N_4824,N_5582);
and U6402 (N_6402,N_5540,N_5987);
and U6403 (N_6403,N_3252,N_5801);
and U6404 (N_6404,N_4322,N_4306);
or U6405 (N_6405,N_3241,N_5636);
and U6406 (N_6406,N_4637,N_6214);
and U6407 (N_6407,N_4118,N_3383);
and U6408 (N_6408,N_3417,N_5363);
nand U6409 (N_6409,N_4851,N_5868);
xnor U6410 (N_6410,N_4352,N_6064);
xnor U6411 (N_6411,N_4538,N_6240);
nor U6412 (N_6412,N_5847,N_4498);
nand U6413 (N_6413,N_4486,N_5464);
and U6414 (N_6414,N_3525,N_3404);
and U6415 (N_6415,N_5428,N_5581);
nand U6416 (N_6416,N_4013,N_3405);
xor U6417 (N_6417,N_3953,N_5016);
nand U6418 (N_6418,N_5643,N_3268);
nor U6419 (N_6419,N_4286,N_4648);
or U6420 (N_6420,N_3975,N_4197);
nor U6421 (N_6421,N_5945,N_4396);
nor U6422 (N_6422,N_5154,N_4859);
and U6423 (N_6423,N_4050,N_3860);
nor U6424 (N_6424,N_6205,N_5782);
and U6425 (N_6425,N_6150,N_5058);
nor U6426 (N_6426,N_3236,N_5999);
or U6427 (N_6427,N_3683,N_3210);
or U6428 (N_6428,N_4857,N_6155);
and U6429 (N_6429,N_5035,N_5354);
xnor U6430 (N_6430,N_5532,N_6018);
and U6431 (N_6431,N_5209,N_5890);
nor U6432 (N_6432,N_5810,N_4220);
nor U6433 (N_6433,N_5693,N_4886);
nand U6434 (N_6434,N_3577,N_4492);
nand U6435 (N_6435,N_4644,N_5683);
nand U6436 (N_6436,N_5312,N_4612);
nor U6437 (N_6437,N_3612,N_5853);
or U6438 (N_6438,N_5099,N_6025);
nor U6439 (N_6439,N_5013,N_3354);
nand U6440 (N_6440,N_6243,N_5689);
and U6441 (N_6441,N_4879,N_3695);
nand U6442 (N_6442,N_5742,N_3973);
and U6443 (N_6443,N_5008,N_3674);
nand U6444 (N_6444,N_3408,N_4592);
and U6445 (N_6445,N_5766,N_4201);
nand U6446 (N_6446,N_4019,N_5130);
xor U6447 (N_6447,N_4558,N_3432);
nor U6448 (N_6448,N_4547,N_4975);
and U6449 (N_6449,N_4324,N_4271);
or U6450 (N_6450,N_4048,N_4591);
and U6451 (N_6451,N_6124,N_4246);
or U6452 (N_6452,N_4786,N_4020);
xor U6453 (N_6453,N_6041,N_4989);
nor U6454 (N_6454,N_5619,N_5727);
or U6455 (N_6455,N_5029,N_6237);
nor U6456 (N_6456,N_5655,N_3258);
nand U6457 (N_6457,N_3930,N_5806);
xnor U6458 (N_6458,N_5171,N_5599);
nand U6459 (N_6459,N_3822,N_3591);
or U6460 (N_6460,N_5646,N_3493);
xnor U6461 (N_6461,N_4571,N_5318);
or U6462 (N_6462,N_4825,N_4138);
nor U6463 (N_6463,N_5059,N_5375);
nor U6464 (N_6464,N_5829,N_3232);
or U6465 (N_6465,N_3495,N_4009);
and U6466 (N_6466,N_4051,N_4139);
xnor U6467 (N_6467,N_5483,N_5435);
or U6468 (N_6468,N_3561,N_4316);
or U6469 (N_6469,N_6196,N_4793);
and U6470 (N_6470,N_4785,N_4598);
nand U6471 (N_6471,N_4045,N_5184);
and U6472 (N_6472,N_3378,N_4948);
and U6473 (N_6473,N_5506,N_3566);
and U6474 (N_6474,N_5571,N_3915);
or U6475 (N_6475,N_5461,N_3626);
or U6476 (N_6476,N_4258,N_4546);
xor U6477 (N_6477,N_6054,N_5086);
and U6478 (N_6478,N_4716,N_5298);
and U6479 (N_6479,N_5063,N_3363);
and U6480 (N_6480,N_4844,N_4100);
nand U6481 (N_6481,N_5542,N_5271);
or U6482 (N_6482,N_4875,N_4718);
nand U6483 (N_6483,N_4705,N_4759);
xor U6484 (N_6484,N_3445,N_6047);
and U6485 (N_6485,N_6191,N_4841);
nor U6486 (N_6486,N_5952,N_4094);
xnor U6487 (N_6487,N_4327,N_3506);
and U6488 (N_6488,N_4878,N_3798);
nor U6489 (N_6489,N_5843,N_5826);
and U6490 (N_6490,N_5794,N_3682);
and U6491 (N_6491,N_3658,N_4908);
or U6492 (N_6492,N_3950,N_5832);
nor U6493 (N_6493,N_5388,N_4383);
or U6494 (N_6494,N_5528,N_5178);
and U6495 (N_6495,N_3468,N_4457);
and U6496 (N_6496,N_3430,N_4707);
nor U6497 (N_6497,N_5028,N_4907);
nand U6498 (N_6498,N_3247,N_6028);
and U6499 (N_6499,N_4536,N_5068);
nand U6500 (N_6500,N_3429,N_4231);
nand U6501 (N_6501,N_4378,N_4052);
nand U6502 (N_6502,N_3681,N_4022);
nand U6503 (N_6503,N_4938,N_4951);
or U6504 (N_6504,N_4656,N_5923);
nand U6505 (N_6505,N_5155,N_4853);
or U6506 (N_6506,N_4305,N_5197);
nand U6507 (N_6507,N_4524,N_4000);
nor U6508 (N_6508,N_5295,N_3868);
and U6509 (N_6509,N_3829,N_6198);
xnor U6510 (N_6510,N_6031,N_4884);
nor U6511 (N_6511,N_5454,N_6088);
nand U6512 (N_6512,N_5373,N_3441);
nand U6513 (N_6513,N_5451,N_4706);
nand U6514 (N_6514,N_4910,N_5419);
xor U6515 (N_6515,N_4942,N_3180);
or U6516 (N_6516,N_5252,N_3839);
or U6517 (N_6517,N_3697,N_4451);
nand U6518 (N_6518,N_4583,N_5495);
nor U6519 (N_6519,N_3585,N_5698);
or U6520 (N_6520,N_5681,N_5336);
and U6521 (N_6521,N_3280,N_5122);
nand U6522 (N_6522,N_4922,N_5860);
nor U6523 (N_6523,N_4804,N_5262);
nor U6524 (N_6524,N_3801,N_3913);
and U6525 (N_6525,N_3818,N_4595);
nor U6526 (N_6526,N_3856,N_6003);
nor U6527 (N_6527,N_5019,N_5045);
nor U6528 (N_6528,N_3294,N_3963);
and U6529 (N_6529,N_4200,N_4784);
nand U6530 (N_6530,N_5344,N_5211);
and U6531 (N_6531,N_5979,N_5588);
and U6532 (N_6532,N_3132,N_5232);
nand U6533 (N_6533,N_6046,N_3148);
nand U6534 (N_6534,N_3789,N_5052);
or U6535 (N_6535,N_5862,N_4335);
or U6536 (N_6536,N_5938,N_3277);
xnor U6537 (N_6537,N_5445,N_3825);
or U6538 (N_6538,N_5394,N_5265);
and U6539 (N_6539,N_5198,N_4573);
xor U6540 (N_6540,N_3836,N_5205);
nor U6541 (N_6541,N_4395,N_3684);
nor U6542 (N_6542,N_3336,N_5709);
nand U6543 (N_6543,N_3712,N_3945);
nand U6544 (N_6544,N_5513,N_4668);
or U6545 (N_6545,N_4389,N_4869);
nand U6546 (N_6546,N_5760,N_4276);
or U6547 (N_6547,N_5544,N_3216);
nor U6548 (N_6548,N_5338,N_3667);
nor U6549 (N_6549,N_4817,N_3473);
nand U6550 (N_6550,N_3185,N_3738);
nand U6551 (N_6551,N_5508,N_4638);
and U6552 (N_6552,N_4461,N_4628);
and U6553 (N_6553,N_3496,N_4653);
xor U6554 (N_6554,N_4004,N_5201);
and U6555 (N_6555,N_4982,N_4413);
and U6556 (N_6556,N_3941,N_3136);
and U6557 (N_6557,N_6199,N_4128);
and U6558 (N_6558,N_5680,N_5820);
or U6559 (N_6559,N_4137,N_5380);
and U6560 (N_6560,N_4544,N_4846);
nor U6561 (N_6561,N_4713,N_5592);
nand U6562 (N_6562,N_5635,N_3528);
nor U6563 (N_6563,N_5768,N_3666);
nand U6564 (N_6564,N_3979,N_5595);
or U6565 (N_6565,N_3641,N_4959);
nor U6566 (N_6566,N_5561,N_6200);
and U6567 (N_6567,N_6234,N_3958);
or U6568 (N_6568,N_5196,N_5095);
nor U6569 (N_6569,N_5956,N_4868);
nand U6570 (N_6570,N_4528,N_5022);
nand U6571 (N_6571,N_3625,N_3332);
or U6572 (N_6572,N_4710,N_5522);
nor U6573 (N_6573,N_6084,N_4015);
and U6574 (N_6574,N_4277,N_6011);
and U6575 (N_6575,N_4570,N_3164);
or U6576 (N_6576,N_6177,N_3174);
nor U6577 (N_6577,N_6192,N_4297);
or U6578 (N_6578,N_5191,N_4292);
xnor U6579 (N_6579,N_5988,N_5856);
and U6580 (N_6580,N_3578,N_5447);
nand U6581 (N_6581,N_5071,N_5092);
nor U6582 (N_6582,N_5414,N_4319);
nand U6583 (N_6583,N_5219,N_4323);
nand U6584 (N_6584,N_5431,N_4752);
xor U6585 (N_6585,N_5401,N_4655);
nor U6586 (N_6586,N_5170,N_5400);
nor U6587 (N_6587,N_5926,N_4732);
nor U6588 (N_6588,N_3313,N_5093);
nor U6589 (N_6589,N_3864,N_3501);
nor U6590 (N_6590,N_3821,N_4545);
nand U6591 (N_6591,N_3899,N_4079);
and U6592 (N_6592,N_4650,N_5409);
nand U6593 (N_6593,N_6140,N_5442);
nand U6594 (N_6594,N_4066,N_6143);
nand U6595 (N_6595,N_5053,N_3371);
or U6596 (N_6596,N_5216,N_6212);
or U6597 (N_6597,N_3325,N_3978);
nor U6598 (N_6598,N_5966,N_4755);
nand U6599 (N_6599,N_5725,N_5563);
nor U6600 (N_6600,N_4363,N_5724);
nor U6601 (N_6601,N_3316,N_5207);
nand U6602 (N_6602,N_4725,N_4860);
nor U6603 (N_6603,N_4454,N_3838);
and U6604 (N_6604,N_6135,N_5111);
nand U6605 (N_6605,N_3853,N_4863);
and U6606 (N_6606,N_4957,N_6089);
nor U6607 (N_6607,N_4935,N_4429);
nor U6608 (N_6608,N_4789,N_4763);
nand U6609 (N_6609,N_5867,N_6201);
xor U6610 (N_6610,N_4465,N_3396);
and U6611 (N_6611,N_5402,N_4039);
nor U6612 (N_6612,N_3618,N_3147);
and U6613 (N_6613,N_5152,N_4411);
or U6614 (N_6614,N_4155,N_4534);
nor U6615 (N_6615,N_3673,N_3192);
or U6616 (N_6616,N_4792,N_4767);
or U6617 (N_6617,N_4620,N_5448);
nand U6618 (N_6618,N_4476,N_6105);
and U6619 (N_6619,N_3139,N_5270);
or U6620 (N_6620,N_3706,N_6204);
or U6621 (N_6621,N_4254,N_5456);
and U6622 (N_6622,N_5714,N_5160);
xor U6623 (N_6623,N_5751,N_5930);
and U6624 (N_6624,N_4296,N_3725);
and U6625 (N_6625,N_5285,N_5175);
or U6626 (N_6626,N_6208,N_4114);
nor U6627 (N_6627,N_4597,N_6217);
nand U6628 (N_6628,N_3568,N_5737);
nand U6629 (N_6629,N_4123,N_3734);
nand U6630 (N_6630,N_5379,N_5505);
nor U6631 (N_6631,N_6231,N_5747);
nor U6632 (N_6632,N_6171,N_4587);
nor U6633 (N_6633,N_5772,N_6023);
nand U6634 (N_6634,N_4689,N_3352);
nor U6635 (N_6635,N_3645,N_5096);
and U6636 (N_6636,N_3348,N_3345);
or U6637 (N_6637,N_5236,N_4679);
or U6638 (N_6638,N_4663,N_3576);
and U6639 (N_6639,N_6049,N_3535);
or U6640 (N_6640,N_3351,N_5533);
and U6641 (N_6641,N_4428,N_6189);
nand U6642 (N_6642,N_4293,N_4144);
nor U6643 (N_6643,N_4420,N_3203);
or U6644 (N_6644,N_4235,N_3878);
nor U6645 (N_6645,N_3522,N_6014);
and U6646 (N_6646,N_5586,N_4988);
xor U6647 (N_6647,N_6167,N_3942);
xor U6648 (N_6648,N_5632,N_4607);
or U6649 (N_6649,N_5072,N_4388);
and U6650 (N_6650,N_5857,N_4783);
nand U6651 (N_6651,N_3521,N_4130);
nor U6652 (N_6652,N_4112,N_5376);
nand U6653 (N_6653,N_3589,N_3135);
nor U6654 (N_6654,N_4207,N_3637);
nand U6655 (N_6655,N_5254,N_3154);
nor U6656 (N_6656,N_5904,N_3259);
xor U6657 (N_6657,N_4820,N_4405);
nand U6658 (N_6658,N_6193,N_3540);
nor U6659 (N_6659,N_4012,N_3765);
and U6660 (N_6660,N_5341,N_5667);
nor U6661 (N_6661,N_5873,N_5281);
nor U6662 (N_6662,N_5535,N_3448);
nor U6663 (N_6663,N_4209,N_5504);
and U6664 (N_6664,N_4680,N_4801);
and U6665 (N_6665,N_4176,N_5311);
or U6666 (N_6666,N_5629,N_4055);
nor U6667 (N_6667,N_4240,N_3957);
or U6668 (N_6668,N_3776,N_5185);
nand U6669 (N_6669,N_3288,N_3145);
and U6670 (N_6670,N_5009,N_4414);
or U6671 (N_6671,N_6233,N_4581);
nor U6672 (N_6672,N_5734,N_5605);
nor U6673 (N_6673,N_3377,N_3692);
nand U6674 (N_6674,N_5974,N_6081);
xor U6675 (N_6675,N_4683,N_5077);
nand U6676 (N_6676,N_5434,N_5036);
nand U6677 (N_6677,N_4794,N_3791);
nor U6678 (N_6678,N_5534,N_6239);
nand U6679 (N_6679,N_3687,N_4101);
nand U6680 (N_6680,N_4195,N_4192);
and U6681 (N_6681,N_5415,N_4699);
or U6682 (N_6682,N_5962,N_3179);
nor U6683 (N_6683,N_5131,N_4781);
nor U6684 (N_6684,N_4893,N_4236);
xor U6685 (N_6685,N_3832,N_3982);
or U6686 (N_6686,N_5031,N_6245);
and U6687 (N_6687,N_4661,N_4387);
or U6688 (N_6688,N_5443,N_3533);
and U6689 (N_6689,N_3908,N_4269);
nand U6690 (N_6690,N_3537,N_3927);
nand U6691 (N_6691,N_5750,N_5079);
nor U6692 (N_6692,N_4473,N_5280);
or U6693 (N_6693,N_5673,N_3954);
nand U6694 (N_6694,N_3219,N_6063);
and U6695 (N_6695,N_6077,N_3235);
xor U6696 (N_6696,N_3701,N_3349);
nand U6697 (N_6697,N_3249,N_3993);
or U6698 (N_6698,N_4175,N_3873);
or U6699 (N_6699,N_3848,N_5288);
and U6700 (N_6700,N_3660,N_4247);
and U6701 (N_6701,N_3949,N_3367);
nor U6702 (N_6702,N_4828,N_3470);
nand U6703 (N_6703,N_3169,N_3205);
nand U6704 (N_6704,N_4603,N_5195);
nor U6705 (N_6705,N_3436,N_5991);
and U6706 (N_6706,N_4651,N_4253);
or U6707 (N_6707,N_3196,N_4564);
nand U6708 (N_6708,N_3994,N_3851);
nand U6709 (N_6709,N_4483,N_5366);
and U6710 (N_6710,N_5549,N_5320);
nor U6711 (N_6711,N_5973,N_3321);
nor U6712 (N_6712,N_3159,N_4448);
or U6713 (N_6713,N_5929,N_6129);
nand U6714 (N_6714,N_5602,N_3601);
or U6715 (N_6715,N_4168,N_4987);
nand U6716 (N_6716,N_5324,N_4918);
xnor U6717 (N_6717,N_3977,N_3184);
and U6718 (N_6718,N_5514,N_5253);
nand U6719 (N_6719,N_4030,N_5963);
nor U6720 (N_6720,N_5142,N_5692);
nor U6721 (N_6721,N_6148,N_5446);
and U6722 (N_6722,N_4614,N_6033);
and U6723 (N_6723,N_3879,N_4998);
nor U6724 (N_6724,N_5422,N_4810);
nor U6725 (N_6725,N_3523,N_3382);
and U6726 (N_6726,N_4517,N_5881);
nand U6727 (N_6727,N_5112,N_3976);
and U6728 (N_6728,N_4764,N_5243);
and U6729 (N_6729,N_5007,N_3140);
or U6730 (N_6730,N_3199,N_6137);
and U6731 (N_6731,N_5116,N_3240);
nand U6732 (N_6732,N_6184,N_5613);
or U6733 (N_6733,N_6158,N_4185);
nor U6734 (N_6734,N_4173,N_5361);
nor U6735 (N_6735,N_3338,N_3855);
and U6736 (N_6736,N_5510,N_5181);
or U6737 (N_6737,N_4212,N_5215);
nor U6738 (N_6738,N_6224,N_4031);
or U6739 (N_6739,N_6165,N_5327);
nand U6740 (N_6740,N_5701,N_4179);
or U6741 (N_6741,N_3213,N_4894);
and U6742 (N_6742,N_5299,N_5905);
nor U6743 (N_6743,N_3328,N_5752);
nor U6744 (N_6744,N_4096,N_3391);
and U6745 (N_6745,N_4295,N_5630);
nor U6746 (N_6746,N_4646,N_3425);
nor U6747 (N_6747,N_4374,N_4234);
and U6748 (N_6748,N_4575,N_6249);
and U6749 (N_6749,N_3892,N_4649);
or U6750 (N_6750,N_6006,N_4471);
and U6751 (N_6751,N_4809,N_5033);
and U6752 (N_6752,N_4180,N_4954);
xnor U6753 (N_6753,N_3127,N_4080);
xnor U6754 (N_6754,N_5664,N_4289);
xor U6755 (N_6755,N_4880,N_5957);
nand U6756 (N_6756,N_6119,N_5168);
xnor U6757 (N_6757,N_3492,N_3156);
nor U6758 (N_6758,N_5302,N_3865);
nand U6759 (N_6759,N_3342,N_5239);
xor U6760 (N_6760,N_3676,N_4540);
or U6761 (N_6761,N_4916,N_4895);
or U6762 (N_6762,N_3546,N_4756);
nor U6763 (N_6763,N_5828,N_4010);
or U6764 (N_6764,N_3901,N_3916);
and U6765 (N_6765,N_3974,N_5049);
and U6766 (N_6766,N_5060,N_4730);
nor U6767 (N_6767,N_3551,N_5863);
nand U6768 (N_6768,N_5392,N_4437);
or U6769 (N_6769,N_4660,N_5964);
nor U6770 (N_6770,N_5432,N_5656);
nor U6771 (N_6771,N_5649,N_3722);
or U6772 (N_6772,N_4059,N_3481);
nand U6773 (N_6773,N_6176,N_5329);
or U6774 (N_6774,N_5055,N_4812);
nor U6775 (N_6775,N_4842,N_4610);
nand U6776 (N_6776,N_3592,N_5246);
and U6777 (N_6777,N_5659,N_5719);
nand U6778 (N_6778,N_3446,N_5740);
and U6779 (N_6779,N_4127,N_3413);
or U6780 (N_6780,N_3452,N_5560);
or U6781 (N_6781,N_5162,N_6042);
and U6782 (N_6782,N_5547,N_4394);
nand U6783 (N_6783,N_5995,N_3301);
and U6784 (N_6784,N_5064,N_5965);
nor U6785 (N_6785,N_6228,N_4866);
and U6786 (N_6786,N_4091,N_3906);
or U6787 (N_6787,N_5950,N_4688);
nor U6788 (N_6788,N_5165,N_6220);
xnor U6789 (N_6789,N_3264,N_4214);
nand U6790 (N_6790,N_5705,N_3903);
nor U6791 (N_6791,N_5140,N_5367);
nor U6792 (N_6792,N_3743,N_5347);
and U6793 (N_6793,N_4830,N_6229);
nand U6794 (N_6794,N_5308,N_5256);
nor U6795 (N_6795,N_4334,N_5303);
nor U6796 (N_6796,N_5654,N_4381);
and U6797 (N_6797,N_4206,N_4708);
nor U6798 (N_6798,N_4172,N_5796);
and U6799 (N_6799,N_6218,N_4417);
xor U6800 (N_6800,N_5517,N_5416);
nor U6801 (N_6801,N_4480,N_3372);
or U6802 (N_6802,N_3295,N_5578);
xnor U6803 (N_6803,N_5226,N_4596);
nand U6804 (N_6804,N_3557,N_5437);
and U6805 (N_6805,N_3990,N_4599);
nand U6806 (N_6806,N_3266,N_5770);
nand U6807 (N_6807,N_4141,N_4858);
and U6808 (N_6808,N_4108,N_4574);
nand U6809 (N_6809,N_4924,N_5405);
nor U6810 (N_6810,N_5272,N_4382);
nand U6811 (N_6811,N_6096,N_4372);
xor U6812 (N_6812,N_3395,N_3777);
nand U6813 (N_6813,N_5488,N_4242);
or U6814 (N_6814,N_4117,N_5889);
nor U6815 (N_6815,N_4881,N_5369);
and U6816 (N_6816,N_5946,N_5384);
nand U6817 (N_6817,N_5206,N_3727);
nand U6818 (N_6818,N_4565,N_4548);
nand U6819 (N_6819,N_4419,N_4474);
nor U6820 (N_6820,N_5066,N_4736);
nor U6821 (N_6821,N_3679,N_5903);
or U6822 (N_6822,N_4937,N_3705);
and U6823 (N_6823,N_6238,N_3439);
nand U6824 (N_6824,N_3239,N_5700);
and U6825 (N_6825,N_4479,N_4072);
or U6826 (N_6826,N_4229,N_5675);
and U6827 (N_6827,N_3587,N_3702);
nand U6828 (N_6828,N_3940,N_5633);
nand U6829 (N_6829,N_4341,N_5982);
or U6830 (N_6830,N_3790,N_4645);
and U6831 (N_6831,N_3284,N_4704);
and U6832 (N_6832,N_3733,N_5217);
nand U6833 (N_6833,N_4182,N_6072);
nor U6834 (N_6834,N_5877,N_3428);
nand U6835 (N_6835,N_5792,N_3753);
nand U6836 (N_6836,N_5237,N_3575);
nand U6837 (N_6837,N_3293,N_5555);
nor U6838 (N_6838,N_4537,N_5221);
or U6839 (N_6839,N_5614,N_3289);
nand U6840 (N_6840,N_4726,N_5610);
nor U6841 (N_6841,N_3877,N_5678);
nor U6842 (N_6842,N_3898,N_3245);
and U6843 (N_6843,N_3897,N_3794);
and U6844 (N_6844,N_3314,N_5529);
and U6845 (N_6845,N_4349,N_4053);
and U6846 (N_6846,N_5525,N_5580);
nand U6847 (N_6847,N_4379,N_4862);
or U6848 (N_6848,N_6130,N_4751);
or U6849 (N_6849,N_3911,N_4762);
and U6850 (N_6850,N_6186,N_3850);
and U6851 (N_6851,N_3444,N_6114);
nor U6852 (N_6852,N_3584,N_5240);
and U6853 (N_6853,N_4035,N_4626);
or U6854 (N_6854,N_4997,N_6187);
or U6855 (N_6855,N_4990,N_3893);
or U6856 (N_6856,N_5470,N_5020);
or U6857 (N_6857,N_5389,N_6020);
and U6858 (N_6858,N_3206,N_5921);
nand U6859 (N_6859,N_5378,N_5048);
or U6860 (N_6860,N_3385,N_3541);
and U6861 (N_6861,N_5969,N_3171);
xnor U6862 (N_6862,N_3785,N_4882);
nor U6863 (N_6863,N_3558,N_5440);
nor U6864 (N_6864,N_4829,N_5735);
nor U6865 (N_6865,N_3426,N_5866);
nand U6866 (N_6866,N_4818,N_3221);
or U6867 (N_6867,N_3891,N_5744);
and U6868 (N_6868,N_5476,N_5666);
xnor U6869 (N_6869,N_6179,N_3552);
or U6870 (N_6870,N_3871,N_3677);
or U6871 (N_6871,N_4971,N_4129);
nor U6872 (N_6872,N_4686,N_5481);
nor U6873 (N_6873,N_5972,N_4131);
or U6874 (N_6874,N_5027,N_3390);
nor U6875 (N_6875,N_3876,N_6211);
or U6876 (N_6876,N_5557,N_5951);
nand U6877 (N_6877,N_4520,N_5305);
or U6878 (N_6878,N_3675,N_5047);
and U6879 (N_6879,N_3661,N_6182);
xnor U6880 (N_6880,N_4360,N_4719);
nand U6881 (N_6881,N_5455,N_5598);
nor U6882 (N_6882,N_4738,N_3594);
or U6883 (N_6883,N_5541,N_6163);
nand U6884 (N_6884,N_5519,N_3852);
nand U6885 (N_6885,N_5014,N_3654);
nand U6886 (N_6886,N_3526,N_3731);
nor U6887 (N_6887,N_5838,N_3715);
or U6888 (N_6888,N_3431,N_4016);
nor U6889 (N_6889,N_3513,N_5286);
and U6890 (N_6890,N_5706,N_4188);
nor U6891 (N_6891,N_4037,N_4855);
and U6892 (N_6892,N_5642,N_3779);
nand U6893 (N_6893,N_5566,N_5350);
and U6894 (N_6894,N_6087,N_5644);
nand U6895 (N_6895,N_4946,N_5377);
nand U6896 (N_6896,N_3613,N_3157);
or U6897 (N_6897,N_5235,N_3630);
nor U6898 (N_6898,N_5842,N_4518);
nand U6899 (N_6899,N_3988,N_5977);
or U6900 (N_6900,N_5682,N_3303);
nand U6901 (N_6901,N_4819,N_4761);
nor U6902 (N_6902,N_3814,N_6085);
nor U6903 (N_6903,N_3549,N_3772);
nor U6904 (N_6904,N_6108,N_5314);
and U6905 (N_6905,N_4594,N_5761);
nand U6906 (N_6906,N_3420,N_3711);
and U6907 (N_6907,N_3388,N_5387);
or U6908 (N_6908,N_5583,N_5471);
xnor U6909 (N_6909,N_5564,N_4265);
xor U6910 (N_6910,N_5763,N_6181);
and U6911 (N_6911,N_5948,N_5040);
nor U6912 (N_6912,N_5886,N_4554);
and U6913 (N_6913,N_4913,N_4338);
nand U6914 (N_6914,N_3780,N_4038);
xnor U6915 (N_6915,N_5485,N_3636);
xor U6916 (N_6916,N_3971,N_5699);
and U6917 (N_6917,N_6083,N_4056);
and U6918 (N_6918,N_5370,N_3629);
xnor U6919 (N_6919,N_3357,N_6195);
nor U6920 (N_6920,N_5840,N_5998);
or U6921 (N_6921,N_4664,N_5831);
xor U6922 (N_6922,N_5815,N_5231);
and U6923 (N_6923,N_6078,N_6131);
nand U6924 (N_6924,N_4058,N_6127);
nand U6925 (N_6925,N_5715,N_5939);
and U6926 (N_6926,N_4044,N_5624);
nand U6927 (N_6927,N_5527,N_4731);
or U6928 (N_6928,N_3263,N_6111);
nor U6929 (N_6929,N_6159,N_3620);
and U6930 (N_6930,N_3846,N_5559);
nor U6931 (N_6931,N_4864,N_5545);
nor U6932 (N_6932,N_5509,N_4418);
xnor U6933 (N_6933,N_3745,N_5425);
nand U6934 (N_6934,N_5397,N_3224);
xnor U6935 (N_6935,N_3161,N_3748);
nand U6936 (N_6936,N_4635,N_3341);
and U6937 (N_6937,N_4616,N_4104);
nand U6938 (N_6938,N_4996,N_5148);
xnor U6939 (N_6939,N_5855,N_5453);
or U6940 (N_6940,N_4399,N_4203);
or U6941 (N_6941,N_4758,N_4945);
or U6942 (N_6942,N_4225,N_5885);
nand U6943 (N_6943,N_5386,N_3544);
nor U6944 (N_6944,N_5739,N_4776);
and U6945 (N_6945,N_4215,N_4239);
or U6946 (N_6946,N_5138,N_5604);
or U6947 (N_6947,N_3218,N_6222);
xnor U6948 (N_6948,N_4559,N_4024);
xnor U6949 (N_6949,N_3732,N_5596);
nor U6950 (N_6950,N_5671,N_3296);
and U6951 (N_6951,N_4712,N_3646);
or U6952 (N_6952,N_4521,N_4373);
and U6953 (N_6953,N_3969,N_5468);
nand U6954 (N_6954,N_4733,N_3796);
nand U6955 (N_6955,N_4248,N_5620);
or U6956 (N_6956,N_4143,N_6065);
or U6957 (N_6957,N_4541,N_3168);
nor U6958 (N_6958,N_5565,N_3735);
nand U6959 (N_6959,N_3176,N_3703);
and U6960 (N_6960,N_4124,N_6038);
xor U6961 (N_6961,N_4157,N_5021);
nand U6962 (N_6962,N_3844,N_3872);
nor U6963 (N_6963,N_5827,N_6190);
or U6964 (N_6964,N_5406,N_3479);
nand U6965 (N_6965,N_4282,N_4561);
and U6966 (N_6966,N_5242,N_6112);
nand U6967 (N_6967,N_5748,N_6227);
nand U6968 (N_6968,N_3686,N_4532);
nor U6969 (N_6969,N_3421,N_6097);
nand U6970 (N_6970,N_6132,N_6101);
nand U6971 (N_6971,N_5776,N_4202);
and U6972 (N_6972,N_4769,N_3680);
xnor U6973 (N_6973,N_4826,N_4299);
and U6974 (N_6974,N_3920,N_5685);
nand U6975 (N_6975,N_5762,N_5393);
or U6976 (N_6976,N_3787,N_5487);
and U6977 (N_6977,N_4146,N_4519);
nand U6978 (N_6978,N_4533,N_3274);
nand U6979 (N_6979,N_3305,N_5164);
or U6980 (N_6980,N_5084,N_3884);
and U6981 (N_6981,N_5627,N_4727);
xor U6982 (N_6982,N_6247,N_5621);
or U6983 (N_6983,N_5004,N_6009);
xnor U6984 (N_6984,N_5944,N_4555);
or U6985 (N_6985,N_5186,N_5467);
xor U6986 (N_6986,N_3992,N_5358);
nor U6987 (N_6987,N_4386,N_3397);
nand U6988 (N_6988,N_6056,N_6043);
nor U6989 (N_6989,N_4151,N_4357);
or U6990 (N_6990,N_6244,N_6216);
nand U6991 (N_6991,N_5225,N_4566);
xnor U6992 (N_6992,N_5273,N_3138);
or U6993 (N_6993,N_4968,N_3996);
and U6994 (N_6994,N_4264,N_3505);
and U6995 (N_6995,N_5107,N_5833);
nor U6996 (N_6996,N_5247,N_3964);
nor U6997 (N_6997,N_6080,N_4071);
and U6998 (N_6998,N_3931,N_6029);
nand U6999 (N_6999,N_5591,N_4443);
nand U7000 (N_7000,N_5125,N_3519);
nor U7001 (N_7001,N_5543,N_5218);
nor U7002 (N_7002,N_6030,N_4260);
nand U7003 (N_7003,N_5928,N_5512);
nor U7004 (N_7004,N_5641,N_6067);
and U7005 (N_7005,N_4284,N_4364);
or U7006 (N_7006,N_5315,N_5825);
nand U7007 (N_7007,N_4032,N_3833);
xor U7008 (N_7008,N_5996,N_5105);
and U7009 (N_7009,N_5420,N_4190);
and U7010 (N_7010,N_4962,N_3195);
xor U7011 (N_7011,N_4452,N_5078);
or U7012 (N_7012,N_6053,N_5769);
and U7013 (N_7013,N_3644,N_3804);
nor U7014 (N_7014,N_5970,N_3602);
xnor U7015 (N_7015,N_4890,N_5249);
nor U7016 (N_7016,N_4963,N_5038);
xor U7017 (N_7017,N_5932,N_4743);
xnor U7018 (N_7018,N_6197,N_4148);
nand U7019 (N_7019,N_4950,N_4618);
nor U7020 (N_7020,N_3634,N_5672);
nor U7021 (N_7021,N_5301,N_5947);
xor U7022 (N_7022,N_5670,N_4613);
and U7023 (N_7023,N_5579,N_6138);
nand U7024 (N_7024,N_4216,N_5124);
xor U7025 (N_7025,N_5333,N_5918);
or U7026 (N_7026,N_3403,N_4799);
nor U7027 (N_7027,N_4011,N_3150);
nand U7028 (N_7028,N_3243,N_5469);
or U7029 (N_7029,N_3137,N_6062);
nand U7030 (N_7030,N_5764,N_4061);
nand U7031 (N_7031,N_5010,N_3361);
xor U7032 (N_7032,N_3271,N_4442);
nor U7033 (N_7033,N_5845,N_4835);
or U7034 (N_7034,N_5292,N_4978);
or U7035 (N_7035,N_4427,N_5989);
and U7036 (N_7036,N_5458,N_3693);
xnor U7037 (N_7037,N_3633,N_5959);
xor U7038 (N_7038,N_3512,N_3300);
or U7039 (N_7039,N_4026,N_6113);
nand U7040 (N_7040,N_5346,N_4659);
nand U7041 (N_7041,N_3869,N_4721);
and U7042 (N_7042,N_6126,N_5661);
nor U7043 (N_7043,N_3610,N_4074);
nand U7044 (N_7044,N_6050,N_5188);
or U7045 (N_7045,N_5738,N_5500);
nor U7046 (N_7046,N_5051,N_5878);
and U7047 (N_7047,N_4008,N_3883);
nand U7048 (N_7048,N_3770,N_3217);
and U7049 (N_7049,N_6160,N_4078);
nand U7050 (N_7050,N_4255,N_5882);
and U7051 (N_7051,N_4606,N_5390);
nand U7052 (N_7052,N_5323,N_4463);
or U7053 (N_7053,N_5901,N_5713);
nand U7054 (N_7054,N_5896,N_5234);
xnor U7055 (N_7055,N_5733,N_4243);
nor U7056 (N_7056,N_4976,N_4780);
nor U7057 (N_7057,N_3509,N_4149);
nor U7058 (N_7058,N_3374,N_5259);
nor U7059 (N_7059,N_4934,N_6156);
and U7060 (N_7060,N_4876,N_3380);
xnor U7061 (N_7061,N_3623,N_5859);
and U7062 (N_7062,N_3582,N_4087);
nand U7063 (N_7063,N_3816,N_4459);
xnor U7064 (N_7064,N_4109,N_5612);
nor U7065 (N_7065,N_4515,N_4525);
and U7066 (N_7066,N_4385,N_5173);
nor U7067 (N_7067,N_3728,N_5823);
or U7068 (N_7068,N_4837,N_5611);
and U7069 (N_7069,N_3767,N_5474);
and U7070 (N_7070,N_5482,N_3197);
nand U7071 (N_7071,N_4692,N_6004);
nor U7072 (N_7072,N_3466,N_3989);
or U7073 (N_7073,N_3754,N_6141);
xor U7074 (N_7074,N_5497,N_6117);
nor U7075 (N_7075,N_6142,N_3364);
nor U7076 (N_7076,N_5712,N_4979);
and U7077 (N_7077,N_3595,N_5902);
nand U7078 (N_7078,N_4915,N_3857);
or U7079 (N_7079,N_4539,N_6145);
nor U7080 (N_7080,N_3398,N_6209);
and U7081 (N_7081,N_4036,N_3488);
and U7082 (N_7082,N_4623,N_3647);
nand U7083 (N_7083,N_6215,N_5005);
or U7084 (N_7084,N_5608,N_5584);
xnor U7085 (N_7085,N_3152,N_5802);
nor U7086 (N_7086,N_3607,N_5372);
and U7087 (N_7087,N_3980,N_5108);
nand U7088 (N_7088,N_5102,N_5880);
nor U7089 (N_7089,N_3387,N_5716);
nor U7090 (N_7090,N_4169,N_3283);
nand U7091 (N_7091,N_3968,N_5741);
nor U7092 (N_7092,N_4723,N_5658);
or U7093 (N_7093,N_4346,N_3478);
nor U7094 (N_7094,N_4393,N_4888);
and U7095 (N_7095,N_3570,N_6005);
nand U7096 (N_7096,N_5711,N_3991);
nor U7097 (N_7097,N_5787,N_3786);
and U7098 (N_7098,N_3460,N_3921);
nand U7099 (N_7099,N_3455,N_3986);
and U7100 (N_7100,N_5082,N_6144);
nor U7101 (N_7101,N_4156,N_4167);
and U7102 (N_7102,N_3511,N_4550);
or U7103 (N_7103,N_3847,N_3830);
nor U7104 (N_7104,N_5294,N_4244);
nor U7105 (N_7105,N_5001,N_5348);
and U7106 (N_7106,N_3807,N_6060);
and U7107 (N_7107,N_3178,N_4313);
or U7108 (N_7108,N_4321,N_5203);
and U7109 (N_7109,N_3485,N_3163);
nor U7110 (N_7110,N_3502,N_3803);
and U7111 (N_7111,N_6070,N_4115);
and U7112 (N_7112,N_4634,N_5278);
nand U7113 (N_7113,N_5858,N_6173);
or U7114 (N_7114,N_5167,N_5618);
nor U7115 (N_7115,N_4069,N_3225);
nand U7116 (N_7116,N_3598,N_3747);
and U7117 (N_7117,N_4062,N_3359);
or U7118 (N_7118,N_3464,N_5771);
and U7119 (N_7119,N_6032,N_5911);
nor U7120 (N_7120,N_4135,N_5567);
xor U7121 (N_7121,N_5793,N_5494);
and U7122 (N_7122,N_4586,N_5704);
or U7123 (N_7123,N_5399,N_4064);
nor U7124 (N_7124,N_4832,N_3534);
nand U7125 (N_7125,N_5985,N_3318);
xnor U7126 (N_7126,N_6236,N_4252);
nand U7127 (N_7127,N_3929,N_4552);
xor U7128 (N_7128,N_4939,N_4081);
and U7129 (N_7129,N_4605,N_5933);
and U7130 (N_7130,N_4579,N_4972);
and U7131 (N_7131,N_3966,N_5465);
nor U7132 (N_7132,N_4506,N_4375);
xor U7133 (N_7133,N_5492,N_4986);
nand U7134 (N_7134,N_5289,N_6154);
or U7135 (N_7135,N_5351,N_4183);
nor U7136 (N_7136,N_4477,N_3447);
nor U7137 (N_7137,N_3628,N_3758);
and U7138 (N_7138,N_4779,N_5332);
or U7139 (N_7139,N_3424,N_5268);
nand U7140 (N_7140,N_3543,N_4270);
nand U7141 (N_7141,N_3574,N_6123);
xnor U7142 (N_7142,N_5695,N_3984);
nor U7143 (N_7143,N_5914,N_5163);
and U7144 (N_7144,N_4693,N_4370);
nand U7145 (N_7145,N_5954,N_4082);
nand U7146 (N_7146,N_4162,N_5157);
and U7147 (N_7147,N_4800,N_5238);
nand U7148 (N_7148,N_4873,N_3375);
nor U7149 (N_7149,N_5789,N_4729);
or U7150 (N_7150,N_4681,N_4585);
or U7151 (N_7151,N_5147,N_5953);
nand U7152 (N_7152,N_5331,N_5149);
nand U7153 (N_7153,N_3355,N_4956);
nor U7154 (N_7154,N_5073,N_3409);
and U7155 (N_7155,N_4654,N_4676);
nor U7156 (N_7156,N_5779,N_5753);
and U7157 (N_7157,N_6207,N_5981);
or U7158 (N_7158,N_4912,N_4193);
nor U7159 (N_7159,N_3972,N_4308);
xor U7160 (N_7160,N_3917,N_5128);
and U7161 (N_7161,N_4865,N_3659);
nor U7162 (N_7162,N_4872,N_5745);
or U7163 (N_7163,N_4099,N_4136);
nor U7164 (N_7164,N_4850,N_3890);
and U7165 (N_7165,N_5213,N_5851);
or U7166 (N_7166,N_3649,N_3465);
nor U7167 (N_7167,N_4808,N_4631);
or U7168 (N_7168,N_4791,N_4088);
or U7169 (N_7169,N_6008,N_5382);
nand U7170 (N_7170,N_4991,N_3256);
xor U7171 (N_7171,N_4194,N_4740);
and U7172 (N_7172,N_4073,N_5362);
or U7173 (N_7173,N_4134,N_4969);
nand U7174 (N_7174,N_5025,N_6094);
or U7175 (N_7175,N_6068,N_3141);
nand U7176 (N_7176,N_5936,N_4930);
nor U7177 (N_7177,N_3442,N_4224);
nand U7178 (N_7178,N_5174,N_3343);
xor U7179 (N_7179,N_3854,N_6175);
xor U7180 (N_7180,N_6136,N_5730);
or U7181 (N_7181,N_3617,N_5244);
and U7182 (N_7182,N_5615,N_4238);
or U7183 (N_7183,N_5097,N_3932);
and U7184 (N_7184,N_5531,N_4140);
nand U7185 (N_7185,N_3368,N_5080);
nand U7186 (N_7186,N_4588,N_4981);
xor U7187 (N_7187,N_5874,N_5967);
and U7188 (N_7188,N_3952,N_3308);
or U7189 (N_7189,N_3153,N_3183);
nand U7190 (N_7190,N_3329,N_3202);
and U7191 (N_7191,N_3773,N_4952);
or U7192 (N_7192,N_5403,N_4633);
nor U7193 (N_7193,N_5879,N_4456);
nor U7194 (N_7194,N_4665,N_5156);
and U7195 (N_7195,N_3961,N_5199);
nand U7196 (N_7196,N_5821,N_3741);
and U7197 (N_7197,N_5797,N_5245);
or U7198 (N_7198,N_4690,N_4353);
nand U7199 (N_7199,N_4931,N_3718);
or U7200 (N_7200,N_5044,N_4677);
nor U7201 (N_7201,N_4132,N_4490);
and U7202 (N_7202,N_6147,N_3704);
and U7203 (N_7203,N_5260,N_5837);
nand U7204 (N_7204,N_4018,N_4701);
xnor U7205 (N_7205,N_4350,N_3862);
or U7206 (N_7206,N_4511,N_3443);
nor U7207 (N_7207,N_4516,N_3333);
nor U7208 (N_7208,N_3642,N_4641);
and U7209 (N_7209,N_4439,N_4687);
nor U7210 (N_7210,N_3322,N_5018);
xor U7211 (N_7211,N_5410,N_5279);
and U7212 (N_7212,N_5407,N_6092);
and U7213 (N_7213,N_5631,N_3820);
nor U7214 (N_7214,N_5136,N_4926);
nand U7215 (N_7215,N_5208,N_4892);
or U7216 (N_7216,N_4120,N_5912);
and U7217 (N_7217,N_3516,N_5848);
and U7218 (N_7218,N_4805,N_5736);
or U7219 (N_7219,N_4086,N_3453);
or U7220 (N_7220,N_5888,N_4847);
xnor U7221 (N_7221,N_4943,N_3726);
or U7222 (N_7222,N_3782,N_5412);
or U7223 (N_7223,N_5204,N_5927);
or U7224 (N_7224,N_5002,N_6230);
nor U7225 (N_7225,N_5310,N_4715);
or U7226 (N_7226,N_4126,N_5117);
or U7227 (N_7227,N_6241,N_6206);
nor U7228 (N_7228,N_3867,N_5942);
xnor U7229 (N_7229,N_5083,N_5085);
nor U7230 (N_7230,N_4891,N_4845);
nand U7231 (N_7231,N_5809,N_5227);
nand U7232 (N_7232,N_5562,N_4189);
nor U7233 (N_7233,N_5150,N_5220);
or U7234 (N_7234,N_4076,N_5269);
nand U7235 (N_7235,N_4315,N_3334);
or U7236 (N_7236,N_3542,N_3177);
and U7237 (N_7237,N_4150,N_5651);
and U7238 (N_7238,N_5523,N_3414);
or U7239 (N_7239,N_3837,N_5463);
and U7240 (N_7240,N_3746,N_5728);
or U7241 (N_7241,N_3547,N_5293);
nor U7242 (N_7242,N_6178,N_4770);
nand U7243 (N_7243,N_5708,N_4110);
nor U7244 (N_7244,N_3563,N_5439);
nor U7245 (N_7245,N_3507,N_3651);
nor U7246 (N_7246,N_6012,N_5807);
xnor U7247 (N_7247,N_3616,N_3774);
nor U7248 (N_7248,N_5460,N_5365);
nand U7249 (N_7249,N_5328,N_5577);
xnor U7250 (N_7250,N_4611,N_4839);
nand U7251 (N_7251,N_4911,N_5480);
nand U7252 (N_7252,N_4241,N_3730);
or U7253 (N_7253,N_5898,N_5839);
nor U7254 (N_7254,N_4992,N_3556);
nor U7255 (N_7255,N_5484,N_4803);
and U7256 (N_7256,N_4049,N_3737);
or U7257 (N_7257,N_4105,N_3751);
nor U7258 (N_7258,N_6002,N_5805);
nor U7259 (N_7259,N_4542,N_4266);
or U7260 (N_7260,N_4491,N_3309);
or U7261 (N_7261,N_5300,N_4054);
and U7262 (N_7262,N_4033,N_6074);
nand U7263 (N_7263,N_5732,N_4569);
xor U7264 (N_7264,N_5039,N_4582);
xnor U7265 (N_7265,N_4093,N_4042);
or U7266 (N_7266,N_3131,N_4469);
and U7267 (N_7267,N_4339,N_4410);
or U7268 (N_7268,N_5087,N_3189);
nand U7269 (N_7269,N_5127,N_5276);
nor U7270 (N_7270,N_4259,N_5767);
nor U7271 (N_7271,N_5429,N_4478);
or U7272 (N_7272,N_5267,N_4694);
or U7273 (N_7273,N_3713,N_5703);
or U7274 (N_7274,N_3394,N_5997);
nor U7275 (N_7275,N_6055,N_5287);
nor U7276 (N_7276,N_5261,N_3222);
and U7277 (N_7277,N_4181,N_5819);
nor U7278 (N_7278,N_6168,N_5104);
nand U7279 (N_7279,N_3440,N_5349);
and U7280 (N_7280,N_5490,N_5993);
nor U7281 (N_7281,N_3571,N_5841);
or U7282 (N_7282,N_6232,N_4262);
and U7283 (N_7283,N_5343,N_3228);
or U7284 (N_7284,N_3508,N_3160);
nor U7285 (N_7285,N_4927,N_4489);
or U7286 (N_7286,N_3874,N_3970);
nor U7287 (N_7287,N_4807,N_6086);
or U7288 (N_7288,N_4102,N_5118);
or U7289 (N_7289,N_3946,N_3834);
nor U7290 (N_7290,N_4640,N_5958);
and U7291 (N_7291,N_3656,N_5574);
or U7292 (N_7292,N_3624,N_5552);
nand U7293 (N_7293,N_4453,N_3450);
nand U7294 (N_7294,N_5723,N_4040);
and U7295 (N_7295,N_3840,N_5830);
and U7296 (N_7296,N_4288,N_4802);
nor U7297 (N_7297,N_3744,N_3842);
nor U7298 (N_7298,N_3476,N_5854);
xor U7299 (N_7299,N_5835,N_6213);
and U7300 (N_7300,N_5790,N_5870);
xor U7301 (N_7301,N_6115,N_5074);
or U7302 (N_7302,N_4902,N_5626);
nand U7303 (N_7303,N_5919,N_4980);
nor U7304 (N_7304,N_4174,N_4083);
nor U7305 (N_7305,N_5182,N_4161);
and U7306 (N_7306,N_5153,N_4508);
and U7307 (N_7307,N_4291,N_4312);
and U7308 (N_7308,N_4095,N_5501);
nand U7309 (N_7309,N_3902,N_5250);
nor U7310 (N_7310,N_4424,N_3909);
nand U7311 (N_7311,N_5098,N_6226);
nor U7312 (N_7312,N_5940,N_4342);
or U7313 (N_7313,N_6021,N_4298);
nand U7314 (N_7314,N_4014,N_5551);
nand U7315 (N_7315,N_5450,N_5371);
and U7316 (N_7316,N_5101,N_3604);
and U7317 (N_7317,N_5120,N_3900);
nor U7318 (N_7318,N_5696,N_4261);
nor U7319 (N_7319,N_4330,N_4233);
and U7320 (N_7320,N_3234,N_3652);
or U7321 (N_7321,N_5473,N_5834);
or U7322 (N_7322,N_4447,N_5662);
nor U7323 (N_7323,N_3226,N_3319);
nor U7324 (N_7324,N_3480,N_3826);
nor U7325 (N_7325,N_3379,N_3463);
xnor U7326 (N_7326,N_6090,N_4709);
nand U7327 (N_7327,N_5255,N_4746);
nand U7328 (N_7328,N_3299,N_4920);
or U7329 (N_7329,N_6061,N_6221);
and U7330 (N_7330,N_5941,N_5546);
or U7331 (N_7331,N_3895,N_6162);
or U7332 (N_7332,N_5746,N_5773);
and U7333 (N_7333,N_4896,N_5030);
nor U7334 (N_7334,N_3928,N_4697);
and U7335 (N_7335,N_5975,N_5980);
nand U7336 (N_7336,N_5385,N_4090);
or U7337 (N_7337,N_3270,N_4993);
and U7338 (N_7338,N_6194,N_3914);
nand U7339 (N_7339,N_4748,N_5786);
and U7340 (N_7340,N_4325,N_6103);
nand U7341 (N_7341,N_4223,N_4584);
nor U7342 (N_7342,N_5360,N_3962);
nor U7343 (N_7343,N_5475,N_5106);
or U7344 (N_7344,N_5491,N_5493);
nand U7345 (N_7345,N_3560,N_4287);
and U7346 (N_7346,N_4929,N_5335);
nor U7347 (N_7347,N_5754,N_5931);
or U7348 (N_7348,N_5983,N_4133);
nand U7349 (N_7349,N_3215,N_5949);
and U7350 (N_7350,N_4556,N_5266);
nor U7351 (N_7351,N_5822,N_3491);
nand U7352 (N_7352,N_5968,N_3700);
nand U7353 (N_7353,N_3810,N_5417);
nand U7354 (N_7354,N_6040,N_5193);
and U7355 (N_7355,N_5326,N_3619);
nor U7356 (N_7356,N_3331,N_3172);
or U7357 (N_7357,N_4371,N_5717);
nand U7358 (N_7358,N_4682,N_3707);
xnor U7359 (N_7359,N_3882,N_3538);
xor U7360 (N_7360,N_3490,N_4512);
or U7361 (N_7361,N_3627,N_5411);
and U7362 (N_7362,N_3362,N_5143);
or U7363 (N_7363,N_4021,N_3723);
nor U7364 (N_7364,N_3524,N_6036);
xnor U7365 (N_7365,N_3517,N_3194);
or U7366 (N_7366,N_4122,N_3212);
and U7367 (N_7367,N_6118,N_5496);
xor U7368 (N_7368,N_5818,N_3317);
nor U7369 (N_7369,N_5992,N_4691);
nand U7370 (N_7370,N_3399,N_5884);
nand U7371 (N_7371,N_3761,N_5258);
nor U7372 (N_7372,N_3435,N_5594);
or U7373 (N_7373,N_4734,N_5121);
nand U7374 (N_7374,N_3366,N_3880);
nand U7375 (N_7375,N_5426,N_5189);
or U7376 (N_7376,N_4487,N_4380);
nor U7377 (N_7377,N_3944,N_4795);
or U7378 (N_7378,N_6149,N_3151);
nor U7379 (N_7379,N_3951,N_4158);
nor U7380 (N_7380,N_5067,N_4580);
nand U7381 (N_7381,N_4909,N_4914);
nor U7382 (N_7382,N_4885,N_3515);
nand U7383 (N_7383,N_4749,N_3422);
nand U7384 (N_7384,N_5263,N_4999);
or U7385 (N_7385,N_3583,N_6058);
nand U7386 (N_7386,N_4604,N_5637);
nor U7387 (N_7387,N_4831,N_3648);
and U7388 (N_7388,N_4422,N_3467);
nand U7389 (N_7389,N_4590,N_6102);
and U7390 (N_7390,N_3162,N_3823);
nor U7391 (N_7391,N_5759,N_5657);
nand U7392 (N_7392,N_5961,N_3797);
and U7393 (N_7393,N_5960,N_5264);
xnor U7394 (N_7394,N_4333,N_3373);
and U7395 (N_7395,N_4778,N_4027);
and U7396 (N_7396,N_5042,N_4356);
and U7397 (N_7397,N_4170,N_3672);
nor U7398 (N_7398,N_5202,N_4531);
and U7399 (N_7399,N_4273,N_3717);
xor U7400 (N_7400,N_4772,N_4503);
nor U7401 (N_7401,N_5395,N_5804);
nor U7402 (N_7402,N_5123,N_5585);
or U7403 (N_7403,N_4790,N_4964);
or U7404 (N_7404,N_4329,N_3134);
or U7405 (N_7405,N_4145,N_5503);
nor U7406 (N_7406,N_4601,N_6100);
xor U7407 (N_7407,N_5282,N_4944);
or U7408 (N_7408,N_4458,N_4774);
nand U7409 (N_7409,N_5046,N_3170);
and U7410 (N_7410,N_4499,N_5616);
xor U7411 (N_7411,N_3956,N_5090);
or U7412 (N_7412,N_4821,N_4210);
and U7413 (N_7413,N_3708,N_3910);
and U7414 (N_7414,N_3600,N_3337);
nor U7415 (N_7415,N_3934,N_4739);
and U7416 (N_7416,N_4098,N_5798);
and U7417 (N_7417,N_5159,N_3344);
and U7418 (N_7418,N_5934,N_3461);
or U7419 (N_7419,N_4685,N_4482);
and U7420 (N_7420,N_5617,N_4034);
and U7421 (N_7421,N_5200,N_3292);
nand U7422 (N_7422,N_4446,N_5812);
nand U7423 (N_7423,N_3251,N_5444);
nor U7424 (N_7424,N_4089,N_5307);
xnor U7425 (N_7425,N_5526,N_4068);
or U7426 (N_7426,N_5135,N_4251);
and U7427 (N_7427,N_5575,N_5006);
and U7428 (N_7428,N_3499,N_3454);
nand U7429 (N_7429,N_5603,N_6152);
nor U7430 (N_7430,N_5486,N_6027);
nor U7431 (N_7431,N_4608,N_4502);
and U7432 (N_7432,N_6223,N_4481);
or U7433 (N_7433,N_5808,N_3437);
or U7434 (N_7434,N_5536,N_3254);
or U7435 (N_7435,N_4889,N_3384);
and U7436 (N_7436,N_3858,N_5146);
nor U7437 (N_7437,N_5306,N_4187);
or U7438 (N_7438,N_3919,N_5043);
or U7439 (N_7439,N_5775,N_4814);
or U7440 (N_7440,N_3597,N_3841);
nor U7441 (N_7441,N_5554,N_4065);
nand U7442 (N_7442,N_3392,N_6024);
or U7443 (N_7443,N_3298,N_5248);
or U7444 (N_7444,N_4493,N_4007);
and U7445 (N_7445,N_4376,N_3207);
and U7446 (N_7446,N_4745,N_6091);
nor U7447 (N_7447,N_5521,N_3451);
xnor U7448 (N_7448,N_3843,N_4627);
nand U7449 (N_7449,N_5284,N_4435);
and U7450 (N_7450,N_3198,N_4320);
nand U7451 (N_7451,N_4092,N_5906);
or U7452 (N_7452,N_5457,N_3752);
and U7453 (N_7453,N_3981,N_3459);
and U7454 (N_7454,N_5894,N_4415);
and U7455 (N_7455,N_5814,N_4629);
nand U7456 (N_7456,N_6185,N_4404);
nor U7457 (N_7457,N_3918,N_3458);
xor U7458 (N_7458,N_5511,N_5190);
and U7459 (N_7459,N_4823,N_5625);
nor U7460 (N_7460,N_5907,N_4906);
or U7461 (N_7461,N_4294,N_4529);
nand U7462 (N_7462,N_4326,N_6010);
and U7463 (N_7463,N_3407,N_3845);
and U7464 (N_7464,N_5339,N_3905);
nor U7465 (N_7465,N_5172,N_3144);
and U7466 (N_7466,N_4468,N_4861);
xnor U7467 (N_7467,N_3639,N_5623);
or U7468 (N_7468,N_4728,N_4275);
or U7469 (N_7469,N_4589,N_3719);
xnor U7470 (N_7470,N_4301,N_3955);
or U7471 (N_7471,N_3581,N_5553);
and U7472 (N_7472,N_4787,N_4003);
nor U7473 (N_7473,N_4625,N_5925);
nor U7474 (N_7474,N_3350,N_3449);
nand U7475 (N_7475,N_3227,N_5459);
and U7476 (N_7476,N_4624,N_5421);
nand U7477 (N_7477,N_6022,N_3569);
xor U7478 (N_7478,N_4815,N_6169);
and U7479 (N_7479,N_4899,N_6034);
nand U7480 (N_7480,N_3376,N_4672);
or U7481 (N_7481,N_4675,N_3762);
nor U7482 (N_7482,N_5976,N_3242);
nand U7483 (N_7483,N_3503,N_5607);
or U7484 (N_7484,N_4196,N_5887);
nand U7485 (N_7485,N_5569,N_5353);
and U7486 (N_7486,N_4615,N_3330);
nand U7487 (N_7487,N_4900,N_3593);
nand U7488 (N_7488,N_4510,N_3638);
and U7489 (N_7489,N_4221,N_6057);
nand U7490 (N_7490,N_4245,N_5669);
or U7491 (N_7491,N_3678,N_5041);
and U7492 (N_7492,N_4507,N_4159);
or U7493 (N_7493,N_3809,N_3655);
and U7494 (N_7494,N_3831,N_4834);
and U7495 (N_7495,N_4449,N_4813);
xnor U7496 (N_7496,N_5011,N_4116);
and U7497 (N_7497,N_3889,N_3130);
nor U7498 (N_7498,N_5955,N_5145);
and U7499 (N_7499,N_4432,N_5688);
nor U7500 (N_7500,N_3611,N_3875);
and U7501 (N_7501,N_3771,N_5291);
or U7502 (N_7502,N_5436,N_4464);
nand U7503 (N_7503,N_4966,N_4213);
nand U7504 (N_7504,N_3186,N_4412);
nor U7505 (N_7505,N_3456,N_3282);
and U7506 (N_7506,N_4798,N_4355);
or U7507 (N_7507,N_3795,N_3805);
and U7508 (N_7508,N_4619,N_3800);
or U7509 (N_7509,N_5702,N_4336);
nand U7510 (N_7510,N_4535,N_4365);
and U7511 (N_7511,N_3764,N_3788);
and U7512 (N_7512,N_3603,N_4029);
nand U7513 (N_7513,N_6146,N_6059);
or U7514 (N_7514,N_3402,N_6121);
or U7515 (N_7515,N_3187,N_3518);
nor U7516 (N_7516,N_3312,N_4811);
and U7517 (N_7517,N_3888,N_3792);
nor U7518 (N_7518,N_3755,N_3685);
or U7519 (N_7519,N_4833,N_3694);
nor U7520 (N_7520,N_3998,N_5590);
and U7521 (N_7521,N_4674,N_3907);
nor U7522 (N_7522,N_4578,N_5994);
and U7523 (N_7523,N_4006,N_3768);
nor U7524 (N_7524,N_4949,N_3393);
or U7525 (N_7525,N_4667,N_4366);
nor U7526 (N_7526,N_5897,N_4657);
nand U7527 (N_7527,N_5990,N_3255);
and U7528 (N_7528,N_4407,N_4854);
nor U7529 (N_7529,N_5876,N_3757);
or U7530 (N_7530,N_4852,N_5920);
xnor U7531 (N_7531,N_4025,N_6106);
or U7532 (N_7532,N_5313,N_6026);
and U7533 (N_7533,N_4696,N_4423);
xor U7534 (N_7534,N_3586,N_4773);
xnor U7535 (N_7535,N_4955,N_3960);
and U7536 (N_7536,N_3146,N_5697);
nand U7537 (N_7537,N_4199,N_4670);
xor U7538 (N_7538,N_4717,N_4678);
or U7539 (N_7539,N_4472,N_4983);
nand U7540 (N_7540,N_4662,N_3190);
or U7541 (N_7541,N_5986,N_4226);
and U7542 (N_7542,N_3947,N_4332);
nand U7543 (N_7543,N_3760,N_3149);
or U7544 (N_7544,N_3590,N_4636);
nand U7545 (N_7545,N_5133,N_4017);
or U7546 (N_7546,N_4700,N_4205);
nand U7547 (N_7547,N_4921,N_3536);
or U7548 (N_7548,N_5844,N_5317);
and U7549 (N_7549,N_4977,N_3188);
or U7550 (N_7550,N_6098,N_3504);
and U7551 (N_7551,N_4919,N_5462);
nor U7552 (N_7552,N_4343,N_5597);
nor U7553 (N_7553,N_4501,N_3885);
nand U7554 (N_7554,N_4304,N_3688);
and U7555 (N_7555,N_4984,N_5572);
nand U7556 (N_7556,N_5115,N_4186);
nor U7557 (N_7557,N_5297,N_3386);
and U7558 (N_7558,N_5777,N_3457);
nor U7559 (N_7559,N_3229,N_4431);
nor U7560 (N_7560,N_4928,N_3653);
and U7561 (N_7561,N_5054,N_6001);
nand U7562 (N_7562,N_3128,N_5548);
xnor U7563 (N_7563,N_5274,N_4827);
nand U7564 (N_7564,N_3370,N_3406);
and U7565 (N_7565,N_5781,N_4572);
or U7566 (N_7566,N_3936,N_4838);
nor U7567 (N_7567,N_5679,N_6172);
xnor U7568 (N_7568,N_3690,N_4067);
nor U7569 (N_7569,N_4742,N_4397);
and U7570 (N_7570,N_3588,N_4602);
nand U7571 (N_7571,N_4425,N_3310);
nor U7572 (N_7572,N_4227,N_3912);
or U7573 (N_7573,N_4075,N_5183);
and U7574 (N_7574,N_4348,N_5026);
nor U7575 (N_7575,N_5765,N_4217);
nor U7576 (N_7576,N_3279,N_5015);
or U7577 (N_7577,N_3346,N_4300);
xnor U7578 (N_7578,N_3427,N_5799);
and U7579 (N_7579,N_4228,N_4402);
nand U7580 (N_7580,N_4307,N_3775);
and U7581 (N_7581,N_4897,N_4562);
or U7582 (N_7582,N_5935,N_5665);
nand U7583 (N_7583,N_3191,N_4560);
nor U7584 (N_7584,N_4496,N_5161);
nor U7585 (N_7585,N_5089,N_3887);
nor U7586 (N_7586,N_3484,N_3510);
nor U7587 (N_7587,N_5340,N_5883);
xnor U7588 (N_7588,N_3419,N_4485);
and U7589 (N_7589,N_4666,N_3866);
and U7590 (N_7590,N_3631,N_3806);
xnor U7591 (N_7591,N_5334,N_5075);
or U7592 (N_7592,N_3253,N_5892);
and U7593 (N_7593,N_5477,N_5639);
nand U7594 (N_7594,N_4290,N_6180);
nand U7595 (N_7595,N_4416,N_6219);
nor U7596 (N_7596,N_5922,N_5634);
or U7597 (N_7597,N_3415,N_5277);
xnor U7598 (N_7598,N_5423,N_5139);
nor U7599 (N_7599,N_5441,N_6188);
and U7600 (N_7600,N_4953,N_3997);
nand U7601 (N_7601,N_5758,N_3411);
or U7602 (N_7602,N_4445,N_5034);
nand U7603 (N_7603,N_3276,N_4669);
nor U7604 (N_7604,N_3290,N_4002);
or U7605 (N_7605,N_3347,N_4328);
nor U7606 (N_7606,N_4500,N_3668);
and U7607 (N_7607,N_5129,N_3579);
xnor U7608 (N_7608,N_6007,N_4714);
and U7609 (N_7609,N_5785,N_6164);
nor U7610 (N_7610,N_5850,N_5391);
and U7611 (N_7611,N_3287,N_3696);
or U7612 (N_7612,N_3573,N_3548);
xor U7613 (N_7613,N_5056,N_4377);
and U7614 (N_7614,N_5062,N_4219);
and U7615 (N_7615,N_4494,N_4441);
nand U7616 (N_7616,N_3793,N_6039);
nand U7617 (N_7617,N_3423,N_5126);
nand U7618 (N_7618,N_5707,N_4450);
xnor U7619 (N_7619,N_3922,N_3182);
nand U7620 (N_7620,N_4467,N_3285);
and U7621 (N_7621,N_4263,N_3133);
or U7622 (N_7622,N_5648,N_4430);
nor U7623 (N_7623,N_5852,N_4557);
or U7624 (N_7624,N_4741,N_6110);
and U7625 (N_7625,N_4085,N_3143);
nor U7626 (N_7626,N_5050,N_6107);
nand U7627 (N_7627,N_6225,N_5330);
xor U7628 (N_7628,N_5499,N_5144);
and U7629 (N_7629,N_3269,N_4836);
and U7630 (N_7630,N_5489,N_4771);
nand U7631 (N_7631,N_3204,N_4765);
or U7632 (N_7632,N_4406,N_6170);
nand U7633 (N_7633,N_3742,N_3514);
nor U7634 (N_7634,N_4513,N_4735);
nand U7635 (N_7635,N_4639,N_6128);
or U7636 (N_7636,N_4153,N_5539);
or U7637 (N_7637,N_3181,N_6093);
and U7638 (N_7638,N_5743,N_5210);
nand U7639 (N_7639,N_5788,N_4961);
xor U7640 (N_7640,N_4960,N_6079);
and U7641 (N_7641,N_4843,N_5103);
xor U7642 (N_7642,N_5869,N_4840);
or U7643 (N_7643,N_5187,N_5900);
nand U7644 (N_7644,N_3320,N_5383);
nor U7645 (N_7645,N_3302,N_6125);
nor U7646 (N_7646,N_3489,N_4318);
or U7647 (N_7647,N_3267,N_4806);
and U7648 (N_7648,N_3572,N_5430);
nand U7649 (N_7649,N_4822,N_5325);
or U7650 (N_7650,N_3863,N_4788);
nor U7651 (N_7651,N_5916,N_4398);
or U7652 (N_7652,N_5359,N_3959);
nand U7653 (N_7653,N_3749,N_5817);
and U7654 (N_7654,N_4958,N_4204);
nor U7655 (N_7655,N_4268,N_3306);
xnor U7656 (N_7656,N_3663,N_4257);
and U7657 (N_7657,N_4232,N_5479);
or U7658 (N_7658,N_5910,N_3261);
or U7659 (N_7659,N_3608,N_4433);
and U7660 (N_7660,N_5194,N_5587);
nand U7661 (N_7661,N_3967,N_4877);
nor U7662 (N_7662,N_6104,N_6073);
or U7663 (N_7663,N_5652,N_5424);
and U7664 (N_7664,N_3497,N_4514);
nand U7665 (N_7665,N_4125,N_4211);
nor U7666 (N_7666,N_5000,N_3849);
nand U7667 (N_7667,N_6019,N_3763);
and U7668 (N_7668,N_3531,N_5653);
and U7669 (N_7669,N_4359,N_5791);
nand U7670 (N_7670,N_3824,N_5638);
or U7671 (N_7671,N_4647,N_5570);
and U7672 (N_7672,N_6051,N_3750);
and U7673 (N_7673,N_4331,N_5721);
nor U7674 (N_7674,N_3539,N_5663);
or U7675 (N_7675,N_4408,N_5357);
nand U7676 (N_7676,N_3248,N_3739);
nand U7677 (N_7677,N_5241,N_3943);
nor U7678 (N_7678,N_3559,N_5222);
nand U7679 (N_7679,N_3622,N_5251);
xnor U7680 (N_7680,N_4867,N_3565);
and U7681 (N_7681,N_3477,N_4369);
or U7682 (N_7682,N_4302,N_4898);
or U7683 (N_7683,N_5861,N_4409);
nand U7684 (N_7684,N_3358,N_4444);
and U7685 (N_7685,N_3220,N_4684);
and U7686 (N_7686,N_3665,N_4106);
nand U7687 (N_7687,N_3389,N_5917);
and U7688 (N_7688,N_3669,N_4436);
nor U7689 (N_7689,N_5355,N_4154);
and U7690 (N_7690,N_3257,N_5438);
and U7691 (N_7691,N_5924,N_3286);
and U7692 (N_7692,N_5668,N_5176);
nor U7693 (N_7693,N_5824,N_3304);
and U7694 (N_7694,N_5069,N_4470);
nand U7695 (N_7695,N_3999,N_4568);
and U7696 (N_7696,N_6122,N_4695);
and U7697 (N_7697,N_6139,N_4280);
nand U7698 (N_7698,N_3643,N_5158);
and U7699 (N_7699,N_3173,N_4526);
or U7700 (N_7700,N_4901,N_3799);
and U7701 (N_7701,N_5356,N_6161);
and U7702 (N_7702,N_3904,N_3200);
nand U7703 (N_7703,N_3720,N_3326);
or U7704 (N_7704,N_3175,N_4593);
and U7705 (N_7705,N_6203,N_3246);
nand U7706 (N_7706,N_4164,N_5478);
nor U7707 (N_7707,N_4191,N_3167);
and U7708 (N_7708,N_4642,N_6082);
and U7709 (N_7709,N_5813,N_3262);
nor U7710 (N_7710,N_4043,N_3657);
or U7711 (N_7711,N_3340,N_4630);
nor U7712 (N_7712,N_3487,N_5290);
and U7713 (N_7713,N_5466,N_3214);
nor U7714 (N_7714,N_3985,N_3311);
nor U7715 (N_7715,N_3935,N_5984);
nor U7716 (N_7716,N_5091,N_6066);
nand U7717 (N_7717,N_5600,N_4368);
and U7718 (N_7718,N_5899,N_4230);
and U7719 (N_7719,N_5229,N_5100);
or U7720 (N_7720,N_4609,N_3896);
and U7721 (N_7721,N_4077,N_6095);
and U7722 (N_7722,N_3238,N_4171);
nor U7723 (N_7723,N_5816,N_3230);
and U7724 (N_7724,N_4567,N_4750);
nand U7725 (N_7725,N_4303,N_4347);
or U7726 (N_7726,N_5180,N_3412);
nor U7727 (N_7727,N_5319,N_4995);
or U7728 (N_7728,N_5647,N_3640);
or U7729 (N_7729,N_4600,N_4317);
nand U7730 (N_7730,N_5674,N_4527);
and U7731 (N_7731,N_3609,N_5516);
nand U7732 (N_7732,N_5449,N_4084);
and U7733 (N_7733,N_4309,N_5937);
and U7734 (N_7734,N_3353,N_4658);
and U7735 (N_7735,N_3335,N_5606);
nor U7736 (N_7736,N_3483,N_5364);
xor U7737 (N_7737,N_5783,N_5756);
or U7738 (N_7738,N_3401,N_4970);
and U7739 (N_7739,N_3532,N_3983);
and U7740 (N_7740,N_5094,N_4504);
or U7741 (N_7741,N_3923,N_4652);
and U7742 (N_7742,N_4797,N_5538);
nand U7743 (N_7743,N_5110,N_5573);
or U7744 (N_7744,N_4848,N_5755);
nor U7745 (N_7745,N_3211,N_3564);
or U7746 (N_7746,N_4870,N_4621);
nor U7747 (N_7747,N_5321,N_3260);
and U7748 (N_7748,N_4107,N_5498);
nand U7749 (N_7749,N_4617,N_6183);
or U7750 (N_7750,N_5452,N_3778);
nand U7751 (N_7751,N_4974,N_5396);
and U7752 (N_7752,N_3471,N_5502);
and U7753 (N_7753,N_6044,N_3562);
nand U7754 (N_7754,N_3275,N_5345);
xor U7755 (N_7755,N_4643,N_5909);
nor U7756 (N_7756,N_4484,N_4936);
and U7757 (N_7757,N_5057,N_4163);
nor U7758 (N_7758,N_4057,N_3827);
and U7759 (N_7759,N_5893,N_4549);
or U7760 (N_7760,N_3433,N_3615);
nor U7761 (N_7761,N_3416,N_5686);
or U7762 (N_7762,N_4166,N_6016);
xnor U7763 (N_7763,N_5645,N_3272);
nand U7764 (N_7764,N_4001,N_4283);
or U7765 (N_7765,N_4237,N_4722);
nand U7766 (N_7766,N_4142,N_6248);
or U7767 (N_7767,N_5433,N_3472);
nand U7768 (N_7768,N_5408,N_4028);
nand U7769 (N_7769,N_4768,N_3938);
nand U7770 (N_7770,N_3527,N_5780);
nand U7771 (N_7771,N_3381,N_5214);
nor U7772 (N_7772,N_4744,N_3265);
nand U7773 (N_7773,N_4754,N_4673);
nand U7774 (N_7774,N_3438,N_4184);
or U7775 (N_7775,N_4403,N_6000);
and U7776 (N_7776,N_3894,N_4760);
nand U7777 (N_7777,N_4932,N_4849);
or U7778 (N_7778,N_3811,N_4816);
xor U7779 (N_7779,N_5726,N_3410);
nor U7780 (N_7780,N_5061,N_3817);
and U7781 (N_7781,N_3530,N_3244);
or U7782 (N_7782,N_5283,N_4967);
nand U7783 (N_7783,N_4391,N_4401);
and U7784 (N_7784,N_5233,N_4871);
or U7785 (N_7785,N_5109,N_5113);
and U7786 (N_7786,N_5037,N_3250);
nor U7787 (N_7787,N_3926,N_4361);
xor U7788 (N_7788,N_5795,N_5628);
and U7789 (N_7789,N_5177,N_4973);
nand U7790 (N_7790,N_3606,N_4198);
nand U7791 (N_7791,N_4796,N_3740);
nand U7792 (N_7792,N_4563,N_4358);
or U7793 (N_7793,N_5368,N_4354);
xnor U7794 (N_7794,N_4509,N_4438);
and U7795 (N_7795,N_4314,N_4753);
xor U7796 (N_7796,N_3729,N_6076);
or U7797 (N_7797,N_5895,N_3766);
and U7798 (N_7798,N_3529,N_5065);
and U7799 (N_7799,N_3434,N_3158);
nor U7800 (N_7800,N_3671,N_4905);
nand U7801 (N_7801,N_4390,N_4249);
nor U7802 (N_7802,N_5589,N_5660);
and U7803 (N_7803,N_4711,N_5720);
and U7804 (N_7804,N_4046,N_3819);
nand U7805 (N_7805,N_4698,N_3691);
or U7806 (N_7806,N_3278,N_4063);
nand U7807 (N_7807,N_4632,N_4097);
nand U7808 (N_7808,N_6157,N_3784);
and U7809 (N_7809,N_3155,N_5296);
and U7810 (N_7810,N_6017,N_4310);
nor U7811 (N_7811,N_5846,N_4147);
nand U7812 (N_7812,N_3418,N_3450);
or U7813 (N_7813,N_5397,N_3522);
and U7814 (N_7814,N_4980,N_5719);
or U7815 (N_7815,N_4413,N_3834);
and U7816 (N_7816,N_4451,N_4480);
xnor U7817 (N_7817,N_6145,N_3430);
nor U7818 (N_7818,N_4624,N_3570);
nor U7819 (N_7819,N_5816,N_4715);
or U7820 (N_7820,N_6015,N_5038);
or U7821 (N_7821,N_6009,N_5622);
xor U7822 (N_7822,N_5963,N_4847);
and U7823 (N_7823,N_3315,N_3376);
or U7824 (N_7824,N_3878,N_4939);
nand U7825 (N_7825,N_5203,N_5995);
nor U7826 (N_7826,N_5190,N_3626);
nand U7827 (N_7827,N_3151,N_6128);
or U7828 (N_7828,N_5440,N_5855);
nand U7829 (N_7829,N_4645,N_3699);
nor U7830 (N_7830,N_4031,N_6090);
or U7831 (N_7831,N_4026,N_3260);
or U7832 (N_7832,N_5370,N_3587);
nand U7833 (N_7833,N_4040,N_3912);
nor U7834 (N_7834,N_5387,N_3423);
nand U7835 (N_7835,N_6151,N_4908);
or U7836 (N_7836,N_4126,N_3853);
nor U7837 (N_7837,N_4244,N_5249);
and U7838 (N_7838,N_4512,N_4325);
nor U7839 (N_7839,N_3308,N_4374);
or U7840 (N_7840,N_4323,N_4034);
nor U7841 (N_7841,N_3214,N_4071);
nor U7842 (N_7842,N_5493,N_4345);
or U7843 (N_7843,N_5343,N_3289);
and U7844 (N_7844,N_4780,N_6222);
xnor U7845 (N_7845,N_6105,N_4358);
nor U7846 (N_7846,N_3496,N_4542);
and U7847 (N_7847,N_3202,N_4764);
nand U7848 (N_7848,N_4349,N_3941);
or U7849 (N_7849,N_3907,N_3933);
or U7850 (N_7850,N_4376,N_6203);
and U7851 (N_7851,N_3202,N_4793);
or U7852 (N_7852,N_5635,N_4725);
and U7853 (N_7853,N_3794,N_4651);
nor U7854 (N_7854,N_3421,N_3587);
and U7855 (N_7855,N_3939,N_3336);
or U7856 (N_7856,N_4052,N_4567);
or U7857 (N_7857,N_3284,N_5247);
or U7858 (N_7858,N_4768,N_5341);
or U7859 (N_7859,N_4161,N_5535);
or U7860 (N_7860,N_4995,N_4822);
and U7861 (N_7861,N_4780,N_4665);
nand U7862 (N_7862,N_5075,N_5888);
nor U7863 (N_7863,N_3594,N_5942);
nand U7864 (N_7864,N_4840,N_4056);
nand U7865 (N_7865,N_3318,N_5317);
or U7866 (N_7866,N_3462,N_3585);
nand U7867 (N_7867,N_4029,N_5991);
and U7868 (N_7868,N_3198,N_5607);
nor U7869 (N_7869,N_3272,N_6238);
nand U7870 (N_7870,N_3973,N_5735);
and U7871 (N_7871,N_4974,N_5520);
nor U7872 (N_7872,N_5163,N_4260);
and U7873 (N_7873,N_5041,N_4770);
nand U7874 (N_7874,N_5504,N_5092);
or U7875 (N_7875,N_3796,N_5612);
or U7876 (N_7876,N_6198,N_5484);
xnor U7877 (N_7877,N_5373,N_3813);
nor U7878 (N_7878,N_3226,N_3568);
xor U7879 (N_7879,N_4760,N_4200);
nor U7880 (N_7880,N_5967,N_5773);
xor U7881 (N_7881,N_4766,N_4850);
and U7882 (N_7882,N_3511,N_3773);
or U7883 (N_7883,N_3975,N_5287);
or U7884 (N_7884,N_4868,N_5399);
nor U7885 (N_7885,N_3466,N_6086);
nand U7886 (N_7886,N_4065,N_5658);
xor U7887 (N_7887,N_4557,N_3877);
or U7888 (N_7888,N_5621,N_5995);
or U7889 (N_7889,N_5205,N_4312);
nand U7890 (N_7890,N_5677,N_3382);
nor U7891 (N_7891,N_5423,N_5865);
nand U7892 (N_7892,N_5088,N_3558);
and U7893 (N_7893,N_3218,N_4576);
and U7894 (N_7894,N_3393,N_4635);
nand U7895 (N_7895,N_3913,N_3917);
nand U7896 (N_7896,N_5546,N_5639);
and U7897 (N_7897,N_4961,N_3224);
and U7898 (N_7898,N_5621,N_3450);
nand U7899 (N_7899,N_3724,N_6185);
and U7900 (N_7900,N_5437,N_5915);
or U7901 (N_7901,N_4835,N_3266);
nor U7902 (N_7902,N_5169,N_5323);
nor U7903 (N_7903,N_4664,N_5721);
nor U7904 (N_7904,N_4637,N_5727);
or U7905 (N_7905,N_5094,N_3547);
nand U7906 (N_7906,N_5720,N_3738);
or U7907 (N_7907,N_4086,N_5241);
nand U7908 (N_7908,N_5415,N_5499);
or U7909 (N_7909,N_4155,N_4608);
xor U7910 (N_7910,N_4659,N_4209);
nor U7911 (N_7911,N_4407,N_6160);
nand U7912 (N_7912,N_3183,N_3833);
and U7913 (N_7913,N_5897,N_5848);
nand U7914 (N_7914,N_5192,N_3990);
nor U7915 (N_7915,N_4642,N_4874);
or U7916 (N_7916,N_5701,N_4025);
or U7917 (N_7917,N_6150,N_3259);
and U7918 (N_7918,N_5293,N_4458);
or U7919 (N_7919,N_4437,N_3530);
or U7920 (N_7920,N_4471,N_4000);
nand U7921 (N_7921,N_5058,N_4861);
or U7922 (N_7922,N_3522,N_5271);
nor U7923 (N_7923,N_5583,N_5237);
and U7924 (N_7924,N_6021,N_4326);
or U7925 (N_7925,N_4475,N_6116);
and U7926 (N_7926,N_4532,N_5453);
or U7927 (N_7927,N_5887,N_5222);
nor U7928 (N_7928,N_5352,N_5233);
nor U7929 (N_7929,N_5792,N_3274);
and U7930 (N_7930,N_6041,N_4350);
and U7931 (N_7931,N_3731,N_3580);
or U7932 (N_7932,N_3419,N_3709);
nor U7933 (N_7933,N_5989,N_3812);
nor U7934 (N_7934,N_4803,N_5953);
and U7935 (N_7935,N_3253,N_5956);
nor U7936 (N_7936,N_4483,N_3530);
nor U7937 (N_7937,N_3921,N_6035);
or U7938 (N_7938,N_3178,N_5167);
and U7939 (N_7939,N_4476,N_3397);
xnor U7940 (N_7940,N_3335,N_4731);
xor U7941 (N_7941,N_6246,N_3968);
or U7942 (N_7942,N_6237,N_4538);
and U7943 (N_7943,N_5581,N_5043);
nor U7944 (N_7944,N_4819,N_4625);
nor U7945 (N_7945,N_4741,N_5046);
nand U7946 (N_7946,N_4515,N_3809);
nor U7947 (N_7947,N_3495,N_5979);
nor U7948 (N_7948,N_3196,N_4996);
nor U7949 (N_7949,N_6205,N_3884);
or U7950 (N_7950,N_5972,N_4883);
nor U7951 (N_7951,N_6210,N_4367);
nor U7952 (N_7952,N_5668,N_3260);
xor U7953 (N_7953,N_3799,N_6128);
xnor U7954 (N_7954,N_4751,N_5667);
nor U7955 (N_7955,N_4244,N_5451);
and U7956 (N_7956,N_3979,N_5435);
or U7957 (N_7957,N_3913,N_3512);
and U7958 (N_7958,N_3283,N_4663);
nand U7959 (N_7959,N_4686,N_4798);
nor U7960 (N_7960,N_5271,N_5526);
nor U7961 (N_7961,N_3665,N_5658);
nor U7962 (N_7962,N_4295,N_3527);
nor U7963 (N_7963,N_3607,N_6082);
nand U7964 (N_7964,N_3310,N_5897);
or U7965 (N_7965,N_5130,N_4608);
and U7966 (N_7966,N_4449,N_4375);
and U7967 (N_7967,N_3962,N_5718);
or U7968 (N_7968,N_3312,N_3420);
and U7969 (N_7969,N_4956,N_6044);
nor U7970 (N_7970,N_5592,N_5407);
nand U7971 (N_7971,N_5798,N_5254);
nor U7972 (N_7972,N_4920,N_4719);
nand U7973 (N_7973,N_5049,N_3824);
nand U7974 (N_7974,N_5993,N_6223);
xor U7975 (N_7975,N_5386,N_6153);
or U7976 (N_7976,N_4270,N_5863);
and U7977 (N_7977,N_4067,N_5847);
nand U7978 (N_7978,N_3691,N_5666);
nand U7979 (N_7979,N_3396,N_4128);
and U7980 (N_7980,N_5453,N_3653);
xor U7981 (N_7981,N_6159,N_4217);
or U7982 (N_7982,N_4969,N_4459);
nor U7983 (N_7983,N_5196,N_4551);
and U7984 (N_7984,N_5054,N_3497);
or U7985 (N_7985,N_6175,N_4565);
nor U7986 (N_7986,N_4113,N_3824);
nand U7987 (N_7987,N_3811,N_3307);
nand U7988 (N_7988,N_4828,N_4739);
nand U7989 (N_7989,N_5028,N_3373);
nor U7990 (N_7990,N_3289,N_3768);
xnor U7991 (N_7991,N_5164,N_4485);
or U7992 (N_7992,N_4169,N_3732);
nor U7993 (N_7993,N_5807,N_5621);
or U7994 (N_7994,N_6013,N_5994);
nand U7995 (N_7995,N_3533,N_6109);
nor U7996 (N_7996,N_6094,N_5936);
or U7997 (N_7997,N_3795,N_4323);
and U7998 (N_7998,N_4381,N_4762);
or U7999 (N_7999,N_4940,N_5560);
nor U8000 (N_8000,N_3491,N_5806);
or U8001 (N_8001,N_5954,N_5525);
and U8002 (N_8002,N_5420,N_5158);
or U8003 (N_8003,N_6202,N_5563);
nor U8004 (N_8004,N_3590,N_3710);
and U8005 (N_8005,N_4927,N_4931);
and U8006 (N_8006,N_4353,N_5303);
and U8007 (N_8007,N_3999,N_6194);
or U8008 (N_8008,N_4924,N_4635);
or U8009 (N_8009,N_4355,N_4895);
nand U8010 (N_8010,N_3750,N_3903);
nand U8011 (N_8011,N_3873,N_5261);
and U8012 (N_8012,N_6120,N_4877);
and U8013 (N_8013,N_5925,N_5961);
and U8014 (N_8014,N_6244,N_6092);
nand U8015 (N_8015,N_5140,N_3132);
nand U8016 (N_8016,N_3526,N_5683);
or U8017 (N_8017,N_5206,N_3259);
nand U8018 (N_8018,N_3710,N_4733);
nand U8019 (N_8019,N_4415,N_3663);
nor U8020 (N_8020,N_5661,N_4337);
or U8021 (N_8021,N_5776,N_5565);
or U8022 (N_8022,N_5135,N_6130);
xor U8023 (N_8023,N_4730,N_5723);
and U8024 (N_8024,N_3178,N_5918);
nand U8025 (N_8025,N_4409,N_4096);
nor U8026 (N_8026,N_4396,N_3820);
or U8027 (N_8027,N_3765,N_5693);
nand U8028 (N_8028,N_4333,N_6183);
and U8029 (N_8029,N_5948,N_4355);
and U8030 (N_8030,N_4183,N_4337);
or U8031 (N_8031,N_5931,N_4863);
or U8032 (N_8032,N_4319,N_5933);
and U8033 (N_8033,N_5716,N_4993);
nand U8034 (N_8034,N_3266,N_4508);
or U8035 (N_8035,N_3423,N_4677);
nand U8036 (N_8036,N_5553,N_5192);
nor U8037 (N_8037,N_4845,N_4302);
xor U8038 (N_8038,N_3266,N_4999);
or U8039 (N_8039,N_4938,N_5287);
and U8040 (N_8040,N_6209,N_4764);
and U8041 (N_8041,N_4703,N_4478);
or U8042 (N_8042,N_4730,N_5347);
and U8043 (N_8043,N_6057,N_6201);
nand U8044 (N_8044,N_4675,N_4978);
and U8045 (N_8045,N_4437,N_3725);
or U8046 (N_8046,N_5895,N_6231);
xor U8047 (N_8047,N_4113,N_3802);
and U8048 (N_8048,N_5161,N_4879);
nor U8049 (N_8049,N_5574,N_5013);
nor U8050 (N_8050,N_5030,N_3630);
nand U8051 (N_8051,N_5866,N_4923);
nor U8052 (N_8052,N_4803,N_4610);
or U8053 (N_8053,N_5433,N_5787);
xor U8054 (N_8054,N_4259,N_4048);
and U8055 (N_8055,N_3983,N_4733);
xor U8056 (N_8056,N_3348,N_3133);
and U8057 (N_8057,N_3994,N_3956);
xnor U8058 (N_8058,N_3610,N_3447);
and U8059 (N_8059,N_3415,N_3781);
nand U8060 (N_8060,N_5579,N_6028);
nand U8061 (N_8061,N_5753,N_5420);
and U8062 (N_8062,N_3826,N_5791);
nor U8063 (N_8063,N_5977,N_4862);
and U8064 (N_8064,N_4065,N_3128);
xnor U8065 (N_8065,N_6218,N_5299);
xnor U8066 (N_8066,N_5215,N_3857);
nand U8067 (N_8067,N_3647,N_5917);
nand U8068 (N_8068,N_4964,N_4938);
or U8069 (N_8069,N_4254,N_5498);
xor U8070 (N_8070,N_3430,N_4831);
nor U8071 (N_8071,N_5366,N_6202);
nor U8072 (N_8072,N_4335,N_5127);
and U8073 (N_8073,N_3226,N_4268);
nor U8074 (N_8074,N_6214,N_4438);
nor U8075 (N_8075,N_6031,N_4930);
and U8076 (N_8076,N_5564,N_5705);
and U8077 (N_8077,N_5656,N_3952);
or U8078 (N_8078,N_5578,N_4273);
nand U8079 (N_8079,N_5092,N_5835);
or U8080 (N_8080,N_5750,N_3867);
and U8081 (N_8081,N_4226,N_4373);
nand U8082 (N_8082,N_3341,N_3146);
or U8083 (N_8083,N_4438,N_4262);
nand U8084 (N_8084,N_5048,N_5012);
or U8085 (N_8085,N_4313,N_3467);
xor U8086 (N_8086,N_5445,N_6037);
and U8087 (N_8087,N_5758,N_3891);
nand U8088 (N_8088,N_5158,N_5021);
and U8089 (N_8089,N_3189,N_4966);
and U8090 (N_8090,N_6125,N_3949);
nand U8091 (N_8091,N_3327,N_3494);
and U8092 (N_8092,N_3168,N_4917);
and U8093 (N_8093,N_6237,N_4412);
nor U8094 (N_8094,N_5068,N_4670);
and U8095 (N_8095,N_5136,N_4589);
nand U8096 (N_8096,N_5599,N_5350);
nand U8097 (N_8097,N_5458,N_3708);
or U8098 (N_8098,N_6001,N_4383);
nand U8099 (N_8099,N_6049,N_4055);
or U8100 (N_8100,N_3996,N_3762);
and U8101 (N_8101,N_3790,N_3464);
nor U8102 (N_8102,N_5143,N_3657);
nand U8103 (N_8103,N_5605,N_5505);
nand U8104 (N_8104,N_3688,N_5094);
xor U8105 (N_8105,N_5965,N_3638);
nor U8106 (N_8106,N_5654,N_3491);
or U8107 (N_8107,N_5387,N_4358);
and U8108 (N_8108,N_5855,N_4856);
and U8109 (N_8109,N_3372,N_3227);
nor U8110 (N_8110,N_6183,N_5584);
xor U8111 (N_8111,N_4795,N_4657);
or U8112 (N_8112,N_3515,N_5118);
and U8113 (N_8113,N_5065,N_3570);
nand U8114 (N_8114,N_5556,N_3171);
nand U8115 (N_8115,N_3970,N_6055);
or U8116 (N_8116,N_3854,N_3467);
nand U8117 (N_8117,N_4538,N_5345);
or U8118 (N_8118,N_4914,N_5480);
and U8119 (N_8119,N_5325,N_4108);
nor U8120 (N_8120,N_3449,N_3772);
nor U8121 (N_8121,N_3126,N_3988);
and U8122 (N_8122,N_6030,N_4616);
or U8123 (N_8123,N_6172,N_3808);
xnor U8124 (N_8124,N_4663,N_3253);
or U8125 (N_8125,N_4540,N_5525);
nand U8126 (N_8126,N_5794,N_5641);
and U8127 (N_8127,N_6152,N_4929);
nor U8128 (N_8128,N_5271,N_4258);
and U8129 (N_8129,N_3180,N_6032);
or U8130 (N_8130,N_4935,N_4714);
and U8131 (N_8131,N_3150,N_5208);
or U8132 (N_8132,N_4172,N_5188);
nor U8133 (N_8133,N_5638,N_5481);
nand U8134 (N_8134,N_5213,N_3456);
nor U8135 (N_8135,N_5641,N_4639);
and U8136 (N_8136,N_3385,N_3686);
xor U8137 (N_8137,N_6038,N_4688);
nand U8138 (N_8138,N_3997,N_4409);
nor U8139 (N_8139,N_3378,N_5736);
or U8140 (N_8140,N_3878,N_4887);
nor U8141 (N_8141,N_4162,N_4906);
nor U8142 (N_8142,N_3670,N_3375);
nor U8143 (N_8143,N_4376,N_3358);
and U8144 (N_8144,N_5680,N_6223);
nand U8145 (N_8145,N_5588,N_4126);
or U8146 (N_8146,N_3597,N_3875);
nand U8147 (N_8147,N_6142,N_3725);
and U8148 (N_8148,N_4161,N_3227);
or U8149 (N_8149,N_6043,N_3978);
nand U8150 (N_8150,N_5664,N_5880);
or U8151 (N_8151,N_3340,N_5371);
xnor U8152 (N_8152,N_3280,N_6142);
nand U8153 (N_8153,N_3293,N_3457);
nand U8154 (N_8154,N_5889,N_6099);
nor U8155 (N_8155,N_6060,N_3660);
nand U8156 (N_8156,N_5466,N_5420);
nor U8157 (N_8157,N_4773,N_3779);
nand U8158 (N_8158,N_5754,N_3933);
or U8159 (N_8159,N_5391,N_5086);
nand U8160 (N_8160,N_6129,N_6084);
nor U8161 (N_8161,N_4339,N_5245);
nand U8162 (N_8162,N_4135,N_4216);
and U8163 (N_8163,N_5270,N_4698);
or U8164 (N_8164,N_3139,N_3704);
nand U8165 (N_8165,N_5028,N_3742);
nand U8166 (N_8166,N_3978,N_3385);
nand U8167 (N_8167,N_5699,N_4192);
or U8168 (N_8168,N_4907,N_4868);
and U8169 (N_8169,N_5324,N_3825);
or U8170 (N_8170,N_5787,N_3456);
and U8171 (N_8171,N_5798,N_4487);
and U8172 (N_8172,N_4671,N_5720);
xor U8173 (N_8173,N_4912,N_6210);
and U8174 (N_8174,N_4752,N_5633);
or U8175 (N_8175,N_3456,N_6130);
and U8176 (N_8176,N_4526,N_4208);
nand U8177 (N_8177,N_6147,N_4792);
xnor U8178 (N_8178,N_3913,N_5140);
or U8179 (N_8179,N_3281,N_5567);
nand U8180 (N_8180,N_4281,N_6040);
xnor U8181 (N_8181,N_3348,N_4314);
nand U8182 (N_8182,N_3370,N_5414);
nor U8183 (N_8183,N_4350,N_3234);
or U8184 (N_8184,N_5408,N_4795);
or U8185 (N_8185,N_4835,N_5808);
or U8186 (N_8186,N_3403,N_5231);
nand U8187 (N_8187,N_3913,N_3740);
and U8188 (N_8188,N_5285,N_4891);
nand U8189 (N_8189,N_5228,N_4717);
nand U8190 (N_8190,N_5915,N_3737);
nand U8191 (N_8191,N_3769,N_5017);
nor U8192 (N_8192,N_4530,N_3921);
or U8193 (N_8193,N_3478,N_3927);
or U8194 (N_8194,N_3165,N_4152);
and U8195 (N_8195,N_4567,N_5690);
nor U8196 (N_8196,N_6156,N_3701);
nand U8197 (N_8197,N_4758,N_3365);
or U8198 (N_8198,N_3948,N_4928);
nor U8199 (N_8199,N_3477,N_5193);
and U8200 (N_8200,N_3697,N_5656);
or U8201 (N_8201,N_4557,N_3845);
nand U8202 (N_8202,N_4867,N_5610);
nand U8203 (N_8203,N_5092,N_3646);
or U8204 (N_8204,N_6011,N_5529);
xnor U8205 (N_8205,N_3158,N_5115);
and U8206 (N_8206,N_5945,N_3785);
nor U8207 (N_8207,N_3788,N_3560);
and U8208 (N_8208,N_4088,N_3835);
or U8209 (N_8209,N_3450,N_5537);
and U8210 (N_8210,N_4807,N_3281);
nand U8211 (N_8211,N_6171,N_3882);
nor U8212 (N_8212,N_4329,N_4833);
nand U8213 (N_8213,N_5487,N_4136);
or U8214 (N_8214,N_3593,N_4015);
xnor U8215 (N_8215,N_3266,N_3933);
nand U8216 (N_8216,N_4394,N_3125);
nor U8217 (N_8217,N_6162,N_6218);
nor U8218 (N_8218,N_3623,N_5375);
xnor U8219 (N_8219,N_3445,N_5332);
xor U8220 (N_8220,N_5426,N_5203);
nor U8221 (N_8221,N_4192,N_6089);
and U8222 (N_8222,N_5201,N_3332);
or U8223 (N_8223,N_5439,N_6129);
nand U8224 (N_8224,N_4071,N_3453);
nand U8225 (N_8225,N_3229,N_4227);
or U8226 (N_8226,N_5060,N_4601);
nand U8227 (N_8227,N_3912,N_5254);
nand U8228 (N_8228,N_3433,N_4060);
nand U8229 (N_8229,N_5402,N_3626);
nor U8230 (N_8230,N_5843,N_3945);
nor U8231 (N_8231,N_5609,N_4666);
and U8232 (N_8232,N_4663,N_4550);
nor U8233 (N_8233,N_3282,N_5075);
or U8234 (N_8234,N_5661,N_5140);
and U8235 (N_8235,N_5813,N_4962);
or U8236 (N_8236,N_4630,N_4115);
xor U8237 (N_8237,N_5127,N_5882);
nand U8238 (N_8238,N_3957,N_3205);
and U8239 (N_8239,N_6172,N_3825);
or U8240 (N_8240,N_6229,N_3251);
nand U8241 (N_8241,N_4178,N_3282);
nand U8242 (N_8242,N_3176,N_4674);
and U8243 (N_8243,N_5634,N_3367);
or U8244 (N_8244,N_4508,N_4908);
nand U8245 (N_8245,N_4840,N_4820);
nor U8246 (N_8246,N_4058,N_3402);
nor U8247 (N_8247,N_5260,N_5411);
nand U8248 (N_8248,N_4484,N_5999);
xor U8249 (N_8249,N_5549,N_3632);
or U8250 (N_8250,N_4095,N_5207);
nor U8251 (N_8251,N_4034,N_5148);
nand U8252 (N_8252,N_4636,N_5280);
nor U8253 (N_8253,N_5862,N_3179);
and U8254 (N_8254,N_3212,N_4948);
xor U8255 (N_8255,N_4392,N_5802);
nand U8256 (N_8256,N_4652,N_4237);
or U8257 (N_8257,N_5262,N_5979);
nor U8258 (N_8258,N_3647,N_4697);
nand U8259 (N_8259,N_5297,N_3431);
or U8260 (N_8260,N_5093,N_5201);
nand U8261 (N_8261,N_4833,N_5002);
nand U8262 (N_8262,N_4315,N_5277);
and U8263 (N_8263,N_4180,N_4268);
and U8264 (N_8264,N_4729,N_5196);
and U8265 (N_8265,N_5831,N_3218);
nor U8266 (N_8266,N_4798,N_3168);
or U8267 (N_8267,N_5109,N_4879);
nand U8268 (N_8268,N_3736,N_4184);
and U8269 (N_8269,N_4718,N_5690);
or U8270 (N_8270,N_4183,N_3438);
xor U8271 (N_8271,N_4920,N_4671);
nor U8272 (N_8272,N_5380,N_5172);
xor U8273 (N_8273,N_3237,N_5966);
or U8274 (N_8274,N_5298,N_4042);
xor U8275 (N_8275,N_4711,N_4579);
and U8276 (N_8276,N_5240,N_3707);
nand U8277 (N_8277,N_5391,N_4351);
nor U8278 (N_8278,N_4406,N_3920);
nand U8279 (N_8279,N_6098,N_3312);
xor U8280 (N_8280,N_4507,N_5380);
and U8281 (N_8281,N_5418,N_4724);
nor U8282 (N_8282,N_4754,N_5550);
nand U8283 (N_8283,N_5032,N_6186);
or U8284 (N_8284,N_4920,N_4366);
nor U8285 (N_8285,N_3788,N_4863);
or U8286 (N_8286,N_4681,N_5387);
and U8287 (N_8287,N_3153,N_5115);
and U8288 (N_8288,N_4947,N_3839);
xor U8289 (N_8289,N_5646,N_5941);
nand U8290 (N_8290,N_4961,N_3953);
and U8291 (N_8291,N_4438,N_5564);
nor U8292 (N_8292,N_4384,N_5028);
and U8293 (N_8293,N_6237,N_4838);
or U8294 (N_8294,N_3461,N_3552);
and U8295 (N_8295,N_4994,N_5986);
and U8296 (N_8296,N_5320,N_3850);
and U8297 (N_8297,N_4934,N_3536);
xnor U8298 (N_8298,N_3249,N_5295);
and U8299 (N_8299,N_4223,N_4525);
nor U8300 (N_8300,N_3270,N_5297);
nor U8301 (N_8301,N_3242,N_6005);
nor U8302 (N_8302,N_4572,N_5648);
xor U8303 (N_8303,N_5547,N_3847);
nand U8304 (N_8304,N_4484,N_5619);
nand U8305 (N_8305,N_6245,N_5826);
nand U8306 (N_8306,N_5595,N_4431);
xor U8307 (N_8307,N_4936,N_5416);
and U8308 (N_8308,N_3308,N_4750);
nand U8309 (N_8309,N_3953,N_4280);
nand U8310 (N_8310,N_4533,N_5333);
xnor U8311 (N_8311,N_4872,N_3824);
nor U8312 (N_8312,N_6116,N_4473);
nor U8313 (N_8313,N_4690,N_4304);
and U8314 (N_8314,N_5873,N_4281);
nand U8315 (N_8315,N_4171,N_3205);
or U8316 (N_8316,N_5604,N_4815);
and U8317 (N_8317,N_6207,N_4533);
nand U8318 (N_8318,N_4449,N_4258);
nand U8319 (N_8319,N_4980,N_4953);
nor U8320 (N_8320,N_3290,N_6108);
nand U8321 (N_8321,N_3751,N_5049);
nor U8322 (N_8322,N_4811,N_5056);
or U8323 (N_8323,N_3733,N_3391);
xor U8324 (N_8324,N_3914,N_3252);
nor U8325 (N_8325,N_5788,N_5974);
and U8326 (N_8326,N_3733,N_3994);
nor U8327 (N_8327,N_3233,N_4982);
or U8328 (N_8328,N_3341,N_3390);
nand U8329 (N_8329,N_4122,N_5898);
nor U8330 (N_8330,N_3628,N_6094);
nor U8331 (N_8331,N_6000,N_5242);
or U8332 (N_8332,N_5572,N_5117);
nand U8333 (N_8333,N_4645,N_4042);
nor U8334 (N_8334,N_5918,N_4351);
or U8335 (N_8335,N_3985,N_4696);
nor U8336 (N_8336,N_3631,N_5637);
and U8337 (N_8337,N_4912,N_5168);
xor U8338 (N_8338,N_5366,N_5143);
nor U8339 (N_8339,N_3580,N_4356);
xor U8340 (N_8340,N_4584,N_3878);
or U8341 (N_8341,N_3848,N_4552);
nor U8342 (N_8342,N_4387,N_5590);
or U8343 (N_8343,N_4538,N_3278);
nor U8344 (N_8344,N_5836,N_3641);
nor U8345 (N_8345,N_3953,N_5066);
or U8346 (N_8346,N_3852,N_5662);
or U8347 (N_8347,N_3231,N_4213);
xor U8348 (N_8348,N_4898,N_3486);
nor U8349 (N_8349,N_4958,N_3311);
nor U8350 (N_8350,N_4857,N_4561);
and U8351 (N_8351,N_3480,N_3538);
and U8352 (N_8352,N_4548,N_5569);
nand U8353 (N_8353,N_3676,N_5933);
nor U8354 (N_8354,N_4701,N_4099);
or U8355 (N_8355,N_3134,N_4358);
nand U8356 (N_8356,N_3907,N_4181);
and U8357 (N_8357,N_4540,N_4726);
and U8358 (N_8358,N_5902,N_4116);
nand U8359 (N_8359,N_5237,N_6072);
nand U8360 (N_8360,N_4822,N_6170);
or U8361 (N_8361,N_3350,N_3844);
and U8362 (N_8362,N_5172,N_3280);
nor U8363 (N_8363,N_5891,N_6011);
and U8364 (N_8364,N_5449,N_5873);
or U8365 (N_8365,N_5790,N_4896);
xor U8366 (N_8366,N_4267,N_5464);
and U8367 (N_8367,N_5131,N_3741);
nand U8368 (N_8368,N_3821,N_4301);
and U8369 (N_8369,N_3289,N_3422);
and U8370 (N_8370,N_5098,N_4632);
and U8371 (N_8371,N_5285,N_4573);
nor U8372 (N_8372,N_6092,N_3968);
or U8373 (N_8373,N_3581,N_5397);
or U8374 (N_8374,N_4248,N_4216);
xor U8375 (N_8375,N_5734,N_3609);
nand U8376 (N_8376,N_5756,N_3356);
and U8377 (N_8377,N_5004,N_5088);
or U8378 (N_8378,N_3380,N_3946);
nor U8379 (N_8379,N_3333,N_5069);
and U8380 (N_8380,N_5362,N_5758);
or U8381 (N_8381,N_3483,N_6001);
and U8382 (N_8382,N_4176,N_5155);
xor U8383 (N_8383,N_5367,N_3313);
nor U8384 (N_8384,N_5576,N_3689);
nand U8385 (N_8385,N_5652,N_3793);
nand U8386 (N_8386,N_5640,N_3783);
and U8387 (N_8387,N_3620,N_3595);
and U8388 (N_8388,N_4195,N_4083);
and U8389 (N_8389,N_3301,N_3192);
nand U8390 (N_8390,N_5969,N_5051);
and U8391 (N_8391,N_3875,N_4923);
and U8392 (N_8392,N_6030,N_6172);
nand U8393 (N_8393,N_6073,N_4507);
nand U8394 (N_8394,N_5052,N_5586);
nand U8395 (N_8395,N_6249,N_5285);
or U8396 (N_8396,N_3977,N_5159);
nor U8397 (N_8397,N_5763,N_4334);
nand U8398 (N_8398,N_4641,N_3500);
and U8399 (N_8399,N_4504,N_3410);
or U8400 (N_8400,N_5547,N_5529);
nand U8401 (N_8401,N_4854,N_3591);
nand U8402 (N_8402,N_5850,N_5632);
xor U8403 (N_8403,N_5838,N_5073);
nand U8404 (N_8404,N_6084,N_5146);
nor U8405 (N_8405,N_4558,N_3350);
nand U8406 (N_8406,N_5676,N_3436);
and U8407 (N_8407,N_4941,N_5636);
xor U8408 (N_8408,N_3391,N_3244);
or U8409 (N_8409,N_5434,N_5601);
xnor U8410 (N_8410,N_3511,N_5376);
nor U8411 (N_8411,N_5378,N_4972);
nor U8412 (N_8412,N_4053,N_3391);
and U8413 (N_8413,N_5282,N_4005);
or U8414 (N_8414,N_4781,N_5615);
nand U8415 (N_8415,N_4537,N_6195);
or U8416 (N_8416,N_5600,N_4878);
nand U8417 (N_8417,N_3254,N_5401);
or U8418 (N_8418,N_3216,N_3310);
and U8419 (N_8419,N_5719,N_5046);
or U8420 (N_8420,N_4354,N_4006);
nand U8421 (N_8421,N_3948,N_4510);
nand U8422 (N_8422,N_5473,N_5114);
nor U8423 (N_8423,N_5723,N_5697);
xor U8424 (N_8424,N_4309,N_5627);
nor U8425 (N_8425,N_5183,N_4105);
nor U8426 (N_8426,N_5060,N_5605);
nand U8427 (N_8427,N_3126,N_3181);
xor U8428 (N_8428,N_6171,N_4450);
or U8429 (N_8429,N_5445,N_6019);
nor U8430 (N_8430,N_4200,N_4219);
xor U8431 (N_8431,N_5916,N_3552);
nor U8432 (N_8432,N_5629,N_5455);
and U8433 (N_8433,N_6243,N_4819);
nor U8434 (N_8434,N_3935,N_5370);
and U8435 (N_8435,N_6128,N_3139);
and U8436 (N_8436,N_3146,N_4138);
nor U8437 (N_8437,N_5786,N_3523);
nor U8438 (N_8438,N_6210,N_3605);
and U8439 (N_8439,N_6089,N_3857);
and U8440 (N_8440,N_3774,N_5404);
or U8441 (N_8441,N_5751,N_5877);
nand U8442 (N_8442,N_3535,N_3363);
xor U8443 (N_8443,N_6033,N_4523);
nor U8444 (N_8444,N_4911,N_4945);
or U8445 (N_8445,N_4074,N_4415);
nand U8446 (N_8446,N_3336,N_4542);
and U8447 (N_8447,N_4837,N_5072);
and U8448 (N_8448,N_6179,N_4007);
nand U8449 (N_8449,N_3330,N_4453);
and U8450 (N_8450,N_5502,N_5148);
nor U8451 (N_8451,N_6113,N_3313);
nor U8452 (N_8452,N_5811,N_3460);
nor U8453 (N_8453,N_6021,N_5176);
and U8454 (N_8454,N_5595,N_5828);
or U8455 (N_8455,N_4608,N_5448);
nand U8456 (N_8456,N_5996,N_3618);
or U8457 (N_8457,N_3280,N_6018);
or U8458 (N_8458,N_5078,N_4365);
nor U8459 (N_8459,N_5502,N_3656);
nor U8460 (N_8460,N_4591,N_3988);
and U8461 (N_8461,N_4911,N_4081);
or U8462 (N_8462,N_4486,N_3603);
nand U8463 (N_8463,N_6162,N_4056);
and U8464 (N_8464,N_6177,N_3758);
nor U8465 (N_8465,N_5446,N_3659);
or U8466 (N_8466,N_3690,N_4079);
nor U8467 (N_8467,N_4151,N_6093);
nor U8468 (N_8468,N_6221,N_6054);
and U8469 (N_8469,N_5977,N_5786);
and U8470 (N_8470,N_5805,N_6005);
nor U8471 (N_8471,N_4293,N_6075);
and U8472 (N_8472,N_3678,N_4153);
nor U8473 (N_8473,N_4825,N_4283);
xor U8474 (N_8474,N_4480,N_4706);
nand U8475 (N_8475,N_4551,N_3985);
and U8476 (N_8476,N_3230,N_3274);
and U8477 (N_8477,N_4568,N_4989);
and U8478 (N_8478,N_4350,N_3950);
xor U8479 (N_8479,N_3548,N_5824);
nor U8480 (N_8480,N_4782,N_4530);
nor U8481 (N_8481,N_5207,N_5895);
xnor U8482 (N_8482,N_6145,N_5686);
or U8483 (N_8483,N_3680,N_3756);
nand U8484 (N_8484,N_3569,N_3813);
nor U8485 (N_8485,N_4984,N_4478);
and U8486 (N_8486,N_6084,N_3379);
and U8487 (N_8487,N_5573,N_4072);
and U8488 (N_8488,N_5713,N_5045);
and U8489 (N_8489,N_5199,N_3453);
nand U8490 (N_8490,N_4340,N_5111);
and U8491 (N_8491,N_5451,N_5552);
or U8492 (N_8492,N_3277,N_4557);
nor U8493 (N_8493,N_3813,N_6024);
nand U8494 (N_8494,N_3416,N_4899);
nor U8495 (N_8495,N_4169,N_4464);
nor U8496 (N_8496,N_6168,N_5768);
xor U8497 (N_8497,N_3353,N_3581);
or U8498 (N_8498,N_3964,N_4234);
nor U8499 (N_8499,N_4181,N_3476);
and U8500 (N_8500,N_4928,N_6195);
nand U8501 (N_8501,N_3385,N_3293);
nand U8502 (N_8502,N_3192,N_3959);
nor U8503 (N_8503,N_6199,N_5615);
nand U8504 (N_8504,N_5351,N_5482);
nand U8505 (N_8505,N_4400,N_4346);
and U8506 (N_8506,N_3365,N_5221);
or U8507 (N_8507,N_4311,N_3828);
or U8508 (N_8508,N_3727,N_4272);
and U8509 (N_8509,N_5925,N_3315);
or U8510 (N_8510,N_3884,N_4080);
nand U8511 (N_8511,N_3753,N_3956);
or U8512 (N_8512,N_5398,N_6098);
or U8513 (N_8513,N_4262,N_4166);
and U8514 (N_8514,N_3806,N_3644);
or U8515 (N_8515,N_4414,N_4273);
nor U8516 (N_8516,N_4914,N_6179);
nor U8517 (N_8517,N_5245,N_6052);
nand U8518 (N_8518,N_4097,N_3192);
and U8519 (N_8519,N_5116,N_5944);
nor U8520 (N_8520,N_4787,N_6200);
or U8521 (N_8521,N_4966,N_3595);
and U8522 (N_8522,N_5198,N_4363);
nand U8523 (N_8523,N_5984,N_5893);
or U8524 (N_8524,N_4177,N_3882);
nand U8525 (N_8525,N_3792,N_3147);
xor U8526 (N_8526,N_4722,N_3322);
and U8527 (N_8527,N_5617,N_4772);
and U8528 (N_8528,N_4845,N_3912);
nand U8529 (N_8529,N_4473,N_4937);
or U8530 (N_8530,N_3816,N_3517);
nand U8531 (N_8531,N_3720,N_6058);
nand U8532 (N_8532,N_4614,N_3861);
and U8533 (N_8533,N_5759,N_4001);
nor U8534 (N_8534,N_3256,N_4963);
or U8535 (N_8535,N_4054,N_5354);
nor U8536 (N_8536,N_3643,N_3927);
and U8537 (N_8537,N_5209,N_5967);
nor U8538 (N_8538,N_4046,N_3540);
xnor U8539 (N_8539,N_3837,N_6217);
xor U8540 (N_8540,N_6090,N_6211);
nor U8541 (N_8541,N_5338,N_4796);
or U8542 (N_8542,N_4003,N_6002);
nand U8543 (N_8543,N_4572,N_5539);
and U8544 (N_8544,N_5252,N_4985);
nand U8545 (N_8545,N_5765,N_4514);
nand U8546 (N_8546,N_3570,N_6082);
and U8547 (N_8547,N_3240,N_4362);
nor U8548 (N_8548,N_3824,N_4564);
or U8549 (N_8549,N_4350,N_4435);
or U8550 (N_8550,N_4670,N_5207);
nor U8551 (N_8551,N_3368,N_3907);
nand U8552 (N_8552,N_4707,N_3719);
nand U8553 (N_8553,N_4903,N_3249);
and U8554 (N_8554,N_4266,N_4665);
or U8555 (N_8555,N_6172,N_5465);
nand U8556 (N_8556,N_3976,N_5989);
nand U8557 (N_8557,N_3414,N_4247);
nor U8558 (N_8558,N_4265,N_5569);
nand U8559 (N_8559,N_3238,N_5116);
and U8560 (N_8560,N_4160,N_4095);
or U8561 (N_8561,N_5487,N_3319);
nor U8562 (N_8562,N_3414,N_5837);
or U8563 (N_8563,N_6017,N_3485);
or U8564 (N_8564,N_5566,N_4128);
nor U8565 (N_8565,N_4702,N_5060);
nand U8566 (N_8566,N_3683,N_6057);
or U8567 (N_8567,N_5167,N_5002);
xnor U8568 (N_8568,N_4458,N_3326);
nand U8569 (N_8569,N_6192,N_5547);
xor U8570 (N_8570,N_5178,N_3351);
nand U8571 (N_8571,N_4863,N_3350);
nand U8572 (N_8572,N_5014,N_6011);
nand U8573 (N_8573,N_4486,N_3555);
or U8574 (N_8574,N_6233,N_4208);
nand U8575 (N_8575,N_3984,N_4220);
and U8576 (N_8576,N_6079,N_4289);
nor U8577 (N_8577,N_6032,N_3985);
nand U8578 (N_8578,N_4248,N_5607);
and U8579 (N_8579,N_4157,N_4871);
or U8580 (N_8580,N_4320,N_5039);
nand U8581 (N_8581,N_3988,N_6032);
xor U8582 (N_8582,N_5328,N_6048);
or U8583 (N_8583,N_4450,N_4136);
xor U8584 (N_8584,N_4599,N_4090);
nor U8585 (N_8585,N_5716,N_5045);
or U8586 (N_8586,N_4297,N_3390);
nand U8587 (N_8587,N_4986,N_5682);
nand U8588 (N_8588,N_4402,N_5752);
or U8589 (N_8589,N_5083,N_5867);
and U8590 (N_8590,N_6110,N_4537);
nor U8591 (N_8591,N_3490,N_3913);
nor U8592 (N_8592,N_5509,N_6032);
nor U8593 (N_8593,N_3811,N_4641);
nor U8594 (N_8594,N_4203,N_4942);
or U8595 (N_8595,N_5739,N_3576);
nand U8596 (N_8596,N_5979,N_5950);
nand U8597 (N_8597,N_3828,N_4757);
xnor U8598 (N_8598,N_5128,N_6190);
nand U8599 (N_8599,N_6003,N_5680);
nand U8600 (N_8600,N_5976,N_4840);
and U8601 (N_8601,N_3407,N_4568);
or U8602 (N_8602,N_5705,N_3519);
nand U8603 (N_8603,N_4822,N_3232);
nand U8604 (N_8604,N_5453,N_5683);
or U8605 (N_8605,N_3964,N_5486);
nand U8606 (N_8606,N_5861,N_4368);
and U8607 (N_8607,N_5117,N_3735);
or U8608 (N_8608,N_3525,N_3521);
nor U8609 (N_8609,N_3255,N_5898);
nor U8610 (N_8610,N_6109,N_4767);
xnor U8611 (N_8611,N_4344,N_4410);
nor U8612 (N_8612,N_5092,N_4941);
nor U8613 (N_8613,N_4804,N_3368);
nand U8614 (N_8614,N_4377,N_3174);
and U8615 (N_8615,N_3145,N_3603);
nand U8616 (N_8616,N_3621,N_5839);
nand U8617 (N_8617,N_6211,N_3921);
and U8618 (N_8618,N_4073,N_5008);
xor U8619 (N_8619,N_4323,N_5214);
xnor U8620 (N_8620,N_5760,N_5564);
nand U8621 (N_8621,N_4803,N_3180);
and U8622 (N_8622,N_6246,N_6023);
nand U8623 (N_8623,N_4047,N_3636);
and U8624 (N_8624,N_4212,N_3688);
nand U8625 (N_8625,N_5446,N_5140);
nand U8626 (N_8626,N_5549,N_5103);
or U8627 (N_8627,N_5524,N_3318);
nand U8628 (N_8628,N_4571,N_5297);
xor U8629 (N_8629,N_4404,N_4515);
nor U8630 (N_8630,N_5326,N_4338);
nand U8631 (N_8631,N_5345,N_3501);
and U8632 (N_8632,N_4528,N_3680);
nor U8633 (N_8633,N_6068,N_5850);
nand U8634 (N_8634,N_3315,N_5842);
nor U8635 (N_8635,N_5963,N_5888);
or U8636 (N_8636,N_5426,N_5936);
nor U8637 (N_8637,N_5587,N_3538);
nand U8638 (N_8638,N_3283,N_5000);
nand U8639 (N_8639,N_4929,N_3922);
or U8640 (N_8640,N_5011,N_5326);
or U8641 (N_8641,N_5834,N_5231);
nor U8642 (N_8642,N_4084,N_6177);
and U8643 (N_8643,N_5659,N_3377);
nand U8644 (N_8644,N_4912,N_4013);
or U8645 (N_8645,N_5341,N_3915);
nor U8646 (N_8646,N_4213,N_6003);
or U8647 (N_8647,N_4713,N_5313);
or U8648 (N_8648,N_3933,N_4716);
and U8649 (N_8649,N_5283,N_4697);
nand U8650 (N_8650,N_3726,N_4466);
and U8651 (N_8651,N_4377,N_4738);
nor U8652 (N_8652,N_4405,N_5154);
and U8653 (N_8653,N_4883,N_5277);
and U8654 (N_8654,N_6064,N_3794);
nand U8655 (N_8655,N_4775,N_3506);
nand U8656 (N_8656,N_5228,N_3575);
nor U8657 (N_8657,N_5667,N_5193);
or U8658 (N_8658,N_4668,N_4201);
xor U8659 (N_8659,N_5485,N_4898);
nor U8660 (N_8660,N_5667,N_4425);
xnor U8661 (N_8661,N_5442,N_5368);
xor U8662 (N_8662,N_4319,N_3802);
xnor U8663 (N_8663,N_3982,N_4577);
nor U8664 (N_8664,N_5961,N_4078);
and U8665 (N_8665,N_6106,N_4609);
or U8666 (N_8666,N_3227,N_4727);
and U8667 (N_8667,N_3171,N_4242);
or U8668 (N_8668,N_5962,N_4579);
and U8669 (N_8669,N_4290,N_5866);
nand U8670 (N_8670,N_4419,N_3548);
nand U8671 (N_8671,N_4794,N_4568);
nor U8672 (N_8672,N_5316,N_3598);
or U8673 (N_8673,N_5349,N_5435);
or U8674 (N_8674,N_3907,N_6219);
nand U8675 (N_8675,N_3992,N_4976);
nor U8676 (N_8676,N_4156,N_3676);
or U8677 (N_8677,N_3980,N_4895);
nand U8678 (N_8678,N_4273,N_6096);
nand U8679 (N_8679,N_3938,N_5776);
nor U8680 (N_8680,N_3244,N_3866);
nand U8681 (N_8681,N_5895,N_4370);
and U8682 (N_8682,N_3993,N_5822);
nor U8683 (N_8683,N_3140,N_5347);
nor U8684 (N_8684,N_3628,N_5331);
and U8685 (N_8685,N_4124,N_3239);
and U8686 (N_8686,N_5259,N_3525);
xnor U8687 (N_8687,N_4348,N_5900);
xor U8688 (N_8688,N_5269,N_3449);
nor U8689 (N_8689,N_6138,N_3918);
xor U8690 (N_8690,N_4144,N_3240);
nor U8691 (N_8691,N_5206,N_5313);
or U8692 (N_8692,N_4520,N_5459);
and U8693 (N_8693,N_4641,N_5021);
and U8694 (N_8694,N_4158,N_5672);
or U8695 (N_8695,N_5616,N_5790);
nor U8696 (N_8696,N_4258,N_4701);
nand U8697 (N_8697,N_5893,N_5094);
nand U8698 (N_8698,N_6221,N_4432);
or U8699 (N_8699,N_4419,N_3593);
nor U8700 (N_8700,N_3887,N_3284);
and U8701 (N_8701,N_4551,N_4719);
nand U8702 (N_8702,N_5242,N_3812);
nand U8703 (N_8703,N_5986,N_4582);
nand U8704 (N_8704,N_4471,N_4933);
nand U8705 (N_8705,N_5058,N_5495);
nand U8706 (N_8706,N_3495,N_5514);
nand U8707 (N_8707,N_4752,N_4557);
nand U8708 (N_8708,N_3271,N_4979);
nor U8709 (N_8709,N_3209,N_4558);
and U8710 (N_8710,N_4649,N_4429);
and U8711 (N_8711,N_6086,N_6026);
and U8712 (N_8712,N_4396,N_4582);
or U8713 (N_8713,N_5510,N_5468);
and U8714 (N_8714,N_4635,N_3831);
or U8715 (N_8715,N_4334,N_5244);
and U8716 (N_8716,N_6134,N_6202);
and U8717 (N_8717,N_4300,N_4265);
and U8718 (N_8718,N_5214,N_4449);
nand U8719 (N_8719,N_3163,N_5469);
or U8720 (N_8720,N_5482,N_4857);
nand U8721 (N_8721,N_5856,N_3813);
xnor U8722 (N_8722,N_4051,N_6177);
xnor U8723 (N_8723,N_3833,N_3600);
xor U8724 (N_8724,N_5901,N_3212);
xor U8725 (N_8725,N_6173,N_5660);
and U8726 (N_8726,N_4039,N_5361);
nand U8727 (N_8727,N_4219,N_3731);
nand U8728 (N_8728,N_5490,N_4803);
nand U8729 (N_8729,N_3390,N_5149);
nor U8730 (N_8730,N_3511,N_4400);
xnor U8731 (N_8731,N_4312,N_3651);
or U8732 (N_8732,N_5369,N_5108);
or U8733 (N_8733,N_5390,N_3614);
nor U8734 (N_8734,N_4594,N_5355);
nand U8735 (N_8735,N_4862,N_4278);
nand U8736 (N_8736,N_5555,N_4275);
or U8737 (N_8737,N_4258,N_5927);
xor U8738 (N_8738,N_3237,N_3529);
nor U8739 (N_8739,N_6054,N_5275);
xnor U8740 (N_8740,N_4286,N_4824);
nor U8741 (N_8741,N_5829,N_3985);
nand U8742 (N_8742,N_3923,N_6195);
and U8743 (N_8743,N_4674,N_5349);
xor U8744 (N_8744,N_3165,N_3694);
nand U8745 (N_8745,N_3140,N_3519);
nor U8746 (N_8746,N_5185,N_4688);
or U8747 (N_8747,N_3346,N_5213);
xor U8748 (N_8748,N_3777,N_3164);
nor U8749 (N_8749,N_4787,N_3137);
nand U8750 (N_8750,N_4940,N_4250);
or U8751 (N_8751,N_4290,N_6192);
nand U8752 (N_8752,N_5722,N_4354);
or U8753 (N_8753,N_4046,N_3375);
or U8754 (N_8754,N_4183,N_5492);
nand U8755 (N_8755,N_4291,N_5498);
nand U8756 (N_8756,N_3411,N_4543);
or U8757 (N_8757,N_4804,N_3911);
and U8758 (N_8758,N_3160,N_5541);
and U8759 (N_8759,N_4397,N_6191);
and U8760 (N_8760,N_4307,N_5000);
nand U8761 (N_8761,N_3974,N_4561);
nor U8762 (N_8762,N_5140,N_4836);
and U8763 (N_8763,N_5949,N_5057);
or U8764 (N_8764,N_4851,N_3169);
or U8765 (N_8765,N_4409,N_5175);
or U8766 (N_8766,N_4933,N_3359);
nor U8767 (N_8767,N_3744,N_3694);
or U8768 (N_8768,N_3243,N_4519);
nand U8769 (N_8769,N_4417,N_3954);
nand U8770 (N_8770,N_3245,N_4705);
and U8771 (N_8771,N_4987,N_5785);
and U8772 (N_8772,N_4518,N_3851);
nand U8773 (N_8773,N_5977,N_3152);
nand U8774 (N_8774,N_3827,N_4702);
nor U8775 (N_8775,N_4725,N_4484);
or U8776 (N_8776,N_6191,N_4319);
nor U8777 (N_8777,N_5625,N_4523);
nor U8778 (N_8778,N_4093,N_4958);
or U8779 (N_8779,N_5995,N_3911);
nor U8780 (N_8780,N_4030,N_5957);
nor U8781 (N_8781,N_5013,N_6125);
or U8782 (N_8782,N_3533,N_4227);
nor U8783 (N_8783,N_4747,N_3446);
nand U8784 (N_8784,N_5384,N_5825);
and U8785 (N_8785,N_4691,N_5705);
nor U8786 (N_8786,N_5691,N_3547);
xor U8787 (N_8787,N_4806,N_3782);
or U8788 (N_8788,N_3785,N_5743);
xnor U8789 (N_8789,N_4690,N_3936);
or U8790 (N_8790,N_5910,N_3286);
nand U8791 (N_8791,N_3250,N_5730);
or U8792 (N_8792,N_3721,N_4627);
or U8793 (N_8793,N_5244,N_4500);
and U8794 (N_8794,N_4017,N_3661);
and U8795 (N_8795,N_5643,N_3147);
nand U8796 (N_8796,N_6004,N_4070);
xor U8797 (N_8797,N_4098,N_4649);
nand U8798 (N_8798,N_4147,N_4301);
and U8799 (N_8799,N_3823,N_4938);
nor U8800 (N_8800,N_3827,N_3850);
nor U8801 (N_8801,N_5785,N_5481);
xnor U8802 (N_8802,N_5467,N_6135);
or U8803 (N_8803,N_5251,N_5381);
or U8804 (N_8804,N_3865,N_5643);
and U8805 (N_8805,N_4081,N_5954);
and U8806 (N_8806,N_3200,N_3652);
and U8807 (N_8807,N_3586,N_5006);
and U8808 (N_8808,N_6068,N_5847);
nor U8809 (N_8809,N_3506,N_3189);
nor U8810 (N_8810,N_3803,N_4620);
nor U8811 (N_8811,N_4491,N_6047);
xor U8812 (N_8812,N_3506,N_4469);
nand U8813 (N_8813,N_5258,N_3862);
and U8814 (N_8814,N_4636,N_5783);
xor U8815 (N_8815,N_4348,N_4714);
nor U8816 (N_8816,N_6141,N_3904);
or U8817 (N_8817,N_5909,N_3671);
nor U8818 (N_8818,N_4887,N_5944);
nand U8819 (N_8819,N_4039,N_5913);
and U8820 (N_8820,N_5291,N_4276);
or U8821 (N_8821,N_5631,N_3944);
nor U8822 (N_8822,N_3225,N_5530);
nand U8823 (N_8823,N_3600,N_5025);
and U8824 (N_8824,N_5497,N_5174);
and U8825 (N_8825,N_3506,N_4352);
or U8826 (N_8826,N_4972,N_3936);
nand U8827 (N_8827,N_4347,N_4170);
nand U8828 (N_8828,N_5598,N_3226);
nand U8829 (N_8829,N_5378,N_5485);
nor U8830 (N_8830,N_4752,N_6186);
nand U8831 (N_8831,N_4608,N_4952);
nor U8832 (N_8832,N_4493,N_5024);
and U8833 (N_8833,N_4147,N_3745);
nand U8834 (N_8834,N_5933,N_5995);
xnor U8835 (N_8835,N_6123,N_5274);
or U8836 (N_8836,N_4813,N_6005);
nand U8837 (N_8837,N_4317,N_4530);
or U8838 (N_8838,N_4102,N_5502);
xor U8839 (N_8839,N_4326,N_3530);
nand U8840 (N_8840,N_4163,N_3879);
nand U8841 (N_8841,N_5252,N_3894);
and U8842 (N_8842,N_3876,N_3575);
and U8843 (N_8843,N_5748,N_3475);
nor U8844 (N_8844,N_5232,N_4975);
nand U8845 (N_8845,N_4587,N_4439);
or U8846 (N_8846,N_3477,N_4939);
or U8847 (N_8847,N_4988,N_5224);
or U8848 (N_8848,N_5905,N_3703);
nor U8849 (N_8849,N_3156,N_5785);
and U8850 (N_8850,N_4296,N_4182);
nor U8851 (N_8851,N_5198,N_6218);
nor U8852 (N_8852,N_6196,N_5892);
nor U8853 (N_8853,N_4470,N_4908);
and U8854 (N_8854,N_6070,N_5034);
or U8855 (N_8855,N_5978,N_4073);
nor U8856 (N_8856,N_4698,N_4089);
or U8857 (N_8857,N_3354,N_5867);
and U8858 (N_8858,N_4582,N_5925);
nor U8859 (N_8859,N_5331,N_4233);
and U8860 (N_8860,N_3602,N_5762);
nor U8861 (N_8861,N_5097,N_3575);
or U8862 (N_8862,N_3228,N_3800);
nand U8863 (N_8863,N_3181,N_4794);
nor U8864 (N_8864,N_3889,N_5519);
nor U8865 (N_8865,N_5489,N_5470);
nor U8866 (N_8866,N_5032,N_5672);
and U8867 (N_8867,N_5028,N_5141);
xor U8868 (N_8868,N_4535,N_4832);
nand U8869 (N_8869,N_5937,N_4532);
and U8870 (N_8870,N_5056,N_5892);
nor U8871 (N_8871,N_4155,N_5691);
xnor U8872 (N_8872,N_4848,N_6085);
xnor U8873 (N_8873,N_4932,N_4536);
nand U8874 (N_8874,N_3334,N_5347);
or U8875 (N_8875,N_4493,N_5756);
xor U8876 (N_8876,N_6067,N_5300);
xnor U8877 (N_8877,N_5943,N_4683);
xor U8878 (N_8878,N_3792,N_3759);
nor U8879 (N_8879,N_6055,N_4034);
and U8880 (N_8880,N_4992,N_6091);
and U8881 (N_8881,N_5714,N_3800);
or U8882 (N_8882,N_5126,N_4762);
or U8883 (N_8883,N_4165,N_5550);
nand U8884 (N_8884,N_4563,N_4895);
nor U8885 (N_8885,N_3307,N_5773);
and U8886 (N_8886,N_5179,N_4921);
and U8887 (N_8887,N_4221,N_5955);
or U8888 (N_8888,N_5326,N_3902);
or U8889 (N_8889,N_6113,N_3620);
or U8890 (N_8890,N_5793,N_5303);
and U8891 (N_8891,N_3524,N_4239);
or U8892 (N_8892,N_3365,N_3177);
nor U8893 (N_8893,N_3528,N_5860);
nor U8894 (N_8894,N_3690,N_3687);
or U8895 (N_8895,N_5819,N_5627);
or U8896 (N_8896,N_3177,N_5640);
nand U8897 (N_8897,N_4318,N_4033);
xnor U8898 (N_8898,N_5444,N_3953);
or U8899 (N_8899,N_4855,N_4038);
or U8900 (N_8900,N_5637,N_5962);
nand U8901 (N_8901,N_4885,N_4058);
and U8902 (N_8902,N_4894,N_6120);
nand U8903 (N_8903,N_4850,N_5827);
and U8904 (N_8904,N_4039,N_3195);
nor U8905 (N_8905,N_4489,N_5279);
or U8906 (N_8906,N_5660,N_3304);
nand U8907 (N_8907,N_5424,N_4689);
nor U8908 (N_8908,N_5723,N_6071);
or U8909 (N_8909,N_4026,N_4491);
and U8910 (N_8910,N_3855,N_5741);
or U8911 (N_8911,N_6118,N_3559);
xnor U8912 (N_8912,N_4410,N_4621);
nand U8913 (N_8913,N_4874,N_4477);
or U8914 (N_8914,N_6195,N_5440);
or U8915 (N_8915,N_5987,N_5048);
and U8916 (N_8916,N_5460,N_3938);
or U8917 (N_8917,N_5412,N_6002);
nor U8918 (N_8918,N_4952,N_4353);
nand U8919 (N_8919,N_5974,N_5164);
and U8920 (N_8920,N_4080,N_4664);
nor U8921 (N_8921,N_5416,N_3127);
nand U8922 (N_8922,N_6141,N_5053);
xnor U8923 (N_8923,N_4380,N_4917);
or U8924 (N_8924,N_6056,N_4350);
and U8925 (N_8925,N_5564,N_5418);
xor U8926 (N_8926,N_5942,N_6105);
nor U8927 (N_8927,N_5598,N_3961);
and U8928 (N_8928,N_5267,N_4235);
nand U8929 (N_8929,N_6141,N_5914);
and U8930 (N_8930,N_3590,N_5958);
and U8931 (N_8931,N_4564,N_5000);
nor U8932 (N_8932,N_4625,N_4071);
nor U8933 (N_8933,N_3876,N_3701);
or U8934 (N_8934,N_3783,N_4487);
and U8935 (N_8935,N_3928,N_3724);
nand U8936 (N_8936,N_4095,N_5431);
nor U8937 (N_8937,N_3763,N_3268);
nand U8938 (N_8938,N_4303,N_5547);
nor U8939 (N_8939,N_5980,N_3628);
nor U8940 (N_8940,N_5509,N_3476);
nand U8941 (N_8941,N_3835,N_6242);
or U8942 (N_8942,N_5804,N_4174);
nand U8943 (N_8943,N_3935,N_3171);
and U8944 (N_8944,N_4393,N_5662);
xor U8945 (N_8945,N_3426,N_5200);
xor U8946 (N_8946,N_4836,N_5908);
xnor U8947 (N_8947,N_3992,N_3161);
and U8948 (N_8948,N_5135,N_5807);
xor U8949 (N_8949,N_4880,N_4533);
and U8950 (N_8950,N_3827,N_5757);
nor U8951 (N_8951,N_5681,N_6012);
nand U8952 (N_8952,N_4554,N_3330);
nor U8953 (N_8953,N_6063,N_4671);
and U8954 (N_8954,N_3897,N_5638);
nor U8955 (N_8955,N_4829,N_3628);
nand U8956 (N_8956,N_5841,N_3286);
nand U8957 (N_8957,N_4323,N_3773);
or U8958 (N_8958,N_5093,N_3395);
or U8959 (N_8959,N_3739,N_3646);
or U8960 (N_8960,N_3271,N_5832);
nor U8961 (N_8961,N_3568,N_3554);
nor U8962 (N_8962,N_5051,N_4100);
nand U8963 (N_8963,N_5110,N_4265);
nand U8964 (N_8964,N_3174,N_4945);
and U8965 (N_8965,N_5863,N_5190);
or U8966 (N_8966,N_3357,N_6244);
and U8967 (N_8967,N_4776,N_6206);
and U8968 (N_8968,N_4373,N_6161);
nand U8969 (N_8969,N_3151,N_4696);
nor U8970 (N_8970,N_4005,N_4768);
xnor U8971 (N_8971,N_3142,N_4343);
nor U8972 (N_8972,N_3285,N_4754);
and U8973 (N_8973,N_4819,N_5689);
nand U8974 (N_8974,N_3209,N_3788);
nor U8975 (N_8975,N_3233,N_5542);
nor U8976 (N_8976,N_5349,N_3164);
or U8977 (N_8977,N_6159,N_3350);
or U8978 (N_8978,N_3845,N_3800);
nor U8979 (N_8979,N_3258,N_6229);
and U8980 (N_8980,N_5459,N_6032);
or U8981 (N_8981,N_5957,N_3372);
nor U8982 (N_8982,N_4279,N_5507);
or U8983 (N_8983,N_4817,N_3336);
or U8984 (N_8984,N_5799,N_4162);
and U8985 (N_8985,N_4835,N_4887);
and U8986 (N_8986,N_3573,N_3287);
nand U8987 (N_8987,N_5802,N_5990);
nor U8988 (N_8988,N_4289,N_3898);
and U8989 (N_8989,N_4835,N_4647);
xnor U8990 (N_8990,N_3328,N_3425);
xor U8991 (N_8991,N_4818,N_5149);
and U8992 (N_8992,N_5667,N_5662);
nor U8993 (N_8993,N_4385,N_4405);
or U8994 (N_8994,N_3985,N_5192);
and U8995 (N_8995,N_6146,N_3255);
nand U8996 (N_8996,N_5061,N_4744);
nand U8997 (N_8997,N_3731,N_4019);
xnor U8998 (N_8998,N_4225,N_5255);
and U8999 (N_8999,N_4690,N_5609);
or U9000 (N_9000,N_3852,N_5745);
or U9001 (N_9001,N_3617,N_5992);
nor U9002 (N_9002,N_5965,N_5918);
nand U9003 (N_9003,N_4628,N_3447);
or U9004 (N_9004,N_3945,N_5201);
and U9005 (N_9005,N_3972,N_4201);
and U9006 (N_9006,N_3836,N_3760);
nor U9007 (N_9007,N_5881,N_5609);
and U9008 (N_9008,N_3854,N_4641);
or U9009 (N_9009,N_4211,N_4405);
nand U9010 (N_9010,N_5621,N_5462);
or U9011 (N_9011,N_4953,N_4188);
nand U9012 (N_9012,N_5837,N_5186);
nand U9013 (N_9013,N_4682,N_5270);
and U9014 (N_9014,N_4525,N_6175);
nand U9015 (N_9015,N_3877,N_3761);
or U9016 (N_9016,N_4767,N_4736);
or U9017 (N_9017,N_5606,N_3219);
or U9018 (N_9018,N_3598,N_3724);
and U9019 (N_9019,N_5447,N_4201);
nand U9020 (N_9020,N_5503,N_4961);
or U9021 (N_9021,N_6218,N_5239);
and U9022 (N_9022,N_4484,N_3669);
and U9023 (N_9023,N_5052,N_5423);
and U9024 (N_9024,N_5416,N_3879);
nand U9025 (N_9025,N_5825,N_3244);
xnor U9026 (N_9026,N_5592,N_5427);
or U9027 (N_9027,N_5504,N_5702);
xnor U9028 (N_9028,N_5282,N_5152);
or U9029 (N_9029,N_3181,N_5505);
nor U9030 (N_9030,N_5597,N_4387);
or U9031 (N_9031,N_6144,N_5761);
nand U9032 (N_9032,N_3704,N_3739);
and U9033 (N_9033,N_3918,N_5197);
xnor U9034 (N_9034,N_3485,N_4746);
or U9035 (N_9035,N_6114,N_3183);
xnor U9036 (N_9036,N_6164,N_5921);
nand U9037 (N_9037,N_4367,N_3966);
nand U9038 (N_9038,N_3702,N_6080);
xnor U9039 (N_9039,N_5790,N_5431);
and U9040 (N_9040,N_6143,N_5927);
nand U9041 (N_9041,N_5843,N_4969);
or U9042 (N_9042,N_3655,N_5986);
or U9043 (N_9043,N_4707,N_6035);
nor U9044 (N_9044,N_5200,N_3356);
xnor U9045 (N_9045,N_4964,N_4987);
or U9046 (N_9046,N_3568,N_3603);
nor U9047 (N_9047,N_5293,N_3404);
or U9048 (N_9048,N_5757,N_3385);
nand U9049 (N_9049,N_5523,N_5955);
nand U9050 (N_9050,N_3824,N_3628);
and U9051 (N_9051,N_5593,N_5112);
nor U9052 (N_9052,N_5040,N_5850);
nand U9053 (N_9053,N_5189,N_4052);
or U9054 (N_9054,N_4769,N_3233);
and U9055 (N_9055,N_6152,N_5063);
or U9056 (N_9056,N_3849,N_5200);
and U9057 (N_9057,N_4517,N_3633);
nor U9058 (N_9058,N_4061,N_5985);
nand U9059 (N_9059,N_5660,N_4231);
xnor U9060 (N_9060,N_4144,N_3648);
nor U9061 (N_9061,N_4533,N_4196);
and U9062 (N_9062,N_4819,N_3269);
and U9063 (N_9063,N_4245,N_4606);
and U9064 (N_9064,N_5598,N_3274);
or U9065 (N_9065,N_5475,N_5419);
or U9066 (N_9066,N_5161,N_5650);
or U9067 (N_9067,N_4376,N_5732);
or U9068 (N_9068,N_5351,N_4586);
nor U9069 (N_9069,N_5299,N_5788);
xor U9070 (N_9070,N_4484,N_4908);
or U9071 (N_9071,N_4423,N_3617);
and U9072 (N_9072,N_4181,N_6025);
or U9073 (N_9073,N_3870,N_6053);
xor U9074 (N_9074,N_3666,N_5012);
or U9075 (N_9075,N_3803,N_5046);
xnor U9076 (N_9076,N_5382,N_6192);
xor U9077 (N_9077,N_4143,N_3919);
or U9078 (N_9078,N_4150,N_4828);
or U9079 (N_9079,N_3570,N_3360);
nor U9080 (N_9080,N_4171,N_3422);
nor U9081 (N_9081,N_5207,N_5157);
nand U9082 (N_9082,N_4929,N_3226);
nor U9083 (N_9083,N_5852,N_3415);
nand U9084 (N_9084,N_3490,N_5841);
or U9085 (N_9085,N_3923,N_3786);
and U9086 (N_9086,N_4684,N_4472);
nand U9087 (N_9087,N_4302,N_4025);
nor U9088 (N_9088,N_5098,N_3957);
or U9089 (N_9089,N_5047,N_5198);
or U9090 (N_9090,N_3822,N_6149);
nor U9091 (N_9091,N_4102,N_3993);
xnor U9092 (N_9092,N_4610,N_4410);
nor U9093 (N_9093,N_5550,N_3976);
or U9094 (N_9094,N_5022,N_3755);
or U9095 (N_9095,N_5263,N_3154);
nand U9096 (N_9096,N_4308,N_6034);
and U9097 (N_9097,N_4832,N_3649);
nand U9098 (N_9098,N_5647,N_6063);
nor U9099 (N_9099,N_3792,N_4718);
nand U9100 (N_9100,N_5789,N_4395);
nand U9101 (N_9101,N_3578,N_4625);
or U9102 (N_9102,N_3417,N_6007);
and U9103 (N_9103,N_5513,N_4284);
or U9104 (N_9104,N_4625,N_5512);
and U9105 (N_9105,N_3437,N_4235);
nor U9106 (N_9106,N_4505,N_4673);
nand U9107 (N_9107,N_5208,N_5012);
nor U9108 (N_9108,N_3511,N_4052);
nand U9109 (N_9109,N_6096,N_5086);
or U9110 (N_9110,N_5918,N_5951);
xnor U9111 (N_9111,N_4945,N_3198);
nor U9112 (N_9112,N_3804,N_4159);
nand U9113 (N_9113,N_5625,N_4697);
and U9114 (N_9114,N_3967,N_5547);
or U9115 (N_9115,N_3700,N_3226);
and U9116 (N_9116,N_3871,N_3799);
and U9117 (N_9117,N_5576,N_3715);
nand U9118 (N_9118,N_6089,N_5282);
and U9119 (N_9119,N_3227,N_5354);
nand U9120 (N_9120,N_6211,N_4625);
nor U9121 (N_9121,N_6039,N_5735);
or U9122 (N_9122,N_4344,N_3921);
nand U9123 (N_9123,N_5049,N_4398);
nor U9124 (N_9124,N_5268,N_5483);
and U9125 (N_9125,N_5544,N_3774);
and U9126 (N_9126,N_3966,N_4613);
nor U9127 (N_9127,N_5179,N_5937);
nand U9128 (N_9128,N_3943,N_3342);
xor U9129 (N_9129,N_4860,N_5209);
nand U9130 (N_9130,N_4551,N_6124);
nor U9131 (N_9131,N_4874,N_3663);
or U9132 (N_9132,N_4329,N_5321);
and U9133 (N_9133,N_4565,N_3919);
xor U9134 (N_9134,N_4943,N_5175);
nor U9135 (N_9135,N_5390,N_5510);
nor U9136 (N_9136,N_4096,N_3482);
nor U9137 (N_9137,N_4229,N_5310);
or U9138 (N_9138,N_4628,N_5694);
or U9139 (N_9139,N_5986,N_5985);
or U9140 (N_9140,N_3188,N_4010);
and U9141 (N_9141,N_4393,N_5062);
and U9142 (N_9142,N_5702,N_4620);
or U9143 (N_9143,N_3216,N_4343);
nand U9144 (N_9144,N_4303,N_4423);
and U9145 (N_9145,N_5917,N_5570);
nor U9146 (N_9146,N_3554,N_5038);
nand U9147 (N_9147,N_5089,N_5780);
and U9148 (N_9148,N_3377,N_4493);
or U9149 (N_9149,N_3461,N_4414);
and U9150 (N_9150,N_5562,N_4917);
nand U9151 (N_9151,N_5835,N_5684);
or U9152 (N_9152,N_5236,N_4911);
nand U9153 (N_9153,N_5555,N_3465);
nand U9154 (N_9154,N_6211,N_6197);
and U9155 (N_9155,N_5479,N_5119);
nor U9156 (N_9156,N_6231,N_4129);
and U9157 (N_9157,N_3156,N_3518);
or U9158 (N_9158,N_5803,N_3412);
or U9159 (N_9159,N_5212,N_4515);
and U9160 (N_9160,N_3158,N_4415);
or U9161 (N_9161,N_4505,N_4527);
or U9162 (N_9162,N_3150,N_4446);
nor U9163 (N_9163,N_5921,N_5535);
or U9164 (N_9164,N_5516,N_5867);
or U9165 (N_9165,N_5638,N_4772);
nand U9166 (N_9166,N_3671,N_4210);
and U9167 (N_9167,N_5565,N_3718);
xnor U9168 (N_9168,N_3702,N_5617);
xor U9169 (N_9169,N_5124,N_4410);
and U9170 (N_9170,N_5332,N_3698);
nand U9171 (N_9171,N_4099,N_4592);
or U9172 (N_9172,N_5371,N_4279);
nand U9173 (N_9173,N_3763,N_5881);
nand U9174 (N_9174,N_4855,N_5910);
or U9175 (N_9175,N_3313,N_3554);
nand U9176 (N_9176,N_4172,N_4013);
nand U9177 (N_9177,N_5168,N_5995);
and U9178 (N_9178,N_6228,N_4603);
nand U9179 (N_9179,N_4157,N_4851);
and U9180 (N_9180,N_5572,N_4053);
nor U9181 (N_9181,N_3278,N_3322);
or U9182 (N_9182,N_4656,N_3958);
and U9183 (N_9183,N_5233,N_4741);
nand U9184 (N_9184,N_4632,N_5171);
and U9185 (N_9185,N_5367,N_3901);
nor U9186 (N_9186,N_5033,N_6029);
nand U9187 (N_9187,N_4778,N_3948);
or U9188 (N_9188,N_3464,N_3811);
nor U9189 (N_9189,N_5452,N_4472);
and U9190 (N_9190,N_5064,N_5345);
or U9191 (N_9191,N_3697,N_3261);
nand U9192 (N_9192,N_4772,N_3416);
nand U9193 (N_9193,N_4999,N_5007);
and U9194 (N_9194,N_4798,N_5824);
and U9195 (N_9195,N_3372,N_3144);
nand U9196 (N_9196,N_3790,N_4151);
or U9197 (N_9197,N_4055,N_5527);
nor U9198 (N_9198,N_4486,N_3775);
nor U9199 (N_9199,N_3613,N_3917);
nand U9200 (N_9200,N_3901,N_4321);
and U9201 (N_9201,N_4547,N_5136);
nor U9202 (N_9202,N_3426,N_5225);
nor U9203 (N_9203,N_3621,N_4433);
and U9204 (N_9204,N_3195,N_3249);
or U9205 (N_9205,N_4822,N_5647);
nand U9206 (N_9206,N_3776,N_4184);
nor U9207 (N_9207,N_3173,N_5625);
or U9208 (N_9208,N_5535,N_5951);
and U9209 (N_9209,N_4537,N_4272);
nand U9210 (N_9210,N_6160,N_4020);
and U9211 (N_9211,N_3129,N_6133);
xor U9212 (N_9212,N_5820,N_3795);
and U9213 (N_9213,N_3390,N_3932);
nor U9214 (N_9214,N_4484,N_5365);
nand U9215 (N_9215,N_4900,N_3590);
and U9216 (N_9216,N_4661,N_4899);
and U9217 (N_9217,N_4565,N_5187);
xnor U9218 (N_9218,N_4211,N_5917);
nand U9219 (N_9219,N_5525,N_3799);
or U9220 (N_9220,N_4718,N_4927);
and U9221 (N_9221,N_5826,N_4476);
and U9222 (N_9222,N_3541,N_6007);
and U9223 (N_9223,N_5363,N_5375);
nor U9224 (N_9224,N_6200,N_3849);
xor U9225 (N_9225,N_4494,N_3503);
and U9226 (N_9226,N_3919,N_5488);
or U9227 (N_9227,N_5189,N_3216);
xnor U9228 (N_9228,N_4111,N_4404);
nor U9229 (N_9229,N_5329,N_3825);
or U9230 (N_9230,N_3932,N_5126);
nand U9231 (N_9231,N_6086,N_6121);
nand U9232 (N_9232,N_5895,N_4097);
or U9233 (N_9233,N_4408,N_6023);
nand U9234 (N_9234,N_5144,N_4675);
and U9235 (N_9235,N_4027,N_3708);
and U9236 (N_9236,N_6204,N_5340);
nor U9237 (N_9237,N_6025,N_3182);
nand U9238 (N_9238,N_5499,N_3768);
nor U9239 (N_9239,N_4070,N_5848);
and U9240 (N_9240,N_6249,N_4950);
nand U9241 (N_9241,N_3780,N_3299);
nor U9242 (N_9242,N_4918,N_3200);
nor U9243 (N_9243,N_5488,N_5834);
nor U9244 (N_9244,N_5891,N_5176);
and U9245 (N_9245,N_6082,N_6137);
and U9246 (N_9246,N_4611,N_5184);
and U9247 (N_9247,N_3812,N_5371);
nor U9248 (N_9248,N_5152,N_5507);
nor U9249 (N_9249,N_4939,N_4197);
xor U9250 (N_9250,N_4440,N_3769);
nor U9251 (N_9251,N_4810,N_3603);
nand U9252 (N_9252,N_4207,N_3137);
and U9253 (N_9253,N_5419,N_5025);
or U9254 (N_9254,N_4310,N_4242);
nand U9255 (N_9255,N_3620,N_3693);
xor U9256 (N_9256,N_3200,N_4764);
and U9257 (N_9257,N_6160,N_4070);
nand U9258 (N_9258,N_5618,N_4111);
nor U9259 (N_9259,N_5490,N_4202);
nor U9260 (N_9260,N_5621,N_3604);
xnor U9261 (N_9261,N_5657,N_5043);
or U9262 (N_9262,N_3294,N_5505);
nor U9263 (N_9263,N_4024,N_5799);
and U9264 (N_9264,N_3254,N_4090);
or U9265 (N_9265,N_4710,N_4000);
nor U9266 (N_9266,N_5738,N_3575);
nand U9267 (N_9267,N_4287,N_3610);
and U9268 (N_9268,N_3686,N_3429);
nor U9269 (N_9269,N_3665,N_5085);
or U9270 (N_9270,N_3300,N_6076);
xor U9271 (N_9271,N_5877,N_4116);
xor U9272 (N_9272,N_5224,N_3290);
nand U9273 (N_9273,N_5756,N_3455);
nor U9274 (N_9274,N_3257,N_4888);
nand U9275 (N_9275,N_4759,N_4645);
and U9276 (N_9276,N_6202,N_3570);
and U9277 (N_9277,N_6025,N_5825);
nor U9278 (N_9278,N_3435,N_4155);
or U9279 (N_9279,N_5410,N_5404);
nor U9280 (N_9280,N_4725,N_3695);
nor U9281 (N_9281,N_4144,N_4421);
nand U9282 (N_9282,N_5931,N_3592);
or U9283 (N_9283,N_5799,N_5406);
nor U9284 (N_9284,N_5641,N_4436);
or U9285 (N_9285,N_5435,N_6030);
or U9286 (N_9286,N_4627,N_4274);
nor U9287 (N_9287,N_5157,N_3697);
nand U9288 (N_9288,N_5802,N_3433);
or U9289 (N_9289,N_6131,N_5643);
nand U9290 (N_9290,N_5739,N_6036);
and U9291 (N_9291,N_4237,N_5761);
nor U9292 (N_9292,N_3185,N_4961);
or U9293 (N_9293,N_6161,N_5092);
or U9294 (N_9294,N_5608,N_4442);
or U9295 (N_9295,N_4665,N_3799);
xor U9296 (N_9296,N_3786,N_4654);
or U9297 (N_9297,N_4754,N_5773);
or U9298 (N_9298,N_5783,N_3728);
nor U9299 (N_9299,N_4357,N_4472);
nor U9300 (N_9300,N_5509,N_5589);
nor U9301 (N_9301,N_3505,N_5921);
nand U9302 (N_9302,N_5019,N_3390);
and U9303 (N_9303,N_4868,N_4309);
nand U9304 (N_9304,N_3185,N_4753);
and U9305 (N_9305,N_6023,N_3681);
or U9306 (N_9306,N_4533,N_5145);
nor U9307 (N_9307,N_6168,N_4423);
and U9308 (N_9308,N_4799,N_5705);
nand U9309 (N_9309,N_6053,N_5164);
or U9310 (N_9310,N_3501,N_6218);
nand U9311 (N_9311,N_3820,N_3530);
xor U9312 (N_9312,N_5999,N_3882);
or U9313 (N_9313,N_5192,N_4601);
nor U9314 (N_9314,N_3398,N_3504);
and U9315 (N_9315,N_3492,N_3409);
or U9316 (N_9316,N_5009,N_4537);
or U9317 (N_9317,N_3324,N_4505);
and U9318 (N_9318,N_5523,N_3684);
and U9319 (N_9319,N_3427,N_5047);
nor U9320 (N_9320,N_5914,N_5428);
nand U9321 (N_9321,N_3592,N_3518);
nor U9322 (N_9322,N_5866,N_5906);
nand U9323 (N_9323,N_3825,N_5571);
or U9324 (N_9324,N_3363,N_5349);
or U9325 (N_9325,N_3401,N_4740);
and U9326 (N_9326,N_5635,N_3173);
nor U9327 (N_9327,N_4278,N_5983);
and U9328 (N_9328,N_4886,N_4481);
xnor U9329 (N_9329,N_5148,N_5601);
xor U9330 (N_9330,N_4097,N_5713);
nand U9331 (N_9331,N_5481,N_5747);
nor U9332 (N_9332,N_5917,N_5048);
nor U9333 (N_9333,N_4006,N_4289);
nand U9334 (N_9334,N_4640,N_4995);
or U9335 (N_9335,N_5242,N_4460);
nand U9336 (N_9336,N_5147,N_5661);
nor U9337 (N_9337,N_5187,N_4661);
and U9338 (N_9338,N_3344,N_5538);
or U9339 (N_9339,N_5401,N_6237);
nor U9340 (N_9340,N_5384,N_4766);
nor U9341 (N_9341,N_3172,N_5288);
nand U9342 (N_9342,N_4678,N_4584);
and U9343 (N_9343,N_3180,N_3925);
nand U9344 (N_9344,N_3477,N_4614);
or U9345 (N_9345,N_6228,N_4775);
or U9346 (N_9346,N_5898,N_6095);
and U9347 (N_9347,N_5190,N_5165);
nor U9348 (N_9348,N_4170,N_3867);
xnor U9349 (N_9349,N_4423,N_3248);
nand U9350 (N_9350,N_4118,N_5654);
nand U9351 (N_9351,N_5925,N_4150);
and U9352 (N_9352,N_4279,N_5585);
or U9353 (N_9353,N_4811,N_5059);
and U9354 (N_9354,N_3644,N_4605);
and U9355 (N_9355,N_4141,N_3189);
xnor U9356 (N_9356,N_5310,N_3496);
xnor U9357 (N_9357,N_5779,N_5411);
nand U9358 (N_9358,N_4444,N_5770);
nor U9359 (N_9359,N_4699,N_4999);
or U9360 (N_9360,N_3778,N_3937);
nand U9361 (N_9361,N_5068,N_3730);
and U9362 (N_9362,N_3229,N_5204);
nand U9363 (N_9363,N_6173,N_3574);
xor U9364 (N_9364,N_5532,N_3259);
and U9365 (N_9365,N_3358,N_5218);
nand U9366 (N_9366,N_4950,N_5494);
and U9367 (N_9367,N_3975,N_5396);
nor U9368 (N_9368,N_5984,N_3584);
xor U9369 (N_9369,N_3207,N_5383);
or U9370 (N_9370,N_4686,N_4257);
or U9371 (N_9371,N_3446,N_4246);
nand U9372 (N_9372,N_4269,N_5851);
nor U9373 (N_9373,N_4119,N_4425);
or U9374 (N_9374,N_4182,N_4228);
nor U9375 (N_9375,N_8860,N_7114);
or U9376 (N_9376,N_8298,N_8516);
and U9377 (N_9377,N_7898,N_7514);
nand U9378 (N_9378,N_6444,N_7750);
nor U9379 (N_9379,N_6305,N_7987);
nand U9380 (N_9380,N_8544,N_8972);
nor U9381 (N_9381,N_9104,N_6303);
nor U9382 (N_9382,N_8553,N_8607);
and U9383 (N_9383,N_7092,N_6621);
xor U9384 (N_9384,N_8128,N_7058);
nor U9385 (N_9385,N_9274,N_6952);
and U9386 (N_9386,N_7233,N_7256);
nor U9387 (N_9387,N_7464,N_8865);
or U9388 (N_9388,N_6709,N_6357);
nor U9389 (N_9389,N_8229,N_8275);
xor U9390 (N_9390,N_7866,N_9123);
and U9391 (N_9391,N_8041,N_8347);
xnor U9392 (N_9392,N_8631,N_7002);
or U9393 (N_9393,N_9210,N_9325);
and U9394 (N_9394,N_7166,N_9354);
or U9395 (N_9395,N_6359,N_8751);
and U9396 (N_9396,N_6437,N_8778);
nand U9397 (N_9397,N_6711,N_7201);
or U9398 (N_9398,N_6984,N_7271);
and U9399 (N_9399,N_6351,N_8098);
or U9400 (N_9400,N_7786,N_8345);
nand U9401 (N_9401,N_6646,N_8620);
nand U9402 (N_9402,N_6917,N_6833);
or U9403 (N_9403,N_8710,N_8821);
nand U9404 (N_9404,N_6591,N_6710);
nor U9405 (N_9405,N_8195,N_8102);
or U9406 (N_9406,N_9027,N_6254);
or U9407 (N_9407,N_7616,N_6502);
nor U9408 (N_9408,N_6265,N_8331);
and U9409 (N_9409,N_7422,N_8154);
and U9410 (N_9410,N_6471,N_8076);
or U9411 (N_9411,N_7590,N_7810);
nand U9412 (N_9412,N_7081,N_7352);
and U9413 (N_9413,N_6697,N_9072);
xnor U9414 (N_9414,N_8449,N_6275);
and U9415 (N_9415,N_7158,N_6630);
nand U9416 (N_9416,N_7951,N_9288);
nand U9417 (N_9417,N_9300,N_9146);
and U9418 (N_9418,N_7922,N_7751);
xor U9419 (N_9419,N_8312,N_6823);
or U9420 (N_9420,N_7797,N_7875);
and U9421 (N_9421,N_8953,N_8501);
nand U9422 (N_9422,N_8922,N_6671);
or U9423 (N_9423,N_7394,N_6329);
nor U9424 (N_9424,N_6512,N_8100);
or U9425 (N_9425,N_8358,N_8720);
and U9426 (N_9426,N_8882,N_7443);
and U9427 (N_9427,N_7530,N_6935);
nor U9428 (N_9428,N_8061,N_7504);
and U9429 (N_9429,N_7222,N_8563);
or U9430 (N_9430,N_8589,N_6448);
or U9431 (N_9431,N_9307,N_7802);
nand U9432 (N_9432,N_8227,N_7149);
nor U9433 (N_9433,N_9235,N_9362);
and U9434 (N_9434,N_9247,N_8459);
or U9435 (N_9435,N_7791,N_7240);
nor U9436 (N_9436,N_8392,N_7568);
or U9437 (N_9437,N_6724,N_7363);
nor U9438 (N_9438,N_8899,N_9172);
or U9439 (N_9439,N_6676,N_8914);
or U9440 (N_9440,N_9074,N_6566);
nor U9441 (N_9441,N_8852,N_7093);
nor U9442 (N_9442,N_8595,N_7237);
nor U9443 (N_9443,N_7812,N_8156);
or U9444 (N_9444,N_7206,N_7047);
and U9445 (N_9445,N_7565,N_8601);
and U9446 (N_9446,N_8220,N_8605);
nand U9447 (N_9447,N_9233,N_6844);
and U9448 (N_9448,N_6576,N_8513);
and U9449 (N_9449,N_8107,N_7526);
nand U9450 (N_9450,N_7887,N_9046);
nand U9451 (N_9451,N_7692,N_8646);
nor U9452 (N_9452,N_7708,N_6445);
and U9453 (N_9453,N_9187,N_8293);
and U9454 (N_9454,N_8350,N_7929);
or U9455 (N_9455,N_6947,N_6936);
and U9456 (N_9456,N_9251,N_7752);
nor U9457 (N_9457,N_9149,N_8702);
and U9458 (N_9458,N_6853,N_8583);
and U9459 (N_9459,N_7417,N_8269);
nor U9460 (N_9460,N_8713,N_8341);
or U9461 (N_9461,N_7931,N_7889);
nor U9462 (N_9462,N_6633,N_8127);
and U9463 (N_9463,N_7524,N_9353);
and U9464 (N_9464,N_8448,N_6541);
or U9465 (N_9465,N_7978,N_8876);
nand U9466 (N_9466,N_6775,N_8669);
nand U9467 (N_9467,N_9335,N_7562);
and U9468 (N_9468,N_6883,N_6687);
and U9469 (N_9469,N_9250,N_7971);
and U9470 (N_9470,N_8433,N_8185);
nand U9471 (N_9471,N_7336,N_7434);
xnor U9472 (N_9472,N_7532,N_6438);
and U9473 (N_9473,N_6705,N_8259);
nand U9474 (N_9474,N_8169,N_7442);
and U9475 (N_9475,N_8733,N_8321);
nand U9476 (N_9476,N_8307,N_6930);
nand U9477 (N_9477,N_8840,N_8153);
or U9478 (N_9478,N_7566,N_6718);
or U9479 (N_9479,N_8579,N_7415);
xor U9480 (N_9480,N_7426,N_8097);
xor U9481 (N_9481,N_8013,N_6252);
or U9482 (N_9482,N_8581,N_8388);
or U9483 (N_9483,N_8394,N_8330);
nand U9484 (N_9484,N_6458,N_8164);
and U9485 (N_9485,N_6260,N_8479);
nor U9486 (N_9486,N_6764,N_8763);
or U9487 (N_9487,N_7662,N_7075);
xnor U9488 (N_9488,N_9010,N_9317);
nor U9489 (N_9489,N_7247,N_6565);
and U9490 (N_9490,N_9209,N_9183);
and U9491 (N_9491,N_7461,N_9238);
nor U9492 (N_9492,N_7681,N_9135);
nor U9493 (N_9493,N_8343,N_8382);
nand U9494 (N_9494,N_6339,N_8724);
nand U9495 (N_9495,N_6267,N_6350);
nor U9496 (N_9496,N_8706,N_7414);
and U9497 (N_9497,N_9330,N_7212);
and U9498 (N_9498,N_6452,N_6500);
nor U9499 (N_9499,N_7881,N_8356);
nor U9500 (N_9500,N_6868,N_8971);
and U9501 (N_9501,N_6542,N_8215);
and U9502 (N_9502,N_7132,N_7517);
nor U9503 (N_9503,N_6349,N_6663);
nand U9504 (N_9504,N_6561,N_6478);
nor U9505 (N_9505,N_9269,N_6372);
nand U9506 (N_9506,N_6376,N_6672);
or U9507 (N_9507,N_7963,N_8122);
nand U9508 (N_9508,N_8494,N_6348);
or U9509 (N_9509,N_7079,N_6944);
or U9510 (N_9510,N_6825,N_8217);
nor U9511 (N_9511,N_8611,N_8892);
or U9512 (N_9512,N_8768,N_8189);
nand U9513 (N_9513,N_7339,N_8874);
or U9514 (N_9514,N_6501,N_8214);
nor U9515 (N_9515,N_7762,N_8488);
nand U9516 (N_9516,N_7354,N_9013);
nor U9517 (N_9517,N_7159,N_8858);
and U9518 (N_9518,N_8912,N_6874);
and U9519 (N_9519,N_7445,N_7539);
nor U9520 (N_9520,N_7669,N_7969);
nor U9521 (N_9521,N_6666,N_9161);
or U9522 (N_9522,N_8963,N_8253);
or U9523 (N_9523,N_7962,N_8309);
nand U9524 (N_9524,N_7968,N_6963);
xnor U9525 (N_9525,N_8979,N_8788);
nor U9526 (N_9526,N_8523,N_7450);
nor U9527 (N_9527,N_7956,N_7747);
nor U9528 (N_9528,N_8032,N_7757);
nand U9529 (N_9529,N_8784,N_8905);
and U9530 (N_9530,N_8091,N_9184);
xnor U9531 (N_9531,N_9345,N_9266);
xnor U9532 (N_9532,N_9014,N_6774);
or U9533 (N_9533,N_7936,N_6263);
nand U9534 (N_9534,N_7519,N_6923);
nor U9535 (N_9535,N_7553,N_8042);
or U9536 (N_9536,N_8604,N_6755);
xor U9537 (N_9537,N_8813,N_6848);
nand U9538 (N_9538,N_6993,N_9240);
xnor U9539 (N_9539,N_8211,N_7537);
and U9540 (N_9540,N_8552,N_7481);
nor U9541 (N_9541,N_8365,N_8994);
or U9542 (N_9542,N_8908,N_6530);
nor U9543 (N_9543,N_8691,N_6706);
or U9544 (N_9544,N_6946,N_6776);
nor U9545 (N_9545,N_8430,N_7477);
or U9546 (N_9546,N_7003,N_7295);
and U9547 (N_9547,N_7226,N_6827);
nor U9548 (N_9548,N_6735,N_9285);
xnor U9549 (N_9549,N_9218,N_6943);
or U9550 (N_9550,N_7389,N_8477);
nand U9551 (N_9551,N_7470,N_8791);
or U9552 (N_9552,N_7953,N_8888);
and U9553 (N_9553,N_8960,N_7794);
xnor U9554 (N_9554,N_6434,N_7637);
nor U9555 (N_9555,N_6745,N_8342);
nor U9556 (N_9556,N_9009,N_7246);
or U9557 (N_9557,N_9136,N_7959);
nand U9558 (N_9558,N_8149,N_7941);
or U9559 (N_9559,N_6343,N_6538);
nor U9560 (N_9560,N_9153,N_7948);
xnor U9561 (N_9561,N_6955,N_7588);
or U9562 (N_9562,N_6696,N_7419);
nor U9563 (N_9563,N_7650,N_6781);
and U9564 (N_9564,N_8773,N_6713);
nand U9565 (N_9565,N_7239,N_7264);
nand U9566 (N_9566,N_7975,N_8679);
nor U9567 (N_9567,N_8825,N_7670);
or U9568 (N_9568,N_7925,N_7111);
nand U9569 (N_9569,N_9331,N_8173);
xor U9570 (N_9570,N_6763,N_7583);
xnor U9571 (N_9571,N_6345,N_7998);
nor U9572 (N_9572,N_8664,N_9348);
nor U9573 (N_9573,N_7703,N_7260);
nor U9574 (N_9574,N_8588,N_8411);
and U9575 (N_9575,N_8105,N_7973);
nor U9576 (N_9576,N_6392,N_7143);
nor U9577 (N_9577,N_9308,N_8661);
nor U9578 (N_9578,N_7314,N_7014);
nand U9579 (N_9579,N_8935,N_6995);
and U9580 (N_9580,N_7800,N_9350);
or U9581 (N_9581,N_8842,N_6627);
or U9582 (N_9582,N_9359,N_7454);
and U9583 (N_9583,N_6894,N_9207);
nand U9584 (N_9584,N_7917,N_7360);
nor U9585 (N_9585,N_8171,N_6669);
and U9586 (N_9586,N_6980,N_7387);
nor U9587 (N_9587,N_8961,N_8817);
nand U9588 (N_9588,N_8668,N_6596);
nor U9589 (N_9589,N_8367,N_9260);
or U9590 (N_9590,N_7269,N_7779);
nand U9591 (N_9591,N_7677,N_7636);
and U9592 (N_9592,N_7932,N_6751);
and U9593 (N_9593,N_6460,N_6987);
nor U9594 (N_9594,N_7997,N_6909);
nor U9595 (N_9595,N_8058,N_7639);
or U9596 (N_9596,N_7217,N_7198);
nand U9597 (N_9597,N_6712,N_6961);
or U9598 (N_9598,N_7839,N_9164);
or U9599 (N_9599,N_9217,N_9206);
and U9600 (N_9600,N_9143,N_9065);
nor U9601 (N_9601,N_7515,N_6908);
nor U9602 (N_9602,N_7983,N_6581);
and U9603 (N_9603,N_9196,N_9031);
or U9604 (N_9604,N_7057,N_7262);
nand U9605 (N_9605,N_8542,N_7439);
nand U9606 (N_9606,N_7469,N_7717);
or U9607 (N_9607,N_9316,N_8471);
or U9608 (N_9608,N_7543,N_8879);
and U9609 (N_9609,N_8292,N_7243);
or U9610 (N_9610,N_6859,N_7766);
or U9611 (N_9611,N_7251,N_7273);
or U9612 (N_9612,N_7996,N_6284);
xor U9613 (N_9613,N_8268,N_6867);
and U9614 (N_9614,N_8534,N_8803);
nor U9615 (N_9615,N_8028,N_7410);
and U9616 (N_9616,N_6954,N_8155);
or U9617 (N_9617,N_7596,N_7268);
xor U9618 (N_9618,N_8396,N_8561);
and U9619 (N_9619,N_7857,N_7687);
nor U9620 (N_9620,N_7207,N_8666);
nor U9621 (N_9621,N_6887,N_6360);
nor U9622 (N_9622,N_7741,N_8231);
xor U9623 (N_9623,N_9119,N_7924);
or U9624 (N_9624,N_8018,N_7690);
xnor U9625 (N_9625,N_8194,N_8886);
nor U9626 (N_9626,N_7508,N_7761);
nor U9627 (N_9627,N_7034,N_6948);
nand U9628 (N_9628,N_7817,N_7625);
nand U9629 (N_9629,N_9025,N_6695);
nor U9630 (N_9630,N_7068,N_6994);
and U9631 (N_9631,N_8921,N_7249);
and U9632 (N_9632,N_8066,N_6570);
nand U9633 (N_9633,N_7876,N_9114);
nand U9634 (N_9634,N_6513,N_8123);
nor U9635 (N_9635,N_8775,N_8806);
nand U9636 (N_9636,N_6784,N_6582);
nand U9637 (N_9637,N_6432,N_8366);
nand U9638 (N_9638,N_6898,N_7328);
nand U9639 (N_9639,N_7016,N_7686);
nand U9640 (N_9640,N_9177,N_9182);
xnor U9641 (N_9641,N_9091,N_6311);
nor U9642 (N_9642,N_7116,N_8257);
nand U9643 (N_9643,N_7044,N_7187);
xnor U9644 (N_9644,N_7611,N_7282);
nand U9645 (N_9645,N_8311,N_8457);
nor U9646 (N_9646,N_7831,N_7758);
nor U9647 (N_9647,N_9234,N_6336);
or U9648 (N_9648,N_6545,N_9075);
nand U9649 (N_9649,N_9085,N_9191);
or U9650 (N_9650,N_7402,N_8805);
or U9651 (N_9651,N_8295,N_8877);
nand U9652 (N_9652,N_7858,N_7476);
nor U9653 (N_9653,N_8585,N_9340);
or U9654 (N_9654,N_6721,N_8749);
or U9655 (N_9655,N_7641,N_6273);
nor U9656 (N_9656,N_6686,N_7164);
nor U9657 (N_9657,N_9367,N_6474);
nor U9658 (N_9658,N_9276,N_6315);
nor U9659 (N_9659,N_6777,N_7468);
nor U9660 (N_9660,N_9272,N_7862);
nand U9661 (N_9661,N_8081,N_7404);
nand U9662 (N_9662,N_8244,N_6620);
and U9663 (N_9663,N_8204,N_8810);
or U9664 (N_9664,N_6855,N_7474);
or U9665 (N_9665,N_6655,N_6966);
nand U9666 (N_9666,N_8282,N_8873);
and U9667 (N_9667,N_8654,N_8325);
xor U9668 (N_9668,N_9159,N_7663);
nand U9669 (N_9669,N_7311,N_7266);
and U9670 (N_9670,N_9295,N_6266);
nor U9671 (N_9671,N_7696,N_8029);
and U9672 (N_9672,N_6599,N_8864);
or U9673 (N_9673,N_8500,N_8671);
nor U9674 (N_9674,N_6255,N_8684);
nor U9675 (N_9675,N_7946,N_6251);
or U9676 (N_9676,N_6536,N_7091);
nor U9677 (N_9677,N_7706,N_6272);
nand U9678 (N_9678,N_8497,N_9092);
xor U9679 (N_9679,N_7790,N_8125);
nor U9680 (N_9680,N_6439,N_8054);
or U9681 (N_9681,N_7406,N_8281);
nand U9682 (N_9682,N_7989,N_8526);
and U9683 (N_9683,N_8381,N_7729);
and U9684 (N_9684,N_6736,N_7277);
and U9685 (N_9685,N_6488,N_6491);
and U9686 (N_9686,N_7901,N_8263);
xnor U9687 (N_9687,N_8902,N_9067);
and U9688 (N_9688,N_9158,N_7679);
and U9689 (N_9689,N_7418,N_8429);
xnor U9690 (N_9690,N_7320,N_6326);
nand U9691 (N_9691,N_9212,N_8792);
nand U9692 (N_9692,N_6321,N_7958);
and U9693 (N_9693,N_7444,N_6647);
nor U9694 (N_9694,N_6824,N_6433);
nor U9695 (N_9695,N_7950,N_6897);
nand U9696 (N_9696,N_7080,N_8610);
nand U9697 (N_9697,N_7617,N_7137);
nand U9698 (N_9698,N_7133,N_7433);
nand U9699 (N_9699,N_7921,N_7748);
and U9700 (N_9700,N_8399,N_9105);
xnor U9701 (N_9701,N_7427,N_9248);
and U9702 (N_9702,N_6957,N_7258);
or U9703 (N_9703,N_6960,N_6972);
nor U9704 (N_9704,N_7868,N_8033);
or U9705 (N_9705,N_6310,N_8019);
and U9706 (N_9706,N_8346,N_9147);
or U9707 (N_9707,N_7803,N_8875);
and U9708 (N_9708,N_7685,N_8602);
and U9709 (N_9709,N_9324,N_9294);
nand U9710 (N_9710,N_6373,N_6401);
or U9711 (N_9711,N_6846,N_9121);
or U9712 (N_9712,N_7411,N_6549);
and U9713 (N_9713,N_9253,N_6328);
and U9714 (N_9714,N_7664,N_7743);
xor U9715 (N_9715,N_6924,N_7825);
nand U9716 (N_9716,N_6370,N_6258);
and U9717 (N_9717,N_6996,N_9116);
and U9718 (N_9718,N_8002,N_6860);
nand U9719 (N_9719,N_6821,N_9093);
nor U9720 (N_9720,N_9277,N_8540);
or U9721 (N_9721,N_6903,N_6685);
nor U9722 (N_9722,N_8243,N_7612);
xor U9723 (N_9723,N_7848,N_8932);
nor U9724 (N_9724,N_7391,N_6933);
or U9725 (N_9725,N_8344,N_6446);
and U9726 (N_9726,N_6816,N_6786);
and U9727 (N_9727,N_7605,N_8898);
or U9728 (N_9728,N_6480,N_7926);
xor U9729 (N_9729,N_7576,N_6340);
nand U9730 (N_9730,N_9355,N_7710);
and U9731 (N_9731,N_8401,N_8831);
and U9732 (N_9732,N_6863,N_7842);
and U9733 (N_9733,N_8168,N_7021);
nand U9734 (N_9734,N_7139,N_7298);
xnor U9735 (N_9735,N_8402,N_8384);
nand U9736 (N_9736,N_8478,N_7011);
nand U9737 (N_9737,N_6973,N_8196);
xnor U9738 (N_9738,N_6603,N_8207);
xnor U9739 (N_9739,N_6274,N_7052);
nand U9740 (N_9740,N_7902,N_8957);
nand U9741 (N_9741,N_9089,N_8393);
nand U9742 (N_9742,N_7373,N_7178);
nand U9743 (N_9743,N_7979,N_7424);
or U9744 (N_9744,N_8562,N_7502);
xnor U9745 (N_9745,N_8147,N_7344);
or U9746 (N_9746,N_8672,N_7742);
nor U9747 (N_9747,N_6733,N_7471);
nor U9748 (N_9748,N_7190,N_6422);
xor U9749 (N_9749,N_6631,N_9363);
nand U9750 (N_9750,N_6363,N_8907);
and U9751 (N_9751,N_8524,N_9168);
nand U9752 (N_9752,N_7465,N_7807);
and U9753 (N_9753,N_6557,N_8612);
and U9754 (N_9754,N_8466,N_8359);
or U9755 (N_9755,N_9108,N_6283);
nor U9756 (N_9756,N_8139,N_8126);
or U9757 (N_9757,N_6590,N_8474);
xor U9758 (N_9758,N_6466,N_8427);
or U9759 (N_9759,N_6919,N_7019);
nand U9760 (N_9760,N_8920,N_9060);
nand U9761 (N_9761,N_8929,N_7304);
nand U9762 (N_9762,N_6312,N_8370);
nand U9763 (N_9763,N_8239,N_8980);
nand U9764 (N_9764,N_8755,N_7064);
nand U9765 (N_9765,N_9045,N_7521);
and U9766 (N_9766,N_9281,N_7118);
nand U9767 (N_9767,N_9117,N_7615);
or U9768 (N_9768,N_7705,N_7121);
nor U9769 (N_9769,N_7491,N_8143);
xor U9770 (N_9770,N_6951,N_8639);
nand U9771 (N_9771,N_8543,N_7867);
xnor U9772 (N_9772,N_6902,N_7230);
or U9773 (N_9773,N_7144,N_7828);
nand U9774 (N_9774,N_7704,N_8044);
xor U9775 (N_9775,N_7972,N_6668);
nor U9776 (N_9776,N_8716,N_9165);
or U9777 (N_9777,N_6366,N_8617);
and U9778 (N_9778,N_9084,N_7787);
or U9779 (N_9779,N_6872,N_8498);
nor U9780 (N_9780,N_8188,N_6375);
and U9781 (N_9781,N_6787,N_8945);
nor U9782 (N_9782,N_6888,N_7265);
nand U9783 (N_9783,N_7903,N_7199);
or U9784 (N_9784,N_6807,N_8571);
and U9785 (N_9785,N_8136,N_8721);
nand U9786 (N_9786,N_8009,N_6945);
and U9787 (N_9787,N_7195,N_6976);
or U9788 (N_9788,N_7899,N_8849);
and U9789 (N_9789,N_7563,N_7241);
nand U9790 (N_9790,N_8868,N_6327);
or U9791 (N_9791,N_8698,N_7560);
xnor U9792 (N_9792,N_8997,N_8390);
nand U9793 (N_9793,N_9337,N_9268);
nand U9794 (N_9794,N_8970,N_8274);
nor U9795 (N_9795,N_7067,N_9349);
nor U9796 (N_9796,N_8145,N_6528);
xnor U9797 (N_9797,N_7236,N_7087);
xor U9798 (N_9798,N_7252,N_7386);
nand U9799 (N_9799,N_6531,N_8469);
and U9800 (N_9800,N_8754,N_9252);
nor U9801 (N_9801,N_9370,N_6814);
or U9802 (N_9802,N_6506,N_7542);
nand U9803 (N_9803,N_7171,N_9140);
nor U9804 (N_9804,N_7744,N_9188);
or U9805 (N_9805,N_8545,N_8736);
or U9806 (N_9806,N_7886,N_9204);
nor U9807 (N_9807,N_6659,N_9373);
nand U9808 (N_9808,N_6342,N_9222);
and U9809 (N_9809,N_6519,N_6598);
nor U9810 (N_9810,N_6358,N_6623);
nand U9811 (N_9811,N_6636,N_9050);
nor U9812 (N_9812,N_6642,N_7040);
and U9813 (N_9813,N_6431,N_8796);
nand U9814 (N_9814,N_6338,N_8911);
xnor U9815 (N_9815,N_6740,N_8374);
nand U9816 (N_9816,N_7510,N_7545);
nand U9817 (N_9817,N_7117,N_7949);
and U9818 (N_9818,N_8655,N_7245);
and U9819 (N_9819,N_6459,N_7362);
and U9820 (N_9820,N_7102,N_7234);
and U9821 (N_9821,N_7169,N_9244);
or U9822 (N_9822,N_7773,N_8592);
or U9823 (N_9823,N_7816,N_8919);
nand U9824 (N_9824,N_7523,N_9166);
nor U9825 (N_9825,N_6464,N_6454);
or U9826 (N_9826,N_8832,N_7208);
nor U9827 (N_9827,N_8111,N_9304);
or U9828 (N_9828,N_9080,N_7781);
nor U9829 (N_9829,N_8385,N_7074);
nor U9830 (N_9830,N_8286,N_8495);
nor U9831 (N_9831,N_7740,N_7235);
nor U9832 (N_9832,N_7645,N_7952);
or U9833 (N_9833,N_6651,N_8528);
nor U9834 (N_9834,N_8237,N_7840);
nand U9835 (N_9835,N_8001,N_7453);
nand U9836 (N_9836,N_6362,N_9041);
and U9837 (N_9837,N_7960,N_8241);
xor U9838 (N_9838,N_6257,N_7897);
and U9839 (N_9839,N_9122,N_7933);
xnor U9840 (N_9840,N_9109,N_9263);
xor U9841 (N_9841,N_6657,N_6836);
and U9842 (N_9842,N_9173,N_7076);
nand U9843 (N_9843,N_6296,N_6495);
xor U9844 (N_9844,N_8063,N_7089);
and U9845 (N_9845,N_7088,N_7316);
nand U9846 (N_9846,N_7115,N_9099);
or U9847 (N_9847,N_8422,N_6467);
nor U9848 (N_9848,N_8262,N_8299);
nor U9849 (N_9849,N_6555,N_9038);
or U9850 (N_9850,N_7824,N_6441);
nor U9851 (N_9851,N_7317,N_8568);
and U9852 (N_9852,N_8939,N_6731);
nor U9853 (N_9853,N_6654,N_8522);
or U9854 (N_9854,N_9280,N_6447);
and U9855 (N_9855,N_8460,N_8677);
and U9856 (N_9856,N_8614,N_7366);
nor U9857 (N_9857,N_8989,N_6813);
nor U9858 (N_9858,N_6288,N_8130);
nor U9859 (N_9859,N_8827,N_7229);
xor U9860 (N_9860,N_7028,N_7110);
nor U9861 (N_9861,N_8795,N_7130);
or U9862 (N_9862,N_6761,N_9321);
and U9863 (N_9863,N_9056,N_8170);
nor U9864 (N_9864,N_7194,N_7765);
and U9865 (N_9865,N_6426,N_7640);
and U9866 (N_9866,N_8538,N_8210);
or U9867 (N_9867,N_7096,N_6490);
nor U9868 (N_9868,N_6927,N_7808);
or U9869 (N_9869,N_9103,N_7993);
or U9870 (N_9870,N_8297,N_6831);
or U9871 (N_9871,N_7700,N_8548);
and U9872 (N_9872,N_6778,N_9032);
nor U9873 (N_9873,N_6594,N_9326);
nor U9874 (N_9874,N_8567,N_8948);
and U9875 (N_9875,N_7498,N_9303);
nor U9876 (N_9876,N_8378,N_6964);
nor U9877 (N_9877,N_6567,N_7455);
nor U9878 (N_9878,N_9057,N_8043);
nand U9879 (N_9879,N_8079,N_8481);
and U9880 (N_9880,N_8010,N_6399);
or U9881 (N_9881,N_8071,N_8729);
nor U9882 (N_9882,N_7943,N_8737);
or U9883 (N_9883,N_7077,N_7737);
xor U9884 (N_9884,N_6628,N_6293);
or U9885 (N_9885,N_7322,N_8714);
nor U9886 (N_9886,N_7995,N_6568);
xor U9887 (N_9887,N_6809,N_7084);
or U9888 (N_9888,N_7200,N_7837);
nand U9889 (N_9889,N_7863,N_7732);
nand U9890 (N_9890,N_8117,N_7204);
and U9891 (N_9891,N_6335,N_6837);
and U9892 (N_9892,N_6881,N_7128);
nor U9893 (N_9893,N_7552,N_7365);
nor U9894 (N_9894,N_8256,N_7313);
nand U9895 (N_9895,N_9357,N_7334);
and U9896 (N_9896,N_7147,N_7676);
and U9897 (N_9897,N_7292,N_8072);
nor U9898 (N_9898,N_9298,N_7179);
nor U9899 (N_9899,N_7497,N_8951);
nand U9900 (N_9900,N_9064,N_7355);
nand U9901 (N_9901,N_8856,N_9088);
or U9902 (N_9902,N_6870,N_6779);
nor U9903 (N_9903,N_8333,N_6574);
nor U9904 (N_9904,N_6470,N_8822);
nor U9905 (N_9905,N_6986,N_7397);
and U9906 (N_9906,N_7036,N_7894);
and U9907 (N_9907,N_8407,N_6732);
nor U9908 (N_9908,N_8065,N_7407);
nor U9909 (N_9909,N_6918,N_8405);
nand U9910 (N_9910,N_8352,N_7712);
nand U9911 (N_9911,N_6532,N_7835);
nand U9912 (N_9912,N_8383,N_7638);
or U9913 (N_9913,N_8166,N_6920);
nand U9914 (N_9914,N_8981,N_6958);
or U9915 (N_9915,N_8369,N_7283);
or U9916 (N_9916,N_6269,N_9297);
nor U9917 (N_9917,N_8308,N_8348);
nand U9918 (N_9918,N_7927,N_7721);
nor U9919 (N_9919,N_7719,N_7880);
xnor U9920 (N_9920,N_8978,N_7378);
and U9921 (N_9921,N_9139,N_7900);
or U9922 (N_9922,N_8004,N_7872);
nand U9923 (N_9923,N_9054,N_7874);
nand U9924 (N_9924,N_8057,N_8506);
and U9925 (N_9925,N_8869,N_6835);
or U9926 (N_9926,N_6704,N_6670);
or U9927 (N_9927,N_7870,N_7736);
nor U9928 (N_9928,N_6597,N_8692);
and U9929 (N_9929,N_9264,N_9195);
nand U9930 (N_9930,N_6742,N_7430);
and U9931 (N_9931,N_7738,N_7162);
and U9932 (N_9932,N_9180,N_8444);
or U9933 (N_9933,N_7479,N_9199);
nor U9934 (N_9934,N_7338,N_7184);
xnor U9935 (N_9935,N_8480,N_8465);
and U9936 (N_9936,N_7216,N_8848);
xor U9937 (N_9937,N_7448,N_7668);
nor U9938 (N_9938,N_8515,N_6760);
and U9939 (N_9939,N_7610,N_8199);
and U9940 (N_9940,N_7871,N_7970);
or U9941 (N_9941,N_7473,N_8435);
and U9942 (N_9942,N_7367,N_6880);
nand U9943 (N_9943,N_8104,N_6320);
and U9944 (N_9944,N_6997,N_8688);
and U9945 (N_9945,N_8767,N_8739);
nand U9946 (N_9946,N_8600,N_8866);
and U9947 (N_9947,N_6465,N_7403);
nand U9948 (N_9948,N_7346,N_8575);
or U9949 (N_9949,N_8240,N_6864);
and U9950 (N_9950,N_7533,N_6602);
and U9951 (N_9951,N_7205,N_6417);
or U9952 (N_9952,N_7789,N_6741);
and U9953 (N_9953,N_7049,N_8151);
and U9954 (N_9954,N_6611,N_9299);
and U9955 (N_9955,N_8566,N_6692);
nor U9956 (N_9956,N_7210,N_8255);
and U9957 (N_9957,N_9006,N_8783);
and U9958 (N_9958,N_8909,N_8228);
and U9959 (N_9959,N_6523,N_6295);
nor U9960 (N_9960,N_8316,N_7321);
xnor U9961 (N_9961,N_7945,N_8723);
and U9962 (N_9962,N_6609,N_7935);
nor U9963 (N_9963,N_7733,N_9291);
xnor U9964 (N_9964,N_6476,N_7695);
xnor U9965 (N_9965,N_8025,N_8450);
and U9966 (N_9966,N_6483,N_6517);
and U9967 (N_9967,N_7227,N_7401);
xnor U9968 (N_9968,N_6632,N_8144);
or U9969 (N_9969,N_6508,N_6766);
nor U9970 (N_9970,N_7270,N_7659);
or U9971 (N_9971,N_7323,N_8045);
or U9972 (N_9972,N_8421,N_7529);
nand U9973 (N_9973,N_7535,N_7548);
nand U9974 (N_9974,N_8993,N_8068);
nand U9975 (N_9975,N_7584,N_6616);
nand U9976 (N_9976,N_6479,N_8722);
xor U9977 (N_9977,N_6891,N_8603);
and U9978 (N_9978,N_7974,N_7018);
or U9979 (N_9979,N_8703,N_9022);
xor U9980 (N_9980,N_8974,N_7838);
nor U9981 (N_9981,N_7672,N_6884);
or U9982 (N_9982,N_9309,N_8090);
and U9983 (N_9983,N_6699,N_6842);
nand U9984 (N_9984,N_8861,N_6412);
or U9985 (N_9985,N_9347,N_9258);
nor U9986 (N_9986,N_9352,N_8927);
nor U9987 (N_9987,N_8386,N_8901);
or U9988 (N_9988,N_9170,N_8455);
or U9989 (N_9989,N_6613,N_7186);
nand U9990 (N_9990,N_6906,N_9339);
nor U9991 (N_9991,N_9035,N_8683);
or U9992 (N_9992,N_8254,N_6660);
nand U9993 (N_9993,N_6526,N_6728);
nor U9994 (N_9994,N_6757,N_6334);
nand U9995 (N_9995,N_6989,N_8142);
nand U9996 (N_9996,N_9020,N_7777);
and U9997 (N_9997,N_6382,N_8680);
and U9998 (N_9998,N_7213,N_6681);
or U9999 (N_9999,N_8828,N_7854);
xor U10000 (N_10000,N_9220,N_6408);
and U10001 (N_10001,N_8628,N_7833);
or U10002 (N_10002,N_9079,N_7674);
nor U10003 (N_10003,N_8777,N_9215);
and U10004 (N_10004,N_9000,N_9137);
nor U10005 (N_10005,N_7923,N_7920);
or U10006 (N_10006,N_6684,N_6420);
or U10007 (N_10007,N_6308,N_8815);
nand U10008 (N_10008,N_7601,N_8572);
and U10009 (N_10009,N_6332,N_9005);
nor U10010 (N_10010,N_8486,N_6378);
or U10011 (N_10011,N_8670,N_9219);
or U10012 (N_10012,N_6866,N_7324);
or U10013 (N_10013,N_8250,N_6518);
and U10014 (N_10014,N_7452,N_7832);
and U10015 (N_10015,N_8745,N_7882);
and U10016 (N_10016,N_8760,N_8493);
or U10017 (N_10017,N_8797,N_7845);
or U10018 (N_10018,N_7627,N_6497);
or U10019 (N_10019,N_6851,N_7420);
nand U10020 (N_10020,N_9225,N_9179);
and U10021 (N_10021,N_8011,N_7774);
or U10022 (N_10022,N_8017,N_9126);
nor U10023 (N_10023,N_9230,N_9176);
and U10024 (N_10024,N_8837,N_6932);
and U10025 (N_10025,N_7168,N_8823);
and U10026 (N_10026,N_6489,N_7811);
nor U10027 (N_10027,N_7805,N_6978);
xor U10028 (N_10028,N_8418,N_8133);
and U10029 (N_10029,N_7735,N_8119);
and U10030 (N_10030,N_7371,N_7368);
xor U10031 (N_10031,N_7528,N_7852);
or U10032 (N_10032,N_6806,N_8326);
and U10033 (N_10033,N_9229,N_8847);
xnor U10034 (N_10034,N_7054,N_7033);
or U10035 (N_10035,N_7531,N_8584);
xor U10036 (N_10036,N_8836,N_7988);
or U10037 (N_10037,N_8108,N_7098);
nand U10038 (N_10038,N_9197,N_8387);
nand U10039 (N_10039,N_9211,N_6525);
nand U10040 (N_10040,N_8461,N_6394);
xor U10041 (N_10041,N_8362,N_6788);
nor U10042 (N_10042,N_7534,N_7326);
nor U10043 (N_10043,N_7821,N_6810);
nand U10044 (N_10044,N_6650,N_6970);
nor U10045 (N_10045,N_8955,N_6588);
and U10046 (N_10046,N_7232,N_7379);
nand U10047 (N_10047,N_6522,N_7869);
nand U10048 (N_10048,N_6383,N_6834);
or U10049 (N_10049,N_7038,N_9312);
and U10050 (N_10050,N_9012,N_9071);
and U10051 (N_10051,N_8665,N_6965);
nand U10052 (N_10052,N_8811,N_7622);
nor U10053 (N_10053,N_7916,N_6316);
nor U10054 (N_10054,N_7912,N_8964);
or U10055 (N_10055,N_7048,N_6270);
nor U10056 (N_10056,N_6661,N_8520);
nor U10057 (N_10057,N_8287,N_7660);
nand U10058 (N_10058,N_7457,N_8900);
nand U10059 (N_10059,N_7175,N_7603);
and U10060 (N_10060,N_6979,N_6652);
and U10061 (N_10061,N_7745,N_6499);
nand U10062 (N_10062,N_9073,N_7486);
nor U10063 (N_10063,N_7634,N_8530);
or U10064 (N_10064,N_6912,N_8681);
nand U10065 (N_10065,N_8718,N_7557);
nand U10066 (N_10066,N_8034,N_8699);
or U10067 (N_10067,N_6701,N_7384);
nor U10068 (N_10068,N_6940,N_7393);
xor U10069 (N_10069,N_8030,N_8328);
or U10070 (N_10070,N_8024,N_6361);
or U10071 (N_10071,N_7796,N_6907);
and U10072 (N_10072,N_9034,N_6850);
nor U10073 (N_10073,N_7460,N_8503);
or U10074 (N_10074,N_7231,N_6605);
or U10075 (N_10075,N_7849,N_8659);
and U10076 (N_10076,N_7830,N_6754);
and U10077 (N_10077,N_8786,N_8110);
nor U10078 (N_10078,N_9343,N_7157);
nor U10079 (N_10079,N_7182,N_7223);
nand U10080 (N_10080,N_6463,N_6279);
nand U10081 (N_10081,N_6304,N_7575);
and U10082 (N_10082,N_7039,N_8674);
nand U10083 (N_10083,N_9290,N_8512);
and U10084 (N_10084,N_8616,N_9292);
and U10085 (N_10085,N_7855,N_7072);
and U10086 (N_10086,N_8531,N_7595);
xor U10087 (N_10087,N_6649,N_7146);
and U10088 (N_10088,N_6707,N_7348);
nand U10089 (N_10089,N_6595,N_6610);
nand U10090 (N_10090,N_7984,N_6414);
or U10091 (N_10091,N_7302,N_7225);
nor U10092 (N_10092,N_6729,N_8658);
xnor U10093 (N_10093,N_6743,N_8787);
or U10094 (N_10094,N_8288,N_7466);
nand U10095 (N_10095,N_7701,N_7678);
nand U10096 (N_10096,N_6556,N_7127);
and U10097 (N_10097,N_7859,N_7599);
nor U10098 (N_10098,N_8193,N_6292);
nor U10099 (N_10099,N_8060,N_9001);
or U10100 (N_10100,N_8491,N_8705);
nand U10101 (N_10101,N_7022,N_8559);
or U10102 (N_10102,N_6614,N_8678);
or U10103 (N_10103,N_9070,N_6737);
and U10104 (N_10104,N_7398,N_6999);
nand U10105 (N_10105,N_8649,N_7183);
and U10106 (N_10106,N_6969,N_7546);
xor U10107 (N_10107,N_8570,N_6758);
or U10108 (N_10108,N_6573,N_8410);
nor U10109 (N_10109,N_6808,N_8735);
nand U10110 (N_10110,N_7561,N_7718);
or U10111 (N_10111,N_6507,N_9145);
nor U10112 (N_10112,N_7877,N_8404);
and U10113 (N_10113,N_9118,N_8246);
and U10114 (N_10114,N_8137,N_8959);
and U10115 (N_10115,N_8468,N_7731);
or U10116 (N_10116,N_6896,N_7405);
nor U10117 (N_10117,N_8517,N_9059);
nand U10118 (N_10118,N_8950,N_8915);
or U10119 (N_10119,N_7437,N_7671);
or U10120 (N_10120,N_9151,N_6739);
nor U10121 (N_10121,N_7499,N_8413);
nand U10122 (N_10122,N_8590,N_6876);
xor U10123 (N_10123,N_8653,N_8890);
nor U10124 (N_10124,N_7944,N_7890);
nand U10125 (N_10125,N_6865,N_7522);
nand U10126 (N_10126,N_7209,N_7846);
nand U10127 (N_10127,N_7181,N_6691);
xor U10128 (N_10128,N_8756,N_8276);
or U10129 (N_10129,N_7904,N_8551);
nand U10130 (N_10130,N_7632,N_8361);
nor U10131 (N_10131,N_8965,N_8412);
or U10132 (N_10132,N_6256,N_6839);
and U10133 (N_10133,N_9021,N_8967);
nor U10134 (N_10134,N_8839,N_7381);
nand U10135 (N_10135,N_8202,N_9076);
and U10136 (N_10136,N_6750,N_8546);
and U10137 (N_10137,N_7573,N_8315);
nor U10138 (N_10138,N_8558,N_8400);
nand U10139 (N_10139,N_7250,N_7913);
nand U10140 (N_10140,N_6277,N_8555);
or U10141 (N_10141,N_7581,N_7644);
nand U10142 (N_10142,N_6698,N_6396);
nand U10143 (N_10143,N_8431,N_8859);
nor U10144 (N_10144,N_6820,N_6496);
nand U10145 (N_10145,N_7412,N_6539);
nor U10146 (N_10146,N_7915,N_6854);
xnor U10147 (N_10147,N_8163,N_8055);
and U10148 (N_10148,N_7284,N_8008);
xor U10149 (N_10149,N_6811,N_8473);
or U10150 (N_10150,N_8966,N_6803);
nand U10151 (N_10151,N_8991,N_8793);
or U10152 (N_10152,N_6406,N_7278);
and U10153 (N_10153,N_7488,N_7428);
nand U10154 (N_10154,N_6593,N_6450);
nand U10155 (N_10155,N_6625,N_9236);
or U10156 (N_10156,N_6829,N_9201);
nand U10157 (N_10157,N_7112,N_9364);
nand U10158 (N_10158,N_7327,N_6586);
and U10159 (N_10159,N_8285,N_8206);
xnor U10160 (N_10160,N_9332,N_7793);
nor U10161 (N_10161,N_8897,N_7594);
and U10162 (N_10162,N_6645,N_8036);
or U10163 (N_10163,N_8537,N_6794);
or U10164 (N_10164,N_8476,N_8092);
and U10165 (N_10165,N_8624,N_9267);
and U10166 (N_10166,N_9155,N_9051);
nand U10167 (N_10167,N_6875,N_8818);
xnor U10168 (N_10168,N_8667,N_7286);
or U10169 (N_10169,N_8596,N_8015);
nor U10170 (N_10170,N_7097,N_8986);
and U10171 (N_10171,N_8947,N_7160);
nand U10172 (N_10172,N_6843,N_8930);
or U10173 (N_10173,N_6302,N_6484);
and U10174 (N_10174,N_7172,N_8245);
or U10175 (N_10175,N_7630,N_7050);
nand U10176 (N_10176,N_6877,N_9261);
nand U10177 (N_10177,N_9322,N_6899);
nor U10178 (N_10178,N_7720,N_6826);
and U10179 (N_10179,N_7860,N_6510);
xnor U10180 (N_10180,N_8694,N_6330);
or U10181 (N_10181,N_6901,N_6857);
xor U10182 (N_10182,N_9366,N_8985);
or U10183 (N_10183,N_8916,N_8021);
or U10184 (N_10184,N_6416,N_7619);
nand U10185 (N_10185,N_8853,N_7888);
nor U10186 (N_10186,N_8462,N_7287);
or U10187 (N_10187,N_6485,N_7577);
nor U10188 (N_10188,N_7103,N_7907);
nor U10189 (N_10189,N_6905,N_8765);
or U10190 (N_10190,N_7319,N_8541);
nor U10191 (N_10191,N_7069,N_9213);
nand U10192 (N_10192,N_7541,N_7728);
and U10193 (N_10193,N_8944,N_6916);
and U10194 (N_10194,N_8271,N_8695);
or U10195 (N_10195,N_7620,N_6579);
nor U10196 (N_10196,N_6323,N_7734);
xnor U10197 (N_10197,N_8048,N_7683);
and U10198 (N_10198,N_7220,N_6325);
and U10199 (N_10199,N_6716,N_7306);
nor U10200 (N_10200,N_8124,N_7551);
nand U10201 (N_10201,N_8373,N_6456);
and U10202 (N_10202,N_7883,N_9259);
or U10203 (N_10203,N_8844,N_8499);
or U10204 (N_10204,N_7156,N_6847);
or U10205 (N_10205,N_8926,N_7844);
or U10206 (N_10206,N_6815,N_8406);
or U10207 (N_10207,N_7836,N_9090);
nor U10208 (N_10208,N_6537,N_7255);
nand U10209 (N_10209,N_8264,N_8310);
xnor U10210 (N_10210,N_8789,N_8483);
and U10211 (N_10211,N_7281,N_7513);
xor U10212 (N_10212,N_6804,N_9120);
nor U10213 (N_10213,N_6795,N_8436);
nor U10214 (N_10214,N_8379,N_8650);
and U10215 (N_10215,N_6309,N_7248);
nand U10216 (N_10216,N_8634,N_9152);
nor U10217 (N_10217,N_8843,N_6675);
or U10218 (N_10218,N_8109,N_8711);
xor U10219 (N_10219,N_6415,N_6276);
nor U10220 (N_10220,N_7374,N_7211);
nand U10221 (N_10221,N_9186,N_8580);
and U10222 (N_10222,N_8304,N_6547);
or U10223 (N_10223,N_8038,N_6962);
or U10224 (N_10224,N_7043,N_8931);
and U10225 (N_10225,N_6773,N_7459);
nor U10226 (N_10226,N_8016,N_8161);
or U10227 (N_10227,N_7120,N_9096);
nand U10228 (N_10228,N_7792,N_8946);
and U10229 (N_10229,N_8801,N_8442);
nand U10230 (N_10230,N_8417,N_9163);
nand U10231 (N_10231,N_6770,N_9110);
nand U10232 (N_10232,N_8968,N_7153);
xnor U10233 (N_10233,N_6353,N_8734);
and U10234 (N_10234,N_8870,N_6511);
nor U10235 (N_10235,N_7063,N_7041);
and U10236 (N_10236,N_7574,N_9323);
nor U10237 (N_10237,N_8425,N_9053);
nand U10238 (N_10238,N_9242,N_6428);
and U10239 (N_10239,N_6515,N_8663);
or U10240 (N_10240,N_9271,N_8956);
nand U10241 (N_10241,N_6637,N_8279);
nor U10242 (N_10242,N_6554,N_6981);
or U10243 (N_10243,N_6475,N_6407);
xor U10244 (N_10244,N_8800,N_6747);
and U10245 (N_10245,N_9239,N_7356);
and U10246 (N_10246,N_8779,N_8645);
or U10247 (N_10247,N_8363,N_8180);
nor U10248 (N_10248,N_9275,N_8556);
nor U10249 (N_10249,N_9192,N_9302);
nand U10250 (N_10250,N_6643,N_6690);
nor U10251 (N_10251,N_8988,N_8355);
xor U10252 (N_10252,N_8007,N_7801);
and U10253 (N_10253,N_7682,N_7778);
nand U10254 (N_10254,N_6324,N_6405);
nand U10255 (N_10255,N_8129,N_8160);
xor U10256 (N_10256,N_8829,N_6259);
and U10257 (N_10257,N_8414,N_8376);
nor U10258 (N_10258,N_8265,N_8235);
or U10259 (N_10259,N_9036,N_8741);
nor U10260 (N_10260,N_7775,N_6818);
and U10261 (N_10261,N_7017,N_8424);
nand U10262 (N_10262,N_8889,N_6291);
nor U10263 (N_10263,N_7485,N_6744);
and U10264 (N_10264,N_9142,N_6845);
or U10265 (N_10265,N_7878,N_7046);
or U10266 (N_10266,N_8484,N_6841);
nand U10267 (N_10267,N_7342,N_8162);
nand U10268 (N_10268,N_8338,N_9154);
nor U10269 (N_10269,N_8191,N_8447);
nand U10270 (N_10270,N_6856,N_6797);
nand U10271 (N_10271,N_6442,N_7030);
nand U10272 (N_10272,N_7105,N_6424);
nand U10273 (N_10273,N_8690,N_7604);
nand U10274 (N_10274,N_6410,N_9002);
nand U10275 (N_10275,N_6271,N_8707);
nand U10276 (N_10276,N_8937,N_6977);
nor U10277 (N_10277,N_8080,N_7307);
or U10278 (N_10278,N_8440,N_8761);
nor U10279 (N_10279,N_6791,N_7289);
and U10280 (N_10280,N_9226,N_7254);
or U10281 (N_10281,N_6516,N_8197);
nand U10282 (N_10282,N_9214,N_8284);
nand U10283 (N_10283,N_9086,N_6756);
and U10284 (N_10284,N_7739,N_6524);
nand U10285 (N_10285,N_6578,N_9049);
and U10286 (N_10286,N_9241,N_7001);
nor U10287 (N_10287,N_7990,N_9224);
or U10288 (N_10288,N_6674,N_6398);
and U10289 (N_10289,N_7606,N_9017);
or U10290 (N_10290,N_6369,N_8527);
and U10291 (N_10291,N_8083,N_7730);
nor U10292 (N_10292,N_7345,N_7746);
and U10293 (N_10293,N_7628,N_9245);
xor U10294 (N_10294,N_8676,N_7905);
or U10295 (N_10295,N_7083,N_7806);
nand U10296 (N_10296,N_7349,N_8012);
or U10297 (N_10297,N_7853,N_9115);
and U10298 (N_10298,N_8183,N_7942);
and U10299 (N_10299,N_8159,N_9270);
xnor U10300 (N_10300,N_6992,N_8764);
and U10301 (N_10301,N_9069,N_6849);
nor U10302 (N_10302,N_8657,N_8327);
nor U10303 (N_10303,N_9334,N_8428);
xor U10304 (N_10304,N_7413,N_8095);
nand U10305 (N_10305,N_9368,N_7015);
and U10306 (N_10306,N_7148,N_6462);
and U10307 (N_10307,N_8807,N_8039);
nand U10308 (N_10308,N_7496,N_9282);
xor U10309 (N_10309,N_8582,N_8172);
nor U10310 (N_10310,N_8863,N_7582);
or U10311 (N_10311,N_8205,N_8230);
or U10312 (N_10312,N_8135,N_6727);
nor U10313 (N_10313,N_8704,N_8887);
and U10314 (N_10314,N_8232,N_8357);
nor U10315 (N_10315,N_6387,N_7818);
nand U10316 (N_10316,N_7451,N_7467);
nor U10317 (N_10317,N_8933,N_7493);
nor U10318 (N_10318,N_8731,N_8280);
or U10319 (N_10319,N_7908,N_8423);
or U10320 (N_10320,N_8249,N_6268);
nand U10321 (N_10321,N_9287,N_7294);
nand U10322 (N_10322,N_8434,N_8408);
nand U10323 (N_10323,N_7315,N_8896);
nor U10324 (N_10324,N_7059,N_7425);
nand U10325 (N_10325,N_8586,N_8996);
and U10326 (N_10326,N_7713,N_8432);
nand U10327 (N_10327,N_6388,N_7056);
nand U10328 (N_10328,N_9185,N_6900);
xor U10329 (N_10329,N_6926,N_7965);
and U10330 (N_10330,N_6583,N_7487);
nand U10331 (N_10331,N_9133,N_9190);
xor U10332 (N_10332,N_8872,N_8216);
nor U10333 (N_10333,N_6558,N_8132);
nor U10334 (N_10334,N_6560,N_8662);
and U10335 (N_10335,N_9042,N_7843);
or U10336 (N_10336,N_7856,N_8740);
nand U10337 (N_10337,N_6922,N_6347);
and U10338 (N_10338,N_8314,N_8652);
and U10339 (N_10339,N_7763,N_8623);
and U10340 (N_10340,N_9171,N_8685);
or U10341 (N_10341,N_9255,N_8093);
nand U10342 (N_10342,N_8040,N_9061);
or U10343 (N_10343,N_7567,N_9351);
and U10344 (N_10344,N_8182,N_9228);
nand U10345 (N_10345,N_8893,N_7108);
nand U10346 (N_10346,N_8715,N_7090);
nand U10347 (N_10347,N_8336,N_7895);
nand U10348 (N_10348,N_8846,N_8064);
nor U10349 (N_10349,N_7966,N_9128);
and U10350 (N_10350,N_7891,N_6753);
nand U10351 (N_10351,N_8809,N_8732);
nand U10352 (N_10352,N_8131,N_8682);
xor U10353 (N_10353,N_6402,N_9157);
and U10354 (N_10354,N_8458,N_8332);
or U10355 (N_10355,N_8878,N_7815);
and U10356 (N_10356,N_7085,N_6562);
xor U10357 (N_10357,N_6680,N_7122);
or U10358 (N_10358,N_7073,N_7847);
or U10359 (N_10359,N_8027,N_9249);
xor U10360 (N_10360,N_6949,N_9130);
and U10361 (N_10361,N_8037,N_6600);
or U10362 (N_10362,N_6921,N_6985);
and U10363 (N_10363,N_7261,N_7027);
and U10364 (N_10364,N_7490,N_6862);
and U10365 (N_10365,N_6893,N_7655);
and U10366 (N_10366,N_8841,N_7711);
and U10367 (N_10367,N_8134,N_6626);
nand U10368 (N_10368,N_9127,N_6693);
nand U10369 (N_10369,N_6634,N_8184);
and U10370 (N_10370,N_6601,N_8851);
and U10371 (N_10371,N_7214,N_8389);
or U10372 (N_10372,N_6640,N_7994);
nand U10373 (N_10373,N_8673,N_8114);
xnor U10374 (N_10374,N_6959,N_8941);
nand U10375 (N_10375,N_7520,N_8391);
and U10376 (N_10376,N_7176,N_8923);
or U10377 (N_10377,N_8814,N_8798);
nor U10378 (N_10378,N_7633,N_6801);
nor U10379 (N_10379,N_8727,N_8977);
nor U10380 (N_10380,N_8942,N_6664);
nor U10381 (N_10381,N_6882,N_6689);
or U10382 (N_10382,N_6929,N_6381);
and U10383 (N_10383,N_8774,N_7753);
or U10384 (N_10384,N_7238,N_6341);
nand U10385 (N_10385,N_8999,N_8272);
or U10386 (N_10386,N_6451,N_7930);
xnor U10387 (N_10387,N_9336,N_7020);
xnor U10388 (N_10388,N_8190,N_8470);
nand U10389 (N_10389,N_7060,N_9342);
nor U10390 (N_10390,N_8320,N_8635);
nor U10391 (N_10391,N_8816,N_9284);
or U10392 (N_10392,N_6822,N_6722);
and U10393 (N_10393,N_6344,N_7986);
or U10394 (N_10394,N_8140,N_8181);
and U10395 (N_10395,N_9082,N_7221);
nor U10396 (N_10396,N_9040,N_7196);
or U10397 (N_10397,N_7377,N_8696);
nand U10398 (N_10398,N_6404,N_6571);
and U10399 (N_10399,N_6789,N_6800);
or U10400 (N_10400,N_7569,N_8504);
xor U10401 (N_10401,N_6910,N_8519);
and U10402 (N_10402,N_8998,N_8179);
nand U10403 (N_10403,N_8047,N_8576);
or U10404 (N_10404,N_9315,N_7301);
and U10405 (N_10405,N_7131,N_8419);
nor U10406 (N_10406,N_6799,N_8799);
xnor U10407 (N_10407,N_9044,N_7106);
nand U10408 (N_10408,N_6494,N_7955);
nor U10409 (N_10409,N_6253,N_7957);
or U10410 (N_10410,N_8633,N_6472);
nor U10411 (N_10411,N_6830,N_7961);
nor U10412 (N_10412,N_8415,N_7509);
nor U10413 (N_10413,N_7123,N_7654);
and U10414 (N_10414,N_8757,N_7267);
nand U10415 (N_10415,N_8354,N_6393);
xor U10416 (N_10416,N_7934,N_7478);
nand U10417 (N_10417,N_7980,N_6298);
or U10418 (N_10418,N_7119,N_7305);
nand U10419 (N_10419,N_6617,N_6607);
nand U10420 (N_10420,N_6469,N_8804);
and U10421 (N_10421,N_8492,N_8221);
and U10422 (N_10422,N_8507,N_6869);
or U10423 (N_10423,N_8557,N_8403);
xor U10424 (N_10424,N_7755,N_7244);
nor U10425 (N_10425,N_8317,N_8115);
nand U10426 (N_10426,N_7525,N_8782);
nor U10427 (N_10427,N_8200,N_6572);
nand U10428 (N_10428,N_8686,N_9341);
nand U10429 (N_10429,N_8834,N_7372);
nor U10430 (N_10430,N_7138,N_6385);
and U10431 (N_10431,N_7285,N_8536);
or U10432 (N_10432,N_8454,N_6384);
nor U10433 (N_10433,N_9077,N_9055);
nor U10434 (N_10434,N_7191,N_9169);
and U10435 (N_10435,N_7383,N_6931);
and U10436 (N_10436,N_7495,N_9174);
or U10437 (N_10437,N_8708,N_6730);
nand U10438 (N_10438,N_7333,N_7928);
xnor U10439 (N_10439,N_9329,N_6768);
nor U10440 (N_10440,N_8175,N_8748);
nand U10441 (N_10441,N_8303,N_7275);
or U10442 (N_10442,N_6585,N_8186);
and U10443 (N_10443,N_7598,N_9265);
nor U10444 (N_10444,N_8416,N_7642);
xor U10445 (N_10445,N_6656,N_7197);
nand U10446 (N_10446,N_6250,N_8075);
or U10447 (N_10447,N_8074,N_8187);
or U10448 (N_10448,N_7505,N_8564);
xnor U10449 (N_10449,N_9346,N_9374);
nand U10450 (N_10450,N_8626,N_6380);
and U10451 (N_10451,N_8360,N_6746);
nor U10452 (N_10452,N_7768,N_8819);
or U10453 (N_10453,N_7850,N_8371);
xor U10454 (N_10454,N_6374,N_7400);
or U10455 (N_10455,N_7697,N_6667);
xor U10456 (N_10456,N_8490,N_7135);
and U10457 (N_10457,N_6285,N_7597);
or U10458 (N_10458,N_8772,N_8467);
and U10459 (N_10459,N_7369,N_7518);
or U10460 (N_10460,N_6819,N_8693);
nand U10461 (N_10461,N_9193,N_8627);
nor U10462 (N_10462,N_6313,N_8880);
and U10463 (N_10463,N_8719,N_6606);
or U10464 (N_10464,N_8456,N_7029);
or U10465 (N_10465,N_8973,N_9372);
and U10466 (N_10466,N_8554,N_7375);
or U10467 (N_10467,N_8656,N_7299);
or U10468 (N_10468,N_6914,N_8850);
or U10469 (N_10469,N_6622,N_9156);
nor U10470 (N_10470,N_6975,N_8918);
nor U10471 (N_10471,N_7767,N_8050);
nand U10472 (N_10472,N_6759,N_7608);
nor U10473 (N_10473,N_6780,N_7547);
or U10474 (N_10474,N_8291,N_8894);
and U10475 (N_10475,N_6619,N_6941);
or U10476 (N_10476,N_7109,N_7296);
nand U10477 (N_10477,N_8643,N_6956);
and U10478 (N_10478,N_6796,N_6678);
nor U10479 (N_10479,N_7940,N_7829);
nand U10480 (N_10480,N_8992,N_8176);
and U10481 (N_10481,N_7771,N_9327);
or U10482 (N_10482,N_8689,N_7684);
nor U10483 (N_10483,N_7673,N_7822);
or U10484 (N_10484,N_9227,N_9024);
or U10485 (N_10485,N_8717,N_7228);
nor U10486 (N_10486,N_8547,N_7274);
and U10487 (N_10487,N_8177,N_8730);
nand U10488 (N_10488,N_6486,N_6832);
nand U10489 (N_10489,N_8954,N_7819);
nand U10490 (N_10490,N_7279,N_6748);
nand U10491 (N_10491,N_9048,N_8201);
or U10492 (N_10492,N_6641,N_6771);
nand U10493 (N_10493,N_9371,N_6679);
xnor U10494 (N_10494,N_7010,N_7025);
xnor U10495 (N_10495,N_8313,N_8238);
and U10496 (N_10496,N_7380,N_9202);
xnor U10497 (N_10497,N_7303,N_8082);
nor U10498 (N_10498,N_6367,N_7032);
and U10499 (N_10499,N_8463,N_6421);
nand U10500 (N_10500,N_7009,N_8521);
or U10501 (N_10501,N_6455,N_9125);
and U10502 (N_10502,N_7707,N_7082);
and U10503 (N_10503,N_6783,N_7101);
nand U10504 (N_10504,N_7357,N_8855);
and U10505 (N_10505,N_6419,N_7104);
nand U10506 (N_10506,N_7841,N_7554);
nand U10507 (N_10507,N_8917,N_7572);
or U10508 (N_10508,N_8632,N_7263);
and U10509 (N_10509,N_8762,N_8482);
and U10510 (N_10510,N_7834,N_8854);
and U10511 (N_10511,N_8152,N_8372);
nor U10512 (N_10512,N_8270,N_6615);
nor U10513 (N_10513,N_8995,N_7396);
and U10514 (N_10514,N_6928,N_8023);
nor U10515 (N_10515,N_7722,N_8867);
nand U10516 (N_10516,N_6717,N_6261);
xor U10517 (N_10517,N_8726,N_9138);
and U10518 (N_10518,N_7621,N_6354);
nand U10519 (N_10519,N_8334,N_8062);
nor U10520 (N_10520,N_6726,N_7480);
nand U10521 (N_10521,N_8438,N_8103);
nor U10522 (N_10522,N_8560,N_8910);
nand U10523 (N_10523,N_8446,N_6988);
and U10524 (N_10524,N_6752,N_9313);
nand U10525 (N_10525,N_6790,N_8226);
or U10526 (N_10526,N_7202,N_6390);
and U10527 (N_10527,N_7154,N_7585);
and U10528 (N_10528,N_9314,N_6443);
or U10529 (N_10529,N_9333,N_8451);
nor U10530 (N_10530,N_6473,N_6950);
nor U10531 (N_10531,N_7188,N_9216);
or U10532 (N_10532,N_9150,N_6371);
nor U10533 (N_10533,N_8514,N_8148);
nand U10534 (N_10534,N_6604,N_7134);
and U10535 (N_10535,N_7602,N_8278);
nand U10536 (N_10536,N_9203,N_7618);
nand U10537 (N_10537,N_9023,N_6487);
nand U10538 (N_10538,N_8031,N_6653);
and U10539 (N_10539,N_7600,N_9019);
xnor U10540 (N_10540,N_7783,N_7555);
or U10541 (N_10541,N_8752,N_9283);
nor U10542 (N_10542,N_7113,N_9243);
or U10543 (N_10543,N_9039,N_8112);
nor U10544 (N_10544,N_8983,N_7432);
or U10545 (N_10545,N_8398,N_7218);
nand U10546 (N_10546,N_7586,N_9081);
nor U10547 (N_10547,N_7421,N_6307);
nor U10548 (N_10548,N_6425,N_8535);
nor U10549 (N_10549,N_7035,N_7648);
nand U10550 (N_10550,N_7409,N_7331);
nor U10551 (N_10551,N_8660,N_7173);
or U10552 (N_10552,N_6400,N_6673);
nor U10553 (N_10553,N_6942,N_9129);
nand U10554 (N_10554,N_7885,N_7399);
or U10555 (N_10555,N_7688,N_7395);
and U10556 (N_10556,N_6769,N_7749);
nor U10557 (N_10557,N_7702,N_9033);
or U10558 (N_10558,N_8077,N_8591);
nor U10559 (N_10559,N_8157,N_7325);
xor U10560 (N_10560,N_7462,N_6527);
nor U10561 (N_10561,N_7012,N_6287);
or U10562 (N_10562,N_7724,N_8086);
nand U10563 (N_10563,N_8223,N_6629);
or U10564 (N_10564,N_9112,N_7353);
nand U10565 (N_10565,N_6477,N_7438);
and U10566 (N_10566,N_7492,N_7538);
nand U10567 (N_10567,N_6575,N_9124);
and U10568 (N_10568,N_8452,N_7140);
nor U10569 (N_10569,N_7981,N_7964);
or U10570 (N_10570,N_7657,N_9004);
and U10571 (N_10571,N_8618,N_7107);
xor U10572 (N_10572,N_8049,N_8059);
xnor U10573 (N_10573,N_8885,N_9198);
nand U10574 (N_10574,N_7714,N_8014);
nand U10575 (N_10575,N_8790,N_8984);
or U10576 (N_10576,N_9178,N_7124);
or U10577 (N_10577,N_6429,N_7095);
or U10578 (N_10578,N_6301,N_8397);
or U10579 (N_10579,N_9369,N_7780);
nand U10580 (N_10580,N_9231,N_8022);
nand U10581 (N_10581,N_9360,N_6584);
nor U10582 (N_10582,N_9043,N_6662);
nor U10583 (N_10583,N_6635,N_9318);
xnor U10584 (N_10584,N_6889,N_7219);
xor U10585 (N_10585,N_7804,N_8770);
and U10586 (N_10586,N_9134,N_8349);
nand U10587 (N_10587,N_9062,N_7516);
nand U10588 (N_10588,N_6352,N_8924);
or U10589 (N_10589,N_7587,N_6550);
and U10590 (N_10590,N_8089,N_7653);
or U10591 (N_10591,N_7785,N_7408);
nor U10592 (N_10592,N_7449,N_8785);
nor U10593 (N_10593,N_8300,N_7564);
or U10594 (N_10594,N_9037,N_8085);
nand U10595 (N_10595,N_6793,N_7795);
nor U10596 (N_10596,N_7006,N_7776);
or U10597 (N_10597,N_8962,N_8952);
and U10598 (N_10598,N_8395,N_9113);
nand U10599 (N_10599,N_7165,N_8445);
nor U10600 (N_10600,N_7813,N_7861);
nand U10601 (N_10601,N_7155,N_7656);
nand U10602 (N_10602,N_7024,N_6968);
nor U10603 (N_10603,N_7297,N_8871);
nand U10604 (N_10604,N_8771,N_8335);
or U10605 (N_10605,N_6314,N_7180);
nor U10606 (N_10606,N_9015,N_8697);
nand U10607 (N_10607,N_8005,N_8743);
or U10608 (N_10608,N_8578,N_7992);
and U10609 (N_10609,N_8742,N_6934);
xor U10610 (N_10610,N_7651,N_8094);
xor U10611 (N_10611,N_7982,N_8121);
or U10612 (N_10612,N_6682,N_6300);
and U10613 (N_10613,N_7004,N_8242);
nor U10614 (N_10614,N_7435,N_7643);
nand U10615 (N_10615,N_8812,N_7631);
nor U10616 (N_10616,N_9047,N_7579);
xor U10617 (N_10617,N_7330,N_6365);
nand U10618 (N_10618,N_8565,N_7329);
or U10619 (N_10619,N_8857,N_7005);
or U10620 (N_10620,N_7589,N_8324);
nand U10621 (N_10621,N_7873,N_7358);
and U10622 (N_10622,N_8218,N_8808);
nor U10623 (N_10623,N_6890,N_6873);
or U10624 (N_10624,N_8409,N_6534);
and U10625 (N_10625,N_8675,N_8368);
or U10626 (N_10626,N_9194,N_6503);
and U10627 (N_10627,N_6983,N_7544);
or U10628 (N_10628,N_6535,N_9262);
or U10629 (N_10629,N_8642,N_6772);
nand U10630 (N_10630,N_7061,N_9132);
nor U10631 (N_10631,N_9018,N_7335);
or U10632 (N_10632,N_7351,N_6878);
nor U10633 (N_10633,N_8165,N_9098);
nand U10634 (N_10634,N_6913,N_8820);
nand U10635 (N_10635,N_8573,N_7340);
or U10636 (N_10636,N_8845,N_6498);
nor U10637 (N_10637,N_7799,N_7693);
nand U10638 (N_10638,N_7820,N_6289);
nor U10639 (N_10639,N_7416,N_6461);
nand U10640 (N_10640,N_7694,N_8934);
nand U10641 (N_10641,N_8485,N_6278);
nor U10642 (N_10642,N_8593,N_7665);
xor U10643 (N_10643,N_8638,N_7359);
nand U10644 (N_10644,N_8574,N_9254);
or U10645 (N_10645,N_6838,N_7062);
nor U10646 (N_10646,N_6306,N_6798);
nor U10647 (N_10647,N_6413,N_8982);
or U10648 (N_10648,N_6782,N_8826);
xor U10649 (N_10649,N_7726,N_7456);
or U10650 (N_10650,N_8587,N_7991);
xor U10651 (N_10651,N_8577,N_6694);
nor U10652 (N_10652,N_7272,N_7031);
nand U10653 (N_10653,N_7167,N_8150);
and U10654 (N_10654,N_9279,N_8539);
and U10655 (N_10655,N_8099,N_9078);
xnor U10656 (N_10656,N_8936,N_8651);
or U10657 (N_10657,N_7343,N_8750);
nor U10658 (N_10658,N_7308,N_6436);
or U10659 (N_10659,N_6564,N_6861);
and U10660 (N_10660,N_8464,N_8294);
and U10661 (N_10661,N_6665,N_6828);
nor U10662 (N_10662,N_6520,N_8453);
and U10663 (N_10663,N_7613,N_6457);
or U10664 (N_10664,N_8234,N_8213);
nor U10665 (N_10665,N_7341,N_8525);
xor U10666 (N_10666,N_7646,N_6879);
and U10667 (N_10667,N_8830,N_8026);
nand U10668 (N_10668,N_6423,N_8510);
or U10669 (N_10669,N_6802,N_8305);
and U10670 (N_10670,N_6852,N_8273);
nor U10671 (N_10671,N_7954,N_7431);
or U10672 (N_10672,N_6683,N_8728);
nand U10673 (N_10673,N_7125,N_6563);
or U10674 (N_10674,N_7007,N_7463);
xor U10675 (N_10675,N_9289,N_6529);
and U10676 (N_10676,N_9296,N_6397);
or U10677 (N_10677,N_8267,N_9008);
nor U10678 (N_10678,N_7652,N_6552);
or U10679 (N_10679,N_8146,N_6492);
and U10680 (N_10680,N_8949,N_8509);
or U10681 (N_10681,N_8746,N_7055);
or U10682 (N_10682,N_8630,N_8266);
nor U10683 (N_10683,N_7809,N_6389);
and U10684 (N_10684,N_7647,N_6409);
or U10685 (N_10685,N_8606,N_6493);
nand U10686 (N_10686,N_8712,N_8701);
nor U10687 (N_10687,N_8158,N_9131);
nand U10688 (N_10688,N_7675,N_6280);
nor U10689 (N_10689,N_7447,N_6319);
and U10690 (N_10690,N_7276,N_7177);
or U10691 (N_10691,N_8212,N_7145);
nor U10692 (N_10692,N_6715,N_7309);
or U10693 (N_10693,N_8106,N_7614);
or U10694 (N_10694,N_7772,N_8375);
nand U10695 (N_10695,N_6723,N_8594);
nand U10696 (N_10696,N_7938,N_8340);
nor U10697 (N_10697,N_8987,N_8940);
nor U10698 (N_10698,N_8198,N_7203);
nor U10699 (N_10699,N_7310,N_9365);
or U10700 (N_10700,N_6551,N_6904);
or U10701 (N_10701,N_6892,N_7257);
xor U10702 (N_10702,N_7851,N_9305);
and U10703 (N_10703,N_9160,N_8337);
or U10704 (N_10704,N_8622,N_8069);
nor U10705 (N_10705,N_6688,N_8301);
nand U10706 (N_10706,N_7013,N_8302);
nand U10707 (N_10707,N_7376,N_6282);
nor U10708 (N_10708,N_6356,N_6953);
nand U10709 (N_10709,N_7623,N_7280);
nor U10710 (N_10710,N_8078,N_7288);
or U10711 (N_10711,N_6708,N_7347);
and U10712 (N_10712,N_9095,N_8225);
nand U10713 (N_10713,N_7666,N_8619);
or U10714 (N_10714,N_6785,N_7472);
or U10715 (N_10715,N_8508,N_6765);
xnor U10716 (N_10716,N_8261,N_8838);
or U10717 (N_10717,N_7725,N_7893);
or U10718 (N_10718,N_7446,N_7100);
nand U10719 (N_10719,N_8549,N_7769);
and U10720 (N_10720,N_7879,N_8637);
and U10721 (N_10721,N_6440,N_7591);
or U10722 (N_10722,N_8780,N_8318);
nor U10723 (N_10723,N_6895,N_6925);
or U10724 (N_10724,N_7680,N_6974);
or U10725 (N_10725,N_7370,N_7580);
nor U10726 (N_10726,N_8046,N_7026);
nor U10727 (N_10727,N_6368,N_7300);
or U10728 (N_10728,N_7592,N_7507);
or U10729 (N_10729,N_7170,N_7152);
nor U10730 (N_10730,N_8141,N_8518);
and U10731 (N_10731,N_8475,N_8319);
nand U10732 (N_10732,N_6553,N_6971);
or U10733 (N_10733,N_8052,N_6521);
nand U10734 (N_10734,N_9029,N_7185);
or U10735 (N_10735,N_6991,N_7756);
xor U10736 (N_10736,N_8087,N_9223);
and U10737 (N_10737,N_7784,N_7008);
and U10738 (N_10738,N_6427,N_8687);
nor U10739 (N_10739,N_7550,N_6990);
xnor U10740 (N_10740,N_9237,N_7192);
and U10741 (N_10741,N_9338,N_8209);
and U10742 (N_10742,N_9205,N_7593);
nor U10743 (N_10743,N_9101,N_7698);
nor U10744 (N_10744,N_8323,N_7126);
and U10745 (N_10745,N_7136,N_7290);
nor U10746 (N_10746,N_8420,N_9100);
or U10747 (N_10747,N_8505,N_7163);
and U10748 (N_10748,N_7506,N_7578);
and U10749 (N_10749,N_6569,N_8906);
and U10750 (N_10750,N_9083,N_6505);
nand U10751 (N_10751,N_8835,N_6589);
or U10752 (N_10752,N_7441,N_7066);
nand U10753 (N_10753,N_7193,N_7536);
nand U10754 (N_10754,N_7078,N_6725);
nor U10755 (N_10755,N_7967,N_7350);
and U10756 (N_10756,N_7392,N_8802);
and U10757 (N_10757,N_8236,N_8222);
xor U10758 (N_10758,N_6281,N_8120);
and U10759 (N_10759,N_8339,N_8598);
nand U10760 (N_10760,N_6403,N_8322);
and U10761 (N_10761,N_7390,N_8441);
nor U10762 (N_10762,N_9328,N_7512);
xor U10763 (N_10763,N_7318,N_6886);
nand U10764 (N_10764,N_6817,N_7364);
nand U10765 (N_10765,N_6937,N_8747);
and U10766 (N_10766,N_6592,N_8975);
nor U10767 (N_10767,N_7161,N_9030);
and U10768 (N_10768,N_9007,N_8738);
or U10769 (N_10769,N_7689,N_9111);
nor U10770 (N_10770,N_8881,N_9246);
and U10771 (N_10771,N_7626,N_8290);
or U10772 (N_10772,N_7661,N_6812);
nand U10773 (N_10773,N_8609,N_6871);
nand U10774 (N_10774,N_7042,N_7559);
nor U10775 (N_10775,N_7382,N_7142);
or U10776 (N_10776,N_9148,N_7000);
nor U10777 (N_10777,N_7823,N_7649);
or U10778 (N_10778,N_9141,N_7937);
and U10779 (N_10779,N_6762,N_8753);
or U10780 (N_10780,N_7782,N_8608);
nor U10781 (N_10781,N_6677,N_6540);
nand U10782 (N_10782,N_8533,N_6559);
nand U10783 (N_10783,N_7023,N_8113);
nand U10784 (N_10784,N_7071,N_8006);
and U10785 (N_10785,N_7909,N_7667);
or U10786 (N_10786,N_7051,N_6386);
or U10787 (N_10787,N_8615,N_6317);
nor U10788 (N_10788,N_7715,N_7070);
nand U10789 (N_10789,N_8020,N_8700);
or U10790 (N_10790,N_7947,N_8067);
nand U10791 (N_10791,N_8233,N_9257);
nand U10792 (N_10792,N_7482,N_6911);
and U10793 (N_10793,N_7976,N_6840);
or U10794 (N_10794,N_6355,N_8496);
or U10795 (N_10795,N_9003,N_9208);
nand U10796 (N_10796,N_6767,N_6418);
and U10797 (N_10797,N_7910,N_7503);
nor U10798 (N_10798,N_9232,N_8903);
nor U10799 (N_10799,N_7150,N_6468);
and U10800 (N_10800,N_7770,N_9344);
nor U10801 (N_10801,N_8003,N_7332);
nor U10802 (N_10802,N_8056,N_8260);
and U10803 (N_10803,N_8625,N_8088);
nand U10804 (N_10804,N_9311,N_9273);
nand U10805 (N_10805,N_8096,N_7919);
nor U10806 (N_10806,N_7635,N_7558);
nor U10807 (N_10807,N_8895,N_9011);
nor U10808 (N_10808,N_7527,N_8380);
or U10809 (N_10809,N_9087,N_8174);
nor U10810 (N_10810,N_6286,N_7484);
nand U10811 (N_10811,N_7293,N_8437);
nor U10812 (N_10812,N_6938,N_7788);
xor U10813 (N_10813,N_9162,N_9016);
and U10814 (N_10814,N_6734,N_7884);
nand U10815 (N_10815,N_8306,N_7242);
or U10816 (N_10816,N_8487,N_8824);
or U10817 (N_10817,N_6738,N_7999);
and U10818 (N_10818,N_7141,N_6379);
and U10819 (N_10819,N_8532,N_8439);
or U10820 (N_10820,N_8247,N_6377);
nor U10821 (N_10821,N_8224,N_8636);
or U10822 (N_10822,N_8766,N_8938);
and U10823 (N_10823,N_8621,N_9200);
xor U10824 (N_10824,N_8629,N_8958);
xnor U10825 (N_10825,N_8709,N_6648);
nor U10826 (N_10826,N_7483,N_6792);
nand U10827 (N_10827,N_6639,N_6411);
nor U10828 (N_10828,N_8364,N_7151);
nor U10829 (N_10829,N_8597,N_7607);
nand U10830 (N_10830,N_7094,N_7699);
nand U10831 (N_10831,N_8641,N_7814);
nand U10832 (N_10832,N_8776,N_7037);
and U10833 (N_10833,N_6624,N_8640);
xnor U10834 (N_10834,N_8053,N_7429);
nand U10835 (N_10835,N_7337,N_6858);
or U10836 (N_10836,N_7629,N_8990);
xnor U10837 (N_10837,N_6577,N_7549);
or U10838 (N_10838,N_7609,N_9278);
nor U10839 (N_10839,N_8904,N_6322);
and U10840 (N_10840,N_6719,N_6264);
nand U10841 (N_10841,N_7458,N_6700);
and U10842 (N_10842,N_7259,N_8283);
or U10843 (N_10843,N_6587,N_9221);
and U10844 (N_10844,N_6885,N_6514);
and U10845 (N_10845,N_9167,N_7571);
xnor U10846 (N_10846,N_8251,N_9028);
nand U10847 (N_10847,N_8073,N_9106);
xnor U10848 (N_10848,N_6364,N_6395);
or U10849 (N_10849,N_6702,N_8178);
or U10850 (N_10850,N_8426,N_8913);
or U10851 (N_10851,N_8289,N_7896);
xor U10852 (N_10852,N_7865,N_8167);
nor U10853 (N_10853,N_8101,N_8489);
and U10854 (N_10854,N_7985,N_9256);
nand U10855 (N_10855,N_7053,N_9026);
xor U10856 (N_10856,N_7798,N_6967);
nor U10857 (N_10857,N_8252,N_6509);
and U10858 (N_10858,N_7086,N_7494);
nand U10859 (N_10859,N_8070,N_6982);
and U10860 (N_10860,N_8511,N_7570);
xnor U10861 (N_10861,N_7436,N_8443);
and U10862 (N_10862,N_7977,N_7475);
or U10863 (N_10863,N_7727,N_9301);
or U10864 (N_10864,N_8258,N_7624);
or U10865 (N_10865,N_8928,N_7892);
and U10866 (N_10866,N_9102,N_6644);
nand U10867 (N_10867,N_8502,N_8472);
nor U10868 (N_10868,N_8208,N_9175);
or U10869 (N_10869,N_6612,N_6449);
and U10870 (N_10870,N_8051,N_7489);
or U10871 (N_10871,N_8116,N_6504);
nor U10872 (N_10872,N_8118,N_6391);
or U10873 (N_10873,N_9320,N_9063);
and U10874 (N_10874,N_6638,N_9358);
and U10875 (N_10875,N_8613,N_9181);
nand U10876 (N_10876,N_6297,N_7918);
nor U10877 (N_10877,N_6453,N_7939);
nor U10878 (N_10878,N_8550,N_6658);
xor U10879 (N_10879,N_9361,N_6618);
and U10880 (N_10880,N_6580,N_7759);
or U10881 (N_10881,N_7864,N_8647);
xor U10882 (N_10882,N_8758,N_9068);
nor U10883 (N_10883,N_8744,N_7423);
and U10884 (N_10884,N_9310,N_8862);
or U10885 (N_10885,N_7500,N_6262);
or U10886 (N_10886,N_6318,N_7709);
xnor U10887 (N_10887,N_8203,N_8976);
nor U10888 (N_10888,N_6333,N_7099);
nand U10889 (N_10889,N_8569,N_8035);
or U10890 (N_10890,N_7658,N_8329);
and U10891 (N_10891,N_6915,N_8769);
or U10892 (N_10892,N_7045,N_9094);
nand U10893 (N_10893,N_7906,N_6939);
or U10894 (N_10894,N_7385,N_7911);
and U10895 (N_10895,N_8529,N_7253);
and U10896 (N_10896,N_6435,N_9058);
and U10897 (N_10897,N_7189,N_8794);
nor U10898 (N_10898,N_6805,N_9286);
or U10899 (N_10899,N_9293,N_6331);
xor U10900 (N_10900,N_7215,N_8884);
or U10901 (N_10901,N_7914,N_6998);
or U10902 (N_10902,N_6481,N_6548);
and U10903 (N_10903,N_8219,N_7129);
nand U10904 (N_10904,N_7291,N_8644);
or U10905 (N_10905,N_7760,N_7556);
nand U10906 (N_10906,N_8248,N_8084);
nor U10907 (N_10907,N_8891,N_6546);
and U10908 (N_10908,N_9319,N_7826);
xnor U10909 (N_10909,N_6299,N_7065);
or U10910 (N_10910,N_9066,N_9107);
nor U10911 (N_10911,N_6703,N_8759);
nand U10912 (N_10912,N_8277,N_7501);
xnor U10913 (N_10913,N_7754,N_7716);
nand U10914 (N_10914,N_8883,N_6544);
nor U10915 (N_10915,N_6482,N_6290);
and U10916 (N_10916,N_8138,N_7440);
or U10917 (N_10917,N_8000,N_8351);
nor U10918 (N_10918,N_6749,N_8353);
and U10919 (N_10919,N_7540,N_9052);
and U10920 (N_10920,N_8833,N_9306);
or U10921 (N_10921,N_7361,N_6430);
nand U10922 (N_10922,N_9097,N_8296);
or U10923 (N_10923,N_7723,N_6543);
xor U10924 (N_10924,N_6294,N_9144);
and U10925 (N_10925,N_7174,N_7764);
nor U10926 (N_10926,N_8925,N_6608);
and U10927 (N_10927,N_6337,N_7312);
or U10928 (N_10928,N_6714,N_8377);
nor U10929 (N_10929,N_7827,N_9356);
nor U10930 (N_10930,N_6533,N_8969);
or U10931 (N_10931,N_8192,N_7511);
and U10932 (N_10932,N_8648,N_6720);
nor U10933 (N_10933,N_9189,N_7224);
and U10934 (N_10934,N_8943,N_7691);
or U10935 (N_10935,N_8781,N_7388);
nor U10936 (N_10936,N_6346,N_8599);
nor U10937 (N_10937,N_8725,N_9161);
nor U10938 (N_10938,N_6955,N_6824);
nor U10939 (N_10939,N_7331,N_7226);
or U10940 (N_10940,N_8678,N_7894);
or U10941 (N_10941,N_7802,N_9102);
nand U10942 (N_10942,N_7174,N_8889);
nand U10943 (N_10943,N_8008,N_6422);
nor U10944 (N_10944,N_6886,N_6674);
or U10945 (N_10945,N_7782,N_8903);
and U10946 (N_10946,N_9330,N_7046);
and U10947 (N_10947,N_6981,N_6676);
nand U10948 (N_10948,N_9162,N_7431);
nand U10949 (N_10949,N_6479,N_6320);
and U10950 (N_10950,N_6587,N_7085);
or U10951 (N_10951,N_8145,N_6976);
nand U10952 (N_10952,N_6760,N_8134);
xnor U10953 (N_10953,N_6389,N_7556);
nor U10954 (N_10954,N_8868,N_9224);
and U10955 (N_10955,N_6517,N_7883);
and U10956 (N_10956,N_6693,N_8291);
nand U10957 (N_10957,N_6322,N_6895);
nand U10958 (N_10958,N_8242,N_8470);
and U10959 (N_10959,N_7335,N_8337);
or U10960 (N_10960,N_9372,N_6349);
nand U10961 (N_10961,N_8463,N_8722);
or U10962 (N_10962,N_9351,N_8270);
and U10963 (N_10963,N_8641,N_7955);
nand U10964 (N_10964,N_6827,N_6651);
and U10965 (N_10965,N_9119,N_6725);
or U10966 (N_10966,N_7261,N_8654);
and U10967 (N_10967,N_9338,N_9036);
or U10968 (N_10968,N_8692,N_9084);
or U10969 (N_10969,N_6650,N_9155);
nand U10970 (N_10970,N_8120,N_7310);
nor U10971 (N_10971,N_6496,N_7204);
and U10972 (N_10972,N_9042,N_8447);
or U10973 (N_10973,N_8205,N_8312);
nand U10974 (N_10974,N_9067,N_8924);
or U10975 (N_10975,N_8546,N_7093);
or U10976 (N_10976,N_7505,N_6414);
and U10977 (N_10977,N_8470,N_9073);
or U10978 (N_10978,N_8753,N_8417);
nor U10979 (N_10979,N_8255,N_7660);
nor U10980 (N_10980,N_8860,N_8361);
nor U10981 (N_10981,N_7440,N_7642);
or U10982 (N_10982,N_6647,N_6723);
or U10983 (N_10983,N_7704,N_6373);
nand U10984 (N_10984,N_8138,N_7969);
nand U10985 (N_10985,N_7620,N_9077);
and U10986 (N_10986,N_6956,N_9114);
or U10987 (N_10987,N_6985,N_6745);
and U10988 (N_10988,N_7663,N_8295);
xnor U10989 (N_10989,N_7987,N_6511);
and U10990 (N_10990,N_7159,N_7646);
or U10991 (N_10991,N_9277,N_9003);
and U10992 (N_10992,N_8472,N_8246);
and U10993 (N_10993,N_9048,N_7636);
and U10994 (N_10994,N_8300,N_6777);
and U10995 (N_10995,N_6469,N_6672);
nand U10996 (N_10996,N_8629,N_8252);
and U10997 (N_10997,N_9200,N_7063);
or U10998 (N_10998,N_6556,N_9009);
and U10999 (N_10999,N_6318,N_8821);
nand U11000 (N_11000,N_8036,N_7399);
and U11001 (N_11001,N_6326,N_8807);
nand U11002 (N_11002,N_8193,N_6851);
nor U11003 (N_11003,N_8716,N_6896);
nand U11004 (N_11004,N_8304,N_8464);
nand U11005 (N_11005,N_8766,N_7588);
and U11006 (N_11006,N_6544,N_6372);
nand U11007 (N_11007,N_7438,N_9317);
nand U11008 (N_11008,N_7473,N_7764);
and U11009 (N_11009,N_7863,N_7850);
nand U11010 (N_11010,N_8826,N_6542);
or U11011 (N_11011,N_9115,N_7540);
nor U11012 (N_11012,N_7933,N_8880);
nand U11013 (N_11013,N_8625,N_6442);
or U11014 (N_11014,N_6844,N_7350);
or U11015 (N_11015,N_6937,N_8440);
nor U11016 (N_11016,N_8223,N_6558);
nor U11017 (N_11017,N_6686,N_7881);
nor U11018 (N_11018,N_8784,N_8341);
nor U11019 (N_11019,N_6687,N_7657);
nand U11020 (N_11020,N_7917,N_9191);
and U11021 (N_11021,N_9334,N_6798);
and U11022 (N_11022,N_8731,N_9148);
nor U11023 (N_11023,N_8867,N_7211);
or U11024 (N_11024,N_9156,N_8451);
nand U11025 (N_11025,N_9155,N_7921);
and U11026 (N_11026,N_6290,N_8442);
nor U11027 (N_11027,N_8634,N_6519);
nor U11028 (N_11028,N_9024,N_9094);
nor U11029 (N_11029,N_8167,N_8817);
and U11030 (N_11030,N_7670,N_6401);
nor U11031 (N_11031,N_8939,N_8129);
nor U11032 (N_11032,N_7188,N_7180);
nor U11033 (N_11033,N_8448,N_9241);
or U11034 (N_11034,N_8373,N_6971);
or U11035 (N_11035,N_7224,N_9314);
nor U11036 (N_11036,N_7656,N_6447);
nor U11037 (N_11037,N_9365,N_8994);
xor U11038 (N_11038,N_7138,N_8372);
xnor U11039 (N_11039,N_9101,N_7237);
nand U11040 (N_11040,N_8741,N_7567);
nor U11041 (N_11041,N_8665,N_7299);
xor U11042 (N_11042,N_9141,N_6849);
and U11043 (N_11043,N_6355,N_7197);
or U11044 (N_11044,N_8777,N_9271);
nor U11045 (N_11045,N_7871,N_6623);
nor U11046 (N_11046,N_7271,N_7034);
nand U11047 (N_11047,N_7136,N_8009);
nand U11048 (N_11048,N_7269,N_6571);
nand U11049 (N_11049,N_8086,N_8090);
nand U11050 (N_11050,N_7293,N_8688);
nor U11051 (N_11051,N_6692,N_8578);
and U11052 (N_11052,N_8967,N_9057);
and U11053 (N_11053,N_7608,N_7802);
xnor U11054 (N_11054,N_7885,N_6984);
or U11055 (N_11055,N_6432,N_8984);
and U11056 (N_11056,N_6579,N_6348);
or U11057 (N_11057,N_7474,N_7494);
and U11058 (N_11058,N_8242,N_9282);
and U11059 (N_11059,N_9053,N_9220);
or U11060 (N_11060,N_7288,N_8848);
nor U11061 (N_11061,N_7749,N_8462);
nand U11062 (N_11062,N_8597,N_6745);
and U11063 (N_11063,N_8081,N_7514);
nand U11064 (N_11064,N_7385,N_8160);
or U11065 (N_11065,N_8823,N_7458);
or U11066 (N_11066,N_8806,N_6806);
xnor U11067 (N_11067,N_7515,N_6881);
nand U11068 (N_11068,N_9177,N_8604);
nor U11069 (N_11069,N_6557,N_8646);
and U11070 (N_11070,N_8911,N_7088);
or U11071 (N_11071,N_8041,N_9206);
and U11072 (N_11072,N_8799,N_7437);
nor U11073 (N_11073,N_8731,N_7203);
and U11074 (N_11074,N_9005,N_7384);
nand U11075 (N_11075,N_7552,N_7193);
or U11076 (N_11076,N_9327,N_9119);
nand U11077 (N_11077,N_9267,N_7805);
nor U11078 (N_11078,N_8932,N_7051);
or U11079 (N_11079,N_7575,N_6525);
nor U11080 (N_11080,N_6793,N_6452);
or U11081 (N_11081,N_7661,N_8937);
nand U11082 (N_11082,N_6864,N_8067);
xnor U11083 (N_11083,N_7282,N_8365);
nand U11084 (N_11084,N_7525,N_7164);
nor U11085 (N_11085,N_7689,N_7305);
nor U11086 (N_11086,N_6960,N_9178);
nand U11087 (N_11087,N_7608,N_9316);
and U11088 (N_11088,N_6867,N_6798);
or U11089 (N_11089,N_8250,N_8892);
nand U11090 (N_11090,N_6390,N_6380);
and U11091 (N_11091,N_6268,N_7805);
nor U11092 (N_11092,N_9079,N_6547);
nand U11093 (N_11093,N_6251,N_7534);
and U11094 (N_11094,N_7450,N_8930);
xor U11095 (N_11095,N_8223,N_6408);
or U11096 (N_11096,N_6426,N_6855);
or U11097 (N_11097,N_9114,N_9207);
nand U11098 (N_11098,N_7326,N_7086);
nand U11099 (N_11099,N_6767,N_8644);
nand U11100 (N_11100,N_8563,N_8594);
and U11101 (N_11101,N_8596,N_6872);
nor U11102 (N_11102,N_6752,N_8729);
or U11103 (N_11103,N_8670,N_6714);
or U11104 (N_11104,N_7379,N_6650);
nand U11105 (N_11105,N_8609,N_6374);
and U11106 (N_11106,N_9031,N_6507);
and U11107 (N_11107,N_7231,N_6680);
xnor U11108 (N_11108,N_6848,N_7700);
or U11109 (N_11109,N_8114,N_8974);
nor U11110 (N_11110,N_9129,N_8577);
and U11111 (N_11111,N_9297,N_6441);
nand U11112 (N_11112,N_7289,N_8759);
or U11113 (N_11113,N_9107,N_8738);
xnor U11114 (N_11114,N_7264,N_9321);
nor U11115 (N_11115,N_8270,N_7485);
and U11116 (N_11116,N_7605,N_8142);
and U11117 (N_11117,N_9081,N_9282);
nand U11118 (N_11118,N_7649,N_8742);
and U11119 (N_11119,N_8867,N_8172);
and U11120 (N_11120,N_6340,N_6487);
and U11121 (N_11121,N_8726,N_8763);
and U11122 (N_11122,N_6514,N_6580);
or U11123 (N_11123,N_8907,N_7189);
nor U11124 (N_11124,N_8921,N_8654);
or U11125 (N_11125,N_6407,N_6356);
nor U11126 (N_11126,N_7217,N_6727);
or U11127 (N_11127,N_6495,N_8367);
xor U11128 (N_11128,N_7984,N_7763);
or U11129 (N_11129,N_8442,N_7253);
nand U11130 (N_11130,N_8525,N_7237);
nor U11131 (N_11131,N_8394,N_8273);
nand U11132 (N_11132,N_6911,N_6955);
or U11133 (N_11133,N_8098,N_7421);
or U11134 (N_11134,N_7333,N_9350);
nand U11135 (N_11135,N_8198,N_6405);
nand U11136 (N_11136,N_9178,N_7615);
nor U11137 (N_11137,N_6367,N_8707);
and U11138 (N_11138,N_9098,N_8562);
xnor U11139 (N_11139,N_7246,N_7804);
and U11140 (N_11140,N_8589,N_8368);
and U11141 (N_11141,N_7833,N_7947);
xor U11142 (N_11142,N_8215,N_8709);
nor U11143 (N_11143,N_7200,N_7214);
nor U11144 (N_11144,N_8191,N_6942);
or U11145 (N_11145,N_7370,N_7723);
nor U11146 (N_11146,N_8118,N_9048);
or U11147 (N_11147,N_8332,N_8745);
and U11148 (N_11148,N_6328,N_6912);
or U11149 (N_11149,N_6849,N_6592);
nand U11150 (N_11150,N_9067,N_7909);
or U11151 (N_11151,N_7817,N_8547);
and U11152 (N_11152,N_7288,N_7971);
and U11153 (N_11153,N_7916,N_6759);
or U11154 (N_11154,N_8674,N_7087);
and U11155 (N_11155,N_7365,N_9298);
nor U11156 (N_11156,N_7877,N_7329);
or U11157 (N_11157,N_7426,N_8959);
and U11158 (N_11158,N_7490,N_6270);
and U11159 (N_11159,N_7978,N_7742);
xor U11160 (N_11160,N_6481,N_7375);
or U11161 (N_11161,N_8260,N_8457);
and U11162 (N_11162,N_8729,N_6950);
and U11163 (N_11163,N_6664,N_7760);
nand U11164 (N_11164,N_7152,N_6820);
nor U11165 (N_11165,N_8420,N_8107);
and U11166 (N_11166,N_7872,N_7842);
and U11167 (N_11167,N_7991,N_8927);
and U11168 (N_11168,N_9288,N_8724);
nor U11169 (N_11169,N_6330,N_8634);
nor U11170 (N_11170,N_8336,N_7890);
and U11171 (N_11171,N_9246,N_7344);
and U11172 (N_11172,N_6400,N_7435);
nand U11173 (N_11173,N_7504,N_8347);
and U11174 (N_11174,N_7701,N_9146);
nand U11175 (N_11175,N_8468,N_7854);
and U11176 (N_11176,N_8600,N_8247);
nand U11177 (N_11177,N_7961,N_8734);
or U11178 (N_11178,N_7057,N_7784);
or U11179 (N_11179,N_9147,N_7227);
nand U11180 (N_11180,N_7686,N_7627);
or U11181 (N_11181,N_7786,N_9280);
or U11182 (N_11182,N_6252,N_7496);
and U11183 (N_11183,N_9168,N_8926);
and U11184 (N_11184,N_7107,N_8078);
nor U11185 (N_11185,N_9227,N_6552);
or U11186 (N_11186,N_8769,N_8042);
nand U11187 (N_11187,N_6517,N_6444);
or U11188 (N_11188,N_6781,N_7023);
nor U11189 (N_11189,N_8833,N_8727);
nor U11190 (N_11190,N_6453,N_9035);
and U11191 (N_11191,N_7111,N_7764);
nor U11192 (N_11192,N_9066,N_6688);
or U11193 (N_11193,N_8818,N_7939);
or U11194 (N_11194,N_8632,N_7109);
nand U11195 (N_11195,N_6514,N_8602);
nand U11196 (N_11196,N_6768,N_8701);
and U11197 (N_11197,N_7572,N_8391);
or U11198 (N_11198,N_8998,N_6314);
or U11199 (N_11199,N_6927,N_8677);
and U11200 (N_11200,N_8617,N_8818);
nand U11201 (N_11201,N_8223,N_8023);
and U11202 (N_11202,N_8393,N_6273);
nand U11203 (N_11203,N_8599,N_6592);
and U11204 (N_11204,N_6980,N_6853);
nand U11205 (N_11205,N_8965,N_8069);
and U11206 (N_11206,N_7433,N_7148);
nor U11207 (N_11207,N_6539,N_7534);
and U11208 (N_11208,N_8619,N_6444);
nand U11209 (N_11209,N_6966,N_7375);
nor U11210 (N_11210,N_8026,N_6979);
nor U11211 (N_11211,N_9085,N_8154);
and U11212 (N_11212,N_8974,N_8078);
nand U11213 (N_11213,N_7234,N_8120);
or U11214 (N_11214,N_7405,N_9254);
or U11215 (N_11215,N_8449,N_6657);
nor U11216 (N_11216,N_6507,N_8748);
and U11217 (N_11217,N_8781,N_8244);
nand U11218 (N_11218,N_7443,N_6811);
and U11219 (N_11219,N_6853,N_7093);
xnor U11220 (N_11220,N_6275,N_7750);
or U11221 (N_11221,N_8168,N_7702);
nor U11222 (N_11222,N_8920,N_9250);
and U11223 (N_11223,N_7717,N_7323);
and U11224 (N_11224,N_6419,N_8848);
xor U11225 (N_11225,N_8349,N_7382);
and U11226 (N_11226,N_7440,N_8103);
and U11227 (N_11227,N_9313,N_7978);
nand U11228 (N_11228,N_6819,N_6255);
or U11229 (N_11229,N_8620,N_7214);
and U11230 (N_11230,N_8749,N_8194);
or U11231 (N_11231,N_8776,N_8567);
nand U11232 (N_11232,N_7517,N_7964);
nor U11233 (N_11233,N_6580,N_7398);
and U11234 (N_11234,N_7620,N_8967);
or U11235 (N_11235,N_7371,N_9255);
nand U11236 (N_11236,N_7055,N_6936);
and U11237 (N_11237,N_7652,N_7230);
or U11238 (N_11238,N_7044,N_7434);
nor U11239 (N_11239,N_8836,N_8706);
or U11240 (N_11240,N_9353,N_9106);
xor U11241 (N_11241,N_6664,N_6405);
nor U11242 (N_11242,N_6835,N_7425);
nand U11243 (N_11243,N_9267,N_8871);
and U11244 (N_11244,N_7776,N_6971);
or U11245 (N_11245,N_8285,N_8811);
nand U11246 (N_11246,N_8044,N_6749);
nor U11247 (N_11247,N_6516,N_9105);
nor U11248 (N_11248,N_7319,N_8693);
nor U11249 (N_11249,N_7567,N_7926);
and U11250 (N_11250,N_6306,N_7130);
nand U11251 (N_11251,N_6378,N_7359);
and U11252 (N_11252,N_8777,N_6275);
xnor U11253 (N_11253,N_9250,N_9142);
nor U11254 (N_11254,N_9373,N_7185);
nor U11255 (N_11255,N_8449,N_8520);
nand U11256 (N_11256,N_8752,N_8912);
nand U11257 (N_11257,N_9137,N_9369);
and U11258 (N_11258,N_7768,N_7496);
or U11259 (N_11259,N_8748,N_8957);
nor U11260 (N_11260,N_8852,N_8134);
nand U11261 (N_11261,N_8269,N_8604);
and U11262 (N_11262,N_6864,N_7852);
or U11263 (N_11263,N_6552,N_9088);
nor U11264 (N_11264,N_8528,N_6357);
nand U11265 (N_11265,N_7152,N_6807);
and U11266 (N_11266,N_7850,N_7529);
nand U11267 (N_11267,N_7107,N_7791);
nor U11268 (N_11268,N_8849,N_6988);
nor U11269 (N_11269,N_9346,N_6967);
or U11270 (N_11270,N_6472,N_7736);
and U11271 (N_11271,N_8907,N_7912);
xor U11272 (N_11272,N_8192,N_7954);
or U11273 (N_11273,N_8382,N_6858);
xor U11274 (N_11274,N_8165,N_7681);
nor U11275 (N_11275,N_7908,N_7543);
nor U11276 (N_11276,N_8331,N_9170);
nand U11277 (N_11277,N_8869,N_7987);
xnor U11278 (N_11278,N_8632,N_8877);
nand U11279 (N_11279,N_7593,N_8258);
nand U11280 (N_11280,N_7374,N_8851);
nand U11281 (N_11281,N_7606,N_7711);
nor U11282 (N_11282,N_6674,N_8175);
xnor U11283 (N_11283,N_9138,N_9167);
or U11284 (N_11284,N_7053,N_7218);
and U11285 (N_11285,N_7444,N_8790);
nand U11286 (N_11286,N_8298,N_7241);
xor U11287 (N_11287,N_7395,N_8786);
nor U11288 (N_11288,N_7652,N_8402);
xor U11289 (N_11289,N_9097,N_9052);
nand U11290 (N_11290,N_9325,N_7872);
or U11291 (N_11291,N_6889,N_6798);
or U11292 (N_11292,N_6910,N_7085);
and U11293 (N_11293,N_7316,N_8060);
or U11294 (N_11294,N_8365,N_6312);
nand U11295 (N_11295,N_9176,N_8545);
nor U11296 (N_11296,N_9171,N_8540);
nor U11297 (N_11297,N_6541,N_8651);
and U11298 (N_11298,N_9110,N_6956);
or U11299 (N_11299,N_8705,N_6366);
nand U11300 (N_11300,N_6322,N_7455);
nand U11301 (N_11301,N_7870,N_6803);
and U11302 (N_11302,N_7564,N_7714);
nand U11303 (N_11303,N_6672,N_7284);
nor U11304 (N_11304,N_7066,N_6727);
nor U11305 (N_11305,N_8900,N_9213);
and U11306 (N_11306,N_6353,N_8440);
nor U11307 (N_11307,N_7801,N_8902);
or U11308 (N_11308,N_8484,N_6700);
nand U11309 (N_11309,N_7657,N_8816);
and U11310 (N_11310,N_6851,N_7799);
xor U11311 (N_11311,N_7317,N_7642);
nor U11312 (N_11312,N_9086,N_6500);
and U11313 (N_11313,N_8668,N_8433);
nand U11314 (N_11314,N_7747,N_7948);
and U11315 (N_11315,N_7723,N_8129);
nor U11316 (N_11316,N_7779,N_9197);
nand U11317 (N_11317,N_6756,N_8927);
or U11318 (N_11318,N_9014,N_9194);
or U11319 (N_11319,N_9367,N_6779);
nor U11320 (N_11320,N_6262,N_7644);
nor U11321 (N_11321,N_6265,N_7645);
nor U11322 (N_11322,N_8666,N_8317);
or U11323 (N_11323,N_9266,N_6863);
nand U11324 (N_11324,N_8081,N_7865);
or U11325 (N_11325,N_7665,N_8556);
nand U11326 (N_11326,N_6678,N_8468);
nand U11327 (N_11327,N_7648,N_6919);
or U11328 (N_11328,N_9365,N_8753);
and U11329 (N_11329,N_6358,N_9005);
nor U11330 (N_11330,N_8669,N_7654);
and U11331 (N_11331,N_8619,N_8603);
nor U11332 (N_11332,N_7919,N_6328);
nand U11333 (N_11333,N_8501,N_7220);
xnor U11334 (N_11334,N_7405,N_9093);
nand U11335 (N_11335,N_6724,N_7307);
and U11336 (N_11336,N_8273,N_8321);
or U11337 (N_11337,N_8766,N_9046);
and U11338 (N_11338,N_9127,N_7485);
nor U11339 (N_11339,N_9031,N_7736);
xnor U11340 (N_11340,N_8313,N_8427);
nand U11341 (N_11341,N_7978,N_8744);
or U11342 (N_11342,N_8228,N_7582);
nor U11343 (N_11343,N_8405,N_9200);
or U11344 (N_11344,N_9032,N_6803);
or U11345 (N_11345,N_8458,N_6600);
and U11346 (N_11346,N_8866,N_6434);
nand U11347 (N_11347,N_6560,N_8566);
nand U11348 (N_11348,N_8439,N_6548);
nor U11349 (N_11349,N_7869,N_7322);
or U11350 (N_11350,N_8686,N_6535);
xnor U11351 (N_11351,N_9290,N_7821);
nor U11352 (N_11352,N_8200,N_8909);
nand U11353 (N_11353,N_7274,N_7340);
or U11354 (N_11354,N_6536,N_8026);
nand U11355 (N_11355,N_8971,N_7739);
nand U11356 (N_11356,N_7325,N_8685);
and U11357 (N_11357,N_6988,N_6283);
and U11358 (N_11358,N_6408,N_7743);
and U11359 (N_11359,N_8428,N_8842);
nor U11360 (N_11360,N_6564,N_7862);
or U11361 (N_11361,N_7922,N_8515);
xor U11362 (N_11362,N_7149,N_6673);
xor U11363 (N_11363,N_8103,N_8339);
and U11364 (N_11364,N_7165,N_8723);
or U11365 (N_11365,N_7970,N_9217);
nor U11366 (N_11366,N_7955,N_7649);
or U11367 (N_11367,N_6605,N_9029);
and U11368 (N_11368,N_8594,N_7424);
and U11369 (N_11369,N_6978,N_9123);
nor U11370 (N_11370,N_9092,N_8314);
xnor U11371 (N_11371,N_8973,N_8678);
xor U11372 (N_11372,N_6683,N_6845);
or U11373 (N_11373,N_6610,N_8423);
nor U11374 (N_11374,N_6476,N_7382);
and U11375 (N_11375,N_6269,N_7745);
nor U11376 (N_11376,N_9186,N_6828);
or U11377 (N_11377,N_9324,N_9315);
and U11378 (N_11378,N_6367,N_6651);
nor U11379 (N_11379,N_8420,N_7924);
xor U11380 (N_11380,N_7372,N_7378);
and U11381 (N_11381,N_6907,N_8915);
nand U11382 (N_11382,N_7977,N_7612);
or U11383 (N_11383,N_7095,N_7294);
nand U11384 (N_11384,N_6636,N_7863);
nor U11385 (N_11385,N_6668,N_8773);
and U11386 (N_11386,N_7763,N_8907);
and U11387 (N_11387,N_9170,N_6409);
xnor U11388 (N_11388,N_6565,N_9262);
and U11389 (N_11389,N_7523,N_7380);
nor U11390 (N_11390,N_8720,N_9085);
nand U11391 (N_11391,N_6455,N_6614);
or U11392 (N_11392,N_8673,N_6742);
and U11393 (N_11393,N_7791,N_8196);
or U11394 (N_11394,N_7687,N_9230);
or U11395 (N_11395,N_7048,N_6512);
and U11396 (N_11396,N_7492,N_8480);
nand U11397 (N_11397,N_8178,N_7123);
or U11398 (N_11398,N_8165,N_6529);
and U11399 (N_11399,N_6541,N_6796);
xor U11400 (N_11400,N_8750,N_7793);
or U11401 (N_11401,N_8128,N_6522);
nand U11402 (N_11402,N_7415,N_6489);
and U11403 (N_11403,N_9216,N_6635);
or U11404 (N_11404,N_9250,N_9330);
and U11405 (N_11405,N_8317,N_6598);
nor U11406 (N_11406,N_7349,N_9048);
or U11407 (N_11407,N_7337,N_7087);
nor U11408 (N_11408,N_6562,N_7397);
nor U11409 (N_11409,N_8345,N_6284);
and U11410 (N_11410,N_6308,N_7840);
nand U11411 (N_11411,N_9163,N_9018);
and U11412 (N_11412,N_7010,N_7568);
nor U11413 (N_11413,N_9201,N_7069);
nand U11414 (N_11414,N_7339,N_6648);
and U11415 (N_11415,N_8970,N_6336);
nand U11416 (N_11416,N_7695,N_8165);
and U11417 (N_11417,N_8707,N_7384);
or U11418 (N_11418,N_6941,N_8227);
or U11419 (N_11419,N_8956,N_7571);
xnor U11420 (N_11420,N_6373,N_6743);
or U11421 (N_11421,N_6902,N_6377);
nor U11422 (N_11422,N_8529,N_7883);
xnor U11423 (N_11423,N_9168,N_6886);
nor U11424 (N_11424,N_8072,N_8526);
nor U11425 (N_11425,N_9091,N_8410);
and U11426 (N_11426,N_6919,N_8434);
nor U11427 (N_11427,N_7859,N_6380);
nor U11428 (N_11428,N_6704,N_8022);
nor U11429 (N_11429,N_9359,N_7336);
nand U11430 (N_11430,N_7988,N_7962);
or U11431 (N_11431,N_8662,N_6473);
or U11432 (N_11432,N_6735,N_9315);
and U11433 (N_11433,N_7905,N_8912);
or U11434 (N_11434,N_8473,N_8573);
nor U11435 (N_11435,N_8451,N_8067);
or U11436 (N_11436,N_8235,N_8175);
and U11437 (N_11437,N_8390,N_7934);
nand U11438 (N_11438,N_7837,N_7067);
nand U11439 (N_11439,N_7669,N_6566);
nand U11440 (N_11440,N_9067,N_7325);
xnor U11441 (N_11441,N_8329,N_7805);
nor U11442 (N_11442,N_7323,N_6759);
nand U11443 (N_11443,N_6365,N_8689);
or U11444 (N_11444,N_8550,N_6290);
nand U11445 (N_11445,N_6911,N_8240);
nand U11446 (N_11446,N_8389,N_7906);
nand U11447 (N_11447,N_7957,N_7489);
nor U11448 (N_11448,N_7371,N_7959);
xnor U11449 (N_11449,N_8097,N_8419);
or U11450 (N_11450,N_9137,N_9331);
nor U11451 (N_11451,N_9015,N_9074);
and U11452 (N_11452,N_7592,N_9341);
xnor U11453 (N_11453,N_8872,N_8661);
and U11454 (N_11454,N_8648,N_7280);
and U11455 (N_11455,N_9014,N_6956);
nand U11456 (N_11456,N_6482,N_6896);
nor U11457 (N_11457,N_7977,N_7072);
xor U11458 (N_11458,N_8268,N_8898);
nor U11459 (N_11459,N_8312,N_7296);
and U11460 (N_11460,N_7210,N_6993);
and U11461 (N_11461,N_6725,N_6686);
nor U11462 (N_11462,N_8105,N_8174);
nand U11463 (N_11463,N_6886,N_9058);
or U11464 (N_11464,N_7712,N_8945);
xnor U11465 (N_11465,N_7515,N_7026);
nor U11466 (N_11466,N_8443,N_8729);
nor U11467 (N_11467,N_7947,N_6797);
and U11468 (N_11468,N_7676,N_8388);
or U11469 (N_11469,N_7176,N_8565);
nor U11470 (N_11470,N_9311,N_6801);
and U11471 (N_11471,N_6464,N_7950);
xnor U11472 (N_11472,N_6588,N_8236);
nor U11473 (N_11473,N_6726,N_7950);
nand U11474 (N_11474,N_6664,N_7065);
and U11475 (N_11475,N_8050,N_8758);
or U11476 (N_11476,N_8225,N_6631);
or U11477 (N_11477,N_8197,N_6538);
nor U11478 (N_11478,N_8985,N_7615);
or U11479 (N_11479,N_7998,N_7513);
or U11480 (N_11480,N_7192,N_6285);
nand U11481 (N_11481,N_9023,N_8123);
and U11482 (N_11482,N_9361,N_8896);
or U11483 (N_11483,N_8871,N_8662);
or U11484 (N_11484,N_6771,N_8499);
and U11485 (N_11485,N_6823,N_7171);
nand U11486 (N_11486,N_7680,N_9172);
nand U11487 (N_11487,N_6889,N_7022);
xor U11488 (N_11488,N_8046,N_9226);
xor U11489 (N_11489,N_6829,N_7860);
nand U11490 (N_11490,N_6724,N_8568);
or U11491 (N_11491,N_6753,N_8639);
or U11492 (N_11492,N_8540,N_7864);
or U11493 (N_11493,N_6422,N_6454);
nand U11494 (N_11494,N_8534,N_7869);
nand U11495 (N_11495,N_8959,N_8792);
and U11496 (N_11496,N_6869,N_7982);
nand U11497 (N_11497,N_7956,N_6844);
xnor U11498 (N_11498,N_7827,N_8629);
and U11499 (N_11499,N_8483,N_8662);
and U11500 (N_11500,N_9351,N_7939);
nand U11501 (N_11501,N_7413,N_7053);
or U11502 (N_11502,N_8345,N_6473);
xor U11503 (N_11503,N_8760,N_7376);
nor U11504 (N_11504,N_7290,N_8346);
xnor U11505 (N_11505,N_8725,N_7054);
and U11506 (N_11506,N_8101,N_8934);
or U11507 (N_11507,N_8887,N_9254);
and U11508 (N_11508,N_9207,N_8159);
and U11509 (N_11509,N_6303,N_8922);
nand U11510 (N_11510,N_7146,N_8422);
and U11511 (N_11511,N_6394,N_8999);
nor U11512 (N_11512,N_9160,N_8121);
nor U11513 (N_11513,N_8192,N_8643);
nand U11514 (N_11514,N_6574,N_6592);
or U11515 (N_11515,N_6806,N_9287);
nor U11516 (N_11516,N_9072,N_6291);
nand U11517 (N_11517,N_8812,N_8342);
and U11518 (N_11518,N_6279,N_6411);
nor U11519 (N_11519,N_6527,N_8006);
nand U11520 (N_11520,N_8666,N_9083);
xor U11521 (N_11521,N_8062,N_8727);
xor U11522 (N_11522,N_7093,N_7158);
or U11523 (N_11523,N_8296,N_6428);
nand U11524 (N_11524,N_6481,N_6822);
xor U11525 (N_11525,N_7892,N_6824);
and U11526 (N_11526,N_6354,N_8186);
nand U11527 (N_11527,N_9128,N_8576);
and U11528 (N_11528,N_8745,N_8619);
nor U11529 (N_11529,N_7278,N_8283);
nor U11530 (N_11530,N_6592,N_8711);
and U11531 (N_11531,N_7289,N_8017);
or U11532 (N_11532,N_6364,N_8754);
and U11533 (N_11533,N_8577,N_6546);
nand U11534 (N_11534,N_9318,N_7466);
and U11535 (N_11535,N_7820,N_6430);
nand U11536 (N_11536,N_6825,N_9196);
nor U11537 (N_11537,N_8491,N_7485);
and U11538 (N_11538,N_7215,N_7668);
and U11539 (N_11539,N_6583,N_7345);
or U11540 (N_11540,N_7112,N_7225);
nand U11541 (N_11541,N_8438,N_6827);
or U11542 (N_11542,N_8704,N_8163);
nor U11543 (N_11543,N_8261,N_8777);
and U11544 (N_11544,N_7670,N_9293);
and U11545 (N_11545,N_9214,N_7273);
or U11546 (N_11546,N_6884,N_6652);
nor U11547 (N_11547,N_8445,N_7824);
and U11548 (N_11548,N_7522,N_8370);
nor U11549 (N_11549,N_6332,N_7969);
and U11550 (N_11550,N_8180,N_8789);
and U11551 (N_11551,N_7232,N_8475);
nand U11552 (N_11552,N_8681,N_9223);
xnor U11553 (N_11553,N_8547,N_6405);
nor U11554 (N_11554,N_6885,N_6797);
nor U11555 (N_11555,N_8227,N_9031);
or U11556 (N_11556,N_7932,N_8042);
nor U11557 (N_11557,N_8100,N_8901);
and U11558 (N_11558,N_7834,N_6780);
nor U11559 (N_11559,N_6255,N_8937);
or U11560 (N_11560,N_8681,N_8106);
and U11561 (N_11561,N_9233,N_9295);
nor U11562 (N_11562,N_6337,N_7812);
nand U11563 (N_11563,N_7755,N_7609);
or U11564 (N_11564,N_9138,N_8786);
or U11565 (N_11565,N_8899,N_7723);
nand U11566 (N_11566,N_8736,N_7005);
xnor U11567 (N_11567,N_7933,N_6254);
or U11568 (N_11568,N_6762,N_9317);
or U11569 (N_11569,N_9307,N_6580);
and U11570 (N_11570,N_9098,N_6489);
nand U11571 (N_11571,N_6338,N_7731);
nand U11572 (N_11572,N_9209,N_6341);
and U11573 (N_11573,N_8453,N_8473);
or U11574 (N_11574,N_6987,N_8470);
xnor U11575 (N_11575,N_7915,N_8106);
nand U11576 (N_11576,N_6297,N_7867);
or U11577 (N_11577,N_6638,N_8293);
or U11578 (N_11578,N_8315,N_8303);
nor U11579 (N_11579,N_7150,N_8787);
and U11580 (N_11580,N_8047,N_6304);
nor U11581 (N_11581,N_9329,N_7644);
or U11582 (N_11582,N_9352,N_7546);
nand U11583 (N_11583,N_8516,N_8163);
and U11584 (N_11584,N_9086,N_6391);
or U11585 (N_11585,N_7987,N_8578);
and U11586 (N_11586,N_9174,N_6319);
nand U11587 (N_11587,N_7992,N_7953);
and U11588 (N_11588,N_7093,N_7267);
nor U11589 (N_11589,N_7115,N_7028);
or U11590 (N_11590,N_6262,N_8933);
nor U11591 (N_11591,N_7521,N_9353);
nor U11592 (N_11592,N_6981,N_8704);
or U11593 (N_11593,N_9219,N_8024);
xor U11594 (N_11594,N_8705,N_7824);
nand U11595 (N_11595,N_8519,N_7315);
and U11596 (N_11596,N_6414,N_7623);
nand U11597 (N_11597,N_8345,N_7025);
or U11598 (N_11598,N_6424,N_7202);
and U11599 (N_11599,N_8977,N_9297);
nor U11600 (N_11600,N_8429,N_7435);
or U11601 (N_11601,N_7474,N_9091);
or U11602 (N_11602,N_6894,N_8968);
xor U11603 (N_11603,N_7791,N_6517);
nand U11604 (N_11604,N_7452,N_8545);
nor U11605 (N_11605,N_9300,N_7849);
and U11606 (N_11606,N_6462,N_7600);
and U11607 (N_11607,N_8084,N_9152);
nor U11608 (N_11608,N_7456,N_6267);
or U11609 (N_11609,N_7824,N_8785);
and U11610 (N_11610,N_7348,N_9074);
or U11611 (N_11611,N_6410,N_9210);
nand U11612 (N_11612,N_8110,N_6884);
xnor U11613 (N_11613,N_7653,N_6722);
and U11614 (N_11614,N_7528,N_8581);
or U11615 (N_11615,N_8970,N_8497);
and U11616 (N_11616,N_9075,N_8095);
or U11617 (N_11617,N_6632,N_8788);
nand U11618 (N_11618,N_7530,N_6798);
or U11619 (N_11619,N_7654,N_8453);
nand U11620 (N_11620,N_8141,N_8217);
nand U11621 (N_11621,N_6316,N_8193);
or U11622 (N_11622,N_6453,N_8009);
and U11623 (N_11623,N_6445,N_7200);
nand U11624 (N_11624,N_8757,N_6759);
nand U11625 (N_11625,N_8787,N_9200);
nor U11626 (N_11626,N_6283,N_9371);
xor U11627 (N_11627,N_9077,N_7732);
and U11628 (N_11628,N_8631,N_7184);
xor U11629 (N_11629,N_6465,N_7067);
or U11630 (N_11630,N_6934,N_7055);
and U11631 (N_11631,N_9033,N_6453);
nand U11632 (N_11632,N_7298,N_7701);
nor U11633 (N_11633,N_7455,N_7473);
nand U11634 (N_11634,N_7948,N_7329);
or U11635 (N_11635,N_8663,N_8866);
and U11636 (N_11636,N_6860,N_9360);
nor U11637 (N_11637,N_9128,N_7562);
or U11638 (N_11638,N_9138,N_6711);
nor U11639 (N_11639,N_8069,N_6327);
and U11640 (N_11640,N_7167,N_7312);
and U11641 (N_11641,N_7973,N_8502);
or U11642 (N_11642,N_7415,N_8108);
nor U11643 (N_11643,N_8761,N_7909);
xor U11644 (N_11644,N_7346,N_7780);
nor U11645 (N_11645,N_6735,N_8534);
nand U11646 (N_11646,N_8337,N_6514);
or U11647 (N_11647,N_7819,N_6370);
nand U11648 (N_11648,N_7599,N_8739);
nor U11649 (N_11649,N_6440,N_7767);
nor U11650 (N_11650,N_8659,N_8086);
and U11651 (N_11651,N_8807,N_6619);
and U11652 (N_11652,N_8358,N_6441);
nor U11653 (N_11653,N_7746,N_9319);
nand U11654 (N_11654,N_6885,N_8089);
xor U11655 (N_11655,N_9247,N_9214);
nand U11656 (N_11656,N_9176,N_7903);
nor U11657 (N_11657,N_9356,N_6916);
or U11658 (N_11658,N_6773,N_8066);
or U11659 (N_11659,N_6486,N_9242);
and U11660 (N_11660,N_8583,N_8840);
and U11661 (N_11661,N_8354,N_8800);
nor U11662 (N_11662,N_7566,N_6872);
nand U11663 (N_11663,N_8915,N_8230);
xor U11664 (N_11664,N_6470,N_6568);
or U11665 (N_11665,N_7411,N_7635);
and U11666 (N_11666,N_6971,N_7173);
nand U11667 (N_11667,N_9289,N_6363);
nor U11668 (N_11668,N_7116,N_9233);
or U11669 (N_11669,N_7776,N_6832);
nand U11670 (N_11670,N_9050,N_8839);
and U11671 (N_11671,N_7332,N_8186);
nor U11672 (N_11672,N_8056,N_8240);
nand U11673 (N_11673,N_6624,N_8981);
nand U11674 (N_11674,N_7371,N_7030);
and U11675 (N_11675,N_9253,N_6582);
nand U11676 (N_11676,N_7987,N_7724);
nand U11677 (N_11677,N_6846,N_7214);
nor U11678 (N_11678,N_8685,N_9348);
nand U11679 (N_11679,N_9206,N_9315);
nor U11680 (N_11680,N_6345,N_8666);
or U11681 (N_11681,N_6594,N_7673);
xnor U11682 (N_11682,N_7787,N_8467);
xnor U11683 (N_11683,N_6469,N_6649);
and U11684 (N_11684,N_7414,N_8459);
and U11685 (N_11685,N_8708,N_8302);
nor U11686 (N_11686,N_8461,N_6398);
nand U11687 (N_11687,N_8452,N_8956);
nor U11688 (N_11688,N_9133,N_6805);
nor U11689 (N_11689,N_8416,N_6766);
and U11690 (N_11690,N_7255,N_6863);
nand U11691 (N_11691,N_7504,N_7774);
nor U11692 (N_11692,N_9305,N_8842);
xnor U11693 (N_11693,N_8490,N_8834);
xnor U11694 (N_11694,N_6319,N_6545);
xor U11695 (N_11695,N_7866,N_6435);
nand U11696 (N_11696,N_8671,N_9123);
nor U11697 (N_11697,N_6256,N_9291);
xor U11698 (N_11698,N_7316,N_7134);
or U11699 (N_11699,N_6635,N_9275);
xnor U11700 (N_11700,N_8299,N_7471);
or U11701 (N_11701,N_6330,N_8558);
nand U11702 (N_11702,N_8365,N_8477);
nand U11703 (N_11703,N_7855,N_7092);
or U11704 (N_11704,N_9120,N_9049);
or U11705 (N_11705,N_8643,N_6740);
or U11706 (N_11706,N_6487,N_6938);
and U11707 (N_11707,N_8713,N_7342);
xor U11708 (N_11708,N_7027,N_6372);
or U11709 (N_11709,N_8195,N_7188);
nor U11710 (N_11710,N_7853,N_7539);
nor U11711 (N_11711,N_6955,N_6458);
or U11712 (N_11712,N_8911,N_8548);
nor U11713 (N_11713,N_7074,N_7208);
and U11714 (N_11714,N_9210,N_7741);
and U11715 (N_11715,N_8766,N_8967);
nor U11716 (N_11716,N_8788,N_6992);
or U11717 (N_11717,N_9069,N_7644);
nor U11718 (N_11718,N_9302,N_8412);
and U11719 (N_11719,N_6471,N_7952);
xnor U11720 (N_11720,N_8334,N_7369);
or U11721 (N_11721,N_8813,N_6418);
xor U11722 (N_11722,N_7094,N_8523);
nor U11723 (N_11723,N_8246,N_9091);
xnor U11724 (N_11724,N_8003,N_7275);
and U11725 (N_11725,N_7934,N_9154);
nor U11726 (N_11726,N_8423,N_9126);
xnor U11727 (N_11727,N_7190,N_7591);
nor U11728 (N_11728,N_7533,N_8738);
nor U11729 (N_11729,N_7043,N_6737);
and U11730 (N_11730,N_8342,N_8930);
nand U11731 (N_11731,N_8724,N_8311);
and U11732 (N_11732,N_7738,N_8985);
or U11733 (N_11733,N_6823,N_8827);
or U11734 (N_11734,N_7735,N_6380);
or U11735 (N_11735,N_8065,N_7739);
and U11736 (N_11736,N_8813,N_8506);
and U11737 (N_11737,N_6402,N_8223);
nand U11738 (N_11738,N_8245,N_8156);
nor U11739 (N_11739,N_8120,N_8053);
and U11740 (N_11740,N_8389,N_7489);
nor U11741 (N_11741,N_8777,N_6313);
or U11742 (N_11742,N_7793,N_8093);
and U11743 (N_11743,N_6387,N_8993);
nor U11744 (N_11744,N_6657,N_8170);
nand U11745 (N_11745,N_6862,N_7545);
and U11746 (N_11746,N_6508,N_8447);
nand U11747 (N_11747,N_6917,N_6357);
and U11748 (N_11748,N_7735,N_8166);
or U11749 (N_11749,N_6523,N_7892);
nor U11750 (N_11750,N_8766,N_8174);
xnor U11751 (N_11751,N_8561,N_6281);
nor U11752 (N_11752,N_7864,N_7264);
nand U11753 (N_11753,N_9333,N_7379);
nand U11754 (N_11754,N_7067,N_7694);
nand U11755 (N_11755,N_6580,N_7814);
and U11756 (N_11756,N_6734,N_8142);
or U11757 (N_11757,N_7644,N_7092);
nand U11758 (N_11758,N_9150,N_6339);
nor U11759 (N_11759,N_6419,N_8458);
and U11760 (N_11760,N_7759,N_6343);
nand U11761 (N_11761,N_7173,N_6616);
or U11762 (N_11762,N_8116,N_8012);
or U11763 (N_11763,N_7938,N_6289);
nor U11764 (N_11764,N_9187,N_8365);
or U11765 (N_11765,N_7326,N_9023);
or U11766 (N_11766,N_8049,N_8389);
nand U11767 (N_11767,N_7338,N_8661);
nor U11768 (N_11768,N_7691,N_6422);
nand U11769 (N_11769,N_6492,N_8363);
nand U11770 (N_11770,N_6311,N_6643);
or U11771 (N_11771,N_9000,N_8583);
nor U11772 (N_11772,N_8284,N_8377);
nand U11773 (N_11773,N_9329,N_8488);
and U11774 (N_11774,N_7417,N_7501);
or U11775 (N_11775,N_9130,N_8815);
nand U11776 (N_11776,N_8888,N_6301);
nor U11777 (N_11777,N_6995,N_8133);
nand U11778 (N_11778,N_6976,N_8341);
or U11779 (N_11779,N_9204,N_8252);
or U11780 (N_11780,N_7245,N_7547);
nand U11781 (N_11781,N_7916,N_7688);
nor U11782 (N_11782,N_7760,N_6997);
nor U11783 (N_11783,N_8780,N_8885);
nor U11784 (N_11784,N_7680,N_7095);
or U11785 (N_11785,N_7409,N_7095);
nand U11786 (N_11786,N_7876,N_8756);
nor U11787 (N_11787,N_8800,N_7824);
nor U11788 (N_11788,N_9309,N_7459);
or U11789 (N_11789,N_7388,N_7955);
xor U11790 (N_11790,N_7435,N_8173);
nand U11791 (N_11791,N_7863,N_8769);
nand U11792 (N_11792,N_8969,N_6318);
xor U11793 (N_11793,N_8967,N_7175);
xnor U11794 (N_11794,N_7751,N_6933);
or U11795 (N_11795,N_6351,N_8424);
nor U11796 (N_11796,N_9034,N_6637);
nand U11797 (N_11797,N_6645,N_7456);
xor U11798 (N_11798,N_8949,N_7184);
nand U11799 (N_11799,N_7037,N_7393);
nor U11800 (N_11800,N_6409,N_9049);
and U11801 (N_11801,N_8778,N_9210);
nand U11802 (N_11802,N_7068,N_7366);
nor U11803 (N_11803,N_9193,N_9219);
xnor U11804 (N_11804,N_6346,N_8551);
or U11805 (N_11805,N_9045,N_8633);
nor U11806 (N_11806,N_9282,N_8050);
and U11807 (N_11807,N_8461,N_7856);
or U11808 (N_11808,N_6251,N_6937);
nor U11809 (N_11809,N_9080,N_8979);
nor U11810 (N_11810,N_8378,N_9129);
xnor U11811 (N_11811,N_7199,N_9079);
or U11812 (N_11812,N_8883,N_8784);
and U11813 (N_11813,N_8754,N_8841);
nor U11814 (N_11814,N_8068,N_7033);
nand U11815 (N_11815,N_7540,N_8239);
or U11816 (N_11816,N_8847,N_6622);
and U11817 (N_11817,N_7426,N_6486);
nand U11818 (N_11818,N_6959,N_7206);
or U11819 (N_11819,N_7305,N_8743);
nand U11820 (N_11820,N_8031,N_8017);
and U11821 (N_11821,N_6445,N_8180);
nor U11822 (N_11822,N_7922,N_7518);
xor U11823 (N_11823,N_9073,N_7800);
and U11824 (N_11824,N_8235,N_7039);
nor U11825 (N_11825,N_8961,N_6773);
nand U11826 (N_11826,N_8753,N_8631);
and U11827 (N_11827,N_6875,N_8695);
xnor U11828 (N_11828,N_6555,N_6658);
xor U11829 (N_11829,N_8018,N_9287);
and U11830 (N_11830,N_8672,N_6320);
or U11831 (N_11831,N_9222,N_8317);
or U11832 (N_11832,N_7146,N_9077);
or U11833 (N_11833,N_8511,N_8367);
nor U11834 (N_11834,N_8957,N_7877);
and U11835 (N_11835,N_6769,N_6737);
or U11836 (N_11836,N_6843,N_8511);
and U11837 (N_11837,N_8847,N_7751);
nor U11838 (N_11838,N_9090,N_8209);
xor U11839 (N_11839,N_9282,N_8747);
nor U11840 (N_11840,N_7401,N_9095);
nand U11841 (N_11841,N_8390,N_7792);
and U11842 (N_11842,N_9313,N_6940);
or U11843 (N_11843,N_6735,N_6300);
and U11844 (N_11844,N_7180,N_6269);
xor U11845 (N_11845,N_7321,N_6467);
or U11846 (N_11846,N_7968,N_6692);
nand U11847 (N_11847,N_6794,N_9184);
nand U11848 (N_11848,N_8126,N_8778);
or U11849 (N_11849,N_9274,N_7783);
nor U11850 (N_11850,N_9324,N_8947);
nor U11851 (N_11851,N_7604,N_7413);
xnor U11852 (N_11852,N_9164,N_6674);
and U11853 (N_11853,N_8877,N_9071);
nor U11854 (N_11854,N_8182,N_9321);
and U11855 (N_11855,N_7279,N_9301);
nor U11856 (N_11856,N_7677,N_8825);
nand U11857 (N_11857,N_6419,N_6252);
nand U11858 (N_11858,N_7830,N_7844);
or U11859 (N_11859,N_8807,N_6999);
or U11860 (N_11860,N_8046,N_7712);
nand U11861 (N_11861,N_7477,N_9172);
and U11862 (N_11862,N_8510,N_9318);
or U11863 (N_11863,N_6808,N_7227);
nor U11864 (N_11864,N_8659,N_8802);
nand U11865 (N_11865,N_6282,N_8725);
nor U11866 (N_11866,N_6643,N_7180);
nand U11867 (N_11867,N_8302,N_7391);
and U11868 (N_11868,N_7565,N_8101);
xnor U11869 (N_11869,N_8732,N_7413);
nor U11870 (N_11870,N_8112,N_9252);
and U11871 (N_11871,N_7209,N_7320);
nand U11872 (N_11872,N_7611,N_8527);
nand U11873 (N_11873,N_6925,N_8381);
nor U11874 (N_11874,N_8421,N_8930);
xor U11875 (N_11875,N_7279,N_7108);
xor U11876 (N_11876,N_8550,N_8893);
nor U11877 (N_11877,N_9278,N_7500);
or U11878 (N_11878,N_8561,N_6325);
xor U11879 (N_11879,N_8861,N_9332);
and U11880 (N_11880,N_6857,N_8436);
or U11881 (N_11881,N_7408,N_8190);
and U11882 (N_11882,N_7251,N_9265);
xnor U11883 (N_11883,N_8851,N_6614);
xor U11884 (N_11884,N_6769,N_7490);
nand U11885 (N_11885,N_7883,N_7815);
nand U11886 (N_11886,N_8659,N_8263);
nor U11887 (N_11887,N_8377,N_6632);
nor U11888 (N_11888,N_6423,N_8288);
or U11889 (N_11889,N_8941,N_9369);
nor U11890 (N_11890,N_7742,N_7109);
xor U11891 (N_11891,N_7718,N_9115);
nand U11892 (N_11892,N_7894,N_7291);
nand U11893 (N_11893,N_8843,N_7345);
nor U11894 (N_11894,N_8431,N_8738);
nand U11895 (N_11895,N_8471,N_9161);
xnor U11896 (N_11896,N_9193,N_8722);
nand U11897 (N_11897,N_6897,N_9330);
and U11898 (N_11898,N_8269,N_6918);
nand U11899 (N_11899,N_8647,N_8708);
or U11900 (N_11900,N_8154,N_7466);
or U11901 (N_11901,N_7205,N_6387);
nor U11902 (N_11902,N_6659,N_7858);
nand U11903 (N_11903,N_8576,N_8755);
and U11904 (N_11904,N_8393,N_8830);
or U11905 (N_11905,N_9200,N_6741);
or U11906 (N_11906,N_7388,N_7978);
nor U11907 (N_11907,N_8699,N_8591);
nand U11908 (N_11908,N_7826,N_8065);
nor U11909 (N_11909,N_8057,N_6970);
xnor U11910 (N_11910,N_8294,N_7167);
and U11911 (N_11911,N_8748,N_8291);
nand U11912 (N_11912,N_8203,N_7833);
and U11913 (N_11913,N_6520,N_9243);
xor U11914 (N_11914,N_6355,N_8310);
and U11915 (N_11915,N_7950,N_8680);
nor U11916 (N_11916,N_8020,N_9024);
xor U11917 (N_11917,N_9281,N_6545);
nor U11918 (N_11918,N_7984,N_8188);
and U11919 (N_11919,N_8470,N_7770);
nand U11920 (N_11920,N_6892,N_8855);
nand U11921 (N_11921,N_7321,N_6372);
and U11922 (N_11922,N_6773,N_6850);
and U11923 (N_11923,N_7775,N_7615);
nor U11924 (N_11924,N_8018,N_8926);
or U11925 (N_11925,N_8003,N_6372);
xnor U11926 (N_11926,N_6599,N_8749);
and U11927 (N_11927,N_8399,N_7519);
or U11928 (N_11928,N_8564,N_7468);
or U11929 (N_11929,N_7391,N_6727);
nand U11930 (N_11930,N_7354,N_7987);
nand U11931 (N_11931,N_7608,N_9145);
nor U11932 (N_11932,N_7849,N_9362);
nand U11933 (N_11933,N_8696,N_7529);
nor U11934 (N_11934,N_6254,N_6826);
nand U11935 (N_11935,N_6809,N_7963);
nor U11936 (N_11936,N_8143,N_6633);
and U11937 (N_11937,N_7860,N_8902);
nor U11938 (N_11938,N_7852,N_8127);
nand U11939 (N_11939,N_7534,N_8971);
or U11940 (N_11940,N_7045,N_7470);
nand U11941 (N_11941,N_8539,N_9136);
or U11942 (N_11942,N_6934,N_7384);
xnor U11943 (N_11943,N_6292,N_7701);
and U11944 (N_11944,N_8821,N_7136);
nand U11945 (N_11945,N_8090,N_8451);
and U11946 (N_11946,N_6998,N_7906);
nand U11947 (N_11947,N_7701,N_8549);
nor U11948 (N_11948,N_7860,N_8750);
xor U11949 (N_11949,N_8788,N_8990);
nor U11950 (N_11950,N_6989,N_6760);
and U11951 (N_11951,N_7873,N_8049);
nand U11952 (N_11952,N_9365,N_6449);
and U11953 (N_11953,N_8568,N_7349);
nand U11954 (N_11954,N_8233,N_7451);
nor U11955 (N_11955,N_6335,N_6369);
nand U11956 (N_11956,N_8740,N_7273);
and U11957 (N_11957,N_8740,N_7564);
xor U11958 (N_11958,N_6448,N_7408);
or U11959 (N_11959,N_8576,N_8937);
nand U11960 (N_11960,N_8932,N_7921);
or U11961 (N_11961,N_8999,N_7876);
and U11962 (N_11962,N_7153,N_8730);
and U11963 (N_11963,N_7745,N_7247);
or U11964 (N_11964,N_8879,N_6395);
xnor U11965 (N_11965,N_8367,N_6416);
and U11966 (N_11966,N_6521,N_8954);
or U11967 (N_11967,N_6939,N_7422);
and U11968 (N_11968,N_7418,N_6756);
or U11969 (N_11969,N_9256,N_8070);
or U11970 (N_11970,N_9036,N_6663);
xor U11971 (N_11971,N_9308,N_6827);
nand U11972 (N_11972,N_7113,N_8370);
and U11973 (N_11973,N_8732,N_6411);
or U11974 (N_11974,N_7884,N_7543);
nand U11975 (N_11975,N_7309,N_8972);
or U11976 (N_11976,N_6734,N_8852);
and U11977 (N_11977,N_8441,N_8962);
nand U11978 (N_11978,N_7195,N_6994);
nor U11979 (N_11979,N_7363,N_7193);
or U11980 (N_11980,N_7473,N_8121);
or U11981 (N_11981,N_7349,N_7192);
nand U11982 (N_11982,N_8606,N_7747);
nand U11983 (N_11983,N_7940,N_7137);
nand U11984 (N_11984,N_8506,N_7660);
nand U11985 (N_11985,N_9233,N_7147);
or U11986 (N_11986,N_6440,N_7025);
nand U11987 (N_11987,N_6922,N_7966);
nor U11988 (N_11988,N_7123,N_7976);
nor U11989 (N_11989,N_8634,N_6370);
nor U11990 (N_11990,N_7137,N_7694);
or U11991 (N_11991,N_8366,N_8887);
and U11992 (N_11992,N_7908,N_7640);
nor U11993 (N_11993,N_7522,N_7451);
xnor U11994 (N_11994,N_7123,N_9239);
and U11995 (N_11995,N_7833,N_6629);
or U11996 (N_11996,N_8811,N_7060);
or U11997 (N_11997,N_7104,N_8136);
nand U11998 (N_11998,N_6946,N_9014);
nand U11999 (N_11999,N_8190,N_8589);
xor U12000 (N_12000,N_7990,N_8375);
and U12001 (N_12001,N_8154,N_6913);
and U12002 (N_12002,N_7900,N_6790);
nor U12003 (N_12003,N_8929,N_6359);
or U12004 (N_12004,N_8435,N_8107);
xnor U12005 (N_12005,N_7351,N_8225);
or U12006 (N_12006,N_8094,N_6315);
or U12007 (N_12007,N_8333,N_7635);
and U12008 (N_12008,N_8459,N_7894);
or U12009 (N_12009,N_8361,N_8182);
and U12010 (N_12010,N_6587,N_9184);
and U12011 (N_12011,N_9367,N_8210);
nor U12012 (N_12012,N_8205,N_9132);
or U12013 (N_12013,N_7497,N_7435);
and U12014 (N_12014,N_7884,N_9062);
nor U12015 (N_12015,N_6861,N_7274);
or U12016 (N_12016,N_9230,N_7520);
and U12017 (N_12017,N_8711,N_6711);
and U12018 (N_12018,N_8228,N_9318);
nor U12019 (N_12019,N_6402,N_8215);
nand U12020 (N_12020,N_8707,N_6736);
and U12021 (N_12021,N_7765,N_8905);
nand U12022 (N_12022,N_8972,N_8614);
xor U12023 (N_12023,N_6332,N_7857);
or U12024 (N_12024,N_6528,N_8606);
or U12025 (N_12025,N_6306,N_7068);
nor U12026 (N_12026,N_6679,N_8862);
and U12027 (N_12027,N_6574,N_8054);
nand U12028 (N_12028,N_7079,N_8990);
nor U12029 (N_12029,N_8172,N_6443);
and U12030 (N_12030,N_6964,N_9326);
or U12031 (N_12031,N_8318,N_7610);
or U12032 (N_12032,N_6266,N_8345);
nand U12033 (N_12033,N_6802,N_7022);
nand U12034 (N_12034,N_7249,N_7514);
nand U12035 (N_12035,N_8468,N_7168);
and U12036 (N_12036,N_6303,N_8488);
xor U12037 (N_12037,N_6937,N_8763);
nor U12038 (N_12038,N_9093,N_6351);
nor U12039 (N_12039,N_9242,N_6865);
nand U12040 (N_12040,N_6511,N_6761);
nand U12041 (N_12041,N_8870,N_6252);
nand U12042 (N_12042,N_7090,N_7150);
or U12043 (N_12043,N_6251,N_8958);
xor U12044 (N_12044,N_9169,N_7300);
nand U12045 (N_12045,N_8733,N_6972);
nor U12046 (N_12046,N_7281,N_6366);
xnor U12047 (N_12047,N_8193,N_8257);
nor U12048 (N_12048,N_8764,N_7346);
nand U12049 (N_12049,N_6905,N_7279);
nor U12050 (N_12050,N_8400,N_6301);
nor U12051 (N_12051,N_6888,N_7608);
nor U12052 (N_12052,N_7388,N_7691);
and U12053 (N_12053,N_6924,N_6369);
nand U12054 (N_12054,N_7263,N_8251);
nor U12055 (N_12055,N_6589,N_6669);
nor U12056 (N_12056,N_7838,N_9157);
nand U12057 (N_12057,N_8468,N_7225);
and U12058 (N_12058,N_6837,N_8388);
nor U12059 (N_12059,N_8733,N_7950);
nor U12060 (N_12060,N_9141,N_7317);
and U12061 (N_12061,N_7555,N_7723);
or U12062 (N_12062,N_8811,N_7717);
or U12063 (N_12063,N_8221,N_7089);
or U12064 (N_12064,N_7949,N_7858);
and U12065 (N_12065,N_6900,N_8577);
xor U12066 (N_12066,N_8559,N_8821);
nand U12067 (N_12067,N_8067,N_6616);
and U12068 (N_12068,N_8913,N_6324);
nor U12069 (N_12069,N_8407,N_6474);
and U12070 (N_12070,N_8380,N_6777);
nand U12071 (N_12071,N_7557,N_6598);
nand U12072 (N_12072,N_8766,N_7174);
nor U12073 (N_12073,N_7197,N_7652);
or U12074 (N_12074,N_9276,N_7244);
nand U12075 (N_12075,N_8625,N_6760);
xor U12076 (N_12076,N_8295,N_7689);
and U12077 (N_12077,N_8232,N_7290);
and U12078 (N_12078,N_9181,N_6713);
nor U12079 (N_12079,N_6514,N_6294);
nand U12080 (N_12080,N_9243,N_8936);
xnor U12081 (N_12081,N_7208,N_6495);
nor U12082 (N_12082,N_9099,N_7319);
and U12083 (N_12083,N_8834,N_6333);
or U12084 (N_12084,N_8607,N_8790);
or U12085 (N_12085,N_7468,N_6844);
nor U12086 (N_12086,N_7287,N_9338);
and U12087 (N_12087,N_7748,N_8142);
xnor U12088 (N_12088,N_7031,N_8012);
or U12089 (N_12089,N_9291,N_8056);
xor U12090 (N_12090,N_9090,N_7321);
nor U12091 (N_12091,N_7865,N_8393);
nand U12092 (N_12092,N_6848,N_9270);
or U12093 (N_12093,N_7706,N_6779);
nor U12094 (N_12094,N_8868,N_7141);
and U12095 (N_12095,N_8780,N_8414);
xor U12096 (N_12096,N_8534,N_7785);
nor U12097 (N_12097,N_9294,N_8434);
nand U12098 (N_12098,N_8049,N_6512);
or U12099 (N_12099,N_6662,N_6752);
nand U12100 (N_12100,N_8714,N_8556);
nor U12101 (N_12101,N_8506,N_6261);
nor U12102 (N_12102,N_6379,N_6845);
nor U12103 (N_12103,N_6364,N_7752);
and U12104 (N_12104,N_6738,N_6390);
or U12105 (N_12105,N_7841,N_7995);
and U12106 (N_12106,N_7698,N_9216);
nand U12107 (N_12107,N_8963,N_9087);
or U12108 (N_12108,N_6532,N_6330);
nor U12109 (N_12109,N_8534,N_7367);
nand U12110 (N_12110,N_8970,N_8170);
or U12111 (N_12111,N_6622,N_6430);
nand U12112 (N_12112,N_7735,N_6735);
or U12113 (N_12113,N_7376,N_8188);
and U12114 (N_12114,N_8718,N_7080);
or U12115 (N_12115,N_6708,N_8134);
nand U12116 (N_12116,N_8641,N_7441);
xor U12117 (N_12117,N_7318,N_8991);
nand U12118 (N_12118,N_8490,N_7605);
or U12119 (N_12119,N_8631,N_8922);
nor U12120 (N_12120,N_8510,N_9268);
xor U12121 (N_12121,N_6889,N_9229);
nor U12122 (N_12122,N_7360,N_8921);
and U12123 (N_12123,N_7000,N_8703);
nand U12124 (N_12124,N_6982,N_6467);
and U12125 (N_12125,N_8254,N_9331);
nor U12126 (N_12126,N_8260,N_8163);
or U12127 (N_12127,N_7532,N_6288);
and U12128 (N_12128,N_7188,N_7404);
or U12129 (N_12129,N_6467,N_8594);
xor U12130 (N_12130,N_6337,N_7837);
or U12131 (N_12131,N_8392,N_8881);
and U12132 (N_12132,N_9162,N_8664);
or U12133 (N_12133,N_8258,N_7142);
xor U12134 (N_12134,N_6996,N_9270);
nor U12135 (N_12135,N_7126,N_8404);
xor U12136 (N_12136,N_8350,N_8507);
or U12137 (N_12137,N_8247,N_7091);
nand U12138 (N_12138,N_6748,N_6362);
nand U12139 (N_12139,N_9260,N_7164);
and U12140 (N_12140,N_9213,N_6833);
nor U12141 (N_12141,N_8673,N_6308);
xor U12142 (N_12142,N_9164,N_6819);
nor U12143 (N_12143,N_8386,N_7614);
and U12144 (N_12144,N_7729,N_8033);
nor U12145 (N_12145,N_9264,N_8528);
nor U12146 (N_12146,N_6710,N_8773);
nand U12147 (N_12147,N_7737,N_8694);
and U12148 (N_12148,N_9085,N_7168);
nor U12149 (N_12149,N_8973,N_7219);
or U12150 (N_12150,N_7196,N_8754);
xor U12151 (N_12151,N_9062,N_6809);
and U12152 (N_12152,N_7013,N_7753);
nand U12153 (N_12153,N_8855,N_7547);
nor U12154 (N_12154,N_8787,N_7456);
xnor U12155 (N_12155,N_6336,N_8797);
nor U12156 (N_12156,N_6377,N_8959);
nand U12157 (N_12157,N_7025,N_8780);
and U12158 (N_12158,N_6345,N_7444);
nand U12159 (N_12159,N_6574,N_6495);
nor U12160 (N_12160,N_7085,N_7671);
nand U12161 (N_12161,N_8129,N_6624);
and U12162 (N_12162,N_7094,N_9140);
or U12163 (N_12163,N_7171,N_7704);
and U12164 (N_12164,N_6394,N_7080);
nor U12165 (N_12165,N_8093,N_8247);
or U12166 (N_12166,N_8528,N_8710);
nand U12167 (N_12167,N_9031,N_7384);
xnor U12168 (N_12168,N_9218,N_9356);
or U12169 (N_12169,N_7544,N_8249);
or U12170 (N_12170,N_8195,N_7562);
and U12171 (N_12171,N_7776,N_6309);
or U12172 (N_12172,N_6348,N_6817);
xnor U12173 (N_12173,N_7137,N_9050);
nor U12174 (N_12174,N_7051,N_6885);
xor U12175 (N_12175,N_6331,N_8793);
nand U12176 (N_12176,N_8558,N_6815);
nor U12177 (N_12177,N_8125,N_7886);
xor U12178 (N_12178,N_8840,N_9214);
nor U12179 (N_12179,N_8413,N_8012);
nor U12180 (N_12180,N_7757,N_6801);
nand U12181 (N_12181,N_8408,N_7021);
xor U12182 (N_12182,N_6817,N_7718);
xor U12183 (N_12183,N_7251,N_7362);
and U12184 (N_12184,N_8332,N_8479);
or U12185 (N_12185,N_9269,N_8759);
nand U12186 (N_12186,N_8937,N_6952);
nor U12187 (N_12187,N_8559,N_6391);
nand U12188 (N_12188,N_6339,N_7921);
nor U12189 (N_12189,N_6664,N_6938);
nor U12190 (N_12190,N_6519,N_7814);
nand U12191 (N_12191,N_9214,N_9331);
nand U12192 (N_12192,N_8860,N_8967);
nand U12193 (N_12193,N_7269,N_7796);
xor U12194 (N_12194,N_9207,N_8882);
or U12195 (N_12195,N_6724,N_8828);
or U12196 (N_12196,N_7963,N_6946);
nor U12197 (N_12197,N_7227,N_7858);
xnor U12198 (N_12198,N_7394,N_9311);
nor U12199 (N_12199,N_7901,N_8330);
or U12200 (N_12200,N_8838,N_8966);
xnor U12201 (N_12201,N_9007,N_8580);
and U12202 (N_12202,N_6874,N_7029);
and U12203 (N_12203,N_6311,N_7499);
or U12204 (N_12204,N_7910,N_7502);
and U12205 (N_12205,N_6269,N_7055);
nor U12206 (N_12206,N_8127,N_7642);
nand U12207 (N_12207,N_7328,N_9270);
or U12208 (N_12208,N_7971,N_9348);
nand U12209 (N_12209,N_9215,N_8776);
nand U12210 (N_12210,N_6680,N_9099);
or U12211 (N_12211,N_8978,N_6484);
and U12212 (N_12212,N_7608,N_7957);
nand U12213 (N_12213,N_7790,N_7546);
xor U12214 (N_12214,N_7933,N_7576);
xnor U12215 (N_12215,N_8262,N_8567);
nand U12216 (N_12216,N_7516,N_7789);
xnor U12217 (N_12217,N_6650,N_7212);
nor U12218 (N_12218,N_6913,N_8196);
nand U12219 (N_12219,N_9175,N_8632);
and U12220 (N_12220,N_9327,N_6987);
and U12221 (N_12221,N_8560,N_9085);
nor U12222 (N_12222,N_7410,N_8830);
and U12223 (N_12223,N_6526,N_8110);
nor U12224 (N_12224,N_9013,N_8027);
and U12225 (N_12225,N_8583,N_7083);
and U12226 (N_12226,N_7465,N_8696);
or U12227 (N_12227,N_6851,N_7678);
and U12228 (N_12228,N_8890,N_8769);
or U12229 (N_12229,N_7122,N_7946);
nor U12230 (N_12230,N_8749,N_7655);
nand U12231 (N_12231,N_6532,N_7311);
nand U12232 (N_12232,N_7972,N_8133);
nand U12233 (N_12233,N_7362,N_7614);
nor U12234 (N_12234,N_8089,N_7898);
nor U12235 (N_12235,N_6843,N_7496);
and U12236 (N_12236,N_8991,N_8420);
and U12237 (N_12237,N_9076,N_6540);
nor U12238 (N_12238,N_8177,N_8509);
or U12239 (N_12239,N_8465,N_8220);
or U12240 (N_12240,N_8643,N_8482);
nor U12241 (N_12241,N_8583,N_9186);
or U12242 (N_12242,N_8055,N_8525);
and U12243 (N_12243,N_7123,N_6898);
nand U12244 (N_12244,N_7468,N_7015);
or U12245 (N_12245,N_9020,N_8096);
and U12246 (N_12246,N_8159,N_8525);
nor U12247 (N_12247,N_8592,N_6385);
and U12248 (N_12248,N_8090,N_8144);
and U12249 (N_12249,N_7695,N_7949);
or U12250 (N_12250,N_8069,N_7748);
and U12251 (N_12251,N_7411,N_8444);
nand U12252 (N_12252,N_7999,N_8769);
or U12253 (N_12253,N_7786,N_7618);
nor U12254 (N_12254,N_7864,N_7650);
xnor U12255 (N_12255,N_9339,N_7788);
nand U12256 (N_12256,N_7481,N_7496);
and U12257 (N_12257,N_8403,N_9280);
and U12258 (N_12258,N_6866,N_8180);
nor U12259 (N_12259,N_6528,N_7098);
or U12260 (N_12260,N_9084,N_6498);
nand U12261 (N_12261,N_8091,N_8937);
or U12262 (N_12262,N_6827,N_6896);
nor U12263 (N_12263,N_7818,N_6386);
or U12264 (N_12264,N_7468,N_8394);
nand U12265 (N_12265,N_6840,N_6269);
nor U12266 (N_12266,N_6812,N_6345);
nor U12267 (N_12267,N_6530,N_7535);
or U12268 (N_12268,N_7098,N_7672);
or U12269 (N_12269,N_8725,N_6741);
and U12270 (N_12270,N_7395,N_6739);
and U12271 (N_12271,N_7320,N_7639);
or U12272 (N_12272,N_8305,N_7863);
xor U12273 (N_12273,N_8987,N_8525);
nor U12274 (N_12274,N_7175,N_6959);
and U12275 (N_12275,N_7974,N_7801);
or U12276 (N_12276,N_6483,N_7843);
xor U12277 (N_12277,N_8943,N_7162);
nand U12278 (N_12278,N_7051,N_8513);
xor U12279 (N_12279,N_8455,N_6417);
or U12280 (N_12280,N_6964,N_8815);
nor U12281 (N_12281,N_7329,N_9099);
and U12282 (N_12282,N_6280,N_8184);
nand U12283 (N_12283,N_8135,N_8289);
xnor U12284 (N_12284,N_9040,N_8164);
and U12285 (N_12285,N_9264,N_8906);
xor U12286 (N_12286,N_9181,N_8243);
and U12287 (N_12287,N_6336,N_8229);
nand U12288 (N_12288,N_6748,N_7748);
xor U12289 (N_12289,N_6881,N_7927);
nor U12290 (N_12290,N_8401,N_7387);
nand U12291 (N_12291,N_7938,N_6582);
nand U12292 (N_12292,N_7837,N_9053);
or U12293 (N_12293,N_8230,N_7414);
nor U12294 (N_12294,N_6909,N_6770);
or U12295 (N_12295,N_9365,N_7013);
and U12296 (N_12296,N_8112,N_8154);
and U12297 (N_12297,N_9317,N_8265);
nor U12298 (N_12298,N_8964,N_8561);
or U12299 (N_12299,N_8525,N_8361);
or U12300 (N_12300,N_6518,N_7497);
nand U12301 (N_12301,N_6610,N_8135);
or U12302 (N_12302,N_7158,N_9136);
nor U12303 (N_12303,N_6953,N_8004);
or U12304 (N_12304,N_9239,N_7285);
or U12305 (N_12305,N_6764,N_7717);
nor U12306 (N_12306,N_7452,N_8840);
nand U12307 (N_12307,N_7726,N_9320);
nor U12308 (N_12308,N_9071,N_7809);
nand U12309 (N_12309,N_8031,N_7725);
xnor U12310 (N_12310,N_9073,N_8669);
xor U12311 (N_12311,N_8818,N_7414);
nor U12312 (N_12312,N_8482,N_7469);
and U12313 (N_12313,N_6906,N_8427);
and U12314 (N_12314,N_8360,N_7604);
nor U12315 (N_12315,N_7335,N_8085);
and U12316 (N_12316,N_7802,N_6407);
nor U12317 (N_12317,N_8678,N_8470);
nor U12318 (N_12318,N_8442,N_7277);
nor U12319 (N_12319,N_8134,N_8961);
xor U12320 (N_12320,N_9220,N_7721);
nand U12321 (N_12321,N_8462,N_8064);
nor U12322 (N_12322,N_8185,N_7149);
or U12323 (N_12323,N_7272,N_8207);
nand U12324 (N_12324,N_7097,N_7747);
and U12325 (N_12325,N_7110,N_7045);
xnor U12326 (N_12326,N_8503,N_6402);
or U12327 (N_12327,N_6732,N_7387);
nor U12328 (N_12328,N_8519,N_7682);
or U12329 (N_12329,N_8183,N_9107);
nand U12330 (N_12330,N_9113,N_8094);
and U12331 (N_12331,N_6607,N_7343);
and U12332 (N_12332,N_7147,N_7703);
and U12333 (N_12333,N_8346,N_6580);
xnor U12334 (N_12334,N_7992,N_7437);
nor U12335 (N_12335,N_6921,N_9101);
and U12336 (N_12336,N_9228,N_6641);
or U12337 (N_12337,N_8180,N_6526);
and U12338 (N_12338,N_8190,N_8647);
nor U12339 (N_12339,N_6419,N_6956);
nand U12340 (N_12340,N_6871,N_6291);
or U12341 (N_12341,N_8989,N_8915);
nand U12342 (N_12342,N_6281,N_6816);
xnor U12343 (N_12343,N_9007,N_9221);
and U12344 (N_12344,N_7897,N_7592);
nand U12345 (N_12345,N_9061,N_6329);
or U12346 (N_12346,N_7348,N_9342);
xor U12347 (N_12347,N_8209,N_7887);
nor U12348 (N_12348,N_8513,N_8233);
nor U12349 (N_12349,N_7166,N_9106);
nand U12350 (N_12350,N_9200,N_7608);
or U12351 (N_12351,N_6790,N_6767);
and U12352 (N_12352,N_6895,N_7421);
nor U12353 (N_12353,N_9322,N_8020);
nand U12354 (N_12354,N_7929,N_7378);
or U12355 (N_12355,N_8101,N_8482);
and U12356 (N_12356,N_8677,N_6806);
and U12357 (N_12357,N_8475,N_8519);
or U12358 (N_12358,N_8996,N_8305);
nand U12359 (N_12359,N_6255,N_8338);
or U12360 (N_12360,N_7345,N_9235);
nor U12361 (N_12361,N_6513,N_7177);
xnor U12362 (N_12362,N_8720,N_8317);
nor U12363 (N_12363,N_8819,N_9234);
and U12364 (N_12364,N_8967,N_7143);
or U12365 (N_12365,N_7259,N_6731);
nor U12366 (N_12366,N_7592,N_7628);
nand U12367 (N_12367,N_8499,N_7994);
nand U12368 (N_12368,N_7631,N_9365);
nand U12369 (N_12369,N_7445,N_7692);
and U12370 (N_12370,N_7335,N_7450);
and U12371 (N_12371,N_6704,N_6366);
nand U12372 (N_12372,N_7800,N_7700);
nor U12373 (N_12373,N_7565,N_6392);
nor U12374 (N_12374,N_8965,N_6825);
nand U12375 (N_12375,N_7603,N_7684);
nor U12376 (N_12376,N_8479,N_9002);
nand U12377 (N_12377,N_7214,N_6417);
nand U12378 (N_12378,N_8051,N_9045);
and U12379 (N_12379,N_7067,N_8403);
nand U12380 (N_12380,N_9190,N_8986);
and U12381 (N_12381,N_6587,N_7864);
nor U12382 (N_12382,N_7878,N_8026);
nand U12383 (N_12383,N_9344,N_9126);
or U12384 (N_12384,N_8547,N_8473);
nand U12385 (N_12385,N_6898,N_8850);
or U12386 (N_12386,N_7383,N_6315);
nor U12387 (N_12387,N_7109,N_6702);
nor U12388 (N_12388,N_6931,N_8984);
or U12389 (N_12389,N_8302,N_8538);
nand U12390 (N_12390,N_6677,N_8289);
and U12391 (N_12391,N_8978,N_8574);
xnor U12392 (N_12392,N_8231,N_7865);
xor U12393 (N_12393,N_8978,N_9049);
and U12394 (N_12394,N_7184,N_9115);
nand U12395 (N_12395,N_9177,N_6656);
nor U12396 (N_12396,N_8970,N_9221);
and U12397 (N_12397,N_7211,N_7735);
nand U12398 (N_12398,N_8069,N_8426);
nand U12399 (N_12399,N_8676,N_6768);
nand U12400 (N_12400,N_7928,N_7734);
nand U12401 (N_12401,N_8809,N_9072);
nand U12402 (N_12402,N_9244,N_8842);
nand U12403 (N_12403,N_8427,N_7740);
and U12404 (N_12404,N_6484,N_9137);
xnor U12405 (N_12405,N_7868,N_7442);
or U12406 (N_12406,N_8586,N_6644);
nand U12407 (N_12407,N_6346,N_6826);
nor U12408 (N_12408,N_6445,N_8608);
and U12409 (N_12409,N_7045,N_6927);
or U12410 (N_12410,N_8110,N_7443);
or U12411 (N_12411,N_8980,N_8764);
nand U12412 (N_12412,N_6259,N_7267);
xnor U12413 (N_12413,N_7531,N_7292);
or U12414 (N_12414,N_7506,N_7180);
nor U12415 (N_12415,N_9230,N_7070);
nor U12416 (N_12416,N_8228,N_9185);
nand U12417 (N_12417,N_7830,N_8669);
and U12418 (N_12418,N_7773,N_8371);
nor U12419 (N_12419,N_9114,N_8909);
or U12420 (N_12420,N_7711,N_8756);
nand U12421 (N_12421,N_7283,N_7142);
nand U12422 (N_12422,N_8802,N_6270);
or U12423 (N_12423,N_7300,N_6874);
nor U12424 (N_12424,N_8637,N_8509);
nor U12425 (N_12425,N_7311,N_9211);
nand U12426 (N_12426,N_6380,N_7833);
or U12427 (N_12427,N_6495,N_6731);
nand U12428 (N_12428,N_9176,N_9206);
and U12429 (N_12429,N_9044,N_8468);
nor U12430 (N_12430,N_7018,N_8625);
xor U12431 (N_12431,N_7804,N_6758);
nand U12432 (N_12432,N_8547,N_7552);
and U12433 (N_12433,N_7592,N_7631);
or U12434 (N_12434,N_8186,N_9011);
nor U12435 (N_12435,N_7758,N_7810);
xor U12436 (N_12436,N_8495,N_8740);
nor U12437 (N_12437,N_6411,N_8392);
nor U12438 (N_12438,N_7126,N_6421);
and U12439 (N_12439,N_8031,N_9088);
xnor U12440 (N_12440,N_6960,N_6907);
xor U12441 (N_12441,N_8961,N_7239);
nor U12442 (N_12442,N_6778,N_7793);
nand U12443 (N_12443,N_6859,N_8424);
xnor U12444 (N_12444,N_6309,N_8884);
or U12445 (N_12445,N_6422,N_8209);
nor U12446 (N_12446,N_8044,N_7094);
nand U12447 (N_12447,N_6318,N_9067);
and U12448 (N_12448,N_7313,N_8529);
nand U12449 (N_12449,N_8320,N_7134);
nand U12450 (N_12450,N_7302,N_7355);
nand U12451 (N_12451,N_7067,N_8223);
xnor U12452 (N_12452,N_6755,N_8319);
nand U12453 (N_12453,N_7370,N_7591);
nor U12454 (N_12454,N_7070,N_8666);
xnor U12455 (N_12455,N_6309,N_9339);
nor U12456 (N_12456,N_8254,N_8611);
xnor U12457 (N_12457,N_6386,N_8098);
nand U12458 (N_12458,N_6388,N_7276);
xnor U12459 (N_12459,N_8789,N_6369);
or U12460 (N_12460,N_8862,N_7193);
or U12461 (N_12461,N_8621,N_6290);
and U12462 (N_12462,N_6983,N_6269);
and U12463 (N_12463,N_6537,N_6608);
or U12464 (N_12464,N_7917,N_9043);
nor U12465 (N_12465,N_6524,N_9219);
and U12466 (N_12466,N_8125,N_7304);
or U12467 (N_12467,N_7891,N_7959);
or U12468 (N_12468,N_6975,N_6357);
nand U12469 (N_12469,N_7800,N_6692);
nand U12470 (N_12470,N_8216,N_9002);
or U12471 (N_12471,N_9190,N_9027);
nor U12472 (N_12472,N_7827,N_8375);
and U12473 (N_12473,N_6525,N_7501);
nand U12474 (N_12474,N_7904,N_6669);
nor U12475 (N_12475,N_6499,N_7324);
nand U12476 (N_12476,N_7253,N_6516);
or U12477 (N_12477,N_8539,N_6460);
or U12478 (N_12478,N_6626,N_7721);
or U12479 (N_12479,N_6604,N_6932);
nand U12480 (N_12480,N_9099,N_9171);
nand U12481 (N_12481,N_6622,N_8160);
nand U12482 (N_12482,N_6343,N_8498);
and U12483 (N_12483,N_7496,N_8950);
and U12484 (N_12484,N_7032,N_8067);
and U12485 (N_12485,N_7921,N_6780);
or U12486 (N_12486,N_8387,N_8004);
nor U12487 (N_12487,N_8007,N_8127);
and U12488 (N_12488,N_6573,N_9091);
nor U12489 (N_12489,N_8780,N_7304);
and U12490 (N_12490,N_7934,N_6614);
xor U12491 (N_12491,N_9247,N_7620);
nand U12492 (N_12492,N_6723,N_6396);
nor U12493 (N_12493,N_7828,N_8532);
and U12494 (N_12494,N_9244,N_8113);
nand U12495 (N_12495,N_8540,N_7730);
or U12496 (N_12496,N_8819,N_7089);
and U12497 (N_12497,N_8817,N_8445);
nand U12498 (N_12498,N_9084,N_8683);
nand U12499 (N_12499,N_8306,N_9092);
nor U12500 (N_12500,N_10840,N_9826);
nand U12501 (N_12501,N_9399,N_10077);
and U12502 (N_12502,N_10709,N_10549);
or U12503 (N_12503,N_11104,N_9450);
nor U12504 (N_12504,N_9931,N_9560);
nand U12505 (N_12505,N_12113,N_11648);
nand U12506 (N_12506,N_10906,N_10455);
nand U12507 (N_12507,N_11397,N_9938);
and U12508 (N_12508,N_9472,N_12036);
nand U12509 (N_12509,N_9394,N_11944);
xor U12510 (N_12510,N_10281,N_9829);
nor U12511 (N_12511,N_9867,N_12399);
nand U12512 (N_12512,N_12172,N_11711);
nand U12513 (N_12513,N_12305,N_10762);
and U12514 (N_12514,N_10784,N_9477);
nand U12515 (N_12515,N_12043,N_11151);
nor U12516 (N_12516,N_10988,N_12034);
xor U12517 (N_12517,N_9762,N_12246);
and U12518 (N_12518,N_9856,N_9678);
nand U12519 (N_12519,N_10485,N_11601);
nor U12520 (N_12520,N_10786,N_9433);
and U12521 (N_12521,N_10695,N_10137);
and U12522 (N_12522,N_9887,N_12217);
nand U12523 (N_12523,N_10307,N_11573);
and U12524 (N_12524,N_10778,N_12465);
nor U12525 (N_12525,N_11168,N_10966);
nand U12526 (N_12526,N_9865,N_12134);
and U12527 (N_12527,N_10812,N_12233);
or U12528 (N_12528,N_10846,N_11886);
xor U12529 (N_12529,N_10951,N_10139);
nand U12530 (N_12530,N_10808,N_9504);
or U12531 (N_12531,N_10359,N_12178);
and U12532 (N_12532,N_11914,N_9499);
nor U12533 (N_12533,N_11161,N_11976);
or U12534 (N_12534,N_9387,N_12184);
nor U12535 (N_12535,N_11278,N_10826);
nor U12536 (N_12536,N_10677,N_10970);
or U12537 (N_12537,N_11460,N_10130);
and U12538 (N_12538,N_11584,N_10590);
nand U12539 (N_12539,N_12253,N_9976);
nor U12540 (N_12540,N_9385,N_12224);
or U12541 (N_12541,N_12135,N_10361);
or U12542 (N_12542,N_10004,N_9733);
or U12543 (N_12543,N_9429,N_10327);
and U12544 (N_12544,N_12182,N_10685);
or U12545 (N_12545,N_11348,N_9444);
or U12546 (N_12546,N_11708,N_11712);
nor U12547 (N_12547,N_10201,N_11930);
nand U12548 (N_12548,N_12153,N_10880);
nand U12549 (N_12549,N_11144,N_9841);
and U12550 (N_12550,N_11231,N_11788);
nand U12551 (N_12551,N_11963,N_10664);
nand U12552 (N_12552,N_11051,N_11483);
or U12553 (N_12553,N_10541,N_11787);
nor U12554 (N_12554,N_10204,N_11575);
and U12555 (N_12555,N_11668,N_11453);
or U12556 (N_12556,N_9383,N_9618);
or U12557 (N_12557,N_9899,N_12053);
nor U12558 (N_12558,N_12205,N_9936);
nor U12559 (N_12559,N_11524,N_9481);
or U12560 (N_12560,N_10374,N_11904);
nor U12561 (N_12561,N_11894,N_10122);
and U12562 (N_12562,N_11109,N_10183);
nand U12563 (N_12563,N_11719,N_10551);
xor U12564 (N_12564,N_9777,N_9945);
nand U12565 (N_12565,N_10793,N_9766);
and U12566 (N_12566,N_9807,N_10791);
nor U12567 (N_12567,N_10629,N_9760);
xor U12568 (N_12568,N_12125,N_11991);
xor U12569 (N_12569,N_10819,N_10440);
or U12570 (N_12570,N_9812,N_9833);
and U12571 (N_12571,N_12219,N_10255);
or U12572 (N_12572,N_10010,N_10962);
nand U12573 (N_12573,N_10473,N_10698);
and U12574 (N_12574,N_11841,N_11842);
and U12575 (N_12575,N_9600,N_11451);
nor U12576 (N_12576,N_10048,N_12140);
or U12577 (N_12577,N_12292,N_9602);
nor U12578 (N_12578,N_10087,N_12107);
or U12579 (N_12579,N_10250,N_9451);
nand U12580 (N_12580,N_11866,N_10965);
and U12581 (N_12581,N_10538,N_11375);
and U12582 (N_12582,N_11047,N_11706);
and U12583 (N_12583,N_9836,N_10957);
nand U12584 (N_12584,N_11628,N_11316);
and U12585 (N_12585,N_11924,N_11704);
and U12586 (N_12586,N_11121,N_10895);
nor U12587 (N_12587,N_11385,N_11836);
nand U12588 (N_12588,N_10510,N_10958);
and U12589 (N_12589,N_9495,N_12032);
nor U12590 (N_12590,N_9568,N_10815);
or U12591 (N_12591,N_12128,N_9443);
and U12592 (N_12592,N_10469,N_9420);
nor U12593 (N_12593,N_12151,N_9715);
nor U12594 (N_12594,N_10796,N_11057);
nor U12595 (N_12595,N_10940,N_12346);
nand U12596 (N_12596,N_11175,N_9874);
and U12597 (N_12597,N_11779,N_10712);
nor U12598 (N_12598,N_10305,N_10755);
nor U12599 (N_12599,N_10852,N_11741);
nand U12600 (N_12600,N_10804,N_11245);
nor U12601 (N_12601,N_11891,N_9554);
or U12602 (N_12602,N_10696,N_12270);
xnor U12603 (N_12603,N_11063,N_10902);
xor U12604 (N_12604,N_11188,N_10015);
and U12605 (N_12605,N_9978,N_11631);
nor U12606 (N_12606,N_12022,N_12301);
nand U12607 (N_12607,N_10877,N_12411);
nand U12608 (N_12608,N_9390,N_10302);
or U12609 (N_12609,N_10419,N_10609);
or U12610 (N_12610,N_10739,N_11226);
nand U12611 (N_12611,N_11939,N_10089);
and U12612 (N_12612,N_12384,N_11064);
nand U12613 (N_12613,N_9688,N_10949);
or U12614 (N_12614,N_10269,N_12031);
and U12615 (N_12615,N_11139,N_12244);
nor U12616 (N_12616,N_10956,N_11880);
and U12617 (N_12617,N_9647,N_10758);
or U12618 (N_12618,N_11156,N_11079);
or U12619 (N_12619,N_9778,N_10661);
nand U12620 (N_12620,N_12317,N_12392);
nand U12621 (N_12621,N_10625,N_10272);
nand U12622 (N_12622,N_11496,N_9934);
or U12623 (N_12623,N_10772,N_11958);
xnor U12624 (N_12624,N_10379,N_11693);
or U12625 (N_12625,N_9644,N_9752);
nor U12626 (N_12626,N_10737,N_12453);
xor U12627 (N_12627,N_12241,N_12359);
and U12628 (N_12628,N_12288,N_10224);
nand U12629 (N_12629,N_10330,N_12426);
or U12630 (N_12630,N_9659,N_9658);
nor U12631 (N_12631,N_11464,N_12044);
and U12632 (N_12632,N_11197,N_12327);
nor U12633 (N_12633,N_10760,N_10024);
or U12634 (N_12634,N_12371,N_9475);
nand U12635 (N_12635,N_11776,N_9438);
nor U12636 (N_12636,N_12297,N_12108);
xor U12637 (N_12637,N_11644,N_11086);
xor U12638 (N_12638,N_10433,N_11697);
or U12639 (N_12639,N_10865,N_11810);
or U12640 (N_12640,N_11362,N_9977);
and U12641 (N_12641,N_10557,N_12167);
nand U12642 (N_12642,N_11509,N_11185);
or U12643 (N_12643,N_11258,N_10291);
nand U12644 (N_12644,N_9631,N_11195);
nor U12645 (N_12645,N_11030,N_11123);
nand U12646 (N_12646,N_9657,N_12132);
nand U12647 (N_12647,N_12148,N_9392);
or U12648 (N_12648,N_10173,N_9651);
or U12649 (N_12649,N_10883,N_12454);
nand U12650 (N_12650,N_9538,N_10351);
nand U12651 (N_12651,N_11018,N_9548);
nand U12652 (N_12652,N_10697,N_10171);
and U12653 (N_12653,N_10991,N_12006);
nor U12654 (N_12654,N_12144,N_12499);
xor U12655 (N_12655,N_12204,N_12252);
xor U12656 (N_12656,N_10761,N_10411);
nor U12657 (N_12657,N_11284,N_10052);
nand U12658 (N_12658,N_10336,N_10561);
nand U12659 (N_12659,N_11795,N_9819);
and U12660 (N_12660,N_10532,N_11102);
nor U12661 (N_12661,N_12494,N_11476);
or U12662 (N_12662,N_9754,N_10413);
and U12663 (N_12663,N_10247,N_9787);
and U12664 (N_12664,N_11905,N_10656);
nand U12665 (N_12665,N_10412,N_12061);
nand U12666 (N_12666,N_9736,N_10064);
or U12667 (N_12667,N_9601,N_11837);
or U12668 (N_12668,N_9409,N_9842);
nor U12669 (N_12669,N_11032,N_12290);
xnor U12670 (N_12670,N_11927,N_11539);
nor U12671 (N_12671,N_11877,N_9997);
xor U12672 (N_12672,N_9942,N_9698);
or U12673 (N_12673,N_12177,N_11270);
nand U12674 (N_12674,N_10900,N_10025);
and U12675 (N_12675,N_12459,N_11408);
nand U12676 (N_12676,N_9963,N_11067);
or U12677 (N_12677,N_9671,N_12115);
nor U12678 (N_12678,N_10020,N_11731);
nor U12679 (N_12679,N_9407,N_11224);
nor U12680 (N_12680,N_10981,N_11046);
nor U12681 (N_12681,N_10713,N_9376);
nor U12682 (N_12682,N_11082,N_11178);
nand U12683 (N_12683,N_10873,N_11636);
nand U12684 (N_12684,N_10492,N_10870);
or U12685 (N_12685,N_10471,N_10517);
and U12686 (N_12686,N_9723,N_12079);
and U12687 (N_12687,N_11507,N_12491);
nand U12688 (N_12688,N_9531,N_12187);
nand U12689 (N_12689,N_12446,N_12235);
nor U12690 (N_12690,N_11972,N_9545);
and U12691 (N_12691,N_11140,N_9650);
or U12692 (N_12692,N_9508,N_10205);
and U12693 (N_12693,N_11449,N_11095);
nand U12694 (N_12694,N_11743,N_11753);
nor U12695 (N_12695,N_12183,N_10780);
nor U12696 (N_12696,N_12016,N_10501);
and U12697 (N_12697,N_11860,N_10803);
and U12698 (N_12698,N_10842,N_10134);
nor U12699 (N_12699,N_11638,N_12025);
or U12700 (N_12700,N_11006,N_10095);
nand U12701 (N_12701,N_10421,N_10974);
and U12702 (N_12702,N_12296,N_9608);
xor U12703 (N_12703,N_10820,N_11988);
nor U12704 (N_12704,N_9578,N_9908);
xor U12705 (N_12705,N_12112,N_10719);
nor U12706 (N_12706,N_11026,N_11153);
nor U12707 (N_12707,N_12412,N_12498);
nor U12708 (N_12708,N_10494,N_10216);
and U12709 (N_12709,N_11022,N_12213);
and U12710 (N_12710,N_12341,N_11331);
and U12711 (N_12711,N_11273,N_11968);
or U12712 (N_12712,N_9825,N_10213);
and U12713 (N_12713,N_12497,N_9988);
and U12714 (N_12714,N_10688,N_9948);
or U12715 (N_12715,N_10364,N_10177);
and U12716 (N_12716,N_10443,N_11116);
nor U12717 (N_12717,N_11818,N_9713);
or U12718 (N_12718,N_10898,N_11645);
or U12719 (N_12719,N_11350,N_10582);
nand U12720 (N_12720,N_12478,N_9486);
nand U12721 (N_12721,N_11999,N_11236);
or U12722 (N_12722,N_9432,N_11209);
or U12723 (N_12723,N_10869,N_9772);
and U12724 (N_12724,N_9677,N_12268);
and U12725 (N_12725,N_12082,N_10229);
or U12726 (N_12726,N_10209,N_11410);
or U12727 (N_12727,N_12111,N_10863);
or U12728 (N_12728,N_12228,N_11034);
or U12729 (N_12729,N_10493,N_10588);
or U12730 (N_12730,N_11789,N_10435);
nor U12731 (N_12731,N_9968,N_9750);
or U12732 (N_12732,N_9785,N_12458);
xor U12733 (N_12733,N_9835,N_10766);
nor U12734 (N_12734,N_9881,N_10769);
nand U12735 (N_12735,N_10890,N_12316);
or U12736 (N_12736,N_9714,N_10481);
or U12737 (N_12737,N_9940,N_12332);
or U12738 (N_12738,N_11950,N_10339);
xor U12739 (N_12739,N_11374,N_11757);
and U12740 (N_12740,N_11990,N_9502);
or U12741 (N_12741,N_11322,N_10152);
nor U12742 (N_12742,N_9488,N_9624);
or U12743 (N_12743,N_11778,N_11283);
nand U12744 (N_12744,N_10174,N_12069);
or U12745 (N_12745,N_9463,N_9384);
nor U12746 (N_12746,N_11184,N_11750);
or U12747 (N_12747,N_10867,N_12321);
nor U12748 (N_12748,N_9447,N_10170);
or U12749 (N_12749,N_10601,N_10985);
nor U12750 (N_12750,N_11911,N_11687);
xnor U12751 (N_12751,N_10982,N_11189);
nand U12752 (N_12752,N_11427,N_10559);
and U12753 (N_12753,N_10675,N_12091);
and U12754 (N_12754,N_9434,N_10775);
nand U12755 (N_12755,N_10477,N_12086);
nor U12756 (N_12756,N_10124,N_9871);
and U12757 (N_12757,N_11133,N_11715);
nand U12758 (N_12758,N_10102,N_10117);
nor U12759 (N_12759,N_12188,N_10613);
xor U12760 (N_12760,N_9655,N_10521);
nand U12761 (N_12761,N_11660,N_10511);
xor U12762 (N_12762,N_10508,N_11379);
nor U12763 (N_12763,N_11830,N_9937);
and U12764 (N_12764,N_10905,N_12073);
xor U12765 (N_12765,N_11369,N_9628);
nand U12766 (N_12766,N_11794,N_11237);
and U12767 (N_12767,N_10180,N_11129);
xor U12768 (N_12768,N_12094,N_10763);
or U12769 (N_12769,N_10246,N_10046);
nor U12770 (N_12770,N_11520,N_9813);
and U12771 (N_12771,N_11305,N_10127);
nand U12772 (N_12772,N_11970,N_11850);
and U12773 (N_12773,N_11325,N_11484);
nor U12774 (N_12774,N_10088,N_12189);
nand U12775 (N_12775,N_9416,N_10363);
nand U12776 (N_12776,N_12028,N_9559);
or U12777 (N_12777,N_11790,N_12357);
nand U12778 (N_12778,N_9757,N_10547);
nor U12779 (N_12779,N_9721,N_12354);
xor U12780 (N_12780,N_10810,N_11170);
nor U12781 (N_12781,N_9914,N_10397);
xor U12782 (N_12782,N_9863,N_9898);
or U12783 (N_12783,N_11992,N_10093);
nor U12784 (N_12784,N_10764,N_9431);
nand U12785 (N_12785,N_10200,N_11540);
and U12786 (N_12786,N_9665,N_11160);
nand U12787 (N_12787,N_11678,N_10522);
nand U12788 (N_12788,N_10008,N_12054);
nor U12789 (N_12789,N_12330,N_10251);
or U12790 (N_12790,N_9706,N_12447);
nand U12791 (N_12791,N_10715,N_9410);
or U12792 (N_12792,N_12026,N_10874);
or U12793 (N_12793,N_10674,N_9854);
nand U12794 (N_12794,N_10701,N_12470);
or U12795 (N_12795,N_10202,N_10669);
and U12796 (N_12796,N_11819,N_12008);
or U12797 (N_12797,N_10002,N_11550);
and U12798 (N_12798,N_10520,N_12249);
nand U12799 (N_12799,N_11613,N_12408);
and U12800 (N_12800,N_12019,N_9543);
and U12801 (N_12801,N_10835,N_11382);
nor U12802 (N_12802,N_12331,N_10228);
nor U12803 (N_12803,N_10767,N_9535);
or U12804 (N_12804,N_9975,N_11308);
or U12805 (N_12805,N_10990,N_10938);
nand U12806 (N_12806,N_12419,N_9738);
xor U12807 (N_12807,N_10311,N_10621);
xor U12808 (N_12808,N_12225,N_10646);
nand U12809 (N_12809,N_9523,N_11510);
and U12810 (N_12810,N_12348,N_10959);
or U12811 (N_12811,N_12083,N_10676);
or U12812 (N_12812,N_10257,N_10882);
nand U12813 (N_12813,N_9839,N_10942);
and U12814 (N_12814,N_11376,N_11777);
nor U12815 (N_12815,N_12048,N_10414);
or U12816 (N_12816,N_10892,N_9742);
and U12817 (N_12817,N_10195,N_10231);
nand U12818 (N_12818,N_10463,N_11203);
and U12819 (N_12819,N_12206,N_10222);
or U12820 (N_12820,N_9643,N_9892);
or U12821 (N_12821,N_12245,N_10987);
nand U12822 (N_12822,N_10575,N_9569);
nand U12823 (N_12823,N_10723,N_10537);
or U12824 (N_12824,N_9905,N_9970);
or U12825 (N_12825,N_12401,N_10750);
and U12826 (N_12826,N_11871,N_11647);
xor U12827 (N_12827,N_10451,N_10799);
nor U12828 (N_12828,N_12015,N_9944);
or U12829 (N_12829,N_10556,N_11942);
and U12830 (N_12830,N_12087,N_10554);
nor U12831 (N_12831,N_11492,N_12284);
or U12832 (N_12832,N_11727,N_9556);
nor U12833 (N_12833,N_11782,N_10977);
or U12834 (N_12834,N_9391,N_12492);
and U12835 (N_12835,N_9776,N_10057);
and U12836 (N_12836,N_10875,N_11612);
or U12837 (N_12837,N_11610,N_10703);
nor U12838 (N_12838,N_9705,N_11920);
or U12839 (N_12839,N_10315,N_9403);
nor U12840 (N_12840,N_11497,N_10568);
nor U12841 (N_12841,N_12381,N_12379);
nand U12842 (N_12842,N_11422,N_12431);
nand U12843 (N_12843,N_10078,N_11985);
nand U12844 (N_12844,N_10096,N_11921);
and U12845 (N_12845,N_12363,N_10221);
or U12846 (N_12846,N_11783,N_9642);
xnor U12847 (N_12847,N_10837,N_9806);
nor U12848 (N_12848,N_11558,N_12045);
nor U12849 (N_12849,N_12421,N_11000);
and U12850 (N_12850,N_9586,N_10995);
nor U12851 (N_12851,N_11027,N_11083);
nor U12852 (N_12852,N_10454,N_10060);
and U12853 (N_12853,N_9837,N_12449);
or U12854 (N_12854,N_10964,N_12117);
or U12855 (N_12855,N_11971,N_12385);
or U12856 (N_12856,N_12129,N_12179);
xor U12857 (N_12857,N_11373,N_9720);
or U12858 (N_12858,N_11989,N_12145);
xor U12859 (N_12859,N_11925,N_9389);
or U12860 (N_12860,N_10748,N_12214);
and U12861 (N_12861,N_9425,N_12405);
or U12862 (N_12862,N_12328,N_9497);
nor U12863 (N_12863,N_11766,N_10297);
xnor U12864 (N_12864,N_11402,N_11621);
nor U12865 (N_12865,N_10245,N_12282);
or U12866 (N_12866,N_10155,N_11952);
nor U12867 (N_12867,N_12059,N_11181);
nor U12868 (N_12868,N_9503,N_10774);
or U12869 (N_12869,N_11796,N_9507);
nor U12870 (N_12870,N_11330,N_12308);
and U12871 (N_12871,N_12063,N_11887);
nor U12872 (N_12872,N_11247,N_12425);
and U12873 (N_12873,N_12121,N_10687);
xor U12874 (N_12874,N_11634,N_10371);
and U12875 (N_12875,N_11442,N_11171);
nand U12876 (N_12876,N_11694,N_11380);
or U12877 (N_12877,N_11131,N_10834);
nor U12878 (N_12878,N_10166,N_9426);
or U12879 (N_12879,N_11085,N_9702);
xnor U12880 (N_12880,N_9927,N_9382);
or U12881 (N_12881,N_9693,N_9653);
nor U12882 (N_12882,N_11908,N_10474);
and U12883 (N_12883,N_11142,N_10845);
xnor U12884 (N_12884,N_11831,N_9999);
nor U12885 (N_12885,N_10334,N_10666);
nand U12886 (N_12886,N_10627,N_12234);
and U12887 (N_12887,N_11568,N_10446);
and U12888 (N_12888,N_9449,N_11980);
nand U12889 (N_12889,N_9788,N_11450);
and U12890 (N_12890,N_12383,N_11744);
nand U12891 (N_12891,N_9815,N_12485);
nor U12892 (N_12892,N_9614,N_12027);
nor U12893 (N_12893,N_12414,N_11826);
nor U12894 (N_12894,N_12312,N_10635);
nor U12895 (N_12895,N_10129,N_10939);
and U12896 (N_12896,N_11534,N_10941);
or U12897 (N_12897,N_11407,N_9967);
xor U12898 (N_12898,N_10495,N_9641);
and U12899 (N_12899,N_9795,N_10194);
and U12900 (N_12900,N_11225,N_10770);
and U12901 (N_12901,N_12068,N_10041);
nand U12902 (N_12902,N_9831,N_12152);
or U12903 (N_12903,N_11918,N_9593);
or U12904 (N_12904,N_9627,N_9958);
nand U12905 (N_12905,N_11065,N_11384);
xnor U12906 (N_12906,N_11845,N_9779);
or U12907 (N_12907,N_9879,N_12475);
nand U12908 (N_12908,N_9461,N_11155);
nor U12909 (N_12909,N_11656,N_12436);
xnor U12910 (N_12910,N_10673,N_12238);
nor U12911 (N_12911,N_9660,N_11892);
nand U12912 (N_12912,N_9878,N_9866);
nand U12913 (N_12913,N_9993,N_10104);
nor U12914 (N_12914,N_12099,N_10014);
or U12915 (N_12915,N_10657,N_10430);
nor U12916 (N_12916,N_10891,N_10050);
xor U12917 (N_12917,N_11938,N_10757);
and U12918 (N_12918,N_9524,N_11618);
nand U12919 (N_12919,N_10818,N_9471);
or U12920 (N_12920,N_10742,N_11272);
nand U12921 (N_12921,N_10310,N_10423);
nor U12922 (N_12922,N_11281,N_11791);
nor U12923 (N_12923,N_11249,N_9491);
nand U12924 (N_12924,N_10649,N_11418);
xnor U12925 (N_12925,N_11501,N_10126);
or U12926 (N_12926,N_11301,N_12373);
and U12927 (N_12927,N_10196,N_11199);
nand U12928 (N_12928,N_10026,N_11180);
xor U12929 (N_12929,N_12093,N_9682);
and U12930 (N_12930,N_11070,N_11696);
nor U12931 (N_12931,N_9792,N_11526);
or U12932 (N_12932,N_9902,N_11289);
or U12933 (N_12933,N_9895,N_12433);
and U12934 (N_12934,N_10617,N_9511);
nor U12935 (N_12935,N_11597,N_9689);
nor U12936 (N_12936,N_10868,N_10147);
and U12937 (N_12937,N_11683,N_9408);
nand U12938 (N_12938,N_11293,N_12277);
nand U12939 (N_12939,N_11313,N_11619);
nand U12940 (N_12940,N_11808,N_11220);
and U12941 (N_12941,N_11228,N_9758);
nand U12942 (N_12942,N_10418,N_11468);
nor U12943 (N_12943,N_10540,N_11833);
xor U12944 (N_12944,N_10261,N_9580);
nand U12945 (N_12945,N_10457,N_10543);
and U12946 (N_12946,N_10069,N_11728);
or U12947 (N_12947,N_11061,N_12420);
or U12948 (N_12948,N_11358,N_9687);
xnor U12949 (N_12949,N_10805,N_12166);
nor U12950 (N_12950,N_10011,N_9811);
or U12951 (N_12951,N_12173,N_12198);
nor U12952 (N_12952,N_12209,N_11663);
and U12953 (N_12953,N_10116,N_11726);
nor U12954 (N_12954,N_12102,N_11957);
nor U12955 (N_12955,N_10496,N_10136);
or U12956 (N_12956,N_11239,N_11344);
nor U12957 (N_12957,N_9563,N_9619);
nand U12958 (N_12958,N_10569,N_11486);
and U12959 (N_12959,N_10771,N_11177);
or U12960 (N_12960,N_10145,N_10074);
xnor U12961 (N_12961,N_10146,N_12378);
nor U12962 (N_12962,N_11425,N_10380);
nand U12963 (N_12963,N_11279,N_12266);
nor U12964 (N_12964,N_12413,N_11596);
nand U12965 (N_12965,N_11763,N_11895);
nand U12966 (N_12966,N_10937,N_10086);
nand U12967 (N_12967,N_9917,N_12324);
xor U12968 (N_12968,N_10439,N_11576);
or U12969 (N_12969,N_10047,N_10876);
nand U12970 (N_12970,N_11010,N_10856);
nand U12971 (N_12971,N_10105,N_9396);
or U12972 (N_12972,N_10720,N_10920);
and U12973 (N_12973,N_11589,N_10295);
xor U12974 (N_12974,N_10708,N_11885);
nand U12975 (N_12975,N_12071,N_11309);
or U12976 (N_12976,N_10304,N_12150);
and U12977 (N_12977,N_9756,N_10790);
or U12978 (N_12978,N_11069,N_12139);
xnor U12979 (N_12979,N_10563,N_12260);
or U12980 (N_12980,N_10156,N_10633);
and U12981 (N_12981,N_11196,N_10909);
xor U12982 (N_12982,N_12406,N_11742);
or U12983 (N_12983,N_9685,N_11521);
or U12984 (N_12984,N_9661,N_10097);
and U12985 (N_12985,N_11827,N_11310);
and U12986 (N_12986,N_10141,N_10515);
nand U12987 (N_12987,N_11847,N_9494);
nand U12988 (N_12988,N_12451,N_10753);
and U12989 (N_12989,N_10151,N_9672);
and U12990 (N_12990,N_10045,N_10901);
nor U12991 (N_12991,N_11463,N_12484);
xnor U12992 (N_12992,N_11424,N_11023);
nand U12993 (N_12993,N_11327,N_10500);
nand U12994 (N_12994,N_11775,N_11646);
nand U12995 (N_12995,N_9817,N_9430);
or U12996 (N_12996,N_10284,N_10839);
nand U12997 (N_12997,N_11263,N_12369);
or U12998 (N_12998,N_10357,N_10654);
and U12999 (N_12999,N_10210,N_9943);
or U13000 (N_13000,N_11452,N_9694);
nand U13001 (N_13001,N_11529,N_11730);
and U13002 (N_13002,N_9745,N_11076);
nor U13003 (N_13003,N_9626,N_9667);
and U13004 (N_13004,N_9629,N_12380);
or U13005 (N_13005,N_12356,N_12170);
nand U13006 (N_13006,N_11532,N_9664);
and U13007 (N_13007,N_10352,N_10504);
or U13008 (N_13008,N_9695,N_11685);
or U13009 (N_13009,N_11825,N_10855);
nand U13010 (N_13010,N_12488,N_10066);
or U13011 (N_13011,N_11686,N_10333);
xnor U13012 (N_13012,N_10042,N_10478);
nand U13013 (N_13013,N_11511,N_12432);
nand U13014 (N_13014,N_9558,N_9603);
nand U13015 (N_13015,N_10929,N_11176);
nor U13016 (N_13016,N_11984,N_9838);
and U13017 (N_13017,N_11873,N_12065);
xor U13018 (N_13018,N_11008,N_9395);
nand U13019 (N_13019,N_11435,N_12300);
nor U13020 (N_13020,N_10332,N_11130);
nor U13021 (N_13021,N_10075,N_11765);
and U13022 (N_13022,N_9674,N_11094);
nand U13023 (N_13023,N_12429,N_10090);
nand U13024 (N_13024,N_9956,N_11535);
or U13025 (N_13025,N_9512,N_11024);
or U13026 (N_13026,N_10943,N_9903);
nor U13027 (N_13027,N_12221,N_11752);
nor U13028 (N_13028,N_11525,N_12306);
and U13029 (N_13029,N_10727,N_10640);
or U13030 (N_13030,N_9822,N_10459);
xor U13031 (N_13031,N_11580,N_11716);
nand U13032 (N_13032,N_12314,N_12460);
or U13033 (N_13033,N_11025,N_11115);
nand U13034 (N_13034,N_10684,N_10239);
nand U13035 (N_13035,N_10927,N_11328);
nor U13036 (N_13036,N_10591,N_11933);
and U13037 (N_13037,N_11433,N_10536);
nand U13038 (N_13038,N_9969,N_12042);
or U13039 (N_13039,N_10587,N_11896);
and U13040 (N_13040,N_10662,N_10331);
nor U13041 (N_13041,N_11386,N_11552);
nor U13042 (N_13042,N_9820,N_11213);
nand U13043 (N_13043,N_9557,N_12066);
nand U13044 (N_13044,N_12146,N_12298);
nor U13045 (N_13045,N_9901,N_10605);
or U13046 (N_13046,N_12051,N_10513);
or U13047 (N_13047,N_9572,N_12041);
nand U13048 (N_13048,N_11640,N_9775);
nand U13049 (N_13049,N_11606,N_12143);
or U13050 (N_13050,N_11342,N_12455);
nand U13051 (N_13051,N_10624,N_11412);
nor U13052 (N_13052,N_10479,N_12329);
nor U13053 (N_13053,N_11187,N_10583);
and U13054 (N_13054,N_10482,N_10961);
or U13055 (N_13055,N_11588,N_9949);
or U13056 (N_13056,N_10670,N_10313);
and U13057 (N_13057,N_11876,N_11383);
or U13058 (N_13058,N_10094,N_10301);
and U13059 (N_13059,N_9584,N_11960);
nand U13060 (N_13060,N_9622,N_12386);
nand U13061 (N_13061,N_10338,N_9406);
or U13062 (N_13062,N_9681,N_11997);
xor U13063 (N_13063,N_11429,N_10039);
nor U13064 (N_13064,N_9452,N_9476);
nand U13065 (N_13065,N_11326,N_11729);
and U13066 (N_13066,N_9900,N_9960);
and U13067 (N_13067,N_11341,N_10160);
xnor U13068 (N_13068,N_11814,N_12409);
and U13069 (N_13069,N_12275,N_11100);
nor U13070 (N_13070,N_10277,N_10372);
nor U13071 (N_13071,N_12127,N_11666);
nand U13072 (N_13072,N_10472,N_10296);
nand U13073 (N_13073,N_11519,N_11291);
or U13074 (N_13074,N_10830,N_10342);
nor U13075 (N_13075,N_11844,N_10335);
xnor U13076 (N_13076,N_10467,N_11856);
nand U13077 (N_13077,N_10516,N_10663);
nor U13078 (N_13078,N_11210,N_11840);
nand U13079 (N_13079,N_11246,N_11504);
or U13080 (N_13080,N_11012,N_12365);
nor U13081 (N_13081,N_10400,N_11212);
nor U13082 (N_13082,N_9460,N_9441);
nand U13083 (N_13083,N_11630,N_12215);
nand U13084 (N_13084,N_9546,N_10490);
and U13085 (N_13085,N_10133,N_10458);
and U13086 (N_13086,N_11467,N_12362);
xor U13087 (N_13087,N_10610,N_10226);
nor U13088 (N_13088,N_10040,N_9676);
and U13089 (N_13089,N_9851,N_11564);
or U13090 (N_13090,N_10896,N_12443);
and U13091 (N_13091,N_11569,N_9884);
nand U13092 (N_13092,N_10316,N_11485);
nor U13093 (N_13093,N_10795,N_12169);
xor U13094 (N_13094,N_9793,N_11722);
nand U13095 (N_13095,N_10402,N_9636);
and U13096 (N_13096,N_10756,N_11855);
nor U13097 (N_13097,N_12347,N_11804);
nor U13098 (N_13098,N_11292,N_10801);
or U13099 (N_13099,N_11898,N_10029);
or U13100 (N_13100,N_11413,N_11409);
nor U13101 (N_13101,N_10546,N_12007);
or U13102 (N_13102,N_10322,N_11536);
and U13103 (N_13103,N_11458,N_10789);
nor U13104 (N_13104,N_11592,N_12261);
nor U13105 (N_13105,N_10109,N_10936);
nor U13106 (N_13106,N_12220,N_10054);
nand U13107 (N_13107,N_11616,N_10080);
or U13108 (N_13108,N_10437,N_11084);
nor U13109 (N_13109,N_12142,N_11821);
or U13110 (N_13110,N_9549,N_9703);
and U13111 (N_13111,N_11854,N_12430);
nor U13112 (N_13112,N_10053,N_10132);
or U13113 (N_13113,N_9930,N_9855);
and U13114 (N_13114,N_11150,N_11566);
and U13115 (N_13115,N_11426,N_10736);
nor U13116 (N_13116,N_12000,N_9615);
nand U13117 (N_13117,N_9730,N_11404);
and U13118 (N_13118,N_11378,N_11677);
nor U13119 (N_13119,N_9455,N_11533);
xor U13120 (N_13120,N_11072,N_11701);
nor U13121 (N_13121,N_10405,N_9561);
xor U13122 (N_13122,N_11500,N_9457);
nand U13123 (N_13123,N_10651,N_11068);
nor U13124 (N_13124,N_12452,N_11721);
nor U13125 (N_13125,N_10449,N_11679);
and U13126 (N_13126,N_11637,N_10207);
nor U13127 (N_13127,N_12165,N_11259);
and U13128 (N_13128,N_12040,N_9386);
xnor U13129 (N_13129,N_11352,N_9607);
and U13130 (N_13130,N_11353,N_10392);
or U13131 (N_13131,N_11432,N_9529);
and U13132 (N_13132,N_12162,N_12272);
nor U13133 (N_13133,N_12110,N_11417);
nand U13134 (N_13134,N_10824,N_10630);
and U13135 (N_13135,N_9597,N_11913);
nand U13136 (N_13136,N_10350,N_10632);
nor U13137 (N_13137,N_9711,N_12289);
nand U13138 (N_13138,N_11311,N_11234);
or U13139 (N_13139,N_10993,N_9848);
nand U13140 (N_13140,N_10388,N_11710);
and U13141 (N_13141,N_11319,N_10340);
nor U13142 (N_13142,N_9562,N_10643);
nand U13143 (N_13143,N_11581,N_10448);
or U13144 (N_13144,N_10879,N_10847);
nor U13145 (N_13145,N_11223,N_12210);
or U13146 (N_13146,N_9850,N_11611);
or U13147 (N_13147,N_11267,N_11470);
nor U13148 (N_13148,N_10428,N_11343);
xor U13149 (N_13149,N_9797,N_12052);
nand U13150 (N_13150,N_12311,N_11861);
or U13151 (N_13151,N_11949,N_10984);
nand U13152 (N_13152,N_12240,N_12095);
nand U13153 (N_13153,N_12391,N_10303);
nand U13154 (N_13154,N_10235,N_11423);
and U13155 (N_13155,N_12085,N_11784);
nand U13156 (N_13156,N_10754,N_12076);
nor U13157 (N_13157,N_11733,N_11649);
nor U13158 (N_13158,N_9663,N_10926);
nor U13159 (N_13159,N_11257,N_9805);
nor U13160 (N_13160,N_10809,N_11865);
and U13161 (N_13161,N_11389,N_12164);
nand U13162 (N_13162,N_11770,N_9809);
nand U13163 (N_13163,N_10385,N_9740);
xnor U13164 (N_13164,N_10211,N_10062);
and U13165 (N_13165,N_10487,N_12340);
nand U13166 (N_13166,N_9998,N_11922);
or U13167 (N_13167,N_10608,N_12360);
nand U13168 (N_13168,N_10408,N_10579);
and U13169 (N_13169,N_9852,N_11823);
and U13170 (N_13170,N_10051,N_11875);
or U13171 (N_13171,N_10220,N_11240);
nand U13172 (N_13172,N_11977,N_10759);
or U13173 (N_13173,N_10285,N_12046);
or U13174 (N_13174,N_10461,N_11221);
or U13175 (N_13175,N_11670,N_10996);
or U13176 (N_13176,N_11229,N_12403);
and U13177 (N_13177,N_12456,N_11780);
nand U13178 (N_13178,N_11307,N_10641);
or U13179 (N_13179,N_11186,N_12393);
and U13180 (N_13180,N_10225,N_12160);
and U13181 (N_13181,N_9466,N_12361);
nand U13182 (N_13182,N_9771,N_12376);
or U13183 (N_13183,N_10871,N_11127);
nor U13184 (N_13184,N_9737,N_10950);
and U13185 (N_13185,N_10665,N_10751);
nor U13186 (N_13186,N_10785,N_10282);
and U13187 (N_13187,N_10971,N_11090);
or U13188 (N_13188,N_10244,N_11233);
and U13189 (N_13189,N_10056,N_10735);
or U13190 (N_13190,N_11329,N_11909);
nand U13191 (N_13191,N_11680,N_10098);
nor U13192 (N_13192,N_11961,N_10888);
nor U13193 (N_13193,N_11208,N_12303);
and U13194 (N_13194,N_9582,N_9786);
nor U13195 (N_13195,N_10393,N_11011);
and U13196 (N_13196,N_10682,N_10150);
and U13197 (N_13197,N_10169,N_12029);
or U13198 (N_13198,N_10512,N_10119);
xnor U13199 (N_13199,N_9840,N_11141);
xnor U13200 (N_13200,N_10893,N_9440);
nor U13201 (N_13201,N_9525,N_9824);
nand U13202 (N_13202,N_9480,N_12353);
nand U13203 (N_13203,N_9617,N_11555);
and U13204 (N_13204,N_11642,N_10028);
nand U13205 (N_13205,N_10544,N_11154);
nor U13206 (N_13206,N_10243,N_12304);
and U13207 (N_13207,N_9893,N_11817);
nor U13208 (N_13208,N_11455,N_11849);
or U13209 (N_13209,N_12322,N_10324);
and U13210 (N_13210,N_10131,N_10404);
nand U13211 (N_13211,N_11900,N_10003);
and U13212 (N_13212,N_10252,N_9846);
nor U13213 (N_13213,N_10259,N_10308);
and U13214 (N_13214,N_12352,N_10212);
nand U13215 (N_13215,N_11912,N_12291);
xnor U13216 (N_13216,N_11682,N_11556);
nor U13217 (N_13217,N_11126,N_9621);
and U13218 (N_13218,N_11747,N_12355);
nor U13219 (N_13219,N_10356,N_11956);
nor U13220 (N_13220,N_11699,N_9808);
xnor U13221 (N_13221,N_10614,N_10672);
and U13222 (N_13222,N_9683,N_11522);
or U13223 (N_13223,N_10023,N_10576);
or U13224 (N_13224,N_10230,N_10833);
xor U13225 (N_13225,N_12226,N_9722);
nand U13226 (N_13226,N_10438,N_11347);
or U13227 (N_13227,N_11285,N_9550);
and U13228 (N_13228,N_11761,N_11146);
nor U13229 (N_13229,N_12192,N_10648);
and U13230 (N_13230,N_11060,N_11013);
nor U13231 (N_13231,N_11349,N_9759);
xnor U13232 (N_13232,N_11420,N_10859);
nand U13233 (N_13233,N_11943,N_9830);
nand U13234 (N_13234,N_12375,N_9911);
nand U13235 (N_13235,N_11917,N_10125);
or U13236 (N_13236,N_10578,N_11364);
nand U13237 (N_13237,N_11626,N_11518);
nor U13238 (N_13238,N_9924,N_12136);
or U13239 (N_13239,N_11809,N_10186);
nor U13240 (N_13240,N_12097,N_11490);
and U13241 (N_13241,N_10908,N_10218);
nand U13242 (N_13242,N_10647,N_11148);
and U13243 (N_13243,N_11207,N_10821);
nor U13244 (N_13244,N_9800,N_9918);
and U13245 (N_13245,N_11813,N_10148);
and U13246 (N_13246,N_9565,N_10658);
nand U13247 (N_13247,N_9541,N_11820);
or U13248 (N_13248,N_11639,N_10321);
and U13249 (N_13249,N_10242,N_10986);
nand U13250 (N_13250,N_11297,N_12123);
and U13251 (N_13251,N_11602,N_10860);
and U13252 (N_13252,N_11254,N_11713);
or U13253 (N_13253,N_12149,N_10997);
or U13254 (N_13254,N_11554,N_9456);
nor U13255 (N_13255,N_11946,N_11732);
nor U13256 (N_13256,N_10460,N_12122);
xnor U13257 (N_13257,N_10286,N_11758);
nor U13258 (N_13258,N_10700,N_10178);
and U13259 (N_13259,N_9843,N_12020);
and U13260 (N_13260,N_11062,N_11872);
nand U13261 (N_13261,N_9566,N_9791);
or U13262 (N_13262,N_10975,N_12398);
nor U13263 (N_13263,N_10925,N_9751);
nand U13264 (N_13264,N_10249,N_10827);
nor U13265 (N_13265,N_10717,N_11998);
and U13266 (N_13266,N_9913,N_10889);
xor U13267 (N_13267,N_10783,N_10841);
and U13268 (N_13268,N_11812,N_11966);
nand U13269 (N_13269,N_10525,N_9587);
or U13270 (N_13270,N_10498,N_12468);
nand U13271 (N_13271,N_10667,N_10616);
nor U13272 (N_13272,N_11355,N_10034);
nor U13273 (N_13273,N_11815,N_11250);
nand U13274 (N_13274,N_10919,N_11658);
or U13275 (N_13275,N_10044,N_11659);
and U13276 (N_13276,N_9530,N_9749);
and U13277 (N_13277,N_12471,N_11048);
nand U13278 (N_13278,N_12163,N_10274);
nor U13279 (N_13279,N_9487,N_10172);
nand U13280 (N_13280,N_10223,N_10192);
nor U13281 (N_13281,N_12131,N_10565);
nor U13282 (N_13282,N_12444,N_11945);
or U13283 (N_13283,N_9680,N_12474);
nand U13284 (N_13284,N_12009,N_11702);
or U13285 (N_13285,N_11400,N_9861);
xnor U13286 (N_13286,N_10038,N_12196);
nor U13287 (N_13287,N_9673,N_11414);
and U13288 (N_13288,N_10049,N_12014);
nor U13289 (N_13289,N_10031,N_10886);
nand U13290 (N_13290,N_9790,N_10526);
nand U13291 (N_13291,N_12239,N_9950);
nand U13292 (N_13292,N_9828,N_12124);
and U13293 (N_13293,N_12154,N_11502);
nand U13294 (N_13294,N_11979,N_11799);
or U13295 (N_13295,N_11138,N_11042);
xnor U13296 (N_13296,N_10885,N_10434);
and U13297 (N_13297,N_11738,N_9388);
nor U13298 (N_13298,N_9979,N_9666);
and U13299 (N_13299,N_10843,N_10947);
and U13300 (N_13300,N_10814,N_12473);
xnor U13301 (N_13301,N_10884,N_11862);
nor U13302 (N_13302,N_11864,N_11438);
nand U13303 (N_13303,N_10476,N_12050);
nand U13304 (N_13304,N_10382,N_11530);
and U13305 (N_13305,N_11545,N_12021);
or U13306 (N_13306,N_10163,N_11629);
nand U13307 (N_13307,N_10683,N_9767);
xnor U13308 (N_13308,N_12397,N_10265);
or U13309 (N_13309,N_11045,N_11785);
or U13310 (N_13310,N_11623,N_10615);
xor U13311 (N_13311,N_9485,N_9875);
and U13312 (N_13312,N_11149,N_11169);
or U13313 (N_13313,N_11446,N_12364);
or U13314 (N_13314,N_12463,N_12368);
or U13315 (N_13315,N_10505,N_9501);
nor U13316 (N_13316,N_11262,N_11829);
and U13317 (N_13317,N_11198,N_9980);
or U13318 (N_13318,N_9765,N_11857);
nor U13319 (N_13319,N_9746,N_9575);
xnor U13320 (N_13320,N_9577,N_12418);
or U13321 (N_13321,N_11764,N_12389);
nand U13322 (N_13322,N_12318,N_10918);
nor U13323 (N_13323,N_11360,N_12302);
and U13324 (N_13324,N_10595,N_11834);
and U13325 (N_13325,N_9704,N_10106);
nand U13326 (N_13326,N_11271,N_11551);
and U13327 (N_13327,N_11655,N_9594);
or U13328 (N_13328,N_10073,N_10741);
and U13329 (N_13329,N_9728,N_9964);
and U13330 (N_13330,N_10318,N_12211);
nor U13331 (N_13331,N_10915,N_10866);
xnor U13332 (N_13332,N_12180,N_9727);
nand U13333 (N_13333,N_10140,N_10275);
and U13334 (N_13334,N_10952,N_10572);
nor U13335 (N_13335,N_10597,N_9404);
and U13336 (N_13336,N_10416,N_9735);
nor U13337 (N_13337,N_11947,N_9915);
and U13338 (N_13338,N_11459,N_10897);
and U13339 (N_13339,N_12437,N_10954);
nand U13340 (N_13340,N_11491,N_9870);
or U13341 (N_13341,N_11570,N_10849);
nor U13342 (N_13342,N_10153,N_9929);
or U13343 (N_13343,N_11937,N_11393);
and U13344 (N_13344,N_9748,N_9847);
xnor U13345 (N_13345,N_9454,N_9649);
or U13346 (N_13346,N_9616,N_9780);
and U13347 (N_13347,N_11846,N_9400);
xor U13348 (N_13348,N_9648,N_9613);
xor U13349 (N_13349,N_10288,N_9783);
nor U13350 (N_13350,N_11381,N_11632);
nand U13351 (N_13351,N_9645,N_9862);
xnor U13352 (N_13352,N_11172,N_9470);
and U13353 (N_13353,N_9489,N_10699);
nand U13354 (N_13354,N_11103,N_11605);
xor U13355 (N_13355,N_9876,N_11361);
nand U13356 (N_13356,N_11962,N_9729);
or U13357 (N_13357,N_9731,N_9701);
or U13358 (N_13358,N_9668,N_10921);
nand U13359 (N_13359,N_10729,N_9521);
and U13360 (N_13360,N_11471,N_10969);
nand U13361 (N_13361,N_11388,N_11440);
or U13362 (N_13362,N_11884,N_10298);
and U13363 (N_13363,N_11137,N_10816);
nor U13364 (N_13364,N_10390,N_11222);
or U13365 (N_13365,N_9483,N_11671);
or U13366 (N_13366,N_10110,N_12295);
or U13367 (N_13367,N_11590,N_12278);
or U13368 (N_13368,N_11014,N_10365);
or U13369 (N_13369,N_10552,N_11870);
nor U13370 (N_13370,N_11401,N_11560);
nand U13371 (N_13371,N_10599,N_10972);
xor U13372 (N_13372,N_9662,N_11073);
xor U13373 (N_13373,N_10208,N_10524);
and U13374 (N_13374,N_10564,N_10378);
and U13375 (N_13375,N_12336,N_11681);
or U13376 (N_13376,N_12283,N_11883);
and U13377 (N_13377,N_11620,N_11190);
and U13378 (N_13378,N_10994,N_11321);
nand U13379 (N_13379,N_10535,N_12075);
nand U13380 (N_13380,N_9564,N_11899);
or U13381 (N_13381,N_10158,N_11508);
nor U13382 (N_13382,N_11695,N_12435);
or U13383 (N_13383,N_9973,N_12496);
nand U13384 (N_13384,N_11143,N_10916);
and U13385 (N_13385,N_11897,N_10983);
or U13386 (N_13386,N_10854,N_10637);
and U13387 (N_13387,N_12395,N_11910);
and U13388 (N_13388,N_9955,N_12002);
and U13389 (N_13389,N_10258,N_12477);
nor U13390 (N_13390,N_12147,N_10722);
and U13391 (N_13391,N_11323,N_10844);
nand U13392 (N_13392,N_11227,N_9467);
nor U13393 (N_13393,N_11673,N_11351);
and U13394 (N_13394,N_11274,N_12037);
and U13395 (N_13395,N_10555,N_11561);
and U13396 (N_13396,N_11755,N_10998);
or U13397 (N_13397,N_9536,N_11050);
nand U13398 (N_13398,N_10489,N_11838);
nand U13399 (N_13399,N_9446,N_9378);
or U13400 (N_13400,N_11454,N_11652);
or U13401 (N_13401,N_11926,N_10396);
or U13402 (N_13402,N_10716,N_10592);
or U13403 (N_13403,N_12372,N_10181);
or U13404 (N_13404,N_10409,N_11863);
or U13405 (N_13405,N_10622,N_11599);
or U13406 (N_13406,N_10175,N_11265);
nor U13407 (N_13407,N_10401,N_10410);
and U13408 (N_13408,N_12004,N_11802);
and U13409 (N_13409,N_11295,N_12168);
nor U13410 (N_13410,N_11163,N_11097);
xor U13411 (N_13411,N_12229,N_11041);
nand U13412 (N_13412,N_10973,N_10858);
xor U13413 (N_13413,N_11959,N_11803);
nor U13414 (N_13414,N_10585,N_11004);
nor U13415 (N_13415,N_12081,N_10111);
nand U13416 (N_13416,N_11625,N_11916);
nor U13417 (N_13417,N_9818,N_10179);
nand U13418 (N_13418,N_11537,N_11235);
nor U13419 (N_13419,N_11859,N_11447);
nand U13420 (N_13420,N_11436,N_10671);
and U13421 (N_13421,N_11754,N_10822);
nand U13422 (N_13422,N_10645,N_11527);
nor U13423 (N_13423,N_11314,N_11167);
or U13424 (N_13424,N_10214,N_11981);
or U13425 (N_13425,N_12130,N_11256);
or U13426 (N_13426,N_9474,N_11587);
nor U13427 (N_13427,N_11547,N_10018);
and U13428 (N_13428,N_12001,N_9916);
nor U13429 (N_13429,N_12003,N_10353);
nand U13430 (N_13430,N_10082,N_11919);
nand U13431 (N_13431,N_10114,N_9849);
nand U13432 (N_13432,N_9595,N_12319);
nand U13433 (N_13433,N_11306,N_11978);
and U13434 (N_13434,N_10653,N_10101);
or U13435 (N_13435,N_11302,N_9640);
and U13436 (N_13436,N_11219,N_12011);
nor U13437 (N_13437,N_11553,N_11690);
or U13438 (N_13438,N_10527,N_11567);
nor U13439 (N_13439,N_12106,N_11851);
nand U13440 (N_13440,N_9864,N_10948);
nor U13441 (N_13441,N_10502,N_12344);
nand U13442 (N_13442,N_11517,N_11902);
and U13443 (N_13443,N_10387,N_10907);
nand U13444 (N_13444,N_11595,N_9571);
or U13445 (N_13445,N_12195,N_11122);
xnor U13446 (N_13446,N_11264,N_10328);
nand U13447 (N_13447,N_12273,N_9639);
and U13448 (N_13448,N_9734,N_9724);
nand U13449 (N_13449,N_11266,N_10032);
nand U13450 (N_13450,N_9885,N_11044);
nor U13451 (N_13451,N_11839,N_12416);
nor U13452 (N_13452,N_11403,N_9414);
nor U13453 (N_13453,N_12193,N_11969);
nand U13454 (N_13454,N_12104,N_10326);
or U13455 (N_13455,N_11585,N_11665);
and U13456 (N_13456,N_9996,N_12114);
nand U13457 (N_13457,N_10197,N_9574);
and U13458 (N_13458,N_11858,N_10035);
nor U13459 (N_13459,N_9669,N_10375);
nand U13460 (N_13460,N_11739,N_10253);
nand U13461 (N_13461,N_9464,N_12481);
or U13462 (N_13462,N_9744,N_10475);
nor U13463 (N_13463,N_11816,N_9510);
nand U13464 (N_13464,N_9514,N_9784);
nand U13465 (N_13465,N_11015,N_11542);
or U13466 (N_13466,N_12017,N_12320);
or U13467 (N_13467,N_10260,N_11725);
and U13468 (N_13468,N_10266,N_11304);
or U13469 (N_13469,N_10580,N_10019);
nand U13470 (N_13470,N_11092,N_9609);
and U13471 (N_13471,N_10427,N_11516);
nor U13472 (N_13472,N_10491,N_11445);
and U13473 (N_13473,N_9428,N_11194);
nand U13474 (N_13474,N_10903,N_10823);
nor U13475 (N_13475,N_10740,N_12138);
or U13476 (N_13476,N_9690,N_12285);
or U13477 (N_13477,N_10215,N_10188);
nor U13478 (N_13478,N_11493,N_12126);
and U13479 (N_13479,N_10660,N_12370);
and U13480 (N_13480,N_11786,N_12445);
or U13481 (N_13481,N_11111,N_12055);
or U13482 (N_13482,N_10545,N_11443);
nor U13483 (N_13483,N_11835,N_10001);
or U13484 (N_13484,N_12313,N_12483);
xnor U13485 (N_13485,N_12388,N_9606);
and U13486 (N_13486,N_11200,N_12161);
nor U13487 (N_13487,N_10747,N_9570);
xnor U13488 (N_13488,N_10190,N_9994);
xor U13489 (N_13489,N_11598,N_11058);
nand U13490 (N_13490,N_10273,N_9528);
nor U13491 (N_13491,N_10444,N_10037);
and U13492 (N_13492,N_10933,N_9781);
nand U13493 (N_13493,N_9987,N_11193);
nand U13494 (N_13494,N_10928,N_9755);
nor U13495 (N_13495,N_11852,N_10571);
nor U13496 (N_13496,N_11523,N_9646);
and U13497 (N_13497,N_11482,N_9686);
nor U13498 (N_13498,N_9753,N_12335);
nor U13499 (N_13499,N_9763,N_9610);
nor U13500 (N_13500,N_12338,N_10108);
nand U13501 (N_13501,N_10182,N_11481);
or U13502 (N_13502,N_10623,N_10704);
nor U13503 (N_13503,N_12013,N_11415);
nand U13504 (N_13504,N_10447,N_10294);
and U13505 (N_13505,N_10256,N_11277);
and U13506 (N_13506,N_10497,N_9991);
nand U13507 (N_13507,N_10711,N_9379);
or U13508 (N_13508,N_10021,N_11105);
nor U13509 (N_13509,N_10091,N_10238);
nor U13510 (N_13510,N_11345,N_9981);
nor U13511 (N_13511,N_11367,N_9962);
nand U13512 (N_13512,N_9419,N_10123);
or U13513 (N_13513,N_9789,N_10425);
or U13514 (N_13514,N_12349,N_10306);
and U13515 (N_13515,N_10930,N_11792);
nor U13516 (N_13516,N_11650,N_11505);
nand U13517 (N_13517,N_12157,N_11009);
or U13518 (N_13518,N_10689,N_11182);
or U13519 (N_13519,N_12427,N_9585);
or U13520 (N_13520,N_11120,N_11366);
or U13521 (N_13521,N_10980,N_10731);
nor U13522 (N_13522,N_10370,N_12208);
or U13523 (N_13523,N_11252,N_9773);
or U13524 (N_13524,N_12202,N_11215);
nand U13525 (N_13525,N_10659,N_11033);
nand U13526 (N_13526,N_11132,N_11166);
or U13527 (N_13527,N_11080,N_11269);
and U13528 (N_13528,N_12175,N_10144);
xor U13529 (N_13529,N_12345,N_10738);
nor U13530 (N_13530,N_10872,N_12257);
or U13531 (N_13531,N_10059,N_11489);
and U13532 (N_13532,N_12176,N_10022);
nand U13533 (N_13533,N_10441,N_11276);
nor U13534 (N_13534,N_11867,N_11192);
nor U13535 (N_13535,N_10529,N_11615);
or U13536 (N_13536,N_11574,N_11691);
nand U13537 (N_13537,N_11356,N_10573);
nor U13538 (N_13538,N_9954,N_11066);
xor U13539 (N_13539,N_12394,N_11591);
nand U13540 (N_13540,N_11774,N_11603);
xor U13541 (N_13541,N_12390,N_9907);
nor U13542 (N_13542,N_9493,N_10358);
and U13543 (N_13543,N_12186,N_11441);
or U13544 (N_13544,N_11017,N_10112);
or U13545 (N_13545,N_12156,N_10033);
nor U13546 (N_13546,N_9620,N_12438);
or U13547 (N_13547,N_10781,N_11096);
xnor U13548 (N_13548,N_10612,N_9551);
nor U13549 (N_13549,N_11736,N_11932);
or U13550 (N_13550,N_11411,N_11806);
or U13551 (N_13551,N_10531,N_12158);
nor U13552 (N_13552,N_11218,N_11688);
nor U13553 (N_13553,N_12084,N_11751);
nand U13554 (N_13554,N_12231,N_9983);
and U13555 (N_13555,N_10887,N_11807);
nor U13556 (N_13556,N_11340,N_11993);
nor U13557 (N_13557,N_11572,N_11941);
nor U13558 (N_13558,N_9633,N_10462);
nand U13559 (N_13559,N_9804,N_11515);
xnor U13560 (N_13560,N_12441,N_11390);
or U13561 (N_13561,N_11052,N_11147);
xor U13562 (N_13562,N_11251,N_11579);
or U13563 (N_13563,N_10198,N_10343);
nand U13564 (N_13564,N_10368,N_10271);
or U13565 (N_13565,N_10436,N_11986);
or U13566 (N_13566,N_10912,N_11955);
xor U13567 (N_13567,N_10415,N_10749);
nand U13568 (N_13568,N_10831,N_11363);
nor U13569 (N_13569,N_9696,N_11473);
xnor U13570 (N_13570,N_9401,N_11769);
and U13571 (N_13571,N_12410,N_11475);
and U13572 (N_13572,N_11333,N_10233);
nor U13573 (N_13573,N_9402,N_11800);
xnor U13574 (N_13574,N_10386,N_11020);
nor U13575 (N_13575,N_12294,N_10728);
and U13576 (N_13576,N_9513,N_10176);
nor U13577 (N_13577,N_10618,N_10577);
xor U13578 (N_13578,N_11419,N_10154);
nand U13579 (N_13579,N_9910,N_9623);
and U13580 (N_13580,N_12265,N_12101);
or U13581 (N_13581,N_10165,N_9675);
nand U13582 (N_13582,N_11205,N_10381);
xor U13583 (N_13583,N_12279,N_10562);
and U13584 (N_13584,N_11717,N_12047);
xnor U13585 (N_13585,N_10232,N_10162);
nor U13586 (N_13586,N_9592,N_9770);
nand U13587 (N_13587,N_11824,N_10911);
or U13588 (N_13588,N_11243,N_10219);
nor U13589 (N_13589,N_11748,N_12058);
and U13590 (N_13590,N_12434,N_9832);
nor U13591 (N_13591,N_10417,N_12199);
and U13592 (N_13592,N_12116,N_10362);
and U13593 (N_13593,N_9782,N_10706);
or U13594 (N_13594,N_10185,N_10829);
or U13595 (N_13595,N_11641,N_9448);
nand U13596 (N_13596,N_9932,N_11805);
and U13597 (N_13597,N_9919,N_9553);
nor U13598 (N_13598,N_12251,N_10714);
xor U13599 (N_13599,N_11669,N_10115);
and U13600 (N_13600,N_11035,N_9886);
or U13601 (N_13601,N_12367,N_11538);
nor U13602 (N_13602,N_10752,N_12299);
xnor U13603 (N_13603,N_11346,N_11718);
nor U13604 (N_13604,N_12462,N_11091);
or U13605 (N_13605,N_11206,N_12264);
xnor U13606 (N_13606,N_11931,N_9890);
or U13607 (N_13607,N_12197,N_11334);
or U13608 (N_13608,N_12337,N_11661);
or U13609 (N_13609,N_9482,N_11627);
nand U13610 (N_13610,N_11101,N_11430);
nand U13611 (N_13611,N_10782,N_9634);
or U13612 (N_13612,N_9588,N_10606);
and U13613 (N_13613,N_11299,N_9459);
and U13614 (N_13614,N_10187,N_12402);
nand U13615 (N_13615,N_11723,N_10857);
nand U13616 (N_13616,N_9599,N_11544);
and U13617 (N_13617,N_9544,N_9933);
and U13618 (N_13618,N_12467,N_9802);
nor U13619 (N_13619,N_11179,N_11705);
nand U13620 (N_13620,N_12358,N_11038);
nor U13621 (N_13621,N_11514,N_9518);
and U13622 (N_13622,N_10692,N_9691);
nand U13623 (N_13623,N_10394,N_12480);
or U13624 (N_13624,N_10530,N_10628);
xor U13625 (N_13625,N_12218,N_11202);
xor U13626 (N_13626,N_10914,N_11745);
nand U13627 (N_13627,N_10013,N_11543);
nand U13628 (N_13628,N_12310,N_10067);
nor U13629 (N_13629,N_11280,N_9604);
nor U13630 (N_13630,N_11600,N_11546);
or U13631 (N_13631,N_10777,N_12466);
or U13632 (N_13632,N_9537,N_10548);
nand U13633 (N_13633,N_9853,N_10776);
nand U13634 (N_13634,N_11461,N_11370);
and U13635 (N_13635,N_11029,N_9953);
or U13636 (N_13636,N_11609,N_12323);
xnor U13637 (N_13637,N_12227,N_11622);
or U13638 (N_13638,N_10725,N_11336);
and U13639 (N_13639,N_10745,N_11031);
nor U13640 (N_13640,N_9679,N_11244);
nor U13641 (N_13641,N_10746,N_12476);
and U13642 (N_13642,N_10946,N_11275);
nor U13643 (N_13643,N_11936,N_11288);
and U13644 (N_13644,N_10280,N_9436);
or U13645 (N_13645,N_12450,N_11653);
and U13646 (N_13646,N_10267,N_12342);
and U13647 (N_13647,N_11081,N_12118);
nand U13648 (N_13648,N_11689,N_11136);
nor U13649 (N_13649,N_11434,N_11159);
xnor U13650 (N_13650,N_11811,N_11107);
nor U13651 (N_13651,N_11562,N_10081);
and U13652 (N_13652,N_12236,N_11298);
or U13653 (N_13653,N_11506,N_10802);
xnor U13654 (N_13654,N_10607,N_12060);
or U13655 (N_13655,N_10992,N_9925);
or U13656 (N_13656,N_10832,N_9904);
nor U13657 (N_13657,N_10456,N_9612);
xnor U13658 (N_13658,N_11387,N_11915);
nor U13659 (N_13659,N_10686,N_10203);
or U13660 (N_13660,N_11934,N_10680);
xnor U13661 (N_13661,N_10999,N_9761);
xnor U13662 (N_13662,N_11879,N_11878);
nand U13663 (N_13663,N_10589,N_10509);
nand U13664 (N_13664,N_11211,N_10312);
or U13665 (N_13665,N_9437,N_12033);
nor U13666 (N_13666,N_10945,N_10744);
or U13667 (N_13667,N_10346,N_12064);
nor U13668 (N_13668,N_10724,N_11448);
and U13669 (N_13669,N_9547,N_9986);
or U13670 (N_13670,N_9533,N_9405);
nand U13671 (N_13671,N_10811,N_11907);
and U13672 (N_13672,N_11232,N_11953);
xor U13673 (N_13673,N_11201,N_10292);
nand U13674 (N_13674,N_11557,N_11513);
nand U13675 (N_13675,N_12495,N_11396);
nand U13676 (N_13676,N_12103,N_11735);
nor U13677 (N_13677,N_10005,N_11617);
and U13678 (N_13678,N_9596,N_10934);
nand U13679 (N_13679,N_10345,N_10399);
or U13680 (N_13680,N_10058,N_11714);
nor U13681 (N_13681,N_9520,N_9718);
nor U13682 (N_13682,N_10466,N_12024);
or U13683 (N_13683,N_12174,N_11948);
or U13684 (N_13684,N_10120,N_10634);
nand U13685 (N_13685,N_11577,N_9590);
and U13686 (N_13686,N_10639,N_10566);
or U13687 (N_13687,N_11317,N_12109);
nand U13688 (N_13688,N_10626,N_10118);
nand U13689 (N_13689,N_9637,N_11204);
or U13690 (N_13690,N_10157,N_11054);
nor U13691 (N_13691,N_10278,N_10279);
xnor U13692 (N_13692,N_10836,N_11028);
or U13693 (N_13693,N_11093,N_12190);
nor U13694 (N_13694,N_11158,N_11756);
xor U13695 (N_13695,N_12062,N_9539);
and U13696 (N_13696,N_9869,N_11416);
xnor U13697 (N_13697,N_11983,N_9732);
and U13698 (N_13698,N_11128,N_10848);
or U13699 (N_13699,N_10063,N_11762);
nor U13700 (N_13700,N_9422,N_10344);
nand U13701 (N_13701,N_11498,N_10944);
or U13702 (N_13702,N_10931,N_11287);
nor U13703 (N_13703,N_12350,N_12039);
or U13704 (N_13704,N_11923,N_11499);
and U13705 (N_13705,N_10354,N_9894);
nand U13706 (N_13706,N_11399,N_11586);
nand U13707 (N_13707,N_11318,N_10861);
nor U13708 (N_13708,N_11929,N_10270);
and U13709 (N_13709,N_11368,N_10164);
and U13710 (N_13710,N_11260,N_11007);
xor U13711 (N_13711,N_10955,N_11593);
or U13712 (N_13712,N_11282,N_10968);
nand U13713 (N_13713,N_9411,N_9716);
xnor U13714 (N_13714,N_9965,N_11893);
nand U13715 (N_13715,N_10935,N_12482);
xnor U13716 (N_13716,N_12005,N_11077);
nand U13717 (N_13717,N_9801,N_11882);
and U13718 (N_13718,N_11214,N_10237);
xnor U13719 (N_13719,N_11793,N_10650);
or U13720 (N_13720,N_10574,N_11848);
or U13721 (N_13721,N_9891,N_10199);
and U13722 (N_13722,N_10429,N_10932);
nor U13723 (N_13723,N_10486,N_9527);
nor U13724 (N_13724,N_10594,N_10904);
or U13725 (N_13725,N_9498,N_9469);
and U13726 (N_13726,N_9888,N_10142);
or U13727 (N_13727,N_12185,N_9816);
nor U13728 (N_13728,N_9992,N_11003);
xnor U13729 (N_13729,N_10619,N_11134);
nor U13730 (N_13730,N_9699,N_11675);
xnor U13731 (N_13731,N_11664,N_9576);
nor U13732 (N_13732,N_10264,N_11479);
nor U13733 (N_13733,N_9380,N_10963);
xor U13734 (N_13734,N_9630,N_10604);
nand U13735 (N_13735,N_11951,N_11074);
nand U13736 (N_13736,N_10287,N_10922);
or U13737 (N_13737,N_9700,N_9984);
nor U13738 (N_13738,N_12077,N_11183);
or U13739 (N_13739,N_11371,N_10743);
or U13740 (N_13740,N_9458,N_9573);
and U13741 (N_13741,N_10570,N_10168);
xnor U13742 (N_13742,N_11868,N_11255);
nor U13743 (N_13743,N_9896,N_10442);
or U13744 (N_13744,N_10283,N_9555);
nor U13745 (N_13745,N_11480,N_9868);
or U13746 (N_13746,N_12281,N_12422);
nor U13747 (N_13747,N_11954,N_9478);
nor U13748 (N_13748,N_9670,N_11559);
nand U13749 (N_13749,N_11106,N_11055);
or U13750 (N_13750,N_12096,N_10254);
and U13751 (N_13751,N_12343,N_10241);
nand U13752 (N_13752,N_10317,N_11124);
nor U13753 (N_13753,N_12377,N_10620);
and U13754 (N_13754,N_10788,N_9484);
or U13755 (N_13755,N_11935,N_10655);
nor U13756 (N_13756,N_10083,N_11563);
or U13757 (N_13757,N_10693,N_10431);
nand U13758 (N_13758,N_11853,N_9873);
or U13759 (N_13759,N_10825,N_10507);
nand U13760 (N_13760,N_12100,N_10320);
and U13761 (N_13761,N_9923,N_9375);
xnor U13762 (N_13762,N_12222,N_9654);
or U13763 (N_13763,N_10798,N_11582);
and U13764 (N_13764,N_10193,N_11078);
and U13765 (N_13765,N_10085,N_10691);
or U13766 (N_13766,N_9803,N_11315);
or U13767 (N_13767,N_12274,N_10263);
and U13768 (N_13768,N_12159,N_12287);
and U13769 (N_13769,N_10598,N_11667);
nor U13770 (N_13770,N_10424,N_11469);
and U13771 (N_13771,N_10347,N_11135);
xor U13772 (N_13772,N_11286,N_9747);
and U13773 (N_13773,N_11165,N_10262);
and U13774 (N_13774,N_11474,N_9951);
or U13775 (N_13775,N_11444,N_10329);
xnor U13776 (N_13776,N_11335,N_12088);
xor U13777 (N_13777,N_9542,N_11974);
and U13778 (N_13778,N_9500,N_10503);
and U13779 (N_13779,N_9435,N_11608);
or U13780 (N_13780,N_10084,N_10550);
and U13781 (N_13781,N_10593,N_10690);
nand U13782 (N_13782,N_12280,N_11037);
nand U13783 (N_13783,N_12366,N_11903);
nor U13784 (N_13784,N_10733,N_9823);
nand U13785 (N_13785,N_12070,N_11828);
xor U13786 (N_13786,N_11261,N_12057);
nand U13787 (N_13787,N_10979,N_10293);
and U13788 (N_13788,N_9532,N_9810);
or U13789 (N_13789,N_11405,N_11797);
and U13790 (N_13790,N_11768,N_10072);
and U13791 (N_13791,N_12479,N_10323);
or U13792 (N_13792,N_9989,N_10806);
nand U13793 (N_13793,N_11457,N_11643);
xnor U13794 (N_13794,N_11312,N_11633);
or U13795 (N_13795,N_11217,N_10450);
nor U13796 (N_13796,N_10079,N_11332);
and U13797 (N_13797,N_9897,N_9719);
nand U13798 (N_13798,N_10468,N_12074);
nand U13799 (N_13799,N_10377,N_12464);
or U13800 (N_13800,N_11578,N_10586);
and U13801 (N_13801,N_9926,N_10596);
or U13802 (N_13802,N_9709,N_10227);
nor U13803 (N_13803,N_11512,N_10445);
and U13804 (N_13804,N_12035,N_12232);
nand U13805 (N_13805,N_12030,N_9540);
nand U13806 (N_13806,N_10533,N_10600);
or U13807 (N_13807,N_10403,N_10518);
nor U13808 (N_13808,N_10036,N_11973);
xnor U13809 (N_13809,N_11740,N_10426);
and U13810 (N_13810,N_9393,N_11760);
nand U13811 (N_13811,N_10707,N_12461);
nand U13812 (N_13812,N_11684,N_12105);
or U13813 (N_13813,N_11703,N_11112);
nor U13814 (N_13814,N_11781,N_10652);
and U13815 (N_13815,N_10016,N_10236);
nor U13816 (N_13816,N_9638,N_10678);
or U13817 (N_13817,N_9909,N_10234);
xor U13818 (N_13818,N_12171,N_10924);
nor U13819 (N_13819,N_11594,N_9581);
nor U13820 (N_13820,N_10314,N_9921);
nand U13821 (N_13821,N_12223,N_10581);
nor U13822 (N_13822,N_11881,N_11734);
xnor U13823 (N_13823,N_9515,N_11406);
xnor U13824 (N_13824,N_9534,N_12194);
and U13825 (N_13825,N_12119,N_11039);
nor U13826 (N_13826,N_12315,N_11303);
and U13827 (N_13827,N_12203,N_12216);
nand U13828 (N_13828,N_10465,N_11421);
or U13829 (N_13829,N_12457,N_10558);
or U13830 (N_13830,N_10807,N_12181);
nor U13831 (N_13831,N_11049,N_9799);
nand U13832 (N_13832,N_11088,N_10276);
nand U13833 (N_13833,N_10138,N_12250);
and U13834 (N_13834,N_11967,N_10012);
or U13835 (N_13835,N_11338,N_12493);
or U13836 (N_13836,N_10787,N_9506);
or U13837 (N_13837,N_10910,N_11724);
nor U13838 (N_13838,N_10464,N_12334);
and U13839 (N_13839,N_11431,N_9509);
and U13840 (N_13840,N_9961,N_10800);
or U13841 (N_13841,N_9796,N_10248);
xnor U13842 (N_13842,N_9941,N_10389);
nor U13843 (N_13843,N_11296,N_9445);
or U13844 (N_13844,N_10341,N_10092);
nand U13845 (N_13845,N_11843,N_10065);
nor U13846 (N_13846,N_12056,N_11749);
or U13847 (N_13847,N_12010,N_12230);
xnor U13848 (N_13848,N_11157,N_9625);
nor U13849 (N_13849,N_11676,N_12200);
and U13850 (N_13850,N_11162,N_11928);
nand U13851 (N_13851,N_11099,N_11002);
nand U13852 (N_13852,N_10488,N_9971);
nor U13853 (N_13853,N_9922,N_11996);
and U13854 (N_13854,N_11339,N_9814);
xor U13855 (N_13855,N_10319,N_10523);
xnor U13856 (N_13856,N_12254,N_11624);
nand U13857 (N_13857,N_9377,N_11801);
nand U13858 (N_13858,N_11654,N_10070);
or U13859 (N_13859,N_12133,N_11230);
nor U13860 (N_13860,N_10189,N_12078);
xor U13861 (N_13861,N_11604,N_12442);
nand U13862 (N_13862,N_10071,N_12089);
or U13863 (N_13863,N_10191,N_12448);
nand U13864 (N_13864,N_9598,N_10149);
or U13865 (N_13865,N_9985,N_9635);
and U13866 (N_13866,N_10917,N_9656);
and U13867 (N_13867,N_10128,N_11583);
nand U13868 (N_13868,N_12407,N_10103);
or U13869 (N_13869,N_9465,N_12469);
or U13870 (N_13870,N_12293,N_11394);
xnor U13871 (N_13871,N_9708,N_10528);
nand U13872 (N_13872,N_9872,N_11528);
nor U13873 (N_13873,N_11772,N_11119);
and U13874 (N_13874,N_10560,N_11465);
nand U13875 (N_13875,N_11253,N_11651);
nor U13876 (N_13876,N_11001,N_10779);
nand U13877 (N_13877,N_10484,N_10470);
nor U13878 (N_13878,N_11365,N_12382);
and U13879 (N_13879,N_9652,N_11635);
xor U13880 (N_13880,N_10718,N_9959);
xor U13881 (N_13881,N_11113,N_11964);
or U13882 (N_13882,N_11242,N_11462);
nor U13883 (N_13883,N_9583,N_10730);
and U13884 (N_13884,N_11021,N_9522);
and U13885 (N_13885,N_10240,N_10638);
and U13886 (N_13886,N_9468,N_12098);
nand U13887 (N_13887,N_12396,N_11075);
and U13888 (N_13888,N_10030,N_9397);
nand U13889 (N_13889,N_11767,N_10391);
and U13890 (N_13890,N_11662,N_9398);
and U13891 (N_13891,N_11975,N_11053);
nor U13892 (N_13892,N_10373,N_10184);
and U13893 (N_13893,N_9741,N_10603);
nand U13894 (N_13894,N_9857,N_11300);
nand U13895 (N_13895,N_9413,N_11503);
and U13896 (N_13896,N_12307,N_9591);
and U13897 (N_13897,N_10768,N_9418);
or U13898 (N_13898,N_10631,N_10369);
or U13899 (N_13899,N_10161,N_11477);
nor U13900 (N_13900,N_12207,N_9717);
nor U13901 (N_13901,N_11478,N_9726);
or U13902 (N_13902,N_11737,N_9381);
nand U13903 (N_13903,N_9412,N_9710);
or U13904 (N_13904,N_12137,N_11005);
nand U13905 (N_13905,N_9505,N_11692);
nor U13906 (N_13906,N_11019,N_9912);
nor U13907 (N_13907,N_12201,N_12072);
and U13908 (N_13908,N_11759,N_12237);
nor U13909 (N_13909,N_9725,N_10007);
and U13910 (N_13910,N_10325,N_10894);
nor U13911 (N_13911,N_9611,N_11016);
nor U13912 (N_13912,N_11437,N_10452);
or U13913 (N_13913,N_9845,N_12067);
xnor U13914 (N_13914,N_9552,N_11888);
nand U13915 (N_13915,N_12012,N_9982);
or U13916 (N_13916,N_9632,N_10681);
nand U13917 (N_13917,N_9421,N_11428);
or U13918 (N_13918,N_10773,N_9972);
or U13919 (N_13919,N_9589,N_12092);
or U13920 (N_13920,N_9712,N_11746);
or U13921 (N_13921,N_10953,N_9974);
nand U13922 (N_13922,N_9516,N_9427);
xor U13923 (N_13923,N_10989,N_11357);
and U13924 (N_13924,N_10432,N_12248);
xor U13925 (N_13925,N_10794,N_12286);
or U13926 (N_13926,N_10553,N_11487);
and U13927 (N_13927,N_12141,N_10851);
or U13928 (N_13928,N_12247,N_11391);
xnor U13929 (N_13929,N_11117,N_10017);
nor U13930 (N_13930,N_9692,N_10006);
or U13931 (N_13931,N_9707,N_12267);
or U13932 (N_13932,N_10159,N_10967);
nand U13933 (N_13933,N_10514,N_11700);
or U13934 (N_13934,N_11614,N_9844);
xor U13935 (N_13935,N_12080,N_9579);
nand U13936 (N_13936,N_12023,N_12090);
and U13937 (N_13937,N_9947,N_10913);
xor U13938 (N_13938,N_10862,N_11395);
and U13939 (N_13939,N_10813,N_9697);
nor U13940 (N_13940,N_11238,N_12263);
nand U13941 (N_13941,N_11822,N_12489);
and U13942 (N_13942,N_9492,N_9883);
and U13943 (N_13943,N_11377,N_10960);
and U13944 (N_13944,N_10878,N_11056);
nand U13945 (N_13945,N_12387,N_10797);
or U13946 (N_13946,N_9859,N_10702);
and U13947 (N_13947,N_10864,N_10611);
or U13948 (N_13948,N_11324,N_10113);
nor U13949 (N_13949,N_11548,N_12486);
and U13950 (N_13950,N_10068,N_11494);
or U13951 (N_13951,N_10453,N_11531);
nand U13952 (N_13952,N_10121,N_11869);
nand U13953 (N_13953,N_10483,N_11466);
or U13954 (N_13954,N_11672,N_10043);
or U13955 (N_13955,N_9423,N_10422);
nor U13956 (N_13956,N_11125,N_11901);
nor U13957 (N_13957,N_12256,N_11036);
or U13958 (N_13958,N_12490,N_9479);
or U13959 (N_13959,N_10765,N_10480);
and U13960 (N_13960,N_10539,N_11940);
nor U13961 (N_13961,N_11488,N_11043);
nor U13962 (N_13962,N_10099,N_12276);
or U13963 (N_13963,N_10407,N_10309);
nor U13964 (N_13964,N_12423,N_12259);
nor U13965 (N_13965,N_11707,N_10206);
nand U13966 (N_13966,N_9834,N_11268);
and U13967 (N_13967,N_11607,N_11294);
and U13968 (N_13968,N_9442,N_10567);
or U13969 (N_13969,N_9424,N_9920);
nand U13970 (N_13970,N_10355,N_10143);
xor U13971 (N_13971,N_9490,N_10366);
and U13972 (N_13972,N_9417,N_10923);
nor U13973 (N_13973,N_12417,N_11059);
and U13974 (N_13974,N_10732,N_10734);
and U13975 (N_13975,N_10978,N_10899);
nand U13976 (N_13976,N_11040,N_9990);
or U13977 (N_13977,N_11773,N_10584);
nor U13978 (N_13978,N_10061,N_11798);
or U13979 (N_13979,N_9453,N_9567);
and U13980 (N_13980,N_10167,N_11398);
and U13981 (N_13981,N_11890,N_11674);
or U13982 (N_13982,N_9877,N_12255);
xnor U13983 (N_13983,N_10519,N_9519);
and U13984 (N_13984,N_9966,N_12191);
or U13985 (N_13985,N_10398,N_10506);
nand U13986 (N_13986,N_12269,N_12487);
or U13987 (N_13987,N_10395,N_9880);
or U13988 (N_13988,N_10100,N_11372);
or U13989 (N_13989,N_11216,N_10850);
or U13990 (N_13990,N_9935,N_11098);
nand U13991 (N_13991,N_10534,N_11709);
nand U13992 (N_13992,N_11720,N_11241);
and U13993 (N_13993,N_11771,N_9769);
nor U13994 (N_13994,N_11118,N_9496);
xor U13995 (N_13995,N_11889,N_11354);
nor U13996 (N_13996,N_12339,N_10076);
or U13997 (N_13997,N_12038,N_9605);
or U13998 (N_13998,N_11439,N_11145);
and U13999 (N_13999,N_10542,N_9473);
or U14000 (N_14000,N_12404,N_10406);
nor U14001 (N_14001,N_10694,N_10726);
or U14002 (N_14002,N_10642,N_11248);
nand U14003 (N_14003,N_11320,N_11549);
or U14004 (N_14004,N_11087,N_10360);
nor U14005 (N_14005,N_12326,N_10721);
or U14006 (N_14006,N_12325,N_9889);
or U14007 (N_14007,N_9764,N_12333);
nand U14008 (N_14008,N_10300,N_12309);
and U14009 (N_14009,N_12243,N_10348);
nand U14010 (N_14010,N_11456,N_12049);
nor U14011 (N_14011,N_9768,N_12262);
and U14012 (N_14012,N_9995,N_12440);
or U14013 (N_14013,N_12351,N_10135);
and U14014 (N_14014,N_10499,N_11874);
nand U14015 (N_14015,N_12400,N_9739);
nand U14016 (N_14016,N_9946,N_10009);
or U14017 (N_14017,N_10828,N_9882);
xor U14018 (N_14018,N_11089,N_10027);
nor U14019 (N_14019,N_11174,N_10289);
or U14020 (N_14020,N_11173,N_12472);
and U14021 (N_14021,N_12271,N_12415);
or U14022 (N_14022,N_12242,N_10853);
xor U14023 (N_14023,N_11982,N_11337);
or U14024 (N_14024,N_9743,N_9526);
nand U14025 (N_14025,N_9415,N_12424);
and U14026 (N_14026,N_11472,N_10299);
or U14027 (N_14027,N_11359,N_9858);
nor U14028 (N_14028,N_9821,N_10107);
nor U14029 (N_14029,N_10217,N_10367);
nand U14030 (N_14030,N_12212,N_10817);
nand U14031 (N_14031,N_9462,N_11995);
or U14032 (N_14032,N_10881,N_12428);
nor U14033 (N_14033,N_12258,N_11994);
or U14034 (N_14034,N_10000,N_9928);
nand U14035 (N_14035,N_11987,N_11152);
xnor U14036 (N_14036,N_10376,N_9906);
or U14037 (N_14037,N_10976,N_9439);
and U14038 (N_14038,N_10705,N_11657);
or U14039 (N_14039,N_11832,N_11698);
nor U14040 (N_14040,N_9827,N_10668);
or U14041 (N_14041,N_11164,N_12374);
xnor U14042 (N_14042,N_12120,N_9798);
nand U14043 (N_14043,N_11108,N_10602);
or U14044 (N_14044,N_11906,N_10838);
or U14045 (N_14045,N_10290,N_12439);
or U14046 (N_14046,N_9774,N_10384);
nor U14047 (N_14047,N_11571,N_9860);
or U14048 (N_14048,N_10383,N_9957);
or U14049 (N_14049,N_10349,N_9939);
and U14050 (N_14050,N_11290,N_10636);
xnor U14051 (N_14051,N_9952,N_11541);
and U14052 (N_14052,N_11110,N_9517);
and U14053 (N_14053,N_10337,N_10710);
xor U14054 (N_14054,N_10644,N_11495);
nand U14055 (N_14055,N_12155,N_10268);
and U14056 (N_14056,N_10792,N_10055);
or U14057 (N_14057,N_11392,N_11114);
xor U14058 (N_14058,N_9794,N_11071);
and U14059 (N_14059,N_11565,N_10420);
or U14060 (N_14060,N_12018,N_11191);
or U14061 (N_14061,N_9684,N_11965);
and U14062 (N_14062,N_10679,N_11244);
or U14063 (N_14063,N_12094,N_9793);
and U14064 (N_14064,N_11185,N_11197);
nand U14065 (N_14065,N_9805,N_10784);
nand U14066 (N_14066,N_12377,N_10198);
nand U14067 (N_14067,N_12218,N_11103);
or U14068 (N_14068,N_10421,N_11404);
or U14069 (N_14069,N_11166,N_10532);
nor U14070 (N_14070,N_9927,N_10013);
nand U14071 (N_14071,N_12148,N_10727);
nor U14072 (N_14072,N_11240,N_9379);
and U14073 (N_14073,N_12018,N_9977);
nand U14074 (N_14074,N_12434,N_11985);
nor U14075 (N_14075,N_11998,N_10885);
or U14076 (N_14076,N_9805,N_10613);
xnor U14077 (N_14077,N_12189,N_11357);
and U14078 (N_14078,N_11576,N_12058);
and U14079 (N_14079,N_9743,N_12132);
or U14080 (N_14080,N_11430,N_12063);
nor U14081 (N_14081,N_11962,N_9399);
or U14082 (N_14082,N_9706,N_11085);
and U14083 (N_14083,N_10183,N_12160);
or U14084 (N_14084,N_12211,N_11206);
or U14085 (N_14085,N_10615,N_12235);
nand U14086 (N_14086,N_12004,N_11194);
nand U14087 (N_14087,N_10855,N_9770);
and U14088 (N_14088,N_10039,N_11524);
nor U14089 (N_14089,N_10310,N_10990);
or U14090 (N_14090,N_12410,N_10413);
or U14091 (N_14091,N_12148,N_11739);
xnor U14092 (N_14092,N_12156,N_10310);
and U14093 (N_14093,N_10972,N_9958);
nand U14094 (N_14094,N_11817,N_11684);
and U14095 (N_14095,N_11355,N_10260);
nand U14096 (N_14096,N_9836,N_10655);
nor U14097 (N_14097,N_10008,N_12027);
nor U14098 (N_14098,N_10151,N_11391);
nor U14099 (N_14099,N_11338,N_11255);
xnor U14100 (N_14100,N_10180,N_9954);
or U14101 (N_14101,N_10115,N_11558);
nor U14102 (N_14102,N_10318,N_12312);
nand U14103 (N_14103,N_10339,N_12182);
or U14104 (N_14104,N_10081,N_12472);
or U14105 (N_14105,N_10274,N_12155);
xor U14106 (N_14106,N_9863,N_10617);
or U14107 (N_14107,N_11515,N_9656);
or U14108 (N_14108,N_10517,N_10649);
or U14109 (N_14109,N_11890,N_9736);
nand U14110 (N_14110,N_11680,N_10690);
or U14111 (N_14111,N_10535,N_11131);
nor U14112 (N_14112,N_12437,N_10816);
and U14113 (N_14113,N_10702,N_11950);
xnor U14114 (N_14114,N_9818,N_9635);
nand U14115 (N_14115,N_10204,N_11545);
nor U14116 (N_14116,N_9467,N_9603);
nand U14117 (N_14117,N_10726,N_10944);
nor U14118 (N_14118,N_12129,N_9542);
nor U14119 (N_14119,N_11622,N_11457);
nand U14120 (N_14120,N_12209,N_9673);
and U14121 (N_14121,N_10170,N_11522);
and U14122 (N_14122,N_12018,N_9912);
or U14123 (N_14123,N_11467,N_12475);
or U14124 (N_14124,N_11894,N_9999);
nor U14125 (N_14125,N_12004,N_12089);
xor U14126 (N_14126,N_9814,N_10427);
nand U14127 (N_14127,N_11055,N_9919);
or U14128 (N_14128,N_11641,N_10385);
or U14129 (N_14129,N_11593,N_11529);
nand U14130 (N_14130,N_10166,N_10297);
nand U14131 (N_14131,N_10085,N_10181);
xnor U14132 (N_14132,N_9716,N_10539);
or U14133 (N_14133,N_12441,N_9918);
nor U14134 (N_14134,N_10124,N_12300);
or U14135 (N_14135,N_11296,N_12029);
xor U14136 (N_14136,N_12043,N_12396);
or U14137 (N_14137,N_11535,N_11205);
and U14138 (N_14138,N_12388,N_11706);
nor U14139 (N_14139,N_11570,N_11479);
and U14140 (N_14140,N_10509,N_11427);
nand U14141 (N_14141,N_10451,N_10166);
nor U14142 (N_14142,N_11034,N_12078);
nand U14143 (N_14143,N_11131,N_12339);
or U14144 (N_14144,N_11335,N_12420);
and U14145 (N_14145,N_9487,N_11816);
and U14146 (N_14146,N_9687,N_11408);
nand U14147 (N_14147,N_11386,N_9465);
and U14148 (N_14148,N_11297,N_10282);
and U14149 (N_14149,N_11758,N_12146);
nor U14150 (N_14150,N_10265,N_10393);
or U14151 (N_14151,N_12052,N_9967);
or U14152 (N_14152,N_9380,N_12234);
or U14153 (N_14153,N_10211,N_11869);
or U14154 (N_14154,N_9646,N_11721);
nand U14155 (N_14155,N_9609,N_11653);
nand U14156 (N_14156,N_10114,N_9447);
and U14157 (N_14157,N_11044,N_10948);
or U14158 (N_14158,N_11722,N_11049);
xnor U14159 (N_14159,N_10471,N_11497);
or U14160 (N_14160,N_11239,N_9847);
and U14161 (N_14161,N_11504,N_10937);
and U14162 (N_14162,N_12205,N_12139);
and U14163 (N_14163,N_11055,N_12324);
or U14164 (N_14164,N_10146,N_12469);
and U14165 (N_14165,N_12474,N_12493);
nor U14166 (N_14166,N_10178,N_9586);
and U14167 (N_14167,N_9652,N_11549);
or U14168 (N_14168,N_9805,N_10148);
or U14169 (N_14169,N_10180,N_11442);
or U14170 (N_14170,N_9998,N_11816);
nor U14171 (N_14171,N_11384,N_12096);
and U14172 (N_14172,N_11271,N_10500);
nand U14173 (N_14173,N_11978,N_11810);
nor U14174 (N_14174,N_11468,N_11148);
nor U14175 (N_14175,N_9486,N_10316);
xor U14176 (N_14176,N_11749,N_11534);
nor U14177 (N_14177,N_9986,N_10041);
or U14178 (N_14178,N_11078,N_9825);
nor U14179 (N_14179,N_12077,N_10930);
and U14180 (N_14180,N_10020,N_10198);
or U14181 (N_14181,N_10244,N_11220);
or U14182 (N_14182,N_9681,N_11271);
nand U14183 (N_14183,N_10743,N_10650);
nand U14184 (N_14184,N_11390,N_12424);
and U14185 (N_14185,N_11567,N_11084);
nand U14186 (N_14186,N_11200,N_9793);
or U14187 (N_14187,N_12211,N_11340);
nor U14188 (N_14188,N_10699,N_9481);
nor U14189 (N_14189,N_10525,N_12254);
and U14190 (N_14190,N_11928,N_10849);
nand U14191 (N_14191,N_10880,N_12472);
xnor U14192 (N_14192,N_12471,N_11477);
or U14193 (N_14193,N_10887,N_11440);
nand U14194 (N_14194,N_11450,N_11887);
and U14195 (N_14195,N_11037,N_11360);
or U14196 (N_14196,N_9690,N_11127);
or U14197 (N_14197,N_12024,N_11032);
nor U14198 (N_14198,N_9753,N_10915);
nand U14199 (N_14199,N_11651,N_9452);
nor U14200 (N_14200,N_9759,N_10883);
xor U14201 (N_14201,N_10673,N_9794);
nor U14202 (N_14202,N_10308,N_9966);
nor U14203 (N_14203,N_12233,N_12464);
and U14204 (N_14204,N_11184,N_11514);
or U14205 (N_14205,N_10675,N_9842);
nand U14206 (N_14206,N_10246,N_11444);
nand U14207 (N_14207,N_12175,N_9485);
nor U14208 (N_14208,N_11461,N_11654);
xnor U14209 (N_14209,N_9829,N_11504);
nand U14210 (N_14210,N_10539,N_9512);
xor U14211 (N_14211,N_11241,N_10315);
nand U14212 (N_14212,N_9520,N_9475);
nor U14213 (N_14213,N_11141,N_9804);
xnor U14214 (N_14214,N_9711,N_9780);
and U14215 (N_14215,N_11190,N_9976);
and U14216 (N_14216,N_12450,N_10360);
nand U14217 (N_14217,N_11896,N_10684);
nand U14218 (N_14218,N_9934,N_11830);
xnor U14219 (N_14219,N_11622,N_12441);
nand U14220 (N_14220,N_10637,N_11941);
xor U14221 (N_14221,N_12295,N_11290);
nor U14222 (N_14222,N_9444,N_10213);
nor U14223 (N_14223,N_11078,N_12470);
nor U14224 (N_14224,N_11184,N_10156);
nand U14225 (N_14225,N_10560,N_10033);
nor U14226 (N_14226,N_10564,N_11197);
nand U14227 (N_14227,N_10367,N_11398);
nand U14228 (N_14228,N_10220,N_10052);
and U14229 (N_14229,N_10535,N_12100);
nor U14230 (N_14230,N_10974,N_10130);
and U14231 (N_14231,N_12216,N_10321);
nor U14232 (N_14232,N_10360,N_9989);
or U14233 (N_14233,N_11823,N_11086);
nand U14234 (N_14234,N_9509,N_12469);
and U14235 (N_14235,N_9736,N_11108);
nand U14236 (N_14236,N_11447,N_9771);
and U14237 (N_14237,N_12386,N_11017);
nor U14238 (N_14238,N_11220,N_10490);
or U14239 (N_14239,N_11409,N_11797);
nand U14240 (N_14240,N_11202,N_10458);
xnor U14241 (N_14241,N_11082,N_10508);
and U14242 (N_14242,N_11282,N_12357);
nor U14243 (N_14243,N_10325,N_9752);
nand U14244 (N_14244,N_11032,N_11114);
or U14245 (N_14245,N_11519,N_10598);
nor U14246 (N_14246,N_11698,N_9521);
nand U14247 (N_14247,N_11962,N_12190);
or U14248 (N_14248,N_11000,N_10761);
nor U14249 (N_14249,N_11696,N_9842);
nand U14250 (N_14250,N_10136,N_10233);
nand U14251 (N_14251,N_9555,N_9725);
nand U14252 (N_14252,N_9714,N_11846);
or U14253 (N_14253,N_11459,N_9556);
nand U14254 (N_14254,N_10785,N_10402);
or U14255 (N_14255,N_10290,N_10326);
nor U14256 (N_14256,N_9702,N_10844);
nor U14257 (N_14257,N_9589,N_11267);
nand U14258 (N_14258,N_11982,N_9653);
nor U14259 (N_14259,N_12153,N_10125);
nand U14260 (N_14260,N_10510,N_11027);
or U14261 (N_14261,N_10679,N_9829);
nor U14262 (N_14262,N_10212,N_11783);
and U14263 (N_14263,N_11550,N_10970);
nand U14264 (N_14264,N_11225,N_11970);
or U14265 (N_14265,N_10705,N_11024);
nor U14266 (N_14266,N_12118,N_10212);
and U14267 (N_14267,N_11161,N_10986);
nand U14268 (N_14268,N_9849,N_11830);
xnor U14269 (N_14269,N_11960,N_11297);
xnor U14270 (N_14270,N_10305,N_9401);
and U14271 (N_14271,N_10735,N_12343);
and U14272 (N_14272,N_10234,N_10953);
nand U14273 (N_14273,N_9999,N_9584);
xnor U14274 (N_14274,N_11651,N_11021);
nand U14275 (N_14275,N_10188,N_11109);
nor U14276 (N_14276,N_10634,N_10853);
or U14277 (N_14277,N_9643,N_9380);
or U14278 (N_14278,N_10063,N_11409);
or U14279 (N_14279,N_10182,N_11467);
nor U14280 (N_14280,N_11057,N_9820);
or U14281 (N_14281,N_11710,N_11737);
or U14282 (N_14282,N_10348,N_9426);
nor U14283 (N_14283,N_11298,N_12083);
nor U14284 (N_14284,N_11585,N_9842);
xor U14285 (N_14285,N_12274,N_11351);
nor U14286 (N_14286,N_11779,N_10738);
or U14287 (N_14287,N_12452,N_9827);
nand U14288 (N_14288,N_11831,N_11625);
nor U14289 (N_14289,N_10456,N_12241);
nand U14290 (N_14290,N_11031,N_10424);
nor U14291 (N_14291,N_10173,N_12296);
nor U14292 (N_14292,N_11347,N_9867);
and U14293 (N_14293,N_11524,N_10536);
nand U14294 (N_14294,N_11184,N_9948);
and U14295 (N_14295,N_10599,N_9996);
nor U14296 (N_14296,N_9848,N_10315);
xor U14297 (N_14297,N_10660,N_11112);
and U14298 (N_14298,N_11284,N_12164);
or U14299 (N_14299,N_10767,N_11613);
or U14300 (N_14300,N_9936,N_9767);
and U14301 (N_14301,N_9961,N_11442);
or U14302 (N_14302,N_10199,N_10640);
xnor U14303 (N_14303,N_9734,N_11554);
nor U14304 (N_14304,N_9590,N_12036);
or U14305 (N_14305,N_10805,N_11839);
xnor U14306 (N_14306,N_10839,N_11245);
nor U14307 (N_14307,N_10163,N_11561);
nand U14308 (N_14308,N_11108,N_9901);
and U14309 (N_14309,N_12292,N_12196);
or U14310 (N_14310,N_11914,N_11871);
xnor U14311 (N_14311,N_11249,N_10339);
nand U14312 (N_14312,N_11187,N_12162);
nand U14313 (N_14313,N_9724,N_10865);
nor U14314 (N_14314,N_11458,N_11207);
nor U14315 (N_14315,N_9980,N_11777);
nor U14316 (N_14316,N_11796,N_11594);
nand U14317 (N_14317,N_11227,N_11478);
and U14318 (N_14318,N_11766,N_10370);
or U14319 (N_14319,N_9885,N_11722);
nand U14320 (N_14320,N_10336,N_9844);
nor U14321 (N_14321,N_9848,N_12160);
nor U14322 (N_14322,N_11887,N_10106);
nand U14323 (N_14323,N_10448,N_9672);
xor U14324 (N_14324,N_11383,N_10516);
nor U14325 (N_14325,N_12294,N_11421);
and U14326 (N_14326,N_11182,N_9663);
nor U14327 (N_14327,N_11314,N_10309);
nand U14328 (N_14328,N_9390,N_10717);
nor U14329 (N_14329,N_9798,N_12431);
nand U14330 (N_14330,N_11194,N_10347);
nor U14331 (N_14331,N_10802,N_11426);
nand U14332 (N_14332,N_10832,N_9960);
nor U14333 (N_14333,N_9566,N_9605);
nand U14334 (N_14334,N_12248,N_12469);
xnor U14335 (N_14335,N_9741,N_12135);
or U14336 (N_14336,N_10863,N_11345);
nand U14337 (N_14337,N_10615,N_10662);
and U14338 (N_14338,N_9615,N_11663);
nand U14339 (N_14339,N_9984,N_10472);
nor U14340 (N_14340,N_10201,N_12128);
nand U14341 (N_14341,N_9823,N_10560);
nand U14342 (N_14342,N_9603,N_10824);
and U14343 (N_14343,N_10857,N_12444);
nand U14344 (N_14344,N_9753,N_11672);
or U14345 (N_14345,N_10545,N_12280);
or U14346 (N_14346,N_10673,N_10900);
nor U14347 (N_14347,N_9397,N_12399);
and U14348 (N_14348,N_9799,N_12169);
nor U14349 (N_14349,N_9488,N_10206);
or U14350 (N_14350,N_10809,N_9845);
nor U14351 (N_14351,N_10931,N_11207);
nand U14352 (N_14352,N_11225,N_10721);
xor U14353 (N_14353,N_11892,N_11102);
or U14354 (N_14354,N_10496,N_10611);
and U14355 (N_14355,N_12498,N_10080);
and U14356 (N_14356,N_11383,N_11770);
nor U14357 (N_14357,N_10037,N_11770);
and U14358 (N_14358,N_9972,N_10029);
and U14359 (N_14359,N_10760,N_9492);
nand U14360 (N_14360,N_9963,N_11261);
and U14361 (N_14361,N_11521,N_12086);
xor U14362 (N_14362,N_12300,N_10905);
and U14363 (N_14363,N_10142,N_10649);
nor U14364 (N_14364,N_10884,N_10543);
nor U14365 (N_14365,N_10920,N_10187);
nand U14366 (N_14366,N_12202,N_11869);
or U14367 (N_14367,N_12268,N_9378);
or U14368 (N_14368,N_10479,N_11942);
and U14369 (N_14369,N_10713,N_12453);
nand U14370 (N_14370,N_12437,N_9961);
and U14371 (N_14371,N_10131,N_10862);
nor U14372 (N_14372,N_9709,N_10552);
nor U14373 (N_14373,N_9379,N_10296);
or U14374 (N_14374,N_11989,N_9964);
nand U14375 (N_14375,N_9379,N_9817);
and U14376 (N_14376,N_10996,N_11357);
and U14377 (N_14377,N_12166,N_11439);
nor U14378 (N_14378,N_11762,N_10143);
and U14379 (N_14379,N_10069,N_9904);
xor U14380 (N_14380,N_11666,N_10919);
or U14381 (N_14381,N_10123,N_11235);
nand U14382 (N_14382,N_11442,N_11794);
nor U14383 (N_14383,N_12425,N_11596);
nor U14384 (N_14384,N_12020,N_12485);
nand U14385 (N_14385,N_10953,N_10983);
or U14386 (N_14386,N_12178,N_9582);
or U14387 (N_14387,N_11283,N_10311);
or U14388 (N_14388,N_10053,N_10455);
xnor U14389 (N_14389,N_11989,N_11828);
nand U14390 (N_14390,N_10788,N_12435);
and U14391 (N_14391,N_11000,N_10099);
and U14392 (N_14392,N_12175,N_10926);
and U14393 (N_14393,N_11773,N_9828);
or U14394 (N_14394,N_9558,N_11955);
and U14395 (N_14395,N_12250,N_10959);
and U14396 (N_14396,N_10115,N_11856);
xor U14397 (N_14397,N_11251,N_9929);
nand U14398 (N_14398,N_12295,N_9716);
and U14399 (N_14399,N_9448,N_11893);
nor U14400 (N_14400,N_9575,N_9631);
and U14401 (N_14401,N_10750,N_9816);
nor U14402 (N_14402,N_11009,N_10513);
nor U14403 (N_14403,N_10047,N_12485);
or U14404 (N_14404,N_10328,N_9847);
xor U14405 (N_14405,N_12210,N_10201);
nand U14406 (N_14406,N_11782,N_12470);
and U14407 (N_14407,N_9706,N_11303);
nand U14408 (N_14408,N_11074,N_10055);
nor U14409 (N_14409,N_12183,N_10377);
nor U14410 (N_14410,N_10495,N_10722);
xor U14411 (N_14411,N_10076,N_9483);
and U14412 (N_14412,N_9647,N_11422);
or U14413 (N_14413,N_10898,N_11624);
xor U14414 (N_14414,N_9537,N_10838);
and U14415 (N_14415,N_11389,N_10029);
nand U14416 (N_14416,N_11679,N_12047);
or U14417 (N_14417,N_9706,N_12401);
nand U14418 (N_14418,N_9627,N_12226);
nor U14419 (N_14419,N_9861,N_11630);
nor U14420 (N_14420,N_11724,N_10660);
nand U14421 (N_14421,N_11165,N_11292);
or U14422 (N_14422,N_9471,N_10597);
or U14423 (N_14423,N_12109,N_11462);
or U14424 (N_14424,N_9819,N_10769);
or U14425 (N_14425,N_9466,N_11934);
xor U14426 (N_14426,N_9444,N_12250);
nand U14427 (N_14427,N_10124,N_12463);
nand U14428 (N_14428,N_11157,N_11366);
and U14429 (N_14429,N_11835,N_12433);
or U14430 (N_14430,N_10057,N_11281);
nor U14431 (N_14431,N_10956,N_11719);
and U14432 (N_14432,N_11217,N_9406);
nand U14433 (N_14433,N_10775,N_11382);
or U14434 (N_14434,N_11504,N_10972);
nor U14435 (N_14435,N_11490,N_10025);
or U14436 (N_14436,N_10723,N_12155);
nor U14437 (N_14437,N_10749,N_11055);
nor U14438 (N_14438,N_10197,N_11308);
xor U14439 (N_14439,N_10328,N_12222);
nand U14440 (N_14440,N_12488,N_11951);
nand U14441 (N_14441,N_10664,N_10048);
or U14442 (N_14442,N_11659,N_10808);
and U14443 (N_14443,N_12274,N_9973);
and U14444 (N_14444,N_11435,N_9496);
or U14445 (N_14445,N_11559,N_10737);
or U14446 (N_14446,N_10230,N_11258);
nor U14447 (N_14447,N_10124,N_11832);
or U14448 (N_14448,N_12145,N_10216);
xnor U14449 (N_14449,N_10573,N_10019);
xnor U14450 (N_14450,N_11155,N_11418);
and U14451 (N_14451,N_11054,N_10328);
and U14452 (N_14452,N_10177,N_10217);
xnor U14453 (N_14453,N_12135,N_10058);
xor U14454 (N_14454,N_12494,N_10668);
nand U14455 (N_14455,N_11009,N_11739);
xnor U14456 (N_14456,N_10982,N_10780);
nor U14457 (N_14457,N_9660,N_9976);
and U14458 (N_14458,N_9616,N_12090);
or U14459 (N_14459,N_10684,N_10754);
nor U14460 (N_14460,N_10456,N_10976);
nand U14461 (N_14461,N_9813,N_10983);
or U14462 (N_14462,N_11904,N_9697);
and U14463 (N_14463,N_11685,N_11966);
and U14464 (N_14464,N_12094,N_10436);
or U14465 (N_14465,N_11409,N_10280);
nor U14466 (N_14466,N_11431,N_9936);
or U14467 (N_14467,N_11381,N_12257);
nand U14468 (N_14468,N_9739,N_11437);
nand U14469 (N_14469,N_12111,N_10749);
or U14470 (N_14470,N_11650,N_9551);
or U14471 (N_14471,N_11622,N_11300);
nand U14472 (N_14472,N_11804,N_12427);
or U14473 (N_14473,N_11114,N_11854);
xor U14474 (N_14474,N_12079,N_9811);
nor U14475 (N_14475,N_10730,N_11340);
or U14476 (N_14476,N_9956,N_10135);
xnor U14477 (N_14477,N_12106,N_9858);
xnor U14478 (N_14478,N_9386,N_11737);
nor U14479 (N_14479,N_11449,N_11565);
or U14480 (N_14480,N_10288,N_10745);
or U14481 (N_14481,N_10953,N_11285);
and U14482 (N_14482,N_11073,N_11625);
nand U14483 (N_14483,N_12489,N_10698);
and U14484 (N_14484,N_9640,N_10252);
or U14485 (N_14485,N_11156,N_12390);
nor U14486 (N_14486,N_11415,N_11170);
or U14487 (N_14487,N_11971,N_11675);
nor U14488 (N_14488,N_10739,N_9504);
nor U14489 (N_14489,N_11377,N_11783);
nor U14490 (N_14490,N_11726,N_12224);
or U14491 (N_14491,N_11821,N_11314);
nor U14492 (N_14492,N_9474,N_11276);
nor U14493 (N_14493,N_10904,N_12437);
nor U14494 (N_14494,N_12271,N_11515);
and U14495 (N_14495,N_10680,N_10189);
nor U14496 (N_14496,N_11274,N_10125);
xnor U14497 (N_14497,N_11419,N_10398);
or U14498 (N_14498,N_9861,N_11263);
nand U14499 (N_14499,N_11798,N_9932);
or U14500 (N_14500,N_11889,N_12146);
and U14501 (N_14501,N_11258,N_11528);
and U14502 (N_14502,N_11678,N_12320);
nand U14503 (N_14503,N_10191,N_11215);
nor U14504 (N_14504,N_9432,N_11996);
and U14505 (N_14505,N_10565,N_10006);
or U14506 (N_14506,N_11321,N_12453);
nor U14507 (N_14507,N_10816,N_10590);
and U14508 (N_14508,N_10523,N_12299);
xnor U14509 (N_14509,N_11103,N_11479);
and U14510 (N_14510,N_10571,N_12130);
or U14511 (N_14511,N_9615,N_12214);
xor U14512 (N_14512,N_11227,N_10296);
nand U14513 (N_14513,N_12298,N_10323);
or U14514 (N_14514,N_10429,N_12144);
or U14515 (N_14515,N_11382,N_11130);
and U14516 (N_14516,N_10342,N_10393);
and U14517 (N_14517,N_12107,N_10661);
or U14518 (N_14518,N_10934,N_12427);
xor U14519 (N_14519,N_11132,N_9684);
or U14520 (N_14520,N_10500,N_10679);
nand U14521 (N_14521,N_12471,N_12437);
nor U14522 (N_14522,N_10130,N_9728);
or U14523 (N_14523,N_10604,N_9416);
xnor U14524 (N_14524,N_11119,N_11662);
nor U14525 (N_14525,N_11520,N_10501);
or U14526 (N_14526,N_10444,N_11425);
and U14527 (N_14527,N_10971,N_11769);
or U14528 (N_14528,N_10559,N_11104);
nand U14529 (N_14529,N_10273,N_11556);
and U14530 (N_14530,N_10991,N_11895);
or U14531 (N_14531,N_12222,N_10762);
and U14532 (N_14532,N_10980,N_10179);
nand U14533 (N_14533,N_10795,N_9461);
nor U14534 (N_14534,N_11557,N_11870);
and U14535 (N_14535,N_9883,N_10937);
and U14536 (N_14536,N_11404,N_9463);
or U14537 (N_14537,N_9660,N_10021);
or U14538 (N_14538,N_10842,N_12368);
and U14539 (N_14539,N_12242,N_9670);
and U14540 (N_14540,N_12484,N_9848);
and U14541 (N_14541,N_11035,N_10035);
nand U14542 (N_14542,N_11898,N_10213);
nand U14543 (N_14543,N_10309,N_12428);
and U14544 (N_14544,N_12061,N_12064);
nand U14545 (N_14545,N_11800,N_10812);
or U14546 (N_14546,N_12309,N_11521);
nor U14547 (N_14547,N_12208,N_11815);
nand U14548 (N_14548,N_10126,N_9976);
nand U14549 (N_14549,N_12418,N_12468);
and U14550 (N_14550,N_11099,N_10254);
and U14551 (N_14551,N_11028,N_12448);
nor U14552 (N_14552,N_9649,N_10516);
and U14553 (N_14553,N_9537,N_10885);
nor U14554 (N_14554,N_11482,N_9505);
nand U14555 (N_14555,N_10245,N_11348);
or U14556 (N_14556,N_10967,N_11951);
or U14557 (N_14557,N_11295,N_11607);
nand U14558 (N_14558,N_11943,N_10212);
and U14559 (N_14559,N_9902,N_9786);
and U14560 (N_14560,N_10121,N_11254);
nand U14561 (N_14561,N_9658,N_10620);
nor U14562 (N_14562,N_10084,N_11005);
nor U14563 (N_14563,N_12295,N_10995);
or U14564 (N_14564,N_11723,N_11538);
nor U14565 (N_14565,N_12247,N_9556);
nand U14566 (N_14566,N_11484,N_9531);
and U14567 (N_14567,N_11262,N_11666);
and U14568 (N_14568,N_10270,N_11194);
xor U14569 (N_14569,N_11006,N_11766);
or U14570 (N_14570,N_10811,N_10391);
nor U14571 (N_14571,N_10050,N_10004);
nand U14572 (N_14572,N_10526,N_10072);
nor U14573 (N_14573,N_10236,N_11744);
and U14574 (N_14574,N_10168,N_11576);
and U14575 (N_14575,N_10061,N_10430);
or U14576 (N_14576,N_10480,N_12489);
nor U14577 (N_14577,N_9936,N_9828);
and U14578 (N_14578,N_9407,N_11770);
and U14579 (N_14579,N_10294,N_12339);
and U14580 (N_14580,N_12189,N_11973);
or U14581 (N_14581,N_9663,N_12312);
nor U14582 (N_14582,N_11525,N_10365);
or U14583 (N_14583,N_11912,N_10555);
nand U14584 (N_14584,N_12182,N_9576);
nor U14585 (N_14585,N_12006,N_10492);
nand U14586 (N_14586,N_10477,N_12202);
nand U14587 (N_14587,N_10862,N_9774);
nor U14588 (N_14588,N_10655,N_11138);
nand U14589 (N_14589,N_11589,N_10040);
and U14590 (N_14590,N_10651,N_9889);
xor U14591 (N_14591,N_10991,N_10731);
and U14592 (N_14592,N_12194,N_9584);
or U14593 (N_14593,N_10710,N_10449);
and U14594 (N_14594,N_11095,N_10157);
and U14595 (N_14595,N_10061,N_9421);
nand U14596 (N_14596,N_12114,N_11368);
nor U14597 (N_14597,N_11740,N_10543);
nand U14598 (N_14598,N_12229,N_10439);
and U14599 (N_14599,N_12369,N_9472);
or U14600 (N_14600,N_11259,N_11648);
nor U14601 (N_14601,N_9873,N_10739);
and U14602 (N_14602,N_11730,N_10361);
and U14603 (N_14603,N_9559,N_11395);
nand U14604 (N_14604,N_9911,N_12373);
or U14605 (N_14605,N_10797,N_9507);
xnor U14606 (N_14606,N_10944,N_10563);
nand U14607 (N_14607,N_9872,N_11940);
or U14608 (N_14608,N_10640,N_12100);
nand U14609 (N_14609,N_11573,N_9762);
nor U14610 (N_14610,N_10635,N_12371);
and U14611 (N_14611,N_10342,N_9423);
nand U14612 (N_14612,N_9523,N_11302);
and U14613 (N_14613,N_9523,N_9521);
xor U14614 (N_14614,N_10781,N_11444);
nor U14615 (N_14615,N_11710,N_11909);
or U14616 (N_14616,N_12418,N_12394);
nor U14617 (N_14617,N_9985,N_9545);
nor U14618 (N_14618,N_9770,N_11538);
nor U14619 (N_14619,N_12047,N_11858);
or U14620 (N_14620,N_11586,N_10465);
nand U14621 (N_14621,N_10553,N_9923);
nor U14622 (N_14622,N_11792,N_11294);
or U14623 (N_14623,N_11659,N_10848);
nor U14624 (N_14624,N_9934,N_10940);
or U14625 (N_14625,N_9777,N_11040);
or U14626 (N_14626,N_10465,N_11045);
nor U14627 (N_14627,N_12022,N_11920);
nand U14628 (N_14628,N_12166,N_11755);
nand U14629 (N_14629,N_10250,N_11349);
nor U14630 (N_14630,N_12432,N_9737);
nor U14631 (N_14631,N_10431,N_10446);
nand U14632 (N_14632,N_10846,N_11275);
and U14633 (N_14633,N_10672,N_10800);
nor U14634 (N_14634,N_11668,N_10215);
nand U14635 (N_14635,N_12240,N_11260);
or U14636 (N_14636,N_11996,N_11635);
or U14637 (N_14637,N_11093,N_10421);
nand U14638 (N_14638,N_10056,N_10816);
xor U14639 (N_14639,N_11918,N_12094);
and U14640 (N_14640,N_12007,N_9600);
nand U14641 (N_14641,N_12154,N_9729);
and U14642 (N_14642,N_9977,N_10904);
or U14643 (N_14643,N_12266,N_11413);
or U14644 (N_14644,N_9544,N_11256);
or U14645 (N_14645,N_10147,N_11824);
nand U14646 (N_14646,N_9877,N_11452);
nor U14647 (N_14647,N_10608,N_10091);
nand U14648 (N_14648,N_10065,N_11324);
xor U14649 (N_14649,N_9920,N_12176);
xnor U14650 (N_14650,N_12141,N_11073);
and U14651 (N_14651,N_9938,N_10557);
nor U14652 (N_14652,N_11590,N_10811);
nand U14653 (N_14653,N_12287,N_9579);
nand U14654 (N_14654,N_11171,N_9803);
nand U14655 (N_14655,N_11545,N_11017);
and U14656 (N_14656,N_11975,N_10554);
xnor U14657 (N_14657,N_10368,N_11181);
nand U14658 (N_14658,N_10681,N_11095);
xor U14659 (N_14659,N_10032,N_11561);
nor U14660 (N_14660,N_11333,N_10831);
or U14661 (N_14661,N_10313,N_10688);
or U14662 (N_14662,N_9732,N_9852);
or U14663 (N_14663,N_10090,N_11007);
xor U14664 (N_14664,N_11301,N_9768);
and U14665 (N_14665,N_10191,N_10534);
nand U14666 (N_14666,N_10680,N_11184);
and U14667 (N_14667,N_11966,N_10187);
and U14668 (N_14668,N_10035,N_11658);
nor U14669 (N_14669,N_10890,N_11976);
nor U14670 (N_14670,N_12461,N_10211);
nor U14671 (N_14671,N_9740,N_11565);
and U14672 (N_14672,N_12294,N_10347);
nor U14673 (N_14673,N_10919,N_11597);
xor U14674 (N_14674,N_10311,N_10771);
nor U14675 (N_14675,N_10629,N_12497);
nor U14676 (N_14676,N_11723,N_11676);
and U14677 (N_14677,N_11960,N_10236);
and U14678 (N_14678,N_9525,N_10131);
and U14679 (N_14679,N_10249,N_9903);
nor U14680 (N_14680,N_11480,N_11353);
nor U14681 (N_14681,N_10079,N_12048);
xor U14682 (N_14682,N_11238,N_10206);
nand U14683 (N_14683,N_10218,N_11401);
or U14684 (N_14684,N_11124,N_10414);
nand U14685 (N_14685,N_10800,N_10365);
or U14686 (N_14686,N_10888,N_10916);
or U14687 (N_14687,N_11573,N_11995);
nor U14688 (N_14688,N_10216,N_10879);
nor U14689 (N_14689,N_11220,N_10973);
or U14690 (N_14690,N_11509,N_12154);
nand U14691 (N_14691,N_10453,N_10074);
xnor U14692 (N_14692,N_10919,N_11426);
and U14693 (N_14693,N_11733,N_11899);
or U14694 (N_14694,N_11806,N_11060);
nor U14695 (N_14695,N_9970,N_9548);
nor U14696 (N_14696,N_11171,N_10149);
or U14697 (N_14697,N_10163,N_9650);
xor U14698 (N_14698,N_11435,N_10201);
nand U14699 (N_14699,N_11811,N_10802);
nor U14700 (N_14700,N_11010,N_12495);
nor U14701 (N_14701,N_11244,N_11742);
and U14702 (N_14702,N_10610,N_11710);
and U14703 (N_14703,N_9795,N_9998);
or U14704 (N_14704,N_10044,N_11277);
or U14705 (N_14705,N_9964,N_12111);
nand U14706 (N_14706,N_10842,N_9434);
nand U14707 (N_14707,N_10959,N_11126);
or U14708 (N_14708,N_11966,N_11387);
or U14709 (N_14709,N_11522,N_12282);
and U14710 (N_14710,N_10483,N_10220);
or U14711 (N_14711,N_10780,N_10108);
and U14712 (N_14712,N_9899,N_12315);
or U14713 (N_14713,N_11978,N_11585);
or U14714 (N_14714,N_11014,N_11296);
nor U14715 (N_14715,N_10762,N_11181);
or U14716 (N_14716,N_10773,N_9409);
and U14717 (N_14717,N_9929,N_9681);
or U14718 (N_14718,N_10962,N_11070);
nor U14719 (N_14719,N_10960,N_10774);
nor U14720 (N_14720,N_10617,N_10853);
nor U14721 (N_14721,N_9461,N_12092);
or U14722 (N_14722,N_9448,N_9972);
or U14723 (N_14723,N_11749,N_11247);
nor U14724 (N_14724,N_9989,N_10182);
or U14725 (N_14725,N_10655,N_11498);
nor U14726 (N_14726,N_9439,N_10751);
or U14727 (N_14727,N_9762,N_10851);
nor U14728 (N_14728,N_12011,N_10693);
and U14729 (N_14729,N_9968,N_12000);
nand U14730 (N_14730,N_9747,N_10494);
nor U14731 (N_14731,N_10958,N_9951);
or U14732 (N_14732,N_10125,N_10768);
or U14733 (N_14733,N_11915,N_9737);
nor U14734 (N_14734,N_10130,N_12358);
or U14735 (N_14735,N_9444,N_10552);
nor U14736 (N_14736,N_10404,N_11899);
nand U14737 (N_14737,N_11749,N_11489);
nor U14738 (N_14738,N_11153,N_12048);
nor U14739 (N_14739,N_11697,N_12146);
nor U14740 (N_14740,N_9927,N_9468);
or U14741 (N_14741,N_10730,N_11045);
nor U14742 (N_14742,N_9880,N_12097);
and U14743 (N_14743,N_9499,N_11357);
and U14744 (N_14744,N_10180,N_12329);
and U14745 (N_14745,N_11456,N_11843);
xor U14746 (N_14746,N_10880,N_12279);
nor U14747 (N_14747,N_11723,N_9802);
and U14748 (N_14748,N_12449,N_9785);
xnor U14749 (N_14749,N_10165,N_11644);
and U14750 (N_14750,N_9539,N_9571);
or U14751 (N_14751,N_9468,N_11299);
nand U14752 (N_14752,N_10385,N_10553);
nand U14753 (N_14753,N_11633,N_12338);
nor U14754 (N_14754,N_10327,N_11265);
and U14755 (N_14755,N_9768,N_10181);
nand U14756 (N_14756,N_11125,N_10306);
or U14757 (N_14757,N_11616,N_12080);
nor U14758 (N_14758,N_9749,N_11448);
nand U14759 (N_14759,N_12400,N_9949);
and U14760 (N_14760,N_9551,N_9667);
or U14761 (N_14761,N_10373,N_12187);
or U14762 (N_14762,N_9489,N_9812);
nand U14763 (N_14763,N_12308,N_9630);
nand U14764 (N_14764,N_11355,N_11235);
nor U14765 (N_14765,N_10764,N_12303);
nor U14766 (N_14766,N_11912,N_10540);
and U14767 (N_14767,N_10530,N_11803);
nor U14768 (N_14768,N_9601,N_9807);
and U14769 (N_14769,N_10057,N_12192);
nand U14770 (N_14770,N_10928,N_9653);
nor U14771 (N_14771,N_10966,N_10807);
or U14772 (N_14772,N_10005,N_10417);
or U14773 (N_14773,N_11663,N_11318);
and U14774 (N_14774,N_12132,N_10708);
nor U14775 (N_14775,N_11482,N_12128);
nor U14776 (N_14776,N_12082,N_10508);
and U14777 (N_14777,N_12012,N_11535);
xor U14778 (N_14778,N_10550,N_9464);
and U14779 (N_14779,N_12449,N_10043);
nor U14780 (N_14780,N_10473,N_11464);
and U14781 (N_14781,N_11177,N_11675);
or U14782 (N_14782,N_9414,N_9776);
xor U14783 (N_14783,N_12316,N_11476);
nand U14784 (N_14784,N_11293,N_11027);
nor U14785 (N_14785,N_10067,N_9855);
nor U14786 (N_14786,N_11428,N_12267);
and U14787 (N_14787,N_9669,N_9542);
nor U14788 (N_14788,N_12084,N_12047);
nand U14789 (N_14789,N_11448,N_12272);
or U14790 (N_14790,N_11067,N_12081);
or U14791 (N_14791,N_10130,N_9818);
and U14792 (N_14792,N_10044,N_11469);
nand U14793 (N_14793,N_10558,N_9979);
or U14794 (N_14794,N_10238,N_11821);
nor U14795 (N_14795,N_10892,N_12416);
and U14796 (N_14796,N_10159,N_11942);
or U14797 (N_14797,N_12099,N_10159);
xor U14798 (N_14798,N_10920,N_11436);
nand U14799 (N_14799,N_12061,N_11090);
nor U14800 (N_14800,N_12201,N_11614);
nand U14801 (N_14801,N_10075,N_12435);
and U14802 (N_14802,N_9869,N_10782);
xor U14803 (N_14803,N_10293,N_12059);
nor U14804 (N_14804,N_12150,N_11314);
xor U14805 (N_14805,N_12034,N_9462);
nand U14806 (N_14806,N_11022,N_10498);
and U14807 (N_14807,N_9985,N_12225);
nand U14808 (N_14808,N_10839,N_11849);
nor U14809 (N_14809,N_12222,N_9767);
or U14810 (N_14810,N_11830,N_11174);
xor U14811 (N_14811,N_11452,N_10360);
and U14812 (N_14812,N_11729,N_10870);
xnor U14813 (N_14813,N_11299,N_10344);
nand U14814 (N_14814,N_12248,N_12028);
nand U14815 (N_14815,N_10920,N_11056);
nand U14816 (N_14816,N_10617,N_9845);
or U14817 (N_14817,N_10017,N_9571);
nor U14818 (N_14818,N_11747,N_12380);
and U14819 (N_14819,N_9433,N_10359);
nand U14820 (N_14820,N_9635,N_12207);
xnor U14821 (N_14821,N_9503,N_11739);
and U14822 (N_14822,N_9926,N_10175);
nand U14823 (N_14823,N_11648,N_10488);
and U14824 (N_14824,N_11539,N_11418);
and U14825 (N_14825,N_9594,N_10644);
xnor U14826 (N_14826,N_9820,N_11295);
nand U14827 (N_14827,N_10852,N_9834);
nand U14828 (N_14828,N_9691,N_10660);
nor U14829 (N_14829,N_12489,N_9666);
or U14830 (N_14830,N_9387,N_11761);
nand U14831 (N_14831,N_10359,N_10032);
nand U14832 (N_14832,N_11879,N_10654);
nand U14833 (N_14833,N_9683,N_10197);
and U14834 (N_14834,N_9622,N_10713);
nand U14835 (N_14835,N_10500,N_10656);
nor U14836 (N_14836,N_11910,N_11950);
and U14837 (N_14837,N_9914,N_9530);
xnor U14838 (N_14838,N_11176,N_9949);
or U14839 (N_14839,N_11219,N_11270);
nor U14840 (N_14840,N_9612,N_10687);
xnor U14841 (N_14841,N_11136,N_12227);
or U14842 (N_14842,N_12066,N_11294);
nor U14843 (N_14843,N_11361,N_11420);
nor U14844 (N_14844,N_10997,N_10759);
nand U14845 (N_14845,N_9432,N_9750);
or U14846 (N_14846,N_9943,N_11227);
or U14847 (N_14847,N_11949,N_9554);
and U14848 (N_14848,N_11227,N_10518);
nor U14849 (N_14849,N_10689,N_9994);
nand U14850 (N_14850,N_11342,N_9892);
or U14851 (N_14851,N_11445,N_11131);
or U14852 (N_14852,N_10896,N_9835);
nand U14853 (N_14853,N_10190,N_11635);
xnor U14854 (N_14854,N_12151,N_12304);
nand U14855 (N_14855,N_9771,N_9934);
or U14856 (N_14856,N_11767,N_11811);
and U14857 (N_14857,N_9964,N_10675);
xnor U14858 (N_14858,N_9512,N_11115);
or U14859 (N_14859,N_12075,N_10060);
nand U14860 (N_14860,N_10821,N_10260);
nand U14861 (N_14861,N_10415,N_9973);
and U14862 (N_14862,N_9416,N_12144);
or U14863 (N_14863,N_11008,N_12095);
nor U14864 (N_14864,N_12008,N_11143);
or U14865 (N_14865,N_11742,N_11179);
nor U14866 (N_14866,N_10908,N_10854);
or U14867 (N_14867,N_11096,N_9794);
or U14868 (N_14868,N_10422,N_10982);
or U14869 (N_14869,N_12210,N_10113);
and U14870 (N_14870,N_10365,N_12410);
or U14871 (N_14871,N_12023,N_11162);
and U14872 (N_14872,N_11503,N_10206);
and U14873 (N_14873,N_10447,N_9581);
nand U14874 (N_14874,N_9615,N_11552);
and U14875 (N_14875,N_10299,N_10616);
nor U14876 (N_14876,N_12443,N_11436);
nand U14877 (N_14877,N_12444,N_11752);
and U14878 (N_14878,N_11183,N_10722);
and U14879 (N_14879,N_10911,N_12271);
xnor U14880 (N_14880,N_10723,N_9664);
or U14881 (N_14881,N_12272,N_11406);
xor U14882 (N_14882,N_9543,N_11996);
nand U14883 (N_14883,N_10461,N_10004);
and U14884 (N_14884,N_9376,N_12009);
nor U14885 (N_14885,N_11685,N_12050);
nor U14886 (N_14886,N_12406,N_9769);
and U14887 (N_14887,N_12478,N_11997);
nand U14888 (N_14888,N_10471,N_12060);
nand U14889 (N_14889,N_10279,N_9513);
nor U14890 (N_14890,N_10220,N_11449);
or U14891 (N_14891,N_12418,N_11621);
or U14892 (N_14892,N_11475,N_12129);
nand U14893 (N_14893,N_9643,N_11586);
or U14894 (N_14894,N_9493,N_9735);
nor U14895 (N_14895,N_9963,N_9867);
nand U14896 (N_14896,N_11928,N_12249);
and U14897 (N_14897,N_10602,N_11641);
and U14898 (N_14898,N_9429,N_11878);
and U14899 (N_14899,N_12007,N_12080);
or U14900 (N_14900,N_10227,N_10357);
xnor U14901 (N_14901,N_10387,N_9865);
and U14902 (N_14902,N_12352,N_10145);
nand U14903 (N_14903,N_11559,N_9694);
xnor U14904 (N_14904,N_12124,N_10438);
or U14905 (N_14905,N_11228,N_11199);
xor U14906 (N_14906,N_11960,N_11966);
or U14907 (N_14907,N_10125,N_10815);
or U14908 (N_14908,N_10751,N_10392);
nand U14909 (N_14909,N_12041,N_11881);
nand U14910 (N_14910,N_12040,N_11785);
or U14911 (N_14911,N_11243,N_9921);
nor U14912 (N_14912,N_11121,N_10316);
or U14913 (N_14913,N_12193,N_10394);
nor U14914 (N_14914,N_10377,N_10120);
nor U14915 (N_14915,N_10360,N_11008);
or U14916 (N_14916,N_11921,N_10938);
nand U14917 (N_14917,N_12013,N_11087);
or U14918 (N_14918,N_11758,N_12022);
or U14919 (N_14919,N_9437,N_12435);
or U14920 (N_14920,N_10594,N_9781);
or U14921 (N_14921,N_10637,N_10043);
nand U14922 (N_14922,N_11001,N_9796);
or U14923 (N_14923,N_9745,N_11635);
nor U14924 (N_14924,N_10584,N_11342);
nor U14925 (N_14925,N_11591,N_9394);
and U14926 (N_14926,N_10757,N_10995);
and U14927 (N_14927,N_9429,N_12496);
nor U14928 (N_14928,N_10444,N_11086);
or U14929 (N_14929,N_10235,N_12075);
nor U14930 (N_14930,N_10513,N_10357);
nand U14931 (N_14931,N_10312,N_10246);
xnor U14932 (N_14932,N_9824,N_10127);
nand U14933 (N_14933,N_11422,N_11425);
xnor U14934 (N_14934,N_12310,N_11524);
and U14935 (N_14935,N_10836,N_11201);
or U14936 (N_14936,N_10586,N_10508);
and U14937 (N_14937,N_11103,N_11020);
nor U14938 (N_14938,N_11794,N_12470);
nand U14939 (N_14939,N_11693,N_11957);
nor U14940 (N_14940,N_10283,N_11246);
xor U14941 (N_14941,N_11460,N_12005);
nor U14942 (N_14942,N_12282,N_12164);
nand U14943 (N_14943,N_12391,N_10486);
or U14944 (N_14944,N_12409,N_10501);
nand U14945 (N_14945,N_9922,N_9708);
nor U14946 (N_14946,N_12039,N_10714);
and U14947 (N_14947,N_9712,N_9784);
nand U14948 (N_14948,N_10099,N_11025);
or U14949 (N_14949,N_12226,N_10537);
xnor U14950 (N_14950,N_10788,N_12400);
nand U14951 (N_14951,N_9637,N_10675);
nor U14952 (N_14952,N_11664,N_11840);
and U14953 (N_14953,N_10644,N_10196);
xor U14954 (N_14954,N_10773,N_10909);
nand U14955 (N_14955,N_11110,N_12206);
and U14956 (N_14956,N_12255,N_10750);
or U14957 (N_14957,N_9984,N_12202);
or U14958 (N_14958,N_11670,N_9533);
nand U14959 (N_14959,N_10243,N_12248);
and U14960 (N_14960,N_9923,N_11101);
nand U14961 (N_14961,N_9452,N_10058);
and U14962 (N_14962,N_9464,N_11945);
or U14963 (N_14963,N_10834,N_11030);
nand U14964 (N_14964,N_10031,N_11873);
nor U14965 (N_14965,N_11181,N_10627);
or U14966 (N_14966,N_12428,N_9421);
and U14967 (N_14967,N_9785,N_11018);
nor U14968 (N_14968,N_12098,N_11908);
nor U14969 (N_14969,N_9603,N_11088);
or U14970 (N_14970,N_10204,N_12081);
nand U14971 (N_14971,N_12291,N_10391);
nor U14972 (N_14972,N_11743,N_11132);
and U14973 (N_14973,N_9719,N_9947);
nand U14974 (N_14974,N_12140,N_9957);
nand U14975 (N_14975,N_10596,N_11858);
and U14976 (N_14976,N_10912,N_12014);
or U14977 (N_14977,N_10594,N_11293);
nor U14978 (N_14978,N_11920,N_11257);
nand U14979 (N_14979,N_9471,N_11533);
and U14980 (N_14980,N_10352,N_10784);
xor U14981 (N_14981,N_9633,N_11564);
and U14982 (N_14982,N_11752,N_11594);
or U14983 (N_14983,N_11082,N_11677);
and U14984 (N_14984,N_10240,N_9682);
and U14985 (N_14985,N_11567,N_11861);
nor U14986 (N_14986,N_10628,N_11060);
or U14987 (N_14987,N_11103,N_12108);
nand U14988 (N_14988,N_10008,N_11024);
nand U14989 (N_14989,N_10597,N_9487);
nor U14990 (N_14990,N_11595,N_9716);
nand U14991 (N_14991,N_9665,N_10781);
and U14992 (N_14992,N_11964,N_11082);
and U14993 (N_14993,N_10023,N_11454);
nand U14994 (N_14994,N_9463,N_9870);
and U14995 (N_14995,N_10397,N_10602);
nor U14996 (N_14996,N_11376,N_10791);
and U14997 (N_14997,N_12155,N_10872);
nor U14998 (N_14998,N_11420,N_10929);
or U14999 (N_14999,N_9729,N_11523);
nor U15000 (N_15000,N_9924,N_10057);
nand U15001 (N_15001,N_10802,N_11372);
xnor U15002 (N_15002,N_11180,N_11123);
and U15003 (N_15003,N_9683,N_11009);
nor U15004 (N_15004,N_12383,N_10621);
xnor U15005 (N_15005,N_9815,N_10162);
nand U15006 (N_15006,N_11398,N_11317);
nand U15007 (N_15007,N_12426,N_11781);
nand U15008 (N_15008,N_10228,N_10143);
nand U15009 (N_15009,N_11637,N_12206);
nand U15010 (N_15010,N_11269,N_12251);
nor U15011 (N_15011,N_10073,N_11739);
and U15012 (N_15012,N_9640,N_11439);
nand U15013 (N_15013,N_9907,N_10222);
and U15014 (N_15014,N_12129,N_9430);
or U15015 (N_15015,N_11369,N_9512);
and U15016 (N_15016,N_10107,N_10328);
nor U15017 (N_15017,N_9622,N_9856);
and U15018 (N_15018,N_12383,N_11530);
nand U15019 (N_15019,N_12465,N_11170);
or U15020 (N_15020,N_11602,N_11022);
or U15021 (N_15021,N_11246,N_11180);
or U15022 (N_15022,N_11205,N_10199);
nor U15023 (N_15023,N_12230,N_10392);
xnor U15024 (N_15024,N_10814,N_10860);
or U15025 (N_15025,N_11333,N_11477);
nand U15026 (N_15026,N_12110,N_10322);
nand U15027 (N_15027,N_11590,N_9420);
nor U15028 (N_15028,N_11974,N_11740);
or U15029 (N_15029,N_10504,N_9692);
and U15030 (N_15030,N_10481,N_11380);
xor U15031 (N_15031,N_9934,N_10742);
and U15032 (N_15032,N_10331,N_11740);
or U15033 (N_15033,N_12123,N_10188);
nor U15034 (N_15034,N_10174,N_10605);
nor U15035 (N_15035,N_10862,N_10151);
nand U15036 (N_15036,N_9851,N_11028);
nor U15037 (N_15037,N_9444,N_12489);
or U15038 (N_15038,N_10826,N_11013);
nand U15039 (N_15039,N_10824,N_11740);
nor U15040 (N_15040,N_9454,N_12447);
or U15041 (N_15041,N_9519,N_9816);
xor U15042 (N_15042,N_10204,N_12386);
xor U15043 (N_15043,N_10691,N_10947);
nor U15044 (N_15044,N_11945,N_10914);
or U15045 (N_15045,N_11507,N_10143);
nor U15046 (N_15046,N_10994,N_10752);
nand U15047 (N_15047,N_12055,N_11934);
or U15048 (N_15048,N_9764,N_12218);
and U15049 (N_15049,N_12488,N_11906);
and U15050 (N_15050,N_10645,N_9720);
nand U15051 (N_15051,N_11035,N_11081);
xnor U15052 (N_15052,N_12327,N_10983);
or U15053 (N_15053,N_11613,N_10505);
nand U15054 (N_15054,N_11024,N_10049);
or U15055 (N_15055,N_10757,N_10685);
and U15056 (N_15056,N_10778,N_9456);
or U15057 (N_15057,N_12362,N_11444);
and U15058 (N_15058,N_11024,N_11106);
nand U15059 (N_15059,N_10187,N_11959);
nor U15060 (N_15060,N_9723,N_11317);
nand U15061 (N_15061,N_11939,N_12414);
and U15062 (N_15062,N_12435,N_10874);
xnor U15063 (N_15063,N_12357,N_10450);
nor U15064 (N_15064,N_10494,N_10427);
nand U15065 (N_15065,N_9502,N_10514);
nor U15066 (N_15066,N_11029,N_11863);
and U15067 (N_15067,N_9627,N_11493);
nor U15068 (N_15068,N_11340,N_11855);
or U15069 (N_15069,N_11724,N_10655);
and U15070 (N_15070,N_11663,N_11355);
nand U15071 (N_15071,N_11656,N_9903);
nand U15072 (N_15072,N_11481,N_11534);
or U15073 (N_15073,N_10963,N_10804);
nor U15074 (N_15074,N_11881,N_10688);
nor U15075 (N_15075,N_10029,N_11307);
nand U15076 (N_15076,N_11645,N_9640);
and U15077 (N_15077,N_11645,N_11895);
nor U15078 (N_15078,N_10867,N_9777);
or U15079 (N_15079,N_10366,N_10173);
nand U15080 (N_15080,N_10823,N_10211);
nor U15081 (N_15081,N_9925,N_12084);
xor U15082 (N_15082,N_10502,N_11207);
and U15083 (N_15083,N_9643,N_11658);
nor U15084 (N_15084,N_10654,N_11521);
and U15085 (N_15085,N_11226,N_12121);
or U15086 (N_15086,N_10321,N_10550);
nand U15087 (N_15087,N_9628,N_9753);
or U15088 (N_15088,N_11909,N_10165);
nor U15089 (N_15089,N_11102,N_10869);
and U15090 (N_15090,N_9993,N_9447);
nor U15091 (N_15091,N_10615,N_11660);
xnor U15092 (N_15092,N_9657,N_10270);
nand U15093 (N_15093,N_11987,N_12247);
or U15094 (N_15094,N_11139,N_11182);
and U15095 (N_15095,N_11938,N_10199);
nor U15096 (N_15096,N_11536,N_12074);
nor U15097 (N_15097,N_11629,N_12063);
nand U15098 (N_15098,N_10517,N_12454);
and U15099 (N_15099,N_10139,N_11406);
nor U15100 (N_15100,N_10019,N_9670);
nor U15101 (N_15101,N_10125,N_10959);
nand U15102 (N_15102,N_10605,N_11260);
xor U15103 (N_15103,N_11403,N_11939);
nor U15104 (N_15104,N_9638,N_12052);
nor U15105 (N_15105,N_10307,N_12404);
or U15106 (N_15106,N_9661,N_9431);
nand U15107 (N_15107,N_10662,N_10443);
xnor U15108 (N_15108,N_10299,N_11266);
and U15109 (N_15109,N_9670,N_10362);
and U15110 (N_15110,N_9735,N_11179);
or U15111 (N_15111,N_11574,N_12041);
and U15112 (N_15112,N_12360,N_9629);
or U15113 (N_15113,N_11367,N_12221);
and U15114 (N_15114,N_11491,N_10099);
nor U15115 (N_15115,N_10537,N_10954);
nor U15116 (N_15116,N_10328,N_9741);
nor U15117 (N_15117,N_9484,N_9696);
or U15118 (N_15118,N_11136,N_10767);
xor U15119 (N_15119,N_11183,N_12427);
and U15120 (N_15120,N_11484,N_11541);
or U15121 (N_15121,N_11961,N_12361);
nand U15122 (N_15122,N_11156,N_10059);
nand U15123 (N_15123,N_10510,N_11186);
nand U15124 (N_15124,N_10456,N_10314);
nand U15125 (N_15125,N_10679,N_11297);
and U15126 (N_15126,N_10099,N_9442);
nand U15127 (N_15127,N_10355,N_9843);
and U15128 (N_15128,N_11836,N_11320);
nand U15129 (N_15129,N_10318,N_10129);
or U15130 (N_15130,N_10584,N_9804);
nand U15131 (N_15131,N_10772,N_9428);
nand U15132 (N_15132,N_9905,N_9708);
nand U15133 (N_15133,N_11465,N_10407);
and U15134 (N_15134,N_11965,N_12259);
nor U15135 (N_15135,N_9375,N_9585);
and U15136 (N_15136,N_12334,N_11873);
or U15137 (N_15137,N_11970,N_11460);
or U15138 (N_15138,N_9681,N_9736);
nor U15139 (N_15139,N_11856,N_9722);
nand U15140 (N_15140,N_11595,N_9717);
nand U15141 (N_15141,N_11157,N_12294);
nor U15142 (N_15142,N_11823,N_11310);
nand U15143 (N_15143,N_11180,N_9670);
xor U15144 (N_15144,N_10464,N_9849);
nand U15145 (N_15145,N_11498,N_10031);
and U15146 (N_15146,N_9812,N_11339);
or U15147 (N_15147,N_10183,N_10066);
nand U15148 (N_15148,N_11443,N_10428);
and U15149 (N_15149,N_10649,N_10128);
nor U15150 (N_15150,N_10659,N_10640);
xor U15151 (N_15151,N_9586,N_12376);
or U15152 (N_15152,N_10282,N_9496);
or U15153 (N_15153,N_10051,N_10332);
nor U15154 (N_15154,N_10677,N_12092);
nand U15155 (N_15155,N_11004,N_12391);
nand U15156 (N_15156,N_12128,N_12215);
and U15157 (N_15157,N_12281,N_11192);
nor U15158 (N_15158,N_10991,N_9700);
nand U15159 (N_15159,N_10177,N_12234);
nor U15160 (N_15160,N_11381,N_10247);
nor U15161 (N_15161,N_9633,N_10066);
nand U15162 (N_15162,N_11017,N_11903);
or U15163 (N_15163,N_10003,N_10565);
and U15164 (N_15164,N_11397,N_10916);
xnor U15165 (N_15165,N_12296,N_11343);
nor U15166 (N_15166,N_11796,N_9955);
or U15167 (N_15167,N_10207,N_12339);
xor U15168 (N_15168,N_11094,N_12118);
and U15169 (N_15169,N_12316,N_12074);
and U15170 (N_15170,N_12273,N_9895);
or U15171 (N_15171,N_10212,N_10190);
xor U15172 (N_15172,N_10511,N_9571);
nand U15173 (N_15173,N_9621,N_10487);
nor U15174 (N_15174,N_11572,N_10103);
nand U15175 (N_15175,N_10948,N_10647);
nor U15176 (N_15176,N_12170,N_11681);
nand U15177 (N_15177,N_11148,N_10922);
and U15178 (N_15178,N_11783,N_10167);
nor U15179 (N_15179,N_11108,N_12338);
and U15180 (N_15180,N_12390,N_10893);
or U15181 (N_15181,N_10532,N_12429);
nand U15182 (N_15182,N_11766,N_11858);
nor U15183 (N_15183,N_12376,N_10219);
or U15184 (N_15184,N_10927,N_11321);
xnor U15185 (N_15185,N_9988,N_12349);
nor U15186 (N_15186,N_9865,N_10959);
nor U15187 (N_15187,N_9816,N_10215);
xnor U15188 (N_15188,N_11017,N_11032);
or U15189 (N_15189,N_12135,N_11085);
and U15190 (N_15190,N_10872,N_10064);
or U15191 (N_15191,N_10183,N_12269);
nor U15192 (N_15192,N_11007,N_10662);
nand U15193 (N_15193,N_11296,N_12246);
xnor U15194 (N_15194,N_10236,N_10908);
or U15195 (N_15195,N_10373,N_10993);
nor U15196 (N_15196,N_10079,N_10811);
and U15197 (N_15197,N_10192,N_9712);
nor U15198 (N_15198,N_11175,N_10408);
nand U15199 (N_15199,N_11895,N_9811);
xor U15200 (N_15200,N_9886,N_10664);
nor U15201 (N_15201,N_12100,N_10976);
xnor U15202 (N_15202,N_9506,N_12129);
or U15203 (N_15203,N_12442,N_9919);
and U15204 (N_15204,N_10945,N_11508);
nor U15205 (N_15205,N_9830,N_10673);
or U15206 (N_15206,N_11947,N_12330);
or U15207 (N_15207,N_11154,N_11348);
and U15208 (N_15208,N_11728,N_12122);
and U15209 (N_15209,N_10883,N_11285);
nand U15210 (N_15210,N_11898,N_9837);
nand U15211 (N_15211,N_10282,N_10387);
xnor U15212 (N_15212,N_9748,N_11459);
nand U15213 (N_15213,N_11638,N_11784);
nor U15214 (N_15214,N_10835,N_11011);
nor U15215 (N_15215,N_10129,N_12257);
xor U15216 (N_15216,N_10323,N_9534);
nand U15217 (N_15217,N_11579,N_9702);
nand U15218 (N_15218,N_12076,N_11444);
and U15219 (N_15219,N_10636,N_11480);
and U15220 (N_15220,N_11195,N_9557);
or U15221 (N_15221,N_11297,N_10085);
and U15222 (N_15222,N_10356,N_11049);
nand U15223 (N_15223,N_11522,N_10012);
nor U15224 (N_15224,N_9414,N_11010);
nor U15225 (N_15225,N_12383,N_10991);
and U15226 (N_15226,N_10620,N_10492);
nor U15227 (N_15227,N_12485,N_10864);
nor U15228 (N_15228,N_9829,N_9642);
nand U15229 (N_15229,N_10447,N_12288);
or U15230 (N_15230,N_10573,N_9718);
or U15231 (N_15231,N_11063,N_11578);
nor U15232 (N_15232,N_12039,N_12161);
or U15233 (N_15233,N_10314,N_11777);
or U15234 (N_15234,N_12304,N_11753);
and U15235 (N_15235,N_10644,N_10271);
nor U15236 (N_15236,N_12330,N_10863);
and U15237 (N_15237,N_12227,N_12115);
nor U15238 (N_15238,N_11732,N_9869);
nor U15239 (N_15239,N_12333,N_11893);
and U15240 (N_15240,N_10739,N_12161);
or U15241 (N_15241,N_11815,N_11442);
or U15242 (N_15242,N_12075,N_11622);
or U15243 (N_15243,N_9402,N_9858);
xor U15244 (N_15244,N_12429,N_10662);
and U15245 (N_15245,N_10148,N_12095);
nand U15246 (N_15246,N_10723,N_10358);
nor U15247 (N_15247,N_10175,N_10902);
nor U15248 (N_15248,N_10454,N_10592);
nand U15249 (N_15249,N_10294,N_9461);
xnor U15250 (N_15250,N_9424,N_9713);
nand U15251 (N_15251,N_12019,N_11599);
or U15252 (N_15252,N_11912,N_11192);
nand U15253 (N_15253,N_9791,N_11921);
nand U15254 (N_15254,N_11279,N_9598);
nor U15255 (N_15255,N_11554,N_10392);
nor U15256 (N_15256,N_10586,N_10482);
nand U15257 (N_15257,N_10194,N_10648);
or U15258 (N_15258,N_11139,N_11222);
xnor U15259 (N_15259,N_10366,N_11978);
nor U15260 (N_15260,N_10370,N_11945);
nor U15261 (N_15261,N_10122,N_12215);
and U15262 (N_15262,N_12441,N_9816);
and U15263 (N_15263,N_9585,N_9638);
xor U15264 (N_15264,N_9378,N_9570);
xor U15265 (N_15265,N_11000,N_9800);
xor U15266 (N_15266,N_9880,N_10137);
and U15267 (N_15267,N_10452,N_10381);
nand U15268 (N_15268,N_11644,N_11430);
nor U15269 (N_15269,N_12017,N_9422);
xor U15270 (N_15270,N_9787,N_9999);
nor U15271 (N_15271,N_12038,N_9490);
nor U15272 (N_15272,N_9956,N_9556);
nor U15273 (N_15273,N_10142,N_11608);
xnor U15274 (N_15274,N_10790,N_11485);
xor U15275 (N_15275,N_10268,N_12492);
nand U15276 (N_15276,N_10611,N_9704);
or U15277 (N_15277,N_10273,N_10980);
nand U15278 (N_15278,N_10454,N_10439);
and U15279 (N_15279,N_12016,N_10823);
and U15280 (N_15280,N_10711,N_12197);
nand U15281 (N_15281,N_9530,N_12260);
and U15282 (N_15282,N_10835,N_9525);
xnor U15283 (N_15283,N_10703,N_12078);
nand U15284 (N_15284,N_10967,N_12488);
nand U15285 (N_15285,N_10641,N_10815);
nand U15286 (N_15286,N_9952,N_12444);
xor U15287 (N_15287,N_11574,N_12190);
nand U15288 (N_15288,N_11556,N_12073);
nand U15289 (N_15289,N_11604,N_12237);
nand U15290 (N_15290,N_11973,N_11551);
and U15291 (N_15291,N_12381,N_10476);
nand U15292 (N_15292,N_11166,N_10354);
and U15293 (N_15293,N_11691,N_10605);
nand U15294 (N_15294,N_10442,N_11810);
nand U15295 (N_15295,N_11388,N_11396);
nor U15296 (N_15296,N_11231,N_11911);
and U15297 (N_15297,N_12104,N_11236);
nor U15298 (N_15298,N_11708,N_9442);
or U15299 (N_15299,N_11979,N_12143);
nand U15300 (N_15300,N_11000,N_10001);
or U15301 (N_15301,N_10839,N_9648);
nand U15302 (N_15302,N_9529,N_12319);
nor U15303 (N_15303,N_10491,N_9797);
and U15304 (N_15304,N_9947,N_9573);
nand U15305 (N_15305,N_11317,N_12195);
and U15306 (N_15306,N_9830,N_10839);
nand U15307 (N_15307,N_11897,N_10146);
or U15308 (N_15308,N_10639,N_11934);
nand U15309 (N_15309,N_9864,N_12107);
nand U15310 (N_15310,N_12259,N_10291);
or U15311 (N_15311,N_12002,N_11535);
and U15312 (N_15312,N_11842,N_10611);
nand U15313 (N_15313,N_10280,N_10826);
and U15314 (N_15314,N_10411,N_11381);
and U15315 (N_15315,N_12437,N_9631);
nor U15316 (N_15316,N_9832,N_11200);
nand U15317 (N_15317,N_11391,N_11276);
nor U15318 (N_15318,N_12165,N_9611);
or U15319 (N_15319,N_9694,N_9761);
or U15320 (N_15320,N_11658,N_12435);
nand U15321 (N_15321,N_11742,N_12051);
or U15322 (N_15322,N_9584,N_9654);
nand U15323 (N_15323,N_11153,N_10913);
xor U15324 (N_15324,N_9747,N_12230);
or U15325 (N_15325,N_10483,N_10705);
or U15326 (N_15326,N_10023,N_11223);
nand U15327 (N_15327,N_11638,N_11601);
xor U15328 (N_15328,N_11866,N_11277);
nor U15329 (N_15329,N_11250,N_12416);
or U15330 (N_15330,N_10364,N_10890);
nor U15331 (N_15331,N_10081,N_10555);
nand U15332 (N_15332,N_10551,N_11098);
and U15333 (N_15333,N_10031,N_9694);
nor U15334 (N_15334,N_9659,N_9911);
nand U15335 (N_15335,N_11129,N_11913);
and U15336 (N_15336,N_10395,N_10820);
nor U15337 (N_15337,N_12343,N_9503);
xnor U15338 (N_15338,N_11364,N_10756);
nand U15339 (N_15339,N_10501,N_10650);
nor U15340 (N_15340,N_11282,N_11765);
and U15341 (N_15341,N_11776,N_10187);
and U15342 (N_15342,N_11954,N_9941);
nor U15343 (N_15343,N_9789,N_12241);
nor U15344 (N_15344,N_10312,N_11322);
or U15345 (N_15345,N_10335,N_11476);
nand U15346 (N_15346,N_12425,N_11505);
nand U15347 (N_15347,N_10297,N_12399);
or U15348 (N_15348,N_11557,N_10086);
or U15349 (N_15349,N_11451,N_12105);
nor U15350 (N_15350,N_10022,N_12174);
and U15351 (N_15351,N_11450,N_9381);
and U15352 (N_15352,N_10131,N_10739);
or U15353 (N_15353,N_10613,N_9773);
nor U15354 (N_15354,N_12220,N_11292);
xnor U15355 (N_15355,N_11013,N_11508);
nor U15356 (N_15356,N_11819,N_11559);
nor U15357 (N_15357,N_9798,N_10512);
and U15358 (N_15358,N_9563,N_10814);
or U15359 (N_15359,N_12455,N_11532);
nor U15360 (N_15360,N_10196,N_11415);
nor U15361 (N_15361,N_10485,N_10522);
and U15362 (N_15362,N_12214,N_10261);
nand U15363 (N_15363,N_11370,N_10051);
or U15364 (N_15364,N_12228,N_12298);
or U15365 (N_15365,N_9823,N_12410);
or U15366 (N_15366,N_11347,N_12343);
xor U15367 (N_15367,N_9827,N_12351);
nor U15368 (N_15368,N_11261,N_12120);
nand U15369 (N_15369,N_12476,N_11202);
xor U15370 (N_15370,N_11835,N_11840);
and U15371 (N_15371,N_10801,N_11487);
nand U15372 (N_15372,N_10762,N_12064);
xnor U15373 (N_15373,N_10275,N_12213);
or U15374 (N_15374,N_9522,N_9562);
and U15375 (N_15375,N_12268,N_10349);
nor U15376 (N_15376,N_11469,N_11456);
nand U15377 (N_15377,N_11538,N_9615);
and U15378 (N_15378,N_10832,N_12421);
or U15379 (N_15379,N_11003,N_10798);
or U15380 (N_15380,N_11750,N_12222);
or U15381 (N_15381,N_11236,N_9723);
nor U15382 (N_15382,N_9695,N_10658);
nor U15383 (N_15383,N_10196,N_11498);
or U15384 (N_15384,N_9770,N_10961);
and U15385 (N_15385,N_12218,N_9851);
and U15386 (N_15386,N_11707,N_11541);
and U15387 (N_15387,N_11282,N_12258);
and U15388 (N_15388,N_12383,N_10705);
or U15389 (N_15389,N_12019,N_10170);
nand U15390 (N_15390,N_11114,N_9573);
xnor U15391 (N_15391,N_10293,N_10969);
and U15392 (N_15392,N_12136,N_11564);
xnor U15393 (N_15393,N_12097,N_10440);
nand U15394 (N_15394,N_10735,N_12256);
or U15395 (N_15395,N_12020,N_12107);
or U15396 (N_15396,N_9497,N_12033);
or U15397 (N_15397,N_9694,N_11208);
and U15398 (N_15398,N_9779,N_11186);
nor U15399 (N_15399,N_10403,N_10471);
nand U15400 (N_15400,N_10532,N_10767);
nor U15401 (N_15401,N_11000,N_9725);
nor U15402 (N_15402,N_9918,N_10290);
nor U15403 (N_15403,N_11951,N_9778);
and U15404 (N_15404,N_11094,N_9989);
or U15405 (N_15405,N_9637,N_11783);
and U15406 (N_15406,N_11528,N_11910);
nand U15407 (N_15407,N_9578,N_12374);
nor U15408 (N_15408,N_11467,N_11191);
xnor U15409 (N_15409,N_10465,N_11489);
or U15410 (N_15410,N_12436,N_11204);
nor U15411 (N_15411,N_10572,N_11194);
nand U15412 (N_15412,N_10149,N_9568);
or U15413 (N_15413,N_10924,N_11044);
or U15414 (N_15414,N_11228,N_9607);
nand U15415 (N_15415,N_9481,N_10438);
nor U15416 (N_15416,N_9754,N_12117);
nor U15417 (N_15417,N_11061,N_10050);
or U15418 (N_15418,N_11432,N_10951);
or U15419 (N_15419,N_10261,N_12282);
nor U15420 (N_15420,N_11122,N_11432);
xor U15421 (N_15421,N_9847,N_11379);
nor U15422 (N_15422,N_10818,N_11684);
and U15423 (N_15423,N_10910,N_10011);
nor U15424 (N_15424,N_10317,N_11556);
nor U15425 (N_15425,N_9708,N_10258);
nand U15426 (N_15426,N_10491,N_12117);
nand U15427 (N_15427,N_12359,N_9688);
and U15428 (N_15428,N_11820,N_10749);
xnor U15429 (N_15429,N_11472,N_9520);
nand U15430 (N_15430,N_9880,N_12438);
or U15431 (N_15431,N_10429,N_9569);
xor U15432 (N_15432,N_12415,N_10715);
or U15433 (N_15433,N_10295,N_11904);
and U15434 (N_15434,N_12029,N_10971);
and U15435 (N_15435,N_9978,N_11575);
and U15436 (N_15436,N_11053,N_10103);
nor U15437 (N_15437,N_12073,N_11788);
and U15438 (N_15438,N_12032,N_9499);
and U15439 (N_15439,N_10352,N_11212);
nand U15440 (N_15440,N_12040,N_11657);
and U15441 (N_15441,N_9554,N_10580);
nor U15442 (N_15442,N_11285,N_11309);
and U15443 (N_15443,N_9816,N_11361);
nor U15444 (N_15444,N_12452,N_10866);
xnor U15445 (N_15445,N_9612,N_10614);
nor U15446 (N_15446,N_11395,N_11879);
nor U15447 (N_15447,N_11121,N_12431);
xnor U15448 (N_15448,N_9761,N_11478);
nand U15449 (N_15449,N_10274,N_12432);
or U15450 (N_15450,N_11498,N_9850);
or U15451 (N_15451,N_10008,N_9657);
or U15452 (N_15452,N_12021,N_11699);
or U15453 (N_15453,N_10358,N_11504);
nor U15454 (N_15454,N_10865,N_10274);
or U15455 (N_15455,N_10557,N_10131);
or U15456 (N_15456,N_9950,N_12196);
and U15457 (N_15457,N_12414,N_11025);
and U15458 (N_15458,N_12432,N_10267);
or U15459 (N_15459,N_11718,N_12238);
nor U15460 (N_15460,N_10781,N_11673);
nand U15461 (N_15461,N_10928,N_10918);
nand U15462 (N_15462,N_12167,N_9641);
or U15463 (N_15463,N_12183,N_9649);
and U15464 (N_15464,N_12210,N_9996);
xnor U15465 (N_15465,N_11926,N_11978);
or U15466 (N_15466,N_10726,N_9591);
nand U15467 (N_15467,N_11385,N_11680);
nand U15468 (N_15468,N_11721,N_9973);
or U15469 (N_15469,N_9837,N_9811);
nor U15470 (N_15470,N_10394,N_10833);
nand U15471 (N_15471,N_9900,N_10578);
nand U15472 (N_15472,N_10573,N_10449);
or U15473 (N_15473,N_12420,N_9945);
xor U15474 (N_15474,N_12471,N_10189);
nor U15475 (N_15475,N_11261,N_12281);
nand U15476 (N_15476,N_10995,N_11041);
nand U15477 (N_15477,N_9823,N_12337);
xor U15478 (N_15478,N_11697,N_10445);
nand U15479 (N_15479,N_10646,N_12203);
or U15480 (N_15480,N_9391,N_11291);
nand U15481 (N_15481,N_9663,N_12008);
and U15482 (N_15482,N_10922,N_9511);
nor U15483 (N_15483,N_9881,N_12036);
nor U15484 (N_15484,N_10845,N_10403);
or U15485 (N_15485,N_11860,N_10833);
nand U15486 (N_15486,N_9982,N_11355);
and U15487 (N_15487,N_10114,N_9891);
or U15488 (N_15488,N_12105,N_11185);
or U15489 (N_15489,N_10533,N_9976);
and U15490 (N_15490,N_11473,N_10330);
nand U15491 (N_15491,N_9965,N_12141);
nor U15492 (N_15492,N_11070,N_10239);
nand U15493 (N_15493,N_9749,N_9969);
nor U15494 (N_15494,N_11113,N_10751);
and U15495 (N_15495,N_12274,N_9718);
xnor U15496 (N_15496,N_9422,N_9580);
nor U15497 (N_15497,N_11494,N_10185);
nand U15498 (N_15498,N_12434,N_10507);
nand U15499 (N_15499,N_12233,N_11442);
and U15500 (N_15500,N_10753,N_10308);
nor U15501 (N_15501,N_9697,N_12103);
or U15502 (N_15502,N_10693,N_9563);
or U15503 (N_15503,N_11819,N_10152);
nand U15504 (N_15504,N_12319,N_10564);
nor U15505 (N_15505,N_11530,N_11591);
nor U15506 (N_15506,N_10497,N_10134);
nor U15507 (N_15507,N_11989,N_9805);
nand U15508 (N_15508,N_11276,N_9810);
and U15509 (N_15509,N_11141,N_10173);
xor U15510 (N_15510,N_9839,N_10592);
nor U15511 (N_15511,N_12332,N_12055);
and U15512 (N_15512,N_10361,N_11970);
nor U15513 (N_15513,N_11849,N_11672);
nand U15514 (N_15514,N_9550,N_11939);
or U15515 (N_15515,N_9766,N_12233);
and U15516 (N_15516,N_11034,N_11328);
or U15517 (N_15517,N_11567,N_10846);
and U15518 (N_15518,N_11128,N_11985);
xor U15519 (N_15519,N_11942,N_12035);
or U15520 (N_15520,N_11046,N_9935);
or U15521 (N_15521,N_10652,N_10993);
nor U15522 (N_15522,N_9463,N_11078);
nor U15523 (N_15523,N_12396,N_11986);
or U15524 (N_15524,N_9650,N_12161);
and U15525 (N_15525,N_9990,N_9925);
nor U15526 (N_15526,N_10879,N_11811);
or U15527 (N_15527,N_11361,N_11076);
and U15528 (N_15528,N_11271,N_9546);
nor U15529 (N_15529,N_10737,N_11887);
or U15530 (N_15530,N_9483,N_11141);
nor U15531 (N_15531,N_11530,N_10732);
xor U15532 (N_15532,N_12473,N_10250);
nor U15533 (N_15533,N_10170,N_10827);
and U15534 (N_15534,N_9690,N_11216);
nor U15535 (N_15535,N_11670,N_9693);
or U15536 (N_15536,N_10401,N_9974);
nand U15537 (N_15537,N_9516,N_11677);
nand U15538 (N_15538,N_11382,N_9874);
xnor U15539 (N_15539,N_10547,N_11722);
xor U15540 (N_15540,N_10200,N_12068);
nand U15541 (N_15541,N_9855,N_9463);
nand U15542 (N_15542,N_11896,N_10012);
xor U15543 (N_15543,N_11610,N_11341);
nor U15544 (N_15544,N_10058,N_12209);
nor U15545 (N_15545,N_9789,N_9563);
nand U15546 (N_15546,N_11450,N_12464);
nor U15547 (N_15547,N_9757,N_11443);
nand U15548 (N_15548,N_10541,N_12378);
and U15549 (N_15549,N_9700,N_11925);
nor U15550 (N_15550,N_9681,N_11048);
and U15551 (N_15551,N_11765,N_10067);
nor U15552 (N_15552,N_9593,N_10631);
or U15553 (N_15553,N_10366,N_10039);
or U15554 (N_15554,N_10628,N_10160);
or U15555 (N_15555,N_10188,N_11655);
and U15556 (N_15556,N_11618,N_10223);
nand U15557 (N_15557,N_10355,N_10395);
nand U15558 (N_15558,N_10697,N_10207);
and U15559 (N_15559,N_11398,N_12182);
nor U15560 (N_15560,N_9961,N_10624);
nand U15561 (N_15561,N_9559,N_11138);
or U15562 (N_15562,N_9899,N_9550);
and U15563 (N_15563,N_12413,N_11733);
nor U15564 (N_15564,N_12248,N_11288);
nand U15565 (N_15565,N_9811,N_11278);
nand U15566 (N_15566,N_9514,N_9478);
nor U15567 (N_15567,N_10672,N_12075);
xor U15568 (N_15568,N_9847,N_9413);
xor U15569 (N_15569,N_11671,N_9635);
nand U15570 (N_15570,N_10723,N_11865);
nor U15571 (N_15571,N_12141,N_11090);
nand U15572 (N_15572,N_9823,N_11601);
xnor U15573 (N_15573,N_9995,N_10920);
nand U15574 (N_15574,N_11825,N_9911);
and U15575 (N_15575,N_12074,N_11244);
or U15576 (N_15576,N_11411,N_12369);
and U15577 (N_15577,N_10624,N_11307);
nor U15578 (N_15578,N_11688,N_9636);
and U15579 (N_15579,N_10044,N_9552);
and U15580 (N_15580,N_9507,N_9935);
nor U15581 (N_15581,N_9995,N_12137);
nand U15582 (N_15582,N_9474,N_12300);
or U15583 (N_15583,N_10222,N_11345);
or U15584 (N_15584,N_10722,N_11698);
nand U15585 (N_15585,N_11351,N_12237);
nor U15586 (N_15586,N_9849,N_11154);
or U15587 (N_15587,N_10932,N_10826);
nand U15588 (N_15588,N_10583,N_11473);
xor U15589 (N_15589,N_9425,N_11963);
or U15590 (N_15590,N_11206,N_10465);
nand U15591 (N_15591,N_11268,N_12251);
or U15592 (N_15592,N_9659,N_11953);
nor U15593 (N_15593,N_11776,N_12444);
nand U15594 (N_15594,N_10578,N_11408);
nand U15595 (N_15595,N_11738,N_11762);
and U15596 (N_15596,N_10653,N_10500);
and U15597 (N_15597,N_11572,N_9508);
or U15598 (N_15598,N_12193,N_11967);
or U15599 (N_15599,N_11458,N_12380);
nand U15600 (N_15600,N_11685,N_12386);
nand U15601 (N_15601,N_11345,N_11004);
nand U15602 (N_15602,N_9811,N_10915);
or U15603 (N_15603,N_11335,N_11223);
and U15604 (N_15604,N_12028,N_11708);
or U15605 (N_15605,N_10742,N_11376);
or U15606 (N_15606,N_11917,N_12043);
nor U15607 (N_15607,N_9737,N_9939);
or U15608 (N_15608,N_10549,N_10070);
and U15609 (N_15609,N_10071,N_11396);
nor U15610 (N_15610,N_12148,N_12101);
or U15611 (N_15611,N_12161,N_10839);
or U15612 (N_15612,N_10827,N_12267);
and U15613 (N_15613,N_9864,N_10474);
and U15614 (N_15614,N_10602,N_12106);
nor U15615 (N_15615,N_10444,N_11343);
or U15616 (N_15616,N_11722,N_10743);
xor U15617 (N_15617,N_10546,N_12054);
nor U15618 (N_15618,N_10483,N_11273);
nand U15619 (N_15619,N_10140,N_11616);
or U15620 (N_15620,N_10553,N_10454);
nand U15621 (N_15621,N_10168,N_12353);
xor U15622 (N_15622,N_12267,N_10873);
or U15623 (N_15623,N_10857,N_11438);
nand U15624 (N_15624,N_10345,N_11427);
and U15625 (N_15625,N_14366,N_13071);
nand U15626 (N_15626,N_14298,N_15588);
or U15627 (N_15627,N_13922,N_14467);
xnor U15628 (N_15628,N_12781,N_13285);
nand U15629 (N_15629,N_12961,N_14392);
nand U15630 (N_15630,N_14306,N_14312);
nor U15631 (N_15631,N_13727,N_15227);
nor U15632 (N_15632,N_13560,N_13959);
xor U15633 (N_15633,N_13620,N_13091);
xor U15634 (N_15634,N_12905,N_15578);
nor U15635 (N_15635,N_15048,N_15323);
nand U15636 (N_15636,N_12741,N_14864);
nor U15637 (N_15637,N_14035,N_13739);
or U15638 (N_15638,N_15601,N_14985);
or U15639 (N_15639,N_13543,N_14477);
and U15640 (N_15640,N_14523,N_13849);
nand U15641 (N_15641,N_13733,N_14791);
nand U15642 (N_15642,N_15326,N_13114);
and U15643 (N_15643,N_14607,N_15416);
and U15644 (N_15644,N_15112,N_14400);
nor U15645 (N_15645,N_14234,N_14066);
nor U15646 (N_15646,N_13540,N_13130);
nor U15647 (N_15647,N_14857,N_15447);
nor U15648 (N_15648,N_14819,N_13466);
nor U15649 (N_15649,N_13144,N_14484);
nor U15650 (N_15650,N_12582,N_14970);
nand U15651 (N_15651,N_14310,N_13578);
or U15652 (N_15652,N_14920,N_15493);
nand U15653 (N_15653,N_14517,N_13497);
nor U15654 (N_15654,N_15267,N_15296);
nor U15655 (N_15655,N_12856,N_12873);
and U15656 (N_15656,N_14789,N_13155);
xor U15657 (N_15657,N_13451,N_13381);
nor U15658 (N_15658,N_15341,N_15579);
nand U15659 (N_15659,N_14180,N_13268);
or U15660 (N_15660,N_15616,N_14759);
or U15661 (N_15661,N_12798,N_14058);
and U15662 (N_15662,N_14449,N_15314);
xnor U15663 (N_15663,N_13587,N_14338);
and U15664 (N_15664,N_14506,N_13845);
nand U15665 (N_15665,N_14629,N_13800);
nor U15666 (N_15666,N_14089,N_14596);
and U15667 (N_15667,N_14303,N_14588);
nor U15668 (N_15668,N_13713,N_13378);
nand U15669 (N_15669,N_15433,N_13397);
and U15670 (N_15670,N_14544,N_14918);
or U15671 (N_15671,N_13404,N_14377);
nor U15672 (N_15672,N_15014,N_13994);
or U15673 (N_15673,N_13810,N_15020);
xnor U15674 (N_15674,N_14885,N_14704);
nor U15675 (N_15675,N_12806,N_14228);
nor U15676 (N_15676,N_14829,N_13399);
nand U15677 (N_15677,N_14961,N_13847);
and U15678 (N_15678,N_15371,N_13401);
or U15679 (N_15679,N_13259,N_15186);
and U15680 (N_15680,N_13423,N_13140);
nand U15681 (N_15681,N_13177,N_13691);
and U15682 (N_15682,N_13877,N_14127);
and U15683 (N_15683,N_13914,N_12545);
nor U15684 (N_15684,N_13472,N_15556);
xnor U15685 (N_15685,N_12510,N_14581);
nand U15686 (N_15686,N_14179,N_15000);
nand U15687 (N_15687,N_13638,N_14602);
or U15688 (N_15688,N_12758,N_13671);
nand U15689 (N_15689,N_14094,N_14685);
or U15690 (N_15690,N_15511,N_14714);
and U15691 (N_15691,N_14380,N_15080);
and U15692 (N_15692,N_14945,N_15127);
or U15693 (N_15693,N_14824,N_14924);
or U15694 (N_15694,N_13848,N_14748);
or U15695 (N_15695,N_14069,N_14221);
and U15696 (N_15696,N_14988,N_13860);
nor U15697 (N_15697,N_14986,N_12503);
and U15698 (N_15698,N_14171,N_12818);
xnor U15699 (N_15699,N_15120,N_14135);
nor U15700 (N_15700,N_12943,N_13505);
or U15701 (N_15701,N_15185,N_15404);
nand U15702 (N_15702,N_14099,N_13106);
and U15703 (N_15703,N_14963,N_13371);
and U15704 (N_15704,N_14726,N_15161);
and U15705 (N_15705,N_14078,N_14816);
or U15706 (N_15706,N_15031,N_13115);
and U15707 (N_15707,N_14663,N_13876);
or U15708 (N_15708,N_13100,N_15436);
nand U15709 (N_15709,N_12765,N_15612);
nor U15710 (N_15710,N_13450,N_14440);
xnor U15711 (N_15711,N_14778,N_12524);
or U15712 (N_15712,N_14785,N_14533);
xor U15713 (N_15713,N_14060,N_14594);
and U15714 (N_15714,N_13042,N_15373);
nor U15715 (N_15715,N_13081,N_12960);
or U15716 (N_15716,N_12920,N_15295);
nor U15717 (N_15717,N_14508,N_13480);
nand U15718 (N_15718,N_14693,N_15402);
and U15719 (N_15719,N_14279,N_14855);
nor U15720 (N_15720,N_13495,N_15397);
nor U15721 (N_15721,N_13963,N_13303);
nor U15722 (N_15722,N_14048,N_14055);
xnor U15723 (N_15723,N_13416,N_13471);
xor U15724 (N_15724,N_12519,N_14503);
nand U15725 (N_15725,N_14110,N_15481);
nand U15726 (N_15726,N_13232,N_15568);
xor U15727 (N_15727,N_14585,N_14518);
xor U15728 (N_15728,N_14561,N_13723);
or U15729 (N_15729,N_15083,N_14223);
nand U15730 (N_15730,N_13324,N_15182);
nand U15731 (N_15731,N_12535,N_14790);
or U15732 (N_15732,N_15026,N_13946);
nand U15733 (N_15733,N_13536,N_13904);
and U15734 (N_15734,N_13780,N_14804);
nor U15735 (N_15735,N_14199,N_13169);
and U15736 (N_15736,N_14957,N_13007);
and U15737 (N_15737,N_14519,N_15223);
nor U15738 (N_15738,N_12608,N_15400);
or U15739 (N_15739,N_14765,N_14435);
or U15740 (N_15740,N_13768,N_15339);
nor U15741 (N_15741,N_15212,N_12505);
nor U15742 (N_15742,N_15074,N_13278);
nand U15743 (N_15743,N_15215,N_12542);
nor U15744 (N_15744,N_14619,N_13582);
xor U15745 (N_15745,N_14879,N_13917);
or U15746 (N_15746,N_15559,N_12565);
or U15747 (N_15747,N_15510,N_14526);
nand U15748 (N_15748,N_12755,N_13247);
and U15749 (N_15749,N_14631,N_13271);
xnor U15750 (N_15750,N_15123,N_12587);
and U15751 (N_15751,N_13297,N_13427);
nor U15752 (N_15752,N_14591,N_12773);
nand U15753 (N_15753,N_13288,N_14742);
and U15754 (N_15754,N_13193,N_13526);
or U15755 (N_15755,N_15265,N_13094);
and U15756 (N_15756,N_13120,N_13932);
xnor U15757 (N_15757,N_14256,N_14735);
nor U15758 (N_15758,N_13402,N_14948);
nor U15759 (N_15759,N_13788,N_14481);
xor U15760 (N_15760,N_12734,N_12779);
nor U15761 (N_15761,N_14955,N_12832);
or U15762 (N_15762,N_14427,N_12974);
and U15763 (N_15763,N_13892,N_13150);
xnor U15764 (N_15764,N_13444,N_14443);
xnor U15765 (N_15765,N_15624,N_12547);
or U15766 (N_15766,N_14661,N_13426);
xnor U15767 (N_15767,N_15505,N_15050);
nor U15768 (N_15768,N_14373,N_15130);
nand U15769 (N_15769,N_14243,N_14311);
or U15770 (N_15770,N_14401,N_14350);
xor U15771 (N_15771,N_14068,N_13327);
nor U15772 (N_15772,N_14067,N_14669);
xnor U15773 (N_15773,N_13901,N_15032);
nand U15774 (N_15774,N_15379,N_15536);
and U15775 (N_15775,N_14383,N_15527);
nand U15776 (N_15776,N_12944,N_14112);
nor U15777 (N_15777,N_13153,N_12667);
and U15778 (N_15778,N_12549,N_14091);
and U15779 (N_15779,N_13342,N_13368);
and U15780 (N_15780,N_13147,N_14173);
xor U15781 (N_15781,N_12539,N_15610);
nor U15782 (N_15782,N_13338,N_13846);
nand U15783 (N_15783,N_14198,N_15428);
and U15784 (N_15784,N_12924,N_14808);
nor U15785 (N_15785,N_15238,N_14903);
nor U15786 (N_15786,N_14584,N_13966);
and U15787 (N_15787,N_13189,N_13314);
nor U15788 (N_15788,N_12836,N_14321);
or U15789 (N_15789,N_14758,N_14784);
or U15790 (N_15790,N_15125,N_14387);
or U15791 (N_15791,N_13843,N_14589);
and U15792 (N_15792,N_15160,N_13119);
and U15793 (N_15793,N_12824,N_15446);
nand U15794 (N_15794,N_15158,N_14912);
nor U15795 (N_15795,N_13839,N_12704);
xnor U15796 (N_15796,N_14466,N_14910);
nand U15797 (N_15797,N_12727,N_13550);
or U15798 (N_15798,N_13801,N_13499);
nand U15799 (N_15799,N_14250,N_12701);
nor U15800 (N_15800,N_14160,N_15248);
nor U15801 (N_15801,N_14239,N_14844);
nor U15802 (N_15802,N_13601,N_12629);
nand U15803 (N_15803,N_12828,N_13659);
xor U15804 (N_15804,N_13011,N_14936);
xnor U15805 (N_15805,N_14488,N_14109);
and U15806 (N_15806,N_14026,N_14915);
or U15807 (N_15807,N_13136,N_12649);
nand U15808 (N_15808,N_13107,N_15514);
nor U15809 (N_15809,N_12590,N_13789);
nand U15810 (N_15810,N_13525,N_13139);
nor U15811 (N_15811,N_14952,N_15262);
and U15812 (N_15812,N_15599,N_14654);
and U15813 (N_15813,N_13455,N_14658);
xnor U15814 (N_15814,N_13750,N_14452);
nor U15815 (N_15815,N_15426,N_14143);
nand U15816 (N_15816,N_13057,N_13686);
and U15817 (N_15817,N_14231,N_13819);
and U15818 (N_15818,N_13977,N_13085);
or U15819 (N_15819,N_15487,N_14848);
xor U15820 (N_15820,N_14802,N_13175);
nand U15821 (N_15821,N_12511,N_15528);
and U15822 (N_15822,N_15051,N_12651);
xor U15823 (N_15823,N_13793,N_14153);
or U15824 (N_15824,N_13385,N_14684);
nor U15825 (N_15825,N_14429,N_14334);
or U15826 (N_15826,N_14733,N_13447);
and U15827 (N_15827,N_14932,N_13595);
nand U15828 (N_15828,N_14529,N_14140);
nor U15829 (N_15829,N_13369,N_14189);
and U15830 (N_15830,N_12558,N_13772);
nor U15831 (N_15831,N_14453,N_14556);
or U15832 (N_15832,N_13212,N_14299);
or U15833 (N_15833,N_14462,N_14005);
or U15834 (N_15834,N_13361,N_13850);
nand U15835 (N_15835,N_14079,N_14301);
nand U15836 (N_15836,N_12592,N_14723);
and U15837 (N_15837,N_14034,N_13056);
nor U15838 (N_15838,N_13710,N_15370);
or U15839 (N_15839,N_13571,N_14770);
nor U15840 (N_15840,N_13261,N_14624);
or U15841 (N_15841,N_14605,N_14205);
nand U15842 (N_15842,N_12949,N_13955);
or U15843 (N_15843,N_15219,N_12909);
nor U15844 (N_15844,N_15228,N_13448);
xnor U15845 (N_15845,N_15299,N_12866);
xor U15846 (N_15846,N_15623,N_13316);
xnor U15847 (N_15847,N_14761,N_15138);
nand U15848 (N_15848,N_14448,N_15194);
nor U15849 (N_15849,N_14725,N_14376);
and U15850 (N_15850,N_13438,N_13196);
nor U15851 (N_15851,N_15537,N_14323);
and U15852 (N_15852,N_15191,N_14870);
xnor U15853 (N_15853,N_13837,N_12712);
and U15854 (N_15854,N_14954,N_13317);
and U15855 (N_15855,N_13289,N_14768);
and U15856 (N_15856,N_12981,N_14474);
nor U15857 (N_15857,N_14928,N_12703);
nand U15858 (N_15858,N_12843,N_13854);
or U15859 (N_15859,N_15049,N_14973);
and U15860 (N_15860,N_14043,N_15438);
or U15861 (N_15861,N_14215,N_12681);
or U15862 (N_15862,N_13030,N_14064);
nor U15863 (N_15863,N_14989,N_13163);
nand U15864 (N_15864,N_14168,N_15357);
or U15865 (N_15865,N_13818,N_12795);
nor U15866 (N_15866,N_15254,N_14480);
and U15867 (N_15867,N_14357,N_13200);
and U15868 (N_15868,N_13320,N_14013);
nor U15869 (N_15869,N_14266,N_14015);
nand U15870 (N_15870,N_14465,N_14971);
nand U15871 (N_15871,N_14420,N_15259);
nand U15872 (N_15872,N_13964,N_14740);
nand U15873 (N_15873,N_15414,N_12994);
xnor U15874 (N_15874,N_15230,N_13015);
nor U15875 (N_15875,N_12841,N_14431);
nor U15876 (N_15876,N_15088,N_15427);
or U15877 (N_15877,N_12738,N_15022);
and U15878 (N_15878,N_14202,N_13240);
and U15879 (N_15879,N_14616,N_15177);
and U15880 (N_15880,N_14741,N_15021);
and U15881 (N_15881,N_15619,N_15197);
nor U15882 (N_15882,N_13012,N_13019);
nand U15883 (N_15883,N_12604,N_13044);
or U15884 (N_15884,N_15224,N_14317);
and U15885 (N_15885,N_14272,N_13611);
or U15886 (N_15886,N_13174,N_15434);
nor U15887 (N_15887,N_14563,N_14597);
nand U15888 (N_15888,N_15542,N_12840);
xnor U15889 (N_15889,N_13118,N_14627);
and U15890 (N_15890,N_12674,N_14391);
nand U15891 (N_15891,N_12713,N_12637);
nand U15892 (N_15892,N_14297,N_15007);
or U15893 (N_15893,N_14807,N_13386);
and U15894 (N_15894,N_12775,N_14913);
nor U15895 (N_15895,N_15270,N_12954);
or U15896 (N_15896,N_15498,N_13413);
nand U15897 (N_15897,N_12769,N_14536);
and U15898 (N_15898,N_13396,N_13952);
nand U15899 (N_15899,N_14100,N_13731);
and U15900 (N_15900,N_14372,N_15200);
nor U15901 (N_15901,N_14336,N_13476);
or U15902 (N_15902,N_15471,N_13999);
or U15903 (N_15903,N_14586,N_14660);
and U15904 (N_15904,N_15593,N_12751);
nand U15905 (N_15905,N_15236,N_14116);
or U15906 (N_15906,N_15253,N_12695);
nand U15907 (N_15907,N_15338,N_15569);
xor U15908 (N_15908,N_14417,N_14081);
and U15909 (N_15909,N_15024,N_13142);
and U15910 (N_15910,N_12710,N_15523);
xor U15911 (N_15911,N_15389,N_14780);
nor U15912 (N_15912,N_12980,N_15001);
or U15913 (N_15913,N_15363,N_15564);
nand U15914 (N_15914,N_14520,N_14224);
or U15915 (N_15915,N_12572,N_13421);
nor U15916 (N_15916,N_12585,N_14300);
and U15917 (N_15917,N_15199,N_14318);
or U15918 (N_15918,N_15292,N_14219);
nand U15919 (N_15919,N_12812,N_14027);
nor U15920 (N_15920,N_13292,N_15243);
nor U15921 (N_15921,N_14821,N_14246);
and U15922 (N_15922,N_14687,N_12569);
nor U15923 (N_15923,N_14138,N_13527);
and U15924 (N_15924,N_15278,N_15406);
nor U15925 (N_15925,N_15285,N_13834);
or U15926 (N_15926,N_15535,N_14502);
nor U15927 (N_15927,N_12707,N_12766);
nor U15928 (N_15928,N_14261,N_14834);
or U15929 (N_15929,N_13003,N_12846);
nand U15930 (N_15930,N_13009,N_12648);
nand U15931 (N_15931,N_14739,N_12692);
xnor U15932 (N_15932,N_13122,N_15480);
xnor U15933 (N_15933,N_14365,N_13254);
and U15934 (N_15934,N_13151,N_15055);
nor U15935 (N_15935,N_12537,N_13925);
or U15936 (N_15936,N_15245,N_13786);
and U15937 (N_15937,N_14269,N_15222);
nand U15938 (N_15938,N_14867,N_13111);
and U15939 (N_15939,N_12715,N_13006);
nand U15940 (N_15940,N_15166,N_13443);
nor U15941 (N_15941,N_13873,N_13300);
and U15942 (N_15942,N_15497,N_14262);
nor U15943 (N_15943,N_12627,N_14217);
xor U15944 (N_15944,N_15086,N_13634);
xor U15945 (N_15945,N_14419,N_14907);
nor U15946 (N_15946,N_13687,N_15269);
and U15947 (N_15947,N_12839,N_13208);
and U15948 (N_15948,N_15333,N_12679);
and U15949 (N_15949,N_15084,N_12670);
and U15950 (N_15950,N_12678,N_15068);
or U15951 (N_15951,N_14990,N_14017);
nand U15952 (N_15952,N_14233,N_13097);
nor U15953 (N_15953,N_14483,N_14032);
nand U15954 (N_15954,N_13531,N_14931);
and U15955 (N_15955,N_14037,N_14793);
nor U15956 (N_15956,N_13935,N_15101);
xnor U15957 (N_15957,N_15018,N_15067);
nand U15958 (N_15958,N_13123,N_13162);
nor U15959 (N_15959,N_13642,N_13102);
nand U15960 (N_15960,N_13522,N_15330);
nand U15961 (N_15961,N_13649,N_14884);
nor U15962 (N_15962,N_13475,N_13485);
and U15963 (N_15963,N_15597,N_14712);
nand U15964 (N_15964,N_14566,N_12928);
or U15965 (N_15965,N_14371,N_13166);
and U15966 (N_15966,N_13652,N_15264);
and U15967 (N_15967,N_13262,N_12984);
nand U15968 (N_15968,N_15283,N_14121);
or U15969 (N_15969,N_12801,N_13067);
nand U15970 (N_15970,N_15091,N_15143);
nand U15971 (N_15971,N_14264,N_14668);
or U15972 (N_15972,N_12906,N_15229);
nor U15973 (N_15973,N_14837,N_12952);
and U15974 (N_15974,N_15249,N_12816);
nand U15975 (N_15975,N_15411,N_15151);
nand U15976 (N_15976,N_14947,N_13812);
nand U15977 (N_15977,N_13370,N_13648);
and U15978 (N_15978,N_14291,N_13305);
nor U15979 (N_15979,N_14580,N_13781);
xor U15980 (N_15980,N_13047,N_12834);
nor U15981 (N_15981,N_12571,N_12730);
nand U15982 (N_15982,N_12936,N_14886);
or U15983 (N_15983,N_13972,N_14552);
nand U15984 (N_15984,N_14152,N_14806);
and U15985 (N_15985,N_12520,N_15211);
and U15986 (N_15986,N_14281,N_12686);
and U15987 (N_15987,N_14666,N_14088);
nor U15988 (N_15988,N_14118,N_13878);
nand U15989 (N_15989,N_15483,N_13243);
xnor U15990 (N_15990,N_13046,N_14252);
nor U15991 (N_15991,N_15316,N_14292);
and U15992 (N_15992,N_14894,N_15502);
nor U15993 (N_15993,N_14249,N_15298);
or U15994 (N_15994,N_15034,N_14274);
xor U15995 (N_15995,N_13830,N_13068);
xnor U15996 (N_15996,N_14329,N_12538);
and U15997 (N_15997,N_14331,N_12719);
xnor U15998 (N_15998,N_13941,N_14163);
or U15999 (N_15999,N_14701,N_14705);
xnor U16000 (N_16000,N_15512,N_13823);
and U16001 (N_16001,N_12525,N_13939);
nand U16002 (N_16002,N_13377,N_14941);
and U16003 (N_16003,N_13523,N_14413);
or U16004 (N_16004,N_15309,N_13950);
or U16005 (N_16005,N_14006,N_13027);
or U16006 (N_16006,N_13911,N_13520);
or U16007 (N_16007,N_15310,N_14286);
and U16008 (N_16008,N_14305,N_14461);
or U16009 (N_16009,N_14548,N_14958);
nand U16010 (N_16010,N_15008,N_15394);
nand U16011 (N_16011,N_13509,N_14113);
nor U16012 (N_16012,N_13753,N_14277);
xnor U16013 (N_16013,N_14464,N_12771);
and U16014 (N_16014,N_12642,N_15417);
and U16015 (N_16015,N_15170,N_15398);
nor U16016 (N_16016,N_12913,N_14782);
and U16017 (N_16017,N_13437,N_14547);
nor U16018 (N_16018,N_13641,N_12516);
and U16019 (N_16019,N_13871,N_14362);
nor U16020 (N_16020,N_15465,N_14996);
nor U16021 (N_16021,N_15079,N_15609);
nor U16022 (N_16022,N_15344,N_13609);
nand U16023 (N_16023,N_15257,N_14237);
nor U16024 (N_16024,N_13462,N_12743);
or U16025 (N_16025,N_12813,N_13050);
xnor U16026 (N_16026,N_14276,N_13429);
xor U16027 (N_16027,N_15365,N_13510);
nand U16028 (N_16028,N_13181,N_13202);
xnor U16029 (N_16029,N_12993,N_13924);
and U16030 (N_16030,N_15304,N_14917);
or U16031 (N_16031,N_13624,N_14630);
and U16032 (N_16032,N_15274,N_13586);
nor U16033 (N_16033,N_15521,N_14085);
nand U16034 (N_16034,N_14007,N_13063);
and U16035 (N_16035,N_15324,N_13422);
or U16036 (N_16036,N_15044,N_12698);
or U16037 (N_16037,N_12854,N_12857);
nor U16038 (N_16038,N_13734,N_14744);
xnor U16039 (N_16039,N_12521,N_14166);
nor U16040 (N_16040,N_12786,N_15146);
or U16041 (N_16041,N_12916,N_14812);
nand U16042 (N_16042,N_14368,N_14156);
xor U16043 (N_16043,N_13717,N_13299);
or U16044 (N_16044,N_13045,N_12646);
nand U16045 (N_16045,N_14516,N_14853);
and U16046 (N_16046,N_14137,N_13866);
or U16047 (N_16047,N_14888,N_15128);
nor U16048 (N_16048,N_12883,N_13746);
nor U16049 (N_16049,N_15327,N_13969);
or U16050 (N_16050,N_13528,N_14141);
and U16051 (N_16051,N_13362,N_15343);
nor U16052 (N_16052,N_14395,N_14841);
xor U16053 (N_16053,N_15477,N_12533);
xnor U16054 (N_16054,N_12838,N_15183);
and U16055 (N_16055,N_13754,N_14339);
or U16056 (N_16056,N_13929,N_14475);
nand U16057 (N_16057,N_12855,N_15155);
nand U16058 (N_16058,N_14571,N_13276);
nor U16059 (N_16059,N_12895,N_14593);
or U16060 (N_16060,N_15376,N_15322);
and U16061 (N_16061,N_14052,N_15572);
or U16062 (N_16062,N_13660,N_12787);
or U16063 (N_16063,N_13555,N_14889);
or U16064 (N_16064,N_13238,N_13726);
nand U16065 (N_16065,N_14460,N_13256);
nor U16066 (N_16066,N_13360,N_15456);
nand U16067 (N_16067,N_14437,N_14904);
and U16068 (N_16068,N_13529,N_15567);
nand U16069 (N_16069,N_13266,N_14218);
xor U16070 (N_16070,N_13055,N_13688);
and U16071 (N_16071,N_14590,N_14599);
nor U16072 (N_16072,N_13465,N_14805);
or U16073 (N_16073,N_14309,N_13542);
and U16074 (N_16074,N_13112,N_13198);
xor U16075 (N_16075,N_14325,N_14149);
nand U16076 (N_16076,N_14559,N_14846);
nor U16077 (N_16077,N_12872,N_14000);
and U16078 (N_16078,N_14105,N_14157);
and U16079 (N_16079,N_13061,N_14745);
nor U16080 (N_16080,N_12564,N_14898);
nand U16081 (N_16081,N_15287,N_13936);
and U16082 (N_16082,N_15172,N_12852);
nor U16083 (N_16083,N_14570,N_14598);
or U16084 (N_16084,N_15041,N_12782);
or U16085 (N_16085,N_13490,N_13249);
and U16086 (N_16086,N_15385,N_13241);
and U16087 (N_16087,N_13352,N_13889);
and U16088 (N_16088,N_14375,N_15149);
nand U16089 (N_16089,N_14746,N_13460);
and U16090 (N_16090,N_13026,N_15239);
or U16091 (N_16091,N_15503,N_14225);
and U16092 (N_16092,N_12939,N_13398);
nand U16093 (N_16093,N_12722,N_14639);
or U16094 (N_16094,N_13127,N_13204);
xor U16095 (N_16095,N_13219,N_12675);
nor U16096 (N_16096,N_14969,N_13530);
xor U16097 (N_16097,N_14956,N_13188);
xnor U16098 (N_16098,N_14022,N_13909);
and U16099 (N_16099,N_13383,N_15081);
or U16100 (N_16100,N_13947,N_14787);
or U16101 (N_16101,N_14978,N_12940);
nor U16102 (N_16102,N_13760,N_14410);
or U16103 (N_16103,N_13138,N_15336);
nor U16104 (N_16104,N_13103,N_12999);
and U16105 (N_16105,N_14489,N_12983);
and U16106 (N_16106,N_13692,N_15435);
nor U16107 (N_16107,N_15036,N_12986);
or U16108 (N_16108,N_15459,N_12885);
xor U16109 (N_16109,N_15378,N_13194);
and U16110 (N_16110,N_15017,N_13816);
or U16111 (N_16111,N_13425,N_12777);
and U16112 (N_16112,N_14749,N_13621);
nand U16113 (N_16113,N_14257,N_14938);
nand U16114 (N_16114,N_13514,N_15331);
nand U16115 (N_16115,N_13803,N_15563);
and U16116 (N_16116,N_12633,N_14734);
nand U16117 (N_16117,N_13956,N_12807);
xor U16118 (N_16118,N_14447,N_14169);
nand U16119 (N_16119,N_13513,N_14408);
and U16120 (N_16120,N_13738,N_12887);
or U16121 (N_16121,N_14470,N_14337);
nor U16122 (N_16122,N_15508,N_14747);
nand U16123 (N_16123,N_13867,N_12870);
nand U16124 (N_16124,N_12631,N_15175);
and U16125 (N_16125,N_14843,N_13137);
nor U16126 (N_16126,N_13814,N_15554);
nand U16127 (N_16127,N_14093,N_14933);
nor U16128 (N_16128,N_15504,N_13394);
nand U16129 (N_16129,N_13420,N_15082);
or U16130 (N_16130,N_14495,N_14942);
xor U16131 (N_16131,N_15190,N_15496);
nor U16132 (N_16132,N_15162,N_13517);
and U16133 (N_16133,N_14743,N_14513);
nand U16134 (N_16134,N_15110,N_14468);
and U16135 (N_16135,N_15256,N_15390);
and U16136 (N_16136,N_12979,N_12778);
nor U16137 (N_16137,N_15103,N_13636);
nand U16138 (N_16138,N_12596,N_14511);
and U16139 (N_16139,N_14111,N_15131);
xor U16140 (N_16140,N_14896,N_14865);
nor U16141 (N_16141,N_15188,N_13379);
and U16142 (N_16142,N_14909,N_13146);
xor U16143 (N_16143,N_12617,N_15543);
and U16144 (N_16144,N_13069,N_15437);
nand U16145 (N_16145,N_13461,N_15046);
xnor U16146 (N_16146,N_13716,N_13028);
xnor U16147 (N_16147,N_14866,N_13336);
or U16148 (N_16148,N_14695,N_13036);
or U16149 (N_16149,N_14409,N_14332);
nor U16150 (N_16150,N_12978,N_14101);
xnor U16151 (N_16151,N_15367,N_14324);
or U16152 (N_16152,N_13156,N_15541);
nand U16153 (N_16153,N_14119,N_12689);
and U16154 (N_16154,N_13680,N_13126);
nand U16155 (N_16155,N_12578,N_14550);
or U16156 (N_16156,N_12625,N_12515);
and U16157 (N_16157,N_12669,N_13173);
xor U16158 (N_16158,N_13874,N_15418);
nor U16159 (N_16159,N_13364,N_14355);
nand U16160 (N_16160,N_15090,N_12823);
or U16161 (N_16161,N_14905,N_14211);
nand U16162 (N_16162,N_13457,N_13318);
or U16163 (N_16163,N_13013,N_14498);
and U16164 (N_16164,N_13248,N_14708);
xnor U16165 (N_16165,N_13516,N_15142);
nand U16166 (N_16166,N_14432,N_14628);
and U16167 (N_16167,N_15028,N_13647);
and U16168 (N_16168,N_13431,N_15057);
or U16169 (N_16169,N_12829,N_15102);
nor U16170 (N_16170,N_12897,N_15405);
or U16171 (N_16171,N_14655,N_15561);
or U16172 (N_16172,N_14386,N_12969);
nand U16173 (N_16173,N_13223,N_12660);
nor U16174 (N_16174,N_15027,N_12507);
xnor U16175 (N_16175,N_13852,N_15126);
nor U16176 (N_16176,N_15509,N_15016);
or U16177 (N_16177,N_14875,N_14651);
nor U16178 (N_16178,N_15312,N_14018);
or U16179 (N_16179,N_13737,N_15425);
nor U16180 (N_16180,N_13694,N_13356);
and U16181 (N_16181,N_15294,N_14103);
nand U16182 (N_16182,N_15075,N_13343);
or U16183 (N_16183,N_12595,N_13617);
and U16184 (N_16184,N_15087,N_14906);
or U16185 (N_16185,N_12898,N_12601);
nand U16186 (N_16186,N_13838,N_13265);
and U16187 (N_16187,N_13868,N_12570);
nand U16188 (N_16188,N_15035,N_13366);
and U16189 (N_16189,N_13228,N_15002);
and U16190 (N_16190,N_15395,N_13294);
nor U16191 (N_16191,N_15407,N_14976);
nor U16192 (N_16192,N_13152,N_13921);
xor U16193 (N_16193,N_13224,N_13477);
nor U16194 (N_16194,N_12780,N_15450);
nor U16195 (N_16195,N_15280,N_14267);
nor U16196 (N_16196,N_13668,N_14681);
nand U16197 (N_16197,N_13575,N_13961);
and U16198 (N_16198,N_13410,N_13086);
nand U16199 (N_16199,N_13728,N_14456);
nand U16200 (N_16200,N_13333,N_13863);
nor U16201 (N_16201,N_13469,N_13785);
and U16202 (N_16202,N_12502,N_14084);
or U16203 (N_16203,N_14194,N_13557);
nor U16204 (N_16204,N_15058,N_13065);
nor U16205 (N_16205,N_15513,N_14186);
nand U16206 (N_16206,N_13905,N_14776);
nor U16207 (N_16207,N_13489,N_15460);
nand U16208 (N_16208,N_15607,N_13991);
and U16209 (N_16209,N_14302,N_14428);
nor U16210 (N_16210,N_14117,N_13931);
nor U16211 (N_16211,N_14540,N_14108);
nand U16212 (N_16212,N_14345,N_13337);
nor U16213 (N_16213,N_14063,N_13987);
or U16214 (N_16214,N_12757,N_15105);
or U16215 (N_16215,N_12725,N_13521);
nor U16216 (N_16216,N_14680,N_14949);
nand U16217 (N_16217,N_14728,N_12517);
and U16218 (N_16218,N_14455,N_13574);
nand U16219 (N_16219,N_15360,N_14263);
nand U16220 (N_16220,N_14679,N_14736);
or U16221 (N_16221,N_14767,N_15488);
and U16222 (N_16222,N_12975,N_14051);
nand U16223 (N_16223,N_13488,N_13709);
or U16224 (N_16224,N_13658,N_14342);
or U16225 (N_16225,N_15251,N_14557);
and U16226 (N_16226,N_13408,N_12788);
and U16227 (N_16227,N_13762,N_14177);
and U16228 (N_16228,N_14213,N_14322);
nor U16229 (N_16229,N_14874,N_14283);
and U16230 (N_16230,N_14568,N_14175);
and U16231 (N_16231,N_14344,N_15121);
nor U16232 (N_16232,N_13957,N_13246);
or U16233 (N_16233,N_14095,N_14703);
nand U16234 (N_16234,N_13888,N_14777);
or U16235 (N_16235,N_13345,N_14147);
or U16236 (N_16236,N_13417,N_14828);
nand U16237 (N_16237,N_15134,N_13831);
and U16238 (N_16238,N_14053,N_12536);
nand U16239 (N_16239,N_13896,N_13724);
nor U16240 (N_16240,N_13664,N_13784);
nor U16241 (N_16241,N_15605,N_14831);
nor U16242 (N_16242,N_12767,N_13295);
nand U16243 (N_16243,N_14772,N_12842);
nor U16244 (N_16244,N_15107,N_14641);
nor U16245 (N_16245,N_13031,N_14878);
and U16246 (N_16246,N_15137,N_14564);
nor U16247 (N_16247,N_13182,N_12877);
nand U16248 (N_16248,N_13275,N_14434);
and U16249 (N_16249,N_13703,N_12563);
or U16250 (N_16250,N_15332,N_14565);
nand U16251 (N_16251,N_15063,N_13811);
xnor U16252 (N_16252,N_14711,N_13842);
nand U16253 (N_16253,N_13206,N_14718);
nand U16254 (N_16254,N_15030,N_13468);
xnor U16255 (N_16255,N_13640,N_14880);
nor U16256 (N_16256,N_13546,N_14307);
and U16257 (N_16257,N_12621,N_15059);
nor U16258 (N_16258,N_12746,N_13197);
or U16259 (N_16259,N_15284,N_13186);
nand U16260 (N_16260,N_14991,N_15250);
nor U16261 (N_16261,N_15468,N_13326);
or U16262 (N_16262,N_12584,N_13190);
and U16263 (N_16263,N_15591,N_14353);
xnor U16264 (N_16264,N_13930,N_12702);
or U16265 (N_16265,N_12759,N_13700);
and U16266 (N_16266,N_14450,N_13832);
xor U16267 (N_16267,N_13655,N_14577);
nor U16268 (N_16268,N_13798,N_13233);
and U16269 (N_16269,N_13938,N_13974);
and U16270 (N_16270,N_13670,N_13765);
or U16271 (N_16271,N_15282,N_14405);
nand U16272 (N_16272,N_15266,N_13143);
and U16273 (N_16273,N_14930,N_14083);
nor U16274 (N_16274,N_13625,N_12619);
and U16275 (N_16275,N_14678,N_12613);
or U16276 (N_16276,N_14531,N_12967);
or U16277 (N_16277,N_12998,N_15551);
nor U16278 (N_16278,N_12546,N_14038);
or U16279 (N_16279,N_14394,N_13752);
or U16280 (N_16280,N_12871,N_12890);
and U16281 (N_16281,N_14525,N_12602);
nor U16282 (N_16282,N_14423,N_15052);
and U16283 (N_16283,N_14553,N_13192);
nor U16284 (N_16284,N_14195,N_13985);
or U16285 (N_16285,N_13833,N_13154);
nand U16286 (N_16286,N_12736,N_15622);
or U16287 (N_16287,N_15095,N_14151);
nor U16288 (N_16288,N_14201,N_13433);
xnor U16289 (N_16289,N_15275,N_15580);
and U16290 (N_16290,N_14126,N_13804);
nor U16291 (N_16291,N_14908,N_13697);
nand U16292 (N_16292,N_14893,N_14754);
or U16293 (N_16293,N_15548,N_15317);
nor U16294 (N_16294,N_13387,N_14359);
xnor U16295 (N_16295,N_15313,N_13092);
and U16296 (N_16296,N_15557,N_13244);
xor U16297 (N_16297,N_15461,N_13319);
or U16298 (N_16298,N_14098,N_15430);
nand U16299 (N_16299,N_12882,N_12745);
nor U16300 (N_16300,N_14493,N_14030);
nor U16301 (N_16301,N_13349,N_14868);
nand U16302 (N_16302,N_13875,N_14964);
or U16303 (N_16303,N_14203,N_12923);
and U16304 (N_16304,N_12900,N_14975);
nor U16305 (N_16305,N_12859,N_13934);
or U16306 (N_16306,N_13644,N_13954);
nor U16307 (N_16307,N_12784,N_15490);
or U16308 (N_16308,N_13598,N_12574);
xor U16309 (N_16309,N_13252,N_15337);
and U16310 (N_16310,N_13148,N_13900);
nand U16311 (N_16311,N_15422,N_15517);
or U16312 (N_16312,N_13979,N_13096);
or U16313 (N_16313,N_14902,N_14532);
nand U16314 (N_16314,N_14826,N_12768);
nand U16315 (N_16315,N_15006,N_12793);
nand U16316 (N_16316,N_14389,N_14161);
and U16317 (N_16317,N_13895,N_13129);
xor U16318 (N_16318,N_15576,N_15594);
or U16319 (N_16319,N_13502,N_14887);
nand U16320 (N_16320,N_12677,N_13588);
and U16321 (N_16321,N_15297,N_14632);
nand U16322 (N_16322,N_13290,N_14165);
and U16323 (N_16323,N_13270,N_12774);
xnor U16324 (N_16324,N_13971,N_15235);
nor U16325 (N_16325,N_15065,N_12849);
and U16326 (N_16326,N_14479,N_14764);
nand U16327 (N_16327,N_15247,N_13706);
and U16328 (N_16328,N_13610,N_15168);
nand U16329 (N_16329,N_14603,N_13770);
and U16330 (N_16330,N_15342,N_13576);
xor U16331 (N_16331,N_14925,N_12931);
or U16332 (N_16332,N_13157,N_15384);
nor U16333 (N_16333,N_13487,N_14131);
nand U16334 (N_16334,N_12802,N_14346);
nor U16335 (N_16335,N_12973,N_12568);
nor U16336 (N_16336,N_13087,N_14115);
nand U16337 (N_16337,N_15147,N_14900);
nand U16338 (N_16338,N_14987,N_14439);
nor U16339 (N_16339,N_12914,N_13942);
nand U16340 (N_16340,N_13747,N_14278);
nand U16341 (N_16341,N_13805,N_13975);
xnor U16342 (N_16342,N_13567,N_14995);
nand U16343 (N_16343,N_13884,N_14004);
nor U16344 (N_16344,N_14814,N_12847);
or U16345 (N_16345,N_15396,N_14096);
or U16346 (N_16346,N_12919,N_13755);
nand U16347 (N_16347,N_12789,N_13347);
and U16348 (N_16348,N_15302,N_12567);
and U16349 (N_16349,N_13211,N_15566);
or U16350 (N_16350,N_15444,N_12552);
or U16351 (N_16351,N_13689,N_15539);
nor U16352 (N_16352,N_13940,N_14862);
or U16353 (N_16353,N_13307,N_15380);
xor U16354 (N_16354,N_15431,N_15300);
and U16355 (N_16355,N_12737,N_15122);
and U16356 (N_16356,N_13229,N_13400);
and U16357 (N_16357,N_12752,N_13821);
nand U16358 (N_16358,N_13599,N_15019);
nor U16359 (N_16359,N_14534,N_15525);
and U16360 (N_16360,N_15045,N_12644);
and U16361 (N_16361,N_12717,N_12965);
nand U16362 (N_16362,N_15119,N_14974);
and U16363 (N_16363,N_14527,N_15413);
nand U16364 (N_16364,N_15148,N_14315);
nand U16365 (N_16365,N_14644,N_14670);
nor U16366 (N_16366,N_13978,N_15484);
nand U16367 (N_16367,N_12509,N_15532);
and U16368 (N_16368,N_12594,N_13185);
or U16369 (N_16369,N_13944,N_15423);
nor U16370 (N_16370,N_13237,N_12831);
nor U16371 (N_16371,N_14029,N_13481);
xor U16372 (N_16372,N_14102,N_12929);
or U16373 (N_16373,N_14795,N_15347);
nor U16374 (N_16374,N_14609,N_14183);
nand U16375 (N_16375,N_14921,N_12728);
nand U16376 (N_16376,N_12561,N_14715);
and U16377 (N_16377,N_14347,N_15062);
nor U16378 (N_16378,N_13902,N_15218);
xor U16379 (N_16379,N_14293,N_13329);
nor U16380 (N_16380,N_14144,N_13537);
nand U16381 (N_16381,N_13054,N_14650);
or U16382 (N_16382,N_15547,N_13141);
or U16383 (N_16383,N_14501,N_14492);
and U16384 (N_16384,N_12576,N_15462);
nor U16385 (N_16385,N_14036,N_12643);
nor U16386 (N_16386,N_13711,N_13570);
and U16387 (N_16387,N_14226,N_14713);
xor U16388 (N_16388,N_12731,N_14504);
xor U16389 (N_16389,N_14494,N_13017);
xor U16390 (N_16390,N_13251,N_14608);
and U16391 (N_16391,N_13021,N_12817);
nor U16392 (N_16392,N_14209,N_13405);
and U16393 (N_16393,N_14500,N_12544);
nor U16394 (N_16394,N_13040,N_14046);
and U16395 (N_16395,N_14158,N_14999);
nor U16396 (N_16396,N_14319,N_15025);
nand U16397 (N_16397,N_12904,N_14025);
nand U16398 (N_16398,N_13698,N_12876);
nand U16399 (N_16399,N_13562,N_15448);
or U16400 (N_16400,N_14314,N_13735);
or U16401 (N_16401,N_13908,N_14251);
nor U16402 (N_16402,N_12889,N_15364);
and U16403 (N_16403,N_15410,N_13885);
nand U16404 (N_16404,N_12697,N_12783);
and U16405 (N_16405,N_12996,N_12672);
and U16406 (N_16406,N_14129,N_13435);
nand U16407 (N_16407,N_14214,N_14451);
or U16408 (N_16408,N_14981,N_15073);
nor U16409 (N_16409,N_15369,N_12611);
or U16410 (N_16410,N_12868,N_14914);
and U16411 (N_16411,N_15522,N_14539);
xor U16412 (N_16412,N_14188,N_14923);
xor U16413 (N_16413,N_14459,N_15221);
and U16414 (N_16414,N_14800,N_12551);
xor U16415 (N_16415,N_12687,N_14381);
nor U16416 (N_16416,N_13906,N_14799);
and U16417 (N_16417,N_15258,N_12735);
and U16418 (N_16418,N_13332,N_15518);
nand U16419 (N_16419,N_14621,N_14065);
or U16420 (N_16420,N_12671,N_14717);
nand U16421 (N_16421,N_12880,N_13623);
and U16422 (N_16422,N_14304,N_13663);
nand U16423 (N_16423,N_13109,N_13277);
and U16424 (N_16424,N_15321,N_14876);
nand U16425 (N_16425,N_14751,N_12977);
nor U16426 (N_16426,N_14295,N_15150);
and U16427 (N_16427,N_12518,N_15463);
nand U16428 (N_16428,N_14469,N_12638);
and U16429 (N_16429,N_15070,N_14771);
and U16430 (N_16430,N_13340,N_13605);
and U16431 (N_16431,N_14935,N_12723);
nand U16432 (N_16432,N_13441,N_15289);
and U16433 (N_16433,N_12696,N_15399);
and U16434 (N_16434,N_13541,N_13943);
and U16435 (N_16435,N_14206,N_14159);
nand U16436 (N_16436,N_13260,N_13287);
or U16437 (N_16437,N_12555,N_15526);
and U16438 (N_16438,N_13432,N_15387);
or U16439 (N_16439,N_14997,N_13628);
and U16440 (N_16440,N_15524,N_13631);
or U16441 (N_16441,N_15353,N_12875);
nor U16442 (N_16442,N_14691,N_12910);
and U16443 (N_16443,N_14688,N_12653);
or U16444 (N_16444,N_14327,N_12809);
or U16445 (N_16445,N_12513,N_13235);
and U16446 (N_16446,N_15208,N_15473);
or U16447 (N_16447,N_14021,N_13580);
nand U16448 (N_16448,N_12941,N_14287);
or U16449 (N_16449,N_14579,N_14045);
and U16450 (N_16450,N_14803,N_13415);
nor U16451 (N_16451,N_14755,N_14558);
nor U16452 (N_16452,N_14729,N_13172);
nand U16453 (N_16453,N_13593,N_13125);
or U16454 (N_16454,N_14946,N_13795);
xor U16455 (N_16455,N_13373,N_13841);
nor U16456 (N_16456,N_13484,N_15216);
or U16457 (N_16457,N_15009,N_12803);
and U16458 (N_16458,N_14653,N_13699);
nor U16459 (N_16459,N_15520,N_14769);
or U16460 (N_16460,N_13590,N_15334);
nor U16461 (N_16461,N_14124,N_13350);
and U16462 (N_16462,N_13627,N_15204);
nand U16463 (N_16463,N_15421,N_12937);
and U16464 (N_16464,N_14351,N_13330);
or U16465 (N_16465,N_15129,N_14738);
or U16466 (N_16466,N_15351,N_13145);
or U16467 (N_16467,N_13357,N_14567);
nor U16468 (N_16468,N_14721,N_13682);
xor U16469 (N_16469,N_12668,N_15043);
nor U16470 (N_16470,N_14061,N_14248);
and U16471 (N_16471,N_13504,N_12655);
or U16472 (N_16472,N_12706,N_14361);
nor U16473 (N_16473,N_13088,N_14546);
or U16474 (N_16474,N_14273,N_13493);
and U16475 (N_16475,N_15375,N_13651);
or U16476 (N_16476,N_13077,N_14646);
nor U16477 (N_16477,N_15485,N_15457);
or U16478 (N_16478,N_12761,N_13014);
nand U16479 (N_16479,N_12685,N_13583);
or U16480 (N_16480,N_13579,N_12899);
or U16481 (N_16481,N_14402,N_12988);
and U16482 (N_16482,N_13534,N_13822);
and U16483 (N_16483,N_12995,N_14348);
nor U16484 (N_16484,N_13351,N_15281);
nand U16485 (N_16485,N_15176,N_12884);
nor U16486 (N_16486,N_13661,N_14123);
nor U16487 (N_16487,N_15506,N_14659);
nor U16488 (N_16488,N_14254,N_12690);
and U16489 (N_16489,N_12921,N_15620);
nand U16490 (N_16490,N_14216,N_13763);
and U16491 (N_16491,N_13715,N_14172);
and U16492 (N_16492,N_14953,N_12799);
xnor U16493 (N_16493,N_15608,N_15201);
nand U16494 (N_16494,N_15047,N_13222);
nand U16495 (N_16495,N_12609,N_14192);
and U16496 (N_16496,N_15544,N_12650);
xor U16497 (N_16497,N_15054,N_12947);
nand U16498 (N_16498,N_14881,N_12501);
nor U16499 (N_16499,N_15596,N_14541);
or U16500 (N_16500,N_15113,N_13160);
nor U16501 (N_16501,N_12800,N_13945);
and U16502 (N_16502,N_15583,N_12911);
nor U16503 (N_16503,N_13023,N_14491);
and U16504 (N_16504,N_14370,N_13380);
and U16505 (N_16505,N_15167,N_13730);
nand U16506 (N_16506,N_13732,N_15077);
nor U16507 (N_16507,N_12721,N_14148);
nand U16508 (N_16508,N_12860,N_13856);
and U16509 (N_16509,N_14521,N_15180);
or U16510 (N_16510,N_12654,N_13159);
and U16511 (N_16511,N_15584,N_15196);
nand U16512 (N_16512,N_14430,N_15482);
xor U16513 (N_16513,N_13643,N_13656);
or U16514 (N_16514,N_15135,N_13532);
xnor U16515 (N_16515,N_14982,N_14260);
nand U16516 (N_16516,N_12664,N_13614);
or U16517 (N_16517,N_15362,N_13073);
nand U16518 (N_16518,N_14702,N_12711);
or U16519 (N_16519,N_12634,N_12639);
and U16520 (N_16520,N_13059,N_15093);
nor U16521 (N_16521,N_13569,N_14994);
or U16522 (N_16522,N_15189,N_13807);
nand U16523 (N_16523,N_13809,N_13996);
and U16524 (N_16524,N_14967,N_14757);
or U16525 (N_16525,N_13538,N_14709);
nand U16526 (N_16526,N_15429,N_13865);
or U16527 (N_16527,N_12647,N_13064);
nand U16528 (N_16528,N_15154,N_12794);
nor U16529 (N_16529,N_13191,N_14404);
nand U16530 (N_16530,N_12907,N_14817);
nor U16531 (N_16531,N_12822,N_13524);
nor U16532 (N_16532,N_15441,N_14162);
and U16533 (N_16533,N_14476,N_12716);
nand U16534 (N_16534,N_15319,N_12636);
nor U16535 (N_16535,N_15089,N_15117);
xor U16536 (N_16536,N_14926,N_12861);
or U16537 (N_16537,N_15318,N_13980);
and U16538 (N_16538,N_14320,N_13482);
or U16539 (N_16539,N_15301,N_12992);
and U16540 (N_16540,N_13308,N_13131);
nand U16541 (N_16541,N_13511,N_13207);
nor U16542 (N_16542,N_14050,N_13808);
or U16543 (N_16543,N_12918,N_13296);
nand U16544 (N_16544,N_13216,N_15530);
and U16545 (N_16545,N_14424,N_12753);
nand U16546 (N_16546,N_15419,N_12694);
nor U16547 (N_16547,N_12580,N_14692);
nor U16548 (N_16548,N_15470,N_15241);
nor U16549 (N_16549,N_13683,N_13078);
xnor U16550 (N_16550,N_15615,N_14497);
or U16551 (N_16551,N_13676,N_15534);
nor U16552 (N_16552,N_14255,N_15368);
and U16553 (N_16553,N_13677,N_13861);
or U16554 (N_16554,N_12896,N_12747);
nor U16555 (N_16555,N_13354,N_13005);
and U16556 (N_16556,N_13913,N_14706);
and U16557 (N_16557,N_15225,N_14178);
and U16558 (N_16558,N_14208,N_14150);
nor U16559 (N_16559,N_13214,N_13826);
nor U16560 (N_16560,N_13486,N_14164);
or U16561 (N_16561,N_14235,N_15374);
nor U16562 (N_16562,N_15076,N_13335);
xor U16563 (N_16563,N_14524,N_13227);
or U16564 (N_16564,N_14601,N_14583);
nand U16565 (N_16565,N_13802,N_12500);
or U16566 (N_16566,N_15377,N_13779);
and U16567 (N_16567,N_13751,N_12797);
or U16568 (N_16568,N_13973,N_14259);
xor U16569 (N_16569,N_13907,N_12851);
nor U16570 (N_16570,N_13568,N_15209);
nand U16571 (N_16571,N_13891,N_13496);
and U16572 (N_16572,N_13110,N_15210);
and U16573 (N_16573,N_12749,N_13828);
and U16574 (N_16574,N_13390,N_14620);
nand U16575 (N_16575,N_15244,N_14720);
or U16576 (N_16576,N_12591,N_15604);
nor U16577 (N_16577,N_12724,N_13257);
or U16578 (N_16578,N_13452,N_14762);
or U16579 (N_16579,N_14326,N_13549);
nand U16580 (N_16580,N_12506,N_14024);
nand U16581 (N_16581,N_14700,N_15206);
nor U16582 (N_16582,N_12744,N_13650);
nor U16583 (N_16583,N_15349,N_15492);
and U16584 (N_16584,N_13581,N_13391);
or U16585 (N_16585,N_14775,N_14191);
nand U16586 (N_16586,N_14760,N_14604);
and U16587 (N_16587,N_12645,N_12934);
and U16588 (N_16588,N_14090,N_13684);
or U16589 (N_16589,N_13965,N_14019);
or U16590 (N_16590,N_13778,N_13113);
nor U16591 (N_16591,N_15346,N_12893);
and U16592 (N_16592,N_13782,N_14554);
and U16593 (N_16593,N_14860,N_13678);
xor U16594 (N_16594,N_15359,N_13820);
nor U16595 (N_16595,N_15553,N_13291);
nor U16596 (N_16596,N_15069,N_12573);
and U16597 (N_16597,N_14393,N_14562);
nor U16598 (N_16598,N_14545,N_13403);
and U16599 (N_16599,N_13657,N_13815);
and U16600 (N_16600,N_13507,N_13167);
or U16601 (N_16601,N_14683,N_12814);
nor U16602 (N_16602,N_14667,N_13239);
nor U16603 (N_16603,N_13245,N_15305);
nor U16604 (N_16604,N_14514,N_15181);
or U16605 (N_16605,N_14699,N_15479);
or U16606 (N_16606,N_14551,N_14284);
and U16607 (N_16607,N_13806,N_15023);
or U16608 (N_16608,N_15015,N_13467);
or U16609 (N_16609,N_13777,N_14397);
nand U16610 (N_16610,N_12556,N_13279);
nand U16611 (N_16611,N_13787,N_13339);
or U16612 (N_16612,N_13221,N_12632);
nand U16613 (N_16613,N_15061,N_12772);
and U16614 (N_16614,N_15260,N_13512);
or U16615 (N_16615,N_13535,N_14399);
and U16616 (N_16616,N_13840,N_15315);
nor U16617 (N_16617,N_14031,N_13076);
nor U16618 (N_16618,N_12902,N_13328);
or U16619 (N_16619,N_14763,N_13864);
xor U16620 (N_16620,N_14854,N_13264);
nor U16621 (N_16621,N_14049,N_13967);
nand U16622 (N_16622,N_14827,N_13436);
or U16623 (N_16623,N_15237,N_14809);
nand U16624 (N_16624,N_12966,N_15173);
nand U16625 (N_16625,N_13375,N_14170);
nor U16626 (N_16626,N_15621,N_15570);
and U16627 (N_16627,N_13195,N_13311);
nand U16628 (N_16628,N_13702,N_15529);
nor U16629 (N_16629,N_13693,N_13890);
or U16630 (N_16630,N_15603,N_13213);
or U16631 (N_16631,N_14471,N_13857);
or U16632 (N_16632,N_14222,N_13757);
nor U16633 (N_16633,N_15124,N_15100);
or U16634 (N_16634,N_13104,N_12942);
or U16635 (N_16635,N_14042,N_15582);
or U16636 (N_16636,N_13853,N_15242);
nor U16637 (N_16637,N_14433,N_12865);
nand U16638 (N_16638,N_13033,N_15531);
and U16639 (N_16639,N_13164,N_13048);
and U16640 (N_16640,N_13695,N_14227);
xnor U16641 (N_16641,N_14333,N_13072);
nand U16642 (N_16642,N_15038,N_12523);
nor U16643 (N_16643,N_15164,N_14849);
nor U16644 (N_16644,N_14230,N_14294);
or U16645 (N_16645,N_13862,N_12869);
nand U16646 (N_16646,N_13790,N_13696);
nor U16647 (N_16647,N_15145,N_13740);
xor U16648 (N_16648,N_13001,N_13679);
and U16649 (N_16649,N_13672,N_14645);
nor U16650 (N_16650,N_13714,N_14240);
or U16651 (N_16651,N_13414,N_13392);
nand U16652 (N_16652,N_12575,N_14573);
or U16653 (N_16653,N_13272,N_15071);
or U16654 (N_16654,N_14833,N_13701);
nor U16655 (N_16655,N_14008,N_14070);
nand U16656 (N_16656,N_12531,N_13479);
or U16657 (N_16657,N_13912,N_12560);
and U16658 (N_16658,N_12881,N_13594);
nor U16659 (N_16659,N_14530,N_13989);
xor U16660 (N_16660,N_14818,N_14106);
nor U16661 (N_16661,N_15187,N_14241);
xor U16662 (N_16662,N_15358,N_14077);
and U16663 (N_16663,N_14075,N_15207);
and U16664 (N_16664,N_14842,N_13704);
xor U16665 (N_16665,N_14107,N_15165);
nand U16666 (N_16666,N_15328,N_13412);
nand U16667 (N_16667,N_13365,N_15574);
nand U16668 (N_16668,N_15614,N_14363);
xnor U16669 (N_16669,N_12858,N_15383);
nor U16670 (N_16670,N_13263,N_15415);
or U16671 (N_16671,N_14349,N_14810);
and U16672 (N_16672,N_13927,N_13395);
nand U16673 (N_16673,N_15540,N_14830);
nand U16674 (N_16674,N_13108,N_14811);
and U16675 (N_16675,N_15495,N_13619);
and U16676 (N_16676,N_12862,N_12968);
nor U16677 (N_16677,N_13551,N_15381);
nand U16678 (N_16678,N_14937,N_13205);
nor U16679 (N_16679,N_12607,N_13654);
and U16680 (N_16680,N_14244,N_14288);
or U16681 (N_16681,N_14697,N_13669);
and U16682 (N_16682,N_14792,N_15501);
and U16683 (N_16683,N_14840,N_13209);
nor U16684 (N_16684,N_14965,N_14384);
nor U16685 (N_16685,N_15246,N_15291);
nor U16686 (N_16686,N_14622,N_12930);
nor U16687 (N_16687,N_13049,N_13869);
and U16688 (N_16688,N_14635,N_14611);
nor U16689 (N_16689,N_13116,N_13769);
or U16690 (N_16690,N_12989,N_14290);
nor U16691 (N_16691,N_14039,N_14040);
or U16692 (N_16692,N_13034,N_14574);
nand U16693 (N_16693,N_14379,N_13255);
xor U16694 (N_16694,N_13388,N_13492);
or U16695 (N_16695,N_13745,N_14801);
or U16696 (N_16696,N_14983,N_13090);
nand U16697 (N_16697,N_14634,N_14001);
and U16698 (N_16698,N_12720,N_13503);
nand U16699 (N_16699,N_14582,N_13775);
nor U16700 (N_16700,N_13564,N_15585);
or U16701 (N_16701,N_13491,N_12791);
or U16702 (N_16702,N_13829,N_12593);
and U16703 (N_16703,N_14352,N_13813);
nand U16704 (N_16704,N_15271,N_15311);
nand U16705 (N_16705,N_14576,N_14054);
nand U16706 (N_16706,N_14617,N_13916);
nor U16707 (N_16707,N_14415,N_13158);
xnor U16708 (N_16708,N_14242,N_12659);
nand U16709 (N_16709,N_14296,N_12922);
and U16710 (N_16710,N_14690,N_15606);
nand U16711 (N_16711,N_15549,N_13066);
xnor U16712 (N_16712,N_13022,N_14145);
nand U16713 (N_16713,N_13367,N_14280);
nand U16714 (N_16714,N_14356,N_12532);
nand U16715 (N_16715,N_14505,N_14815);
or U16716 (N_16716,N_13577,N_12935);
nor U16717 (N_16717,N_13995,N_12709);
xnor U16718 (N_16718,N_14535,N_13618);
and U16719 (N_16719,N_14139,N_14929);
and U16720 (N_16720,N_13872,N_13844);
nand U16721 (N_16721,N_14560,N_13098);
or U16722 (N_16722,N_15205,N_14838);
nor U16723 (N_16723,N_15263,N_13500);
nor U16724 (N_16724,N_14737,N_13442);
and U16725 (N_16725,N_14731,N_14872);
and U16726 (N_16726,N_14247,N_13242);
xnor U16727 (N_16727,N_13615,N_14398);
or U16728 (N_16728,N_15458,N_14538);
and U16729 (N_16729,N_12559,N_12938);
nor U16730 (N_16730,N_12951,N_12693);
nand U16731 (N_16731,N_14869,N_13720);
and U16732 (N_16732,N_13722,N_14134);
nor U16733 (N_16733,N_14167,N_14966);
and U16734 (N_16734,N_14649,N_12739);
and U16735 (N_16735,N_14258,N_13859);
nand U16736 (N_16736,N_12971,N_12819);
nand U16737 (N_16737,N_14122,N_15590);
nand U16738 (N_16738,N_14891,N_13302);
nand U16739 (N_16739,N_12957,N_13029);
and U16740 (N_16740,N_14472,N_13183);
nor U16741 (N_16741,N_14057,N_13603);
nor U16742 (N_16742,N_13079,N_13894);
nand U16743 (N_16743,N_12708,N_13773);
nand U16744 (N_16744,N_14457,N_14972);
or U16745 (N_16745,N_14056,N_13082);
nor U16746 (N_16746,N_13304,N_14543);
nand U16747 (N_16747,N_14074,N_14041);
nand U16748 (N_16748,N_12540,N_15354);
xnor U16749 (N_16749,N_14674,N_15562);
nor U16750 (N_16750,N_13796,N_12597);
nor U16751 (N_16751,N_12529,N_15252);
xor U16752 (N_16752,N_15445,N_13960);
and U16753 (N_16753,N_14082,N_12583);
or U16754 (N_16754,N_12776,N_15600);
or U16755 (N_16755,N_15555,N_12864);
nor U16756 (N_16756,N_13331,N_15478);
nand U16757 (N_16757,N_14207,N_14696);
nor U16758 (N_16758,N_13674,N_15064);
and U16759 (N_16759,N_15303,N_13776);
or U16760 (N_16760,N_14643,N_15366);
xnor U16761 (N_16761,N_14656,N_12683);
or U16762 (N_16762,N_12997,N_14572);
nor U16763 (N_16763,N_14652,N_12811);
and U16764 (N_16764,N_13882,N_12714);
nor U16765 (N_16765,N_14335,N_15467);
nand U16766 (N_16766,N_13881,N_13592);
nand U16767 (N_16767,N_13220,N_15592);
nand U16768 (N_16768,N_13135,N_14783);
nor U16769 (N_16769,N_13584,N_13218);
nand U16770 (N_16770,N_15096,N_14647);
and U16771 (N_16771,N_13606,N_14984);
or U16772 (N_16772,N_13498,N_15361);
nand U16773 (N_16773,N_15320,N_14979);
and U16774 (N_16774,N_14625,N_13767);
or U16775 (N_16775,N_14473,N_13418);
xor U16776 (N_16776,N_14210,N_12754);
xnor U16777 (N_16777,N_15491,N_12541);
or U16778 (N_16778,N_14672,N_15329);
and U16779 (N_16779,N_13708,N_13612);
nand U16780 (N_16780,N_15116,N_14187);
or U16781 (N_16781,N_13725,N_13382);
and U16782 (N_16782,N_14023,N_15042);
nand U16783 (N_16783,N_12620,N_13016);
or U16784 (N_16784,N_14839,N_12612);
nor U16785 (N_16785,N_13411,N_13958);
or U16786 (N_16786,N_13756,N_14358);
or U16787 (N_16787,N_14664,N_14014);
nand U16788 (N_16788,N_15010,N_13301);
or U16789 (N_16789,N_13736,N_14245);
nor U16790 (N_16790,N_13759,N_15132);
or U16791 (N_16791,N_14686,N_14486);
and U16792 (N_16792,N_15408,N_14507);
nor U16793 (N_16793,N_15586,N_12948);
nand U16794 (N_16794,N_14512,N_14403);
xnor U16795 (N_16795,N_15004,N_15056);
nand U16796 (N_16796,N_13613,N_12630);
nand U16797 (N_16797,N_14968,N_12796);
and U16798 (N_16798,N_13341,N_14673);
nor U16799 (N_16799,N_13983,N_13666);
xor U16800 (N_16800,N_12891,N_14047);
xnor U16801 (N_16801,N_14606,N_14275);
and U16802 (N_16802,N_13134,N_14753);
or U16803 (N_16803,N_14515,N_12666);
and U16804 (N_16804,N_15403,N_13282);
nor U16805 (N_16805,N_15340,N_14960);
and U16806 (N_16806,N_14774,N_12963);
xnor U16807 (N_16807,N_12764,N_12946);
nand U16808 (N_16808,N_12763,N_14340);
nand U16809 (N_16809,N_14781,N_14642);
and U16810 (N_16810,N_14916,N_15372);
xnor U16811 (N_16811,N_15464,N_12663);
nor U16812 (N_16812,N_15178,N_14436);
or U16813 (N_16813,N_12673,N_12548);
nor U16814 (N_16814,N_12825,N_13920);
nor U16815 (N_16815,N_12550,N_15033);
nand U16816 (N_16816,N_15442,N_14062);
or U16817 (N_16817,N_13719,N_13231);
nor U16818 (N_16818,N_14382,N_12622);
and U16819 (N_16819,N_14626,N_14939);
nor U16820 (N_16820,N_13236,N_12927);
and U16821 (N_16821,N_13993,N_12808);
nor U16822 (N_16822,N_12821,N_14204);
or U16823 (N_16823,N_14719,N_14528);
xor U16824 (N_16824,N_15053,N_12732);
and U16825 (N_16825,N_15109,N_14253);
nor U16826 (N_16826,N_14441,N_13565);
nor U16827 (N_16827,N_14773,N_13948);
nor U16828 (N_16828,N_14899,N_14020);
and U16829 (N_16829,N_13903,N_15577);
and U16830 (N_16830,N_12589,N_13766);
nand U16831 (N_16831,N_13128,N_15108);
and U16832 (N_16832,N_13515,N_13685);
nand U16833 (N_16833,N_13928,N_14675);
or U16834 (N_16834,N_13440,N_13315);
or U16835 (N_16835,N_15515,N_13559);
or U16836 (N_16836,N_13083,N_12534);
nand U16837 (N_16837,N_13041,N_15500);
nand U16838 (N_16838,N_14977,N_12729);
nor U16839 (N_16839,N_13075,N_15489);
nand U16840 (N_16840,N_13774,N_15013);
nor U16841 (N_16841,N_12656,N_13667);
and U16842 (N_16842,N_13171,N_13990);
nand U16843 (N_16843,N_14637,N_13986);
or U16844 (N_16844,N_12756,N_13199);
or U16845 (N_16845,N_14087,N_14059);
nand U16846 (N_16846,N_15575,N_13020);
nand U16847 (N_16847,N_15550,N_14677);
and U16848 (N_16848,N_13556,N_14406);
nand U16849 (N_16849,N_13446,N_15273);
and U16850 (N_16850,N_13070,N_12581);
and U16851 (N_16851,N_12553,N_13284);
nor U16852 (N_16852,N_14390,N_14482);
or U16853 (N_16853,N_14856,N_13794);
or U16854 (N_16854,N_15538,N_15140);
nand U16855 (N_16855,N_14425,N_14418);
nand U16856 (N_16856,N_14756,N_14012);
and U16857 (N_16857,N_12733,N_13984);
nor U16858 (N_16858,N_14220,N_14289);
or U16859 (N_16859,N_15198,N_13645);
xor U16860 (N_16860,N_15060,N_14076);
nand U16861 (N_16861,N_13306,N_14592);
nand U16862 (N_16862,N_14490,N_15494);
xor U16863 (N_16863,N_13074,N_13170);
nand U16864 (N_16864,N_14496,N_13554);
xnor U16865 (N_16865,N_15533,N_13035);
nor U16866 (N_16866,N_13458,N_15163);
and U16867 (N_16867,N_13548,N_12987);
xnor U16868 (N_16868,N_13622,N_13002);
or U16869 (N_16869,N_13817,N_15099);
nor U16870 (N_16870,N_13464,N_13742);
nand U16871 (N_16871,N_13258,N_13981);
and U16872 (N_16872,N_14412,N_13552);
xnor U16873 (N_16873,N_15595,N_13675);
nand U16874 (N_16874,N_12844,N_13321);
xor U16875 (N_16875,N_12624,N_14682);
and U16876 (N_16876,N_15136,N_13970);
or U16877 (N_16877,N_14750,N_13880);
nor U16878 (N_16878,N_15454,N_12955);
nor U16879 (N_16879,N_13483,N_14033);
nand U16880 (N_16880,N_14374,N_15240);
or U16881 (N_16881,N_12815,N_14154);
or U16882 (N_16882,N_14097,N_14863);
and U16883 (N_16883,N_12684,N_14633);
nor U16884 (N_16884,N_14522,N_13626);
or U16885 (N_16885,N_13372,N_12742);
nand U16886 (N_16886,N_14892,N_14407);
or U16887 (N_16887,N_13953,N_12562);
nor U16888 (N_16888,N_13226,N_14950);
nor U16889 (N_16889,N_15356,N_13635);
nand U16890 (N_16890,N_13089,N_13053);
and U16891 (N_16891,N_13792,N_14752);
nand U16892 (N_16892,N_13629,N_13897);
nor U16893 (N_16893,N_13217,N_13353);
or U16894 (N_16894,N_13430,N_15560);
or U16895 (N_16895,N_12628,N_13825);
nor U16896 (N_16896,N_13741,N_12700);
and U16897 (N_16897,N_12970,N_15519);
or U16898 (N_16898,N_12982,N_12835);
nor U16899 (N_16899,N_14128,N_12863);
nand U16900 (N_16900,N_13585,N_13454);
nor U16901 (N_16901,N_14859,N_13453);
and U16902 (N_16902,N_14612,N_15232);
and U16903 (N_16903,N_15388,N_14993);
and U16904 (N_16904,N_12635,N_13591);
or U16905 (N_16905,N_14360,N_13473);
nand U16906 (N_16906,N_12623,N_13743);
nand U16907 (N_16907,N_12894,N_13099);
and U16908 (N_16908,N_15097,N_13004);
and U16909 (N_16909,N_13434,N_13910);
nor U16910 (N_16910,N_15157,N_15382);
or U16911 (N_16911,N_12726,N_15261);
nand U16912 (N_16912,N_14010,N_13545);
or U16913 (N_16913,N_14285,N_14016);
or U16914 (N_16914,N_13589,N_13607);
nor U16915 (N_16915,N_14028,N_14132);
xor U16916 (N_16916,N_13051,N_14146);
nor U16917 (N_16917,N_13835,N_12586);
nand U16918 (N_16918,N_15286,N_13616);
or U16919 (N_16919,N_12514,N_14610);
or U16920 (N_16920,N_14959,N_12688);
and U16921 (N_16921,N_14142,N_12972);
nand U16922 (N_16922,N_13165,N_15115);
or U16923 (N_16923,N_15602,N_13744);
nor U16924 (N_16924,N_12579,N_12915);
or U16925 (N_16925,N_14873,N_13992);
and U16926 (N_16926,N_14176,N_13313);
nor U16927 (N_16927,N_14174,N_12912);
nand U16928 (N_16928,N_14270,N_13836);
or U16929 (N_16929,N_15293,N_13783);
nand U16930 (N_16930,N_13133,N_12959);
nand U16931 (N_16931,N_14689,N_13718);
and U16932 (N_16932,N_15474,N_12618);
and U16933 (N_16933,N_14133,N_13389);
xor U16934 (N_16934,N_14182,N_14438);
nor U16935 (N_16935,N_15476,N_14537);
or U16936 (N_16936,N_13374,N_13573);
and U16937 (N_16937,N_13707,N_13879);
and U16938 (N_16938,N_14343,N_14890);
or U16939 (N_16939,N_12554,N_12956);
and U16940 (N_16940,N_15159,N_14354);
or U16941 (N_16941,N_13234,N_12577);
and U16942 (N_16942,N_12770,N_13043);
and U16943 (N_16943,N_15558,N_13149);
and U16944 (N_16944,N_13602,N_12662);
and U16945 (N_16945,N_13749,N_13348);
nor U16946 (N_16946,N_14578,N_15193);
and U16947 (N_16947,N_12874,N_12626);
nand U16948 (N_16948,N_13976,N_13000);
nor U16949 (N_16949,N_13203,N_14962);
and U16950 (N_16950,N_15133,N_13025);
and U16951 (N_16951,N_14002,N_13178);
and U16952 (N_16952,N_14388,N_13662);
nor U16953 (N_16953,N_12901,N_12926);
nand U16954 (N_16954,N_13267,N_12879);
xnor U16955 (N_16955,N_15589,N_12886);
xor U16956 (N_16956,N_13637,N_12830);
and U16957 (N_16957,N_13293,N_15037);
and U16958 (N_16958,N_14716,N_15573);
xnor U16959 (N_16959,N_14114,N_13384);
xnor U16960 (N_16960,N_15276,N_14445);
nor U16961 (N_16961,N_13346,N_12528);
or U16962 (N_16962,N_15546,N_12588);
nand U16963 (N_16963,N_15106,N_15152);
nor U16964 (N_16964,N_12792,N_12945);
and U16965 (N_16965,N_12953,N_15486);
nand U16966 (N_16966,N_15156,N_12837);
xor U16967 (N_16967,N_13463,N_14851);
nor U16968 (N_16968,N_14727,N_12962);
or U16969 (N_16969,N_14011,N_12805);
or U16970 (N_16970,N_13997,N_13363);
nand U16971 (N_16971,N_13533,N_14575);
nor U16972 (N_16972,N_14569,N_13393);
nand U16973 (N_16973,N_14003,N_12878);
nand U16974 (N_16974,N_13508,N_14080);
nor U16975 (N_16975,N_14798,N_13093);
or U16976 (N_16976,N_15598,N_13951);
or U16977 (N_16977,N_12566,N_12762);
or U16978 (N_16978,N_15452,N_13407);
nand U16979 (N_16979,N_14951,N_14614);
nor U16980 (N_16980,N_15466,N_15012);
and U16981 (N_16981,N_14998,N_13923);
nor U16982 (N_16982,N_12790,N_13596);
or U16983 (N_16983,N_14442,N_13105);
or U16984 (N_16984,N_15141,N_12543);
or U16985 (N_16985,N_15153,N_13325);
or U16986 (N_16986,N_15066,N_13309);
nor U16987 (N_16987,N_15192,N_13312);
or U16988 (N_16988,N_14229,N_13286);
nand U16989 (N_16989,N_13187,N_14416);
and U16990 (N_16990,N_12661,N_15453);
nor U16991 (N_16991,N_12658,N_15306);
nor U16992 (N_16992,N_14414,N_15029);
nor U16993 (N_16993,N_13915,N_13630);
nor U16994 (N_16994,N_13544,N_15393);
nor U16995 (N_16995,N_15255,N_15268);
nor U16996 (N_16996,N_14623,N_14232);
and U16997 (N_16997,N_13184,N_15571);
nor U16998 (N_16998,N_14671,N_13281);
nand U16999 (N_16999,N_14184,N_13566);
xnor U17000 (N_17000,N_12699,N_13558);
and U17001 (N_17001,N_13424,N_13225);
and U17002 (N_17002,N_13998,N_15111);
or U17003 (N_17003,N_13705,N_14190);
nand U17004 (N_17004,N_12748,N_13918);
nand U17005 (N_17005,N_14788,N_15352);
nand U17006 (N_17006,N_12833,N_13052);
nor U17007 (N_17007,N_14378,N_13721);
nor U17008 (N_17008,N_12603,N_13761);
and U17009 (N_17009,N_13506,N_15451);
or U17010 (N_17010,N_13547,N_12760);
nand U17011 (N_17011,N_14444,N_14282);
or U17012 (N_17012,N_12932,N_12950);
or U17013 (N_17013,N_13933,N_15092);
and U17014 (N_17014,N_13937,N_14943);
nand U17015 (N_17015,N_14092,N_13201);
nand U17016 (N_17016,N_14600,N_14835);
nand U17017 (N_17017,N_13665,N_15613);
nor U17018 (N_17018,N_13494,N_14730);
or U17019 (N_17019,N_14992,N_15272);
nand U17020 (N_17020,N_15335,N_13101);
nand U17021 (N_17021,N_14732,N_15348);
nor U17022 (N_17022,N_15587,N_14845);
or U17023 (N_17023,N_13855,N_12903);
nand U17024 (N_17024,N_13632,N_14638);
nand U17025 (N_17025,N_15552,N_13883);
nor U17026 (N_17026,N_14422,N_14196);
nor U17027 (N_17027,N_14328,N_15475);
nor U17028 (N_17028,N_14193,N_15401);
xnor U17029 (N_17029,N_12933,N_13653);
xor U17030 (N_17030,N_15203,N_14009);
and U17031 (N_17031,N_12853,N_14722);
and U17032 (N_17032,N_12892,N_15139);
xnor U17033 (N_17033,N_13553,N_13791);
and U17034 (N_17034,N_13919,N_15507);
nor U17035 (N_17035,N_14615,N_12522);
xnor U17036 (N_17036,N_13008,N_13764);
nand U17037 (N_17037,N_15040,N_12867);
xor U17038 (N_17038,N_13161,N_13084);
nor U17039 (N_17039,N_12615,N_14236);
nor U17040 (N_17040,N_15409,N_12991);
or U17041 (N_17041,N_15581,N_13018);
nand U17042 (N_17042,N_13121,N_13690);
or U17043 (N_17043,N_14341,N_15455);
xnor U17044 (N_17044,N_14385,N_13474);
or U17045 (N_17045,N_15345,N_15195);
nor U17046 (N_17046,N_15231,N_12530);
nand U17047 (N_17047,N_13428,N_13253);
and U17048 (N_17048,N_14895,N_14980);
nor U17049 (N_17049,N_14130,N_15449);
or U17050 (N_17050,N_15003,N_12917);
nor U17051 (N_17051,N_13449,N_14613);
or U17052 (N_17052,N_12908,N_15290);
xor U17053 (N_17053,N_13470,N_12508);
xor U17054 (N_17054,N_15472,N_12985);
nor U17055 (N_17055,N_13712,N_15202);
nand U17056 (N_17056,N_13600,N_14823);
nor U17057 (N_17057,N_15011,N_15098);
and U17058 (N_17058,N_15565,N_12598);
nor U17059 (N_17059,N_15617,N_14825);
xnor U17060 (N_17060,N_14927,N_14421);
nor U17061 (N_17061,N_13478,N_13038);
nor U17062 (N_17062,N_15307,N_12826);
xor U17063 (N_17063,N_13358,N_12925);
nor U17064 (N_17064,N_13539,N_15499);
nand U17065 (N_17065,N_15085,N_14446);
or U17066 (N_17066,N_12804,N_12680);
nand U17067 (N_17067,N_12705,N_15169);
nand U17068 (N_17068,N_15288,N_13758);
or U17069 (N_17069,N_14934,N_13344);
and U17070 (N_17070,N_14197,N_15618);
or U17071 (N_17071,N_12606,N_15277);
xnor U17072 (N_17072,N_14411,N_13597);
nand U17073 (N_17073,N_14454,N_13893);
nor U17074 (N_17074,N_13179,N_13322);
or U17075 (N_17075,N_14265,N_12990);
or U17076 (N_17076,N_14911,N_13376);
xor U17077 (N_17077,N_14648,N_15325);
and U17078 (N_17078,N_14072,N_15386);
nor U17079 (N_17079,N_13824,N_14676);
nor U17080 (N_17080,N_13334,N_12810);
xnor U17081 (N_17081,N_13439,N_14882);
and U17082 (N_17082,N_15072,N_13283);
or U17083 (N_17083,N_12676,N_13988);
and U17084 (N_17084,N_12691,N_15420);
or U17085 (N_17085,N_15217,N_12820);
nand U17086 (N_17086,N_15144,N_13604);
nand U17087 (N_17087,N_14155,N_13827);
and U17088 (N_17088,N_12976,N_13310);
nand U17089 (N_17089,N_13926,N_15114);
or U17090 (N_17090,N_15424,N_14587);
or U17091 (N_17091,N_13572,N_13982);
xnor U17092 (N_17092,N_13633,N_13176);
and U17093 (N_17093,N_13886,N_14330);
nand U17094 (N_17094,N_14796,N_14104);
and U17095 (N_17095,N_14922,N_15391);
nor U17096 (N_17096,N_14822,N_15545);
and U17097 (N_17097,N_15104,N_15440);
nand U17098 (N_17098,N_15432,N_14883);
nor U17099 (N_17099,N_13851,N_13274);
xor U17100 (N_17100,N_14120,N_14871);
nand U17101 (N_17101,N_13639,N_14858);
and U17102 (N_17102,N_14698,N_14820);
nand U17103 (N_17103,N_15308,N_14832);
nand U17104 (N_17104,N_13519,N_15094);
and U17105 (N_17105,N_14200,N_14786);
xnor U17106 (N_17106,N_13899,N_13024);
nor U17107 (N_17107,N_12616,N_14662);
xor U17108 (N_17108,N_15355,N_12964);
and U17109 (N_17109,N_14549,N_15078);
and U17110 (N_17110,N_14396,N_15469);
nand U17111 (N_17111,N_14463,N_12599);
or U17112 (N_17112,N_14181,N_15213);
and U17113 (N_17113,N_14271,N_15179);
nand U17114 (N_17114,N_12785,N_15279);
nor U17115 (N_17115,N_14766,N_14313);
or U17116 (N_17116,N_14901,N_12750);
or U17117 (N_17117,N_13355,N_13646);
nor U17118 (N_17118,N_14919,N_13968);
xnor U17119 (N_17119,N_14555,N_13210);
and U17120 (N_17120,N_13962,N_14595);
and U17121 (N_17121,N_13681,N_12605);
xor U17122 (N_17122,N_12657,N_12850);
nand U17123 (N_17123,N_14694,N_15439);
and U17124 (N_17124,N_14238,N_12665);
xnor U17125 (N_17125,N_15174,N_14364);
xor U17126 (N_17126,N_12827,N_15214);
nor U17127 (N_17127,N_13887,N_13409);
nand U17128 (N_17128,N_13037,N_14073);
nand U17129 (N_17129,N_14707,N_14071);
nor U17130 (N_17130,N_13729,N_14136);
nand U17131 (N_17131,N_14852,N_15226);
and U17132 (N_17132,N_12888,N_14797);
nand U17133 (N_17133,N_13095,N_14369);
and U17134 (N_17134,N_13058,N_14185);
and U17135 (N_17135,N_14044,N_13406);
and U17136 (N_17136,N_15412,N_14794);
nand U17137 (N_17137,N_12557,N_14657);
and U17138 (N_17138,N_14487,N_12958);
xnor U17139 (N_17139,N_13419,N_14940);
and U17140 (N_17140,N_13456,N_13501);
nand U17141 (N_17141,N_15233,N_13608);
nand U17142 (N_17142,N_14836,N_13280);
nand U17143 (N_17143,N_12526,N_12512);
and U17144 (N_17144,N_12640,N_13673);
or U17145 (N_17145,N_14268,N_14618);
nor U17146 (N_17146,N_14509,N_14724);
nor U17147 (N_17147,N_12504,N_12682);
nor U17148 (N_17148,N_15118,N_13273);
and U17149 (N_17149,N_12652,N_14367);
nand U17150 (N_17150,N_15611,N_15171);
or U17151 (N_17151,N_14847,N_15443);
and U17152 (N_17152,N_12600,N_14861);
nor U17153 (N_17153,N_13771,N_14510);
nor U17154 (N_17154,N_13117,N_12610);
nor U17155 (N_17155,N_14944,N_13215);
and U17156 (N_17156,N_15516,N_13563);
nand U17157 (N_17157,N_15039,N_15392);
and U17158 (N_17158,N_14640,N_13858);
and U17159 (N_17159,N_14779,N_13010);
xnor U17160 (N_17160,N_12527,N_14308);
or U17161 (N_17161,N_13230,N_13039);
nor U17162 (N_17162,N_13459,N_14086);
nand U17163 (N_17163,N_13032,N_14813);
or U17164 (N_17164,N_13080,N_13062);
xnor U17165 (N_17165,N_13445,N_12740);
nor U17166 (N_17166,N_15350,N_13797);
and U17167 (N_17167,N_14458,N_15005);
nor U17168 (N_17168,N_14125,N_14426);
or U17169 (N_17169,N_13124,N_14478);
nor U17170 (N_17170,N_13180,N_12845);
xor U17171 (N_17171,N_14636,N_13269);
and U17172 (N_17172,N_12614,N_15184);
nand U17173 (N_17173,N_14485,N_15220);
and U17174 (N_17174,N_13132,N_13898);
and U17175 (N_17175,N_14850,N_14665);
or U17176 (N_17176,N_14316,N_13949);
nor U17177 (N_17177,N_13323,N_14499);
or U17178 (N_17178,N_13518,N_13250);
nand U17179 (N_17179,N_12848,N_13561);
nor U17180 (N_17180,N_14212,N_13748);
and U17181 (N_17181,N_13060,N_14542);
nor U17182 (N_17182,N_13168,N_12718);
or U17183 (N_17183,N_13870,N_13799);
nor U17184 (N_17184,N_13298,N_15234);
nand U17185 (N_17185,N_14877,N_13359);
xor U17186 (N_17186,N_12641,N_14897);
and U17187 (N_17187,N_14710,N_13391);
or U17188 (N_17188,N_13003,N_13635);
nor U17189 (N_17189,N_15110,N_13735);
or U17190 (N_17190,N_13295,N_15544);
and U17191 (N_17191,N_15199,N_14625);
nor U17192 (N_17192,N_15214,N_14052);
or U17193 (N_17193,N_14212,N_15392);
or U17194 (N_17194,N_15005,N_13909);
nand U17195 (N_17195,N_12536,N_15606);
and U17196 (N_17196,N_15395,N_14074);
nor U17197 (N_17197,N_14562,N_15197);
or U17198 (N_17198,N_12627,N_14571);
nor U17199 (N_17199,N_14388,N_12924);
nand U17200 (N_17200,N_13368,N_12898);
and U17201 (N_17201,N_13780,N_12551);
and U17202 (N_17202,N_15219,N_13783);
or U17203 (N_17203,N_13493,N_12835);
and U17204 (N_17204,N_14603,N_13312);
or U17205 (N_17205,N_14543,N_12759);
nand U17206 (N_17206,N_13277,N_14780);
or U17207 (N_17207,N_13874,N_15543);
and U17208 (N_17208,N_15072,N_15451);
nand U17209 (N_17209,N_14238,N_14037);
or U17210 (N_17210,N_14816,N_13671);
nor U17211 (N_17211,N_14494,N_12658);
nand U17212 (N_17212,N_13220,N_13714);
nor U17213 (N_17213,N_15085,N_12588);
and U17214 (N_17214,N_13600,N_15112);
or U17215 (N_17215,N_12628,N_15273);
and U17216 (N_17216,N_12852,N_14068);
nor U17217 (N_17217,N_14797,N_13517);
nor U17218 (N_17218,N_12786,N_14056);
and U17219 (N_17219,N_15083,N_14839);
or U17220 (N_17220,N_15424,N_14714);
xor U17221 (N_17221,N_13719,N_15505);
nor U17222 (N_17222,N_14476,N_13658);
nor U17223 (N_17223,N_15169,N_13600);
xnor U17224 (N_17224,N_14858,N_12694);
nor U17225 (N_17225,N_14367,N_14305);
and U17226 (N_17226,N_14140,N_13424);
nand U17227 (N_17227,N_13895,N_14115);
nand U17228 (N_17228,N_13637,N_15192);
or U17229 (N_17229,N_13260,N_15561);
or U17230 (N_17230,N_14314,N_14820);
or U17231 (N_17231,N_13799,N_15589);
and U17232 (N_17232,N_13165,N_13783);
xnor U17233 (N_17233,N_13174,N_13061);
or U17234 (N_17234,N_14538,N_14649);
xnor U17235 (N_17235,N_13595,N_14360);
xnor U17236 (N_17236,N_14792,N_14300);
or U17237 (N_17237,N_14393,N_13037);
nor U17238 (N_17238,N_14859,N_14012);
nand U17239 (N_17239,N_13163,N_12767);
xor U17240 (N_17240,N_12982,N_12514);
or U17241 (N_17241,N_13189,N_15415);
nand U17242 (N_17242,N_13711,N_12976);
nor U17243 (N_17243,N_15438,N_15117);
nand U17244 (N_17244,N_13625,N_12573);
nor U17245 (N_17245,N_15317,N_14159);
xnor U17246 (N_17246,N_14951,N_15605);
nor U17247 (N_17247,N_12515,N_13807);
nand U17248 (N_17248,N_13443,N_14206);
or U17249 (N_17249,N_12886,N_13332);
or U17250 (N_17250,N_13437,N_14912);
or U17251 (N_17251,N_15269,N_13270);
and U17252 (N_17252,N_14089,N_14032);
nand U17253 (N_17253,N_15387,N_13386);
or U17254 (N_17254,N_15442,N_13845);
nand U17255 (N_17255,N_13152,N_14679);
or U17256 (N_17256,N_14089,N_13971);
nand U17257 (N_17257,N_13192,N_13531);
nand U17258 (N_17258,N_15339,N_14992);
or U17259 (N_17259,N_14984,N_12783);
nor U17260 (N_17260,N_13933,N_13683);
nand U17261 (N_17261,N_13860,N_15517);
nor U17262 (N_17262,N_13130,N_13662);
and U17263 (N_17263,N_15368,N_13848);
nand U17264 (N_17264,N_15018,N_15232);
and U17265 (N_17265,N_14197,N_15564);
nand U17266 (N_17266,N_14578,N_13526);
xnor U17267 (N_17267,N_14895,N_14512);
nor U17268 (N_17268,N_12681,N_12548);
and U17269 (N_17269,N_14434,N_13637);
nor U17270 (N_17270,N_14685,N_14897);
or U17271 (N_17271,N_14444,N_14834);
and U17272 (N_17272,N_15083,N_14859);
nand U17273 (N_17273,N_15097,N_13865);
nor U17274 (N_17274,N_14370,N_15045);
and U17275 (N_17275,N_13616,N_14566);
or U17276 (N_17276,N_12718,N_12519);
nand U17277 (N_17277,N_13341,N_15105);
and U17278 (N_17278,N_15343,N_14855);
or U17279 (N_17279,N_14431,N_15394);
nor U17280 (N_17280,N_15566,N_15193);
nand U17281 (N_17281,N_14109,N_14141);
or U17282 (N_17282,N_15143,N_15078);
and U17283 (N_17283,N_14663,N_13572);
nand U17284 (N_17284,N_14641,N_15180);
nand U17285 (N_17285,N_13949,N_15300);
nor U17286 (N_17286,N_13815,N_14039);
nand U17287 (N_17287,N_13561,N_14390);
nor U17288 (N_17288,N_14727,N_13380);
or U17289 (N_17289,N_12775,N_15431);
nor U17290 (N_17290,N_13776,N_15608);
nor U17291 (N_17291,N_13730,N_13653);
and U17292 (N_17292,N_13687,N_13959);
nor U17293 (N_17293,N_12824,N_12666);
or U17294 (N_17294,N_14482,N_14398);
nor U17295 (N_17295,N_13939,N_13800);
or U17296 (N_17296,N_13901,N_13212);
and U17297 (N_17297,N_15228,N_13544);
xor U17298 (N_17298,N_13368,N_15369);
xnor U17299 (N_17299,N_15371,N_13929);
and U17300 (N_17300,N_13544,N_14685);
nand U17301 (N_17301,N_13798,N_13406);
and U17302 (N_17302,N_14327,N_15162);
nand U17303 (N_17303,N_14011,N_13447);
xnor U17304 (N_17304,N_12872,N_13777);
or U17305 (N_17305,N_13630,N_14754);
nand U17306 (N_17306,N_13139,N_13466);
or U17307 (N_17307,N_14939,N_15622);
and U17308 (N_17308,N_13215,N_13634);
nand U17309 (N_17309,N_12789,N_13824);
nor U17310 (N_17310,N_13787,N_13302);
nor U17311 (N_17311,N_14806,N_13223);
or U17312 (N_17312,N_15504,N_14753);
or U17313 (N_17313,N_12515,N_13546);
xor U17314 (N_17314,N_14896,N_14166);
or U17315 (N_17315,N_13620,N_13779);
or U17316 (N_17316,N_13360,N_12893);
or U17317 (N_17317,N_12958,N_13787);
or U17318 (N_17318,N_12506,N_12771);
nand U17319 (N_17319,N_13958,N_14033);
or U17320 (N_17320,N_14202,N_14289);
or U17321 (N_17321,N_13659,N_14423);
and U17322 (N_17322,N_13575,N_14906);
or U17323 (N_17323,N_14345,N_13935);
and U17324 (N_17324,N_15317,N_14703);
and U17325 (N_17325,N_15254,N_12979);
and U17326 (N_17326,N_12815,N_14166);
nor U17327 (N_17327,N_12942,N_14666);
nor U17328 (N_17328,N_14499,N_14902);
or U17329 (N_17329,N_13592,N_14456);
or U17330 (N_17330,N_15303,N_14758);
nand U17331 (N_17331,N_14514,N_13501);
nand U17332 (N_17332,N_12524,N_14578);
nor U17333 (N_17333,N_15196,N_15295);
nor U17334 (N_17334,N_13306,N_14840);
and U17335 (N_17335,N_15177,N_13700);
nand U17336 (N_17336,N_12972,N_14050);
nand U17337 (N_17337,N_13875,N_15421);
nor U17338 (N_17338,N_12663,N_14763);
and U17339 (N_17339,N_14407,N_14383);
nor U17340 (N_17340,N_14962,N_14528);
nand U17341 (N_17341,N_12901,N_14668);
nor U17342 (N_17342,N_13083,N_13108);
nor U17343 (N_17343,N_15450,N_12827);
or U17344 (N_17344,N_15295,N_14672);
xor U17345 (N_17345,N_13667,N_14822);
or U17346 (N_17346,N_13444,N_13874);
or U17347 (N_17347,N_12997,N_15090);
and U17348 (N_17348,N_12982,N_14777);
and U17349 (N_17349,N_15154,N_13899);
and U17350 (N_17350,N_12668,N_14281);
nor U17351 (N_17351,N_14483,N_14255);
nand U17352 (N_17352,N_15078,N_13683);
and U17353 (N_17353,N_15155,N_13740);
and U17354 (N_17354,N_13257,N_13379);
nand U17355 (N_17355,N_15090,N_14315);
nor U17356 (N_17356,N_14681,N_13720);
nand U17357 (N_17357,N_13380,N_14556);
xnor U17358 (N_17358,N_15310,N_15569);
nand U17359 (N_17359,N_14368,N_14877);
and U17360 (N_17360,N_14494,N_12821);
and U17361 (N_17361,N_13485,N_14359);
nand U17362 (N_17362,N_14582,N_15338);
and U17363 (N_17363,N_15149,N_14962);
nand U17364 (N_17364,N_13941,N_13392);
and U17365 (N_17365,N_13425,N_14765);
nor U17366 (N_17366,N_14225,N_12561);
and U17367 (N_17367,N_12777,N_15600);
nor U17368 (N_17368,N_13518,N_15493);
nor U17369 (N_17369,N_12857,N_13928);
or U17370 (N_17370,N_13676,N_14300);
xor U17371 (N_17371,N_15552,N_13753);
nor U17372 (N_17372,N_13290,N_13036);
nor U17373 (N_17373,N_15196,N_13808);
nand U17374 (N_17374,N_14610,N_15138);
nand U17375 (N_17375,N_13192,N_13689);
nand U17376 (N_17376,N_13393,N_14514);
nand U17377 (N_17377,N_13348,N_15064);
nand U17378 (N_17378,N_15167,N_12547);
nand U17379 (N_17379,N_13142,N_13022);
or U17380 (N_17380,N_13300,N_13212);
nand U17381 (N_17381,N_14004,N_15074);
nand U17382 (N_17382,N_14662,N_15484);
nor U17383 (N_17383,N_14257,N_13259);
and U17384 (N_17384,N_15341,N_14624);
nor U17385 (N_17385,N_13765,N_15440);
or U17386 (N_17386,N_14193,N_13951);
xnor U17387 (N_17387,N_13594,N_14924);
and U17388 (N_17388,N_12630,N_14079);
or U17389 (N_17389,N_14938,N_12738);
nand U17390 (N_17390,N_15431,N_14462);
nand U17391 (N_17391,N_13342,N_12500);
nand U17392 (N_17392,N_13968,N_14299);
nor U17393 (N_17393,N_13535,N_14384);
xor U17394 (N_17394,N_14514,N_15016);
or U17395 (N_17395,N_15123,N_14525);
nand U17396 (N_17396,N_15114,N_14070);
nand U17397 (N_17397,N_12518,N_13781);
or U17398 (N_17398,N_15570,N_14583);
xnor U17399 (N_17399,N_14919,N_13700);
and U17400 (N_17400,N_12885,N_13830);
or U17401 (N_17401,N_13419,N_13110);
nor U17402 (N_17402,N_15561,N_14002);
or U17403 (N_17403,N_13758,N_13780);
nand U17404 (N_17404,N_14441,N_15536);
or U17405 (N_17405,N_15002,N_13279);
nand U17406 (N_17406,N_14235,N_15323);
nor U17407 (N_17407,N_12686,N_14653);
or U17408 (N_17408,N_14906,N_12764);
and U17409 (N_17409,N_15129,N_13316);
nor U17410 (N_17410,N_13493,N_15250);
nand U17411 (N_17411,N_12821,N_14362);
and U17412 (N_17412,N_13199,N_14190);
nor U17413 (N_17413,N_14698,N_15410);
or U17414 (N_17414,N_14706,N_15082);
nand U17415 (N_17415,N_14341,N_13032);
and U17416 (N_17416,N_13347,N_14438);
nand U17417 (N_17417,N_13504,N_15216);
and U17418 (N_17418,N_14589,N_14062);
or U17419 (N_17419,N_13252,N_13573);
and U17420 (N_17420,N_12939,N_14065);
nor U17421 (N_17421,N_13516,N_13902);
nand U17422 (N_17422,N_14264,N_14168);
nor U17423 (N_17423,N_13009,N_14469);
and U17424 (N_17424,N_15015,N_14734);
nor U17425 (N_17425,N_13346,N_12532);
xnor U17426 (N_17426,N_13318,N_14865);
or U17427 (N_17427,N_12732,N_15311);
xnor U17428 (N_17428,N_15523,N_14439);
or U17429 (N_17429,N_13698,N_15096);
nand U17430 (N_17430,N_14259,N_15165);
and U17431 (N_17431,N_14017,N_14063);
and U17432 (N_17432,N_12702,N_14183);
and U17433 (N_17433,N_14836,N_14113);
nor U17434 (N_17434,N_13593,N_13945);
and U17435 (N_17435,N_13760,N_15219);
nor U17436 (N_17436,N_12859,N_13162);
and U17437 (N_17437,N_14482,N_14905);
or U17438 (N_17438,N_13330,N_14276);
or U17439 (N_17439,N_13914,N_13407);
or U17440 (N_17440,N_13448,N_14048);
and U17441 (N_17441,N_12662,N_13323);
or U17442 (N_17442,N_14417,N_14036);
and U17443 (N_17443,N_15374,N_12956);
and U17444 (N_17444,N_12939,N_14969);
and U17445 (N_17445,N_13344,N_14541);
nor U17446 (N_17446,N_13038,N_15301);
and U17447 (N_17447,N_14418,N_14419);
nor U17448 (N_17448,N_13180,N_13549);
xnor U17449 (N_17449,N_14367,N_14604);
and U17450 (N_17450,N_12816,N_13812);
and U17451 (N_17451,N_15342,N_13519);
nand U17452 (N_17452,N_12978,N_14651);
and U17453 (N_17453,N_13901,N_12828);
xor U17454 (N_17454,N_13599,N_15286);
or U17455 (N_17455,N_13465,N_13662);
and U17456 (N_17456,N_13284,N_15588);
and U17457 (N_17457,N_15548,N_12510);
nor U17458 (N_17458,N_15502,N_13843);
nor U17459 (N_17459,N_14127,N_13270);
or U17460 (N_17460,N_14720,N_14234);
and U17461 (N_17461,N_14577,N_12607);
xnor U17462 (N_17462,N_13673,N_12501);
and U17463 (N_17463,N_13317,N_12589);
nor U17464 (N_17464,N_14553,N_12503);
xnor U17465 (N_17465,N_15207,N_14601);
nor U17466 (N_17466,N_15110,N_14927);
or U17467 (N_17467,N_14557,N_12817);
xor U17468 (N_17468,N_13662,N_14082);
xnor U17469 (N_17469,N_14495,N_13366);
nand U17470 (N_17470,N_14516,N_13266);
nand U17471 (N_17471,N_13028,N_14177);
nand U17472 (N_17472,N_15237,N_14270);
nand U17473 (N_17473,N_14729,N_13089);
nor U17474 (N_17474,N_13105,N_15484);
nor U17475 (N_17475,N_15523,N_15487);
or U17476 (N_17476,N_12501,N_12787);
xnor U17477 (N_17477,N_13868,N_15617);
xor U17478 (N_17478,N_12518,N_13363);
nand U17479 (N_17479,N_13555,N_12758);
xor U17480 (N_17480,N_14068,N_15149);
and U17481 (N_17481,N_13115,N_12755);
or U17482 (N_17482,N_15475,N_15556);
and U17483 (N_17483,N_15237,N_15077);
and U17484 (N_17484,N_14906,N_14037);
nand U17485 (N_17485,N_14436,N_14179);
nor U17486 (N_17486,N_14055,N_14093);
or U17487 (N_17487,N_15147,N_14397);
nor U17488 (N_17488,N_12618,N_14632);
nand U17489 (N_17489,N_12938,N_14252);
and U17490 (N_17490,N_15502,N_14033);
and U17491 (N_17491,N_13316,N_12758);
and U17492 (N_17492,N_14545,N_14379);
nand U17493 (N_17493,N_15130,N_13440);
and U17494 (N_17494,N_14170,N_12877);
nor U17495 (N_17495,N_13531,N_14150);
nand U17496 (N_17496,N_12856,N_14680);
or U17497 (N_17497,N_14201,N_15533);
and U17498 (N_17498,N_14293,N_15126);
or U17499 (N_17499,N_13548,N_13063);
or U17500 (N_17500,N_15607,N_14082);
nand U17501 (N_17501,N_15615,N_15299);
or U17502 (N_17502,N_15197,N_13249);
nor U17503 (N_17503,N_13495,N_14843);
nand U17504 (N_17504,N_15316,N_13825);
or U17505 (N_17505,N_13349,N_13383);
and U17506 (N_17506,N_14249,N_14287);
and U17507 (N_17507,N_13764,N_12897);
or U17508 (N_17508,N_12743,N_14148);
and U17509 (N_17509,N_14010,N_12720);
nor U17510 (N_17510,N_13631,N_13667);
or U17511 (N_17511,N_14802,N_14540);
xor U17512 (N_17512,N_14788,N_14573);
nand U17513 (N_17513,N_15141,N_12918);
nor U17514 (N_17514,N_12973,N_13747);
nor U17515 (N_17515,N_15433,N_13251);
or U17516 (N_17516,N_14955,N_13816);
nand U17517 (N_17517,N_13958,N_13977);
or U17518 (N_17518,N_14286,N_13015);
nor U17519 (N_17519,N_13275,N_12650);
or U17520 (N_17520,N_14989,N_13485);
or U17521 (N_17521,N_12903,N_14029);
and U17522 (N_17522,N_15233,N_14134);
or U17523 (N_17523,N_13732,N_14757);
nor U17524 (N_17524,N_12795,N_13908);
and U17525 (N_17525,N_14642,N_13684);
nand U17526 (N_17526,N_13095,N_13443);
nor U17527 (N_17527,N_14748,N_13972);
and U17528 (N_17528,N_14814,N_14056);
nor U17529 (N_17529,N_14122,N_13849);
or U17530 (N_17530,N_14705,N_14049);
or U17531 (N_17531,N_15441,N_13791);
or U17532 (N_17532,N_14159,N_14118);
nor U17533 (N_17533,N_15016,N_14458);
nand U17534 (N_17534,N_14476,N_14183);
xnor U17535 (N_17535,N_12538,N_14903);
nand U17536 (N_17536,N_15002,N_14715);
nor U17537 (N_17537,N_14238,N_12885);
xnor U17538 (N_17538,N_14142,N_14043);
and U17539 (N_17539,N_14307,N_13734);
and U17540 (N_17540,N_14229,N_13145);
nor U17541 (N_17541,N_15281,N_13605);
nand U17542 (N_17542,N_12559,N_13673);
xor U17543 (N_17543,N_15060,N_13371);
or U17544 (N_17544,N_13198,N_15296);
nand U17545 (N_17545,N_15416,N_13647);
and U17546 (N_17546,N_13713,N_13040);
nand U17547 (N_17547,N_14776,N_13322);
or U17548 (N_17548,N_13486,N_12632);
nand U17549 (N_17549,N_12670,N_15274);
and U17550 (N_17550,N_14650,N_14553);
or U17551 (N_17551,N_15406,N_12641);
nor U17552 (N_17552,N_14980,N_12645);
nor U17553 (N_17553,N_13521,N_12611);
or U17554 (N_17554,N_14966,N_13886);
or U17555 (N_17555,N_13794,N_12787);
nor U17556 (N_17556,N_15334,N_14414);
and U17557 (N_17557,N_14102,N_13402);
nor U17558 (N_17558,N_14469,N_12707);
or U17559 (N_17559,N_14510,N_13229);
xnor U17560 (N_17560,N_13993,N_14745);
nor U17561 (N_17561,N_15390,N_13298);
or U17562 (N_17562,N_13972,N_14874);
xnor U17563 (N_17563,N_12848,N_13625);
xor U17564 (N_17564,N_14851,N_14146);
and U17565 (N_17565,N_13473,N_14429);
xor U17566 (N_17566,N_14738,N_14122);
or U17567 (N_17567,N_14594,N_13936);
nor U17568 (N_17568,N_12954,N_13921);
xnor U17569 (N_17569,N_12524,N_12813);
or U17570 (N_17570,N_15475,N_13680);
or U17571 (N_17571,N_13574,N_14915);
or U17572 (N_17572,N_15349,N_13843);
nand U17573 (N_17573,N_14250,N_14203);
or U17574 (N_17574,N_14428,N_14365);
or U17575 (N_17575,N_13358,N_15116);
nand U17576 (N_17576,N_13855,N_15227);
nor U17577 (N_17577,N_14681,N_12865);
and U17578 (N_17578,N_15461,N_13246);
nand U17579 (N_17579,N_15336,N_14884);
or U17580 (N_17580,N_12840,N_13122);
or U17581 (N_17581,N_14244,N_13670);
nor U17582 (N_17582,N_13632,N_14093);
and U17583 (N_17583,N_14463,N_12533);
nand U17584 (N_17584,N_13539,N_15316);
nor U17585 (N_17585,N_14410,N_13834);
xnor U17586 (N_17586,N_12509,N_14671);
nand U17587 (N_17587,N_15478,N_13283);
and U17588 (N_17588,N_14371,N_12621);
nand U17589 (N_17589,N_13042,N_14557);
or U17590 (N_17590,N_12503,N_13325);
nand U17591 (N_17591,N_13579,N_12875);
nor U17592 (N_17592,N_15104,N_14607);
nor U17593 (N_17593,N_13885,N_13586);
or U17594 (N_17594,N_14428,N_14931);
or U17595 (N_17595,N_13591,N_15471);
xor U17596 (N_17596,N_12788,N_14590);
nand U17597 (N_17597,N_12623,N_12835);
nand U17598 (N_17598,N_14184,N_15352);
or U17599 (N_17599,N_13990,N_13616);
or U17600 (N_17600,N_13319,N_13248);
and U17601 (N_17601,N_12660,N_15007);
or U17602 (N_17602,N_14910,N_12618);
and U17603 (N_17603,N_14867,N_13906);
or U17604 (N_17604,N_13585,N_12930);
and U17605 (N_17605,N_15581,N_13431);
nand U17606 (N_17606,N_13719,N_14359);
or U17607 (N_17607,N_13087,N_13547);
nand U17608 (N_17608,N_14016,N_13178);
nor U17609 (N_17609,N_13764,N_15410);
or U17610 (N_17610,N_12837,N_15386);
and U17611 (N_17611,N_15541,N_15462);
nor U17612 (N_17612,N_15573,N_13657);
or U17613 (N_17613,N_12722,N_14944);
nor U17614 (N_17614,N_12831,N_14393);
and U17615 (N_17615,N_15224,N_14135);
and U17616 (N_17616,N_12858,N_15555);
and U17617 (N_17617,N_14356,N_14167);
and U17618 (N_17618,N_14796,N_15512);
nand U17619 (N_17619,N_12512,N_13896);
or U17620 (N_17620,N_12745,N_15490);
nand U17621 (N_17621,N_14519,N_14461);
nand U17622 (N_17622,N_13265,N_13683);
nor U17623 (N_17623,N_15414,N_15003);
or U17624 (N_17624,N_14368,N_14042);
xor U17625 (N_17625,N_14627,N_13610);
and U17626 (N_17626,N_13208,N_15457);
and U17627 (N_17627,N_14567,N_13364);
xnor U17628 (N_17628,N_14177,N_14943);
xor U17629 (N_17629,N_12748,N_12782);
and U17630 (N_17630,N_14034,N_13605);
or U17631 (N_17631,N_15113,N_14374);
nor U17632 (N_17632,N_13876,N_14473);
and U17633 (N_17633,N_14142,N_13715);
nor U17634 (N_17634,N_15265,N_12668);
xor U17635 (N_17635,N_12555,N_14507);
nand U17636 (N_17636,N_13791,N_13350);
xnor U17637 (N_17637,N_13631,N_13563);
or U17638 (N_17638,N_13576,N_13925);
xor U17639 (N_17639,N_13961,N_13238);
and U17640 (N_17640,N_13432,N_13819);
and U17641 (N_17641,N_12934,N_15369);
or U17642 (N_17642,N_15277,N_14959);
and U17643 (N_17643,N_13059,N_12597);
and U17644 (N_17644,N_12626,N_13054);
or U17645 (N_17645,N_14451,N_12755);
or U17646 (N_17646,N_14339,N_13632);
or U17647 (N_17647,N_15192,N_13585);
or U17648 (N_17648,N_15077,N_15133);
nor U17649 (N_17649,N_14335,N_13170);
nor U17650 (N_17650,N_13833,N_14484);
and U17651 (N_17651,N_12849,N_12577);
and U17652 (N_17652,N_12953,N_14189);
xor U17653 (N_17653,N_13301,N_14650);
nand U17654 (N_17654,N_15066,N_14874);
nand U17655 (N_17655,N_13092,N_14796);
nor U17656 (N_17656,N_15350,N_13685);
or U17657 (N_17657,N_13616,N_13789);
or U17658 (N_17658,N_13103,N_13612);
and U17659 (N_17659,N_14396,N_13749);
or U17660 (N_17660,N_13470,N_15321);
nand U17661 (N_17661,N_13860,N_15554);
nand U17662 (N_17662,N_12764,N_12519);
or U17663 (N_17663,N_14220,N_13045);
nand U17664 (N_17664,N_12671,N_12558);
or U17665 (N_17665,N_14419,N_14469);
nor U17666 (N_17666,N_14942,N_12501);
nor U17667 (N_17667,N_13786,N_13975);
xor U17668 (N_17668,N_14385,N_14064);
nand U17669 (N_17669,N_14764,N_14783);
and U17670 (N_17670,N_14040,N_14706);
nand U17671 (N_17671,N_12817,N_14875);
nor U17672 (N_17672,N_13794,N_13312);
nor U17673 (N_17673,N_14744,N_15252);
nand U17674 (N_17674,N_14430,N_12628);
nor U17675 (N_17675,N_15165,N_14885);
nand U17676 (N_17676,N_14095,N_13281);
nand U17677 (N_17677,N_13387,N_15175);
or U17678 (N_17678,N_15372,N_13914);
or U17679 (N_17679,N_13960,N_12552);
and U17680 (N_17680,N_15443,N_15015);
or U17681 (N_17681,N_12800,N_14535);
or U17682 (N_17682,N_13852,N_15176);
nor U17683 (N_17683,N_13093,N_15352);
nand U17684 (N_17684,N_15239,N_14784);
nor U17685 (N_17685,N_12692,N_13127);
nor U17686 (N_17686,N_14532,N_14251);
nand U17687 (N_17687,N_15465,N_15289);
nor U17688 (N_17688,N_13969,N_14149);
nand U17689 (N_17689,N_14992,N_13572);
or U17690 (N_17690,N_12685,N_13129);
or U17691 (N_17691,N_14369,N_14197);
and U17692 (N_17692,N_15029,N_13460);
xor U17693 (N_17693,N_15041,N_13348);
or U17694 (N_17694,N_14947,N_13546);
nor U17695 (N_17695,N_14004,N_15228);
xnor U17696 (N_17696,N_14180,N_13692);
nand U17697 (N_17697,N_15085,N_13094);
or U17698 (N_17698,N_14623,N_14752);
nor U17699 (N_17699,N_13004,N_12564);
nor U17700 (N_17700,N_14522,N_13649);
and U17701 (N_17701,N_15516,N_15559);
or U17702 (N_17702,N_14163,N_15251);
nand U17703 (N_17703,N_15108,N_13011);
and U17704 (N_17704,N_14664,N_12566);
nor U17705 (N_17705,N_15124,N_13487);
xor U17706 (N_17706,N_14490,N_14210);
nor U17707 (N_17707,N_15355,N_13416);
and U17708 (N_17708,N_14433,N_12968);
nor U17709 (N_17709,N_14066,N_13198);
or U17710 (N_17710,N_13432,N_15088);
and U17711 (N_17711,N_13214,N_15240);
xnor U17712 (N_17712,N_14989,N_12579);
nor U17713 (N_17713,N_14913,N_12532);
and U17714 (N_17714,N_12534,N_15479);
or U17715 (N_17715,N_14341,N_12905);
and U17716 (N_17716,N_14479,N_14878);
nor U17717 (N_17717,N_13844,N_14455);
or U17718 (N_17718,N_12680,N_15613);
or U17719 (N_17719,N_14832,N_13114);
nand U17720 (N_17720,N_13415,N_13671);
or U17721 (N_17721,N_14839,N_15129);
and U17722 (N_17722,N_13748,N_15378);
nand U17723 (N_17723,N_12895,N_13167);
nand U17724 (N_17724,N_12823,N_14585);
or U17725 (N_17725,N_13772,N_14667);
or U17726 (N_17726,N_15143,N_14427);
or U17727 (N_17727,N_12869,N_14477);
nand U17728 (N_17728,N_15422,N_15288);
or U17729 (N_17729,N_12787,N_13735);
or U17730 (N_17730,N_15125,N_12867);
and U17731 (N_17731,N_15433,N_12709);
nor U17732 (N_17732,N_12564,N_14991);
or U17733 (N_17733,N_12639,N_12713);
nand U17734 (N_17734,N_14291,N_15119);
nand U17735 (N_17735,N_13877,N_12514);
or U17736 (N_17736,N_13490,N_12577);
and U17737 (N_17737,N_13901,N_13716);
and U17738 (N_17738,N_13066,N_13314);
nand U17739 (N_17739,N_13961,N_13950);
nor U17740 (N_17740,N_14131,N_13881);
and U17741 (N_17741,N_14451,N_13177);
or U17742 (N_17742,N_13186,N_13366);
and U17743 (N_17743,N_12982,N_14049);
nand U17744 (N_17744,N_15315,N_15153);
nor U17745 (N_17745,N_15377,N_15329);
and U17746 (N_17746,N_13009,N_13545);
and U17747 (N_17747,N_15587,N_14705);
nor U17748 (N_17748,N_12648,N_14286);
nor U17749 (N_17749,N_13096,N_15190);
nand U17750 (N_17750,N_14752,N_14022);
nor U17751 (N_17751,N_13957,N_14179);
nor U17752 (N_17752,N_14784,N_14077);
nand U17753 (N_17753,N_14002,N_13614);
or U17754 (N_17754,N_15327,N_15076);
or U17755 (N_17755,N_13761,N_13640);
xor U17756 (N_17756,N_15183,N_15068);
and U17757 (N_17757,N_14429,N_13813);
or U17758 (N_17758,N_12818,N_13257);
nand U17759 (N_17759,N_13020,N_14354);
nand U17760 (N_17760,N_14607,N_15101);
and U17761 (N_17761,N_14850,N_15509);
and U17762 (N_17762,N_13175,N_12918);
xor U17763 (N_17763,N_15513,N_15424);
xnor U17764 (N_17764,N_15469,N_14651);
and U17765 (N_17765,N_12572,N_14989);
nor U17766 (N_17766,N_13707,N_15366);
or U17767 (N_17767,N_12689,N_14773);
nor U17768 (N_17768,N_12723,N_14535);
nor U17769 (N_17769,N_15244,N_13370);
nor U17770 (N_17770,N_15357,N_12792);
or U17771 (N_17771,N_13513,N_15581);
or U17772 (N_17772,N_13725,N_13359);
nor U17773 (N_17773,N_14398,N_14925);
and U17774 (N_17774,N_13813,N_13314);
nor U17775 (N_17775,N_12738,N_14247);
nand U17776 (N_17776,N_14913,N_14473);
or U17777 (N_17777,N_13685,N_14540);
nand U17778 (N_17778,N_15206,N_14437);
nor U17779 (N_17779,N_14442,N_14463);
and U17780 (N_17780,N_14484,N_14566);
nor U17781 (N_17781,N_13461,N_13644);
nor U17782 (N_17782,N_14033,N_14428);
xnor U17783 (N_17783,N_14347,N_14515);
xor U17784 (N_17784,N_13021,N_12629);
or U17785 (N_17785,N_13213,N_14631);
nand U17786 (N_17786,N_14385,N_14735);
nand U17787 (N_17787,N_14089,N_14336);
or U17788 (N_17788,N_14889,N_13861);
and U17789 (N_17789,N_12946,N_14517);
nand U17790 (N_17790,N_14929,N_15076);
nand U17791 (N_17791,N_15528,N_13768);
nand U17792 (N_17792,N_14267,N_13647);
and U17793 (N_17793,N_15489,N_15206);
nand U17794 (N_17794,N_14435,N_14471);
nand U17795 (N_17795,N_12713,N_13140);
or U17796 (N_17796,N_15065,N_15274);
xnor U17797 (N_17797,N_14480,N_13692);
and U17798 (N_17798,N_14834,N_14644);
nor U17799 (N_17799,N_12882,N_13865);
or U17800 (N_17800,N_12548,N_15235);
nand U17801 (N_17801,N_12812,N_12588);
or U17802 (N_17802,N_12962,N_14849);
nor U17803 (N_17803,N_14577,N_14868);
nand U17804 (N_17804,N_14663,N_12620);
nand U17805 (N_17805,N_13351,N_14557);
and U17806 (N_17806,N_13050,N_14239);
xnor U17807 (N_17807,N_14749,N_14283);
nand U17808 (N_17808,N_12958,N_13856);
or U17809 (N_17809,N_14173,N_14509);
xnor U17810 (N_17810,N_13518,N_13616);
or U17811 (N_17811,N_12582,N_14851);
and U17812 (N_17812,N_13424,N_13775);
nand U17813 (N_17813,N_14160,N_13157);
nor U17814 (N_17814,N_13340,N_12563);
nor U17815 (N_17815,N_13872,N_12506);
nor U17816 (N_17816,N_14925,N_14893);
or U17817 (N_17817,N_14952,N_14586);
and U17818 (N_17818,N_15196,N_15311);
or U17819 (N_17819,N_13809,N_14905);
or U17820 (N_17820,N_14854,N_12965);
nand U17821 (N_17821,N_12867,N_13621);
or U17822 (N_17822,N_15570,N_13461);
and U17823 (N_17823,N_15245,N_15135);
nand U17824 (N_17824,N_13519,N_13040);
nand U17825 (N_17825,N_14263,N_12737);
nor U17826 (N_17826,N_13669,N_13808);
xnor U17827 (N_17827,N_12833,N_14379);
and U17828 (N_17828,N_13598,N_14958);
nor U17829 (N_17829,N_14997,N_15539);
or U17830 (N_17830,N_13010,N_15598);
and U17831 (N_17831,N_15329,N_12953);
and U17832 (N_17832,N_13900,N_13377);
xnor U17833 (N_17833,N_15410,N_15622);
xnor U17834 (N_17834,N_15202,N_14273);
and U17835 (N_17835,N_13700,N_14334);
nor U17836 (N_17836,N_15552,N_13835);
xnor U17837 (N_17837,N_13012,N_14278);
xor U17838 (N_17838,N_13127,N_13934);
or U17839 (N_17839,N_14750,N_14239);
or U17840 (N_17840,N_13831,N_15093);
nor U17841 (N_17841,N_12851,N_15299);
or U17842 (N_17842,N_15104,N_14226);
or U17843 (N_17843,N_13431,N_12568);
or U17844 (N_17844,N_14011,N_13080);
or U17845 (N_17845,N_13421,N_14996);
or U17846 (N_17846,N_14011,N_12571);
or U17847 (N_17847,N_12630,N_13636);
nand U17848 (N_17848,N_12888,N_14144);
or U17849 (N_17849,N_12704,N_12557);
nor U17850 (N_17850,N_12557,N_13610);
nor U17851 (N_17851,N_13820,N_13071);
or U17852 (N_17852,N_15492,N_14213);
or U17853 (N_17853,N_13156,N_15380);
or U17854 (N_17854,N_13698,N_12989);
and U17855 (N_17855,N_15594,N_13419);
and U17856 (N_17856,N_12543,N_13892);
nor U17857 (N_17857,N_13896,N_12865);
nand U17858 (N_17858,N_14131,N_14165);
nor U17859 (N_17859,N_14097,N_12907);
xnor U17860 (N_17860,N_13653,N_12768);
and U17861 (N_17861,N_14010,N_13064);
and U17862 (N_17862,N_14950,N_14563);
nand U17863 (N_17863,N_15207,N_13147);
and U17864 (N_17864,N_14227,N_12947);
nand U17865 (N_17865,N_15584,N_15264);
nand U17866 (N_17866,N_13856,N_15512);
and U17867 (N_17867,N_13614,N_13587);
or U17868 (N_17868,N_14929,N_15337);
nand U17869 (N_17869,N_14208,N_14404);
nor U17870 (N_17870,N_12779,N_14352);
and U17871 (N_17871,N_13659,N_14297);
nand U17872 (N_17872,N_14245,N_12620);
xor U17873 (N_17873,N_13493,N_12682);
xor U17874 (N_17874,N_12860,N_14440);
nand U17875 (N_17875,N_13341,N_14452);
or U17876 (N_17876,N_15357,N_12595);
or U17877 (N_17877,N_13108,N_14300);
and U17878 (N_17878,N_15193,N_15043);
nor U17879 (N_17879,N_13884,N_12978);
nor U17880 (N_17880,N_14263,N_13312);
and U17881 (N_17881,N_12955,N_14014);
and U17882 (N_17882,N_14060,N_15422);
nand U17883 (N_17883,N_13737,N_15156);
and U17884 (N_17884,N_13710,N_12693);
or U17885 (N_17885,N_13559,N_13893);
nand U17886 (N_17886,N_13179,N_15193);
nor U17887 (N_17887,N_14118,N_15476);
or U17888 (N_17888,N_13713,N_12972);
and U17889 (N_17889,N_15487,N_14939);
nor U17890 (N_17890,N_12556,N_12635);
or U17891 (N_17891,N_13060,N_13911);
nand U17892 (N_17892,N_12896,N_14545);
nor U17893 (N_17893,N_12557,N_15131);
nand U17894 (N_17894,N_13434,N_15464);
xnor U17895 (N_17895,N_13918,N_12963);
nor U17896 (N_17896,N_14801,N_13502);
and U17897 (N_17897,N_14102,N_15148);
nor U17898 (N_17898,N_15072,N_12797);
or U17899 (N_17899,N_15298,N_13515);
and U17900 (N_17900,N_15222,N_13660);
or U17901 (N_17901,N_13356,N_12933);
nor U17902 (N_17902,N_15389,N_12751);
or U17903 (N_17903,N_14494,N_14593);
and U17904 (N_17904,N_13611,N_13169);
or U17905 (N_17905,N_12769,N_14391);
nor U17906 (N_17906,N_13108,N_14606);
or U17907 (N_17907,N_13752,N_12817);
or U17908 (N_17908,N_13651,N_15298);
and U17909 (N_17909,N_13868,N_15051);
nand U17910 (N_17910,N_12732,N_14340);
nand U17911 (N_17911,N_13731,N_15350);
or U17912 (N_17912,N_13201,N_15175);
nand U17913 (N_17913,N_15492,N_14239);
nand U17914 (N_17914,N_13379,N_12953);
and U17915 (N_17915,N_14517,N_15068);
nor U17916 (N_17916,N_14259,N_14040);
xor U17917 (N_17917,N_13544,N_14634);
or U17918 (N_17918,N_14856,N_13805);
xnor U17919 (N_17919,N_13497,N_13336);
or U17920 (N_17920,N_13331,N_13803);
nand U17921 (N_17921,N_13903,N_12776);
and U17922 (N_17922,N_12832,N_14217);
nor U17923 (N_17923,N_14407,N_14544);
or U17924 (N_17924,N_12611,N_14706);
or U17925 (N_17925,N_15441,N_12595);
xor U17926 (N_17926,N_13388,N_12508);
nor U17927 (N_17927,N_14933,N_13139);
nor U17928 (N_17928,N_13692,N_14091);
nor U17929 (N_17929,N_13045,N_14754);
and U17930 (N_17930,N_13164,N_15273);
nand U17931 (N_17931,N_14935,N_13326);
and U17932 (N_17932,N_12823,N_12858);
xor U17933 (N_17933,N_15391,N_12705);
or U17934 (N_17934,N_15549,N_13515);
xnor U17935 (N_17935,N_13045,N_13190);
xnor U17936 (N_17936,N_13591,N_13135);
or U17937 (N_17937,N_14617,N_13259);
and U17938 (N_17938,N_12865,N_12618);
nand U17939 (N_17939,N_15169,N_12978);
and U17940 (N_17940,N_12770,N_12710);
xnor U17941 (N_17941,N_13233,N_12772);
nand U17942 (N_17942,N_13964,N_13325);
and U17943 (N_17943,N_13651,N_14324);
nor U17944 (N_17944,N_14378,N_13992);
nor U17945 (N_17945,N_15135,N_14656);
or U17946 (N_17946,N_12654,N_14090);
nand U17947 (N_17947,N_12742,N_13890);
nor U17948 (N_17948,N_13614,N_13849);
and U17949 (N_17949,N_15401,N_13228);
nand U17950 (N_17950,N_13189,N_15607);
nand U17951 (N_17951,N_13235,N_13867);
or U17952 (N_17952,N_14014,N_13385);
nand U17953 (N_17953,N_12676,N_14947);
nand U17954 (N_17954,N_13853,N_14853);
nand U17955 (N_17955,N_13419,N_15545);
nand U17956 (N_17956,N_15170,N_14007);
or U17957 (N_17957,N_14347,N_15218);
or U17958 (N_17958,N_13204,N_15039);
nor U17959 (N_17959,N_14280,N_13553);
nand U17960 (N_17960,N_13506,N_15612);
or U17961 (N_17961,N_12669,N_14350);
or U17962 (N_17962,N_15161,N_14865);
nor U17963 (N_17963,N_14648,N_14466);
nand U17964 (N_17964,N_13598,N_13482);
nand U17965 (N_17965,N_13419,N_13537);
nor U17966 (N_17966,N_13945,N_12772);
or U17967 (N_17967,N_14970,N_14895);
and U17968 (N_17968,N_15517,N_15119);
or U17969 (N_17969,N_13412,N_14431);
and U17970 (N_17970,N_12996,N_14559);
nor U17971 (N_17971,N_15523,N_12617);
xor U17972 (N_17972,N_13879,N_14626);
nor U17973 (N_17973,N_13323,N_12731);
nor U17974 (N_17974,N_14138,N_14850);
and U17975 (N_17975,N_12828,N_12603);
xor U17976 (N_17976,N_15599,N_13461);
xor U17977 (N_17977,N_14633,N_14770);
nor U17978 (N_17978,N_14437,N_15143);
and U17979 (N_17979,N_14212,N_14668);
or U17980 (N_17980,N_14632,N_14918);
or U17981 (N_17981,N_13900,N_13197);
nand U17982 (N_17982,N_14864,N_14450);
nand U17983 (N_17983,N_15224,N_14379);
or U17984 (N_17984,N_14424,N_15085);
and U17985 (N_17985,N_13352,N_13464);
or U17986 (N_17986,N_13732,N_13585);
nor U17987 (N_17987,N_14385,N_13452);
and U17988 (N_17988,N_14889,N_12926);
and U17989 (N_17989,N_13463,N_12837);
nand U17990 (N_17990,N_14566,N_15205);
nand U17991 (N_17991,N_12851,N_15243);
nor U17992 (N_17992,N_13636,N_14276);
nor U17993 (N_17993,N_13525,N_13359);
xor U17994 (N_17994,N_14278,N_14966);
xor U17995 (N_17995,N_14055,N_12968);
nor U17996 (N_17996,N_14756,N_14131);
and U17997 (N_17997,N_13132,N_15038);
nand U17998 (N_17998,N_13725,N_14520);
nand U17999 (N_17999,N_15522,N_13635);
or U18000 (N_18000,N_15084,N_12980);
nand U18001 (N_18001,N_12706,N_13277);
or U18002 (N_18002,N_13936,N_14947);
xnor U18003 (N_18003,N_13578,N_15359);
nor U18004 (N_18004,N_12884,N_12890);
and U18005 (N_18005,N_14016,N_13685);
or U18006 (N_18006,N_14332,N_14473);
or U18007 (N_18007,N_15014,N_13868);
and U18008 (N_18008,N_13923,N_14298);
and U18009 (N_18009,N_14426,N_13682);
nand U18010 (N_18010,N_13898,N_14478);
or U18011 (N_18011,N_12939,N_13223);
xor U18012 (N_18012,N_13227,N_13172);
or U18013 (N_18013,N_12555,N_13726);
or U18014 (N_18014,N_12809,N_15072);
nor U18015 (N_18015,N_13347,N_12687);
and U18016 (N_18016,N_14091,N_15483);
and U18017 (N_18017,N_15547,N_14091);
nor U18018 (N_18018,N_15231,N_14215);
nand U18019 (N_18019,N_13119,N_12516);
nand U18020 (N_18020,N_13947,N_13903);
nand U18021 (N_18021,N_12921,N_12658);
xnor U18022 (N_18022,N_13211,N_14664);
and U18023 (N_18023,N_14712,N_13623);
or U18024 (N_18024,N_15003,N_13438);
nand U18025 (N_18025,N_14104,N_12941);
and U18026 (N_18026,N_14862,N_15401);
or U18027 (N_18027,N_15472,N_15306);
nor U18028 (N_18028,N_13357,N_14042);
or U18029 (N_18029,N_14962,N_14848);
and U18030 (N_18030,N_13338,N_13063);
nor U18031 (N_18031,N_13034,N_14413);
xor U18032 (N_18032,N_12560,N_14746);
and U18033 (N_18033,N_13755,N_13930);
or U18034 (N_18034,N_13205,N_14279);
nand U18035 (N_18035,N_13041,N_14326);
nand U18036 (N_18036,N_12976,N_12831);
and U18037 (N_18037,N_14346,N_13982);
xnor U18038 (N_18038,N_14605,N_13080);
nor U18039 (N_18039,N_13648,N_12763);
and U18040 (N_18040,N_15463,N_13390);
and U18041 (N_18041,N_14284,N_14531);
nand U18042 (N_18042,N_13278,N_12836);
nand U18043 (N_18043,N_13691,N_15249);
nand U18044 (N_18044,N_12678,N_14266);
or U18045 (N_18045,N_15449,N_14898);
xor U18046 (N_18046,N_13458,N_14913);
and U18047 (N_18047,N_12530,N_13378);
nand U18048 (N_18048,N_12857,N_13474);
and U18049 (N_18049,N_15162,N_15027);
and U18050 (N_18050,N_12697,N_14972);
xnor U18051 (N_18051,N_13729,N_14843);
nand U18052 (N_18052,N_13731,N_13213);
and U18053 (N_18053,N_14208,N_13791);
or U18054 (N_18054,N_14057,N_13855);
and U18055 (N_18055,N_12629,N_13966);
nor U18056 (N_18056,N_12992,N_14361);
xnor U18057 (N_18057,N_15329,N_15558);
nand U18058 (N_18058,N_12568,N_12592);
or U18059 (N_18059,N_14342,N_14267);
nor U18060 (N_18060,N_14789,N_15447);
and U18061 (N_18061,N_14371,N_14080);
and U18062 (N_18062,N_14406,N_12510);
or U18063 (N_18063,N_13184,N_13269);
or U18064 (N_18064,N_15275,N_13143);
xor U18065 (N_18065,N_15406,N_13609);
nand U18066 (N_18066,N_14859,N_14858);
nor U18067 (N_18067,N_15038,N_12883);
nand U18068 (N_18068,N_14734,N_13932);
and U18069 (N_18069,N_15605,N_15359);
nor U18070 (N_18070,N_15558,N_15521);
xor U18071 (N_18071,N_14647,N_13064);
or U18072 (N_18072,N_15113,N_13822);
nand U18073 (N_18073,N_13433,N_14576);
nand U18074 (N_18074,N_15247,N_12857);
xnor U18075 (N_18075,N_13033,N_15249);
and U18076 (N_18076,N_12991,N_12731);
xor U18077 (N_18077,N_14889,N_14018);
and U18078 (N_18078,N_14348,N_12856);
and U18079 (N_18079,N_13530,N_12885);
nand U18080 (N_18080,N_14037,N_13206);
or U18081 (N_18081,N_14581,N_14616);
or U18082 (N_18082,N_13108,N_14455);
nor U18083 (N_18083,N_14931,N_12721);
or U18084 (N_18084,N_15450,N_15513);
xnor U18085 (N_18085,N_14704,N_12625);
nand U18086 (N_18086,N_12554,N_13561);
nand U18087 (N_18087,N_12837,N_13217);
or U18088 (N_18088,N_15027,N_13708);
and U18089 (N_18089,N_14790,N_12978);
or U18090 (N_18090,N_15075,N_13264);
or U18091 (N_18091,N_13421,N_14429);
or U18092 (N_18092,N_12971,N_15429);
or U18093 (N_18093,N_13692,N_13617);
nand U18094 (N_18094,N_14188,N_13685);
nand U18095 (N_18095,N_15421,N_13504);
or U18096 (N_18096,N_13758,N_15538);
or U18097 (N_18097,N_13315,N_12643);
or U18098 (N_18098,N_14353,N_15441);
nor U18099 (N_18099,N_14004,N_12852);
or U18100 (N_18100,N_15402,N_13666);
nor U18101 (N_18101,N_13081,N_15424);
or U18102 (N_18102,N_15028,N_14756);
and U18103 (N_18103,N_13682,N_14301);
nand U18104 (N_18104,N_14137,N_13490);
and U18105 (N_18105,N_15599,N_13799);
xnor U18106 (N_18106,N_14556,N_14417);
or U18107 (N_18107,N_14061,N_14912);
and U18108 (N_18108,N_14782,N_14382);
or U18109 (N_18109,N_15364,N_14345);
nor U18110 (N_18110,N_15210,N_14722);
and U18111 (N_18111,N_12829,N_13504);
nand U18112 (N_18112,N_15182,N_12662);
xnor U18113 (N_18113,N_14315,N_13959);
xor U18114 (N_18114,N_14106,N_14362);
nand U18115 (N_18115,N_14919,N_12999);
and U18116 (N_18116,N_14074,N_14720);
nor U18117 (N_18117,N_14887,N_14833);
or U18118 (N_18118,N_12785,N_15260);
nand U18119 (N_18119,N_13633,N_12538);
and U18120 (N_18120,N_13894,N_15521);
xor U18121 (N_18121,N_14373,N_12639);
nor U18122 (N_18122,N_14405,N_14796);
and U18123 (N_18123,N_15009,N_14220);
or U18124 (N_18124,N_15038,N_15388);
and U18125 (N_18125,N_14259,N_13397);
nand U18126 (N_18126,N_14689,N_13452);
nor U18127 (N_18127,N_12651,N_15400);
and U18128 (N_18128,N_12944,N_14959);
nor U18129 (N_18129,N_12596,N_13750);
nor U18130 (N_18130,N_15283,N_13783);
xor U18131 (N_18131,N_13321,N_13697);
or U18132 (N_18132,N_12840,N_15106);
nor U18133 (N_18133,N_14984,N_14488);
and U18134 (N_18134,N_13686,N_14556);
xnor U18135 (N_18135,N_12598,N_12616);
or U18136 (N_18136,N_13161,N_13414);
nor U18137 (N_18137,N_13318,N_14118);
nor U18138 (N_18138,N_12761,N_14909);
xnor U18139 (N_18139,N_15518,N_14606);
and U18140 (N_18140,N_14636,N_14579);
nand U18141 (N_18141,N_13032,N_13758);
nand U18142 (N_18142,N_14266,N_15024);
nand U18143 (N_18143,N_14927,N_13772);
nor U18144 (N_18144,N_14281,N_12970);
nand U18145 (N_18145,N_13222,N_14634);
nor U18146 (N_18146,N_13152,N_13752);
or U18147 (N_18147,N_14284,N_14757);
xor U18148 (N_18148,N_14739,N_14997);
nor U18149 (N_18149,N_14783,N_13112);
and U18150 (N_18150,N_14118,N_14374);
nor U18151 (N_18151,N_14963,N_13382);
nor U18152 (N_18152,N_12796,N_12776);
or U18153 (N_18153,N_14999,N_13484);
or U18154 (N_18154,N_12577,N_14931);
xor U18155 (N_18155,N_14858,N_14715);
or U18156 (N_18156,N_13833,N_15456);
nand U18157 (N_18157,N_13586,N_14625);
nor U18158 (N_18158,N_14171,N_14495);
and U18159 (N_18159,N_12990,N_15458);
xnor U18160 (N_18160,N_15063,N_14745);
nor U18161 (N_18161,N_15358,N_13361);
nor U18162 (N_18162,N_14523,N_14919);
nor U18163 (N_18163,N_13005,N_14146);
and U18164 (N_18164,N_14724,N_14264);
or U18165 (N_18165,N_12926,N_15387);
or U18166 (N_18166,N_14392,N_14709);
or U18167 (N_18167,N_12551,N_14283);
nand U18168 (N_18168,N_14640,N_15231);
or U18169 (N_18169,N_12615,N_13836);
and U18170 (N_18170,N_12757,N_13907);
and U18171 (N_18171,N_13097,N_15459);
and U18172 (N_18172,N_15193,N_12970);
xor U18173 (N_18173,N_14795,N_13025);
nand U18174 (N_18174,N_12983,N_14023);
nor U18175 (N_18175,N_12833,N_15065);
nand U18176 (N_18176,N_14410,N_14488);
nand U18177 (N_18177,N_12587,N_13284);
nor U18178 (N_18178,N_13193,N_13184);
nor U18179 (N_18179,N_13992,N_14773);
nor U18180 (N_18180,N_15349,N_13553);
nand U18181 (N_18181,N_13965,N_14074);
nand U18182 (N_18182,N_12700,N_15108);
or U18183 (N_18183,N_14612,N_13282);
and U18184 (N_18184,N_14077,N_12729);
and U18185 (N_18185,N_12858,N_13967);
nand U18186 (N_18186,N_15201,N_12935);
nor U18187 (N_18187,N_13232,N_12616);
nor U18188 (N_18188,N_13572,N_12882);
nand U18189 (N_18189,N_13913,N_13998);
nand U18190 (N_18190,N_14329,N_14980);
or U18191 (N_18191,N_14640,N_13336);
and U18192 (N_18192,N_12775,N_12609);
nand U18193 (N_18193,N_13814,N_13668);
or U18194 (N_18194,N_13702,N_13067);
and U18195 (N_18195,N_13301,N_13972);
nor U18196 (N_18196,N_14337,N_12542);
or U18197 (N_18197,N_14678,N_14483);
or U18198 (N_18198,N_15226,N_14368);
and U18199 (N_18199,N_14654,N_13479);
or U18200 (N_18200,N_15424,N_12668);
nand U18201 (N_18201,N_12949,N_15177);
and U18202 (N_18202,N_13156,N_14731);
nand U18203 (N_18203,N_15022,N_13339);
or U18204 (N_18204,N_14588,N_12507);
xor U18205 (N_18205,N_12839,N_13425);
nor U18206 (N_18206,N_14637,N_13673);
nor U18207 (N_18207,N_13573,N_13558);
nand U18208 (N_18208,N_15476,N_12546);
and U18209 (N_18209,N_12650,N_14924);
nand U18210 (N_18210,N_14144,N_14539);
xnor U18211 (N_18211,N_12929,N_13877);
and U18212 (N_18212,N_14286,N_12595);
nand U18213 (N_18213,N_14946,N_13847);
and U18214 (N_18214,N_14499,N_14791);
or U18215 (N_18215,N_13677,N_15393);
nand U18216 (N_18216,N_13616,N_14968);
nor U18217 (N_18217,N_13558,N_12778);
xor U18218 (N_18218,N_15299,N_12631);
or U18219 (N_18219,N_13497,N_14635);
nor U18220 (N_18220,N_15216,N_15497);
or U18221 (N_18221,N_13965,N_13966);
xor U18222 (N_18222,N_13954,N_15336);
or U18223 (N_18223,N_14405,N_13559);
and U18224 (N_18224,N_13477,N_14464);
xnor U18225 (N_18225,N_15063,N_13153);
and U18226 (N_18226,N_12591,N_12632);
xnor U18227 (N_18227,N_13791,N_13423);
nand U18228 (N_18228,N_13264,N_13729);
and U18229 (N_18229,N_14506,N_15188);
nor U18230 (N_18230,N_13698,N_15601);
and U18231 (N_18231,N_12828,N_12879);
or U18232 (N_18232,N_15375,N_14369);
nand U18233 (N_18233,N_14078,N_13514);
or U18234 (N_18234,N_14270,N_13056);
and U18235 (N_18235,N_15025,N_15242);
nor U18236 (N_18236,N_14564,N_14783);
and U18237 (N_18237,N_13983,N_14963);
or U18238 (N_18238,N_14592,N_14051);
and U18239 (N_18239,N_13771,N_13232);
and U18240 (N_18240,N_12688,N_13089);
nor U18241 (N_18241,N_13377,N_15555);
and U18242 (N_18242,N_12519,N_14594);
or U18243 (N_18243,N_15468,N_12605);
and U18244 (N_18244,N_14195,N_12783);
nand U18245 (N_18245,N_13558,N_13440);
and U18246 (N_18246,N_13608,N_13284);
nand U18247 (N_18247,N_12819,N_13011);
nor U18248 (N_18248,N_15370,N_12593);
or U18249 (N_18249,N_13045,N_14787);
nand U18250 (N_18250,N_13155,N_15110);
nand U18251 (N_18251,N_15261,N_14014);
and U18252 (N_18252,N_13381,N_12926);
xnor U18253 (N_18253,N_13108,N_12872);
and U18254 (N_18254,N_14591,N_14114);
or U18255 (N_18255,N_13443,N_15196);
nor U18256 (N_18256,N_15006,N_13569);
nand U18257 (N_18257,N_13288,N_13843);
xor U18258 (N_18258,N_14542,N_12783);
and U18259 (N_18259,N_14663,N_14803);
nor U18260 (N_18260,N_13653,N_13867);
and U18261 (N_18261,N_14817,N_13923);
xnor U18262 (N_18262,N_13677,N_14047);
or U18263 (N_18263,N_15534,N_14320);
nand U18264 (N_18264,N_15400,N_14425);
xnor U18265 (N_18265,N_13895,N_15129);
or U18266 (N_18266,N_15263,N_15470);
or U18267 (N_18267,N_14581,N_15174);
or U18268 (N_18268,N_14711,N_13454);
and U18269 (N_18269,N_13816,N_15484);
or U18270 (N_18270,N_14688,N_12681);
xnor U18271 (N_18271,N_13930,N_13719);
nor U18272 (N_18272,N_13111,N_14382);
nor U18273 (N_18273,N_15312,N_13979);
nor U18274 (N_18274,N_14361,N_14803);
and U18275 (N_18275,N_15552,N_13351);
nand U18276 (N_18276,N_14772,N_13047);
and U18277 (N_18277,N_15283,N_13976);
and U18278 (N_18278,N_14691,N_13493);
and U18279 (N_18279,N_14315,N_12825);
nand U18280 (N_18280,N_14930,N_14846);
or U18281 (N_18281,N_12703,N_13623);
and U18282 (N_18282,N_14668,N_12819);
nand U18283 (N_18283,N_15506,N_15431);
and U18284 (N_18284,N_15028,N_14304);
or U18285 (N_18285,N_12866,N_15443);
and U18286 (N_18286,N_13493,N_12870);
xor U18287 (N_18287,N_14326,N_15411);
xor U18288 (N_18288,N_13003,N_12914);
xor U18289 (N_18289,N_15112,N_15011);
xor U18290 (N_18290,N_14416,N_15478);
nand U18291 (N_18291,N_12677,N_14072);
and U18292 (N_18292,N_15294,N_15056);
and U18293 (N_18293,N_15091,N_14750);
nand U18294 (N_18294,N_14109,N_14189);
nand U18295 (N_18295,N_13231,N_13524);
nand U18296 (N_18296,N_14800,N_15326);
nand U18297 (N_18297,N_14258,N_12763);
nand U18298 (N_18298,N_15248,N_14881);
or U18299 (N_18299,N_15465,N_14262);
and U18300 (N_18300,N_15218,N_13024);
nand U18301 (N_18301,N_14132,N_15560);
nand U18302 (N_18302,N_14863,N_15335);
xor U18303 (N_18303,N_14269,N_13907);
nor U18304 (N_18304,N_14837,N_15316);
nor U18305 (N_18305,N_14816,N_13885);
or U18306 (N_18306,N_15480,N_13135);
nand U18307 (N_18307,N_13172,N_13007);
or U18308 (N_18308,N_13407,N_13841);
and U18309 (N_18309,N_15028,N_15510);
and U18310 (N_18310,N_13380,N_13663);
and U18311 (N_18311,N_12608,N_12980);
and U18312 (N_18312,N_13069,N_14903);
nand U18313 (N_18313,N_14033,N_14774);
and U18314 (N_18314,N_12635,N_15249);
xor U18315 (N_18315,N_13707,N_13721);
nor U18316 (N_18316,N_13845,N_14530);
and U18317 (N_18317,N_15159,N_15220);
or U18318 (N_18318,N_15164,N_12663);
xor U18319 (N_18319,N_14753,N_13076);
or U18320 (N_18320,N_13674,N_15548);
nand U18321 (N_18321,N_14154,N_15617);
nand U18322 (N_18322,N_14283,N_14638);
nand U18323 (N_18323,N_14642,N_14764);
and U18324 (N_18324,N_14396,N_13864);
or U18325 (N_18325,N_13598,N_15599);
nor U18326 (N_18326,N_15498,N_12917);
nand U18327 (N_18327,N_14657,N_15491);
and U18328 (N_18328,N_13710,N_14931);
or U18329 (N_18329,N_15117,N_14648);
and U18330 (N_18330,N_12602,N_14373);
nand U18331 (N_18331,N_13988,N_15189);
or U18332 (N_18332,N_12942,N_12692);
and U18333 (N_18333,N_14470,N_15269);
xor U18334 (N_18334,N_13297,N_14857);
nor U18335 (N_18335,N_13919,N_14816);
nor U18336 (N_18336,N_15186,N_12781);
and U18337 (N_18337,N_13381,N_13305);
nor U18338 (N_18338,N_15162,N_14887);
nor U18339 (N_18339,N_13886,N_14616);
nor U18340 (N_18340,N_13028,N_15452);
nor U18341 (N_18341,N_14649,N_15515);
xnor U18342 (N_18342,N_13140,N_15391);
and U18343 (N_18343,N_15384,N_12572);
nand U18344 (N_18344,N_13266,N_13989);
and U18345 (N_18345,N_13597,N_13183);
and U18346 (N_18346,N_12937,N_12668);
or U18347 (N_18347,N_15447,N_14708);
nor U18348 (N_18348,N_13458,N_14473);
or U18349 (N_18349,N_14900,N_13186);
nor U18350 (N_18350,N_13843,N_13530);
xor U18351 (N_18351,N_14720,N_12729);
xor U18352 (N_18352,N_13421,N_13716);
and U18353 (N_18353,N_13297,N_14796);
and U18354 (N_18354,N_13968,N_14079);
and U18355 (N_18355,N_12707,N_14407);
nor U18356 (N_18356,N_12809,N_14541);
or U18357 (N_18357,N_13697,N_13734);
nand U18358 (N_18358,N_13691,N_15525);
nand U18359 (N_18359,N_12615,N_13819);
or U18360 (N_18360,N_15083,N_14483);
nor U18361 (N_18361,N_13911,N_14288);
and U18362 (N_18362,N_13877,N_15390);
nand U18363 (N_18363,N_14282,N_12855);
nor U18364 (N_18364,N_13882,N_14408);
xor U18365 (N_18365,N_15272,N_15545);
xnor U18366 (N_18366,N_12553,N_15505);
and U18367 (N_18367,N_14674,N_15221);
nand U18368 (N_18368,N_13380,N_15205);
xnor U18369 (N_18369,N_12615,N_14504);
nand U18370 (N_18370,N_13849,N_13440);
nor U18371 (N_18371,N_12818,N_12773);
and U18372 (N_18372,N_14709,N_13427);
and U18373 (N_18373,N_12837,N_15567);
or U18374 (N_18374,N_13465,N_13506);
nand U18375 (N_18375,N_13321,N_13216);
nand U18376 (N_18376,N_13014,N_12521);
and U18377 (N_18377,N_12599,N_15406);
or U18378 (N_18378,N_12749,N_14172);
or U18379 (N_18379,N_12510,N_12713);
nor U18380 (N_18380,N_13027,N_12970);
xor U18381 (N_18381,N_13353,N_15102);
xor U18382 (N_18382,N_14571,N_15494);
nand U18383 (N_18383,N_15098,N_14299);
nand U18384 (N_18384,N_13824,N_15592);
nand U18385 (N_18385,N_12977,N_13853);
or U18386 (N_18386,N_13054,N_14097);
or U18387 (N_18387,N_14459,N_13135);
or U18388 (N_18388,N_15251,N_13371);
nand U18389 (N_18389,N_15508,N_13175);
xor U18390 (N_18390,N_12878,N_14891);
or U18391 (N_18391,N_15227,N_13372);
and U18392 (N_18392,N_14993,N_13959);
and U18393 (N_18393,N_13104,N_15518);
nand U18394 (N_18394,N_15019,N_12991);
nor U18395 (N_18395,N_15411,N_13023);
and U18396 (N_18396,N_13697,N_12713);
nand U18397 (N_18397,N_14974,N_13682);
nor U18398 (N_18398,N_14607,N_13087);
or U18399 (N_18399,N_15376,N_13179);
nand U18400 (N_18400,N_15213,N_12705);
nor U18401 (N_18401,N_13280,N_12792);
or U18402 (N_18402,N_12815,N_13748);
and U18403 (N_18403,N_12543,N_13522);
xnor U18404 (N_18404,N_15465,N_13751);
xnor U18405 (N_18405,N_14665,N_12721);
nand U18406 (N_18406,N_15410,N_12584);
xor U18407 (N_18407,N_12892,N_12636);
or U18408 (N_18408,N_14725,N_12922);
nand U18409 (N_18409,N_12650,N_13892);
nor U18410 (N_18410,N_14646,N_13395);
nor U18411 (N_18411,N_15551,N_13051);
nand U18412 (N_18412,N_13884,N_14792);
or U18413 (N_18413,N_13234,N_14062);
nor U18414 (N_18414,N_14672,N_12717);
and U18415 (N_18415,N_14480,N_15017);
and U18416 (N_18416,N_14818,N_14121);
nor U18417 (N_18417,N_13452,N_15542);
and U18418 (N_18418,N_13174,N_15307);
and U18419 (N_18419,N_14806,N_12684);
nor U18420 (N_18420,N_15574,N_12998);
and U18421 (N_18421,N_13316,N_15158);
or U18422 (N_18422,N_13075,N_14167);
nand U18423 (N_18423,N_12699,N_15126);
or U18424 (N_18424,N_14805,N_14270);
nand U18425 (N_18425,N_15270,N_13959);
and U18426 (N_18426,N_12836,N_14707);
or U18427 (N_18427,N_12599,N_14537);
and U18428 (N_18428,N_12640,N_14700);
nand U18429 (N_18429,N_14958,N_15038);
nor U18430 (N_18430,N_12967,N_15391);
and U18431 (N_18431,N_14029,N_12933);
and U18432 (N_18432,N_14522,N_13708);
and U18433 (N_18433,N_15061,N_15208);
nand U18434 (N_18434,N_15290,N_14828);
nand U18435 (N_18435,N_14934,N_13448);
or U18436 (N_18436,N_13935,N_14723);
nor U18437 (N_18437,N_12974,N_13172);
and U18438 (N_18438,N_15367,N_13676);
or U18439 (N_18439,N_12854,N_13267);
nand U18440 (N_18440,N_13320,N_14782);
and U18441 (N_18441,N_13739,N_12893);
or U18442 (N_18442,N_14563,N_14418);
and U18443 (N_18443,N_12597,N_14114);
nand U18444 (N_18444,N_15356,N_13308);
and U18445 (N_18445,N_15139,N_14171);
nor U18446 (N_18446,N_12767,N_14418);
nand U18447 (N_18447,N_15577,N_12757);
xnor U18448 (N_18448,N_14081,N_12589);
or U18449 (N_18449,N_12809,N_15338);
or U18450 (N_18450,N_15156,N_13459);
nand U18451 (N_18451,N_14106,N_12878);
nor U18452 (N_18452,N_12518,N_13327);
xor U18453 (N_18453,N_13267,N_14119);
or U18454 (N_18454,N_14920,N_14357);
nand U18455 (N_18455,N_14816,N_14744);
nand U18456 (N_18456,N_14226,N_14434);
xnor U18457 (N_18457,N_14508,N_13336);
xor U18458 (N_18458,N_13763,N_14342);
nor U18459 (N_18459,N_13188,N_13147);
nor U18460 (N_18460,N_15344,N_13415);
xor U18461 (N_18461,N_15265,N_13136);
nand U18462 (N_18462,N_14657,N_13055);
nor U18463 (N_18463,N_13861,N_12964);
or U18464 (N_18464,N_15205,N_14492);
nor U18465 (N_18465,N_12978,N_15154);
xnor U18466 (N_18466,N_13638,N_14074);
nand U18467 (N_18467,N_15479,N_12625);
xnor U18468 (N_18468,N_14836,N_14147);
or U18469 (N_18469,N_13896,N_14642);
and U18470 (N_18470,N_15370,N_13698);
nand U18471 (N_18471,N_15048,N_15058);
and U18472 (N_18472,N_15437,N_14022);
xnor U18473 (N_18473,N_14785,N_14509);
nor U18474 (N_18474,N_12708,N_14748);
and U18475 (N_18475,N_15551,N_14793);
nand U18476 (N_18476,N_14066,N_13583);
nor U18477 (N_18477,N_13006,N_13455);
or U18478 (N_18478,N_13590,N_13596);
xnor U18479 (N_18479,N_13923,N_14734);
nand U18480 (N_18480,N_13706,N_14656);
and U18481 (N_18481,N_13867,N_12511);
nand U18482 (N_18482,N_12689,N_12897);
nor U18483 (N_18483,N_15491,N_14516);
nand U18484 (N_18484,N_14043,N_13380);
or U18485 (N_18485,N_14954,N_14725);
and U18486 (N_18486,N_13022,N_15000);
nand U18487 (N_18487,N_13470,N_14720);
xor U18488 (N_18488,N_14028,N_15049);
xnor U18489 (N_18489,N_13152,N_15202);
or U18490 (N_18490,N_12904,N_13759);
nor U18491 (N_18491,N_14721,N_14135);
nand U18492 (N_18492,N_14521,N_13141);
nor U18493 (N_18493,N_13238,N_13131);
nor U18494 (N_18494,N_15051,N_13431);
or U18495 (N_18495,N_14746,N_13679);
nor U18496 (N_18496,N_14195,N_13992);
nor U18497 (N_18497,N_15142,N_13974);
nand U18498 (N_18498,N_13452,N_13476);
nand U18499 (N_18499,N_13169,N_14944);
nand U18500 (N_18500,N_12574,N_15387);
or U18501 (N_18501,N_13294,N_13693);
or U18502 (N_18502,N_14599,N_15083);
or U18503 (N_18503,N_13582,N_15270);
xor U18504 (N_18504,N_13182,N_14142);
and U18505 (N_18505,N_12522,N_12705);
and U18506 (N_18506,N_14807,N_13212);
nor U18507 (N_18507,N_12606,N_12803);
xnor U18508 (N_18508,N_13183,N_13625);
nand U18509 (N_18509,N_14066,N_12993);
nor U18510 (N_18510,N_13621,N_15527);
nor U18511 (N_18511,N_13646,N_14457);
or U18512 (N_18512,N_13249,N_14303);
and U18513 (N_18513,N_13337,N_14974);
or U18514 (N_18514,N_12810,N_13508);
nand U18515 (N_18515,N_14621,N_13847);
or U18516 (N_18516,N_14193,N_15606);
or U18517 (N_18517,N_12621,N_13305);
and U18518 (N_18518,N_14465,N_15479);
nor U18519 (N_18519,N_13413,N_12604);
nor U18520 (N_18520,N_15266,N_14082);
or U18521 (N_18521,N_12686,N_15552);
nand U18522 (N_18522,N_15101,N_13426);
or U18523 (N_18523,N_13096,N_14223);
nor U18524 (N_18524,N_15622,N_15614);
nor U18525 (N_18525,N_12567,N_14255);
nand U18526 (N_18526,N_14393,N_13253);
and U18527 (N_18527,N_14772,N_12957);
nor U18528 (N_18528,N_14147,N_15587);
nand U18529 (N_18529,N_15438,N_13640);
nand U18530 (N_18530,N_13383,N_15103);
and U18531 (N_18531,N_13029,N_14247);
xnor U18532 (N_18532,N_12950,N_12908);
nand U18533 (N_18533,N_13434,N_12546);
or U18534 (N_18534,N_14667,N_13383);
nor U18535 (N_18535,N_15104,N_14445);
xnor U18536 (N_18536,N_14367,N_14892);
nor U18537 (N_18537,N_13944,N_13018);
xor U18538 (N_18538,N_14467,N_15569);
nor U18539 (N_18539,N_15106,N_14355);
and U18540 (N_18540,N_12767,N_15582);
xnor U18541 (N_18541,N_12553,N_13907);
or U18542 (N_18542,N_15539,N_13832);
and U18543 (N_18543,N_12538,N_15013);
xnor U18544 (N_18544,N_14518,N_12838);
xor U18545 (N_18545,N_15001,N_12844);
or U18546 (N_18546,N_12804,N_14134);
or U18547 (N_18547,N_13468,N_13018);
nand U18548 (N_18548,N_12614,N_15391);
xor U18549 (N_18549,N_13516,N_15527);
xnor U18550 (N_18550,N_14963,N_13829);
or U18551 (N_18551,N_12776,N_14159);
xor U18552 (N_18552,N_13160,N_12653);
nand U18553 (N_18553,N_14883,N_14651);
xnor U18554 (N_18554,N_15186,N_13703);
nor U18555 (N_18555,N_13753,N_13556);
nand U18556 (N_18556,N_15344,N_13835);
and U18557 (N_18557,N_13260,N_15563);
xnor U18558 (N_18558,N_15136,N_13649);
and U18559 (N_18559,N_12837,N_14969);
and U18560 (N_18560,N_14455,N_14565);
or U18561 (N_18561,N_14685,N_14544);
and U18562 (N_18562,N_13987,N_14198);
nor U18563 (N_18563,N_15465,N_14443);
nand U18564 (N_18564,N_13569,N_13986);
nand U18565 (N_18565,N_14824,N_12597);
and U18566 (N_18566,N_13219,N_14713);
xnor U18567 (N_18567,N_14898,N_13931);
nor U18568 (N_18568,N_12730,N_13049);
nor U18569 (N_18569,N_13978,N_13341);
or U18570 (N_18570,N_15105,N_13667);
or U18571 (N_18571,N_14999,N_14860);
and U18572 (N_18572,N_14361,N_14129);
and U18573 (N_18573,N_14521,N_14511);
or U18574 (N_18574,N_13223,N_15218);
nor U18575 (N_18575,N_12870,N_13978);
nand U18576 (N_18576,N_12943,N_14037);
nor U18577 (N_18577,N_15236,N_13388);
nor U18578 (N_18578,N_13980,N_14529);
nor U18579 (N_18579,N_12807,N_13658);
and U18580 (N_18580,N_15610,N_13505);
nand U18581 (N_18581,N_13293,N_13988);
and U18582 (N_18582,N_12576,N_13804);
or U18583 (N_18583,N_14135,N_13715);
nand U18584 (N_18584,N_15509,N_13455);
nand U18585 (N_18585,N_13605,N_13868);
nor U18586 (N_18586,N_14240,N_14195);
or U18587 (N_18587,N_15608,N_13515);
nand U18588 (N_18588,N_13073,N_12610);
nand U18589 (N_18589,N_13395,N_15072);
and U18590 (N_18590,N_15171,N_14555);
nor U18591 (N_18591,N_12500,N_15496);
and U18592 (N_18592,N_12866,N_12882);
or U18593 (N_18593,N_12979,N_14492);
nor U18594 (N_18594,N_13849,N_13457);
or U18595 (N_18595,N_12529,N_14445);
or U18596 (N_18596,N_15119,N_13780);
or U18597 (N_18597,N_14317,N_13797);
or U18598 (N_18598,N_15142,N_15366);
nor U18599 (N_18599,N_14419,N_13786);
nor U18600 (N_18600,N_13336,N_13154);
xnor U18601 (N_18601,N_14985,N_15067);
nand U18602 (N_18602,N_14153,N_15120);
and U18603 (N_18603,N_13632,N_13435);
and U18604 (N_18604,N_14906,N_15623);
nand U18605 (N_18605,N_12790,N_14129);
nand U18606 (N_18606,N_13263,N_14288);
or U18607 (N_18607,N_12824,N_13175);
nor U18608 (N_18608,N_14528,N_14842);
or U18609 (N_18609,N_14133,N_15018);
or U18610 (N_18610,N_13738,N_14257);
nor U18611 (N_18611,N_13034,N_13497);
and U18612 (N_18612,N_15196,N_15227);
or U18613 (N_18613,N_13444,N_15019);
xnor U18614 (N_18614,N_14598,N_13741);
and U18615 (N_18615,N_13910,N_15155);
and U18616 (N_18616,N_13328,N_14338);
and U18617 (N_18617,N_14504,N_13849);
nor U18618 (N_18618,N_15464,N_14316);
nand U18619 (N_18619,N_14948,N_15072);
nor U18620 (N_18620,N_15406,N_14688);
xor U18621 (N_18621,N_13363,N_12769);
nand U18622 (N_18622,N_13536,N_13849);
nor U18623 (N_18623,N_15530,N_12956);
or U18624 (N_18624,N_13072,N_14771);
nand U18625 (N_18625,N_13856,N_14118);
and U18626 (N_18626,N_13917,N_15272);
and U18627 (N_18627,N_12774,N_15472);
or U18628 (N_18628,N_14895,N_13472);
nor U18629 (N_18629,N_14086,N_13661);
and U18630 (N_18630,N_15091,N_14286);
or U18631 (N_18631,N_13335,N_13053);
nand U18632 (N_18632,N_13433,N_12754);
nor U18633 (N_18633,N_13582,N_14609);
nor U18634 (N_18634,N_12713,N_12786);
or U18635 (N_18635,N_14841,N_13605);
nor U18636 (N_18636,N_13917,N_14755);
nor U18637 (N_18637,N_15396,N_15203);
nor U18638 (N_18638,N_14374,N_12505);
or U18639 (N_18639,N_13757,N_15136);
nor U18640 (N_18640,N_15129,N_15410);
nor U18641 (N_18641,N_15050,N_13762);
or U18642 (N_18642,N_12876,N_14783);
nor U18643 (N_18643,N_14879,N_13642);
nand U18644 (N_18644,N_13602,N_12502);
nor U18645 (N_18645,N_13749,N_14826);
and U18646 (N_18646,N_12816,N_13938);
nand U18647 (N_18647,N_13733,N_14263);
nand U18648 (N_18648,N_14959,N_14724);
or U18649 (N_18649,N_13125,N_13908);
nor U18650 (N_18650,N_14833,N_13634);
or U18651 (N_18651,N_13198,N_13840);
and U18652 (N_18652,N_13149,N_14122);
and U18653 (N_18653,N_12614,N_13312);
xor U18654 (N_18654,N_15318,N_15002);
nand U18655 (N_18655,N_14230,N_15369);
or U18656 (N_18656,N_15178,N_15059);
xnor U18657 (N_18657,N_13139,N_14386);
nand U18658 (N_18658,N_12632,N_12906);
nand U18659 (N_18659,N_13918,N_13441);
and U18660 (N_18660,N_13227,N_13566);
nand U18661 (N_18661,N_13042,N_13102);
nor U18662 (N_18662,N_15390,N_15219);
nor U18663 (N_18663,N_14839,N_15187);
nor U18664 (N_18664,N_13543,N_15029);
nor U18665 (N_18665,N_14364,N_12549);
nand U18666 (N_18666,N_13931,N_13262);
and U18667 (N_18667,N_14792,N_14745);
or U18668 (N_18668,N_12857,N_14010);
and U18669 (N_18669,N_14790,N_13744);
nor U18670 (N_18670,N_15386,N_14013);
xnor U18671 (N_18671,N_14538,N_14286);
xnor U18672 (N_18672,N_14112,N_14144);
or U18673 (N_18673,N_14692,N_14932);
nor U18674 (N_18674,N_14926,N_13249);
xor U18675 (N_18675,N_13415,N_14472);
nand U18676 (N_18676,N_13361,N_15275);
nand U18677 (N_18677,N_13452,N_14568);
nand U18678 (N_18678,N_13864,N_12625);
nand U18679 (N_18679,N_13139,N_14099);
nor U18680 (N_18680,N_14304,N_15347);
nor U18681 (N_18681,N_15127,N_14632);
or U18682 (N_18682,N_13212,N_14552);
or U18683 (N_18683,N_14112,N_15605);
xor U18684 (N_18684,N_14549,N_12710);
and U18685 (N_18685,N_14390,N_13879);
xnor U18686 (N_18686,N_15468,N_13947);
or U18687 (N_18687,N_14578,N_14331);
and U18688 (N_18688,N_14301,N_13332);
and U18689 (N_18689,N_12580,N_13439);
or U18690 (N_18690,N_13865,N_12895);
nand U18691 (N_18691,N_12697,N_12724);
nand U18692 (N_18692,N_13720,N_13779);
nor U18693 (N_18693,N_12780,N_13811);
or U18694 (N_18694,N_14943,N_15553);
or U18695 (N_18695,N_13731,N_13652);
and U18696 (N_18696,N_12670,N_15211);
nor U18697 (N_18697,N_15410,N_14757);
nor U18698 (N_18698,N_13630,N_12506);
nand U18699 (N_18699,N_13853,N_13721);
or U18700 (N_18700,N_14286,N_15574);
and U18701 (N_18701,N_12511,N_13143);
and U18702 (N_18702,N_14323,N_14231);
or U18703 (N_18703,N_14397,N_13123);
or U18704 (N_18704,N_15295,N_12654);
or U18705 (N_18705,N_14738,N_13914);
nand U18706 (N_18706,N_12614,N_14810);
and U18707 (N_18707,N_13927,N_13792);
xnor U18708 (N_18708,N_14698,N_13621);
nand U18709 (N_18709,N_15129,N_13381);
and U18710 (N_18710,N_13902,N_13974);
and U18711 (N_18711,N_13553,N_14126);
and U18712 (N_18712,N_12979,N_15089);
nor U18713 (N_18713,N_13856,N_13396);
and U18714 (N_18714,N_13092,N_12729);
nand U18715 (N_18715,N_13199,N_12868);
or U18716 (N_18716,N_14830,N_12675);
nand U18717 (N_18717,N_12779,N_15450);
and U18718 (N_18718,N_12936,N_12884);
nand U18719 (N_18719,N_12524,N_13325);
nor U18720 (N_18720,N_13576,N_13464);
or U18721 (N_18721,N_14285,N_13490);
or U18722 (N_18722,N_14933,N_14705);
or U18723 (N_18723,N_13786,N_14481);
xnor U18724 (N_18724,N_14709,N_13717);
nand U18725 (N_18725,N_13876,N_15505);
nand U18726 (N_18726,N_13989,N_14815);
or U18727 (N_18727,N_13015,N_14770);
and U18728 (N_18728,N_14789,N_13949);
nand U18729 (N_18729,N_13369,N_13645);
nor U18730 (N_18730,N_14799,N_14293);
or U18731 (N_18731,N_14658,N_15086);
or U18732 (N_18732,N_13606,N_12927);
nor U18733 (N_18733,N_13360,N_13724);
nor U18734 (N_18734,N_13505,N_14820);
nand U18735 (N_18735,N_12527,N_13552);
nand U18736 (N_18736,N_15421,N_12944);
nand U18737 (N_18737,N_14978,N_13386);
nor U18738 (N_18738,N_13769,N_14524);
nand U18739 (N_18739,N_14140,N_13875);
xor U18740 (N_18740,N_13409,N_12724);
and U18741 (N_18741,N_14945,N_13776);
and U18742 (N_18742,N_15483,N_15386);
xnor U18743 (N_18743,N_12586,N_14425);
nor U18744 (N_18744,N_13521,N_13102);
xor U18745 (N_18745,N_15609,N_13952);
nand U18746 (N_18746,N_15061,N_13205);
or U18747 (N_18747,N_12925,N_15475);
nand U18748 (N_18748,N_13779,N_12967);
and U18749 (N_18749,N_13378,N_14210);
nor U18750 (N_18750,N_16275,N_16019);
xnor U18751 (N_18751,N_17947,N_17302);
nor U18752 (N_18752,N_17264,N_17709);
or U18753 (N_18753,N_16771,N_16029);
xnor U18754 (N_18754,N_17899,N_16893);
nor U18755 (N_18755,N_16245,N_17426);
nor U18756 (N_18756,N_16325,N_15752);
and U18757 (N_18757,N_16194,N_16673);
nand U18758 (N_18758,N_17390,N_16686);
nor U18759 (N_18759,N_17854,N_15710);
or U18760 (N_18760,N_16196,N_18577);
and U18761 (N_18761,N_18022,N_17469);
xnor U18762 (N_18762,N_17950,N_18486);
nor U18763 (N_18763,N_17253,N_17819);
nand U18764 (N_18764,N_18465,N_17946);
xnor U18765 (N_18765,N_18714,N_17943);
and U18766 (N_18766,N_16662,N_17746);
nor U18767 (N_18767,N_15878,N_15750);
and U18768 (N_18768,N_16649,N_18189);
nand U18769 (N_18769,N_18359,N_16391);
nor U18770 (N_18770,N_18507,N_16084);
and U18771 (N_18771,N_15704,N_16707);
nand U18772 (N_18772,N_18047,N_18171);
or U18773 (N_18773,N_16743,N_17763);
nand U18774 (N_18774,N_16976,N_17648);
nor U18775 (N_18775,N_17149,N_18588);
nand U18776 (N_18776,N_17631,N_17157);
nand U18777 (N_18777,N_17432,N_16972);
or U18778 (N_18778,N_16313,N_16967);
or U18779 (N_18779,N_17090,N_15656);
or U18780 (N_18780,N_16920,N_15879);
or U18781 (N_18781,N_16692,N_16484);
or U18782 (N_18782,N_18062,N_15918);
nand U18783 (N_18783,N_17225,N_16906);
nor U18784 (N_18784,N_17425,N_15856);
nand U18785 (N_18785,N_18529,N_16682);
nor U18786 (N_18786,N_16570,N_18457);
xnor U18787 (N_18787,N_18553,N_17133);
or U18788 (N_18788,N_17798,N_17224);
xnor U18789 (N_18789,N_16027,N_17686);
xnor U18790 (N_18790,N_16427,N_15821);
or U18791 (N_18791,N_18075,N_16980);
or U18792 (N_18792,N_17918,N_16031);
xor U18793 (N_18793,N_18254,N_16942);
xor U18794 (N_18794,N_17377,N_17927);
nand U18795 (N_18795,N_17681,N_16741);
and U18796 (N_18796,N_15733,N_15913);
nor U18797 (N_18797,N_18408,N_16362);
or U18798 (N_18798,N_17628,N_16536);
nor U18799 (N_18799,N_17705,N_16260);
xor U18800 (N_18800,N_17052,N_18098);
nor U18801 (N_18801,N_15994,N_18340);
or U18802 (N_18802,N_18721,N_17239);
and U18803 (N_18803,N_18327,N_16929);
or U18804 (N_18804,N_16677,N_16343);
nor U18805 (N_18805,N_17944,N_17385);
nand U18806 (N_18806,N_18664,N_16552);
nor U18807 (N_18807,N_17067,N_16255);
and U18808 (N_18808,N_16957,N_18459);
nand U18809 (N_18809,N_17732,N_18630);
nand U18810 (N_18810,N_18099,N_17679);
nand U18811 (N_18811,N_17036,N_18618);
nand U18812 (N_18812,N_18474,N_16602);
or U18813 (N_18813,N_18228,N_17735);
and U18814 (N_18814,N_16907,N_16804);
and U18815 (N_18815,N_18449,N_18334);
or U18816 (N_18816,N_17362,N_15977);
or U18817 (N_18817,N_18259,N_17363);
and U18818 (N_18818,N_18127,N_16795);
and U18819 (N_18819,N_17552,N_16699);
or U18820 (N_18820,N_16849,N_15953);
and U18821 (N_18821,N_17751,N_15708);
and U18822 (N_18822,N_16721,N_18628);
xnor U18823 (N_18823,N_15754,N_15844);
xnor U18824 (N_18824,N_16598,N_16955);
or U18825 (N_18825,N_15991,N_16358);
nand U18826 (N_18826,N_17372,N_16985);
or U18827 (N_18827,N_16149,N_15712);
and U18828 (N_18828,N_15843,N_17139);
and U18829 (N_18829,N_18199,N_18051);
nand U18830 (N_18830,N_16791,N_15764);
and U18831 (N_18831,N_17537,N_18447);
xor U18832 (N_18832,N_18413,N_15912);
and U18833 (N_18833,N_16750,N_17981);
xnor U18834 (N_18834,N_17241,N_15639);
and U18835 (N_18835,N_17146,N_15674);
or U18836 (N_18836,N_17894,N_18412);
or U18837 (N_18837,N_18016,N_16150);
nand U18838 (N_18838,N_16600,N_15812);
and U18839 (N_18839,N_15722,N_15935);
xor U18840 (N_18840,N_16319,N_16553);
nand U18841 (N_18841,N_17250,N_17439);
or U18842 (N_18842,N_17066,N_18702);
or U18843 (N_18843,N_17092,N_17830);
or U18844 (N_18844,N_16114,N_16641);
nand U18845 (N_18845,N_18514,N_16278);
or U18846 (N_18846,N_16695,N_16002);
or U18847 (N_18847,N_18320,N_15634);
nor U18848 (N_18848,N_15841,N_17419);
nand U18849 (N_18849,N_16819,N_16730);
nor U18850 (N_18850,N_18633,N_17243);
nand U18851 (N_18851,N_16198,N_16169);
or U18852 (N_18852,N_16377,N_16748);
nand U18853 (N_18853,N_18742,N_16818);
xor U18854 (N_18854,N_17436,N_16059);
xor U18855 (N_18855,N_17194,N_18673);
xor U18856 (N_18856,N_18530,N_16076);
nor U18857 (N_18857,N_16611,N_16646);
and U18858 (N_18858,N_15881,N_16666);
nand U18859 (N_18859,N_17109,N_16360);
xnor U18860 (N_18860,N_16859,N_18284);
nor U18861 (N_18861,N_17162,N_16307);
nor U18862 (N_18862,N_18521,N_17703);
and U18863 (N_18863,N_17995,N_18406);
nand U18864 (N_18864,N_17599,N_16161);
xnor U18865 (N_18865,N_17482,N_16619);
nand U18866 (N_18866,N_16135,N_18519);
and U18867 (N_18867,N_15740,N_17747);
nand U18868 (N_18868,N_15633,N_15840);
and U18869 (N_18869,N_17008,N_17657);
xnor U18870 (N_18870,N_18677,N_17799);
or U18871 (N_18871,N_15831,N_16527);
nor U18872 (N_18872,N_16235,N_15653);
xnor U18873 (N_18873,N_15728,N_18362);
nor U18874 (N_18874,N_18293,N_15926);
nor U18875 (N_18875,N_17455,N_15797);
or U18876 (N_18876,N_18023,N_18357);
and U18877 (N_18877,N_16020,N_15726);
xor U18878 (N_18878,N_18350,N_18073);
and U18879 (N_18879,N_15786,N_16228);
and U18880 (N_18880,N_17095,N_17204);
nor U18881 (N_18881,N_16668,N_17172);
xor U18882 (N_18882,N_17114,N_17730);
or U18883 (N_18883,N_16414,N_18031);
nor U18884 (N_18884,N_18451,N_17838);
xor U18885 (N_18885,N_17949,N_16894);
and U18886 (N_18886,N_16187,N_18065);
nor U18887 (N_18887,N_15875,N_15650);
and U18888 (N_18888,N_16386,N_17564);
nor U18889 (N_18889,N_18708,N_18580);
or U18890 (N_18890,N_17338,N_17589);
xor U18891 (N_18891,N_17471,N_15915);
and U18892 (N_18892,N_16452,N_17042);
nand U18893 (N_18893,N_17272,N_16921);
nor U18894 (N_18894,N_17260,N_16856);
or U18895 (N_18895,N_18568,N_17293);
and U18896 (N_18896,N_16503,N_16259);
and U18897 (N_18897,N_18114,N_18651);
nor U18898 (N_18898,N_18740,N_17378);
nand U18899 (N_18899,N_15891,N_18040);
and U18900 (N_18900,N_17654,N_18049);
xor U18901 (N_18901,N_15745,N_17930);
nand U18902 (N_18902,N_16191,N_17083);
and U18903 (N_18903,N_17676,N_18623);
nor U18904 (N_18904,N_16803,N_17937);
and U18905 (N_18905,N_16651,N_16069);
nand U18906 (N_18906,N_18272,N_16993);
nand U18907 (N_18907,N_18239,N_16635);
nand U18908 (N_18908,N_17812,N_18037);
nor U18909 (N_18909,N_17341,N_18043);
and U18910 (N_18910,N_17683,N_18123);
or U18911 (N_18911,N_17062,N_17043);
nand U18912 (N_18912,N_17970,N_17179);
or U18913 (N_18913,N_18288,N_15939);
and U18914 (N_18914,N_17847,N_17473);
and U18915 (N_18915,N_18308,N_15942);
and U18916 (N_18916,N_17125,N_18355);
or U18917 (N_18917,N_17326,N_18573);
and U18918 (N_18918,N_17921,N_16720);
or U18919 (N_18919,N_18556,N_16447);
nand U18920 (N_18920,N_18719,N_15852);
nand U18921 (N_18921,N_17101,N_16745);
and U18922 (N_18922,N_16417,N_16107);
nor U18923 (N_18923,N_17639,N_16590);
nand U18924 (N_18924,N_17410,N_18410);
nand U18925 (N_18925,N_16768,N_18059);
nor U18926 (N_18926,N_18369,N_16227);
nand U18927 (N_18927,N_18695,N_17601);
xnor U18928 (N_18928,N_17691,N_15738);
xnor U18929 (N_18929,N_17545,N_17213);
nand U18930 (N_18930,N_17667,N_15743);
or U18931 (N_18931,N_17532,N_17879);
or U18932 (N_18932,N_18068,N_15870);
nor U18933 (N_18933,N_17404,N_18693);
and U18934 (N_18934,N_17459,N_18250);
nand U18935 (N_18935,N_17697,N_16915);
or U18936 (N_18936,N_18496,N_17672);
nor U18937 (N_18937,N_17998,N_18282);
and U18938 (N_18938,N_16616,N_16630);
nand U18939 (N_18939,N_16075,N_17979);
or U18940 (N_18940,N_17767,N_15773);
nand U18941 (N_18941,N_16830,N_17642);
nor U18942 (N_18942,N_16332,N_18076);
xor U18943 (N_18943,N_16369,N_17718);
or U18944 (N_18944,N_16212,N_17619);
nand U18945 (N_18945,N_17489,N_17926);
or U18946 (N_18946,N_16866,N_15690);
nand U18947 (N_18947,N_16410,N_15793);
xnor U18948 (N_18948,N_17766,N_18435);
nand U18949 (N_18949,N_17118,N_16608);
nor U18950 (N_18950,N_17173,N_18650);
or U18951 (N_18951,N_15731,N_18642);
and U18952 (N_18952,N_17587,N_17817);
and U18953 (N_18953,N_17030,N_18038);
or U18954 (N_18954,N_15895,N_16058);
and U18955 (N_18955,N_15698,N_17959);
xor U18956 (N_18956,N_17165,N_17576);
and U18957 (N_18957,N_18088,N_17216);
nand U18958 (N_18958,N_16612,N_17184);
nand U18959 (N_18959,N_15958,N_18488);
nand U18960 (N_18960,N_15635,N_16806);
or U18961 (N_18961,N_16786,N_16537);
xor U18962 (N_18962,N_15869,N_17917);
nor U18963 (N_18963,N_16432,N_16565);
nor U18964 (N_18964,N_18417,N_17571);
and U18965 (N_18965,N_16204,N_16658);
or U18966 (N_18966,N_18376,N_18313);
nor U18967 (N_18967,N_18668,N_17491);
or U18968 (N_18968,N_15996,N_18363);
and U18969 (N_18969,N_15969,N_16374);
or U18970 (N_18970,N_18626,N_16437);
nand U18971 (N_18971,N_17063,N_18559);
nand U18972 (N_18972,N_16665,N_16688);
or U18973 (N_18973,N_18331,N_17038);
and U18974 (N_18974,N_16863,N_16162);
or U18975 (N_18975,N_17591,N_16130);
and U18976 (N_18976,N_17784,N_17574);
xor U18977 (N_18977,N_16816,N_16626);
nor U18978 (N_18978,N_17650,N_16798);
nand U18979 (N_18979,N_16861,N_18686);
or U18980 (N_18980,N_18211,N_16435);
or U18981 (N_18981,N_18318,N_17600);
nand U18982 (N_18982,N_15686,N_17230);
or U18983 (N_18983,N_15850,N_16039);
nand U18984 (N_18984,N_17311,N_17242);
nor U18985 (N_18985,N_15678,N_17866);
nand U18986 (N_18986,N_17181,N_16405);
xor U18987 (N_18987,N_16778,N_17147);
nand U18988 (N_18988,N_17586,N_16583);
or U18989 (N_18989,N_17986,N_17796);
nand U18990 (N_18990,N_17901,N_17595);
nor U18991 (N_18991,N_15711,N_16642);
nand U18992 (N_18992,N_17444,N_17609);
or U18993 (N_18993,N_18289,N_17757);
or U18994 (N_18994,N_15974,N_16463);
nand U18995 (N_18995,N_16564,N_15857);
nor U18996 (N_18996,N_16109,N_18011);
and U18997 (N_18997,N_18545,N_18205);
and U18998 (N_18998,N_16329,N_16389);
or U18999 (N_18999,N_17973,N_18006);
nand U19000 (N_19000,N_15887,N_16850);
or U19001 (N_19001,N_17261,N_18394);
and U19002 (N_19002,N_16505,N_18180);
and U19003 (N_19003,N_15748,N_16314);
nand U19004 (N_19004,N_17785,N_16787);
and U19005 (N_19005,N_18203,N_17441);
or U19006 (N_19006,N_16070,N_17256);
or U19007 (N_19007,N_15964,N_18213);
and U19008 (N_19008,N_18347,N_17025);
or U19009 (N_19009,N_17675,N_15871);
xnor U19010 (N_19010,N_18454,N_16013);
and U19011 (N_19011,N_18540,N_16961);
and U19012 (N_19012,N_16534,N_17288);
or U19013 (N_19013,N_18079,N_16296);
nand U19014 (N_19014,N_15819,N_16017);
nor U19015 (N_19015,N_16354,N_16821);
nand U19016 (N_19016,N_17312,N_17435);
nand U19017 (N_19017,N_15898,N_16025);
xor U19018 (N_19018,N_16148,N_17266);
or U19019 (N_19019,N_18492,N_16182);
nor U19020 (N_19020,N_16078,N_16831);
or U19021 (N_19021,N_16953,N_17662);
nor U19022 (N_19022,N_17400,N_16810);
xor U19023 (N_19023,N_16220,N_17327);
nor U19024 (N_19024,N_16004,N_17249);
nand U19025 (N_19025,N_18300,N_17374);
nor U19026 (N_19026,N_17989,N_16223);
or U19027 (N_19027,N_16835,N_15890);
nand U19028 (N_19028,N_16740,N_16108);
or U19029 (N_19029,N_17132,N_17904);
or U19030 (N_19030,N_18298,N_17105);
and U19031 (N_19031,N_18297,N_16346);
or U19032 (N_19032,N_15669,N_17702);
and U19033 (N_19033,N_16136,N_18166);
nor U19034 (N_19034,N_15968,N_16226);
or U19035 (N_19035,N_17647,N_15874);
and U19036 (N_19036,N_18498,N_17097);
xnor U19037 (N_19037,N_15792,N_16874);
nand U19038 (N_19038,N_18629,N_16011);
or U19039 (N_19039,N_18683,N_15769);
nand U19040 (N_19040,N_16497,N_18636);
nor U19041 (N_19041,N_15908,N_17658);
or U19042 (N_19042,N_18685,N_17047);
and U19043 (N_19043,N_18008,N_18129);
nand U19044 (N_19044,N_18523,N_16522);
and U19045 (N_19045,N_18306,N_15734);
xor U19046 (N_19046,N_16691,N_16573);
or U19047 (N_19047,N_16008,N_18341);
xnor U19048 (N_19048,N_16186,N_16322);
or U19049 (N_19049,N_16378,N_16962);
nor U19050 (N_19050,N_15700,N_15693);
nor U19051 (N_19051,N_17049,N_18130);
nand U19052 (N_19052,N_18305,N_16726);
or U19053 (N_19053,N_18030,N_18572);
nand U19054 (N_19054,N_17701,N_18366);
and U19055 (N_19055,N_18360,N_16916);
or U19056 (N_19056,N_16170,N_17726);
nor U19057 (N_19057,N_15956,N_18167);
nand U19058 (N_19058,N_18344,N_16395);
nor U19059 (N_19059,N_16206,N_17403);
or U19060 (N_19060,N_16218,N_18632);
and U19061 (N_19061,N_15791,N_17684);
or U19062 (N_19062,N_16940,N_18328);
nand U19063 (N_19063,N_17834,N_17508);
xor U19064 (N_19064,N_17512,N_17916);
nand U19065 (N_19065,N_18562,N_18330);
or U19066 (N_19066,N_17493,N_17237);
and U19067 (N_19067,N_16678,N_16670);
or U19068 (N_19068,N_16241,N_18440);
nor U19069 (N_19069,N_16345,N_16842);
nor U19070 (N_19070,N_17258,N_16142);
or U19071 (N_19071,N_16053,N_16034);
nand U19072 (N_19072,N_15709,N_16979);
nor U19073 (N_19073,N_17211,N_16763);
nand U19074 (N_19074,N_17855,N_15940);
nor U19075 (N_19075,N_16828,N_17106);
nor U19076 (N_19076,N_16003,N_18491);
or U19077 (N_19077,N_15910,N_16257);
or U19078 (N_19078,N_16939,N_16949);
xor U19079 (N_19079,N_18072,N_16023);
or U19080 (N_19080,N_18617,N_16706);
nand U19081 (N_19081,N_17723,N_16769);
or U19082 (N_19082,N_16569,N_15729);
and U19083 (N_19083,N_16301,N_16634);
or U19084 (N_19084,N_16383,N_17696);
and U19085 (N_19085,N_15685,N_17310);
or U19086 (N_19086,N_17706,N_17023);
and U19087 (N_19087,N_16637,N_17993);
nand U19088 (N_19088,N_17168,N_18225);
nand U19089 (N_19089,N_16363,N_18042);
nor U19090 (N_19090,N_17623,N_17058);
and U19091 (N_19091,N_15882,N_18212);
nand U19092 (N_19092,N_16290,N_17883);
and U19093 (N_19093,N_18120,N_18220);
xor U19094 (N_19094,N_17020,N_16254);
and U19095 (N_19095,N_17728,N_18728);
or U19096 (N_19096,N_17939,N_16772);
and U19097 (N_19097,N_17368,N_17167);
and U19098 (N_19098,N_15931,N_16625);
nand U19099 (N_19099,N_16101,N_16411);
nand U19100 (N_19100,N_16617,N_16126);
nor U19101 (N_19101,N_17221,N_16057);
or U19102 (N_19102,N_17543,N_15691);
nand U19103 (N_19103,N_18713,N_16247);
nor U19104 (N_19104,N_18625,N_16782);
or U19105 (N_19105,N_16171,N_17206);
xor U19106 (N_19106,N_17313,N_16917);
xor U19107 (N_19107,N_18733,N_18661);
or U19108 (N_19108,N_17274,N_15664);
xnor U19109 (N_19109,N_18218,N_17014);
or U19110 (N_19110,N_15855,N_17197);
nor U19111 (N_19111,N_17547,N_17100);
or U19112 (N_19112,N_17559,N_16994);
or U19113 (N_19113,N_16765,N_17890);
or U19114 (N_19114,N_16216,N_16181);
and U19115 (N_19115,N_17273,N_17254);
nor U19116 (N_19116,N_17123,N_18247);
and U19117 (N_19117,N_18301,N_18467);
and U19118 (N_19118,N_18196,N_17613);
nand U19119 (N_19119,N_16016,N_17096);
and U19120 (N_19120,N_16908,N_16252);
and U19121 (N_19121,N_17522,N_16337);
or U19122 (N_19122,N_17467,N_16521);
nor U19123 (N_19123,N_16041,N_18471);
or U19124 (N_19124,N_17652,N_17526);
or U19125 (N_19125,N_17081,N_18525);
and U19126 (N_19126,N_17695,N_16457);
nand U19127 (N_19127,N_17490,N_16511);
and U19128 (N_19128,N_17958,N_18444);
and U19129 (N_19129,N_15695,N_16280);
or U19130 (N_19130,N_16103,N_17850);
xnor U19131 (N_19131,N_18278,N_16758);
nor U19132 (N_19132,N_16281,N_16334);
or U19133 (N_19133,N_17379,N_16871);
and U19134 (N_19134,N_16456,N_18416);
or U19135 (N_19135,N_18383,N_17091);
nand U19136 (N_19136,N_15846,N_18063);
or U19137 (N_19137,N_17335,N_16284);
or U19138 (N_19138,N_15950,N_16586);
or U19139 (N_19139,N_17257,N_18161);
nor U19140 (N_19140,N_15767,N_18690);
nand U19141 (N_19141,N_18653,N_18624);
nor U19142 (N_19142,N_18108,N_16288);
nor U19143 (N_19143,N_17663,N_18361);
nand U19144 (N_19144,N_18245,N_17016);
nand U19145 (N_19145,N_15725,N_16555);
or U19146 (N_19146,N_18044,N_18512);
nand U19147 (N_19147,N_15981,N_18370);
or U19148 (N_19148,N_18005,N_18490);
nand U19149 (N_19149,N_18419,N_18185);
nor U19150 (N_19150,N_15658,N_16424);
nand U19151 (N_19151,N_18688,N_18662);
or U19152 (N_19152,N_18154,N_18267);
and U19153 (N_19153,N_15759,N_16530);
and U19154 (N_19154,N_17656,N_16685);
nand U19155 (N_19155,N_16163,N_16141);
nor U19156 (N_19156,N_18158,N_17578);
or U19157 (N_19157,N_18548,N_17321);
and U19158 (N_19158,N_15842,N_15679);
xnor U19159 (N_19159,N_18299,N_17307);
xor U19160 (N_19160,N_18578,N_16467);
nand U19161 (N_19161,N_18339,N_16326);
and U19162 (N_19162,N_18443,N_17568);
nor U19163 (N_19163,N_16793,N_17720);
nand U19164 (N_19164,N_16300,N_18382);
or U19165 (N_19165,N_17107,N_17810);
nor U19166 (N_19166,N_16895,N_15798);
or U19167 (N_19167,N_17655,N_18277);
and U19168 (N_19168,N_18433,N_17597);
xnor U19169 (N_19169,N_15696,N_16415);
or U19170 (N_19170,N_16507,N_16622);
and U19171 (N_19171,N_18329,N_15860);
nand U19172 (N_19172,N_17861,N_15957);
and U19173 (N_19173,N_16614,N_17622);
and U19174 (N_19174,N_15736,N_15825);
nand U19175 (N_19175,N_16200,N_18101);
and U19176 (N_19176,N_15744,N_18132);
or U19177 (N_19177,N_17160,N_17427);
nand U19178 (N_19178,N_16797,N_17217);
and U19179 (N_19179,N_16509,N_18058);
or U19180 (N_19180,N_15967,N_17821);
nor U19181 (N_19181,N_18506,N_17113);
xor U19182 (N_19182,N_16838,N_17477);
or U19183 (N_19183,N_18082,N_16705);
xor U19184 (N_19184,N_16618,N_16207);
nor U19185 (N_19185,N_16267,N_16251);
and U19186 (N_19186,N_17053,N_17178);
nand U19187 (N_19187,N_18711,N_18106);
nor U19188 (N_19188,N_15681,N_18258);
nor U19189 (N_19189,N_17382,N_18025);
nor U19190 (N_19190,N_17409,N_17928);
nor U19191 (N_19191,N_17610,N_17069);
and U19192 (N_19192,N_17964,N_16698);
or U19193 (N_19193,N_17128,N_17028);
or U19194 (N_19194,N_18224,N_18012);
or U19195 (N_19195,N_17953,N_16192);
nor U19196 (N_19196,N_17833,N_16572);
nand U19197 (N_19197,N_15801,N_17465);
nor U19198 (N_19198,N_16195,N_17389);
nor U19199 (N_19199,N_18694,N_16533);
nand U19200 (N_19200,N_18178,N_18381);
nand U19201 (N_19201,N_16128,N_17176);
nand U19202 (N_19202,N_17494,N_18671);
nor U19203 (N_19203,N_17910,N_17187);
nor U19204 (N_19204,N_15946,N_17102);
nor U19205 (N_19205,N_16203,N_18179);
nor U19206 (N_19206,N_15641,N_16609);
and U19207 (N_19207,N_16860,N_16119);
and U19208 (N_19208,N_17451,N_16621);
and U19209 (N_19209,N_17521,N_17867);
nor U19210 (N_19210,N_18215,N_16802);
nand U19211 (N_19211,N_18276,N_17740);
nand U19212 (N_19212,N_17129,N_17297);
xnor U19213 (N_19213,N_18173,N_16018);
nand U19214 (N_19214,N_16975,N_16134);
and U19215 (N_19215,N_17431,N_15659);
and U19216 (N_19216,N_17772,N_18269);
xor U19217 (N_19217,N_15781,N_18738);
nand U19218 (N_19218,N_17764,N_17698);
nand U19219 (N_19219,N_16106,N_16843);
nand U19220 (N_19220,N_18372,N_16129);
nand U19221 (N_19221,N_16291,N_16164);
nor U19222 (N_19222,N_16814,N_15989);
and U19223 (N_19223,N_17103,N_16143);
nand U19224 (N_19224,N_17802,N_17486);
and U19225 (N_19225,N_18152,N_16471);
and U19226 (N_19226,N_16189,N_15911);
or U19227 (N_19227,N_17787,N_18516);
or U19228 (N_19228,N_17836,N_15719);
or U19229 (N_19229,N_17112,N_16111);
nor U19230 (N_19230,N_18232,N_17888);
nand U19231 (N_19231,N_17487,N_16233);
and U19232 (N_19232,N_16661,N_18703);
or U19233 (N_19233,N_18549,N_18183);
or U19234 (N_19234,N_16948,N_16954);
and U19235 (N_19235,N_17715,N_17267);
and U19236 (N_19236,N_18319,N_16178);
nor U19237 (N_19237,N_18397,N_18071);
nand U19238 (N_19238,N_17792,N_18122);
and U19239 (N_19239,N_17054,N_16669);
and U19240 (N_19240,N_18260,N_18718);
and U19241 (N_19241,N_18256,N_18579);
or U19242 (N_19242,N_15809,N_18332);
nand U19243 (N_19243,N_18274,N_16501);
nand U19244 (N_19244,N_16478,N_17566);
and U19245 (N_19245,N_15803,N_18565);
nor U19246 (N_19246,N_16425,N_17605);
and U19247 (N_19247,N_15697,N_18286);
and U19248 (N_19248,N_16919,N_16969);
nand U19249 (N_19249,N_18292,N_17670);
and U19250 (N_19250,N_18066,N_16146);
nor U19251 (N_19251,N_16010,N_15742);
and U19252 (N_19252,N_15999,N_18036);
and U19253 (N_19253,N_16393,N_17397);
nand U19254 (N_19254,N_15859,N_17882);
and U19255 (N_19255,N_17422,N_16050);
and U19256 (N_19256,N_16640,N_16671);
nand U19257 (N_19257,N_18725,N_17627);
and U19258 (N_19258,N_17134,N_17572);
and U19259 (N_19259,N_15770,N_16878);
or U19260 (N_19260,N_16581,N_17891);
nor U19261 (N_19261,N_16468,N_15984);
or U19262 (N_19262,N_17219,N_18188);
nor U19263 (N_19263,N_17629,N_17474);
nor U19264 (N_19264,N_17753,N_16742);
nand U19265 (N_19265,N_15675,N_15929);
and U19266 (N_19266,N_15862,N_16366);
and U19267 (N_19267,N_16951,N_17806);
and U19268 (N_19268,N_15902,N_17366);
xor U19269 (N_19269,N_16829,N_18145);
xor U19270 (N_19270,N_18124,N_16090);
nand U19271 (N_19271,N_17453,N_16382);
or U19272 (N_19272,N_16327,N_17721);
and U19273 (N_19273,N_15783,N_18197);
xnor U19274 (N_19274,N_17634,N_17665);
and U19275 (N_19275,N_16451,N_17398);
and U19276 (N_19276,N_16924,N_15796);
or U19277 (N_19277,N_16987,N_16493);
and U19278 (N_19278,N_18316,N_18706);
nand U19279 (N_19279,N_15927,N_17438);
nand U19280 (N_19280,N_16629,N_16836);
or U19281 (N_19281,N_17196,N_16304);
or U19282 (N_19282,N_16780,N_18091);
xor U19283 (N_19283,N_16855,N_18448);
or U19284 (N_19284,N_15990,N_16180);
and U19285 (N_19285,N_18162,N_17170);
xnor U19286 (N_19286,N_17837,N_16077);
or U19287 (N_19287,N_15788,N_15919);
xor U19288 (N_19288,N_18547,N_18494);
and U19289 (N_19289,N_15776,N_17548);
and U19290 (N_19290,N_16239,N_18317);
and U19291 (N_19291,N_15626,N_17089);
or U19292 (N_19292,N_17978,N_17068);
and U19293 (N_19293,N_17189,N_15732);
nand U19294 (N_19294,N_16356,N_18140);
or U19295 (N_19295,N_18561,N_17447);
or U19296 (N_19296,N_17611,N_16238);
nand U19297 (N_19297,N_16599,N_17166);
or U19298 (N_19298,N_18414,N_16545);
and U19299 (N_19299,N_16097,N_17514);
or U19300 (N_19300,N_18726,N_16124);
xnor U19301 (N_19301,N_16561,N_15807);
nor U19302 (N_19302,N_15627,N_18396);
nand U19303 (N_19303,N_16439,N_15917);
nand U19304 (N_19304,N_16429,N_18312);
or U19305 (N_19305,N_17843,N_17516);
xnor U19306 (N_19306,N_17470,N_16690);
and U19307 (N_19307,N_18112,N_18182);
and U19308 (N_19308,N_17885,N_16152);
nor U19309 (N_19309,N_16335,N_17614);
nor U19310 (N_19310,N_16294,N_18614);
or U19311 (N_19311,N_17872,N_15665);
nor U19312 (N_19312,N_18520,N_16406);
or U19313 (N_19313,N_18655,N_18364);
or U19314 (N_19314,N_16909,N_18594);
nor U19315 (N_19315,N_16494,N_18131);
nand U19316 (N_19316,N_15921,N_18248);
and U19317 (N_19317,N_16689,N_18153);
xnor U19318 (N_19318,N_16455,N_18337);
xnor U19319 (N_19319,N_18736,N_18654);
nor U19320 (N_19320,N_16479,N_17569);
nand U19321 (N_19321,N_16991,N_16444);
nand U19322 (N_19322,N_17524,N_17413);
or U19323 (N_19323,N_18460,N_15723);
nand U19324 (N_19324,N_16263,N_17278);
nor U19325 (N_19325,N_17011,N_18453);
nor U19326 (N_19326,N_16202,N_16460);
nor U19327 (N_19327,N_16585,N_16234);
nand U19328 (N_19328,N_17719,N_17355);
nor U19329 (N_19329,N_17280,N_17277);
nand U19330 (N_19330,N_16805,N_17895);
and U19331 (N_19331,N_18024,N_18349);
nand U19332 (N_19332,N_17227,N_16535);
and U19333 (N_19333,N_18184,N_17015);
and U19334 (N_19334,N_17955,N_18209);
or U19335 (N_19335,N_15955,N_17004);
nor U19336 (N_19336,N_18583,N_16096);
nor U19337 (N_19337,N_16639,N_18064);
and U19338 (N_19338,N_17298,N_18169);
xnor U19339 (N_19339,N_17231,N_18518);
nand U19340 (N_19340,N_18281,N_15947);
or U19341 (N_19341,N_15998,N_18354);
and U19342 (N_19342,N_16399,N_17897);
and U19343 (N_19343,N_17974,N_17561);
nor U19344 (N_19344,N_16309,N_18659);
nor U19345 (N_19345,N_17775,N_17632);
or U19346 (N_19346,N_18119,N_18658);
and U19347 (N_19347,N_15972,N_17161);
nand U19348 (N_19348,N_16531,N_16384);
and U19349 (N_19349,N_18021,N_17037);
nand U19350 (N_19350,N_16711,N_17558);
or U19351 (N_19351,N_16205,N_15787);
and U19352 (N_19352,N_17394,N_18696);
xor U19353 (N_19353,N_18027,N_16990);
nand U19354 (N_19354,N_15834,N_16001);
and U19355 (N_19355,N_16638,N_18377);
or U19356 (N_19356,N_18729,N_17649);
or U19357 (N_19357,N_17805,N_15986);
nand U19358 (N_19358,N_18724,N_16099);
and U19359 (N_19359,N_17760,N_18151);
nand U19360 (N_19360,N_18590,N_15824);
xnor U19361 (N_19361,N_16714,N_17992);
nor U19362 (N_19362,N_17517,N_18165);
or U19363 (N_19363,N_18502,N_18242);
nor U19364 (N_19364,N_16352,N_17301);
nor U19365 (N_19365,N_18170,N_16038);
nand U19366 (N_19366,N_17737,N_18265);
and U19367 (N_19367,N_18141,N_16775);
nand U19368 (N_19368,N_16490,N_17815);
nand U19369 (N_19369,N_17878,N_17971);
nand U19370 (N_19370,N_17961,N_17940);
or U19371 (N_19371,N_15800,N_17829);
nor U19372 (N_19372,N_16965,N_17148);
or U19373 (N_19373,N_17433,N_17164);
nand U19374 (N_19374,N_17626,N_17511);
or U19375 (N_19375,N_16529,N_15720);
nand U19376 (N_19376,N_18136,N_15886);
nor U19377 (N_19377,N_16330,N_17428);
nor U19378 (N_19378,N_15717,N_15960);
nor U19379 (N_19379,N_17434,N_16502);
and U19380 (N_19380,N_17130,N_17457);
or U19381 (N_19381,N_17346,N_17045);
nor U19382 (N_19382,N_17527,N_16062);
or U19383 (N_19383,N_16672,N_17804);
and U19384 (N_19384,N_16005,N_17975);
nor U19385 (N_19385,N_15993,N_16177);
or U19386 (N_19386,N_18380,N_18296);
or U19387 (N_19387,N_18351,N_17606);
or U19388 (N_19388,N_17500,N_16421);
xor U19389 (N_19389,N_16824,N_17761);
nor U19390 (N_19390,N_17716,N_16952);
nor U19391 (N_19391,N_17445,N_17383);
or U19392 (N_19392,N_16576,N_18020);
nand U19393 (N_19393,N_18094,N_17556);
or U19394 (N_19394,N_17013,N_17329);
or U19395 (N_19395,N_17956,N_16890);
or U19396 (N_19396,N_18148,N_16100);
or U19397 (N_19397,N_18035,N_15845);
nand U19398 (N_19398,N_17304,N_17859);
nor U19399 (N_19399,N_18747,N_16209);
and U19400 (N_19400,N_17604,N_18616);
nor U19401 (N_19401,N_16681,N_16823);
nor U19402 (N_19402,N_17314,N_17027);
nand U19403 (N_19403,N_16557,N_17592);
and U19404 (N_19404,N_18698,N_17188);
nand U19405 (N_19405,N_17932,N_16837);
nand U19406 (N_19406,N_17271,N_15768);
and U19407 (N_19407,N_16213,N_15706);
nand U19408 (N_19408,N_18200,N_18398);
nor U19409 (N_19409,N_17029,N_15692);
nor U19410 (N_19410,N_17777,N_18236);
or U19411 (N_19411,N_16458,N_18214);
nor U19412 (N_19412,N_16744,N_16368);
and U19413 (N_19413,N_16562,N_17481);
and U19414 (N_19414,N_17464,N_17198);
and U19415 (N_19415,N_16873,N_15643);
or U19416 (N_19416,N_17158,N_16801);
and U19417 (N_19417,N_18660,N_17593);
xor U19418 (N_19418,N_16515,N_16470);
nor U19419 (N_19419,N_18393,N_16597);
and U19420 (N_19420,N_18303,N_15963);
and U19421 (N_19421,N_17531,N_17156);
nor U19422 (N_19422,N_15737,N_17443);
nand U19423 (N_19423,N_18699,N_17065);
nor U19424 (N_19424,N_16350,N_18202);
and U19425 (N_19425,N_18386,N_18257);
nor U19426 (N_19426,N_17240,N_16081);
nor U19427 (N_19427,N_18420,N_18640);
or U19428 (N_19428,N_17440,N_18504);
nand U19429 (N_19429,N_16500,N_15657);
and U19430 (N_19430,N_16925,N_16443);
nand U19431 (N_19431,N_18587,N_16604);
nor U19432 (N_19432,N_18111,N_17286);
xnor U19433 (N_19433,N_18230,N_16766);
xnor U19434 (N_19434,N_15925,N_16506);
or U19435 (N_19435,N_16904,N_16541);
nand U19436 (N_19436,N_16400,N_15866);
or U19437 (N_19437,N_16118,N_17907);
and U19438 (N_19438,N_15761,N_17332);
nor U19439 (N_19439,N_15985,N_18532);
nand U19440 (N_19440,N_16409,N_17839);
nand U19441 (N_19441,N_17842,N_18600);
nor U19442 (N_19442,N_17873,N_17152);
or U19443 (N_19443,N_16032,N_17050);
and U19444 (N_19444,N_17220,N_16913);
nor U19445 (N_19445,N_18458,N_18589);
and U19446 (N_19446,N_15804,N_16093);
or U19447 (N_19447,N_18712,N_17497);
nand U19448 (N_19448,N_16657,N_16000);
nor U19449 (N_19449,N_16933,N_17690);
nor U19450 (N_19450,N_15982,N_15785);
nor U19451 (N_19451,N_16885,N_16243);
nor U19452 (N_19452,N_17660,N_18375);
xnor U19453 (N_19453,N_16922,N_17538);
nor U19454 (N_19454,N_16560,N_18056);
xnor U19455 (N_19455,N_16250,N_18493);
nor U19456 (N_19456,N_17209,N_18746);
or U19457 (N_19457,N_17922,N_16396);
nor U19458 (N_19458,N_17699,N_18418);
or U19459 (N_19459,N_16485,N_16588);
nor U19460 (N_19460,N_18426,N_18596);
and U19461 (N_19461,N_16174,N_16813);
and U19462 (N_19462,N_18749,N_16796);
xor U19463 (N_19463,N_18595,N_18385);
xnor U19464 (N_19464,N_18591,N_17789);
or U19465 (N_19465,N_18680,N_15835);
xor U19466 (N_19466,N_16722,N_17825);
nor U19467 (N_19467,N_17294,N_17263);
nor U19468 (N_19468,N_17929,N_17039);
and U19469 (N_19469,N_16727,N_16728);
nor U19470 (N_19470,N_16516,N_17229);
or U19471 (N_19471,N_17768,N_17640);
nand U19472 (N_19472,N_18472,N_17952);
or U19473 (N_19473,N_16297,N_18544);
or U19474 (N_19474,N_16655,N_18684);
nor U19475 (N_19475,N_16870,N_15688);
nand U19476 (N_19476,N_16935,N_18424);
xor U19477 (N_19477,N_16168,N_16089);
or U19478 (N_19478,N_17594,N_17339);
or U19479 (N_19479,N_15885,N_16615);
and U19480 (N_19480,N_18422,N_17247);
or U19481 (N_19481,N_16977,N_18470);
nand U19482 (N_19482,N_16353,N_18222);
nor U19483 (N_19483,N_17215,N_16342);
or U19484 (N_19484,N_16268,N_18552);
nor U19485 (N_19485,N_17416,N_16249);
or U19486 (N_19486,N_16660,N_15839);
or U19487 (N_19487,N_16115,N_18048);
or U19488 (N_19488,N_17071,N_18261);
and U19489 (N_19489,N_16310,N_17463);
or U19490 (N_19490,N_16215,N_16858);
xor U19491 (N_19491,N_16402,N_18116);
nand U19492 (N_19492,N_15705,N_15873);
nor U19493 (N_19493,N_16684,N_17319);
and U19494 (N_19494,N_18275,N_16088);
nand U19495 (N_19495,N_17121,N_17519);
and U19496 (N_19496,N_16809,N_17205);
or U19497 (N_19497,N_17340,N_16208);
nand U19498 (N_19498,N_17533,N_18262);
nor U19499 (N_19499,N_15655,N_16499);
or U19500 (N_19500,N_15640,N_16375);
nor U19501 (N_19501,N_17391,N_18061);
nor U19502 (N_19502,N_16882,N_16755);
and U19503 (N_19503,N_18569,N_18113);
nand U19504 (N_19504,N_15823,N_18400);
xor U19505 (N_19505,N_17429,N_16139);
and U19506 (N_19506,N_17962,N_16927);
and U19507 (N_19507,N_15863,N_15739);
nand U19508 (N_19508,N_18026,N_16548);
or U19509 (N_19509,N_17603,N_17317);
nand U19510 (N_19510,N_16276,N_16887);
nor U19511 (N_19511,N_15880,N_16958);
nand U19512 (N_19512,N_18194,N_16155);
or U19513 (N_19513,N_17175,N_15684);
and U19514 (N_19514,N_16418,N_17581);
xor U19515 (N_19515,N_17750,N_17908);
nand U19516 (N_19516,N_16015,N_16983);
or U19517 (N_19517,N_17567,N_17057);
and U19518 (N_19518,N_18374,N_16733);
and U19519 (N_19519,N_17823,N_18700);
or U19520 (N_19520,N_18315,N_17159);
xnor U19521 (N_19521,N_17646,N_17779);
or U19522 (N_19522,N_17040,N_15822);
and U19523 (N_19523,N_18602,N_17722);
nand U19524 (N_19524,N_15746,N_16550);
nor U19525 (N_19525,N_18574,N_15909);
and U19526 (N_19526,N_16584,N_16504);
nor U19527 (N_19527,N_17583,N_16080);
or U19528 (N_19528,N_18584,N_18430);
xor U19529 (N_19529,N_18001,N_17303);
nand U19530 (N_19530,N_17997,N_18147);
nor U19531 (N_19531,N_17807,N_15888);
nor U19532 (N_19532,N_17295,N_16989);
nand U19533 (N_19533,N_18070,N_17458);
or U19534 (N_19534,N_17137,N_17886);
nor U19535 (N_19535,N_18709,N_16580);
nand U19536 (N_19536,N_17064,N_15638);
and U19537 (N_19537,N_17275,N_16464);
or U19538 (N_19538,N_16944,N_17911);
or U19539 (N_19539,N_15753,N_16664);
nor U19540 (N_19540,N_16394,N_18034);
xnor U19541 (N_19541,N_18599,N_18295);
xnor U19542 (N_19542,N_17342,N_15699);
or U19543 (N_19543,N_17315,N_16946);
xnor U19544 (N_19544,N_16792,N_18644);
xnor U19545 (N_19545,N_16926,N_16361);
nor U19546 (N_19546,N_16269,N_16122);
nand U19547 (N_19547,N_16784,N_18388);
nand U19548 (N_19548,N_15721,N_16514);
nand U19549 (N_19549,N_18285,N_17153);
nand U19550 (N_19550,N_17174,N_17098);
nor U19551 (N_19551,N_18450,N_16133);
xor U19552 (N_19552,N_17865,N_16312);
nor U19553 (N_19553,N_18495,N_16659);
xor U19554 (N_19554,N_17046,N_15795);
or U19555 (N_19555,N_17505,N_17442);
nand U19556 (N_19556,N_17708,N_16610);
nand U19557 (N_19557,N_18681,N_15983);
nor U19558 (N_19558,N_16007,N_16035);
and U19559 (N_19559,N_17305,N_18456);
and U19560 (N_19560,N_18007,N_16292);
and U19561 (N_19561,N_15892,N_15630);
nor U19562 (N_19562,N_17612,N_17248);
nand U19563 (N_19563,N_17233,N_17523);
nor U19564 (N_19564,N_18368,N_16092);
and U19565 (N_19565,N_15661,N_16481);
nand U19566 (N_19566,N_16082,N_17831);
nand U19567 (N_19567,N_17857,N_16132);
or U19568 (N_19568,N_15905,N_18311);
or U19569 (N_19569,N_17108,N_18566);
or U19570 (N_19570,N_16071,N_18446);
and U19571 (N_19571,N_17226,N_18325);
nand U19572 (N_19572,N_18053,N_18353);
nor U19573 (N_19573,N_17762,N_16419);
nand U19574 (N_19574,N_16518,N_18367);
nor U19575 (N_19575,N_17641,N_18032);
nand U19576 (N_19576,N_17557,N_16624);
nand U19577 (N_19577,N_16526,N_16603);
nand U19578 (N_19578,N_17456,N_15757);
or U19579 (N_19579,N_15811,N_16336);
xor U19580 (N_19580,N_16911,N_18135);
nand U19581 (N_19581,N_17835,N_16528);
nand U19582 (N_19582,N_16982,N_17948);
xnor U19583 (N_19583,N_15673,N_15995);
nand U19584 (N_19584,N_15779,N_15799);
nand U19585 (N_19585,N_18157,N_17353);
nand U19586 (N_19586,N_18647,N_18323);
nand U19587 (N_19587,N_16480,N_18358);
or U19588 (N_19588,N_15671,N_16116);
xor U19589 (N_19589,N_16153,N_16285);
or U19590 (N_19590,N_15782,N_17700);
nor U19591 (N_19591,N_16397,N_17373);
nor U19592 (N_19592,N_18270,N_18666);
or U19593 (N_19593,N_16482,N_16848);
nor U19594 (N_19594,N_17573,N_17687);
xor U19595 (N_19595,N_16270,N_16700);
xor U19596 (N_19596,N_18528,N_16862);
and U19597 (N_19597,N_17783,N_16434);
nor U19598 (N_19598,N_17420,N_18139);
nand U19599 (N_19599,N_15660,N_18739);
and U19600 (N_19600,N_16138,N_16365);
xnor U19601 (N_19601,N_17544,N_16715);
nand U19602 (N_19602,N_17418,N_18050);
xnor U19603 (N_19603,N_16654,N_18604);
xor U19604 (N_19604,N_17841,N_18732);
xnor U19605 (N_19605,N_17078,N_16320);
nor U19606 (N_19606,N_17462,N_17881);
or U19607 (N_19607,N_16477,N_16466);
or U19608 (N_19608,N_18177,N_15682);
nand U19609 (N_19609,N_17941,N_17299);
nand U19610 (N_19610,N_18253,N_16995);
xnor U19611 (N_19611,N_17669,N_16589);
nor U19612 (N_19612,N_16201,N_16224);
xor U19613 (N_19613,N_18345,N_16112);
nand U19614 (N_19614,N_15802,N_18084);
nand U19615 (N_19615,N_17534,N_16520);
and U19616 (N_19616,N_17673,N_17554);
and U19617 (N_19617,N_16773,N_15867);
nand U19618 (N_19618,N_17704,N_15930);
or U19619 (N_19619,N_16800,N_18192);
nand U19620 (N_19620,N_17048,N_16087);
xor U19621 (N_19621,N_16188,N_16045);
or U19622 (N_19622,N_16538,N_18054);
nand U19623 (N_19623,N_17893,N_16543);
or U19624 (N_19624,N_16749,N_18399);
and U19625 (N_19625,N_16879,N_17688);
nand U19626 (N_19626,N_16757,N_17912);
nand U19627 (N_19627,N_17437,N_17724);
or U19628 (N_19628,N_18144,N_16303);
nand U19629 (N_19629,N_17963,N_18627);
or U19630 (N_19630,N_17803,N_17495);
or U19631 (N_19631,N_16338,N_16794);
xnor U19632 (N_19632,N_17635,N_17369);
nor U19633 (N_19633,N_16172,N_18610);
and U19634 (N_19634,N_17144,N_17848);
xnor U19635 (N_19635,N_16311,N_18631);
nor U19636 (N_19636,N_18455,N_16446);
nor U19637 (N_19637,N_17844,N_17323);
nand U19638 (N_19638,N_15938,N_18142);
or U19639 (N_19639,N_18181,N_15952);
and U19640 (N_19640,N_15900,N_17086);
and U19641 (N_19641,N_15934,N_17320);
and U19642 (N_19642,N_16702,N_16453);
and U19643 (N_19643,N_17744,N_18302);
nand U19644 (N_19644,N_18500,N_15945);
nor U19645 (N_19645,N_18401,N_17513);
nor U19646 (N_19646,N_16854,N_15662);
or U19647 (N_19647,N_16052,N_16065);
and U19648 (N_19648,N_17991,N_16696);
or U19649 (N_19649,N_17423,N_17077);
nand U19650 (N_19650,N_16880,N_17392);
and U19651 (N_19651,N_15756,N_15973);
nor U19652 (N_19652,N_18674,N_18606);
and U19653 (N_19653,N_16851,N_18527);
and U19654 (N_19654,N_17478,N_17485);
xnor U19655 (N_19655,N_18509,N_17270);
or U19656 (N_19656,N_18710,N_18226);
and U19657 (N_19657,N_16667,N_17896);
and U19658 (N_19658,N_17060,N_16620);
nand U19659 (N_19659,N_16910,N_17851);
nand U19660 (N_19660,N_18705,N_17736);
and U19661 (N_19661,N_17330,N_17001);
and U19662 (N_19662,N_15631,N_17005);
nor U19663 (N_19663,N_16724,N_17801);
or U19664 (N_19664,N_16596,N_16554);
or U19665 (N_19665,N_18321,N_18510);
nor U19666 (N_19666,N_16373,N_18077);
and U19667 (N_19667,N_16864,N_18240);
or U19668 (N_19668,N_18191,N_16959);
or U19669 (N_19669,N_18052,N_18309);
nand U19670 (N_19670,N_18146,N_15978);
and U19671 (N_19671,N_17154,N_16892);
nor U19672 (N_19672,N_16877,N_17421);
nor U19673 (N_19673,N_18691,N_17507);
and U19674 (N_19674,N_16759,N_17238);
or U19675 (N_19675,N_18538,N_15980);
nand U19676 (N_19676,N_18597,N_17415);
or U19677 (N_19677,N_15741,N_17365);
or U19678 (N_19678,N_17006,N_17645);
nand U19679 (N_19679,N_17920,N_17529);
nand U19680 (N_19680,N_16754,N_17245);
or U19681 (N_19681,N_15965,N_18687);
and U19682 (N_19682,N_18638,N_18537);
and U19683 (N_19683,N_15814,N_16986);
xor U19684 (N_19684,N_16872,N_16197);
and U19685 (N_19685,N_18227,N_15636);
nand U19686 (N_19686,N_17283,N_18121);
nor U19687 (N_19687,N_18551,N_18670);
nor U19688 (N_19688,N_16708,N_17009);
nor U19689 (N_19689,N_17653,N_16046);
or U19690 (N_19690,N_16779,N_17010);
nor U19691 (N_19691,N_17200,N_18168);
and U19692 (N_19692,N_17727,N_16416);
nor U19693 (N_19693,N_18432,N_17909);
nor U19694 (N_19694,N_16299,N_17717);
nor U19695 (N_19695,N_17671,N_18542);
or U19696 (N_19696,N_16712,N_16328);
nand U19697 (N_19697,N_16433,N_16653);
and U19698 (N_19698,N_18338,N_18263);
or U19699 (N_19699,N_16380,N_17289);
and U19700 (N_19700,N_15941,N_17689);
and U19701 (N_19701,N_17793,N_17210);
or U19702 (N_19702,N_17965,N_17472);
nand U19703 (N_19703,N_17985,N_18234);
and U19704 (N_19704,N_18365,N_18571);
or U19705 (N_19705,N_17430,N_18387);
and U19706 (N_19706,N_18723,N_16486);
and U19707 (N_19707,N_18000,N_15907);
nor U19708 (N_19708,N_17520,N_16592);
nor U19709 (N_19709,N_16996,N_16357);
or U19710 (N_19710,N_15827,N_17682);
or U19711 (N_19711,N_16376,N_17070);
and U19712 (N_19712,N_18138,N_16315);
nand U19713 (N_19713,N_18483,N_17448);
nand U19714 (N_19714,N_18002,N_18335);
nand U19715 (N_19715,N_18028,N_18324);
and U19716 (N_19716,N_17228,N_16072);
or U19717 (N_19717,N_16388,N_16710);
and U19718 (N_19718,N_18010,N_15832);
and U19719 (N_19719,N_17333,N_16834);
and U19720 (N_19720,N_17692,N_15687);
or U19721 (N_19721,N_16747,N_18403);
and U19722 (N_19722,N_18238,N_17637);
xnor U19723 (N_19723,N_17351,N_17781);
nor U19724 (N_19724,N_16230,N_17002);
or U19725 (N_19725,N_15771,N_16914);
nor U19726 (N_19726,N_17541,N_15893);
nand U19727 (N_19727,N_15899,N_17193);
or U19728 (N_19728,N_16694,N_17117);
nor U19729 (N_19729,N_17291,N_18601);
nor U19730 (N_19730,N_16318,N_16988);
nor U19731 (N_19731,N_16091,N_18217);
or U19732 (N_19732,N_18499,N_15897);
nand U19733 (N_19733,N_15830,N_16868);
xnor U19734 (N_19734,N_16938,N_16900);
nand U19735 (N_19735,N_17143,N_17232);
and U19736 (N_19736,N_18080,N_18307);
nand U19737 (N_19737,N_18223,N_17832);
or U19738 (N_19738,N_17900,N_15922);
nand U19739 (N_19739,N_16687,N_16703);
nand U19740 (N_19740,N_17364,N_18159);
or U19741 (N_19741,N_16807,N_16055);
nand U19742 (N_19742,N_17936,N_15987);
nand U19743 (N_19743,N_18156,N_16283);
xnor U19744 (N_19744,N_18641,N_18046);
or U19745 (N_19745,N_18029,N_17354);
nor U19746 (N_19746,N_15780,N_16293);
nand U19747 (N_19747,N_17155,N_16154);
and U19748 (N_19748,N_18117,N_18273);
and U19749 (N_19749,N_17300,N_17749);
xnor U19750 (N_19750,N_16127,N_17131);
nor U19751 (N_19751,N_18110,N_18343);
or U19752 (N_19752,N_18701,N_17555);
nand U19753 (N_19753,N_16884,N_18041);
and U19754 (N_19754,N_18264,N_16079);
nor U19755 (N_19755,N_16398,N_17150);
nor U19756 (N_19756,N_17367,N_16853);
or U19757 (N_19757,N_15853,N_16512);
nor U19758 (N_19758,N_18198,N_16014);
and U19759 (N_19759,N_16876,N_17791);
nand U19760 (N_19760,N_17334,N_18193);
or U19761 (N_19761,N_17889,N_18207);
or U19762 (N_19762,N_17546,N_15628);
or U19763 (N_19763,N_16556,N_17140);
nor U19764 (N_19764,N_15672,N_17733);
nor U19765 (N_19765,N_16523,N_16567);
or U19766 (N_19766,N_18304,N_18622);
nor U19767 (N_19767,N_18395,N_16381);
nand U19768 (N_19768,N_16158,N_16647);
nor U19769 (N_19769,N_18134,N_16492);
or U19770 (N_19770,N_16559,N_18186);
nand U19771 (N_19771,N_17082,N_16709);
or U19772 (N_19772,N_16289,N_18085);
or U19773 (N_19773,N_16412,N_17984);
or U19774 (N_19774,N_16999,N_17488);
nand U19775 (N_19775,N_15701,N_15971);
nand U19776 (N_19776,N_16372,N_18294);
xnor U19777 (N_19777,N_18204,N_17933);
and U19778 (N_19778,N_17268,N_16491);
nor U19779 (N_19779,N_17287,N_18102);
xnor U19780 (N_19780,N_18081,N_17424);
nor U19781 (N_19781,N_16341,N_17212);
nor U19782 (N_19782,N_15645,N_15760);
or U19783 (N_19783,N_17279,N_17235);
and U19784 (N_19784,N_16753,N_16676);
and U19785 (N_19785,N_17951,N_15755);
nor U19786 (N_19786,N_17119,N_16558);
nand U19787 (N_19787,N_16295,N_18392);
and U19788 (N_19788,N_16074,N_18423);
xnor U19789 (N_19789,N_17510,N_17621);
and U19790 (N_19790,N_18603,N_18096);
nor U19791 (N_19791,N_17852,N_15966);
nand U19792 (N_19792,N_17395,N_16783);
or U19793 (N_19793,N_18593,N_15868);
and U19794 (N_19794,N_16488,N_16426);
xor U19795 (N_19795,N_17528,N_17811);
and U19796 (N_19796,N_17074,N_16287);
nor U19797 (N_19797,N_18100,N_17384);
nand U19798 (N_19798,N_16508,N_15789);
and U19799 (N_19799,N_18244,N_16734);
nand U19800 (N_19800,N_17826,N_16852);
xor U19801 (N_19801,N_17386,N_16881);
or U19802 (N_19802,N_17498,N_17496);
or U19803 (N_19803,N_16812,N_15872);
and U19804 (N_19804,N_18692,N_18216);
xor U19805 (N_19805,N_16422,N_18715);
nor U19806 (N_19806,N_18125,N_18415);
nand U19807 (N_19807,N_17085,N_17012);
and U19808 (N_19808,N_16790,N_16960);
nor U19809 (N_19809,N_17141,N_16067);
and U19810 (N_19810,N_18557,N_16563);
xor U19811 (N_19811,N_17871,N_17625);
nor U19812 (N_19812,N_16064,N_16006);
xor U19813 (N_19813,N_18533,N_16817);
nor U19814 (N_19814,N_16277,N_16966);
and U19815 (N_19815,N_16984,N_16385);
nand U19816 (N_19816,N_16051,N_15647);
or U19817 (N_19817,N_16815,N_18646);
nor U19818 (N_19818,N_17022,N_17738);
or U19819 (N_19819,N_17713,N_16832);
and U19820 (N_19820,N_15901,N_17401);
or U19821 (N_19821,N_16971,N_18014);
and U19822 (N_19822,N_16857,N_17773);
nor U19823 (N_19823,N_17255,N_17680);
and U19824 (N_19824,N_16408,N_15774);
or U19825 (N_19825,N_15959,N_17475);
nand U19826 (N_19826,N_17694,N_17731);
nand U19827 (N_19827,N_17380,N_16184);
xnor U19828 (N_19828,N_18013,N_16454);
nor U19829 (N_19829,N_16918,N_17575);
and U19830 (N_19830,N_16650,N_16594);
nand U19831 (N_19831,N_18582,N_15828);
or U19832 (N_19832,N_17502,N_17183);
or U19833 (N_19833,N_17643,N_16085);
nand U19834 (N_19834,N_17492,N_16888);
or U19835 (N_19835,N_17966,N_16519);
nor U19836 (N_19836,N_16883,N_15689);
and U19837 (N_19837,N_15928,N_16140);
and U19838 (N_19838,N_17925,N_17530);
nor U19839 (N_19839,N_17638,N_17560);
nand U19840 (N_19840,N_15826,N_16542);
and U19841 (N_19841,N_18689,N_15790);
and U19842 (N_19842,N_16351,N_16774);
nor U19843 (N_19843,N_17845,N_17820);
nand U19844 (N_19844,N_15715,N_17542);
nor U19845 (N_19845,N_17282,N_16981);
nor U19846 (N_19846,N_15794,N_15992);
and U19847 (N_19847,N_17515,N_15749);
nor U19848 (N_19848,N_16036,N_18501);
nand U19849 (N_19849,N_16222,N_18045);
or U19850 (N_19850,N_16157,N_18221);
nand U19851 (N_19851,N_17651,N_17827);
nand U19852 (N_19852,N_18463,N_15727);
nor U19853 (N_19853,N_17754,N_18104);
nand U19854 (N_19854,N_18731,N_18268);
or U19855 (N_19855,N_16808,N_16321);
and U19856 (N_19856,N_16513,N_16117);
or U19857 (N_19857,N_18735,N_18720);
nor U19858 (N_19858,N_16407,N_17931);
nand U19859 (N_19859,N_17774,N_17816);
nor U19860 (N_19860,N_16012,N_18676);
or U19861 (N_19861,N_16903,N_18469);
nor U19862 (N_19862,N_17246,N_17110);
nand U19863 (N_19863,N_17136,N_17003);
nand U19864 (N_19864,N_15954,N_16173);
nand U19865 (N_19865,N_15858,N_16054);
nor U19866 (N_19866,N_17553,N_15914);
or U19867 (N_19867,N_18722,N_16675);
or U19868 (N_19868,N_16367,N_18667);
nor U19869 (N_19869,N_17381,N_16575);
nor U19870 (N_19870,N_16693,N_18513);
nand U19871 (N_19871,N_18290,N_17905);
nand U19872 (N_19872,N_17906,N_17506);
nand U19873 (N_19873,N_16237,N_16595);
and U19874 (N_19874,N_16997,N_18555);
and U19875 (N_19875,N_17758,N_18074);
nor U19876 (N_19876,N_16193,N_16094);
or U19877 (N_19877,N_17618,N_16546);
and U19878 (N_19878,N_16923,N_16056);
nand U19879 (N_19879,N_17743,N_17967);
nand U19880 (N_19880,N_17756,N_16956);
nor U19881 (N_19881,N_17115,N_17032);
nand U19882 (N_19882,N_16770,N_18475);
and U19883 (N_19883,N_16968,N_18643);
nand U19884 (N_19884,N_15707,N_16532);
nand U19885 (N_19885,N_18235,N_16905);
nand U19886 (N_19886,N_17755,N_18150);
and U19887 (N_19887,N_17408,N_16970);
xnor U19888 (N_19888,N_18003,N_17877);
nand U19889 (N_19889,N_18246,N_15865);
and U19890 (N_19890,N_17480,N_16631);
or U19891 (N_19891,N_17898,N_15818);
or U19892 (N_19892,N_18473,N_17661);
nor U19893 (N_19893,N_15652,N_16030);
and U19894 (N_19894,N_16998,N_17518);
or U19895 (N_19895,N_15735,N_16349);
or U19896 (N_19896,N_16440,N_17972);
xor U19897 (N_19897,N_18621,N_16472);
xor U19898 (N_19898,N_16305,N_17582);
and U19899 (N_19899,N_17185,N_16021);
xnor U19900 (N_19900,N_18461,N_18378);
or U19901 (N_19901,N_15680,N_18241);
nand U19902 (N_19902,N_16028,N_17414);
xor U19903 (N_19903,N_15970,N_17358);
xor U19904 (N_19904,N_17190,N_16459);
nand U19905 (N_19905,N_17284,N_16992);
nor U19906 (N_19906,N_17725,N_15836);
xor U19907 (N_19907,N_17536,N_18409);
or U19908 (N_19908,N_16061,N_17461);
nor U19909 (N_19909,N_17376,N_16899);
or U19910 (N_19910,N_16469,N_18564);
and U19911 (N_19911,N_17659,N_15949);
and U19912 (N_19912,N_16156,N_16286);
and U19913 (N_19913,N_18137,N_18505);
nand U19914 (N_19914,N_16544,N_18550);
nand U19915 (N_19915,N_18744,N_17588);
nand U19916 (N_19916,N_16867,N_17262);
and U19917 (N_19917,N_17449,N_17142);
nor U19918 (N_19918,N_15988,N_16428);
xor U19919 (N_19919,N_16060,N_17607);
nor U19920 (N_19920,N_17375,N_15894);
nand U19921 (N_19921,N_18371,N_18517);
or U19922 (N_19922,N_16928,N_18437);
or U19923 (N_19923,N_17860,N_17797);
or U19924 (N_19924,N_18704,N_17269);
xnor U19925 (N_19925,N_16217,N_16009);
nor U19926 (N_19926,N_16272,N_17707);
or U19927 (N_19927,N_17056,N_17584);
xor U19928 (N_19928,N_17000,N_16605);
nor U19929 (N_19929,N_16390,N_18682);
or U19930 (N_19930,N_18133,N_18649);
nand U19931 (N_19931,N_17624,N_18607);
xor U19932 (N_19932,N_17771,N_16847);
nor U19933 (N_19933,N_16540,N_18477);
xnor U19934 (N_19934,N_18620,N_17479);
or U19935 (N_19935,N_16839,N_18515);
and U19936 (N_19936,N_16735,N_18431);
and U19937 (N_19937,N_16176,N_15702);
and U19938 (N_19938,N_16674,N_17892);
nand U19939 (N_19939,N_15816,N_17214);
nand U19940 (N_19940,N_16788,N_16934);
or U19941 (N_19941,N_16652,N_17822);
and U19942 (N_19942,N_17192,N_16606);
nand U19943 (N_19943,N_18322,N_18149);
or U19944 (N_19944,N_16049,N_16865);
xnor U19945 (N_19945,N_16756,N_16190);
nand U19946 (N_19946,N_15775,N_17550);
and U19947 (N_19947,N_17292,N_17387);
nand U19948 (N_19948,N_17729,N_16104);
nor U19949 (N_19949,N_17087,N_16761);
or U19950 (N_19950,N_17203,N_16214);
or U19951 (N_19951,N_18389,N_17862);
or U19952 (N_19952,N_15962,N_18480);
nand U19953 (N_19953,N_17446,N_16232);
nor U19954 (N_19954,N_17880,N_16683);
xnor U19955 (N_19955,N_16760,N_17938);
xor U19956 (N_19956,N_17163,N_16306);
nor U19957 (N_19957,N_16145,N_17999);
nand U19958 (N_19958,N_17509,N_18748);
nor U19959 (N_19959,N_17417,N_17565);
nor U19960 (N_19960,N_17636,N_16364);
and U19961 (N_19961,N_17501,N_16841);
xor U19962 (N_19962,N_18511,N_17285);
or U19963 (N_19963,N_17504,N_17924);
and U19964 (N_19964,N_18485,N_15694);
xnor U19965 (N_19965,N_17251,N_17186);
nand U19966 (N_19966,N_15896,N_16680);
and U19967 (N_19967,N_16739,N_16510);
nor U19968 (N_19968,N_16591,N_17349);
nand U19969 (N_19969,N_15937,N_17356);
or U19970 (N_19970,N_17876,N_18487);
or U19971 (N_19971,N_18251,N_18536);
nand U19972 (N_19972,N_18271,N_16449);
nand U19973 (N_19973,N_17752,N_18476);
and U19974 (N_19974,N_18608,N_16648);
nand U19975 (N_19975,N_16370,N_16902);
or U19976 (N_19976,N_17182,N_16371);
or U19977 (N_19977,N_16308,N_15936);
xor U19978 (N_19978,N_17824,N_17099);
or U19979 (N_19979,N_18233,N_17942);
and U19980 (N_19980,N_17864,N_15815);
and U19981 (N_19981,N_17808,N_18466);
and U19982 (N_19982,N_17073,N_16137);
nor U19983 (N_19983,N_17539,N_17800);
and U19984 (N_19984,N_15877,N_17608);
nand U19985 (N_19985,N_18637,N_18429);
or U19986 (N_19986,N_18103,N_17617);
or U19987 (N_19987,N_18336,N_15667);
and U19988 (N_19988,N_16167,N_15923);
or U19989 (N_19989,N_16211,N_15663);
nand U19990 (N_19990,N_18201,N_18428);
nor U19991 (N_19991,N_17124,N_16387);
or U19992 (N_19992,N_17598,N_18585);
nand U19993 (N_19993,N_16846,N_18730);
or U19994 (N_19994,N_16253,N_16261);
and U19995 (N_19995,N_16461,N_16886);
and U19996 (N_19996,N_17201,N_18652);
and U19997 (N_19997,N_17742,N_18567);
nand U19998 (N_19998,N_18237,N_18356);
xnor U19999 (N_19999,N_17818,N_17745);
and U20000 (N_20000,N_16086,N_16474);
and U20001 (N_20001,N_18060,N_16331);
nor U20002 (N_20002,N_17923,N_16438);
nand U20003 (N_20003,N_17080,N_17990);
and U20004 (N_20004,N_16827,N_17788);
nor U20005 (N_20005,N_18634,N_16912);
xor U20006 (N_20006,N_16339,N_17169);
xor U20007 (N_20007,N_16125,N_16256);
or U20008 (N_20008,N_16582,N_15718);
nor U20009 (N_20009,N_18663,N_17957);
or U20010 (N_20010,N_16875,N_16495);
nand U20011 (N_20011,N_17044,N_17406);
xor U20012 (N_20012,N_15861,N_17348);
and U20013 (N_20013,N_18163,N_17399);
and U20014 (N_20014,N_16645,N_18669);
xor U20015 (N_20015,N_16945,N_18592);
and U20016 (N_20016,N_17858,N_17976);
and U20017 (N_20017,N_18411,N_17236);
or U20018 (N_20018,N_17306,N_15632);
nand U20019 (N_20019,N_15976,N_16121);
nand U20020 (N_20020,N_18243,N_17711);
and U20021 (N_20021,N_15642,N_17324);
or U20022 (N_20022,N_15932,N_17265);
and U20023 (N_20023,N_15778,N_17685);
and U20024 (N_20024,N_16423,N_16392);
and U20025 (N_20025,N_17954,N_16231);
or U20026 (N_20026,N_16551,N_17856);
and U20027 (N_20027,N_17616,N_16033);
nor U20028 (N_20028,N_17079,N_17846);
and U20029 (N_20029,N_16732,N_16159);
and U20030 (N_20030,N_15903,N_17739);
nand U20031 (N_20031,N_15751,N_15714);
and U20032 (N_20032,N_16316,N_15784);
and U20033 (N_20033,N_15961,N_18436);
or U20034 (N_20034,N_16822,N_15772);
nor U20035 (N_20035,N_15820,N_17328);
and U20036 (N_20036,N_15851,N_17795);
xnor U20037 (N_20037,N_16436,N_16811);
nor U20038 (N_20038,N_16729,N_18390);
and U20039 (N_20039,N_15637,N_16048);
nand U20040 (N_20040,N_15847,N_18252);
nand U20041 (N_20041,N_17712,N_18526);
or U20042 (N_20042,N_17388,N_17296);
nand U20043 (N_20043,N_18155,N_17244);
nand U20044 (N_20044,N_18210,N_17902);
xnor U20045 (N_20045,N_16413,N_16713);
and U20046 (N_20046,N_16601,N_16401);
or U20047 (N_20047,N_17360,N_17180);
and U20048 (N_20048,N_16937,N_16448);
nor U20049 (N_20049,N_15730,N_18543);
nand U20050 (N_20050,N_17208,N_16737);
nand U20051 (N_20051,N_17778,N_17770);
or U20052 (N_20052,N_16340,N_16936);
nor U20053 (N_20053,N_16896,N_16978);
nand U20054 (N_20054,N_18554,N_17563);
and U20055 (N_20055,N_16024,N_18438);
or U20056 (N_20056,N_17344,N_16183);
nor U20057 (N_20057,N_17551,N_18055);
xnor U20058 (N_20058,N_18017,N_17347);
or U20059 (N_20059,N_16404,N_16113);
nor U20060 (N_20060,N_15683,N_16420);
and U20061 (N_20061,N_17714,N_17223);
nor U20062 (N_20062,N_17828,N_16047);
or U20063 (N_20063,N_16964,N_16517);
nand U20064 (N_20064,N_17887,N_18581);
nor U20065 (N_20065,N_17919,N_18716);
or U20066 (N_20066,N_18373,N_18391);
nor U20067 (N_20067,N_16679,N_17868);
or U20068 (N_20068,N_17151,N_17849);
nor U20069 (N_20069,N_15666,N_15724);
nand U20070 (N_20070,N_17468,N_16578);
or U20071 (N_20071,N_15763,N_15837);
xor U20072 (N_20072,N_16240,N_17034);
xnor U20073 (N_20073,N_16613,N_17666);
or U20074 (N_20074,N_18266,N_17710);
nand U20075 (N_20075,N_17076,N_17094);
or U20076 (N_20076,N_17357,N_18727);
xnor U20077 (N_20077,N_15649,N_17934);
nor U20078 (N_20078,N_18707,N_17316);
or U20079 (N_20079,N_16462,N_17290);
or U20080 (N_20080,N_17884,N_15808);
nor U20081 (N_20081,N_15849,N_16974);
or U20082 (N_20082,N_17988,N_16487);
nor U20083 (N_20083,N_17630,N_18384);
and U20084 (N_20084,N_18576,N_17127);
nor U20085 (N_20085,N_16752,N_18160);
and U20086 (N_20086,N_16704,N_18176);
and U20087 (N_20087,N_16144,N_16244);
and U20088 (N_20088,N_16043,N_17620);
or U20089 (N_20089,N_16762,N_15948);
xor U20090 (N_20090,N_18619,N_16199);
or U20091 (N_20091,N_16105,N_17370);
or U20092 (N_20092,N_18678,N_17135);
or U20093 (N_20093,N_18187,N_17983);
nor U20094 (N_20094,N_16083,N_17407);
nor U20095 (N_20095,N_16947,N_16151);
or U20096 (N_20096,N_18741,N_18018);
or U20097 (N_20097,N_18069,N_17790);
nor U20098 (N_20098,N_18118,N_17361);
or U20099 (N_20099,N_18280,N_18067);
nor U20100 (N_20100,N_18089,N_15904);
and U20101 (N_20101,N_16889,N_17126);
nand U20102 (N_20102,N_16068,N_17396);
nor U20103 (N_20103,N_18333,N_17945);
and U20104 (N_20104,N_16891,N_17195);
nor U20105 (N_20105,N_16333,N_17041);
or U20106 (N_20106,N_16571,N_18095);
or U20107 (N_20107,N_17466,N_17061);
nor U20108 (N_20108,N_18645,N_17969);
nor U20109 (N_20109,N_18679,N_17596);
nand U20110 (N_20110,N_18004,N_15810);
nand U20111 (N_20111,N_17450,N_17033);
and U20112 (N_20112,N_16623,N_16098);
or U20113 (N_20113,N_16236,N_18489);
xnor U20114 (N_20114,N_18615,N_17460);
or U20115 (N_20115,N_15766,N_18482);
nand U20116 (N_20116,N_15884,N_17019);
or U20117 (N_20117,N_18083,N_17051);
nand U20118 (N_20118,N_17021,N_17668);
nor U20119 (N_20119,N_18484,N_18164);
nand U20120 (N_20120,N_16175,N_15762);
nand U20121 (N_20121,N_16785,N_16539);
nand U20122 (N_20122,N_17644,N_16719);
nor U20123 (N_20123,N_17345,N_18425);
and U20124 (N_20124,N_17913,N_16825);
nor U20125 (N_20125,N_18675,N_18128);
nor U20126 (N_20126,N_16131,N_16941);
nand U20127 (N_20127,N_16282,N_16431);
and U20128 (N_20128,N_17499,N_17580);
nand U20129 (N_20129,N_15833,N_17874);
xor U20130 (N_20130,N_18090,N_18348);
xnor U20131 (N_20131,N_17452,N_16496);
nand U20132 (N_20132,N_18404,N_15654);
or U20133 (N_20133,N_17177,N_18009);
nand U20134 (N_20134,N_16465,N_16628);
nor U20135 (N_20135,N_18174,N_15676);
nor U20136 (N_20136,N_18613,N_16258);
nand U20137 (N_20137,N_15813,N_16248);
nand U20138 (N_20138,N_16445,N_16359);
and U20139 (N_20139,N_16265,N_18109);
and U20140 (N_20140,N_15765,N_17987);
nand U20141 (N_20141,N_15747,N_18478);
or U20142 (N_20142,N_16897,N_16898);
or U20143 (N_20143,N_17318,N_18093);
and U20144 (N_20144,N_16789,N_16095);
nor U20145 (N_20145,N_18558,N_18105);
or U20146 (N_20146,N_17914,N_17579);
or U20147 (N_20147,N_17483,N_16663);
nand U20148 (N_20148,N_15805,N_17863);
nor U20149 (N_20149,N_16298,N_16229);
nand U20150 (N_20150,N_17814,N_15889);
or U20151 (N_20151,N_15703,N_16489);
or U20152 (N_20152,N_17055,N_16179);
or U20153 (N_20153,N_17331,N_18143);
nor U20154 (N_20154,N_15646,N_17350);
nand U20155 (N_20155,N_16820,N_18434);
or U20156 (N_20156,N_16731,N_16026);
nor U20157 (N_20157,N_16225,N_17093);
xnor U20158 (N_20158,N_18445,N_17980);
and U20159 (N_20159,N_16767,N_18115);
or U20160 (N_20160,N_17794,N_18019);
or U20161 (N_20161,N_17104,N_17786);
nand U20162 (N_20162,N_16636,N_15758);
and U20163 (N_20163,N_18405,N_15943);
nor U20164 (N_20164,N_17059,N_16324);
or U20165 (N_20165,N_16347,N_16442);
or U20166 (N_20166,N_16577,N_17024);
nand U20167 (N_20167,N_15651,N_18605);
nor U20168 (N_20168,N_17996,N_18522);
nor U20169 (N_20169,N_17359,N_17677);
and U20170 (N_20170,N_18560,N_16441);
and U20171 (N_20171,N_16627,N_16264);
nand U20172 (N_20172,N_18563,N_18745);
and U20173 (N_20173,N_16473,N_16716);
and U20174 (N_20174,N_16656,N_18665);
nor U20175 (N_20175,N_18539,N_16574);
nand U20176 (N_20176,N_15644,N_17476);
nand U20177 (N_20177,N_17222,N_17935);
and U20178 (N_20178,N_15629,N_16833);
and U20179 (N_20179,N_16302,N_16525);
nor U20180 (N_20180,N_15648,N_18657);
and U20181 (N_20181,N_16781,N_17308);
xnor U20182 (N_20182,N_17759,N_16317);
nand U20183 (N_20183,N_18057,N_18427);
or U20184 (N_20184,N_17402,N_17405);
nand U20185 (N_20185,N_17570,N_17218);
or U20186 (N_20186,N_17322,N_17026);
nor U20187 (N_20187,N_18524,N_17007);
nor U20188 (N_20188,N_18656,N_17122);
nand U20189 (N_20189,N_17352,N_17853);
nor U20190 (N_20190,N_17309,N_18508);
xor U20191 (N_20191,N_17411,N_18639);
nor U20192 (N_20192,N_16751,N_18279);
or U20193 (N_20193,N_16403,N_17968);
nor U20194 (N_20194,N_16736,N_16931);
and U20195 (N_20195,N_17259,N_16475);
nor U20196 (N_20196,N_17412,N_16123);
nor U20197 (N_20197,N_16266,N_16022);
nand U20198 (N_20198,N_16738,N_18586);
or U20199 (N_20199,N_16273,N_18462);
or U20200 (N_20200,N_16271,N_16274);
or U20201 (N_20201,N_17084,N_18287);
or U20202 (N_20202,N_15864,N_16844);
or U20203 (N_20203,N_16633,N_16717);
nor U20204 (N_20204,N_18468,N_17549);
xnor U20205 (N_20205,N_15854,N_18479);
and U20206 (N_20206,N_16063,N_17678);
nand U20207 (N_20207,N_16746,N_15838);
nand U20208 (N_20208,N_17602,N_18481);
nor U20209 (N_20209,N_17769,N_16476);
and U20210 (N_20210,N_16042,N_16110);
xnor U20211 (N_20211,N_17765,N_17336);
or U20212 (N_20212,N_16073,N_16718);
and U20213 (N_20213,N_18175,N_17017);
nand U20214 (N_20214,N_18672,N_17590);
nand U20215 (N_20215,N_16355,N_18092);
xnor U20216 (N_20216,N_16483,N_17281);
xor U20217 (N_20217,N_16826,N_18531);
xnor U20218 (N_20218,N_15677,N_16723);
xor U20219 (N_20219,N_18291,N_15979);
nor U20220 (N_20220,N_18231,N_18249);
and U20221 (N_20221,N_18439,N_15916);
nor U20222 (N_20222,N_15933,N_18635);
nand U20223 (N_20223,N_16524,N_18314);
and U20224 (N_20224,N_18086,N_18078);
nand U20225 (N_20225,N_18598,N_17585);
and U20226 (N_20226,N_16221,N_18172);
xnor U20227 (N_20227,N_16044,N_16549);
or U20228 (N_20228,N_18743,N_16725);
nand U20229 (N_20229,N_16120,N_15625);
or U20230 (N_20230,N_18087,N_18609);
and U20231 (N_20231,N_18441,N_18208);
or U20232 (N_20232,N_17960,N_16930);
or U20233 (N_20233,N_18421,N_17982);
or U20234 (N_20234,N_15716,N_16450);
and U20235 (N_20235,N_18535,N_16901);
nor U20236 (N_20236,N_18611,N_18352);
nor U20237 (N_20237,N_18346,N_17202);
and U20238 (N_20238,N_18195,N_18206);
and U20239 (N_20239,N_16764,N_15997);
or U20240 (N_20240,N_17903,N_17031);
nor U20241 (N_20241,N_17343,N_17577);
nand U20242 (N_20242,N_17138,N_17484);
and U20243 (N_20243,N_18342,N_17337);
or U20244 (N_20244,N_17748,N_17454);
xor U20245 (N_20245,N_16323,N_15951);
and U20246 (N_20246,N_15944,N_17035);
nor U20247 (N_20247,N_15668,N_16697);
nor U20248 (N_20248,N_17734,N_18464);
and U20249 (N_20249,N_17776,N_18407);
xnor U20250 (N_20250,N_15806,N_17870);
and U20251 (N_20251,N_16066,N_16210);
and U20252 (N_20252,N_17111,N_18737);
or U20253 (N_20253,N_17780,N_18126);
nor U20254 (N_20254,N_17371,N_18310);
or U20255 (N_20255,N_16932,N_16776);
nor U20256 (N_20256,N_16869,N_16246);
or U20257 (N_20257,N_15975,N_17145);
nand U20258 (N_20258,N_18503,N_16950);
nand U20259 (N_20259,N_18097,N_17875);
xor U20260 (N_20260,N_16701,N_15817);
nor U20261 (N_20261,N_15777,N_18546);
nand U20262 (N_20262,N_18283,N_17977);
and U20263 (N_20263,N_16644,N_17088);
and U20264 (N_20264,N_17393,N_17633);
or U20265 (N_20265,N_16963,N_18229);
xnor U20266 (N_20266,N_17813,N_16037);
and U20267 (N_20267,N_17199,N_18379);
nand U20268 (N_20268,N_18648,N_16566);
and U20269 (N_20269,N_16242,N_17525);
nor U20270 (N_20270,N_16777,N_17276);
nand U20271 (N_20271,N_16643,N_18442);
or U20272 (N_20272,N_17615,N_15883);
and U20273 (N_20273,N_17994,N_17191);
and U20274 (N_20274,N_16348,N_18697);
nand U20275 (N_20275,N_17018,N_18039);
and U20276 (N_20276,N_15920,N_18190);
nor U20277 (N_20277,N_16547,N_15670);
nand U20278 (N_20278,N_16607,N_16587);
nand U20279 (N_20279,N_17207,N_16262);
or U20280 (N_20280,N_18541,N_15924);
nand U20281 (N_20281,N_15906,N_16185);
and U20282 (N_20282,N_18534,N_18326);
or U20283 (N_20283,N_17072,N_16279);
nor U20284 (N_20284,N_16344,N_17325);
or U20285 (N_20285,N_17915,N_17562);
or U20286 (N_20286,N_17120,N_16379);
xor U20287 (N_20287,N_16147,N_17674);
nand U20288 (N_20288,N_17535,N_16102);
or U20289 (N_20289,N_17503,N_16943);
xnor U20290 (N_20290,N_16498,N_16845);
and U20291 (N_20291,N_17252,N_17741);
and U20292 (N_20292,N_16166,N_16568);
or U20293 (N_20293,N_17809,N_16160);
xnor U20294 (N_20294,N_17869,N_18717);
and U20295 (N_20295,N_16973,N_17664);
and U20296 (N_20296,N_17171,N_16219);
nand U20297 (N_20297,N_15829,N_18107);
or U20298 (N_20298,N_17840,N_18015);
or U20299 (N_20299,N_18452,N_18402);
and U20300 (N_20300,N_16840,N_17782);
xnor U20301 (N_20301,N_18734,N_17234);
or U20302 (N_20302,N_17693,N_16040);
or U20303 (N_20303,N_15848,N_16165);
and U20304 (N_20304,N_18255,N_18033);
nand U20305 (N_20305,N_18612,N_16632);
or U20306 (N_20306,N_18575,N_18570);
or U20307 (N_20307,N_17116,N_17540);
and U20308 (N_20308,N_18497,N_16430);
or U20309 (N_20309,N_15876,N_16579);
or U20310 (N_20310,N_15713,N_16593);
xnor U20311 (N_20311,N_18219,N_16799);
nand U20312 (N_20312,N_17075,N_17260);
xor U20313 (N_20313,N_16812,N_17374);
nor U20314 (N_20314,N_16989,N_16495);
or U20315 (N_20315,N_17661,N_18140);
and U20316 (N_20316,N_16501,N_16479);
and U20317 (N_20317,N_18380,N_16638);
nor U20318 (N_20318,N_16006,N_18748);
nor U20319 (N_20319,N_18230,N_15708);
nor U20320 (N_20320,N_17445,N_17010);
or U20321 (N_20321,N_17347,N_16894);
nand U20322 (N_20322,N_16554,N_16302);
nand U20323 (N_20323,N_16441,N_16589);
nand U20324 (N_20324,N_16532,N_18205);
xnor U20325 (N_20325,N_17051,N_17673);
or U20326 (N_20326,N_17747,N_16889);
or U20327 (N_20327,N_16050,N_16305);
or U20328 (N_20328,N_17535,N_18555);
xor U20329 (N_20329,N_17157,N_18322);
or U20330 (N_20330,N_18011,N_17870);
or U20331 (N_20331,N_17855,N_16724);
nand U20332 (N_20332,N_17095,N_16646);
or U20333 (N_20333,N_17630,N_18484);
or U20334 (N_20334,N_18533,N_18292);
and U20335 (N_20335,N_16974,N_18531);
nor U20336 (N_20336,N_15998,N_17070);
xnor U20337 (N_20337,N_17386,N_17826);
nand U20338 (N_20338,N_16094,N_16442);
xor U20339 (N_20339,N_17155,N_16294);
nand U20340 (N_20340,N_18099,N_18549);
nor U20341 (N_20341,N_18135,N_16718);
nand U20342 (N_20342,N_18431,N_16608);
and U20343 (N_20343,N_17013,N_17803);
nor U20344 (N_20344,N_16402,N_15808);
and U20345 (N_20345,N_16665,N_16148);
nor U20346 (N_20346,N_18620,N_17499);
and U20347 (N_20347,N_17452,N_17747);
xnor U20348 (N_20348,N_16344,N_16170);
nand U20349 (N_20349,N_15701,N_16861);
nand U20350 (N_20350,N_15888,N_16253);
or U20351 (N_20351,N_18540,N_18406);
nand U20352 (N_20352,N_18441,N_17804);
xnor U20353 (N_20353,N_17367,N_18557);
nand U20354 (N_20354,N_18660,N_17275);
or U20355 (N_20355,N_18694,N_18332);
and U20356 (N_20356,N_15785,N_15709);
nor U20357 (N_20357,N_17889,N_17477);
nor U20358 (N_20358,N_16442,N_15821);
and U20359 (N_20359,N_16812,N_18552);
nor U20360 (N_20360,N_18262,N_16514);
nor U20361 (N_20361,N_18122,N_18163);
or U20362 (N_20362,N_18045,N_16594);
or U20363 (N_20363,N_15988,N_16540);
or U20364 (N_20364,N_17666,N_17151);
nand U20365 (N_20365,N_18630,N_17195);
nor U20366 (N_20366,N_15984,N_16017);
nor U20367 (N_20367,N_18304,N_17185);
and U20368 (N_20368,N_17770,N_18550);
nor U20369 (N_20369,N_17588,N_16653);
and U20370 (N_20370,N_18192,N_15768);
xor U20371 (N_20371,N_15895,N_16307);
and U20372 (N_20372,N_17275,N_18240);
or U20373 (N_20373,N_17331,N_18323);
or U20374 (N_20374,N_16812,N_16185);
nand U20375 (N_20375,N_17855,N_18322);
and U20376 (N_20376,N_18454,N_17154);
xnor U20377 (N_20377,N_16228,N_18550);
or U20378 (N_20378,N_15881,N_17768);
nand U20379 (N_20379,N_15980,N_17843);
and U20380 (N_20380,N_17271,N_18232);
or U20381 (N_20381,N_18728,N_17142);
and U20382 (N_20382,N_17624,N_18233);
and U20383 (N_20383,N_17022,N_17501);
or U20384 (N_20384,N_16949,N_16353);
nor U20385 (N_20385,N_17646,N_17181);
and U20386 (N_20386,N_18592,N_18186);
and U20387 (N_20387,N_17947,N_16816);
nor U20388 (N_20388,N_17218,N_15896);
nand U20389 (N_20389,N_16023,N_17729);
nor U20390 (N_20390,N_18069,N_16198);
or U20391 (N_20391,N_17452,N_16815);
and U20392 (N_20392,N_15730,N_17599);
or U20393 (N_20393,N_18536,N_17612);
and U20394 (N_20394,N_18695,N_18665);
and U20395 (N_20395,N_16330,N_16211);
nor U20396 (N_20396,N_17425,N_18115);
nand U20397 (N_20397,N_15917,N_17828);
and U20398 (N_20398,N_17045,N_15746);
xnor U20399 (N_20399,N_17560,N_17980);
and U20400 (N_20400,N_17486,N_16901);
or U20401 (N_20401,N_18082,N_16821);
nand U20402 (N_20402,N_17178,N_18735);
and U20403 (N_20403,N_17628,N_18353);
nor U20404 (N_20404,N_18227,N_16768);
nor U20405 (N_20405,N_17945,N_15730);
nor U20406 (N_20406,N_18159,N_16973);
nor U20407 (N_20407,N_17685,N_18738);
nor U20408 (N_20408,N_18102,N_17665);
or U20409 (N_20409,N_17866,N_15790);
nor U20410 (N_20410,N_17487,N_18136);
xor U20411 (N_20411,N_16368,N_16424);
nand U20412 (N_20412,N_16721,N_16077);
and U20413 (N_20413,N_15946,N_16925);
nor U20414 (N_20414,N_17292,N_17182);
or U20415 (N_20415,N_18098,N_16741);
or U20416 (N_20416,N_18428,N_15661);
and U20417 (N_20417,N_16491,N_16946);
or U20418 (N_20418,N_15949,N_17977);
or U20419 (N_20419,N_17225,N_16949);
and U20420 (N_20420,N_18173,N_17521);
and U20421 (N_20421,N_17988,N_18292);
and U20422 (N_20422,N_17159,N_16308);
and U20423 (N_20423,N_16396,N_16940);
nand U20424 (N_20424,N_16286,N_15842);
nand U20425 (N_20425,N_17494,N_16979);
nor U20426 (N_20426,N_16559,N_16678);
nand U20427 (N_20427,N_17233,N_17536);
or U20428 (N_20428,N_18304,N_18502);
nand U20429 (N_20429,N_16981,N_16761);
nor U20430 (N_20430,N_17611,N_16611);
or U20431 (N_20431,N_18405,N_16973);
and U20432 (N_20432,N_16889,N_18509);
xor U20433 (N_20433,N_17992,N_18122);
nand U20434 (N_20434,N_17715,N_17131);
or U20435 (N_20435,N_16228,N_17712);
and U20436 (N_20436,N_17164,N_16185);
or U20437 (N_20437,N_16324,N_18456);
nor U20438 (N_20438,N_18272,N_16675);
nor U20439 (N_20439,N_15695,N_17786);
or U20440 (N_20440,N_16920,N_17368);
nor U20441 (N_20441,N_18144,N_17098);
nand U20442 (N_20442,N_17381,N_17067);
and U20443 (N_20443,N_17409,N_16813);
nor U20444 (N_20444,N_18025,N_17572);
nand U20445 (N_20445,N_18578,N_15655);
and U20446 (N_20446,N_18498,N_18617);
or U20447 (N_20447,N_16116,N_16583);
nand U20448 (N_20448,N_16543,N_16823);
or U20449 (N_20449,N_18255,N_18618);
nand U20450 (N_20450,N_17613,N_16336);
and U20451 (N_20451,N_17071,N_18199);
nand U20452 (N_20452,N_17253,N_17412);
nor U20453 (N_20453,N_17963,N_16131);
nor U20454 (N_20454,N_17791,N_15927);
or U20455 (N_20455,N_15902,N_16340);
and U20456 (N_20456,N_17181,N_17394);
xnor U20457 (N_20457,N_18718,N_17388);
xor U20458 (N_20458,N_18192,N_16384);
and U20459 (N_20459,N_17669,N_17654);
nand U20460 (N_20460,N_15708,N_16881);
nor U20461 (N_20461,N_17244,N_17547);
or U20462 (N_20462,N_17323,N_15912);
nand U20463 (N_20463,N_16474,N_16731);
xor U20464 (N_20464,N_18673,N_18236);
nor U20465 (N_20465,N_15731,N_18187);
xnor U20466 (N_20466,N_18617,N_16472);
and U20467 (N_20467,N_16520,N_16330);
and U20468 (N_20468,N_16822,N_18643);
nor U20469 (N_20469,N_18739,N_18631);
nor U20470 (N_20470,N_16634,N_15972);
or U20471 (N_20471,N_17884,N_16368);
and U20472 (N_20472,N_17498,N_16367);
nor U20473 (N_20473,N_17845,N_16775);
nor U20474 (N_20474,N_17467,N_17758);
or U20475 (N_20475,N_17920,N_16666);
and U20476 (N_20476,N_16149,N_18103);
and U20477 (N_20477,N_18149,N_15855);
or U20478 (N_20478,N_18078,N_17551);
nand U20479 (N_20479,N_17012,N_18293);
or U20480 (N_20480,N_17804,N_18165);
and U20481 (N_20481,N_17013,N_17425);
or U20482 (N_20482,N_17905,N_15641);
and U20483 (N_20483,N_17295,N_15811);
and U20484 (N_20484,N_18494,N_16627);
nor U20485 (N_20485,N_17727,N_16325);
nor U20486 (N_20486,N_18454,N_17544);
nor U20487 (N_20487,N_18256,N_17358);
and U20488 (N_20488,N_18193,N_16828);
nor U20489 (N_20489,N_17112,N_17607);
and U20490 (N_20490,N_16818,N_17688);
and U20491 (N_20491,N_18194,N_15795);
nor U20492 (N_20492,N_15672,N_18428);
or U20493 (N_20493,N_17885,N_17598);
nand U20494 (N_20494,N_17198,N_17175);
nand U20495 (N_20495,N_18254,N_16939);
nand U20496 (N_20496,N_16305,N_18713);
and U20497 (N_20497,N_17419,N_17303);
nor U20498 (N_20498,N_16047,N_15911);
nand U20499 (N_20499,N_17987,N_16627);
and U20500 (N_20500,N_16159,N_16040);
or U20501 (N_20501,N_18641,N_17890);
and U20502 (N_20502,N_16219,N_15881);
xor U20503 (N_20503,N_16158,N_16721);
nand U20504 (N_20504,N_17192,N_17281);
and U20505 (N_20505,N_16684,N_18577);
nor U20506 (N_20506,N_16127,N_16370);
and U20507 (N_20507,N_15820,N_16129);
and U20508 (N_20508,N_17864,N_17563);
and U20509 (N_20509,N_16982,N_17352);
nand U20510 (N_20510,N_17633,N_18142);
or U20511 (N_20511,N_15920,N_18284);
and U20512 (N_20512,N_16312,N_16640);
and U20513 (N_20513,N_15858,N_16234);
or U20514 (N_20514,N_18696,N_18640);
nand U20515 (N_20515,N_16706,N_18150);
and U20516 (N_20516,N_16572,N_18339);
and U20517 (N_20517,N_16298,N_16511);
nor U20518 (N_20518,N_16668,N_18518);
nor U20519 (N_20519,N_16372,N_17312);
or U20520 (N_20520,N_17574,N_16459);
xnor U20521 (N_20521,N_16969,N_18467);
xnor U20522 (N_20522,N_18162,N_16725);
and U20523 (N_20523,N_18749,N_17663);
and U20524 (N_20524,N_18414,N_18061);
nor U20525 (N_20525,N_18092,N_16963);
and U20526 (N_20526,N_17151,N_17713);
or U20527 (N_20527,N_18359,N_18477);
nand U20528 (N_20528,N_17172,N_16075);
or U20529 (N_20529,N_15927,N_16010);
or U20530 (N_20530,N_17965,N_16851);
nor U20531 (N_20531,N_17967,N_17273);
or U20532 (N_20532,N_17340,N_16907);
nor U20533 (N_20533,N_18368,N_16412);
nor U20534 (N_20534,N_17099,N_16957);
nand U20535 (N_20535,N_17337,N_17815);
and U20536 (N_20536,N_18559,N_17655);
xnor U20537 (N_20537,N_16311,N_18692);
nor U20538 (N_20538,N_16006,N_17714);
nor U20539 (N_20539,N_18153,N_15747);
xor U20540 (N_20540,N_17229,N_16775);
and U20541 (N_20541,N_18267,N_16784);
and U20542 (N_20542,N_17431,N_17453);
and U20543 (N_20543,N_15970,N_18026);
nand U20544 (N_20544,N_16095,N_18167);
or U20545 (N_20545,N_15645,N_16740);
nor U20546 (N_20546,N_17066,N_18686);
nor U20547 (N_20547,N_16004,N_17290);
and U20548 (N_20548,N_16996,N_17026);
nand U20549 (N_20549,N_18136,N_18341);
and U20550 (N_20550,N_18037,N_15715);
or U20551 (N_20551,N_15684,N_18133);
or U20552 (N_20552,N_15962,N_16754);
and U20553 (N_20553,N_18469,N_17487);
or U20554 (N_20554,N_17122,N_17996);
or U20555 (N_20555,N_17373,N_16848);
or U20556 (N_20556,N_17028,N_17834);
or U20557 (N_20557,N_17769,N_16734);
xnor U20558 (N_20558,N_17714,N_17253);
nand U20559 (N_20559,N_17044,N_17996);
nand U20560 (N_20560,N_16480,N_15884);
and U20561 (N_20561,N_16969,N_16018);
nand U20562 (N_20562,N_15742,N_18381);
or U20563 (N_20563,N_15907,N_15741);
xor U20564 (N_20564,N_16131,N_15878);
xor U20565 (N_20565,N_15661,N_15963);
or U20566 (N_20566,N_18256,N_17097);
and U20567 (N_20567,N_16265,N_16709);
nand U20568 (N_20568,N_17755,N_16902);
nor U20569 (N_20569,N_17400,N_16066);
nand U20570 (N_20570,N_18221,N_15784);
nor U20571 (N_20571,N_17745,N_17144);
and U20572 (N_20572,N_17988,N_15769);
nand U20573 (N_20573,N_16477,N_16180);
nand U20574 (N_20574,N_18314,N_16702);
nand U20575 (N_20575,N_16108,N_17222);
nor U20576 (N_20576,N_17568,N_15845);
nand U20577 (N_20577,N_16698,N_17748);
and U20578 (N_20578,N_17865,N_16066);
nand U20579 (N_20579,N_18181,N_18208);
nor U20580 (N_20580,N_18001,N_16773);
xor U20581 (N_20581,N_16675,N_18649);
and U20582 (N_20582,N_17154,N_17250);
and U20583 (N_20583,N_17515,N_15645);
or U20584 (N_20584,N_17406,N_16536);
xnor U20585 (N_20585,N_15713,N_17878);
nor U20586 (N_20586,N_16700,N_17448);
or U20587 (N_20587,N_17114,N_18411);
or U20588 (N_20588,N_16911,N_16579);
nor U20589 (N_20589,N_17830,N_16602);
nand U20590 (N_20590,N_18416,N_16271);
nand U20591 (N_20591,N_18328,N_17216);
nand U20592 (N_20592,N_17438,N_16300);
nand U20593 (N_20593,N_18578,N_17822);
xnor U20594 (N_20594,N_17312,N_18369);
nand U20595 (N_20595,N_18103,N_18703);
nand U20596 (N_20596,N_16443,N_17441);
or U20597 (N_20597,N_18323,N_16672);
or U20598 (N_20598,N_15645,N_17993);
nor U20599 (N_20599,N_17053,N_16682);
nand U20600 (N_20600,N_17995,N_15865);
or U20601 (N_20601,N_16049,N_18152);
and U20602 (N_20602,N_18095,N_16442);
nand U20603 (N_20603,N_17769,N_18468);
and U20604 (N_20604,N_16356,N_15722);
nor U20605 (N_20605,N_16053,N_17506);
and U20606 (N_20606,N_16076,N_18704);
and U20607 (N_20607,N_16069,N_18394);
nand U20608 (N_20608,N_18696,N_18121);
nor U20609 (N_20609,N_18485,N_16714);
and U20610 (N_20610,N_16481,N_16871);
nor U20611 (N_20611,N_18440,N_18004);
nor U20612 (N_20612,N_17377,N_17069);
and U20613 (N_20613,N_17044,N_17753);
or U20614 (N_20614,N_15785,N_18082);
nand U20615 (N_20615,N_18632,N_17705);
xor U20616 (N_20616,N_16943,N_15883);
nor U20617 (N_20617,N_16789,N_16312);
or U20618 (N_20618,N_15744,N_18256);
xnor U20619 (N_20619,N_18347,N_17418);
or U20620 (N_20620,N_16044,N_16020);
nand U20621 (N_20621,N_17377,N_18450);
and U20622 (N_20622,N_15680,N_17808);
or U20623 (N_20623,N_16548,N_16865);
or U20624 (N_20624,N_17193,N_17326);
nand U20625 (N_20625,N_17744,N_16434);
or U20626 (N_20626,N_17820,N_16138);
or U20627 (N_20627,N_15814,N_17314);
nor U20628 (N_20628,N_18018,N_18388);
nor U20629 (N_20629,N_15689,N_17994);
nor U20630 (N_20630,N_18088,N_17119);
or U20631 (N_20631,N_18399,N_17335);
and U20632 (N_20632,N_16718,N_15826);
or U20633 (N_20633,N_15688,N_17078);
and U20634 (N_20634,N_16710,N_18596);
or U20635 (N_20635,N_17684,N_17593);
nand U20636 (N_20636,N_17718,N_17794);
nor U20637 (N_20637,N_16867,N_18153);
nor U20638 (N_20638,N_18373,N_16069);
and U20639 (N_20639,N_17362,N_15880);
or U20640 (N_20640,N_16419,N_18418);
nor U20641 (N_20641,N_18212,N_18118);
or U20642 (N_20642,N_17644,N_18084);
and U20643 (N_20643,N_18401,N_17463);
nor U20644 (N_20644,N_17908,N_17565);
or U20645 (N_20645,N_18124,N_17301);
or U20646 (N_20646,N_18222,N_17462);
and U20647 (N_20647,N_18674,N_18508);
nor U20648 (N_20648,N_15751,N_17439);
or U20649 (N_20649,N_16950,N_17048);
nor U20650 (N_20650,N_17832,N_17780);
nand U20651 (N_20651,N_16764,N_17420);
nor U20652 (N_20652,N_16343,N_17492);
and U20653 (N_20653,N_16982,N_17152);
or U20654 (N_20654,N_16400,N_16299);
nand U20655 (N_20655,N_16598,N_18157);
nand U20656 (N_20656,N_18696,N_17113);
nand U20657 (N_20657,N_16543,N_18463);
or U20658 (N_20658,N_16744,N_18473);
or U20659 (N_20659,N_16785,N_18244);
nor U20660 (N_20660,N_16668,N_18020);
or U20661 (N_20661,N_15719,N_16456);
and U20662 (N_20662,N_18344,N_16878);
and U20663 (N_20663,N_17657,N_16494);
and U20664 (N_20664,N_16868,N_16168);
nand U20665 (N_20665,N_18707,N_16731);
nand U20666 (N_20666,N_16372,N_17993);
xor U20667 (N_20667,N_17348,N_18560);
nor U20668 (N_20668,N_16741,N_15900);
or U20669 (N_20669,N_17337,N_17697);
or U20670 (N_20670,N_18504,N_17318);
xnor U20671 (N_20671,N_17196,N_17821);
and U20672 (N_20672,N_17023,N_16466);
or U20673 (N_20673,N_17596,N_16435);
xnor U20674 (N_20674,N_16817,N_17871);
xnor U20675 (N_20675,N_17544,N_17454);
or U20676 (N_20676,N_18462,N_17061);
and U20677 (N_20677,N_18518,N_18459);
and U20678 (N_20678,N_16905,N_17157);
nand U20679 (N_20679,N_17803,N_16457);
xnor U20680 (N_20680,N_15781,N_17354);
or U20681 (N_20681,N_17555,N_18266);
nor U20682 (N_20682,N_16219,N_18415);
and U20683 (N_20683,N_18302,N_17875);
nand U20684 (N_20684,N_16127,N_18717);
nor U20685 (N_20685,N_18638,N_17008);
or U20686 (N_20686,N_17625,N_15984);
or U20687 (N_20687,N_15969,N_16244);
or U20688 (N_20688,N_16726,N_16136);
nor U20689 (N_20689,N_17770,N_16776);
nand U20690 (N_20690,N_18383,N_17035);
nor U20691 (N_20691,N_17852,N_17548);
and U20692 (N_20692,N_16259,N_16846);
xnor U20693 (N_20693,N_16108,N_17880);
nor U20694 (N_20694,N_17773,N_18280);
xnor U20695 (N_20695,N_17816,N_17312);
or U20696 (N_20696,N_17371,N_17014);
nand U20697 (N_20697,N_15640,N_16386);
xnor U20698 (N_20698,N_17036,N_17655);
and U20699 (N_20699,N_18719,N_15634);
and U20700 (N_20700,N_16908,N_17840);
xor U20701 (N_20701,N_16967,N_16969);
nand U20702 (N_20702,N_18284,N_17218);
xor U20703 (N_20703,N_18678,N_17885);
nand U20704 (N_20704,N_15967,N_16553);
or U20705 (N_20705,N_16673,N_16928);
or U20706 (N_20706,N_17104,N_16031);
or U20707 (N_20707,N_16498,N_16830);
nor U20708 (N_20708,N_15928,N_16725);
nor U20709 (N_20709,N_16984,N_17785);
nor U20710 (N_20710,N_15907,N_16537);
or U20711 (N_20711,N_17864,N_18277);
or U20712 (N_20712,N_16876,N_17669);
nor U20713 (N_20713,N_15736,N_16275);
xnor U20714 (N_20714,N_17209,N_16649);
nand U20715 (N_20715,N_16630,N_18603);
or U20716 (N_20716,N_16303,N_17431);
or U20717 (N_20717,N_16662,N_17160);
or U20718 (N_20718,N_16853,N_16996);
nand U20719 (N_20719,N_18003,N_16852);
or U20720 (N_20720,N_17171,N_18054);
or U20721 (N_20721,N_18270,N_17239);
or U20722 (N_20722,N_17335,N_17955);
nand U20723 (N_20723,N_15625,N_18682);
nand U20724 (N_20724,N_17427,N_16007);
and U20725 (N_20725,N_17071,N_18083);
nor U20726 (N_20726,N_16265,N_17781);
nand U20727 (N_20727,N_17349,N_18640);
nand U20728 (N_20728,N_18242,N_18636);
and U20729 (N_20729,N_18049,N_15961);
nor U20730 (N_20730,N_16026,N_17448);
or U20731 (N_20731,N_15642,N_17617);
xnor U20732 (N_20732,N_18263,N_16055);
xor U20733 (N_20733,N_15974,N_16092);
and U20734 (N_20734,N_15659,N_16277);
and U20735 (N_20735,N_18348,N_16042);
nand U20736 (N_20736,N_17617,N_17581);
nor U20737 (N_20737,N_16873,N_15891);
and U20738 (N_20738,N_18390,N_18255);
and U20739 (N_20739,N_16408,N_18267);
nor U20740 (N_20740,N_17158,N_18296);
nor U20741 (N_20741,N_17646,N_16950);
nand U20742 (N_20742,N_17491,N_16549);
and U20743 (N_20743,N_16086,N_17007);
or U20744 (N_20744,N_17129,N_17572);
or U20745 (N_20745,N_16109,N_16376);
nor U20746 (N_20746,N_16301,N_17927);
nand U20747 (N_20747,N_16150,N_16388);
nor U20748 (N_20748,N_18700,N_16315);
and U20749 (N_20749,N_17034,N_15918);
nor U20750 (N_20750,N_16623,N_16502);
nand U20751 (N_20751,N_16387,N_17438);
nor U20752 (N_20752,N_18110,N_17624);
or U20753 (N_20753,N_18217,N_16510);
and U20754 (N_20754,N_16059,N_18567);
nand U20755 (N_20755,N_17868,N_16822);
and U20756 (N_20756,N_18324,N_18377);
and U20757 (N_20757,N_18506,N_16450);
and U20758 (N_20758,N_17886,N_17345);
and U20759 (N_20759,N_18243,N_15932);
nand U20760 (N_20760,N_16746,N_16108);
and U20761 (N_20761,N_15810,N_18121);
nand U20762 (N_20762,N_16819,N_17794);
nor U20763 (N_20763,N_18137,N_15852);
and U20764 (N_20764,N_18195,N_16164);
nand U20765 (N_20765,N_16973,N_17314);
nand U20766 (N_20766,N_16146,N_17923);
nand U20767 (N_20767,N_18411,N_16503);
nand U20768 (N_20768,N_16618,N_15969);
or U20769 (N_20769,N_17518,N_18708);
and U20770 (N_20770,N_16692,N_18071);
nand U20771 (N_20771,N_17571,N_16956);
or U20772 (N_20772,N_17732,N_16182);
nand U20773 (N_20773,N_16618,N_16685);
and U20774 (N_20774,N_17733,N_17423);
or U20775 (N_20775,N_17086,N_17769);
and U20776 (N_20776,N_16444,N_16567);
nand U20777 (N_20777,N_16875,N_17051);
or U20778 (N_20778,N_15999,N_16959);
or U20779 (N_20779,N_17727,N_16735);
nor U20780 (N_20780,N_18544,N_16968);
and U20781 (N_20781,N_18289,N_15837);
or U20782 (N_20782,N_18039,N_15793);
nand U20783 (N_20783,N_18100,N_16576);
xnor U20784 (N_20784,N_16686,N_16274);
and U20785 (N_20785,N_18580,N_17624);
nand U20786 (N_20786,N_16229,N_15777);
xnor U20787 (N_20787,N_16470,N_16996);
nand U20788 (N_20788,N_16062,N_16325);
nor U20789 (N_20789,N_18540,N_17123);
nand U20790 (N_20790,N_17180,N_18633);
and U20791 (N_20791,N_16698,N_17581);
nor U20792 (N_20792,N_17678,N_17475);
or U20793 (N_20793,N_15889,N_16976);
or U20794 (N_20794,N_18738,N_18109);
and U20795 (N_20795,N_16745,N_18068);
nor U20796 (N_20796,N_17720,N_18265);
or U20797 (N_20797,N_16947,N_17446);
xnor U20798 (N_20798,N_18540,N_16317);
nor U20799 (N_20799,N_17573,N_17342);
nand U20800 (N_20800,N_18523,N_18468);
xor U20801 (N_20801,N_18593,N_16586);
or U20802 (N_20802,N_16155,N_16202);
or U20803 (N_20803,N_16226,N_17439);
and U20804 (N_20804,N_17243,N_16082);
nand U20805 (N_20805,N_16173,N_16485);
or U20806 (N_20806,N_15758,N_17476);
and U20807 (N_20807,N_17942,N_18044);
or U20808 (N_20808,N_18522,N_17522);
xnor U20809 (N_20809,N_17149,N_15806);
nor U20810 (N_20810,N_15803,N_16821);
and U20811 (N_20811,N_18732,N_15660);
nand U20812 (N_20812,N_17306,N_16366);
and U20813 (N_20813,N_16254,N_17306);
and U20814 (N_20814,N_15801,N_17968);
nor U20815 (N_20815,N_16556,N_17384);
and U20816 (N_20816,N_18699,N_15787);
or U20817 (N_20817,N_17611,N_18607);
and U20818 (N_20818,N_17999,N_17334);
nor U20819 (N_20819,N_16540,N_17082);
and U20820 (N_20820,N_17709,N_16060);
nor U20821 (N_20821,N_16535,N_16689);
or U20822 (N_20822,N_16477,N_17712);
nor U20823 (N_20823,N_18365,N_18029);
nor U20824 (N_20824,N_16860,N_18484);
nor U20825 (N_20825,N_17602,N_17098);
and U20826 (N_20826,N_15857,N_18477);
xnor U20827 (N_20827,N_18227,N_16644);
xor U20828 (N_20828,N_17944,N_17879);
and U20829 (N_20829,N_17629,N_17631);
nand U20830 (N_20830,N_16274,N_16084);
or U20831 (N_20831,N_15771,N_18273);
and U20832 (N_20832,N_18699,N_17293);
nand U20833 (N_20833,N_17115,N_16362);
nor U20834 (N_20834,N_18344,N_17124);
nor U20835 (N_20835,N_18536,N_16984);
and U20836 (N_20836,N_17072,N_18047);
or U20837 (N_20837,N_16780,N_15750);
nor U20838 (N_20838,N_18438,N_16427);
nand U20839 (N_20839,N_18395,N_16848);
nor U20840 (N_20840,N_16353,N_15950);
or U20841 (N_20841,N_16700,N_15948);
or U20842 (N_20842,N_18117,N_17543);
or U20843 (N_20843,N_16021,N_17456);
nor U20844 (N_20844,N_17562,N_18099);
and U20845 (N_20845,N_16589,N_15639);
nand U20846 (N_20846,N_16281,N_17950);
and U20847 (N_20847,N_16129,N_18546);
or U20848 (N_20848,N_18391,N_17844);
nand U20849 (N_20849,N_17304,N_16400);
nand U20850 (N_20850,N_16910,N_16951);
nand U20851 (N_20851,N_16065,N_17738);
xnor U20852 (N_20852,N_18016,N_18485);
or U20853 (N_20853,N_16685,N_15806);
or U20854 (N_20854,N_15921,N_18660);
and U20855 (N_20855,N_17446,N_15731);
nor U20856 (N_20856,N_16358,N_17823);
nand U20857 (N_20857,N_17437,N_17280);
nand U20858 (N_20858,N_16717,N_16684);
nand U20859 (N_20859,N_15686,N_16991);
nor U20860 (N_20860,N_15678,N_16819);
or U20861 (N_20861,N_17658,N_16205);
nand U20862 (N_20862,N_17460,N_17577);
nand U20863 (N_20863,N_18616,N_17932);
or U20864 (N_20864,N_18634,N_17681);
nand U20865 (N_20865,N_15705,N_16642);
nor U20866 (N_20866,N_16054,N_17144);
or U20867 (N_20867,N_17380,N_18389);
or U20868 (N_20868,N_16969,N_16742);
xnor U20869 (N_20869,N_16106,N_17748);
nor U20870 (N_20870,N_16113,N_15718);
and U20871 (N_20871,N_17579,N_16588);
or U20872 (N_20872,N_18270,N_15928);
xnor U20873 (N_20873,N_18417,N_18648);
nand U20874 (N_20874,N_17922,N_16362);
nand U20875 (N_20875,N_16553,N_16708);
and U20876 (N_20876,N_15702,N_18276);
or U20877 (N_20877,N_18640,N_16165);
nand U20878 (N_20878,N_16720,N_16957);
or U20879 (N_20879,N_18598,N_18650);
nand U20880 (N_20880,N_16998,N_18030);
and U20881 (N_20881,N_16305,N_17588);
and U20882 (N_20882,N_17599,N_16188);
xor U20883 (N_20883,N_18329,N_16845);
and U20884 (N_20884,N_15837,N_18163);
and U20885 (N_20885,N_17518,N_18050);
or U20886 (N_20886,N_16660,N_15973);
and U20887 (N_20887,N_17320,N_17738);
nand U20888 (N_20888,N_16771,N_18713);
nor U20889 (N_20889,N_16357,N_17034);
or U20890 (N_20890,N_16337,N_16100);
and U20891 (N_20891,N_18095,N_18029);
nand U20892 (N_20892,N_18478,N_18559);
and U20893 (N_20893,N_17901,N_18163);
and U20894 (N_20894,N_17163,N_17979);
and U20895 (N_20895,N_17494,N_16255);
nor U20896 (N_20896,N_17874,N_17312);
or U20897 (N_20897,N_18051,N_17912);
nand U20898 (N_20898,N_17557,N_17126);
nand U20899 (N_20899,N_16552,N_18287);
nor U20900 (N_20900,N_15710,N_18289);
and U20901 (N_20901,N_15863,N_16477);
nand U20902 (N_20902,N_18735,N_17115);
nor U20903 (N_20903,N_18527,N_17070);
xnor U20904 (N_20904,N_17070,N_16804);
nand U20905 (N_20905,N_15699,N_17951);
xor U20906 (N_20906,N_17823,N_17878);
and U20907 (N_20907,N_18117,N_18351);
nand U20908 (N_20908,N_18151,N_16753);
and U20909 (N_20909,N_18651,N_16202);
nor U20910 (N_20910,N_16719,N_16192);
and U20911 (N_20911,N_15652,N_17562);
or U20912 (N_20912,N_15998,N_16288);
nor U20913 (N_20913,N_16437,N_16127);
xor U20914 (N_20914,N_16665,N_17232);
or U20915 (N_20915,N_18190,N_15642);
nor U20916 (N_20916,N_17606,N_16394);
and U20917 (N_20917,N_18528,N_16855);
and U20918 (N_20918,N_16011,N_16436);
nand U20919 (N_20919,N_16506,N_16966);
xnor U20920 (N_20920,N_15970,N_17491);
or U20921 (N_20921,N_16968,N_16298);
and U20922 (N_20922,N_18550,N_16139);
nand U20923 (N_20923,N_16116,N_17881);
xor U20924 (N_20924,N_17723,N_17830);
nand U20925 (N_20925,N_18021,N_16329);
nor U20926 (N_20926,N_16832,N_16501);
and U20927 (N_20927,N_17708,N_18300);
nor U20928 (N_20928,N_16665,N_17287);
nand U20929 (N_20929,N_16692,N_16000);
and U20930 (N_20930,N_17380,N_18310);
xnor U20931 (N_20931,N_17141,N_18200);
or U20932 (N_20932,N_17045,N_18588);
and U20933 (N_20933,N_16104,N_16688);
and U20934 (N_20934,N_17477,N_18230);
and U20935 (N_20935,N_18344,N_18098);
and U20936 (N_20936,N_15652,N_17276);
nor U20937 (N_20937,N_16584,N_18429);
nand U20938 (N_20938,N_16916,N_18183);
and U20939 (N_20939,N_16009,N_16406);
or U20940 (N_20940,N_16439,N_18514);
and U20941 (N_20941,N_17352,N_17845);
and U20942 (N_20942,N_15918,N_17329);
or U20943 (N_20943,N_16021,N_16026);
or U20944 (N_20944,N_18212,N_16088);
or U20945 (N_20945,N_17785,N_17772);
and U20946 (N_20946,N_18628,N_17647);
or U20947 (N_20947,N_17062,N_16958);
nand U20948 (N_20948,N_18593,N_15875);
nor U20949 (N_20949,N_18071,N_15858);
nand U20950 (N_20950,N_16242,N_18231);
and U20951 (N_20951,N_18041,N_17132);
or U20952 (N_20952,N_16889,N_16723);
nand U20953 (N_20953,N_18378,N_18126);
nor U20954 (N_20954,N_16872,N_18079);
nor U20955 (N_20955,N_16029,N_15794);
nor U20956 (N_20956,N_18342,N_16374);
and U20957 (N_20957,N_16148,N_16816);
nand U20958 (N_20958,N_18335,N_16276);
nor U20959 (N_20959,N_16765,N_16646);
and U20960 (N_20960,N_15968,N_17762);
and U20961 (N_20961,N_18713,N_16661);
nand U20962 (N_20962,N_17527,N_18146);
or U20963 (N_20963,N_17951,N_18470);
or U20964 (N_20964,N_18681,N_17689);
or U20965 (N_20965,N_16946,N_18522);
nand U20966 (N_20966,N_18570,N_18097);
and U20967 (N_20967,N_17396,N_17546);
nand U20968 (N_20968,N_16906,N_17929);
and U20969 (N_20969,N_16600,N_17539);
and U20970 (N_20970,N_16509,N_18736);
nand U20971 (N_20971,N_18500,N_16847);
nand U20972 (N_20972,N_17577,N_18306);
and U20973 (N_20973,N_17544,N_16607);
nor U20974 (N_20974,N_16092,N_17056);
and U20975 (N_20975,N_18367,N_18677);
nand U20976 (N_20976,N_18487,N_17426);
nand U20977 (N_20977,N_17364,N_16837);
and U20978 (N_20978,N_16041,N_16762);
nor U20979 (N_20979,N_18465,N_17933);
nand U20980 (N_20980,N_16046,N_17485);
nor U20981 (N_20981,N_18237,N_18691);
nor U20982 (N_20982,N_17220,N_15734);
or U20983 (N_20983,N_17664,N_16398);
xnor U20984 (N_20984,N_17754,N_17281);
and U20985 (N_20985,N_15712,N_16633);
nand U20986 (N_20986,N_17574,N_18257);
and U20987 (N_20987,N_18218,N_17816);
nor U20988 (N_20988,N_17931,N_18507);
and U20989 (N_20989,N_16926,N_18373);
or U20990 (N_20990,N_15697,N_17573);
xor U20991 (N_20991,N_15656,N_18485);
and U20992 (N_20992,N_18220,N_17947);
and U20993 (N_20993,N_18398,N_17886);
and U20994 (N_20994,N_17006,N_18097);
nand U20995 (N_20995,N_17620,N_18353);
and U20996 (N_20996,N_15805,N_18422);
nor U20997 (N_20997,N_17836,N_16318);
or U20998 (N_20998,N_18256,N_18049);
or U20999 (N_20999,N_16492,N_16843);
nand U21000 (N_21000,N_16217,N_18667);
nor U21001 (N_21001,N_18700,N_18098);
nand U21002 (N_21002,N_16003,N_16805);
nor U21003 (N_21003,N_18399,N_15926);
and U21004 (N_21004,N_16272,N_17414);
or U21005 (N_21005,N_16035,N_17664);
nor U21006 (N_21006,N_18357,N_17356);
or U21007 (N_21007,N_17862,N_17798);
nor U21008 (N_21008,N_16506,N_16038);
and U21009 (N_21009,N_18614,N_16488);
nor U21010 (N_21010,N_17838,N_16605);
nor U21011 (N_21011,N_18586,N_18596);
or U21012 (N_21012,N_15656,N_16536);
nand U21013 (N_21013,N_17007,N_17263);
xnor U21014 (N_21014,N_17718,N_15806);
or U21015 (N_21015,N_15990,N_16895);
nor U21016 (N_21016,N_15834,N_15757);
nor U21017 (N_21017,N_17173,N_15811);
or U21018 (N_21018,N_16025,N_16266);
nand U21019 (N_21019,N_18040,N_17711);
nor U21020 (N_21020,N_16913,N_18224);
nor U21021 (N_21021,N_15689,N_16849);
xor U21022 (N_21022,N_15627,N_18262);
nor U21023 (N_21023,N_15928,N_16331);
or U21024 (N_21024,N_18584,N_17835);
and U21025 (N_21025,N_16931,N_16437);
nand U21026 (N_21026,N_15939,N_16696);
or U21027 (N_21027,N_16882,N_17052);
nand U21028 (N_21028,N_17502,N_15912);
and U21029 (N_21029,N_17119,N_18744);
nand U21030 (N_21030,N_16287,N_18236);
or U21031 (N_21031,N_15919,N_18451);
nor U21032 (N_21032,N_17098,N_16609);
nand U21033 (N_21033,N_17240,N_17900);
or U21034 (N_21034,N_16546,N_16362);
nor U21035 (N_21035,N_18129,N_16439);
and U21036 (N_21036,N_18706,N_16755);
nor U21037 (N_21037,N_17168,N_17232);
and U21038 (N_21038,N_16371,N_17080);
nand U21039 (N_21039,N_16196,N_17483);
and U21040 (N_21040,N_16295,N_18095);
nand U21041 (N_21041,N_15645,N_15803);
or U21042 (N_21042,N_15930,N_17177);
nand U21043 (N_21043,N_18418,N_17572);
and U21044 (N_21044,N_16657,N_17585);
or U21045 (N_21045,N_16589,N_17990);
nand U21046 (N_21046,N_15680,N_15788);
and U21047 (N_21047,N_15732,N_18316);
nand U21048 (N_21048,N_16608,N_16285);
nand U21049 (N_21049,N_16526,N_16970);
or U21050 (N_21050,N_16592,N_17402);
xor U21051 (N_21051,N_17265,N_18293);
nor U21052 (N_21052,N_16892,N_17408);
and U21053 (N_21053,N_15665,N_17735);
and U21054 (N_21054,N_17986,N_17425);
nor U21055 (N_21055,N_16714,N_18616);
and U21056 (N_21056,N_17226,N_17178);
nor U21057 (N_21057,N_17618,N_16749);
nor U21058 (N_21058,N_18600,N_18039);
and U21059 (N_21059,N_15639,N_15868);
and U21060 (N_21060,N_15780,N_16112);
or U21061 (N_21061,N_17154,N_16158);
or U21062 (N_21062,N_16455,N_17788);
xnor U21063 (N_21063,N_17152,N_16135);
xor U21064 (N_21064,N_16421,N_16505);
or U21065 (N_21065,N_16788,N_15895);
nor U21066 (N_21066,N_16919,N_15722);
or U21067 (N_21067,N_17768,N_17457);
nand U21068 (N_21068,N_15856,N_18447);
or U21069 (N_21069,N_18077,N_17257);
nor U21070 (N_21070,N_16038,N_17863);
nand U21071 (N_21071,N_18508,N_17274);
nor U21072 (N_21072,N_17248,N_16133);
nor U21073 (N_21073,N_17596,N_17573);
nand U21074 (N_21074,N_17476,N_18146);
and U21075 (N_21075,N_17194,N_17707);
and U21076 (N_21076,N_18670,N_17327);
nor U21077 (N_21077,N_18153,N_17964);
nor U21078 (N_21078,N_17901,N_16711);
or U21079 (N_21079,N_17393,N_17878);
nand U21080 (N_21080,N_16735,N_16464);
and U21081 (N_21081,N_15835,N_15863);
xnor U21082 (N_21082,N_18271,N_17317);
and U21083 (N_21083,N_18558,N_18367);
nand U21084 (N_21084,N_18600,N_16545);
nor U21085 (N_21085,N_16116,N_16072);
or U21086 (N_21086,N_16580,N_16939);
or U21087 (N_21087,N_16985,N_18377);
and U21088 (N_21088,N_17460,N_16843);
or U21089 (N_21089,N_17949,N_18335);
nor U21090 (N_21090,N_18742,N_17357);
and U21091 (N_21091,N_16390,N_17448);
nand U21092 (N_21092,N_16678,N_18376);
and U21093 (N_21093,N_15829,N_16028);
nand U21094 (N_21094,N_16029,N_17210);
or U21095 (N_21095,N_15669,N_17838);
or U21096 (N_21096,N_16899,N_16349);
and U21097 (N_21097,N_16253,N_16857);
or U21098 (N_21098,N_18195,N_15819);
nor U21099 (N_21099,N_16341,N_15890);
and U21100 (N_21100,N_18474,N_18589);
and U21101 (N_21101,N_16244,N_16069);
nand U21102 (N_21102,N_18344,N_15841);
and U21103 (N_21103,N_17192,N_16147);
and U21104 (N_21104,N_16537,N_17476);
nor U21105 (N_21105,N_16919,N_15984);
nand U21106 (N_21106,N_17692,N_16802);
and U21107 (N_21107,N_15889,N_17044);
nand U21108 (N_21108,N_16207,N_17122);
or U21109 (N_21109,N_17146,N_18180);
nand U21110 (N_21110,N_15811,N_17286);
xor U21111 (N_21111,N_17055,N_18129);
nand U21112 (N_21112,N_17536,N_15670);
nand U21113 (N_21113,N_18628,N_17555);
or U21114 (N_21114,N_17158,N_17583);
and U21115 (N_21115,N_17993,N_17496);
nor U21116 (N_21116,N_15759,N_18018);
or U21117 (N_21117,N_17346,N_17956);
nor U21118 (N_21118,N_16854,N_17337);
and U21119 (N_21119,N_17772,N_17988);
and U21120 (N_21120,N_17800,N_16809);
nor U21121 (N_21121,N_17927,N_16910);
nand U21122 (N_21122,N_18676,N_17739);
nand U21123 (N_21123,N_16484,N_15852);
or U21124 (N_21124,N_18081,N_15696);
or U21125 (N_21125,N_16358,N_16655);
nor U21126 (N_21126,N_17203,N_17567);
and U21127 (N_21127,N_16381,N_16715);
nand U21128 (N_21128,N_17705,N_16092);
nand U21129 (N_21129,N_17191,N_18348);
nor U21130 (N_21130,N_16526,N_15942);
and U21131 (N_21131,N_18664,N_15648);
or U21132 (N_21132,N_17834,N_16767);
or U21133 (N_21133,N_18205,N_18030);
xnor U21134 (N_21134,N_18550,N_18506);
nor U21135 (N_21135,N_17816,N_18679);
or U21136 (N_21136,N_16448,N_17234);
xnor U21137 (N_21137,N_17053,N_17317);
nor U21138 (N_21138,N_18093,N_18655);
or U21139 (N_21139,N_16249,N_18512);
and U21140 (N_21140,N_16057,N_17975);
nand U21141 (N_21141,N_15790,N_16870);
and U21142 (N_21142,N_16937,N_16173);
and U21143 (N_21143,N_17106,N_15630);
or U21144 (N_21144,N_18277,N_15704);
nand U21145 (N_21145,N_17932,N_17878);
xnor U21146 (N_21146,N_17005,N_18292);
nor U21147 (N_21147,N_17200,N_17052);
or U21148 (N_21148,N_17795,N_16830);
nand U21149 (N_21149,N_18451,N_16444);
xnor U21150 (N_21150,N_17391,N_17053);
or U21151 (N_21151,N_16974,N_16095);
xor U21152 (N_21152,N_18260,N_16911);
nand U21153 (N_21153,N_18538,N_18720);
nor U21154 (N_21154,N_17015,N_16723);
xnor U21155 (N_21155,N_18567,N_17921);
nor U21156 (N_21156,N_17653,N_18612);
or U21157 (N_21157,N_18246,N_16084);
xor U21158 (N_21158,N_16193,N_16095);
nand U21159 (N_21159,N_15818,N_16155);
or U21160 (N_21160,N_18696,N_17594);
and U21161 (N_21161,N_16937,N_18659);
or U21162 (N_21162,N_17347,N_16478);
nand U21163 (N_21163,N_15881,N_16095);
or U21164 (N_21164,N_16405,N_16166);
nor U21165 (N_21165,N_18574,N_17698);
nor U21166 (N_21166,N_16790,N_16611);
nand U21167 (N_21167,N_18173,N_15941);
or U21168 (N_21168,N_17990,N_18494);
and U21169 (N_21169,N_16670,N_15682);
xnor U21170 (N_21170,N_16953,N_18608);
nor U21171 (N_21171,N_17792,N_16369);
nor U21172 (N_21172,N_16362,N_16487);
nand U21173 (N_21173,N_18605,N_18082);
and U21174 (N_21174,N_17357,N_16760);
and U21175 (N_21175,N_17614,N_16827);
xor U21176 (N_21176,N_15822,N_18445);
nand U21177 (N_21177,N_16143,N_16886);
or U21178 (N_21178,N_16743,N_16623);
nand U21179 (N_21179,N_18520,N_17855);
or U21180 (N_21180,N_18401,N_17281);
nand U21181 (N_21181,N_18600,N_18238);
and U21182 (N_21182,N_16565,N_18177);
nor U21183 (N_21183,N_17813,N_17273);
nor U21184 (N_21184,N_16462,N_17839);
or U21185 (N_21185,N_15634,N_16580);
nand U21186 (N_21186,N_18434,N_16172);
or U21187 (N_21187,N_18412,N_16324);
nand U21188 (N_21188,N_15763,N_18478);
nand U21189 (N_21189,N_15882,N_18168);
nor U21190 (N_21190,N_15756,N_17150);
and U21191 (N_21191,N_17431,N_17805);
nand U21192 (N_21192,N_17294,N_17386);
nor U21193 (N_21193,N_16098,N_18374);
xnor U21194 (N_21194,N_15702,N_18659);
nor U21195 (N_21195,N_18288,N_18003);
or U21196 (N_21196,N_16680,N_18665);
nand U21197 (N_21197,N_17360,N_17341);
nand U21198 (N_21198,N_17915,N_16324);
or U21199 (N_21199,N_18501,N_18150);
nand U21200 (N_21200,N_17242,N_16731);
nor U21201 (N_21201,N_17785,N_17596);
or U21202 (N_21202,N_17610,N_17659);
nor U21203 (N_21203,N_15874,N_18555);
or U21204 (N_21204,N_16909,N_17250);
xor U21205 (N_21205,N_16831,N_16508);
xor U21206 (N_21206,N_15890,N_16261);
nor U21207 (N_21207,N_17113,N_17681);
nand U21208 (N_21208,N_16150,N_17411);
nand U21209 (N_21209,N_17646,N_17408);
nor U21210 (N_21210,N_18050,N_15847);
nand U21211 (N_21211,N_17271,N_16712);
nor U21212 (N_21212,N_16419,N_16311);
nor U21213 (N_21213,N_18498,N_17332);
and U21214 (N_21214,N_17268,N_17856);
xnor U21215 (N_21215,N_17276,N_17996);
nor U21216 (N_21216,N_18385,N_17771);
nor U21217 (N_21217,N_18361,N_17894);
nor U21218 (N_21218,N_16626,N_17220);
and U21219 (N_21219,N_17016,N_18628);
nand U21220 (N_21220,N_15774,N_18356);
nand U21221 (N_21221,N_17328,N_18138);
xor U21222 (N_21222,N_16730,N_16489);
nor U21223 (N_21223,N_18153,N_17367);
nor U21224 (N_21224,N_16162,N_18134);
and U21225 (N_21225,N_17581,N_18474);
or U21226 (N_21226,N_18733,N_16501);
and U21227 (N_21227,N_16606,N_16858);
or U21228 (N_21228,N_16846,N_16638);
nand U21229 (N_21229,N_18719,N_16513);
nor U21230 (N_21230,N_16649,N_17622);
nor U21231 (N_21231,N_16769,N_16137);
nor U21232 (N_21232,N_16836,N_17886);
nand U21233 (N_21233,N_16066,N_15707);
nor U21234 (N_21234,N_15735,N_16586);
nor U21235 (N_21235,N_17778,N_17061);
or U21236 (N_21236,N_17560,N_17405);
or U21237 (N_21237,N_17707,N_17206);
nor U21238 (N_21238,N_16694,N_17947);
nor U21239 (N_21239,N_17871,N_17211);
nand U21240 (N_21240,N_18334,N_16504);
or U21241 (N_21241,N_16941,N_18451);
and U21242 (N_21242,N_18351,N_18423);
nand U21243 (N_21243,N_18502,N_16168);
nor U21244 (N_21244,N_18067,N_18252);
xnor U21245 (N_21245,N_17392,N_17411);
or U21246 (N_21246,N_18535,N_16185);
or U21247 (N_21247,N_18308,N_16961);
or U21248 (N_21248,N_18031,N_18092);
nand U21249 (N_21249,N_18385,N_17088);
nor U21250 (N_21250,N_17994,N_17387);
nor U21251 (N_21251,N_15877,N_16196);
nand U21252 (N_21252,N_15726,N_15636);
nor U21253 (N_21253,N_15720,N_17437);
xor U21254 (N_21254,N_16421,N_18259);
nor U21255 (N_21255,N_16352,N_18167);
xor U21256 (N_21256,N_17518,N_17512);
nor U21257 (N_21257,N_16746,N_16042);
and U21258 (N_21258,N_17974,N_18691);
and U21259 (N_21259,N_16264,N_18167);
nor U21260 (N_21260,N_17913,N_16017);
or U21261 (N_21261,N_18346,N_16257);
xnor U21262 (N_21262,N_16097,N_16716);
nor U21263 (N_21263,N_16452,N_15797);
nand U21264 (N_21264,N_16561,N_15766);
or U21265 (N_21265,N_18592,N_17399);
nand U21266 (N_21266,N_16422,N_16326);
xor U21267 (N_21267,N_17032,N_17564);
nor U21268 (N_21268,N_15829,N_15889);
nand U21269 (N_21269,N_17090,N_17597);
nand U21270 (N_21270,N_17575,N_16638);
nand U21271 (N_21271,N_18364,N_16602);
nor U21272 (N_21272,N_16525,N_17712);
nor U21273 (N_21273,N_15712,N_18201);
nor U21274 (N_21274,N_16156,N_17553);
and U21275 (N_21275,N_16977,N_16756);
or U21276 (N_21276,N_18504,N_16496);
nand U21277 (N_21277,N_18658,N_16364);
and U21278 (N_21278,N_17039,N_17159);
nand U21279 (N_21279,N_16195,N_18218);
and U21280 (N_21280,N_17011,N_17605);
nor U21281 (N_21281,N_15813,N_18630);
nor U21282 (N_21282,N_16279,N_18689);
or U21283 (N_21283,N_17302,N_16998);
and U21284 (N_21284,N_18279,N_18616);
xnor U21285 (N_21285,N_18394,N_16931);
or U21286 (N_21286,N_16956,N_17086);
or U21287 (N_21287,N_16398,N_17675);
nand U21288 (N_21288,N_17724,N_16634);
nand U21289 (N_21289,N_15858,N_16138);
xor U21290 (N_21290,N_16997,N_18641);
and U21291 (N_21291,N_16411,N_17914);
and U21292 (N_21292,N_17237,N_17347);
nor U21293 (N_21293,N_17739,N_15985);
and U21294 (N_21294,N_15734,N_17910);
nand U21295 (N_21295,N_18027,N_17886);
xor U21296 (N_21296,N_16757,N_18089);
nor U21297 (N_21297,N_18251,N_18155);
or U21298 (N_21298,N_16179,N_17967);
or U21299 (N_21299,N_16372,N_16152);
nand U21300 (N_21300,N_15903,N_17458);
nand U21301 (N_21301,N_17127,N_16531);
and U21302 (N_21302,N_17842,N_18738);
or U21303 (N_21303,N_17009,N_16782);
and U21304 (N_21304,N_15644,N_17621);
nor U21305 (N_21305,N_17008,N_18453);
nand U21306 (N_21306,N_16769,N_18111);
and U21307 (N_21307,N_15726,N_18638);
or U21308 (N_21308,N_17754,N_18255);
nor U21309 (N_21309,N_16011,N_17245);
nand U21310 (N_21310,N_16082,N_18230);
xor U21311 (N_21311,N_16058,N_15925);
and U21312 (N_21312,N_15988,N_18027);
and U21313 (N_21313,N_15678,N_17940);
nor U21314 (N_21314,N_18368,N_16583);
nand U21315 (N_21315,N_17249,N_16407);
nand U21316 (N_21316,N_16410,N_18633);
nor U21317 (N_21317,N_16315,N_18166);
nand U21318 (N_21318,N_17251,N_18278);
nand U21319 (N_21319,N_16147,N_15989);
or U21320 (N_21320,N_17521,N_17154);
and U21321 (N_21321,N_16174,N_16146);
xor U21322 (N_21322,N_17356,N_18062);
xnor U21323 (N_21323,N_18049,N_16235);
nor U21324 (N_21324,N_16111,N_18287);
nand U21325 (N_21325,N_16975,N_18375);
xnor U21326 (N_21326,N_15829,N_16057);
nand U21327 (N_21327,N_16713,N_16076);
nor U21328 (N_21328,N_16337,N_16753);
nor U21329 (N_21329,N_16038,N_15794);
or U21330 (N_21330,N_16661,N_15924);
nor U21331 (N_21331,N_15902,N_17330);
xnor U21332 (N_21332,N_16361,N_17073);
nand U21333 (N_21333,N_16425,N_16567);
and U21334 (N_21334,N_17721,N_18262);
nor U21335 (N_21335,N_16515,N_18582);
nor U21336 (N_21336,N_17062,N_17240);
or U21337 (N_21337,N_17554,N_18397);
and U21338 (N_21338,N_18673,N_16057);
nand U21339 (N_21339,N_16147,N_17968);
nor U21340 (N_21340,N_16952,N_18744);
nand U21341 (N_21341,N_16465,N_16359);
or U21342 (N_21342,N_16562,N_17706);
nand U21343 (N_21343,N_16798,N_17148);
and U21344 (N_21344,N_16429,N_16748);
nand U21345 (N_21345,N_15838,N_17933);
nor U21346 (N_21346,N_18039,N_15856);
nand U21347 (N_21347,N_18451,N_17913);
and U21348 (N_21348,N_18351,N_17441);
or U21349 (N_21349,N_16973,N_17974);
xnor U21350 (N_21350,N_17493,N_18128);
xnor U21351 (N_21351,N_18493,N_17042);
nor U21352 (N_21352,N_16730,N_16061);
nor U21353 (N_21353,N_15739,N_17480);
nor U21354 (N_21354,N_15954,N_17829);
nand U21355 (N_21355,N_15650,N_16864);
or U21356 (N_21356,N_16490,N_18263);
xnor U21357 (N_21357,N_17080,N_18253);
nor U21358 (N_21358,N_17368,N_17752);
and U21359 (N_21359,N_15770,N_17303);
nand U21360 (N_21360,N_18547,N_15854);
xor U21361 (N_21361,N_16084,N_18011);
nand U21362 (N_21362,N_17561,N_15995);
or U21363 (N_21363,N_16073,N_18140);
or U21364 (N_21364,N_17859,N_16290);
xor U21365 (N_21365,N_16675,N_18607);
or U21366 (N_21366,N_17537,N_16949);
or U21367 (N_21367,N_17051,N_17387);
or U21368 (N_21368,N_16175,N_17661);
nand U21369 (N_21369,N_18224,N_18718);
or U21370 (N_21370,N_16896,N_15969);
nand U21371 (N_21371,N_16105,N_16300);
and U21372 (N_21372,N_16232,N_18601);
or U21373 (N_21373,N_18403,N_17912);
and U21374 (N_21374,N_17772,N_16333);
nor U21375 (N_21375,N_15822,N_17563);
and U21376 (N_21376,N_16744,N_17686);
nor U21377 (N_21377,N_17934,N_18059);
or U21378 (N_21378,N_17993,N_16573);
xnor U21379 (N_21379,N_17676,N_15997);
or U21380 (N_21380,N_17550,N_18286);
xor U21381 (N_21381,N_16254,N_16505);
nand U21382 (N_21382,N_18057,N_15790);
and U21383 (N_21383,N_16147,N_16345);
or U21384 (N_21384,N_16551,N_17456);
or U21385 (N_21385,N_16857,N_18155);
nor U21386 (N_21386,N_15786,N_17688);
or U21387 (N_21387,N_16253,N_16050);
and U21388 (N_21388,N_16132,N_17962);
xnor U21389 (N_21389,N_16070,N_16191);
and U21390 (N_21390,N_15672,N_17179);
xnor U21391 (N_21391,N_17839,N_16936);
and U21392 (N_21392,N_17784,N_16612);
nand U21393 (N_21393,N_18205,N_16144);
xnor U21394 (N_21394,N_18577,N_16569);
and U21395 (N_21395,N_16723,N_16117);
nand U21396 (N_21396,N_17349,N_16001);
nand U21397 (N_21397,N_17612,N_16201);
or U21398 (N_21398,N_16839,N_18246);
nand U21399 (N_21399,N_16003,N_16651);
nor U21400 (N_21400,N_16317,N_18591);
or U21401 (N_21401,N_18258,N_18050);
nand U21402 (N_21402,N_16770,N_16574);
or U21403 (N_21403,N_18703,N_17619);
or U21404 (N_21404,N_16347,N_17143);
or U21405 (N_21405,N_17326,N_15895);
or U21406 (N_21406,N_18284,N_17629);
nand U21407 (N_21407,N_17383,N_16725);
or U21408 (N_21408,N_18585,N_16839);
xor U21409 (N_21409,N_17435,N_16713);
nor U21410 (N_21410,N_16155,N_17435);
and U21411 (N_21411,N_16427,N_16615);
nand U21412 (N_21412,N_15999,N_15952);
xnor U21413 (N_21413,N_17476,N_17458);
nor U21414 (N_21414,N_16355,N_18517);
nor U21415 (N_21415,N_15734,N_16295);
nor U21416 (N_21416,N_15661,N_18095);
or U21417 (N_21417,N_17455,N_17152);
and U21418 (N_21418,N_16557,N_16262);
nor U21419 (N_21419,N_17258,N_17149);
nand U21420 (N_21420,N_18099,N_18102);
and U21421 (N_21421,N_18245,N_18153);
nand U21422 (N_21422,N_16642,N_17796);
or U21423 (N_21423,N_16138,N_17503);
or U21424 (N_21424,N_16974,N_16682);
and U21425 (N_21425,N_16255,N_17108);
and U21426 (N_21426,N_16089,N_17091);
nor U21427 (N_21427,N_17578,N_17787);
and U21428 (N_21428,N_17099,N_18336);
and U21429 (N_21429,N_17520,N_16328);
and U21430 (N_21430,N_16153,N_16943);
xor U21431 (N_21431,N_16462,N_17020);
nor U21432 (N_21432,N_15814,N_17339);
nand U21433 (N_21433,N_16194,N_15912);
or U21434 (N_21434,N_18284,N_18216);
and U21435 (N_21435,N_18678,N_16550);
nand U21436 (N_21436,N_17310,N_16695);
and U21437 (N_21437,N_15706,N_16468);
xnor U21438 (N_21438,N_15845,N_17181);
and U21439 (N_21439,N_17629,N_16694);
and U21440 (N_21440,N_18320,N_18081);
nor U21441 (N_21441,N_15852,N_15901);
xor U21442 (N_21442,N_18287,N_16799);
nor U21443 (N_21443,N_17429,N_16762);
or U21444 (N_21444,N_16746,N_17152);
nor U21445 (N_21445,N_16799,N_17569);
or U21446 (N_21446,N_16659,N_18608);
nor U21447 (N_21447,N_17894,N_16689);
xnor U21448 (N_21448,N_15929,N_17531);
xor U21449 (N_21449,N_17693,N_17732);
nand U21450 (N_21450,N_17145,N_17662);
and U21451 (N_21451,N_17073,N_17796);
and U21452 (N_21452,N_17010,N_17614);
or U21453 (N_21453,N_18439,N_17470);
xor U21454 (N_21454,N_17692,N_18145);
nor U21455 (N_21455,N_16503,N_16335);
xnor U21456 (N_21456,N_18449,N_16297);
or U21457 (N_21457,N_18055,N_17060);
and U21458 (N_21458,N_18443,N_18446);
nand U21459 (N_21459,N_17777,N_18165);
nand U21460 (N_21460,N_17064,N_18452);
and U21461 (N_21461,N_16237,N_16922);
or U21462 (N_21462,N_15628,N_15680);
nand U21463 (N_21463,N_17799,N_18694);
and U21464 (N_21464,N_18069,N_18617);
or U21465 (N_21465,N_17065,N_18071);
nand U21466 (N_21466,N_15768,N_15837);
nor U21467 (N_21467,N_16751,N_18142);
and U21468 (N_21468,N_17254,N_17747);
nand U21469 (N_21469,N_15716,N_16516);
nor U21470 (N_21470,N_16962,N_16259);
nor U21471 (N_21471,N_16149,N_16529);
xor U21472 (N_21472,N_15810,N_17548);
nand U21473 (N_21473,N_18362,N_17675);
nand U21474 (N_21474,N_17250,N_16730);
nor U21475 (N_21475,N_18421,N_15754);
nand U21476 (N_21476,N_16942,N_16999);
nand U21477 (N_21477,N_16478,N_16994);
and U21478 (N_21478,N_18119,N_18353);
nand U21479 (N_21479,N_16550,N_16446);
or U21480 (N_21480,N_18694,N_18415);
nor U21481 (N_21481,N_18379,N_15855);
nand U21482 (N_21482,N_16761,N_17470);
nand U21483 (N_21483,N_18615,N_16704);
nor U21484 (N_21484,N_16262,N_18608);
or U21485 (N_21485,N_17979,N_17596);
or U21486 (N_21486,N_18127,N_18424);
or U21487 (N_21487,N_18242,N_16079);
and U21488 (N_21488,N_15686,N_16347);
and U21489 (N_21489,N_15782,N_17739);
nor U21490 (N_21490,N_17232,N_17290);
or U21491 (N_21491,N_17167,N_15937);
nand U21492 (N_21492,N_18524,N_18510);
or U21493 (N_21493,N_16188,N_16485);
and U21494 (N_21494,N_16889,N_18413);
and U21495 (N_21495,N_17577,N_18103);
nor U21496 (N_21496,N_16101,N_15703);
or U21497 (N_21497,N_15810,N_16632);
xnor U21498 (N_21498,N_17719,N_18437);
and U21499 (N_21499,N_17862,N_16620);
and U21500 (N_21500,N_18607,N_16463);
or U21501 (N_21501,N_17604,N_17095);
nand U21502 (N_21502,N_16887,N_15736);
nor U21503 (N_21503,N_17303,N_15874);
nand U21504 (N_21504,N_18554,N_16391);
or U21505 (N_21505,N_17158,N_16289);
or U21506 (N_21506,N_16953,N_18054);
and U21507 (N_21507,N_16359,N_16456);
nand U21508 (N_21508,N_18106,N_17399);
and U21509 (N_21509,N_16820,N_16438);
or U21510 (N_21510,N_17988,N_16903);
nand U21511 (N_21511,N_17155,N_18272);
nand U21512 (N_21512,N_17298,N_15799);
nor U21513 (N_21513,N_15845,N_16334);
and U21514 (N_21514,N_18740,N_17648);
nor U21515 (N_21515,N_17932,N_17006);
nand U21516 (N_21516,N_17925,N_18048);
nor U21517 (N_21517,N_16140,N_16063);
and U21518 (N_21518,N_17749,N_17992);
nor U21519 (N_21519,N_15637,N_17928);
or U21520 (N_21520,N_17355,N_15783);
nand U21521 (N_21521,N_15905,N_17156);
nor U21522 (N_21522,N_16929,N_18382);
nand U21523 (N_21523,N_18077,N_17938);
nor U21524 (N_21524,N_17013,N_17021);
and U21525 (N_21525,N_18257,N_17073);
nor U21526 (N_21526,N_17478,N_16967);
and U21527 (N_21527,N_16133,N_15989);
or U21528 (N_21528,N_18157,N_17869);
and U21529 (N_21529,N_17183,N_16923);
nand U21530 (N_21530,N_17321,N_16651);
and U21531 (N_21531,N_18584,N_16573);
and U21532 (N_21532,N_17165,N_18422);
or U21533 (N_21533,N_16796,N_18599);
or U21534 (N_21534,N_17503,N_17526);
or U21535 (N_21535,N_18646,N_17787);
xnor U21536 (N_21536,N_15789,N_17710);
and U21537 (N_21537,N_18345,N_17251);
and U21538 (N_21538,N_16360,N_16126);
nand U21539 (N_21539,N_18714,N_16074);
or U21540 (N_21540,N_15653,N_18049);
nand U21541 (N_21541,N_17569,N_15863);
nand U21542 (N_21542,N_17329,N_17045);
nor U21543 (N_21543,N_15931,N_17294);
nand U21544 (N_21544,N_17867,N_15911);
or U21545 (N_21545,N_16546,N_16251);
nand U21546 (N_21546,N_16815,N_18564);
xor U21547 (N_21547,N_17712,N_17230);
xnor U21548 (N_21548,N_16983,N_17920);
or U21549 (N_21549,N_16163,N_17000);
nor U21550 (N_21550,N_17980,N_18327);
nand U21551 (N_21551,N_18290,N_17230);
and U21552 (N_21552,N_15655,N_16829);
nor U21553 (N_21553,N_16553,N_16186);
and U21554 (N_21554,N_16420,N_15961);
and U21555 (N_21555,N_18368,N_17419);
nand U21556 (N_21556,N_16374,N_15654);
xnor U21557 (N_21557,N_18462,N_18245);
or U21558 (N_21558,N_18740,N_17437);
or U21559 (N_21559,N_17544,N_18076);
xnor U21560 (N_21560,N_17011,N_15838);
nand U21561 (N_21561,N_16016,N_18088);
or U21562 (N_21562,N_15957,N_17464);
nand U21563 (N_21563,N_15852,N_17749);
or U21564 (N_21564,N_16225,N_18713);
nand U21565 (N_21565,N_16655,N_15946);
nor U21566 (N_21566,N_17314,N_16818);
nand U21567 (N_21567,N_16843,N_16695);
or U21568 (N_21568,N_17751,N_18705);
or U21569 (N_21569,N_16761,N_16543);
nor U21570 (N_21570,N_16939,N_17073);
and U21571 (N_21571,N_17427,N_16957);
xor U21572 (N_21572,N_16912,N_17505);
and U21573 (N_21573,N_16920,N_17140);
nor U21574 (N_21574,N_17208,N_18451);
nand U21575 (N_21575,N_17285,N_18189);
or U21576 (N_21576,N_16934,N_17307);
and U21577 (N_21577,N_17086,N_17502);
and U21578 (N_21578,N_16536,N_17860);
nor U21579 (N_21579,N_16695,N_17131);
nor U21580 (N_21580,N_17393,N_16922);
or U21581 (N_21581,N_16995,N_16229);
xnor U21582 (N_21582,N_16767,N_18529);
nor U21583 (N_21583,N_18477,N_17449);
or U21584 (N_21584,N_18578,N_17899);
nand U21585 (N_21585,N_17920,N_17385);
or U21586 (N_21586,N_18551,N_16232);
xnor U21587 (N_21587,N_18450,N_17047);
or U21588 (N_21588,N_17063,N_17598);
or U21589 (N_21589,N_17985,N_18712);
nor U21590 (N_21590,N_16326,N_17923);
nor U21591 (N_21591,N_16037,N_15699);
and U21592 (N_21592,N_17025,N_16104);
and U21593 (N_21593,N_17063,N_17373);
or U21594 (N_21594,N_18213,N_17816);
nor U21595 (N_21595,N_18356,N_18589);
and U21596 (N_21596,N_18464,N_17608);
nand U21597 (N_21597,N_16092,N_18305);
nor U21598 (N_21598,N_16013,N_17507);
nand U21599 (N_21599,N_18276,N_15719);
nor U21600 (N_21600,N_16390,N_16965);
or U21601 (N_21601,N_18451,N_18093);
nor U21602 (N_21602,N_16946,N_18619);
or U21603 (N_21603,N_16230,N_17013);
nor U21604 (N_21604,N_18632,N_15819);
nand U21605 (N_21605,N_18662,N_18079);
and U21606 (N_21606,N_16650,N_18698);
nor U21607 (N_21607,N_16206,N_15873);
nand U21608 (N_21608,N_17249,N_17174);
nor U21609 (N_21609,N_18477,N_18242);
xnor U21610 (N_21610,N_16830,N_16650);
xor U21611 (N_21611,N_16894,N_18615);
nand U21612 (N_21612,N_16733,N_17783);
nand U21613 (N_21613,N_15955,N_17570);
or U21614 (N_21614,N_16626,N_16304);
nor U21615 (N_21615,N_16183,N_18428);
nor U21616 (N_21616,N_16658,N_16606);
nor U21617 (N_21617,N_16395,N_16918);
nor U21618 (N_21618,N_16261,N_16968);
nand U21619 (N_21619,N_18253,N_16344);
nor U21620 (N_21620,N_17589,N_16910);
or U21621 (N_21621,N_15647,N_16795);
nand U21622 (N_21622,N_16938,N_18269);
and U21623 (N_21623,N_16404,N_15998);
xor U21624 (N_21624,N_16356,N_17267);
or U21625 (N_21625,N_17058,N_18009);
xor U21626 (N_21626,N_16678,N_18484);
or U21627 (N_21627,N_17089,N_18728);
and U21628 (N_21628,N_16225,N_16986);
or U21629 (N_21629,N_17108,N_17807);
nand U21630 (N_21630,N_17997,N_18425);
nand U21631 (N_21631,N_18242,N_17039);
or U21632 (N_21632,N_17400,N_18507);
nand U21633 (N_21633,N_18362,N_16114);
nor U21634 (N_21634,N_18251,N_18599);
or U21635 (N_21635,N_15684,N_17252);
or U21636 (N_21636,N_16103,N_16731);
nand U21637 (N_21637,N_15664,N_16777);
nand U21638 (N_21638,N_17598,N_16126);
nor U21639 (N_21639,N_15795,N_17991);
nand U21640 (N_21640,N_18259,N_17191);
or U21641 (N_21641,N_18114,N_17551);
nand U21642 (N_21642,N_15777,N_17494);
nor U21643 (N_21643,N_16559,N_17268);
or U21644 (N_21644,N_17694,N_16823);
and U21645 (N_21645,N_17788,N_18226);
nand U21646 (N_21646,N_18378,N_17528);
or U21647 (N_21647,N_17866,N_18453);
and U21648 (N_21648,N_16395,N_17996);
or U21649 (N_21649,N_16034,N_16665);
nand U21650 (N_21650,N_17476,N_15690);
or U21651 (N_21651,N_16718,N_16604);
nor U21652 (N_21652,N_18196,N_18640);
or U21653 (N_21653,N_16488,N_18319);
nand U21654 (N_21654,N_16858,N_17592);
or U21655 (N_21655,N_18709,N_17859);
nand U21656 (N_21656,N_15852,N_16570);
or U21657 (N_21657,N_15912,N_18001);
or U21658 (N_21658,N_18186,N_17343);
nand U21659 (N_21659,N_16163,N_16834);
and U21660 (N_21660,N_18036,N_16459);
and U21661 (N_21661,N_17518,N_17134);
and U21662 (N_21662,N_15754,N_18675);
nand U21663 (N_21663,N_18442,N_18097);
nor U21664 (N_21664,N_16965,N_16261);
nor U21665 (N_21665,N_16113,N_18470);
nand U21666 (N_21666,N_16728,N_17622);
or U21667 (N_21667,N_18137,N_17523);
and U21668 (N_21668,N_17303,N_17088);
or U21669 (N_21669,N_15953,N_18107);
nor U21670 (N_21670,N_17816,N_17941);
or U21671 (N_21671,N_17992,N_16975);
or U21672 (N_21672,N_16278,N_17339);
nor U21673 (N_21673,N_16069,N_18385);
nand U21674 (N_21674,N_17412,N_17849);
nor U21675 (N_21675,N_16990,N_17815);
xor U21676 (N_21676,N_16092,N_16528);
nand U21677 (N_21677,N_17591,N_18440);
nand U21678 (N_21678,N_17293,N_17240);
xnor U21679 (N_21679,N_16136,N_17348);
nand U21680 (N_21680,N_16974,N_16050);
xor U21681 (N_21681,N_16541,N_17921);
nand U21682 (N_21682,N_16858,N_17083);
nand U21683 (N_21683,N_16739,N_18306);
or U21684 (N_21684,N_18694,N_15733);
or U21685 (N_21685,N_17974,N_15823);
nor U21686 (N_21686,N_18226,N_18405);
and U21687 (N_21687,N_18201,N_16121);
nor U21688 (N_21688,N_15716,N_17429);
nand U21689 (N_21689,N_16984,N_18153);
xnor U21690 (N_21690,N_18223,N_17290);
or U21691 (N_21691,N_16770,N_18385);
and U21692 (N_21692,N_17694,N_16348);
or U21693 (N_21693,N_17264,N_15856);
or U21694 (N_21694,N_17837,N_17608);
or U21695 (N_21695,N_16493,N_16043);
and U21696 (N_21696,N_17169,N_17282);
and U21697 (N_21697,N_17395,N_16677);
or U21698 (N_21698,N_18202,N_18602);
nand U21699 (N_21699,N_16085,N_16481);
xnor U21700 (N_21700,N_17824,N_17466);
nand U21701 (N_21701,N_15834,N_18431);
nand U21702 (N_21702,N_17027,N_17112);
nand U21703 (N_21703,N_16456,N_15761);
or U21704 (N_21704,N_16177,N_16909);
or U21705 (N_21705,N_16737,N_18109);
xor U21706 (N_21706,N_16767,N_17434);
and U21707 (N_21707,N_18630,N_18444);
xnor U21708 (N_21708,N_16715,N_16960);
xor U21709 (N_21709,N_17730,N_16883);
nand U21710 (N_21710,N_17157,N_17442);
and U21711 (N_21711,N_18278,N_18052);
and U21712 (N_21712,N_17129,N_15626);
or U21713 (N_21713,N_17243,N_16711);
xnor U21714 (N_21714,N_16173,N_16569);
nor U21715 (N_21715,N_15777,N_16965);
or U21716 (N_21716,N_17993,N_16485);
or U21717 (N_21717,N_18376,N_18271);
nand U21718 (N_21718,N_15967,N_17820);
nand U21719 (N_21719,N_16579,N_16562);
and U21720 (N_21720,N_15912,N_15961);
and U21721 (N_21721,N_16994,N_15870);
nor U21722 (N_21722,N_17530,N_18504);
xnor U21723 (N_21723,N_17095,N_16347);
nor U21724 (N_21724,N_18078,N_17602);
nand U21725 (N_21725,N_16997,N_15943);
nand U21726 (N_21726,N_16059,N_17141);
nor U21727 (N_21727,N_18633,N_16718);
nand U21728 (N_21728,N_18285,N_15880);
xnor U21729 (N_21729,N_17347,N_16636);
nor U21730 (N_21730,N_18277,N_17057);
nand U21731 (N_21731,N_17580,N_17273);
and U21732 (N_21732,N_16210,N_17071);
nor U21733 (N_21733,N_16755,N_16963);
nor U21734 (N_21734,N_17213,N_16994);
nor U21735 (N_21735,N_16864,N_17269);
or U21736 (N_21736,N_18324,N_18267);
nand U21737 (N_21737,N_15866,N_16878);
and U21738 (N_21738,N_18173,N_15629);
nor U21739 (N_21739,N_18131,N_16511);
nor U21740 (N_21740,N_17359,N_16158);
nor U21741 (N_21741,N_17477,N_15773);
and U21742 (N_21742,N_16236,N_16227);
nor U21743 (N_21743,N_16396,N_17070);
nand U21744 (N_21744,N_17393,N_18646);
nor U21745 (N_21745,N_18251,N_17114);
and U21746 (N_21746,N_16119,N_16201);
or U21747 (N_21747,N_18319,N_16476);
nor U21748 (N_21748,N_18392,N_18334);
and U21749 (N_21749,N_16808,N_17729);
nand U21750 (N_21750,N_17939,N_16233);
nor U21751 (N_21751,N_18118,N_17940);
and U21752 (N_21752,N_16602,N_18290);
and U21753 (N_21753,N_16441,N_16060);
nand U21754 (N_21754,N_18528,N_18212);
and U21755 (N_21755,N_16810,N_18149);
and U21756 (N_21756,N_18239,N_16193);
xor U21757 (N_21757,N_17292,N_17457);
nand U21758 (N_21758,N_18618,N_16031);
or U21759 (N_21759,N_17043,N_18312);
and U21760 (N_21760,N_17910,N_16422);
or U21761 (N_21761,N_17252,N_15907);
and U21762 (N_21762,N_16542,N_17356);
or U21763 (N_21763,N_17131,N_17356);
nor U21764 (N_21764,N_17523,N_15689);
or U21765 (N_21765,N_17724,N_17656);
nor U21766 (N_21766,N_16244,N_17674);
and U21767 (N_21767,N_16861,N_18518);
nor U21768 (N_21768,N_16066,N_18610);
nand U21769 (N_21769,N_17302,N_16905);
or U21770 (N_21770,N_17500,N_16067);
nor U21771 (N_21771,N_15867,N_17390);
nor U21772 (N_21772,N_17177,N_16556);
xor U21773 (N_21773,N_18460,N_17807);
or U21774 (N_21774,N_18359,N_18284);
xnor U21775 (N_21775,N_15887,N_17478);
and U21776 (N_21776,N_16834,N_17598);
or U21777 (N_21777,N_16727,N_18701);
nor U21778 (N_21778,N_18345,N_17376);
or U21779 (N_21779,N_16725,N_17927);
or U21780 (N_21780,N_17557,N_16008);
xnor U21781 (N_21781,N_16741,N_15982);
nand U21782 (N_21782,N_15913,N_16741);
xor U21783 (N_21783,N_16565,N_16906);
nand U21784 (N_21784,N_17730,N_17424);
and U21785 (N_21785,N_16909,N_18427);
nor U21786 (N_21786,N_16245,N_16262);
nand U21787 (N_21787,N_17508,N_16085);
or U21788 (N_21788,N_17075,N_17703);
and U21789 (N_21789,N_17682,N_15954);
xnor U21790 (N_21790,N_18145,N_17038);
nor U21791 (N_21791,N_16516,N_16967);
or U21792 (N_21792,N_17998,N_16438);
xor U21793 (N_21793,N_18234,N_17498);
or U21794 (N_21794,N_16705,N_18027);
and U21795 (N_21795,N_17578,N_17358);
nand U21796 (N_21796,N_17313,N_16188);
or U21797 (N_21797,N_18462,N_17528);
or U21798 (N_21798,N_16969,N_15988);
or U21799 (N_21799,N_17221,N_17268);
and U21800 (N_21800,N_16016,N_16205);
and U21801 (N_21801,N_18096,N_16553);
or U21802 (N_21802,N_17790,N_16977);
nor U21803 (N_21803,N_18586,N_17676);
nor U21804 (N_21804,N_17725,N_18336);
nand U21805 (N_21805,N_17468,N_17841);
nor U21806 (N_21806,N_17316,N_16750);
and U21807 (N_21807,N_17332,N_16884);
nor U21808 (N_21808,N_16801,N_15945);
nand U21809 (N_21809,N_16501,N_16779);
nor U21810 (N_21810,N_16541,N_17946);
and U21811 (N_21811,N_17184,N_17020);
xnor U21812 (N_21812,N_17261,N_18230);
and U21813 (N_21813,N_17083,N_16529);
and U21814 (N_21814,N_15803,N_18142);
xor U21815 (N_21815,N_17667,N_16552);
nand U21816 (N_21816,N_16210,N_15982);
nand U21817 (N_21817,N_15968,N_18223);
or U21818 (N_21818,N_16038,N_16838);
xor U21819 (N_21819,N_17462,N_18433);
xor U21820 (N_21820,N_18668,N_17254);
xor U21821 (N_21821,N_16340,N_17410);
nor U21822 (N_21822,N_16130,N_17068);
or U21823 (N_21823,N_16920,N_16676);
nor U21824 (N_21824,N_17058,N_17782);
and U21825 (N_21825,N_17222,N_16353);
and U21826 (N_21826,N_17467,N_17633);
or U21827 (N_21827,N_16108,N_17078);
or U21828 (N_21828,N_17249,N_18176);
nor U21829 (N_21829,N_17703,N_18173);
nor U21830 (N_21830,N_15865,N_16420);
or U21831 (N_21831,N_18620,N_17383);
nor U21832 (N_21832,N_15944,N_18467);
and U21833 (N_21833,N_17715,N_15655);
nand U21834 (N_21834,N_17674,N_16924);
nor U21835 (N_21835,N_16113,N_16307);
or U21836 (N_21836,N_18587,N_16530);
and U21837 (N_21837,N_18218,N_16855);
or U21838 (N_21838,N_16267,N_15887);
and U21839 (N_21839,N_18399,N_16104);
and U21840 (N_21840,N_18610,N_16462);
nand U21841 (N_21841,N_18594,N_17587);
nand U21842 (N_21842,N_16218,N_17959);
nand U21843 (N_21843,N_15669,N_15711);
nand U21844 (N_21844,N_16585,N_15977);
nand U21845 (N_21845,N_15834,N_18716);
or U21846 (N_21846,N_17204,N_15718);
nor U21847 (N_21847,N_18486,N_16667);
nor U21848 (N_21848,N_18747,N_16021);
and U21849 (N_21849,N_18239,N_17019);
nand U21850 (N_21850,N_16422,N_18570);
xnor U21851 (N_21851,N_17335,N_17351);
xor U21852 (N_21852,N_16433,N_16807);
nor U21853 (N_21853,N_16647,N_17053);
or U21854 (N_21854,N_17231,N_18367);
or U21855 (N_21855,N_16241,N_18594);
or U21856 (N_21856,N_18442,N_17434);
nor U21857 (N_21857,N_16015,N_17700);
nand U21858 (N_21858,N_16636,N_17063);
nand U21859 (N_21859,N_17197,N_17736);
nor U21860 (N_21860,N_18536,N_17115);
and U21861 (N_21861,N_15659,N_17782);
nor U21862 (N_21862,N_16350,N_15906);
and U21863 (N_21863,N_18389,N_15669);
nor U21864 (N_21864,N_15990,N_16059);
nand U21865 (N_21865,N_15787,N_17372);
nand U21866 (N_21866,N_18116,N_16378);
and U21867 (N_21867,N_18191,N_17132);
xor U21868 (N_21868,N_15824,N_16133);
or U21869 (N_21869,N_18199,N_16649);
and U21870 (N_21870,N_18076,N_15817);
and U21871 (N_21871,N_18235,N_15972);
and U21872 (N_21872,N_18357,N_16525);
nand U21873 (N_21873,N_17909,N_16410);
xnor U21874 (N_21874,N_17254,N_18369);
nand U21875 (N_21875,N_20343,N_21592);
nand U21876 (N_21876,N_20589,N_20474);
or U21877 (N_21877,N_18830,N_18858);
nand U21878 (N_21878,N_20385,N_21659);
and U21879 (N_21879,N_19034,N_19317);
nand U21880 (N_21880,N_20441,N_20078);
or U21881 (N_21881,N_20352,N_20550);
or U21882 (N_21882,N_19181,N_21189);
or U21883 (N_21883,N_18838,N_19710);
nand U21884 (N_21884,N_19168,N_19198);
or U21885 (N_21885,N_19142,N_18752);
nand U21886 (N_21886,N_20497,N_20193);
or U21887 (N_21887,N_21551,N_20137);
or U21888 (N_21888,N_20476,N_19328);
and U21889 (N_21889,N_20010,N_21338);
or U21890 (N_21890,N_20307,N_18982);
nor U21891 (N_21891,N_20319,N_21202);
nor U21892 (N_21892,N_20342,N_20825);
and U21893 (N_21893,N_20792,N_21020);
nor U21894 (N_21894,N_18831,N_19174);
nor U21895 (N_21895,N_19291,N_20379);
nor U21896 (N_21896,N_20454,N_20626);
or U21897 (N_21897,N_20644,N_20208);
nand U21898 (N_21898,N_20779,N_21815);
and U21899 (N_21899,N_20052,N_21574);
nand U21900 (N_21900,N_20599,N_21705);
or U21901 (N_21901,N_20676,N_21555);
or U21902 (N_21902,N_19072,N_21049);
or U21903 (N_21903,N_21625,N_21671);
xor U21904 (N_21904,N_21733,N_21023);
and U21905 (N_21905,N_19046,N_21642);
nor U21906 (N_21906,N_18907,N_18800);
xor U21907 (N_21907,N_18879,N_20752);
or U21908 (N_21908,N_20855,N_21250);
xor U21909 (N_21909,N_21639,N_21349);
and U21910 (N_21910,N_21026,N_21088);
nand U21911 (N_21911,N_19708,N_20748);
and U21912 (N_21912,N_21785,N_20255);
and U21913 (N_21913,N_19629,N_18821);
nand U21914 (N_21914,N_19895,N_21304);
or U21915 (N_21915,N_21107,N_21140);
nor U21916 (N_21916,N_21197,N_19082);
and U21917 (N_21917,N_20017,N_21399);
and U21918 (N_21918,N_20219,N_21697);
nand U21919 (N_21919,N_19136,N_19119);
nand U21920 (N_21920,N_21209,N_21110);
nor U21921 (N_21921,N_21097,N_19669);
nor U21922 (N_21922,N_19100,N_20224);
and U21923 (N_21923,N_21254,N_21729);
xnor U21924 (N_21924,N_19321,N_19070);
nand U21925 (N_21925,N_20108,N_21476);
or U21926 (N_21926,N_19149,N_19866);
nor U21927 (N_21927,N_19695,N_20522);
nand U21928 (N_21928,N_19733,N_19686);
nand U21929 (N_21929,N_21242,N_21068);
xor U21930 (N_21930,N_20483,N_21811);
nor U21931 (N_21931,N_20709,N_19165);
nor U21932 (N_21932,N_21211,N_19406);
nor U21933 (N_21933,N_20455,N_20958);
nand U21934 (N_21934,N_21360,N_19863);
xnor U21935 (N_21935,N_19097,N_19263);
and U21936 (N_21936,N_19915,N_18762);
nor U21937 (N_21937,N_20556,N_20396);
nand U21938 (N_21938,N_21104,N_20020);
and U21939 (N_21939,N_19252,N_19022);
or U21940 (N_21940,N_20292,N_21352);
nor U21941 (N_21941,N_21321,N_20911);
or U21942 (N_21942,N_20902,N_19088);
nand U21943 (N_21943,N_18914,N_20096);
and U21944 (N_21944,N_19945,N_19173);
xor U21945 (N_21945,N_21389,N_20510);
nand U21946 (N_21946,N_20138,N_21398);
and U21947 (N_21947,N_20783,N_18897);
nor U21948 (N_21948,N_19880,N_21050);
or U21949 (N_21949,N_19826,N_21220);
and U21950 (N_21950,N_21385,N_20251);
nand U21951 (N_21951,N_20953,N_20828);
and U21952 (N_21952,N_20298,N_19179);
nor U21953 (N_21953,N_21042,N_19290);
nand U21954 (N_21954,N_20140,N_20997);
nand U21955 (N_21955,N_21047,N_20749);
or U21956 (N_21956,N_20566,N_20555);
nand U21957 (N_21957,N_20120,N_19587);
nor U21958 (N_21958,N_21612,N_19466);
nand U21959 (N_21959,N_19287,N_19925);
and U21960 (N_21960,N_19967,N_19690);
nand U21961 (N_21961,N_19676,N_20194);
nand U21962 (N_21962,N_20452,N_19146);
xor U21963 (N_21963,N_21680,N_19738);
nand U21964 (N_21964,N_19527,N_19027);
nand U21965 (N_21965,N_20268,N_19847);
nor U21966 (N_21966,N_20403,N_21771);
or U21967 (N_21967,N_18895,N_20401);
nand U21968 (N_21968,N_20637,N_20025);
nand U21969 (N_21969,N_19790,N_18788);
nand U21970 (N_21970,N_20152,N_20692);
nand U21971 (N_21971,N_21358,N_18966);
or U21972 (N_21972,N_19621,N_20802);
or U21973 (N_21973,N_21062,N_20492);
and U21974 (N_21974,N_20972,N_20619);
xor U21975 (N_21975,N_20728,N_19218);
and U21976 (N_21976,N_19451,N_20593);
or U21977 (N_21977,N_21706,N_20485);
xor U21978 (N_21978,N_21421,N_21069);
nor U21979 (N_21979,N_19354,N_21505);
and U21980 (N_21980,N_20665,N_19151);
and U21981 (N_21981,N_19722,N_19260);
or U21982 (N_21982,N_19449,N_21278);
or U21983 (N_21983,N_21339,N_19481);
nand U21984 (N_21984,N_19023,N_20384);
xor U21985 (N_21985,N_21027,N_21801);
and U21986 (N_21986,N_18983,N_21134);
xor U21987 (N_21987,N_20229,N_19076);
xor U21988 (N_21988,N_21731,N_21786);
nand U21989 (N_21989,N_19414,N_18989);
nor U21990 (N_21990,N_19741,N_20773);
and U21991 (N_21991,N_19012,N_19315);
or U21992 (N_21992,N_21805,N_19734);
or U21993 (N_21993,N_19107,N_20710);
or U21994 (N_21994,N_20428,N_19066);
nor U21995 (N_21995,N_20439,N_20741);
and U21996 (N_21996,N_18969,N_19601);
xnor U21997 (N_21997,N_19721,N_21288);
nor U21998 (N_21998,N_20889,N_19170);
nor U21999 (N_21999,N_20920,N_20357);
nor U22000 (N_22000,N_20734,N_21131);
nand U22001 (N_22001,N_21586,N_21509);
and U22002 (N_22002,N_20252,N_18803);
nand U22003 (N_22003,N_19713,N_19507);
nor U22004 (N_22004,N_20894,N_20829);
xor U22005 (N_22005,N_20793,N_19484);
or U22006 (N_22006,N_20819,N_21116);
xor U22007 (N_22007,N_19110,N_20062);
nand U22008 (N_22008,N_20360,N_19965);
and U22009 (N_22009,N_21487,N_18841);
or U22010 (N_22010,N_20469,N_19843);
nor U22011 (N_22011,N_19247,N_21354);
and U22012 (N_22012,N_19646,N_20797);
or U22013 (N_22013,N_20854,N_21130);
or U22014 (N_22014,N_20071,N_20976);
nand U22015 (N_22015,N_21086,N_20055);
nand U22016 (N_22016,N_19832,N_21825);
or U22017 (N_22017,N_19517,N_19538);
nor U22018 (N_22018,N_19234,N_19467);
nor U22019 (N_22019,N_19586,N_21778);
or U22020 (N_22020,N_21065,N_20533);
nand U22021 (N_22021,N_21739,N_21522);
nor U22022 (N_22022,N_19759,N_19293);
nor U22023 (N_22023,N_18975,N_20707);
and U22024 (N_22024,N_20048,N_19368);
or U22025 (N_22025,N_21411,N_20100);
nand U22026 (N_22026,N_19063,N_20306);
and U22027 (N_22027,N_21529,N_20839);
and U22028 (N_22028,N_21307,N_20316);
and U22029 (N_22029,N_19954,N_20660);
and U22030 (N_22030,N_19374,N_21784);
nand U22031 (N_22031,N_20959,N_18869);
nand U22032 (N_22032,N_20060,N_21040);
nand U22033 (N_22033,N_19966,N_20277);
and U22034 (N_22034,N_20238,N_21206);
xnor U22035 (N_22035,N_21454,N_20930);
nand U22036 (N_22036,N_20568,N_20284);
nor U22037 (N_22037,N_21318,N_21426);
or U22038 (N_22038,N_21783,N_19504);
nand U22039 (N_22039,N_19184,N_19938);
or U22040 (N_22040,N_21275,N_20056);
nand U22041 (N_22041,N_20365,N_19771);
nand U22042 (N_22042,N_19200,N_21830);
and U22043 (N_22043,N_19786,N_20210);
nand U22044 (N_22044,N_19332,N_21851);
nand U22045 (N_22045,N_21565,N_20154);
nor U22046 (N_22046,N_21663,N_20253);
or U22047 (N_22047,N_20367,N_20868);
nand U22048 (N_22048,N_18962,N_21758);
nor U22049 (N_22049,N_18912,N_21618);
and U22050 (N_22050,N_19709,N_20267);
nand U22051 (N_22051,N_19319,N_21376);
nand U22052 (N_22052,N_19750,N_18943);
and U22053 (N_22053,N_18846,N_21218);
or U22054 (N_22054,N_21835,N_19788);
nand U22055 (N_22055,N_20870,N_21840);
and U22056 (N_22056,N_19091,N_19649);
nor U22057 (N_22057,N_20486,N_20076);
nand U22058 (N_22058,N_20195,N_19047);
and U22059 (N_22059,N_21214,N_19421);
xor U22060 (N_22060,N_19588,N_21442);
and U22061 (N_22061,N_21704,N_21256);
nor U22062 (N_22062,N_21407,N_20711);
nand U22063 (N_22063,N_20426,N_21306);
or U22064 (N_22064,N_21543,N_19336);
or U22065 (N_22065,N_21164,N_20961);
xnor U22066 (N_22066,N_19124,N_21446);
and U22067 (N_22067,N_20756,N_21858);
nor U22068 (N_22068,N_21362,N_19192);
and U22069 (N_22069,N_21695,N_18790);
or U22070 (N_22070,N_18786,N_19460);
nor U22071 (N_22071,N_20146,N_19980);
xnor U22072 (N_22072,N_21861,N_21366);
or U22073 (N_22073,N_20898,N_20337);
nand U22074 (N_22074,N_20458,N_21173);
and U22075 (N_22075,N_19246,N_19567);
nand U22076 (N_22076,N_20356,N_20174);
nor U22077 (N_22077,N_18986,N_20329);
or U22078 (N_22078,N_20106,N_21181);
and U22079 (N_22079,N_18900,N_19593);
nand U22080 (N_22080,N_21440,N_18889);
xnor U22081 (N_22081,N_20609,N_20631);
and U22082 (N_22082,N_19267,N_20543);
or U22083 (N_22083,N_20440,N_20823);
nor U22084 (N_22084,N_19465,N_20444);
nand U22085 (N_22085,N_20026,N_19859);
nor U22086 (N_22086,N_20341,N_20024);
and U22087 (N_22087,N_19642,N_21126);
nor U22088 (N_22088,N_19109,N_20842);
and U22089 (N_22089,N_21619,N_21063);
nand U22090 (N_22090,N_19625,N_21029);
or U22091 (N_22091,N_21800,N_20354);
nor U22092 (N_22092,N_19706,N_18911);
nor U22093 (N_22093,N_20318,N_18882);
nand U22094 (N_22094,N_18992,N_20639);
or U22095 (N_22095,N_21806,N_21857);
nor U22096 (N_22096,N_19437,N_19519);
or U22097 (N_22097,N_21244,N_19951);
and U22098 (N_22098,N_19125,N_19453);
or U22099 (N_22099,N_19984,N_18862);
nor U22100 (N_22100,N_20838,N_20808);
and U22101 (N_22101,N_18801,N_18772);
xnor U22102 (N_22102,N_20067,N_19445);
xnor U22103 (N_22103,N_20668,N_21602);
or U22104 (N_22104,N_21191,N_21176);
xor U22105 (N_22105,N_20175,N_20446);
and U22106 (N_22106,N_21195,N_21626);
nor U22107 (N_22107,N_21710,N_20218);
and U22108 (N_22108,N_19787,N_19666);
or U22109 (N_22109,N_20977,N_20513);
or U22110 (N_22110,N_21863,N_21346);
or U22111 (N_22111,N_19054,N_21264);
nor U22112 (N_22112,N_19199,N_20786);
nor U22113 (N_22113,N_21298,N_19755);
nand U22114 (N_22114,N_21143,N_20715);
nand U22115 (N_22115,N_21167,N_18822);
nand U22116 (N_22116,N_19194,N_21644);
and U22117 (N_22117,N_19175,N_19389);
nand U22118 (N_22118,N_21550,N_21258);
nand U22119 (N_22119,N_19090,N_19688);
or U22120 (N_22120,N_19238,N_20005);
xnor U22121 (N_22121,N_21634,N_18981);
or U22122 (N_22122,N_19424,N_19217);
nor U22123 (N_22123,N_20099,N_19419);
nor U22124 (N_22124,N_19021,N_19546);
and U22125 (N_22125,N_20328,N_19186);
or U22126 (N_22126,N_20982,N_21600);
or U22127 (N_22127,N_19740,N_21119);
nor U22128 (N_22128,N_21528,N_21064);
and U22129 (N_22129,N_20917,N_19405);
and U22130 (N_22130,N_21035,N_21432);
nor U22131 (N_22131,N_20289,N_19382);
nand U22132 (N_22132,N_19652,N_21756);
and U22133 (N_22133,N_19691,N_20107);
xnor U22134 (N_22134,N_18894,N_19128);
or U22135 (N_22135,N_20437,N_19906);
and U22136 (N_22136,N_20241,N_20706);
nor U22137 (N_22137,N_20718,N_20260);
or U22138 (N_22138,N_20023,N_20617);
nand U22139 (N_22139,N_18920,N_20874);
nand U22140 (N_22140,N_19462,N_21378);
or U22141 (N_22141,N_20659,N_20420);
nor U22142 (N_22142,N_20523,N_21539);
and U22143 (N_22143,N_21678,N_21235);
and U22144 (N_22144,N_19776,N_19474);
nor U22145 (N_22145,N_20956,N_20355);
or U22146 (N_22146,N_19739,N_21271);
and U22147 (N_22147,N_21396,N_18961);
and U22148 (N_22148,N_19392,N_20456);
nor U22149 (N_22149,N_21030,N_21370);
nand U22150 (N_22150,N_20368,N_20304);
or U22151 (N_22151,N_20349,N_20041);
nand U22152 (N_22152,N_19817,N_20602);
and U22153 (N_22153,N_21567,N_20847);
or U22154 (N_22154,N_21416,N_21356);
and U22155 (N_22155,N_18924,N_21526);
and U22156 (N_22156,N_19638,N_18950);
and U22157 (N_22157,N_21793,N_21841);
xor U22158 (N_22158,N_20700,N_21517);
nand U22159 (N_22159,N_19222,N_20422);
or U22160 (N_22160,N_19502,N_20683);
or U22161 (N_22161,N_21343,N_19767);
and U22162 (N_22162,N_20431,N_20795);
nor U22163 (N_22163,N_21163,N_21577);
nor U22164 (N_22164,N_21460,N_20656);
and U22165 (N_22165,N_18945,N_18782);
and U22166 (N_22166,N_21694,N_19384);
and U22167 (N_22167,N_20197,N_19493);
nand U22168 (N_22168,N_19401,N_21438);
and U22169 (N_22169,N_19777,N_21372);
nand U22170 (N_22170,N_19883,N_19387);
nand U22171 (N_22171,N_21253,N_19461);
or U22172 (N_22172,N_19543,N_19920);
nor U22173 (N_22173,N_20247,N_19028);
nand U22174 (N_22174,N_21078,N_21802);
or U22175 (N_22175,N_19934,N_19431);
nand U22176 (N_22176,N_19842,N_19942);
or U22177 (N_22177,N_19940,N_21781);
or U22178 (N_22178,N_19622,N_21607);
nor U22179 (N_22179,N_20047,N_19641);
xor U22180 (N_22180,N_21673,N_19952);
and U22181 (N_22181,N_20233,N_19112);
xor U22182 (N_22182,N_20430,N_19468);
nand U22183 (N_22183,N_20862,N_18861);
nor U22184 (N_22184,N_20720,N_18832);
or U22185 (N_22185,N_18893,N_21575);
nand U22186 (N_22186,N_19307,N_20986);
nand U22187 (N_22187,N_20995,N_19492);
or U22188 (N_22188,N_21641,N_18939);
nand U22189 (N_22189,N_21445,N_18867);
nor U22190 (N_22190,N_20916,N_19117);
nor U22191 (N_22191,N_21780,N_20151);
nand U22192 (N_22192,N_21412,N_21207);
xor U22193 (N_22193,N_21079,N_20092);
nor U22194 (N_22194,N_20427,N_20340);
xnor U22195 (N_22195,N_19053,N_21601);
or U22196 (N_22196,N_19114,N_21239);
nand U22197 (N_22197,N_20553,N_21716);
nor U22198 (N_22198,N_20559,N_21263);
xor U22199 (N_22199,N_19602,N_20632);
or U22200 (N_22200,N_21590,N_21845);
and U22201 (N_22201,N_19292,N_21359);
nand U22202 (N_22202,N_21558,N_21854);
xor U22203 (N_22203,N_21819,N_21675);
xnor U22204 (N_22204,N_19825,N_21333);
and U22205 (N_22205,N_19308,N_19300);
or U22206 (N_22206,N_19862,N_20757);
and U22207 (N_22207,N_21357,N_21124);
nor U22208 (N_22208,N_20211,N_19541);
and U22209 (N_22209,N_20054,N_21852);
xnor U22210 (N_22210,N_20091,N_21405);
nand U22211 (N_22211,N_19243,N_19647);
and U22212 (N_22212,N_20296,N_20142);
xnor U22213 (N_22213,N_19857,N_20721);
or U22214 (N_22214,N_19775,N_20680);
or U22215 (N_22215,N_19147,N_19829);
xnor U22216 (N_22216,N_21441,N_19403);
or U22217 (N_22217,N_21425,N_19628);
or U22218 (N_22218,N_20851,N_19873);
nor U22219 (N_22219,N_20132,N_18850);
and U22220 (N_22220,N_21827,N_21160);
or U22221 (N_22221,N_18754,N_20913);
and U22222 (N_22222,N_21241,N_21720);
nor U22223 (N_22223,N_21595,N_19081);
nand U22224 (N_22224,N_19285,N_20192);
or U22225 (N_22225,N_21834,N_21483);
nand U22226 (N_22226,N_19067,N_20028);
nor U22227 (N_22227,N_18775,N_20849);
nor U22228 (N_22228,N_18836,N_20971);
nand U22229 (N_22229,N_20627,N_21453);
or U22230 (N_22230,N_19848,N_19483);
and U22231 (N_22231,N_18937,N_19562);
nor U22232 (N_22232,N_20562,N_20696);
nand U22233 (N_22233,N_20480,N_20373);
nor U22234 (N_22234,N_21227,N_19501);
or U22235 (N_22235,N_21380,N_18814);
or U22236 (N_22236,N_21762,N_19298);
xnor U22237 (N_22237,N_20150,N_20772);
and U22238 (N_22238,N_20630,N_19187);
or U22239 (N_22239,N_18818,N_20841);
or U22240 (N_22240,N_21502,N_20136);
and U22241 (N_22241,N_19773,N_18784);
nor U22242 (N_22242,N_19929,N_20664);
nand U22243 (N_22243,N_21294,N_19997);
or U22244 (N_22244,N_21081,N_20811);
nor U22245 (N_22245,N_20830,N_21536);
nand U22246 (N_22246,N_19827,N_20058);
or U22247 (N_22247,N_21132,N_19573);
or U22248 (N_22248,N_21168,N_20202);
nand U22249 (N_22249,N_21790,N_20729);
nand U22250 (N_22250,N_21511,N_19699);
nand U22251 (N_22251,N_21662,N_19903);
nand U22252 (N_22252,N_20988,N_19785);
or U22253 (N_22253,N_20459,N_19428);
nand U22254 (N_22254,N_19803,N_21186);
xnor U22255 (N_22255,N_21584,N_18892);
nor U22256 (N_22256,N_20145,N_20677);
xnor U22257 (N_22257,N_19703,N_20101);
nor U22258 (N_22258,N_20826,N_20726);
nand U22259 (N_22259,N_21099,N_19271);
xnor U22260 (N_22260,N_20438,N_21713);
nand U22261 (N_22261,N_18988,N_19933);
nor U22262 (N_22262,N_21597,N_19594);
nor U22263 (N_22263,N_21685,N_19436);
xor U22264 (N_22264,N_21820,N_19013);
nand U22265 (N_22265,N_19014,N_20176);
and U22266 (N_22266,N_21796,N_19893);
nand U22267 (N_22267,N_19810,N_20733);
nor U22268 (N_22268,N_19080,N_20086);
or U22269 (N_22269,N_19558,N_21744);
nor U22270 (N_22270,N_19167,N_19811);
xnor U22271 (N_22271,N_18828,N_21809);
nand U22272 (N_22272,N_20079,N_21114);
and U22273 (N_22273,N_19892,N_20518);
or U22274 (N_22274,N_19656,N_20186);
xor U22275 (N_22275,N_19060,N_21547);
or U22276 (N_22276,N_20266,N_20133);
nor U22277 (N_22277,N_21424,N_19870);
nor U22278 (N_22278,N_19357,N_20405);
nand U22279 (N_22279,N_19530,N_21179);
nand U22280 (N_22280,N_19229,N_19705);
nand U22281 (N_22281,N_18970,N_20362);
nand U22282 (N_22282,N_20612,N_21464);
nor U22283 (N_22283,N_19375,N_19113);
nor U22284 (N_22284,N_19910,N_21542);
and U22285 (N_22285,N_19960,N_20646);
and U22286 (N_22286,N_21683,N_19745);
nand U22287 (N_22287,N_20163,N_19002);
and U22288 (N_22288,N_19427,N_19655);
nor U22289 (N_22289,N_21393,N_20781);
nor U22290 (N_22290,N_20039,N_21351);
nor U22291 (N_22291,N_19239,N_21664);
or U22292 (N_22292,N_19108,N_21589);
nor U22293 (N_22293,N_20567,N_21839);
or U22294 (N_22294,N_19993,N_20674);
nor U22295 (N_22295,N_21201,N_21125);
nor U22296 (N_22296,N_21645,N_21169);
and U22297 (N_22297,N_20844,N_18972);
or U22298 (N_22298,N_18990,N_21711);
or U22299 (N_22299,N_21344,N_20081);
nor U22300 (N_22300,N_18901,N_19650);
nand U22301 (N_22301,N_21384,N_20763);
or U22302 (N_22302,N_20794,N_21515);
and U22303 (N_22303,N_20269,N_21817);
nand U22304 (N_22304,N_21133,N_19045);
nor U22305 (N_22305,N_18951,N_21871);
nand U22306 (N_22306,N_19563,N_21007);
and U22307 (N_22307,N_20863,N_21072);
nor U22308 (N_22308,N_21165,N_21382);
and U22309 (N_22309,N_19918,N_21410);
xnor U22310 (N_22310,N_21237,N_19425);
or U22311 (N_22311,N_20206,N_21213);
or U22312 (N_22312,N_19927,N_21571);
nor U22313 (N_22313,N_21325,N_21604);
nand U22314 (N_22314,N_18877,N_20124);
nand U22315 (N_22315,N_21491,N_19446);
nand U22316 (N_22316,N_19302,N_20457);
and U22317 (N_22317,N_21455,N_21418);
and U22318 (N_22318,N_21843,N_20558);
nand U22319 (N_22319,N_19220,N_19976);
or U22320 (N_22320,N_21655,N_19349);
or U22321 (N_22321,N_20875,N_19605);
or U22322 (N_22322,N_19106,N_19459);
xor U22323 (N_22323,N_18985,N_19183);
and U22324 (N_22324,N_19216,N_21653);
or U22325 (N_22325,N_21690,N_19597);
nand U22326 (N_22326,N_19654,N_19990);
or U22327 (N_22327,N_21290,N_20046);
nor U22328 (N_22328,N_19099,N_21482);
xor U22329 (N_22329,N_21219,N_21329);
or U22330 (N_22330,N_21628,N_19399);
and U22331 (N_22331,N_19894,N_19907);
nor U22332 (N_22332,N_20003,N_19010);
nor U22333 (N_22333,N_19634,N_18926);
nand U22334 (N_22334,N_20979,N_21870);
nand U22335 (N_22335,N_21015,N_18834);
xnor U22336 (N_22336,N_20400,N_21408);
and U22337 (N_22337,N_19730,N_20204);
nor U22338 (N_22338,N_20472,N_20970);
nor U22339 (N_22339,N_19510,N_20040);
nand U22340 (N_22340,N_20890,N_18770);
nor U22341 (N_22341,N_20248,N_20539);
or U22342 (N_22342,N_19350,N_19849);
or U22343 (N_22343,N_21578,N_21192);
nand U22344 (N_22344,N_21776,N_19207);
or U22345 (N_22345,N_20933,N_20087);
nand U22346 (N_22346,N_20717,N_20236);
nor U22347 (N_22347,N_19751,N_21332);
nand U22348 (N_22348,N_19410,N_20147);
nand U22349 (N_22349,N_21559,N_19277);
and U22350 (N_22350,N_20376,N_21194);
nor U22351 (N_22351,N_21400,N_21363);
nor U22352 (N_22352,N_19905,N_20942);
and U22353 (N_22353,N_20270,N_20366);
and U22354 (N_22354,N_21723,N_19359);
and U22355 (N_22355,N_20111,N_19571);
nand U22356 (N_22356,N_19390,N_21693);
nor U22357 (N_22357,N_21012,N_19269);
nand U22358 (N_22358,N_18875,N_20695);
nand U22359 (N_22359,N_21315,N_18829);
nand U22360 (N_22360,N_20240,N_20732);
or U22361 (N_22361,N_19630,N_20117);
nor U22362 (N_22362,N_19793,N_20944);
nand U22363 (N_22363,N_19670,N_19011);
nor U22364 (N_22364,N_20239,N_21797);
nand U22365 (N_22365,N_19258,N_20790);
nor U22366 (N_22366,N_20528,N_20178);
nand U22367 (N_22367,N_20980,N_19619);
nor U22368 (N_22368,N_20516,N_20130);
xnor U22369 (N_22369,N_21692,N_20921);
and U22370 (N_22370,N_19592,N_19333);
or U22371 (N_22371,N_19257,N_21795);
nand U22372 (N_22372,N_21118,N_19917);
nand U22373 (N_22373,N_20765,N_20027);
or U22374 (N_22374,N_20914,N_20382);
nor U22375 (N_22375,N_18915,N_20827);
nor U22376 (N_22376,N_19888,N_21274);
nand U22377 (N_22377,N_19441,N_21498);
or U22378 (N_22378,N_20380,N_20287);
or U22379 (N_22379,N_21459,N_19073);
nand U22380 (N_22380,N_19720,N_19416);
xnor U22381 (N_22381,N_20613,N_20850);
nand U22382 (N_22382,N_21611,N_20478);
nor U22383 (N_22383,N_19314,N_19763);
and U22384 (N_22384,N_19059,N_19778);
or U22385 (N_22385,N_20671,N_19844);
nor U22386 (N_22386,N_20766,N_19657);
xnor U22387 (N_22387,N_18904,N_21787);
or U22388 (N_22388,N_20407,N_20564);
and U22389 (N_22389,N_21190,N_21198);
or U22390 (N_22390,N_19454,N_19979);
or U22391 (N_22391,N_20125,N_20712);
and U22392 (N_22392,N_20261,N_21153);
nand U22393 (N_22393,N_19208,N_19851);
or U22394 (N_22394,N_18918,N_21748);
nand U22395 (N_22395,N_20820,N_20663);
and U22396 (N_22396,N_20807,N_20776);
or U22397 (N_22397,N_19725,N_19212);
nand U22398 (N_22398,N_18932,N_21868);
and U22399 (N_22399,N_19430,N_21225);
or U22400 (N_22400,N_19001,N_20482);
xor U22401 (N_22401,N_21051,N_19000);
nand U22402 (N_22402,N_20220,N_20297);
nor U22403 (N_22403,N_20777,N_19760);
xor U22404 (N_22404,N_19343,N_21323);
and U22405 (N_22405,N_19228,N_20300);
nor U22406 (N_22406,N_18899,N_21753);
nor U22407 (N_22407,N_21364,N_20166);
nand U22408 (N_22408,N_19371,N_21221);
or U22409 (N_22409,N_20274,N_19623);
nand U22410 (N_22410,N_19089,N_19473);
xor U22411 (N_22411,N_21269,N_20258);
xnor U22412 (N_22412,N_20083,N_21297);
nand U22413 (N_22413,N_19056,N_20905);
and U22414 (N_22414,N_19598,N_20800);
or U22415 (N_22415,N_20201,N_19818);
or U22416 (N_22416,N_20666,N_21563);
xor U22417 (N_22417,N_20075,N_19123);
and U22418 (N_22418,N_20764,N_19660);
nand U22419 (N_22419,N_20569,N_20744);
nor U22420 (N_22420,N_20925,N_21355);
nand U22421 (N_22421,N_20413,N_19286);
xnor U22422 (N_22422,N_19963,N_19364);
nor U22423 (N_22423,N_19831,N_19752);
xnor U22424 (N_22424,N_20481,N_20620);
and U22425 (N_22425,N_20044,N_19780);
or U22426 (N_22426,N_20774,N_19715);
nand U22427 (N_22427,N_19339,N_19254);
and U22428 (N_22428,N_21286,N_20393);
nand U22429 (N_22429,N_20615,N_19415);
nor U22430 (N_22430,N_21730,N_21087);
or U22431 (N_22431,N_21038,N_20903);
and U22432 (N_22432,N_21452,N_20165);
or U22433 (N_22433,N_19037,N_18979);
and U22434 (N_22434,N_21161,N_21303);
xnor U22435 (N_22435,N_20837,N_21319);
and U22436 (N_22436,N_19981,N_20461);
nand U22437 (N_22437,N_20424,N_21474);
nand U22438 (N_22438,N_21243,N_20590);
nor U22439 (N_22439,N_20008,N_21444);
xor U22440 (N_22440,N_21679,N_19182);
nand U22441 (N_22441,N_19753,N_20487);
nand U22442 (N_22442,N_20503,N_18927);
nand U22443 (N_22443,N_20309,N_21810);
and U22444 (N_22444,N_21499,N_20237);
nand U22445 (N_22445,N_19983,N_21032);
and U22446 (N_22446,N_19926,N_20751);
nand U22447 (N_22447,N_21105,N_21866);
and U22448 (N_22448,N_19855,N_19640);
nor U22449 (N_22449,N_18845,N_19276);
and U22450 (N_22450,N_19148,N_19886);
and U22451 (N_22451,N_21122,N_20149);
nor U22452 (N_22452,N_21157,N_21596);
nand U22453 (N_22453,N_19872,N_21745);
and U22454 (N_22454,N_21000,N_20622);
nor U22455 (N_22455,N_20148,N_21461);
or U22456 (N_22456,N_18769,N_21174);
or U22457 (N_22457,N_21500,N_19781);
nand U22458 (N_22458,N_19841,N_20860);
nor U22459 (N_22459,N_20451,N_20596);
or U22460 (N_22460,N_20552,N_21260);
and U22461 (N_22461,N_20623,N_20897);
or U22462 (N_22462,N_20814,N_18812);
nand U22463 (N_22463,N_21622,N_20941);
nor U22464 (N_22464,N_21472,N_20158);
or U22465 (N_22465,N_19505,N_21492);
and U22466 (N_22466,N_21120,N_19673);
or U22467 (N_22467,N_18902,N_19448);
or U22468 (N_22468,N_21651,N_19606);
or U22469 (N_22469,N_19704,N_19400);
xor U22470 (N_22470,N_21470,N_19627);
and U22471 (N_22471,N_21223,N_20818);
nand U22472 (N_22472,N_18987,N_20162);
nand U22473 (N_22473,N_19388,N_21496);
nand U22474 (N_22474,N_20924,N_20471);
and U22475 (N_22475,N_21458,N_21200);
nor U22476 (N_22476,N_20967,N_21831);
nand U22477 (N_22477,N_20638,N_19999);
and U22478 (N_22478,N_21305,N_20595);
or U22479 (N_22479,N_20200,N_21605);
and U22480 (N_22480,N_20938,N_19305);
and U22481 (N_22481,N_21534,N_20169);
or U22482 (N_22482,N_20143,N_19850);
or U22483 (N_22483,N_20189,N_19118);
and U22484 (N_22484,N_19885,N_19177);
nand U22485 (N_22485,N_20722,N_21621);
or U22486 (N_22486,N_21615,N_18955);
or U22487 (N_22487,N_21149,N_19452);
and U22488 (N_22488,N_21273,N_19735);
and U22489 (N_22489,N_21624,N_20742);
and U22490 (N_22490,N_19135,N_18864);
or U22491 (N_22491,N_19618,N_20030);
and U22492 (N_22492,N_19794,N_20377);
or U22493 (N_22493,N_20339,N_19131);
and U22494 (N_22494,N_21646,N_19347);
nor U22495 (N_22495,N_21299,N_19294);
nand U22496 (N_22496,N_20525,N_20080);
nand U22497 (N_22497,N_21117,N_19139);
nor U22498 (N_22498,N_19435,N_19762);
or U22499 (N_22499,N_19418,N_20998);
nand U22500 (N_22500,N_20002,N_19322);
and U22501 (N_22501,N_20398,N_19015);
xnor U22502 (N_22502,N_20885,N_20502);
xnor U22503 (N_22503,N_21080,N_19684);
or U22504 (N_22504,N_20346,N_21648);
or U22505 (N_22505,N_19413,N_19456);
nand U22506 (N_22506,N_20517,N_20689);
nand U22507 (N_22507,N_19909,N_19998);
nor U22508 (N_22508,N_20050,N_20952);
or U22509 (N_22509,N_19991,N_19262);
nand U22510 (N_22510,N_20114,N_19363);
nand U22511 (N_22511,N_19692,N_19409);
or U22512 (N_22512,N_19092,N_21468);
nor U22513 (N_22513,N_19749,N_21643);
nand U22514 (N_22514,N_21422,N_20853);
or U22515 (N_22515,N_20535,N_20743);
and U22516 (N_22516,N_20466,N_19525);
xnor U22517 (N_22517,N_19680,N_21285);
and U22518 (N_22518,N_21415,N_19754);
nand U22519 (N_22519,N_19129,N_19921);
and U22520 (N_22520,N_21856,N_21777);
and U22521 (N_22521,N_18761,N_20592);
nand U22522 (N_22522,N_20037,N_19497);
nor U22523 (N_22523,N_19540,N_20597);
nand U22524 (N_22524,N_20691,N_20824);
nor U22525 (N_22525,N_19615,N_19936);
or U22526 (N_22526,N_18773,N_18957);
nor U22527 (N_22527,N_21636,N_20259);
nor U22528 (N_22528,N_21089,N_20390);
or U22529 (N_22529,N_19423,N_18942);
nand U22530 (N_22530,N_20548,N_21844);
nand U22531 (N_22531,N_21603,N_18794);
nor U22532 (N_22532,N_20470,N_19233);
or U22533 (N_22533,N_18880,N_19898);
or U22534 (N_22534,N_20187,N_20652);
or U22535 (N_22535,N_21572,N_20812);
and U22536 (N_22536,N_20880,N_21021);
or U22537 (N_22537,N_20604,N_19681);
nor U22538 (N_22538,N_20761,N_19696);
or U22539 (N_22539,N_20484,N_19897);
nand U22540 (N_22540,N_19596,N_20937);
and U22541 (N_22541,N_21449,N_21538);
or U22542 (N_22542,N_20272,N_19935);
nor U22543 (N_22543,N_19144,N_20688);
nand U22544 (N_22544,N_19729,N_19858);
nor U22545 (N_22545,N_20217,N_19678);
nor U22546 (N_22546,N_21501,N_19162);
and U22547 (N_22547,N_21292,N_20670);
and U22548 (N_22548,N_21707,N_19973);
nor U22549 (N_22549,N_20650,N_20230);
nand U22550 (N_22550,N_19155,N_21371);
xnor U22551 (N_22551,N_19378,N_20320);
nand U22552 (N_22552,N_20386,N_21524);
nor U22553 (N_22553,N_20434,N_19007);
nand U22554 (N_22554,N_20780,N_20994);
and U22555 (N_22555,N_20372,N_20990);
nor U22556 (N_22556,N_19737,N_19355);
xor U22557 (N_22557,N_21001,N_19901);
nand U22558 (N_22558,N_21342,N_21101);
or U22559 (N_22559,N_19578,N_20344);
nor U22560 (N_22560,N_20408,N_21652);
nor U22561 (N_22561,N_20419,N_18984);
nand U22562 (N_22562,N_21082,N_21135);
and U22563 (N_22563,N_19444,N_18820);
and U22564 (N_22564,N_19969,N_19464);
xnor U22565 (N_22565,N_20433,N_19458);
or U22566 (N_22566,N_20181,N_19457);
or U22567 (N_22567,N_20858,N_21684);
or U22568 (N_22568,N_19316,N_19561);
nor U22569 (N_22569,N_20499,N_20188);
nand U22570 (N_22570,N_18795,N_20699);
nor U22571 (N_22571,N_19697,N_19694);
and U22572 (N_22572,N_21768,N_19805);
nand U22573 (N_22573,N_19856,N_20973);
or U22574 (N_22574,N_21687,N_18865);
nand U22575 (N_22575,N_21674,N_21654);
nor U22576 (N_22576,N_19515,N_21262);
and U22577 (N_22577,N_20322,N_20810);
nand U22578 (N_22578,N_19514,N_19985);
nand U22579 (N_22579,N_20739,N_20127);
nor U22580 (N_22580,N_21044,N_20262);
nor U22581 (N_22581,N_20275,N_20658);
nor U22582 (N_22582,N_19726,N_21721);
or U22583 (N_22583,N_20196,N_21838);
and U22584 (N_22584,N_21490,N_21248);
and U22585 (N_22585,N_19255,N_20996);
nor U22586 (N_22586,N_21738,N_19227);
nand U22587 (N_22587,N_21743,N_20032);
or U22588 (N_22588,N_19471,N_19304);
nor U22589 (N_22589,N_21588,N_21193);
xor U22590 (N_22590,N_20835,N_20969);
and U22591 (N_22591,N_20126,N_20511);
nor U22592 (N_22592,N_19420,N_20038);
or U22593 (N_22593,N_19764,N_20168);
nand U22594 (N_22594,N_19932,N_21004);
nand U22595 (N_22595,N_18798,N_18922);
nand U22596 (N_22596,N_19782,N_20611);
nor U22597 (N_22597,N_19226,N_20006);
nand U22598 (N_22598,N_20435,N_19904);
nor U22599 (N_22599,N_19104,N_21495);
nand U22600 (N_22600,N_18810,N_21368);
and U22601 (N_22601,N_20042,N_21735);
or U22602 (N_22602,N_21277,N_19499);
or U22603 (N_22603,N_18866,N_19679);
nor U22604 (N_22604,N_20265,N_21494);
nor U22605 (N_22605,N_18817,N_20301);
nor U22606 (N_22606,N_20394,N_21148);
or U22607 (N_22607,N_19830,N_20532);
nor U22608 (N_22608,N_19311,N_18756);
nand U22609 (N_22609,N_21656,N_20141);
nor U22610 (N_22610,N_19865,N_20093);
nand U22611 (N_22611,N_19946,N_19283);
and U22612 (N_22612,N_19025,N_21180);
nand U22613 (N_22613,N_19861,N_19911);
nor U22614 (N_22614,N_21024,N_20526);
nand U22615 (N_22615,N_19624,N_20804);
or U22616 (N_22616,N_19923,N_19769);
or U22617 (N_22617,N_21616,N_21252);
nor U22618 (N_22618,N_21807,N_20234);
and U22619 (N_22619,N_21331,N_20974);
and U22620 (N_22620,N_21111,N_20053);
or U22621 (N_22621,N_19432,N_21689);
xor U22622 (N_22622,N_21379,N_20908);
xor U22623 (N_22623,N_20940,N_19801);
or U22624 (N_22624,N_19955,N_21336);
and U22625 (N_22625,N_20180,N_20161);
and U22626 (N_22626,N_19663,N_21255);
or U22627 (N_22627,N_20822,N_19224);
or U22628 (N_22628,N_19644,N_19667);
nand U22629 (N_22629,N_21229,N_19658);
nand U22630 (N_22630,N_19535,N_21847);
and U22631 (N_22631,N_19839,N_21138);
nand U22632 (N_22632,N_19565,N_19518);
xor U22633 (N_22633,N_20001,N_21310);
nand U22634 (N_22634,N_19610,N_20846);
nor U22635 (N_22635,N_20064,N_19172);
or U22636 (N_22636,N_19101,N_19051);
or U22637 (N_22637,N_20227,N_19908);
or U22638 (N_22638,N_20283,N_19672);
and U22639 (N_22639,N_19093,N_20877);
and U22640 (N_22640,N_20264,N_19576);
or U22641 (N_22641,N_19486,N_20782);
xnor U22642 (N_22642,N_20374,N_18760);
or U22643 (N_22643,N_20796,N_21583);
or U22644 (N_22644,N_19306,N_21700);
or U22645 (N_22645,N_21579,N_19823);
and U22646 (N_22646,N_20257,N_20244);
xor U22647 (N_22647,N_21060,N_20687);
nand U22648 (N_22648,N_21216,N_20448);
or U22649 (N_22649,N_18807,N_21272);
and U22650 (N_22650,N_19813,N_19736);
or U22651 (N_22651,N_21508,N_21510);
nor U22652 (N_22652,N_21113,N_21865);
xor U22653 (N_22653,N_20740,N_20789);
xor U22654 (N_22654,N_19358,N_20153);
xnor U22655 (N_22655,N_18941,N_21236);
nor U22656 (N_22656,N_19689,N_19724);
nand U22657 (N_22657,N_19833,N_19373);
xnor U22658 (N_22658,N_21151,N_21521);
nor U22659 (N_22659,N_19900,N_20738);
nor U22660 (N_22660,N_20473,N_21394);
and U22661 (N_22661,N_19916,N_18870);
and U22662 (N_22662,N_21677,N_20778);
and U22663 (N_22663,N_21043,N_20936);
nand U22664 (N_22664,N_18874,N_20488);
and U22665 (N_22665,N_18916,N_21048);
nand U22666 (N_22666,N_20866,N_18934);
or U22667 (N_22667,N_20624,N_19838);
nand U22668 (N_22668,N_20867,N_21002);
and U22669 (N_22669,N_20049,N_18750);
or U22670 (N_22670,N_19232,N_20616);
nor U22671 (N_22671,N_19075,N_20159);
nand U22672 (N_22672,N_20984,N_21701);
nor U22673 (N_22673,N_18923,N_19728);
or U22674 (N_22674,N_20395,N_19041);
nand U22675 (N_22675,N_20330,N_20570);
and U22676 (N_22676,N_21755,N_20068);
xnor U22677 (N_22677,N_19609,N_21185);
and U22678 (N_22678,N_21123,N_21477);
or U22679 (N_22679,N_19245,N_19531);
nand U22680 (N_22680,N_21096,N_19127);
xnor U22681 (N_22681,N_19564,N_20857);
nand U22682 (N_22682,N_21763,N_20584);
and U22683 (N_22683,N_19433,N_21367);
and U22684 (N_22684,N_19038,N_21085);
or U22685 (N_22685,N_21373,N_21484);
xor U22686 (N_22686,N_21821,N_21417);
xnor U22687 (N_22687,N_19632,N_20504);
nor U22688 (N_22688,N_21166,N_19949);
nand U22689 (N_22689,N_20993,N_21594);
nor U22690 (N_22690,N_20768,N_21722);
and U22691 (N_22691,N_18837,N_20336);
and U22692 (N_22692,N_18999,N_20649);
xnor U22693 (N_22693,N_21092,N_21544);
nand U22694 (N_22694,N_21708,N_18847);
xnor U22695 (N_22695,N_20886,N_18826);
nor U22696 (N_22696,N_19806,N_19891);
or U22697 (N_22697,N_21465,N_20363);
or U22698 (N_22698,N_19024,N_20493);
xnor U22699 (N_22699,N_19334,N_20098);
and U22700 (N_22700,N_20411,N_19261);
and U22701 (N_22701,N_21341,N_20369);
xnor U22702 (N_22702,N_20983,N_19522);
nand U22703 (N_22703,N_20191,N_18813);
or U22704 (N_22704,N_21115,N_19837);
and U22705 (N_22705,N_18789,N_19326);
nor U22706 (N_22706,N_18779,N_19930);
nand U22707 (N_22707,N_21519,N_21347);
and U22708 (N_22708,N_21514,N_21187);
nor U22709 (N_22709,N_18852,N_19482);
nand U22710 (N_22710,N_20072,N_21280);
nor U22711 (N_22711,N_20276,N_20642);
xnor U22712 (N_22712,N_21265,N_21862);
or U22713 (N_22713,N_20496,N_19800);
nand U22714 (N_22714,N_19557,N_21598);
or U22715 (N_22715,N_19270,N_21696);
nand U22716 (N_22716,N_19757,N_21717);
xor U22717 (N_22717,N_19568,N_21632);
xor U22718 (N_22718,N_20279,N_20601);
nor U22719 (N_22719,N_20011,N_20762);
nor U22720 (N_22720,N_21251,N_20878);
nor U22721 (N_22721,N_19103,N_20134);
nor U22722 (N_22722,N_18856,N_19160);
nand U22723 (N_22723,N_19820,N_20112);
or U22724 (N_22724,N_20636,N_19868);
nor U22725 (N_22725,N_19487,N_19653);
and U22726 (N_22726,N_20934,N_21150);
nand U22727 (N_22727,N_19821,N_20935);
nor U22728 (N_22728,N_20542,N_20213);
xnor U22729 (N_22729,N_20865,N_21614);
nand U22730 (N_22730,N_19386,N_21016);
nand U22731 (N_22731,N_21549,N_20225);
or U22732 (N_22732,N_18806,N_18777);
nor U22733 (N_22733,N_21867,N_20524);
and U22734 (N_22734,N_20370,N_20549);
nand U22735 (N_22735,N_19600,N_18958);
or U22736 (N_22736,N_19712,N_20754);
xor U22737 (N_22737,N_21537,N_20209);
nand U22738 (N_22738,N_20704,N_18765);
or U22739 (N_22739,N_21312,N_19068);
nor U22740 (N_22740,N_21749,N_20899);
nor U22741 (N_22741,N_20788,N_18787);
or U22742 (N_22742,N_20073,N_20494);
nor U22743 (N_22743,N_18948,N_19582);
nor U22744 (N_22744,N_19323,N_18935);
or U22745 (N_22745,N_19337,N_19693);
xor U22746 (N_22746,N_20640,N_20932);
and U22747 (N_22747,N_19044,N_20563);
and U22748 (N_22748,N_19747,N_19361);
nand U22749 (N_22749,N_21860,N_19717);
and U22750 (N_22750,N_19153,N_21480);
xor U22751 (N_22751,N_19937,N_19899);
or U22752 (N_22752,N_20651,N_21046);
nand U22753 (N_22753,N_20945,N_18823);
nand U22754 (N_22754,N_21561,N_20910);
nand U22755 (N_22755,N_18995,N_19700);
nor U22756 (N_22756,N_20278,N_20074);
nand U22757 (N_22757,N_19477,N_21172);
xnor U22758 (N_22758,N_19408,N_20443);
and U22759 (N_22759,N_20775,N_21155);
or U22760 (N_22760,N_20308,N_21554);
nand U22761 (N_22761,N_19273,N_19521);
nand U22762 (N_22762,N_21010,N_19031);
or U22763 (N_22763,N_20669,N_19366);
or U22764 (N_22764,N_21387,N_21576);
or U22765 (N_22765,N_20009,N_21300);
nor U22766 (N_22766,N_20182,N_19249);
nor U22767 (N_22767,N_19341,N_20397);
and U22768 (N_22768,N_18917,N_18799);
nand U22769 (N_22769,N_21798,N_21146);
nand U22770 (N_22770,N_19284,N_20939);
or U22771 (N_22771,N_19520,N_19132);
or U22772 (N_22772,N_21503,N_21513);
nor U22773 (N_22773,N_21233,N_20170);
nand U22774 (N_22774,N_20273,N_19890);
nand U22775 (N_22775,N_21587,N_19577);
nand U22776 (N_22776,N_20705,N_19039);
xor U22777 (N_22777,N_21075,N_20960);
or U22778 (N_22778,N_19524,N_19840);
and U22779 (N_22779,N_21427,N_21775);
or U22780 (N_22780,N_19896,N_21430);
nor U22781 (N_22781,N_19225,N_20883);
or U22782 (N_22782,N_18967,N_21740);
nor U22783 (N_22783,N_20869,N_19180);
nor U22784 (N_22784,N_21314,N_20212);
nor U22785 (N_22785,N_18946,N_21330);
and U22786 (N_22786,N_19133,N_20951);
and U22787 (N_22787,N_20312,N_19864);
or U22788 (N_22788,N_21580,N_20736);
or U22789 (N_22789,N_20000,N_18963);
nor U22790 (N_22790,N_21836,N_21204);
or U22791 (N_22791,N_19476,N_21406);
nand U22792 (N_22792,N_20545,N_20965);
and U22793 (N_22793,N_20538,N_21608);
and U22794 (N_22794,N_18910,N_18759);
xnor U22795 (N_22795,N_18755,N_19553);
nand U22796 (N_22796,N_21147,N_19881);
nor U22797 (N_22797,N_19197,N_19591);
nor U22798 (N_22798,N_18978,N_20621);
or U22799 (N_22799,N_21404,N_19544);
or U22800 (N_22800,N_20034,N_20966);
nor U22801 (N_22801,N_18977,N_20334);
nand U22802 (N_22802,N_20576,N_20876);
and U22803 (N_22803,N_18888,N_19798);
or U22804 (N_22804,N_20389,N_19549);
nor U22805 (N_22805,N_19005,N_21760);
nor U22806 (N_22806,N_21849,N_20896);
nor U22807 (N_22807,N_21788,N_21056);
and U22808 (N_22808,N_21025,N_19033);
nand U22809 (N_22809,N_19948,N_21413);
and U22810 (N_22810,N_18891,N_20118);
and U22811 (N_22811,N_21725,N_21727);
nand U22812 (N_22812,N_20600,N_19071);
nand U22813 (N_22813,N_20871,N_21128);
or U22814 (N_22814,N_19614,N_19018);
and U22815 (N_22815,N_21516,N_20271);
xnor U22816 (N_22816,N_21098,N_19248);
xnor U22817 (N_22817,N_19633,N_19612);
and U22818 (N_22818,N_19052,N_19391);
or U22819 (N_22819,N_20879,N_20070);
or U22820 (N_22820,N_21736,N_20805);
xor U22821 (N_22821,N_19668,N_19141);
xor U22822 (N_22822,N_21451,N_21361);
and U22823 (N_22823,N_21670,N_18849);
and U22824 (N_22824,N_20282,N_20291);
or U22825 (N_22825,N_21864,N_20872);
nor U22826 (N_22826,N_19190,N_20226);
and U22827 (N_22827,N_20173,N_19161);
nor U22828 (N_22828,N_20964,N_20520);
nand U22829 (N_22829,N_21212,N_20684);
or U22830 (N_22830,N_20164,N_19062);
nor U22831 (N_22831,N_21052,N_19727);
and U22832 (N_22832,N_21279,N_20110);
or U22833 (N_22833,N_21401,N_20537);
nor U22834 (N_22834,N_21709,N_19746);
nor U22835 (N_22835,N_20065,N_21489);
nor U22836 (N_22836,N_21822,N_18851);
nor U22837 (N_22837,N_20978,N_18921);
nor U22838 (N_22838,N_20295,N_21222);
or U22839 (N_22839,N_20156,N_21818);
and U22840 (N_22840,N_21556,N_19301);
nand U22841 (N_22841,N_19707,N_19765);
or U22842 (N_22842,N_19383,N_20105);
nor U22843 (N_22843,N_20661,N_18940);
nand U22844 (N_22844,N_19235,N_20540);
nand U22845 (N_22845,N_21804,N_21183);
and U22846 (N_22846,N_20679,N_21533);
or U22847 (N_22847,N_20922,N_21507);
nand U22848 (N_22848,N_21774,N_19057);
and U22849 (N_22849,N_21093,N_20946);
xnor U22850 (N_22850,N_20453,N_19875);
nor U22851 (N_22851,N_19569,N_20583);
or U22852 (N_22852,N_21545,N_20231);
nand U22853 (N_22853,N_21091,N_18855);
or U22854 (N_22854,N_18804,N_19353);
or U22855 (N_22855,N_19956,N_21627);
nor U22856 (N_22856,N_20325,N_19395);
and U22857 (N_22857,N_18906,N_21869);
and U22858 (N_22858,N_19096,N_19442);
and U22859 (N_22859,N_20333,N_19130);
nor U22860 (N_22860,N_19485,N_19209);
nor U22861 (N_22861,N_19214,N_19231);
and U22862 (N_22862,N_21737,N_21094);
and U22863 (N_22863,N_18936,N_21308);
nor U22864 (N_22864,N_20014,N_18887);
nand U22865 (N_22865,N_19581,N_20228);
and U22866 (N_22866,N_19398,N_21436);
nor U22867 (N_22867,N_20725,N_21145);
xor U22868 (N_22868,N_20031,N_19069);
xnor U22869 (N_22869,N_19206,N_21217);
or U22870 (N_22870,N_20235,N_18808);
or U22871 (N_22871,N_21090,N_21073);
or U22872 (N_22872,N_21606,N_20888);
nor U22873 (N_22873,N_21270,N_19396);
or U22874 (N_22874,N_21320,N_20521);
or U22875 (N_22875,N_19802,N_19617);
and U22876 (N_22876,N_19169,N_21419);
and U22877 (N_22877,N_19377,N_20409);
and U22878 (N_22878,N_18881,N_21061);
nor U22879 (N_22879,N_20834,N_19095);
xor U22880 (N_22880,N_19381,N_20606);
or U22881 (N_22881,N_19369,N_20013);
or U22882 (N_22882,N_21397,N_19017);
and U22883 (N_22883,N_20654,N_20462);
and U22884 (N_22884,N_19019,N_21246);
nor U22885 (N_22885,N_21008,N_19211);
nor U22886 (N_22886,N_19219,N_19178);
nor U22887 (N_22887,N_21564,N_21757);
nand U22888 (N_22888,N_20603,N_19244);
and U22889 (N_22889,N_19438,N_18859);
nand U22890 (N_22890,N_18949,N_19356);
xor U22891 (N_22891,N_20832,N_20392);
and U22892 (N_22892,N_20641,N_21703);
or U22893 (N_22893,N_20097,N_19236);
nand U22894 (N_22894,N_19480,N_19958);
nand U22895 (N_22895,N_20625,N_19250);
and U22896 (N_22896,N_20585,N_19050);
and U22897 (N_22897,N_21669,N_18998);
xor U22898 (N_22898,N_20012,N_19105);
and U22899 (N_22899,N_19978,N_20950);
xor U22900 (N_22900,N_20281,N_20634);
nor U22901 (N_22901,N_20856,N_19506);
or U22902 (N_22902,N_20324,N_18811);
nand U22903 (N_22903,N_19662,N_20598);
nor U22904 (N_22904,N_19185,N_20285);
xor U22905 (N_22905,N_18780,N_20135);
nor U22906 (N_22906,N_20256,N_21794);
nor U22907 (N_22907,N_19164,N_21266);
and U22908 (N_22908,N_21581,N_19537);
nor U22909 (N_22909,N_19256,N_20727);
nor U22910 (N_22910,N_21829,N_19539);
nor U22911 (N_22911,N_20500,N_19121);
nor U22912 (N_22912,N_21289,N_19742);
xnor U22913 (N_22913,N_21658,N_21196);
nor U22914 (N_22914,N_19809,N_19912);
or U22915 (N_22915,N_20250,N_19816);
nor U22916 (N_22916,N_19297,N_19223);
nor U22917 (N_22917,N_20571,N_21283);
and U22918 (N_22918,N_19547,N_21142);
nand U22919 (N_22919,N_19120,N_21084);
nand U22920 (N_22920,N_20184,N_19533);
or U22921 (N_22921,N_21629,N_20579);
and U22922 (N_22922,N_20069,N_18898);
or U22923 (N_22923,N_19977,N_19221);
nor U22924 (N_22924,N_19083,N_20302);
or U22925 (N_22925,N_21506,N_20423);
or U22926 (N_22926,N_21754,N_20560);
xnor U22927 (N_22927,N_19972,N_19772);
nor U22928 (N_22928,N_19079,N_21074);
nor U22929 (N_22929,N_21457,N_20185);
nor U22930 (N_22930,N_20345,N_19496);
and U22931 (N_22931,N_21824,N_18873);
and U22932 (N_22932,N_18843,N_19555);
or U22933 (N_22933,N_21170,N_18953);
and U22934 (N_22934,N_19860,N_19078);
and U22935 (N_22935,N_21317,N_21712);
and U22936 (N_22936,N_20575,N_19030);
nand U22937 (N_22937,N_21013,N_20895);
or U22938 (N_22938,N_20035,N_21792);
or U22939 (N_22939,N_21045,N_20507);
or U22940 (N_22940,N_20215,N_20305);
nor U22941 (N_22941,N_21058,N_20817);
and U22942 (N_22942,N_20450,N_20280);
nand U22943 (N_22943,N_21640,N_19303);
and U22944 (N_22944,N_20724,N_20852);
or U22945 (N_22945,N_21377,N_19887);
nand U22946 (N_22946,N_21803,N_19295);
and U22947 (N_22947,N_19770,N_20992);
or U22948 (N_22948,N_21083,N_20635);
nand U22949 (N_22949,N_20770,N_20221);
nor U22950 (N_22950,N_19417,N_18878);
xnor U22951 (N_22951,N_21141,N_21295);
nand U22952 (N_22952,N_19205,N_20063);
nor U22953 (N_22953,N_19346,N_20317);
nand U22954 (N_22954,N_19061,N_20884);
or U22955 (N_22955,N_20315,N_18996);
xor U22956 (N_22956,N_20183,N_19251);
or U22957 (N_22957,N_20864,N_20955);
nor U22958 (N_22958,N_19040,N_19362);
nand U22959 (N_22959,N_18751,N_19397);
nor U22960 (N_22960,N_21033,N_20614);
nand U22961 (N_22961,N_19607,N_18890);
xnor U22962 (N_22962,N_20358,N_21345);
nand U22963 (N_22963,N_20402,N_21620);
and U22964 (N_22964,N_19370,N_18767);
or U22965 (N_22965,N_21403,N_20019);
or U22966 (N_22966,N_21383,N_18793);
nand U22967 (N_22967,N_21159,N_18857);
nand U22968 (N_22968,N_19324,N_20594);
or U22969 (N_22969,N_18980,N_19020);
nor U22970 (N_22970,N_20882,N_20702);
nand U22971 (N_22971,N_20243,N_19196);
or U22972 (N_22972,N_20755,N_21732);
or U22973 (N_22973,N_20404,N_20321);
nand U22974 (N_22974,N_18993,N_20784);
and U22975 (N_22975,N_20104,N_20985);
nor U22976 (N_22976,N_19784,N_21386);
nand U22977 (N_22977,N_19500,N_20906);
nor U22978 (N_22978,N_20022,N_19137);
or U22979 (N_22979,N_19463,N_19532);
and U22980 (N_22980,N_20246,N_21034);
and U22981 (N_22981,N_20673,N_21773);
and U22982 (N_22982,N_20647,N_21715);
xor U22983 (N_22983,N_21456,N_20310);
or U22984 (N_22984,N_21770,N_21365);
xnor U22985 (N_22985,N_21486,N_19143);
and U22986 (N_22986,N_19913,N_20495);
or U22987 (N_22987,N_21328,N_20949);
xor U22988 (N_22988,N_20682,N_19768);
xor U22989 (N_22989,N_19289,N_19536);
nand U22990 (N_22990,N_18824,N_19516);
xnor U22991 (N_22991,N_20991,N_18776);
nor U22992 (N_22992,N_19274,N_20205);
and U22993 (N_22993,N_19288,N_20508);
or U22994 (N_22994,N_21177,N_21238);
nor U22995 (N_22995,N_20084,N_20077);
nand U22996 (N_22996,N_21095,N_19494);
and U22997 (N_22997,N_21463,N_18758);
and U22998 (N_22998,N_19188,N_19877);
or U22999 (N_22999,N_21532,N_20809);
and U23000 (N_23000,N_20968,N_21431);
nand U23001 (N_23001,N_18819,N_21287);
nor U23002 (N_23002,N_21493,N_19042);
nand U23003 (N_23003,N_19852,N_19440);
nand U23004 (N_23004,N_20445,N_21828);
nor U23005 (N_23005,N_21375,N_19282);
xor U23006 (N_23006,N_21014,N_20415);
and U23007 (N_23007,N_21479,N_21471);
nand U23008 (N_23008,N_20901,N_18938);
xnor U23009 (N_23009,N_21208,N_21374);
nand U23010 (N_23010,N_19924,N_20057);
and U23011 (N_23011,N_21291,N_19922);
nor U23012 (N_23012,N_20843,N_19152);
nor U23013 (N_23013,N_18792,N_21031);
xnor U23014 (N_23014,N_19004,N_21599);
xor U23015 (N_23015,N_21335,N_20190);
and U23016 (N_23016,N_19489,N_19950);
or U23017 (N_23017,N_19215,N_21178);
or U23018 (N_23018,N_19545,N_20581);
nand U23019 (N_23019,N_21391,N_21022);
or U23020 (N_23020,N_21420,N_19714);
or U23021 (N_23021,N_20323,N_20157);
nand U23022 (N_23022,N_19006,N_19970);
or U23023 (N_23023,N_19566,N_19719);
nor U23024 (N_23024,N_20036,N_18842);
nor U23025 (N_23025,N_21301,N_19077);
nor U23026 (N_23026,N_20378,N_21541);
nand U23027 (N_23027,N_18796,N_20179);
nand U23028 (N_23028,N_19171,N_21573);
and U23029 (N_23029,N_20388,N_21261);
nor U23030 (N_23030,N_20144,N_19645);
or U23031 (N_23031,N_19268,N_19281);
xnor U23032 (N_23032,N_20383,N_20633);
nand U23033 (N_23033,N_21293,N_18903);
nand U23034 (N_23034,N_20816,N_21448);
nor U23035 (N_23035,N_21816,N_19016);
xnor U23036 (N_23036,N_21267,N_19791);
nor U23037 (N_23037,N_19902,N_18968);
and U23038 (N_23038,N_19783,N_18885);
nor U23039 (N_23039,N_20629,N_20657);
nor U23040 (N_23040,N_20467,N_20045);
and U23041 (N_23041,N_19156,N_20943);
nor U23042 (N_23042,N_18991,N_20672);
nor U23043 (N_23043,N_18854,N_20311);
or U23044 (N_23044,N_18971,N_21435);
xnor U23045 (N_23045,N_21752,N_19029);
nand U23046 (N_23046,N_19204,N_20335);
or U23047 (N_23047,N_19470,N_20655);
or U23048 (N_23048,N_21568,N_19682);
nand U23049 (N_23049,N_20103,N_18944);
or U23050 (N_23050,N_19154,N_19335);
xor U23051 (N_23051,N_20662,N_19299);
nand U23052 (N_23052,N_21691,N_21003);
and U23053 (N_23053,N_19931,N_20561);
and U23054 (N_23054,N_20587,N_19992);
nor U23055 (N_23055,N_19572,N_19145);
and U23056 (N_23056,N_21276,N_20061);
nor U23057 (N_23057,N_20326,N_20116);
nor U23058 (N_23058,N_19939,N_19675);
and U23059 (N_23059,N_19799,N_21121);
nand U23060 (N_23060,N_20573,N_21661);
nor U23061 (N_23061,N_20286,N_19845);
and U23062 (N_23062,N_21872,N_19351);
and U23063 (N_23063,N_21742,N_20004);
nand U23064 (N_23064,N_20541,N_21103);
and U23065 (N_23065,N_20577,N_20338);
nand U23066 (N_23066,N_19876,N_19964);
and U23067 (N_23067,N_20904,N_19166);
or U23068 (N_23068,N_21766,N_19455);
or U23069 (N_23069,N_18753,N_18848);
nand U23070 (N_23070,N_19404,N_20565);
nor U23071 (N_23071,N_21609,N_19914);
nand U23072 (N_23072,N_21688,N_20442);
nand U23073 (N_23073,N_20848,N_20082);
or U23074 (N_23074,N_20327,N_21657);
or U23075 (N_23075,N_20303,N_21011);
and U23076 (N_23076,N_21395,N_20931);
or U23077 (N_23077,N_21210,N_18783);
nand U23078 (N_23078,N_21037,N_19312);
and U23079 (N_23079,N_19043,N_21837);
xor U23080 (N_23080,N_19702,N_19635);
nand U23081 (N_23081,N_20746,N_20547);
nor U23082 (N_23082,N_19275,N_21350);
nor U23083 (N_23083,N_20840,N_19559);
nand U23084 (N_23084,N_20529,N_21230);
or U23085 (N_23085,N_20515,N_18994);
nor U23086 (N_23086,N_20489,N_19585);
nand U23087 (N_23087,N_21340,N_21108);
and U23088 (N_23088,N_19111,N_19163);
and U23089 (N_23089,N_20501,N_19943);
nor U23090 (N_23090,N_21569,N_18952);
xor U23091 (N_23091,N_20927,N_19342);
nor U23092 (N_23092,N_21548,N_19986);
nor U23093 (N_23093,N_20171,N_19824);
or U23094 (N_23094,N_19264,N_20586);
xor U23095 (N_23095,N_19331,N_19836);
and U23096 (N_23096,N_21224,N_21348);
nor U23097 (N_23097,N_20618,N_20918);
or U23098 (N_23098,N_19620,N_20412);
nor U23099 (N_23099,N_18956,N_19774);
nand U23100 (N_23100,N_21842,N_18913);
or U23101 (N_23101,N_21257,N_19189);
nand U23102 (N_23102,N_20833,N_21812);
nand U23103 (N_23103,N_19542,N_20574);
nor U23104 (N_23104,N_19176,N_20172);
nor U23105 (N_23105,N_19526,N_20293);
nor U23106 (N_23106,N_20750,N_18931);
nand U23107 (N_23107,N_19064,N_21672);
and U23108 (N_23108,N_21650,N_21240);
nor U23109 (N_23109,N_20785,N_20708);
nand U23110 (N_23110,N_21369,N_20745);
or U23111 (N_23111,N_19534,N_21633);
or U23112 (N_23112,N_19879,N_19055);
nor U23113 (N_23113,N_18974,N_20859);
nand U23114 (N_23114,N_19987,N_18883);
or U23115 (N_23115,N_18896,N_20900);
and U23116 (N_23116,N_21245,N_20551);
nand U23117 (N_23117,N_20254,N_19084);
and U23118 (N_23118,N_21268,N_21434);
or U23119 (N_23119,N_21067,N_21311);
nand U23120 (N_23120,N_19279,N_20477);
and U23121 (N_23121,N_20769,N_21228);
nand U23122 (N_23122,N_19878,N_19928);
xnor U23123 (N_23123,N_20418,N_20359);
nand U23124 (N_23124,N_21309,N_20723);
or U23125 (N_23125,N_18947,N_18853);
nand U23126 (N_23126,N_19026,N_20610);
and U23127 (N_23127,N_20534,N_19035);
or U23128 (N_23128,N_19687,N_21215);
nand U23129 (N_23129,N_20787,N_19867);
nand U23130 (N_23130,N_18909,N_20128);
and U23131 (N_23131,N_18827,N_19795);
and U23132 (N_23132,N_19134,N_20160);
nor U23133 (N_23133,N_19814,N_19065);
nand U23134 (N_23134,N_21850,N_18871);
nor U23135 (N_23135,N_19822,N_19379);
nand U23136 (N_23136,N_19944,N_19636);
xor U23137 (N_23137,N_18757,N_21666);
nand U23138 (N_23138,N_19957,N_20348);
nand U23139 (N_23139,N_21779,N_21630);
or U23140 (N_23140,N_20214,N_21203);
nand U23141 (N_23141,N_18835,N_20119);
nor U23142 (N_23142,N_19590,N_21188);
and U23143 (N_23143,N_21682,N_18868);
and U23144 (N_23144,N_18771,N_20546);
nor U23145 (N_23145,N_21552,N_21791);
or U23146 (N_23146,N_19049,N_20758);
nor U23147 (N_23147,N_19138,N_21846);
nand U23148 (N_23148,N_19126,N_20929);
and U23149 (N_23149,N_21302,N_19329);
or U23150 (N_23150,N_21525,N_21582);
nor U23151 (N_23151,N_21259,N_19874);
or U23152 (N_23152,N_19982,N_20113);
and U23153 (N_23153,N_19102,N_20514);
nor U23154 (N_23154,N_20414,N_19551);
and U23155 (N_23155,N_19661,N_20391);
nand U23156 (N_23156,N_19834,N_19394);
and U23157 (N_23157,N_19664,N_20578);
xnor U23158 (N_23158,N_19637,N_20399);
xnor U23159 (N_23159,N_20475,N_19611);
nor U23160 (N_23160,N_20018,N_21070);
nand U23161 (N_23161,N_20007,N_19974);
nand U23162 (N_23162,N_19237,N_21152);
nand U23163 (N_23163,N_18933,N_20831);
or U23164 (N_23164,N_19748,N_20893);
nand U23165 (N_23165,N_20131,N_20530);
or U23166 (N_23166,N_20588,N_19338);
and U23167 (N_23167,N_21668,N_19744);
nor U23168 (N_23168,N_20432,N_19815);
nor U23169 (N_23169,N_20353,N_18763);
xnor U23170 (N_23170,N_21057,N_21018);
nor U23171 (N_23171,N_19779,N_20605);
nor U23172 (N_23172,N_21874,N_18964);
or U23173 (N_23173,N_20572,N_18929);
nor U23174 (N_23174,N_18976,N_20645);
and U23175 (N_23175,N_19280,N_21327);
nand U23176 (N_23176,N_21623,N_19554);
nand U23177 (N_23177,N_20694,N_18840);
and U23178 (N_23178,N_20449,N_18905);
and U23179 (N_23179,N_21036,N_21282);
nor U23180 (N_23180,N_21450,N_21028);
or U23181 (N_23181,N_19723,N_19603);
xnor U23182 (N_23182,N_19523,N_19393);
nor U23183 (N_23183,N_19203,N_19240);
nand U23184 (N_23184,N_20410,N_19407);
nor U23185 (N_23185,N_21184,N_19085);
nor U23186 (N_23186,N_19086,N_19756);
nand U23187 (N_23187,N_21414,N_19193);
or U23188 (N_23188,N_20747,N_19971);
xnor U23189 (N_23189,N_21613,N_21324);
and U23190 (N_23190,N_21485,N_21106);
nor U23191 (N_23191,N_20693,N_18825);
nor U23192 (N_23192,N_20821,N_21231);
nand U23193 (N_23193,N_19094,N_20288);
or U23194 (N_23194,N_21719,N_20232);
nand U23195 (N_23195,N_19961,N_21402);
nand U23196 (N_23196,N_21570,N_19574);
and U23197 (N_23197,N_20954,N_20066);
and U23198 (N_23198,N_20591,N_19512);
nand U23199 (N_23199,N_19604,N_19412);
xnor U23200 (N_23200,N_21055,N_21782);
nand U23201 (N_23201,N_21724,N_20016);
nand U23202 (N_23202,N_21873,N_20681);
nor U23203 (N_23203,N_20803,N_19330);
or U23204 (N_23204,N_19869,N_19988);
xor U23205 (N_23205,N_21226,N_20845);
or U23206 (N_23206,N_20815,N_20421);
nor U23207 (N_23207,N_20981,N_18930);
nor U23208 (N_23208,N_19807,N_20801);
xnor U23209 (N_23209,N_20962,N_21175);
or U23210 (N_23210,N_21540,N_21531);
nand U23211 (N_23211,N_19278,N_20731);
nand U23212 (N_23212,N_19550,N_19087);
nor U23213 (N_23213,N_20753,N_21467);
nand U23214 (N_23214,N_19643,N_19560);
nand U23215 (N_23215,N_19469,N_18863);
and U23216 (N_23216,N_20505,N_21750);
nor U23217 (N_23217,N_21129,N_19731);
nand U23218 (N_23218,N_21813,N_19626);
nand U23219 (N_23219,N_21759,N_21109);
nor U23220 (N_23220,N_21859,N_18809);
xor U23221 (N_23221,N_20667,N_20607);
or U23222 (N_23222,N_21638,N_18815);
nand U23223 (N_23223,N_20090,N_19376);
and U23224 (N_23224,N_21714,N_21182);
and U23225 (N_23225,N_20791,N_19365);
xor U23226 (N_23226,N_20909,N_19595);
nor U23227 (N_23227,N_21698,N_19296);
xnor U23228 (N_23228,N_20887,N_21649);
or U23229 (N_23229,N_19552,N_18965);
nand U23230 (N_23230,N_20675,N_19344);
or U23231 (N_23231,N_19846,N_20294);
and U23232 (N_23232,N_21249,N_21761);
nand U23233 (N_23233,N_20737,N_19975);
nand U23234 (N_23234,N_19758,N_21136);
nor U23235 (N_23235,N_18774,N_19509);
nand U23236 (N_23236,N_19575,N_20643);
nor U23237 (N_23237,N_19472,N_20109);
and U23238 (N_23238,N_21100,N_19996);
nand U23239 (N_23239,N_20678,N_21520);
xor U23240 (N_23240,N_19711,N_21059);
or U23241 (N_23241,N_18960,N_21234);
or U23242 (N_23242,N_19766,N_21530);
xor U23243 (N_23243,N_21823,N_20999);
nand U23244 (N_23244,N_20051,N_21462);
nor U23245 (N_23245,N_21409,N_21699);
nor U23246 (N_23246,N_20685,N_20464);
and U23247 (N_23247,N_21546,N_19479);
nand U23248 (N_23248,N_21005,N_20249);
nor U23249 (N_23249,N_19513,N_20245);
nor U23250 (N_23250,N_20703,N_19989);
xnor U23251 (N_23251,N_21833,N_21557);
and U23252 (N_23252,N_18973,N_21808);
or U23253 (N_23253,N_21039,N_19819);
and U23254 (N_23254,N_19889,N_21429);
or U23255 (N_23255,N_20759,N_19253);
or U23256 (N_23256,N_18886,N_20290);
and U23257 (N_23257,N_21772,N_19036);
nor U23258 (N_23258,N_18785,N_20088);
nand U23259 (N_23259,N_19853,N_21437);
or U23260 (N_23260,N_21447,N_20177);
nand U23261 (N_23261,N_19732,N_18768);
nor U23262 (N_23262,N_21381,N_20361);
and U23263 (N_23263,N_20029,N_21466);
nand U23264 (N_23264,N_19671,N_20928);
and U23265 (N_23265,N_21726,N_19528);
and U23266 (N_23266,N_21281,N_19327);
nand U23267 (N_23267,N_21728,N_21635);
nand U23268 (N_23268,N_18802,N_19116);
and U23269 (N_23269,N_20222,N_20701);
nor U23270 (N_23270,N_19385,N_21316);
and U23271 (N_23271,N_18997,N_19242);
xnor U23272 (N_23272,N_21158,N_18791);
nor U23273 (N_23273,N_20714,N_19556);
or U23274 (N_23274,N_19835,N_20089);
nand U23275 (N_23275,N_21637,N_19266);
nand U23276 (N_23276,N_21617,N_21473);
or U23277 (N_23277,N_19352,N_21077);
nand U23278 (N_23278,N_20021,N_21686);
and U23279 (N_23279,N_19701,N_19309);
nor U23280 (N_23280,N_20331,N_21769);
nand U23281 (N_23281,N_20491,N_21156);
or U23282 (N_23282,N_20719,N_20544);
and U23283 (N_23283,N_20347,N_19570);
xor U23284 (N_23284,N_19685,N_20059);
nor U23285 (N_23285,N_20735,N_21553);
xnor U23286 (N_23286,N_20381,N_20806);
nand U23287 (N_23287,N_21518,N_21665);
and U23288 (N_23288,N_20350,N_18908);
nor U23289 (N_23289,N_19529,N_18833);
nand U23290 (N_23290,N_21512,N_19058);
xor U23291 (N_23291,N_19345,N_21747);
and U23292 (N_23292,N_19488,N_19583);
nand U23293 (N_23293,N_18766,N_20963);
and U23294 (N_23294,N_21504,N_21443);
nor U23295 (N_23295,N_20557,N_18797);
or U23296 (N_23296,N_18928,N_19158);
nor U23297 (N_23297,N_20512,N_21734);
or U23298 (N_23298,N_19683,N_20498);
or U23299 (N_23299,N_19797,N_21562);
or U23300 (N_23300,N_21334,N_20907);
nor U23301 (N_23301,N_21826,N_19718);
nand U23302 (N_23302,N_20095,N_21353);
or U23303 (N_23303,N_20881,N_19808);
nor U23304 (N_23304,N_19677,N_21139);
or U23305 (N_23305,N_20771,N_19259);
nand U23306 (N_23306,N_20203,N_20121);
or U23307 (N_23307,N_20129,N_20730);
and U23308 (N_23308,N_20447,N_18954);
or U23309 (N_23309,N_19953,N_19508);
or U23310 (N_23310,N_21853,N_20436);
or U23311 (N_23311,N_19599,N_20608);
nand U23312 (N_23312,N_19674,N_19210);
nor U23313 (N_23313,N_20094,N_20263);
or U23314 (N_23314,N_20465,N_19348);
and U23315 (N_23315,N_20468,N_20313);
nand U23316 (N_23316,N_20760,N_21855);
and U23317 (N_23317,N_18860,N_21041);
and U23318 (N_23318,N_20861,N_19698);
and U23319 (N_23319,N_20912,N_20314);
and U23320 (N_23320,N_21702,N_20836);
or U23321 (N_23321,N_20207,N_21814);
nor U23322 (N_23322,N_21284,N_20429);
nand U23323 (N_23323,N_20948,N_21337);
nor U23324 (N_23324,N_21751,N_19478);
nand U23325 (N_23325,N_21053,N_19804);
or U23326 (N_23326,N_19743,N_19201);
nor U23327 (N_23327,N_20506,N_19272);
and U23328 (N_23328,N_20989,N_20554);
nand U23329 (N_23329,N_20653,N_20716);
or U23330 (N_23330,N_19475,N_19032);
nor U23331 (N_23331,N_20698,N_19074);
nor U23332 (N_23332,N_19761,N_19584);
xnor U23333 (N_23333,N_20417,N_21162);
nand U23334 (N_23334,N_21523,N_21481);
or U23335 (N_23335,N_21071,N_20987);
nor U23336 (N_23336,N_20015,N_21296);
and U23337 (N_23337,N_19648,N_21322);
xnor U23338 (N_23338,N_19098,N_21144);
nand U23339 (N_23339,N_18781,N_19959);
nand U23340 (N_23340,N_21799,N_21478);
or U23341 (N_23341,N_19789,N_21718);
and U23342 (N_23342,N_20043,N_19140);
xnor U23343 (N_23343,N_19157,N_20915);
nor U23344 (N_23344,N_18764,N_21102);
or U23345 (N_23345,N_18925,N_19411);
nand U23346 (N_23346,N_20085,N_19429);
and U23347 (N_23347,N_21566,N_19241);
and U23348 (N_23348,N_20155,N_19159);
nand U23349 (N_23349,N_18919,N_19265);
xnor U23350 (N_23350,N_19318,N_19230);
nand U23351 (N_23351,N_20767,N_19511);
xor U23352 (N_23352,N_20527,N_19828);
or U23353 (N_23353,N_21390,N_19631);
or U23354 (N_23354,N_19968,N_20299);
xor U23355 (N_23355,N_19422,N_19495);
and U23356 (N_23356,N_19380,N_19548);
nor U23357 (N_23357,N_21610,N_20580);
nand U23358 (N_23358,N_19443,N_21154);
nor U23359 (N_23359,N_20628,N_19447);
and U23360 (N_23360,N_21076,N_20490);
nand U23361 (N_23361,N_19651,N_20199);
nand U23362 (N_23362,N_21127,N_19195);
nand U23363 (N_23363,N_20460,N_21313);
and U23364 (N_23364,N_21789,N_18872);
or U23365 (N_23365,N_19340,N_19008);
or U23366 (N_23366,N_21535,N_21560);
or U23367 (N_23367,N_20351,N_19503);
xor U23368 (N_23368,N_20167,N_19213);
nand U23369 (N_23369,N_20690,N_19426);
nor U23370 (N_23370,N_19947,N_21527);
or U23371 (N_23371,N_20375,N_20957);
or U23372 (N_23372,N_18884,N_20923);
nor U23373 (N_23373,N_21006,N_21660);
nor U23374 (N_23374,N_20799,N_19716);
or U23375 (N_23375,N_19202,N_21054);
or U23376 (N_23376,N_19402,N_19579);
nor U23377 (N_23377,N_21667,N_20033);
or U23378 (N_23378,N_19812,N_21681);
nor U23379 (N_23379,N_20582,N_20648);
nand U23380 (N_23380,N_20223,N_19994);
nor U23381 (N_23381,N_19009,N_19919);
nor U23382 (N_23382,N_19665,N_19491);
nor U23383 (N_23383,N_21199,N_19498);
xnor U23384 (N_23384,N_18805,N_21326);
nand U23385 (N_23385,N_20798,N_20697);
nor U23386 (N_23386,N_20216,N_20364);
nand U23387 (N_23387,N_21631,N_18876);
or U23388 (N_23388,N_21746,N_21469);
and U23389 (N_23389,N_21232,N_18816);
nor U23390 (N_23390,N_20713,N_19320);
xor U23391 (N_23391,N_21137,N_19191);
and U23392 (N_23392,N_21171,N_19439);
and U23393 (N_23393,N_20463,N_21647);
and U23394 (N_23394,N_19048,N_21593);
and U23395 (N_23395,N_19589,N_18839);
nand U23396 (N_23396,N_20387,N_19115);
or U23397 (N_23397,N_21439,N_21676);
and U23398 (N_23398,N_19122,N_21765);
or U23399 (N_23399,N_19490,N_21585);
or U23400 (N_23400,N_20536,N_21764);
nand U23401 (N_23401,N_20926,N_19360);
or U23402 (N_23402,N_20198,N_20139);
nor U23403 (N_23403,N_21497,N_20425);
nor U23404 (N_23404,N_21392,N_19639);
nor U23405 (N_23405,N_20332,N_21388);
nor U23406 (N_23406,N_21741,N_20813);
nor U23407 (N_23407,N_18778,N_21066);
nand U23408 (N_23408,N_19796,N_20919);
and U23409 (N_23409,N_20416,N_19995);
or U23410 (N_23410,N_21488,N_21848);
or U23411 (N_23411,N_19434,N_20947);
nand U23412 (N_23412,N_20509,N_20406);
xor U23413 (N_23413,N_20102,N_19962);
nand U23414 (N_23414,N_21017,N_21475);
nor U23415 (N_23415,N_21423,N_19313);
or U23416 (N_23416,N_19871,N_21009);
nand U23417 (N_23417,N_18844,N_20531);
or U23418 (N_23418,N_19792,N_21767);
and U23419 (N_23419,N_20686,N_20371);
or U23420 (N_23420,N_19367,N_20242);
and U23421 (N_23421,N_19372,N_21428);
xor U23422 (N_23422,N_21591,N_20115);
xor U23423 (N_23423,N_20873,N_20975);
nor U23424 (N_23424,N_19613,N_18959);
xnor U23425 (N_23425,N_19941,N_19580);
nor U23426 (N_23426,N_19616,N_21112);
nor U23427 (N_23427,N_19450,N_20122);
or U23428 (N_23428,N_19882,N_20891);
nor U23429 (N_23429,N_21433,N_19854);
and U23430 (N_23430,N_21205,N_20519);
and U23431 (N_23431,N_19310,N_20892);
xnor U23432 (N_23432,N_19150,N_19325);
nor U23433 (N_23433,N_20479,N_20123);
and U23434 (N_23434,N_21247,N_19884);
and U23435 (N_23435,N_19608,N_19003);
or U23436 (N_23436,N_21832,N_21019);
or U23437 (N_23437,N_19659,N_18886);
and U23438 (N_23438,N_19361,N_21285);
or U23439 (N_23439,N_20655,N_19400);
and U23440 (N_23440,N_21293,N_18961);
and U23441 (N_23441,N_19899,N_21570);
nand U23442 (N_23442,N_20171,N_20708);
nor U23443 (N_23443,N_21257,N_20256);
and U23444 (N_23444,N_20121,N_20528);
or U23445 (N_23445,N_19787,N_19903);
nand U23446 (N_23446,N_21744,N_19059);
and U23447 (N_23447,N_21256,N_19108);
and U23448 (N_23448,N_20981,N_21399);
nand U23449 (N_23449,N_21815,N_19090);
nand U23450 (N_23450,N_21652,N_20849);
xor U23451 (N_23451,N_21006,N_20567);
nand U23452 (N_23452,N_20349,N_21051);
nor U23453 (N_23453,N_20092,N_19195);
nor U23454 (N_23454,N_21616,N_20053);
nand U23455 (N_23455,N_19373,N_19031);
or U23456 (N_23456,N_20801,N_19257);
xnor U23457 (N_23457,N_19788,N_21273);
or U23458 (N_23458,N_20430,N_19406);
nor U23459 (N_23459,N_18966,N_20294);
nor U23460 (N_23460,N_20231,N_21825);
nor U23461 (N_23461,N_19938,N_21317);
or U23462 (N_23462,N_18975,N_20284);
nand U23463 (N_23463,N_19167,N_18795);
nand U23464 (N_23464,N_18955,N_20536);
and U23465 (N_23465,N_21322,N_21065);
or U23466 (N_23466,N_20924,N_21426);
or U23467 (N_23467,N_20580,N_19229);
nor U23468 (N_23468,N_19048,N_20119);
nand U23469 (N_23469,N_19591,N_21860);
or U23470 (N_23470,N_19469,N_20996);
nor U23471 (N_23471,N_18899,N_19584);
or U23472 (N_23472,N_20592,N_21761);
nor U23473 (N_23473,N_19960,N_19574);
and U23474 (N_23474,N_21745,N_20551);
and U23475 (N_23475,N_18925,N_21261);
or U23476 (N_23476,N_19333,N_21680);
or U23477 (N_23477,N_18959,N_19687);
or U23478 (N_23478,N_20186,N_19811);
nor U23479 (N_23479,N_18945,N_18992);
nand U23480 (N_23480,N_19340,N_19688);
or U23481 (N_23481,N_21568,N_21523);
and U23482 (N_23482,N_18792,N_20326);
or U23483 (N_23483,N_19968,N_19757);
or U23484 (N_23484,N_20330,N_18926);
and U23485 (N_23485,N_20160,N_20702);
and U23486 (N_23486,N_18814,N_20730);
nand U23487 (N_23487,N_20370,N_19677);
xnor U23488 (N_23488,N_21154,N_20947);
or U23489 (N_23489,N_19987,N_20808);
and U23490 (N_23490,N_21279,N_19580);
or U23491 (N_23491,N_18937,N_19221);
or U23492 (N_23492,N_20983,N_18792);
nor U23493 (N_23493,N_20586,N_21730);
and U23494 (N_23494,N_21874,N_19637);
and U23495 (N_23495,N_21189,N_21199);
nor U23496 (N_23496,N_21290,N_21846);
or U23497 (N_23497,N_18801,N_21717);
and U23498 (N_23498,N_19421,N_20165);
and U23499 (N_23499,N_21017,N_21104);
nand U23500 (N_23500,N_21846,N_21251);
nand U23501 (N_23501,N_19968,N_21003);
and U23502 (N_23502,N_21196,N_21763);
or U23503 (N_23503,N_20997,N_19253);
and U23504 (N_23504,N_21830,N_21320);
xor U23505 (N_23505,N_20709,N_20973);
and U23506 (N_23506,N_20509,N_21634);
nor U23507 (N_23507,N_20503,N_21520);
or U23508 (N_23508,N_19879,N_19937);
nand U23509 (N_23509,N_18928,N_21005);
or U23510 (N_23510,N_19936,N_21747);
xnor U23511 (N_23511,N_18902,N_21172);
nand U23512 (N_23512,N_18847,N_20686);
and U23513 (N_23513,N_19547,N_21666);
and U23514 (N_23514,N_21071,N_19171);
nand U23515 (N_23515,N_19716,N_21022);
nand U23516 (N_23516,N_21093,N_19858);
or U23517 (N_23517,N_19444,N_21618);
nand U23518 (N_23518,N_20552,N_18887);
or U23519 (N_23519,N_20804,N_20520);
and U23520 (N_23520,N_20808,N_21369);
and U23521 (N_23521,N_20414,N_20185);
nand U23522 (N_23522,N_20633,N_20028);
or U23523 (N_23523,N_20973,N_19678);
nand U23524 (N_23524,N_21583,N_19821);
and U23525 (N_23525,N_21375,N_20960);
or U23526 (N_23526,N_20976,N_20977);
and U23527 (N_23527,N_21217,N_20481);
nand U23528 (N_23528,N_19609,N_19006);
or U23529 (N_23529,N_19458,N_20899);
xor U23530 (N_23530,N_20604,N_19460);
or U23531 (N_23531,N_19118,N_21118);
xor U23532 (N_23532,N_19027,N_19700);
or U23533 (N_23533,N_19412,N_20311);
or U23534 (N_23534,N_19857,N_18960);
and U23535 (N_23535,N_21188,N_19365);
nor U23536 (N_23536,N_20052,N_19914);
and U23537 (N_23537,N_21315,N_21731);
nor U23538 (N_23538,N_19037,N_21809);
nand U23539 (N_23539,N_19260,N_19318);
nand U23540 (N_23540,N_19538,N_20870);
and U23541 (N_23541,N_20965,N_20297);
or U23542 (N_23542,N_19247,N_19639);
and U23543 (N_23543,N_20356,N_21485);
nor U23544 (N_23544,N_21632,N_19070);
nand U23545 (N_23545,N_20644,N_19033);
and U23546 (N_23546,N_18845,N_20615);
or U23547 (N_23547,N_21778,N_20622);
or U23548 (N_23548,N_20763,N_20669);
nor U23549 (N_23549,N_18920,N_21697);
or U23550 (N_23550,N_18750,N_20334);
and U23551 (N_23551,N_19227,N_19925);
or U23552 (N_23552,N_19788,N_21228);
nand U23553 (N_23553,N_21774,N_21603);
nor U23554 (N_23554,N_21448,N_20966);
xor U23555 (N_23555,N_19590,N_21042);
or U23556 (N_23556,N_21221,N_21346);
nor U23557 (N_23557,N_19775,N_18768);
and U23558 (N_23558,N_18898,N_21223);
and U23559 (N_23559,N_21188,N_19213);
or U23560 (N_23560,N_20407,N_21372);
nor U23561 (N_23561,N_19686,N_21317);
nor U23562 (N_23562,N_19002,N_20923);
or U23563 (N_23563,N_19738,N_21571);
nor U23564 (N_23564,N_19831,N_21414);
and U23565 (N_23565,N_19162,N_20339);
and U23566 (N_23566,N_20057,N_18883);
and U23567 (N_23567,N_20730,N_21440);
nand U23568 (N_23568,N_20429,N_19923);
or U23569 (N_23569,N_19811,N_20829);
or U23570 (N_23570,N_21451,N_18806);
xnor U23571 (N_23571,N_20610,N_19518);
or U23572 (N_23572,N_21546,N_20224);
or U23573 (N_23573,N_20520,N_19124);
and U23574 (N_23574,N_19688,N_19042);
nor U23575 (N_23575,N_21734,N_21008);
nand U23576 (N_23576,N_19117,N_21786);
xor U23577 (N_23577,N_19348,N_21248);
nor U23578 (N_23578,N_21741,N_20176);
nand U23579 (N_23579,N_19993,N_20662);
nor U23580 (N_23580,N_19230,N_19377);
or U23581 (N_23581,N_20886,N_19988);
nand U23582 (N_23582,N_20430,N_20412);
nor U23583 (N_23583,N_18776,N_21093);
nand U23584 (N_23584,N_21519,N_21012);
or U23585 (N_23585,N_19625,N_19473);
nand U23586 (N_23586,N_20912,N_19771);
nand U23587 (N_23587,N_20701,N_20574);
xnor U23588 (N_23588,N_20970,N_20314);
or U23589 (N_23589,N_18822,N_19610);
nor U23590 (N_23590,N_21412,N_19877);
and U23591 (N_23591,N_21104,N_19676);
and U23592 (N_23592,N_21572,N_19860);
nor U23593 (N_23593,N_20459,N_21872);
nand U23594 (N_23594,N_18767,N_19943);
nand U23595 (N_23595,N_20445,N_19955);
nor U23596 (N_23596,N_19910,N_19803);
nor U23597 (N_23597,N_20179,N_20172);
or U23598 (N_23598,N_19140,N_21849);
and U23599 (N_23599,N_20543,N_21575);
or U23600 (N_23600,N_21792,N_19379);
xor U23601 (N_23601,N_19644,N_21011);
nor U23602 (N_23602,N_20553,N_21795);
or U23603 (N_23603,N_18837,N_20888);
nand U23604 (N_23604,N_19502,N_20757);
nor U23605 (N_23605,N_19281,N_19136);
nor U23606 (N_23606,N_18891,N_19151);
and U23607 (N_23607,N_19529,N_19427);
nor U23608 (N_23608,N_21268,N_21720);
nor U23609 (N_23609,N_19273,N_21120);
nand U23610 (N_23610,N_21660,N_19048);
and U23611 (N_23611,N_19627,N_19422);
nor U23612 (N_23612,N_18942,N_20141);
nor U23613 (N_23613,N_21271,N_18816);
nor U23614 (N_23614,N_20025,N_19589);
nand U23615 (N_23615,N_19919,N_21594);
or U23616 (N_23616,N_21353,N_21296);
and U23617 (N_23617,N_20489,N_20685);
nor U23618 (N_23618,N_21786,N_19227);
or U23619 (N_23619,N_21225,N_19377);
nor U23620 (N_23620,N_21127,N_20802);
nor U23621 (N_23621,N_21546,N_19088);
and U23622 (N_23622,N_21692,N_20887);
nor U23623 (N_23623,N_19112,N_20665);
and U23624 (N_23624,N_21574,N_20473);
nand U23625 (N_23625,N_21445,N_21280);
nor U23626 (N_23626,N_21193,N_20064);
or U23627 (N_23627,N_21620,N_18958);
and U23628 (N_23628,N_20700,N_21520);
nand U23629 (N_23629,N_19112,N_20245);
nor U23630 (N_23630,N_19605,N_19479);
nor U23631 (N_23631,N_21228,N_20381);
nand U23632 (N_23632,N_20092,N_21157);
and U23633 (N_23633,N_20080,N_21546);
xnor U23634 (N_23634,N_19033,N_19109);
or U23635 (N_23635,N_20313,N_18839);
or U23636 (N_23636,N_19058,N_20683);
xor U23637 (N_23637,N_20703,N_21260);
nor U23638 (N_23638,N_21312,N_19718);
nor U23639 (N_23639,N_19402,N_19158);
nor U23640 (N_23640,N_18853,N_20822);
and U23641 (N_23641,N_20424,N_19663);
xor U23642 (N_23642,N_21363,N_21326);
or U23643 (N_23643,N_21625,N_18754);
xor U23644 (N_23644,N_21855,N_21354);
nor U23645 (N_23645,N_19002,N_21371);
or U23646 (N_23646,N_19742,N_21740);
nand U23647 (N_23647,N_21177,N_21240);
and U23648 (N_23648,N_20081,N_21031);
nor U23649 (N_23649,N_20284,N_20574);
nor U23650 (N_23650,N_18851,N_20395);
or U23651 (N_23651,N_21860,N_20285);
xor U23652 (N_23652,N_21582,N_21766);
nand U23653 (N_23653,N_19312,N_18833);
or U23654 (N_23654,N_21169,N_21349);
nor U23655 (N_23655,N_19493,N_18776);
and U23656 (N_23656,N_19304,N_19779);
nor U23657 (N_23657,N_21255,N_21124);
xor U23658 (N_23658,N_20929,N_21550);
nand U23659 (N_23659,N_21169,N_20365);
or U23660 (N_23660,N_20928,N_20669);
and U23661 (N_23661,N_19352,N_21112);
nand U23662 (N_23662,N_20285,N_19855);
nand U23663 (N_23663,N_20319,N_20370);
or U23664 (N_23664,N_19558,N_20428);
nand U23665 (N_23665,N_19633,N_20436);
nand U23666 (N_23666,N_21457,N_20182);
nand U23667 (N_23667,N_18928,N_19530);
nand U23668 (N_23668,N_21330,N_20928);
or U23669 (N_23669,N_18962,N_19828);
nor U23670 (N_23670,N_19977,N_19676);
nand U23671 (N_23671,N_19046,N_21629);
nor U23672 (N_23672,N_19816,N_20072);
nor U23673 (N_23673,N_19975,N_18802);
nor U23674 (N_23674,N_19513,N_19452);
nor U23675 (N_23675,N_19899,N_19329);
nand U23676 (N_23676,N_20251,N_18915);
or U23677 (N_23677,N_21787,N_19890);
xnor U23678 (N_23678,N_19395,N_21593);
nor U23679 (N_23679,N_21772,N_20124);
and U23680 (N_23680,N_20165,N_20894);
xnor U23681 (N_23681,N_21287,N_18756);
or U23682 (N_23682,N_21656,N_21822);
and U23683 (N_23683,N_19246,N_19853);
nand U23684 (N_23684,N_20841,N_20008);
xnor U23685 (N_23685,N_19610,N_21423);
xor U23686 (N_23686,N_19621,N_21107);
or U23687 (N_23687,N_19798,N_20251);
or U23688 (N_23688,N_20631,N_20574);
or U23689 (N_23689,N_20542,N_18795);
or U23690 (N_23690,N_19568,N_21181);
and U23691 (N_23691,N_20039,N_20852);
xor U23692 (N_23692,N_21619,N_20430);
nand U23693 (N_23693,N_20790,N_21038);
nor U23694 (N_23694,N_20720,N_21740);
nand U23695 (N_23695,N_19620,N_20553);
xor U23696 (N_23696,N_18963,N_20378);
nand U23697 (N_23697,N_20557,N_18921);
xnor U23698 (N_23698,N_19065,N_20724);
or U23699 (N_23699,N_20446,N_19403);
or U23700 (N_23700,N_18984,N_21488);
or U23701 (N_23701,N_18812,N_20233);
and U23702 (N_23702,N_20847,N_19718);
nor U23703 (N_23703,N_21693,N_21665);
or U23704 (N_23704,N_21482,N_21579);
nor U23705 (N_23705,N_21130,N_20025);
and U23706 (N_23706,N_19542,N_20689);
and U23707 (N_23707,N_21442,N_19685);
nor U23708 (N_23708,N_19004,N_20491);
and U23709 (N_23709,N_18813,N_20048);
nor U23710 (N_23710,N_21655,N_20865);
and U23711 (N_23711,N_19706,N_21783);
or U23712 (N_23712,N_20797,N_20218);
and U23713 (N_23713,N_18785,N_20007);
nor U23714 (N_23714,N_20896,N_18982);
nor U23715 (N_23715,N_19693,N_19332);
nor U23716 (N_23716,N_19291,N_20000);
nand U23717 (N_23717,N_19698,N_20179);
or U23718 (N_23718,N_19955,N_21137);
and U23719 (N_23719,N_19304,N_20336);
nand U23720 (N_23720,N_21146,N_19245);
nand U23721 (N_23721,N_19305,N_21612);
nor U23722 (N_23722,N_19323,N_19008);
or U23723 (N_23723,N_21616,N_19802);
nand U23724 (N_23724,N_20503,N_20803);
or U23725 (N_23725,N_20009,N_20917);
nor U23726 (N_23726,N_18806,N_21236);
and U23727 (N_23727,N_20539,N_20607);
nand U23728 (N_23728,N_20085,N_18823);
nor U23729 (N_23729,N_20206,N_18814);
and U23730 (N_23730,N_20085,N_21605);
and U23731 (N_23731,N_19599,N_19762);
nor U23732 (N_23732,N_20559,N_20961);
and U23733 (N_23733,N_19825,N_19385);
or U23734 (N_23734,N_20801,N_19791);
or U23735 (N_23735,N_19337,N_20873);
nor U23736 (N_23736,N_20214,N_20506);
or U23737 (N_23737,N_21595,N_21168);
nor U23738 (N_23738,N_20798,N_21568);
nor U23739 (N_23739,N_20260,N_20692);
xnor U23740 (N_23740,N_19873,N_20075);
nand U23741 (N_23741,N_21572,N_19521);
nand U23742 (N_23742,N_19452,N_20816);
and U23743 (N_23743,N_21195,N_21762);
xnor U23744 (N_23744,N_20047,N_19766);
or U23745 (N_23745,N_20262,N_18865);
or U23746 (N_23746,N_19646,N_20486);
and U23747 (N_23747,N_18794,N_19746);
and U23748 (N_23748,N_20107,N_19086);
and U23749 (N_23749,N_19820,N_21514);
or U23750 (N_23750,N_20783,N_21162);
and U23751 (N_23751,N_19876,N_21593);
xnor U23752 (N_23752,N_20481,N_21456);
or U23753 (N_23753,N_19861,N_21069);
nand U23754 (N_23754,N_18840,N_18975);
and U23755 (N_23755,N_20246,N_19317);
nor U23756 (N_23756,N_20098,N_20813);
and U23757 (N_23757,N_19116,N_21676);
nand U23758 (N_23758,N_19294,N_19329);
xor U23759 (N_23759,N_19442,N_18954);
xor U23760 (N_23760,N_19347,N_20748);
or U23761 (N_23761,N_20718,N_21089);
xor U23762 (N_23762,N_19092,N_21328);
nand U23763 (N_23763,N_20019,N_18887);
and U23764 (N_23764,N_21322,N_18890);
or U23765 (N_23765,N_21600,N_21144);
nand U23766 (N_23766,N_21049,N_20729);
nor U23767 (N_23767,N_20044,N_20640);
xor U23768 (N_23768,N_21472,N_21527);
or U23769 (N_23769,N_20604,N_20069);
nand U23770 (N_23770,N_19457,N_20416);
or U23771 (N_23771,N_19162,N_20684);
and U23772 (N_23772,N_20886,N_20241);
and U23773 (N_23773,N_20885,N_20957);
nand U23774 (N_23774,N_19699,N_21706);
and U23775 (N_23775,N_19326,N_19110);
or U23776 (N_23776,N_21020,N_19723);
xnor U23777 (N_23777,N_20529,N_19074);
or U23778 (N_23778,N_20468,N_18796);
or U23779 (N_23779,N_21087,N_21573);
and U23780 (N_23780,N_20719,N_20818);
nand U23781 (N_23781,N_20091,N_20618);
and U23782 (N_23782,N_19707,N_19010);
nor U23783 (N_23783,N_19976,N_20748);
or U23784 (N_23784,N_20105,N_19347);
or U23785 (N_23785,N_21755,N_18806);
and U23786 (N_23786,N_19165,N_18964);
and U23787 (N_23787,N_21518,N_19542);
nor U23788 (N_23788,N_19648,N_18818);
or U23789 (N_23789,N_19746,N_21012);
nand U23790 (N_23790,N_21637,N_19451);
and U23791 (N_23791,N_20557,N_20949);
and U23792 (N_23792,N_21550,N_20373);
xnor U23793 (N_23793,N_21718,N_20433);
nor U23794 (N_23794,N_20999,N_21090);
and U23795 (N_23795,N_19272,N_21822);
and U23796 (N_23796,N_19624,N_20956);
nand U23797 (N_23797,N_19041,N_21388);
nand U23798 (N_23798,N_20973,N_21349);
nand U23799 (N_23799,N_21394,N_19871);
and U23800 (N_23800,N_21706,N_21125);
or U23801 (N_23801,N_19298,N_21811);
nand U23802 (N_23802,N_21675,N_18933);
and U23803 (N_23803,N_20204,N_20774);
xnor U23804 (N_23804,N_18750,N_19268);
and U23805 (N_23805,N_18937,N_20321);
or U23806 (N_23806,N_19698,N_19056);
nand U23807 (N_23807,N_19751,N_21810);
and U23808 (N_23808,N_18985,N_21707);
and U23809 (N_23809,N_21077,N_20635);
nor U23810 (N_23810,N_19597,N_19127);
nand U23811 (N_23811,N_20698,N_19541);
or U23812 (N_23812,N_20146,N_20298);
nand U23813 (N_23813,N_19130,N_20258);
and U23814 (N_23814,N_21354,N_21674);
nor U23815 (N_23815,N_19172,N_21007);
nand U23816 (N_23816,N_21151,N_21319);
nor U23817 (N_23817,N_21334,N_19825);
xor U23818 (N_23818,N_19935,N_19823);
or U23819 (N_23819,N_18757,N_18814);
or U23820 (N_23820,N_19812,N_21873);
or U23821 (N_23821,N_20491,N_19335);
or U23822 (N_23822,N_19547,N_18927);
nor U23823 (N_23823,N_20135,N_19656);
nand U23824 (N_23824,N_21510,N_21689);
xor U23825 (N_23825,N_19720,N_19197);
and U23826 (N_23826,N_19402,N_20732);
and U23827 (N_23827,N_19849,N_20861);
or U23828 (N_23828,N_19584,N_21639);
nor U23829 (N_23829,N_21504,N_19528);
nor U23830 (N_23830,N_21047,N_19779);
xor U23831 (N_23831,N_18775,N_20646);
or U23832 (N_23832,N_21166,N_19727);
and U23833 (N_23833,N_21423,N_20360);
xor U23834 (N_23834,N_21509,N_19637);
xnor U23835 (N_23835,N_20182,N_20816);
and U23836 (N_23836,N_20073,N_21599);
or U23837 (N_23837,N_20343,N_21599);
and U23838 (N_23838,N_19126,N_19854);
nor U23839 (N_23839,N_20904,N_19744);
or U23840 (N_23840,N_21070,N_21159);
or U23841 (N_23841,N_21247,N_19052);
and U23842 (N_23842,N_21007,N_20905);
nand U23843 (N_23843,N_21409,N_21092);
and U23844 (N_23844,N_19654,N_21837);
xnor U23845 (N_23845,N_21226,N_20495);
and U23846 (N_23846,N_18961,N_21733);
nor U23847 (N_23847,N_19140,N_21794);
nor U23848 (N_23848,N_18945,N_20984);
xor U23849 (N_23849,N_21256,N_20924);
and U23850 (N_23850,N_20991,N_19597);
nand U23851 (N_23851,N_21621,N_21414);
and U23852 (N_23852,N_19083,N_20525);
nand U23853 (N_23853,N_21679,N_18761);
and U23854 (N_23854,N_18906,N_19201);
or U23855 (N_23855,N_21787,N_19701);
or U23856 (N_23856,N_20141,N_19109);
and U23857 (N_23857,N_19096,N_21849);
nor U23858 (N_23858,N_18919,N_19647);
or U23859 (N_23859,N_19217,N_21395);
and U23860 (N_23860,N_20173,N_20218);
nor U23861 (N_23861,N_19271,N_20069);
nand U23862 (N_23862,N_21647,N_18945);
and U23863 (N_23863,N_21079,N_20459);
nand U23864 (N_23864,N_20386,N_19215);
or U23865 (N_23865,N_20043,N_20315);
nand U23866 (N_23866,N_21659,N_18873);
and U23867 (N_23867,N_19943,N_20539);
nand U23868 (N_23868,N_21740,N_19527);
xor U23869 (N_23869,N_20084,N_19698);
or U23870 (N_23870,N_20137,N_19808);
nor U23871 (N_23871,N_20645,N_20238);
nand U23872 (N_23872,N_20513,N_20981);
nor U23873 (N_23873,N_20625,N_19348);
nor U23874 (N_23874,N_18763,N_19187);
nor U23875 (N_23875,N_19074,N_20188);
nor U23876 (N_23876,N_21567,N_20465);
or U23877 (N_23877,N_18994,N_18772);
nor U23878 (N_23878,N_20947,N_19822);
nand U23879 (N_23879,N_21610,N_19595);
xnor U23880 (N_23880,N_19318,N_19793);
or U23881 (N_23881,N_18785,N_21592);
nor U23882 (N_23882,N_19297,N_19562);
nor U23883 (N_23883,N_20123,N_19039);
xor U23884 (N_23884,N_19357,N_19761);
and U23885 (N_23885,N_20794,N_19235);
nand U23886 (N_23886,N_21821,N_20681);
or U23887 (N_23887,N_21644,N_21735);
or U23888 (N_23888,N_20057,N_19679);
nor U23889 (N_23889,N_19400,N_21696);
and U23890 (N_23890,N_21139,N_20887);
nand U23891 (N_23891,N_20094,N_18844);
or U23892 (N_23892,N_21758,N_21781);
nor U23893 (N_23893,N_20799,N_21528);
nand U23894 (N_23894,N_20348,N_20249);
nand U23895 (N_23895,N_19628,N_21368);
and U23896 (N_23896,N_19372,N_19200);
nand U23897 (N_23897,N_21224,N_20522);
or U23898 (N_23898,N_21223,N_19618);
nand U23899 (N_23899,N_20787,N_20100);
nor U23900 (N_23900,N_18911,N_21001);
nand U23901 (N_23901,N_19082,N_21204);
xnor U23902 (N_23902,N_19419,N_18767);
or U23903 (N_23903,N_20429,N_19531);
nor U23904 (N_23904,N_20298,N_19464);
or U23905 (N_23905,N_20288,N_19439);
or U23906 (N_23906,N_21583,N_19237);
nor U23907 (N_23907,N_20265,N_20857);
or U23908 (N_23908,N_20284,N_19196);
nand U23909 (N_23909,N_19073,N_18989);
nor U23910 (N_23910,N_18932,N_19145);
or U23911 (N_23911,N_21788,N_19019);
nor U23912 (N_23912,N_20735,N_19200);
and U23913 (N_23913,N_19458,N_20570);
nand U23914 (N_23914,N_19517,N_21129);
nor U23915 (N_23915,N_18846,N_19969);
or U23916 (N_23916,N_20940,N_19673);
nor U23917 (N_23917,N_21663,N_21856);
or U23918 (N_23918,N_20536,N_20535);
or U23919 (N_23919,N_21809,N_20438);
or U23920 (N_23920,N_19558,N_19687);
or U23921 (N_23921,N_18879,N_21253);
nor U23922 (N_23922,N_20079,N_19570);
or U23923 (N_23923,N_21522,N_20574);
xor U23924 (N_23924,N_21716,N_18931);
or U23925 (N_23925,N_20935,N_18971);
or U23926 (N_23926,N_19061,N_19341);
nand U23927 (N_23927,N_19536,N_21300);
nand U23928 (N_23928,N_21104,N_19622);
or U23929 (N_23929,N_20861,N_21261);
nand U23930 (N_23930,N_21647,N_19461);
and U23931 (N_23931,N_19206,N_18962);
nand U23932 (N_23932,N_20538,N_19079);
nand U23933 (N_23933,N_19076,N_19470);
xor U23934 (N_23934,N_19001,N_21851);
nor U23935 (N_23935,N_19367,N_21659);
and U23936 (N_23936,N_21553,N_20170);
and U23937 (N_23937,N_21248,N_21398);
nand U23938 (N_23938,N_20412,N_20781);
nand U23939 (N_23939,N_20172,N_20041);
nor U23940 (N_23940,N_19711,N_18959);
xor U23941 (N_23941,N_21448,N_21287);
nor U23942 (N_23942,N_20865,N_21293);
and U23943 (N_23943,N_21216,N_20181);
nand U23944 (N_23944,N_21773,N_21799);
nand U23945 (N_23945,N_19548,N_20151);
and U23946 (N_23946,N_18849,N_20722);
nand U23947 (N_23947,N_21700,N_21388);
nand U23948 (N_23948,N_20390,N_21450);
or U23949 (N_23949,N_21734,N_20637);
and U23950 (N_23950,N_20841,N_20239);
and U23951 (N_23951,N_18889,N_19229);
or U23952 (N_23952,N_21450,N_21810);
or U23953 (N_23953,N_21683,N_21722);
nor U23954 (N_23954,N_19445,N_19382);
nor U23955 (N_23955,N_20922,N_20988);
or U23956 (N_23956,N_20828,N_18967);
nand U23957 (N_23957,N_19930,N_21334);
and U23958 (N_23958,N_21155,N_20959);
or U23959 (N_23959,N_20203,N_19705);
nor U23960 (N_23960,N_20350,N_20708);
nand U23961 (N_23961,N_20946,N_20972);
xor U23962 (N_23962,N_19031,N_20302);
nand U23963 (N_23963,N_20505,N_21600);
and U23964 (N_23964,N_20996,N_20983);
nor U23965 (N_23965,N_21461,N_19621);
nand U23966 (N_23966,N_20578,N_21585);
and U23967 (N_23967,N_19172,N_19544);
nor U23968 (N_23968,N_21513,N_20206);
nor U23969 (N_23969,N_19547,N_19234);
nand U23970 (N_23970,N_21849,N_19565);
nand U23971 (N_23971,N_21177,N_21576);
or U23972 (N_23972,N_18934,N_21803);
xor U23973 (N_23973,N_21229,N_21449);
nor U23974 (N_23974,N_19865,N_21176);
and U23975 (N_23975,N_19154,N_21312);
nand U23976 (N_23976,N_19585,N_21332);
nand U23977 (N_23977,N_19259,N_20895);
or U23978 (N_23978,N_21158,N_19725);
and U23979 (N_23979,N_21761,N_20469);
and U23980 (N_23980,N_19341,N_18920);
or U23981 (N_23981,N_20272,N_21470);
xnor U23982 (N_23982,N_21872,N_20274);
nor U23983 (N_23983,N_19078,N_19575);
nand U23984 (N_23984,N_19103,N_21671);
nand U23985 (N_23985,N_20847,N_19214);
xnor U23986 (N_23986,N_19878,N_20188);
or U23987 (N_23987,N_21673,N_21172);
nand U23988 (N_23988,N_20675,N_21465);
nor U23989 (N_23989,N_21044,N_18841);
and U23990 (N_23990,N_19376,N_18942);
and U23991 (N_23991,N_20064,N_19128);
or U23992 (N_23992,N_21507,N_20943);
nand U23993 (N_23993,N_21603,N_20452);
nand U23994 (N_23994,N_20243,N_19366);
or U23995 (N_23995,N_20427,N_21321);
nand U23996 (N_23996,N_21858,N_18841);
nor U23997 (N_23997,N_21584,N_21847);
nor U23998 (N_23998,N_21491,N_20366);
and U23999 (N_23999,N_21372,N_19262);
nand U24000 (N_24000,N_20124,N_19004);
nand U24001 (N_24001,N_20313,N_21371);
or U24002 (N_24002,N_19360,N_21182);
nand U24003 (N_24003,N_21596,N_20710);
or U24004 (N_24004,N_19278,N_20537);
nor U24005 (N_24005,N_18969,N_19376);
nor U24006 (N_24006,N_21821,N_20157);
nor U24007 (N_24007,N_19628,N_21836);
nor U24008 (N_24008,N_20890,N_19592);
and U24009 (N_24009,N_19924,N_20466);
nand U24010 (N_24010,N_20467,N_21709);
or U24011 (N_24011,N_21438,N_21622);
and U24012 (N_24012,N_19813,N_19773);
or U24013 (N_24013,N_18902,N_19864);
or U24014 (N_24014,N_19258,N_18849);
and U24015 (N_24015,N_21855,N_19267);
nor U24016 (N_24016,N_19422,N_21679);
or U24017 (N_24017,N_21226,N_20698);
and U24018 (N_24018,N_21019,N_19201);
nor U24019 (N_24019,N_20381,N_20436);
xor U24020 (N_24020,N_19529,N_19343);
or U24021 (N_24021,N_19247,N_21254);
or U24022 (N_24022,N_21487,N_21204);
nor U24023 (N_24023,N_20956,N_21774);
or U24024 (N_24024,N_20880,N_19958);
or U24025 (N_24025,N_19618,N_21669);
nand U24026 (N_24026,N_19928,N_19605);
xnor U24027 (N_24027,N_21685,N_19699);
xor U24028 (N_24028,N_19372,N_19835);
nor U24029 (N_24029,N_21726,N_18845);
xor U24030 (N_24030,N_19697,N_21668);
xnor U24031 (N_24031,N_20034,N_21536);
nor U24032 (N_24032,N_20890,N_20836);
or U24033 (N_24033,N_20472,N_20128);
or U24034 (N_24034,N_21731,N_20020);
and U24035 (N_24035,N_19095,N_21402);
nand U24036 (N_24036,N_19649,N_19300);
and U24037 (N_24037,N_19178,N_20238);
or U24038 (N_24038,N_20687,N_20827);
nand U24039 (N_24039,N_20879,N_21849);
and U24040 (N_24040,N_21439,N_19620);
nand U24041 (N_24041,N_18859,N_20327);
or U24042 (N_24042,N_19604,N_21830);
and U24043 (N_24043,N_19944,N_19982);
xor U24044 (N_24044,N_21868,N_21002);
nor U24045 (N_24045,N_19281,N_21077);
nor U24046 (N_24046,N_21226,N_20230);
nand U24047 (N_24047,N_21621,N_20844);
nand U24048 (N_24048,N_21046,N_20459);
nand U24049 (N_24049,N_18971,N_20759);
xnor U24050 (N_24050,N_20106,N_20640);
nor U24051 (N_24051,N_20862,N_21691);
and U24052 (N_24052,N_20706,N_21660);
and U24053 (N_24053,N_19241,N_21806);
and U24054 (N_24054,N_21478,N_21275);
and U24055 (N_24055,N_21290,N_20398);
nor U24056 (N_24056,N_21594,N_21335);
or U24057 (N_24057,N_19982,N_19380);
and U24058 (N_24058,N_20941,N_18816);
xor U24059 (N_24059,N_19538,N_21516);
nor U24060 (N_24060,N_20155,N_20862);
nand U24061 (N_24061,N_20559,N_20713);
xor U24062 (N_24062,N_21778,N_21134);
and U24063 (N_24063,N_19257,N_19454);
and U24064 (N_24064,N_20391,N_20846);
or U24065 (N_24065,N_19203,N_20273);
nand U24066 (N_24066,N_20385,N_19562);
nand U24067 (N_24067,N_20156,N_21040);
nand U24068 (N_24068,N_19745,N_20339);
nand U24069 (N_24069,N_20948,N_20259);
and U24070 (N_24070,N_18904,N_20749);
or U24071 (N_24071,N_19850,N_20916);
nand U24072 (N_24072,N_19645,N_18851);
nand U24073 (N_24073,N_20857,N_21726);
or U24074 (N_24074,N_19791,N_20579);
or U24075 (N_24075,N_20853,N_18858);
and U24076 (N_24076,N_20115,N_20114);
or U24077 (N_24077,N_19179,N_19355);
or U24078 (N_24078,N_20018,N_20824);
xnor U24079 (N_24079,N_19857,N_19220);
or U24080 (N_24080,N_21553,N_21736);
nor U24081 (N_24081,N_20923,N_18820);
nor U24082 (N_24082,N_19442,N_20489);
and U24083 (N_24083,N_20451,N_18756);
nor U24084 (N_24084,N_19401,N_21853);
and U24085 (N_24085,N_19593,N_21043);
nand U24086 (N_24086,N_19171,N_18950);
and U24087 (N_24087,N_18846,N_20566);
nor U24088 (N_24088,N_21055,N_18886);
nor U24089 (N_24089,N_21035,N_19396);
and U24090 (N_24090,N_21691,N_19576);
nand U24091 (N_24091,N_21814,N_21725);
and U24092 (N_24092,N_20012,N_19565);
nand U24093 (N_24093,N_19848,N_21732);
or U24094 (N_24094,N_20100,N_18831);
or U24095 (N_24095,N_20808,N_21329);
and U24096 (N_24096,N_20056,N_20142);
nor U24097 (N_24097,N_20198,N_20463);
nand U24098 (N_24098,N_21144,N_18823);
nor U24099 (N_24099,N_19566,N_21743);
and U24100 (N_24100,N_19755,N_21259);
xor U24101 (N_24101,N_21549,N_21402);
nor U24102 (N_24102,N_19651,N_20526);
and U24103 (N_24103,N_21369,N_19326);
nand U24104 (N_24104,N_21783,N_20752);
nor U24105 (N_24105,N_20819,N_21789);
or U24106 (N_24106,N_19868,N_20422);
or U24107 (N_24107,N_20765,N_20460);
xnor U24108 (N_24108,N_18948,N_19678);
nor U24109 (N_24109,N_19637,N_19942);
and U24110 (N_24110,N_21094,N_21862);
nand U24111 (N_24111,N_21229,N_21854);
and U24112 (N_24112,N_19336,N_19657);
nand U24113 (N_24113,N_19419,N_19205);
nand U24114 (N_24114,N_21817,N_19873);
xor U24115 (N_24115,N_19649,N_20067);
nand U24116 (N_24116,N_19273,N_19344);
and U24117 (N_24117,N_21017,N_20620);
and U24118 (N_24118,N_19603,N_20942);
nand U24119 (N_24119,N_18871,N_20731);
and U24120 (N_24120,N_19612,N_20269);
or U24121 (N_24121,N_20907,N_21731);
and U24122 (N_24122,N_21394,N_19819);
nor U24123 (N_24123,N_20756,N_18940);
or U24124 (N_24124,N_21340,N_19498);
xor U24125 (N_24125,N_21342,N_21065);
or U24126 (N_24126,N_20624,N_20605);
xnor U24127 (N_24127,N_19122,N_19258);
xnor U24128 (N_24128,N_21108,N_20230);
nand U24129 (N_24129,N_20810,N_20307);
xor U24130 (N_24130,N_19612,N_20693);
nand U24131 (N_24131,N_21482,N_21384);
nor U24132 (N_24132,N_21727,N_21832);
xor U24133 (N_24133,N_18940,N_19737);
and U24134 (N_24134,N_19850,N_19253);
and U24135 (N_24135,N_20321,N_20536);
or U24136 (N_24136,N_19969,N_20984);
xor U24137 (N_24137,N_19794,N_20781);
nand U24138 (N_24138,N_19236,N_21436);
or U24139 (N_24139,N_21242,N_19380);
and U24140 (N_24140,N_18803,N_20039);
nand U24141 (N_24141,N_18998,N_19006);
nor U24142 (N_24142,N_19230,N_21602);
or U24143 (N_24143,N_18828,N_21651);
nand U24144 (N_24144,N_20877,N_21819);
nor U24145 (N_24145,N_19731,N_19781);
nor U24146 (N_24146,N_18989,N_21592);
or U24147 (N_24147,N_18833,N_21300);
and U24148 (N_24148,N_19266,N_21084);
or U24149 (N_24149,N_20169,N_18817);
nand U24150 (N_24150,N_20638,N_19808);
nand U24151 (N_24151,N_19140,N_20130);
and U24152 (N_24152,N_20176,N_20369);
or U24153 (N_24153,N_18817,N_20722);
or U24154 (N_24154,N_20196,N_21462);
nand U24155 (N_24155,N_20690,N_19808);
xor U24156 (N_24156,N_21163,N_21066);
and U24157 (N_24157,N_19714,N_19156);
nor U24158 (N_24158,N_20709,N_21579);
xor U24159 (N_24159,N_21364,N_21521);
and U24160 (N_24160,N_20044,N_18860);
nor U24161 (N_24161,N_21729,N_19339);
nand U24162 (N_24162,N_21065,N_18934);
nor U24163 (N_24163,N_19174,N_20579);
xnor U24164 (N_24164,N_21591,N_20183);
nor U24165 (N_24165,N_19213,N_20379);
and U24166 (N_24166,N_19244,N_21231);
and U24167 (N_24167,N_20786,N_21646);
and U24168 (N_24168,N_19707,N_20283);
xnor U24169 (N_24169,N_21209,N_19778);
or U24170 (N_24170,N_19793,N_19427);
and U24171 (N_24171,N_21213,N_19988);
xor U24172 (N_24172,N_20573,N_20234);
or U24173 (N_24173,N_20231,N_18967);
nor U24174 (N_24174,N_20133,N_19882);
or U24175 (N_24175,N_19230,N_20180);
or U24176 (N_24176,N_21351,N_20218);
and U24177 (N_24177,N_21002,N_19026);
and U24178 (N_24178,N_18784,N_20288);
or U24179 (N_24179,N_21093,N_19353);
nor U24180 (N_24180,N_21787,N_19272);
nor U24181 (N_24181,N_20330,N_19907);
nor U24182 (N_24182,N_20308,N_19759);
and U24183 (N_24183,N_19338,N_19985);
and U24184 (N_24184,N_18938,N_20621);
nand U24185 (N_24185,N_19270,N_21312);
nand U24186 (N_24186,N_21114,N_19383);
and U24187 (N_24187,N_20532,N_20026);
nor U24188 (N_24188,N_20873,N_19692);
nand U24189 (N_24189,N_19251,N_20477);
or U24190 (N_24190,N_20654,N_19745);
xor U24191 (N_24191,N_19503,N_20038);
or U24192 (N_24192,N_21642,N_21368);
and U24193 (N_24193,N_21500,N_21682);
or U24194 (N_24194,N_20293,N_21017);
or U24195 (N_24195,N_20650,N_19298);
nor U24196 (N_24196,N_18822,N_19946);
nand U24197 (N_24197,N_20042,N_21702);
or U24198 (N_24198,N_18812,N_21196);
and U24199 (N_24199,N_20952,N_19976);
nor U24200 (N_24200,N_19440,N_21747);
nor U24201 (N_24201,N_20716,N_18896);
and U24202 (N_24202,N_19655,N_21442);
nand U24203 (N_24203,N_20663,N_18773);
xnor U24204 (N_24204,N_18822,N_19232);
or U24205 (N_24205,N_19082,N_21268);
nand U24206 (N_24206,N_19850,N_21110);
and U24207 (N_24207,N_21282,N_21232);
xor U24208 (N_24208,N_20223,N_20937);
or U24209 (N_24209,N_20167,N_19547);
and U24210 (N_24210,N_21043,N_19066);
and U24211 (N_24211,N_19617,N_21650);
or U24212 (N_24212,N_21510,N_18795);
or U24213 (N_24213,N_21873,N_21506);
nand U24214 (N_24214,N_20767,N_19947);
nor U24215 (N_24215,N_21777,N_19127);
or U24216 (N_24216,N_21594,N_21755);
and U24217 (N_24217,N_19578,N_21779);
and U24218 (N_24218,N_19199,N_21032);
nand U24219 (N_24219,N_21492,N_19329);
and U24220 (N_24220,N_18815,N_19614);
nor U24221 (N_24221,N_19239,N_19448);
nor U24222 (N_24222,N_21377,N_18789);
and U24223 (N_24223,N_19348,N_21682);
or U24224 (N_24224,N_21558,N_19480);
and U24225 (N_24225,N_20885,N_21693);
nor U24226 (N_24226,N_19732,N_18801);
nand U24227 (N_24227,N_19590,N_20008);
and U24228 (N_24228,N_19535,N_21614);
nor U24229 (N_24229,N_20358,N_20498);
xor U24230 (N_24230,N_19818,N_19711);
and U24231 (N_24231,N_20426,N_21042);
or U24232 (N_24232,N_21410,N_21315);
or U24233 (N_24233,N_19263,N_20834);
nor U24234 (N_24234,N_21462,N_19416);
nor U24235 (N_24235,N_19688,N_20371);
nor U24236 (N_24236,N_20062,N_20885);
and U24237 (N_24237,N_19304,N_20154);
and U24238 (N_24238,N_20974,N_20883);
nand U24239 (N_24239,N_19296,N_20333);
or U24240 (N_24240,N_19708,N_19285);
or U24241 (N_24241,N_21028,N_20837);
and U24242 (N_24242,N_20878,N_18848);
nor U24243 (N_24243,N_20501,N_21418);
nor U24244 (N_24244,N_19022,N_20372);
nand U24245 (N_24245,N_19025,N_18894);
nor U24246 (N_24246,N_21199,N_20033);
and U24247 (N_24247,N_18843,N_20773);
or U24248 (N_24248,N_20305,N_19178);
nor U24249 (N_24249,N_19252,N_19733);
nand U24250 (N_24250,N_19089,N_21339);
nand U24251 (N_24251,N_21496,N_20751);
and U24252 (N_24252,N_19823,N_20412);
and U24253 (N_24253,N_20878,N_19661);
nand U24254 (N_24254,N_20187,N_20069);
nor U24255 (N_24255,N_19127,N_21345);
nand U24256 (N_24256,N_20491,N_21043);
xnor U24257 (N_24257,N_20399,N_21715);
nor U24258 (N_24258,N_20545,N_19683);
or U24259 (N_24259,N_19236,N_21045);
nor U24260 (N_24260,N_20484,N_20912);
xnor U24261 (N_24261,N_21412,N_18901);
nand U24262 (N_24262,N_20818,N_21831);
or U24263 (N_24263,N_19258,N_19196);
nand U24264 (N_24264,N_19342,N_20395);
nor U24265 (N_24265,N_21307,N_21831);
nand U24266 (N_24266,N_21209,N_21380);
and U24267 (N_24267,N_20400,N_18801);
and U24268 (N_24268,N_21735,N_19541);
nand U24269 (N_24269,N_21515,N_20705);
nor U24270 (N_24270,N_20992,N_19402);
and U24271 (N_24271,N_19071,N_21095);
and U24272 (N_24272,N_19552,N_20859);
nand U24273 (N_24273,N_20677,N_19698);
nand U24274 (N_24274,N_19609,N_20358);
and U24275 (N_24275,N_20466,N_19071);
or U24276 (N_24276,N_18912,N_19363);
nand U24277 (N_24277,N_19941,N_19691);
or U24278 (N_24278,N_20001,N_19566);
nand U24279 (N_24279,N_20062,N_19497);
and U24280 (N_24280,N_18750,N_19430);
and U24281 (N_24281,N_19496,N_19548);
nor U24282 (N_24282,N_20714,N_21771);
xor U24283 (N_24283,N_19041,N_19877);
nor U24284 (N_24284,N_19852,N_21750);
and U24285 (N_24285,N_19808,N_21819);
and U24286 (N_24286,N_21298,N_18935);
nand U24287 (N_24287,N_20041,N_21224);
and U24288 (N_24288,N_20766,N_18971);
and U24289 (N_24289,N_21674,N_21804);
nand U24290 (N_24290,N_21860,N_21717);
nand U24291 (N_24291,N_19862,N_19457);
nor U24292 (N_24292,N_21624,N_19391);
and U24293 (N_24293,N_21066,N_20928);
nand U24294 (N_24294,N_18966,N_20482);
and U24295 (N_24295,N_21351,N_18818);
or U24296 (N_24296,N_19418,N_20592);
nand U24297 (N_24297,N_20061,N_19624);
nor U24298 (N_24298,N_19050,N_19612);
nand U24299 (N_24299,N_19485,N_21646);
nand U24300 (N_24300,N_21198,N_18827);
or U24301 (N_24301,N_18770,N_18786);
nor U24302 (N_24302,N_19252,N_19646);
or U24303 (N_24303,N_19007,N_20924);
nor U24304 (N_24304,N_20851,N_20252);
nand U24305 (N_24305,N_18755,N_19160);
nand U24306 (N_24306,N_20277,N_20944);
nand U24307 (N_24307,N_20803,N_21504);
and U24308 (N_24308,N_20691,N_19219);
nor U24309 (N_24309,N_21639,N_21550);
nor U24310 (N_24310,N_21677,N_21405);
nand U24311 (N_24311,N_18772,N_20409);
nand U24312 (N_24312,N_20700,N_20742);
nor U24313 (N_24313,N_19434,N_21842);
or U24314 (N_24314,N_21364,N_19003);
and U24315 (N_24315,N_19116,N_21081);
nand U24316 (N_24316,N_21106,N_21418);
or U24317 (N_24317,N_19193,N_19500);
nand U24318 (N_24318,N_20515,N_21344);
and U24319 (N_24319,N_21367,N_21673);
or U24320 (N_24320,N_20943,N_19524);
and U24321 (N_24321,N_20446,N_21518);
nor U24322 (N_24322,N_20858,N_20824);
nor U24323 (N_24323,N_21795,N_20282);
nor U24324 (N_24324,N_19740,N_20932);
nor U24325 (N_24325,N_21024,N_21772);
or U24326 (N_24326,N_19602,N_20290);
and U24327 (N_24327,N_21256,N_21665);
or U24328 (N_24328,N_19727,N_21377);
or U24329 (N_24329,N_19954,N_19521);
nand U24330 (N_24330,N_19616,N_19433);
and U24331 (N_24331,N_19247,N_20808);
nor U24332 (N_24332,N_21074,N_21251);
nand U24333 (N_24333,N_20755,N_21723);
nand U24334 (N_24334,N_20267,N_21471);
nand U24335 (N_24335,N_19842,N_20492);
or U24336 (N_24336,N_20747,N_19726);
nor U24337 (N_24337,N_21744,N_20383);
nand U24338 (N_24338,N_19478,N_20188);
nor U24339 (N_24339,N_18794,N_20967);
nand U24340 (N_24340,N_20551,N_19332);
xor U24341 (N_24341,N_20614,N_21392);
nor U24342 (N_24342,N_21535,N_18981);
nor U24343 (N_24343,N_20946,N_20397);
or U24344 (N_24344,N_18789,N_19542);
nor U24345 (N_24345,N_21328,N_21262);
nor U24346 (N_24346,N_21838,N_19406);
and U24347 (N_24347,N_20159,N_18952);
nor U24348 (N_24348,N_19121,N_18907);
nand U24349 (N_24349,N_19427,N_20036);
and U24350 (N_24350,N_20311,N_21807);
nor U24351 (N_24351,N_20152,N_20108);
nor U24352 (N_24352,N_21776,N_21609);
nand U24353 (N_24353,N_19731,N_18786);
or U24354 (N_24354,N_20166,N_20369);
nor U24355 (N_24355,N_18907,N_19379);
nor U24356 (N_24356,N_18902,N_21746);
or U24357 (N_24357,N_20054,N_20728);
xnor U24358 (N_24358,N_20593,N_19227);
and U24359 (N_24359,N_21675,N_18990);
nand U24360 (N_24360,N_20024,N_20160);
nand U24361 (N_24361,N_20460,N_19086);
or U24362 (N_24362,N_19102,N_19762);
or U24363 (N_24363,N_19285,N_20262);
xor U24364 (N_24364,N_18979,N_18900);
or U24365 (N_24365,N_20210,N_19674);
nand U24366 (N_24366,N_21407,N_19648);
nand U24367 (N_24367,N_20784,N_20729);
and U24368 (N_24368,N_19976,N_20533);
nor U24369 (N_24369,N_19492,N_19952);
xor U24370 (N_24370,N_19444,N_19148);
nand U24371 (N_24371,N_21369,N_19130);
or U24372 (N_24372,N_19546,N_19016);
nor U24373 (N_24373,N_20385,N_21259);
nand U24374 (N_24374,N_21044,N_20521);
nor U24375 (N_24375,N_20936,N_20450);
nor U24376 (N_24376,N_21234,N_20371);
or U24377 (N_24377,N_19376,N_20984);
nand U24378 (N_24378,N_20439,N_21078);
and U24379 (N_24379,N_21645,N_19541);
xnor U24380 (N_24380,N_18861,N_20314);
nand U24381 (N_24381,N_20976,N_20127);
nor U24382 (N_24382,N_20346,N_21848);
nor U24383 (N_24383,N_18872,N_19036);
or U24384 (N_24384,N_21342,N_20907);
and U24385 (N_24385,N_19512,N_21311);
nand U24386 (N_24386,N_21413,N_21654);
or U24387 (N_24387,N_21607,N_19620);
or U24388 (N_24388,N_21753,N_20930);
or U24389 (N_24389,N_19271,N_19540);
or U24390 (N_24390,N_20076,N_19148);
nand U24391 (N_24391,N_20453,N_21202);
or U24392 (N_24392,N_20388,N_19658);
xnor U24393 (N_24393,N_20410,N_19443);
or U24394 (N_24394,N_20771,N_21543);
nor U24395 (N_24395,N_20661,N_21280);
nor U24396 (N_24396,N_21351,N_18750);
nand U24397 (N_24397,N_20184,N_20221);
nand U24398 (N_24398,N_19192,N_19695);
nand U24399 (N_24399,N_21170,N_19461);
nor U24400 (N_24400,N_21209,N_21153);
nor U24401 (N_24401,N_20455,N_21489);
and U24402 (N_24402,N_21182,N_19099);
xor U24403 (N_24403,N_19881,N_21863);
nand U24404 (N_24404,N_20671,N_20723);
or U24405 (N_24405,N_18842,N_20035);
or U24406 (N_24406,N_19722,N_19366);
xor U24407 (N_24407,N_19658,N_20776);
xor U24408 (N_24408,N_20275,N_19597);
or U24409 (N_24409,N_20659,N_21083);
or U24410 (N_24410,N_19898,N_21017);
nand U24411 (N_24411,N_20584,N_19726);
or U24412 (N_24412,N_21708,N_20048);
or U24413 (N_24413,N_19253,N_21653);
nand U24414 (N_24414,N_19691,N_20593);
nor U24415 (N_24415,N_20110,N_19502);
and U24416 (N_24416,N_21490,N_20936);
nor U24417 (N_24417,N_20776,N_20568);
and U24418 (N_24418,N_21782,N_20695);
and U24419 (N_24419,N_20350,N_19482);
nand U24420 (N_24420,N_19032,N_21722);
nor U24421 (N_24421,N_21740,N_20780);
and U24422 (N_24422,N_21090,N_20321);
nor U24423 (N_24423,N_19914,N_19034);
or U24424 (N_24424,N_20808,N_21551);
or U24425 (N_24425,N_21245,N_20788);
nand U24426 (N_24426,N_21852,N_20775);
nand U24427 (N_24427,N_20775,N_21794);
and U24428 (N_24428,N_19622,N_19159);
and U24429 (N_24429,N_19577,N_18958);
or U24430 (N_24430,N_19488,N_19364);
nor U24431 (N_24431,N_21412,N_20704);
nand U24432 (N_24432,N_21616,N_21674);
nor U24433 (N_24433,N_21622,N_21129);
or U24434 (N_24434,N_21086,N_19612);
or U24435 (N_24435,N_19018,N_19632);
or U24436 (N_24436,N_19720,N_19895);
and U24437 (N_24437,N_21390,N_19370);
nor U24438 (N_24438,N_21684,N_20295);
nand U24439 (N_24439,N_19947,N_19993);
or U24440 (N_24440,N_20525,N_20566);
and U24441 (N_24441,N_18828,N_18893);
and U24442 (N_24442,N_20071,N_19898);
nor U24443 (N_24443,N_20766,N_20865);
or U24444 (N_24444,N_20555,N_21147);
and U24445 (N_24445,N_21675,N_18763);
nand U24446 (N_24446,N_20412,N_18925);
or U24447 (N_24447,N_19507,N_19109);
nand U24448 (N_24448,N_18791,N_20070);
xnor U24449 (N_24449,N_20655,N_21178);
or U24450 (N_24450,N_20303,N_20565);
and U24451 (N_24451,N_20929,N_21595);
or U24452 (N_24452,N_21239,N_20226);
and U24453 (N_24453,N_18814,N_20466);
nand U24454 (N_24454,N_19638,N_19786);
xor U24455 (N_24455,N_18795,N_19484);
xnor U24456 (N_24456,N_19512,N_19393);
xor U24457 (N_24457,N_19631,N_21667);
xnor U24458 (N_24458,N_19405,N_19508);
xor U24459 (N_24459,N_20401,N_19551);
xor U24460 (N_24460,N_20462,N_18975);
or U24461 (N_24461,N_20747,N_19566);
nor U24462 (N_24462,N_19615,N_20602);
nand U24463 (N_24463,N_19126,N_19911);
nand U24464 (N_24464,N_20677,N_20884);
or U24465 (N_24465,N_21645,N_20080);
nor U24466 (N_24466,N_21662,N_20106);
and U24467 (N_24467,N_20954,N_20117);
nand U24468 (N_24468,N_19308,N_20501);
nor U24469 (N_24469,N_21309,N_21335);
xor U24470 (N_24470,N_19460,N_21174);
xnor U24471 (N_24471,N_21869,N_20808);
nor U24472 (N_24472,N_19015,N_18922);
or U24473 (N_24473,N_19075,N_20687);
and U24474 (N_24474,N_19105,N_21273);
or U24475 (N_24475,N_20859,N_19409);
or U24476 (N_24476,N_21768,N_20136);
nand U24477 (N_24477,N_21479,N_20551);
or U24478 (N_24478,N_20413,N_20530);
and U24479 (N_24479,N_19101,N_20363);
or U24480 (N_24480,N_20836,N_19101);
and U24481 (N_24481,N_19757,N_19471);
nor U24482 (N_24482,N_19107,N_20066);
nor U24483 (N_24483,N_21164,N_20053);
or U24484 (N_24484,N_20992,N_20678);
and U24485 (N_24485,N_20853,N_19369);
nand U24486 (N_24486,N_21339,N_19983);
nor U24487 (N_24487,N_20717,N_20876);
xor U24488 (N_24488,N_20343,N_20162);
nor U24489 (N_24489,N_20976,N_20830);
and U24490 (N_24490,N_19346,N_20517);
nand U24491 (N_24491,N_21669,N_19940);
nor U24492 (N_24492,N_21103,N_21251);
xnor U24493 (N_24493,N_20666,N_19439);
and U24494 (N_24494,N_19209,N_20157);
nor U24495 (N_24495,N_19489,N_20702);
nor U24496 (N_24496,N_19979,N_19996);
and U24497 (N_24497,N_19687,N_21403);
xnor U24498 (N_24498,N_19743,N_19502);
or U24499 (N_24499,N_21376,N_18799);
and U24500 (N_24500,N_19395,N_20091);
nand U24501 (N_24501,N_19174,N_19359);
nor U24502 (N_24502,N_19102,N_19127);
and U24503 (N_24503,N_19543,N_20695);
or U24504 (N_24504,N_19444,N_19067);
or U24505 (N_24505,N_19921,N_19210);
nand U24506 (N_24506,N_20004,N_18812);
or U24507 (N_24507,N_20996,N_19905);
and U24508 (N_24508,N_20912,N_20592);
and U24509 (N_24509,N_21048,N_21549);
nand U24510 (N_24510,N_19983,N_21219);
nand U24511 (N_24511,N_19954,N_20328);
xor U24512 (N_24512,N_21474,N_21563);
nor U24513 (N_24513,N_19775,N_21771);
nor U24514 (N_24514,N_21136,N_21019);
or U24515 (N_24515,N_20418,N_18932);
or U24516 (N_24516,N_19387,N_18809);
nand U24517 (N_24517,N_20096,N_21830);
and U24518 (N_24518,N_18977,N_19172);
and U24519 (N_24519,N_20413,N_20325);
nor U24520 (N_24520,N_20382,N_19906);
nand U24521 (N_24521,N_21735,N_19055);
or U24522 (N_24522,N_21089,N_18977);
nor U24523 (N_24523,N_21247,N_20476);
nand U24524 (N_24524,N_20188,N_19538);
nor U24525 (N_24525,N_20656,N_20222);
xnor U24526 (N_24526,N_21471,N_18913);
nor U24527 (N_24527,N_21787,N_20058);
or U24528 (N_24528,N_20616,N_21533);
xnor U24529 (N_24529,N_19823,N_21062);
nor U24530 (N_24530,N_18786,N_18965);
or U24531 (N_24531,N_21614,N_19628);
nand U24532 (N_24532,N_20167,N_21501);
nor U24533 (N_24533,N_20455,N_21389);
nor U24534 (N_24534,N_20707,N_19322);
or U24535 (N_24535,N_21239,N_21839);
and U24536 (N_24536,N_21689,N_20985);
nor U24537 (N_24537,N_21180,N_19499);
nor U24538 (N_24538,N_21179,N_18758);
or U24539 (N_24539,N_21001,N_19160);
nor U24540 (N_24540,N_20420,N_19559);
nand U24541 (N_24541,N_20949,N_21314);
nand U24542 (N_24542,N_20778,N_21695);
nor U24543 (N_24543,N_20640,N_18872);
and U24544 (N_24544,N_19767,N_21406);
nand U24545 (N_24545,N_18755,N_21403);
or U24546 (N_24546,N_20291,N_20091);
xnor U24547 (N_24547,N_19145,N_19236);
nand U24548 (N_24548,N_19190,N_20963);
nor U24549 (N_24549,N_21169,N_20315);
and U24550 (N_24550,N_21643,N_21410);
xnor U24551 (N_24551,N_19214,N_20125);
nor U24552 (N_24552,N_19399,N_19645);
nor U24553 (N_24553,N_21127,N_21216);
or U24554 (N_24554,N_20535,N_20541);
or U24555 (N_24555,N_21150,N_19046);
and U24556 (N_24556,N_20231,N_19190);
nand U24557 (N_24557,N_21410,N_19674);
and U24558 (N_24558,N_19779,N_19848);
or U24559 (N_24559,N_19809,N_19504);
nand U24560 (N_24560,N_19175,N_21292);
nand U24561 (N_24561,N_21154,N_20625);
nor U24562 (N_24562,N_19116,N_19819);
nand U24563 (N_24563,N_21012,N_18896);
nor U24564 (N_24564,N_21656,N_19874);
xnor U24565 (N_24565,N_19994,N_21199);
xor U24566 (N_24566,N_19919,N_19093);
nand U24567 (N_24567,N_20938,N_21226);
nor U24568 (N_24568,N_21075,N_20987);
and U24569 (N_24569,N_20320,N_18932);
nor U24570 (N_24570,N_21571,N_19510);
nand U24571 (N_24571,N_21247,N_19841);
and U24572 (N_24572,N_20576,N_19235);
and U24573 (N_24573,N_19801,N_19076);
nor U24574 (N_24574,N_21589,N_20694);
nor U24575 (N_24575,N_21362,N_21315);
nor U24576 (N_24576,N_21838,N_20457);
or U24577 (N_24577,N_21868,N_20386);
nand U24578 (N_24578,N_19899,N_19380);
nor U24579 (N_24579,N_19812,N_20130);
nor U24580 (N_24580,N_21694,N_21717);
nand U24581 (N_24581,N_20150,N_20563);
nor U24582 (N_24582,N_21007,N_19574);
and U24583 (N_24583,N_20461,N_21554);
nand U24584 (N_24584,N_21078,N_19111);
nor U24585 (N_24585,N_18760,N_19370);
nand U24586 (N_24586,N_19942,N_20209);
nand U24587 (N_24587,N_21232,N_20346);
or U24588 (N_24588,N_19874,N_21006);
and U24589 (N_24589,N_21562,N_20724);
or U24590 (N_24590,N_19350,N_21274);
nand U24591 (N_24591,N_19018,N_20635);
or U24592 (N_24592,N_20398,N_21786);
nor U24593 (N_24593,N_19735,N_20852);
and U24594 (N_24594,N_19984,N_20097);
or U24595 (N_24595,N_21064,N_21767);
and U24596 (N_24596,N_19933,N_21476);
nor U24597 (N_24597,N_20915,N_19949);
or U24598 (N_24598,N_21561,N_20265);
nand U24599 (N_24599,N_21605,N_20314);
nor U24600 (N_24600,N_18999,N_21026);
and U24601 (N_24601,N_18980,N_21760);
nand U24602 (N_24602,N_18846,N_18882);
or U24603 (N_24603,N_20142,N_21584);
nor U24604 (N_24604,N_21813,N_20965);
and U24605 (N_24605,N_20718,N_21310);
and U24606 (N_24606,N_20948,N_20359);
nand U24607 (N_24607,N_19712,N_19252);
or U24608 (N_24608,N_20248,N_19077);
and U24609 (N_24609,N_19486,N_19266);
xor U24610 (N_24610,N_19302,N_19891);
or U24611 (N_24611,N_21578,N_19247);
nor U24612 (N_24612,N_20813,N_19577);
or U24613 (N_24613,N_20599,N_18958);
or U24614 (N_24614,N_19209,N_18838);
or U24615 (N_24615,N_19873,N_19707);
and U24616 (N_24616,N_20543,N_20026);
xnor U24617 (N_24617,N_21457,N_19152);
nand U24618 (N_24618,N_20874,N_20800);
and U24619 (N_24619,N_21658,N_20408);
nand U24620 (N_24620,N_18923,N_19469);
nor U24621 (N_24621,N_19360,N_21723);
and U24622 (N_24622,N_20936,N_21812);
nor U24623 (N_24623,N_20844,N_21873);
or U24624 (N_24624,N_19665,N_19887);
nand U24625 (N_24625,N_20804,N_19466);
xnor U24626 (N_24626,N_18872,N_19501);
nand U24627 (N_24627,N_20911,N_20006);
and U24628 (N_24628,N_20510,N_20155);
nand U24629 (N_24629,N_21296,N_20810);
nand U24630 (N_24630,N_20042,N_20136);
nand U24631 (N_24631,N_20819,N_18829);
or U24632 (N_24632,N_19845,N_18958);
nor U24633 (N_24633,N_19722,N_19042);
nor U24634 (N_24634,N_21131,N_21830);
and U24635 (N_24635,N_19837,N_21503);
or U24636 (N_24636,N_20758,N_20614);
nor U24637 (N_24637,N_19437,N_20758);
nor U24638 (N_24638,N_20501,N_19163);
nor U24639 (N_24639,N_21791,N_21856);
or U24640 (N_24640,N_20676,N_20333);
nor U24641 (N_24641,N_21532,N_20571);
nand U24642 (N_24642,N_19625,N_20119);
or U24643 (N_24643,N_20696,N_20185);
and U24644 (N_24644,N_20938,N_20426);
xor U24645 (N_24645,N_21274,N_20830);
or U24646 (N_24646,N_21768,N_21124);
and U24647 (N_24647,N_18750,N_21238);
nand U24648 (N_24648,N_21785,N_19098);
nand U24649 (N_24649,N_20580,N_20596);
or U24650 (N_24650,N_19021,N_21464);
nand U24651 (N_24651,N_19926,N_21529);
nor U24652 (N_24652,N_21197,N_20724);
and U24653 (N_24653,N_18898,N_21397);
nand U24654 (N_24654,N_21635,N_20525);
or U24655 (N_24655,N_21078,N_20061);
nand U24656 (N_24656,N_20160,N_18825);
or U24657 (N_24657,N_20594,N_20837);
or U24658 (N_24658,N_18815,N_18869);
nand U24659 (N_24659,N_19294,N_21400);
nor U24660 (N_24660,N_21533,N_19962);
nor U24661 (N_24661,N_21424,N_20017);
or U24662 (N_24662,N_19700,N_20787);
nor U24663 (N_24663,N_20653,N_19289);
nor U24664 (N_24664,N_19502,N_18767);
nand U24665 (N_24665,N_21731,N_20216);
nand U24666 (N_24666,N_19025,N_19834);
nor U24667 (N_24667,N_20777,N_20663);
nand U24668 (N_24668,N_20862,N_19473);
or U24669 (N_24669,N_20977,N_20701);
xnor U24670 (N_24670,N_19838,N_19119);
and U24671 (N_24671,N_20395,N_20276);
nor U24672 (N_24672,N_21262,N_19535);
or U24673 (N_24673,N_19629,N_18824);
and U24674 (N_24674,N_19392,N_21148);
nand U24675 (N_24675,N_19584,N_18830);
nand U24676 (N_24676,N_20019,N_21212);
nor U24677 (N_24677,N_20441,N_19027);
nand U24678 (N_24678,N_19243,N_21484);
nand U24679 (N_24679,N_21030,N_21740);
nand U24680 (N_24680,N_20463,N_21143);
or U24681 (N_24681,N_19108,N_19278);
nor U24682 (N_24682,N_21220,N_21442);
nor U24683 (N_24683,N_19107,N_19474);
and U24684 (N_24684,N_21867,N_19954);
and U24685 (N_24685,N_20577,N_21031);
nor U24686 (N_24686,N_20123,N_20111);
nor U24687 (N_24687,N_21109,N_21691);
and U24688 (N_24688,N_18899,N_20872);
and U24689 (N_24689,N_18782,N_21478);
nand U24690 (N_24690,N_21175,N_20345);
and U24691 (N_24691,N_19358,N_20321);
nor U24692 (N_24692,N_19415,N_21688);
nor U24693 (N_24693,N_19529,N_20243);
xor U24694 (N_24694,N_19175,N_19190);
and U24695 (N_24695,N_19343,N_19444);
and U24696 (N_24696,N_20216,N_19794);
and U24697 (N_24697,N_19032,N_19977);
and U24698 (N_24698,N_20527,N_21337);
nand U24699 (N_24699,N_20537,N_21446);
or U24700 (N_24700,N_21064,N_19117);
or U24701 (N_24701,N_21734,N_18792);
or U24702 (N_24702,N_21625,N_20457);
and U24703 (N_24703,N_20425,N_20864);
nor U24704 (N_24704,N_19938,N_19916);
nand U24705 (N_24705,N_21187,N_19550);
nor U24706 (N_24706,N_18890,N_21592);
nor U24707 (N_24707,N_18877,N_20886);
and U24708 (N_24708,N_21778,N_21607);
and U24709 (N_24709,N_21441,N_19937);
and U24710 (N_24710,N_20408,N_21618);
nor U24711 (N_24711,N_21650,N_19878);
nor U24712 (N_24712,N_21742,N_20122);
nand U24713 (N_24713,N_19961,N_19024);
and U24714 (N_24714,N_19754,N_19919);
nor U24715 (N_24715,N_19536,N_19267);
xnor U24716 (N_24716,N_20751,N_18943);
nand U24717 (N_24717,N_19561,N_18840);
nor U24718 (N_24718,N_19175,N_19184);
nor U24719 (N_24719,N_21564,N_20520);
or U24720 (N_24720,N_20351,N_21217);
and U24721 (N_24721,N_19195,N_21817);
nor U24722 (N_24722,N_21099,N_19889);
nand U24723 (N_24723,N_19089,N_20767);
nand U24724 (N_24724,N_20679,N_20155);
and U24725 (N_24725,N_18898,N_19461);
nor U24726 (N_24726,N_21201,N_21463);
nor U24727 (N_24727,N_20004,N_19844);
or U24728 (N_24728,N_18824,N_19626);
and U24729 (N_24729,N_20097,N_20329);
or U24730 (N_24730,N_19081,N_21147);
nor U24731 (N_24731,N_18794,N_20530);
nor U24732 (N_24732,N_19406,N_21536);
nand U24733 (N_24733,N_19766,N_21732);
nand U24734 (N_24734,N_20909,N_20536);
or U24735 (N_24735,N_20958,N_19949);
nor U24736 (N_24736,N_19425,N_19620);
xor U24737 (N_24737,N_21770,N_19603);
or U24738 (N_24738,N_19328,N_20686);
nor U24739 (N_24739,N_19676,N_19735);
xnor U24740 (N_24740,N_19771,N_20542);
nand U24741 (N_24741,N_21213,N_20118);
nand U24742 (N_24742,N_20970,N_20755);
nor U24743 (N_24743,N_21456,N_20826);
nand U24744 (N_24744,N_20360,N_21302);
or U24745 (N_24745,N_21261,N_18807);
and U24746 (N_24746,N_19072,N_21846);
and U24747 (N_24747,N_19783,N_19716);
nand U24748 (N_24748,N_19478,N_21544);
or U24749 (N_24749,N_19562,N_18922);
or U24750 (N_24750,N_19681,N_20946);
or U24751 (N_24751,N_21311,N_21494);
nor U24752 (N_24752,N_19813,N_20824);
or U24753 (N_24753,N_20038,N_20853);
nor U24754 (N_24754,N_19227,N_19613);
nand U24755 (N_24755,N_21153,N_21611);
and U24756 (N_24756,N_20805,N_21363);
or U24757 (N_24757,N_20404,N_21530);
nand U24758 (N_24758,N_20644,N_19843);
and U24759 (N_24759,N_19468,N_19097);
and U24760 (N_24760,N_20342,N_21332);
nand U24761 (N_24761,N_20592,N_21602);
and U24762 (N_24762,N_18757,N_20280);
or U24763 (N_24763,N_19847,N_20514);
nand U24764 (N_24764,N_19445,N_20207);
nand U24765 (N_24765,N_19400,N_19255);
and U24766 (N_24766,N_21132,N_21283);
nor U24767 (N_24767,N_21315,N_21671);
xor U24768 (N_24768,N_20895,N_20722);
or U24769 (N_24769,N_20114,N_19836);
xnor U24770 (N_24770,N_19998,N_20082);
nand U24771 (N_24771,N_20977,N_20330);
or U24772 (N_24772,N_18880,N_19691);
or U24773 (N_24773,N_18796,N_19329);
nor U24774 (N_24774,N_21855,N_18849);
or U24775 (N_24775,N_20274,N_21349);
nand U24776 (N_24776,N_19708,N_19906);
xor U24777 (N_24777,N_21390,N_21209);
and U24778 (N_24778,N_19998,N_21040);
nor U24779 (N_24779,N_18900,N_21167);
or U24780 (N_24780,N_20007,N_20874);
or U24781 (N_24781,N_21604,N_20470);
or U24782 (N_24782,N_19702,N_20713);
and U24783 (N_24783,N_21776,N_18836);
nor U24784 (N_24784,N_21619,N_20504);
and U24785 (N_24785,N_21739,N_21620);
nor U24786 (N_24786,N_19268,N_21187);
or U24787 (N_24787,N_20705,N_20450);
nand U24788 (N_24788,N_21118,N_19656);
nor U24789 (N_24789,N_20479,N_20604);
and U24790 (N_24790,N_20747,N_18934);
xor U24791 (N_24791,N_19029,N_19469);
or U24792 (N_24792,N_21768,N_18786);
nor U24793 (N_24793,N_19025,N_20328);
or U24794 (N_24794,N_19858,N_21568);
nor U24795 (N_24795,N_19047,N_19121);
or U24796 (N_24796,N_19471,N_19899);
nor U24797 (N_24797,N_21053,N_20532);
nor U24798 (N_24798,N_19479,N_19014);
or U24799 (N_24799,N_19752,N_19588);
nand U24800 (N_24800,N_21330,N_18851);
or U24801 (N_24801,N_21721,N_21530);
nand U24802 (N_24802,N_19429,N_20160);
nor U24803 (N_24803,N_21318,N_21475);
nand U24804 (N_24804,N_18898,N_19692);
and U24805 (N_24805,N_21778,N_21319);
nand U24806 (N_24806,N_19435,N_19417);
or U24807 (N_24807,N_20886,N_19359);
and U24808 (N_24808,N_21682,N_20199);
or U24809 (N_24809,N_21483,N_21217);
or U24810 (N_24810,N_20104,N_20000);
xnor U24811 (N_24811,N_18884,N_18942);
or U24812 (N_24812,N_19423,N_21672);
nand U24813 (N_24813,N_21423,N_19048);
nand U24814 (N_24814,N_19135,N_21311);
nor U24815 (N_24815,N_19699,N_20266);
xnor U24816 (N_24816,N_20227,N_21364);
nor U24817 (N_24817,N_21583,N_21782);
nand U24818 (N_24818,N_21695,N_21853);
or U24819 (N_24819,N_20245,N_19849);
nand U24820 (N_24820,N_21396,N_19822);
nand U24821 (N_24821,N_19101,N_19030);
nor U24822 (N_24822,N_19887,N_18884);
and U24823 (N_24823,N_21842,N_19180);
xor U24824 (N_24824,N_20485,N_21270);
or U24825 (N_24825,N_20294,N_21690);
nand U24826 (N_24826,N_21558,N_20605);
nor U24827 (N_24827,N_20523,N_19566);
nor U24828 (N_24828,N_21162,N_21658);
nand U24829 (N_24829,N_21785,N_19527);
nor U24830 (N_24830,N_20428,N_21234);
nor U24831 (N_24831,N_19973,N_20551);
nor U24832 (N_24832,N_21505,N_19363);
and U24833 (N_24833,N_20774,N_18913);
xnor U24834 (N_24834,N_18751,N_20799);
and U24835 (N_24835,N_18910,N_19255);
xnor U24836 (N_24836,N_21385,N_21459);
or U24837 (N_24837,N_21366,N_20699);
or U24838 (N_24838,N_20120,N_21287);
nor U24839 (N_24839,N_20833,N_20334);
nor U24840 (N_24840,N_20462,N_19415);
nor U24841 (N_24841,N_20559,N_21146);
nand U24842 (N_24842,N_21227,N_20993);
nor U24843 (N_24843,N_21135,N_19723);
and U24844 (N_24844,N_18803,N_19236);
nor U24845 (N_24845,N_19109,N_18758);
and U24846 (N_24846,N_20768,N_21492);
xnor U24847 (N_24847,N_20913,N_18890);
or U24848 (N_24848,N_19736,N_18773);
nand U24849 (N_24849,N_20427,N_18772);
xnor U24850 (N_24850,N_20454,N_19196);
and U24851 (N_24851,N_19424,N_21015);
and U24852 (N_24852,N_20406,N_18893);
nand U24853 (N_24853,N_19281,N_21629);
nand U24854 (N_24854,N_20676,N_20257);
and U24855 (N_24855,N_20521,N_20687);
nor U24856 (N_24856,N_20488,N_20845);
nand U24857 (N_24857,N_19589,N_19242);
xor U24858 (N_24858,N_19798,N_21258);
nand U24859 (N_24859,N_18789,N_20800);
or U24860 (N_24860,N_20059,N_20120);
nand U24861 (N_24861,N_21614,N_19980);
and U24862 (N_24862,N_18768,N_21581);
nor U24863 (N_24863,N_19700,N_19056);
or U24864 (N_24864,N_20224,N_21386);
nor U24865 (N_24865,N_21135,N_21505);
nor U24866 (N_24866,N_20253,N_19707);
nor U24867 (N_24867,N_20702,N_20814);
nand U24868 (N_24868,N_21132,N_20067);
or U24869 (N_24869,N_19084,N_21543);
nor U24870 (N_24870,N_21821,N_21541);
and U24871 (N_24871,N_18957,N_20158);
and U24872 (N_24872,N_18891,N_19584);
and U24873 (N_24873,N_19094,N_21112);
nor U24874 (N_24874,N_18901,N_20289);
and U24875 (N_24875,N_20252,N_20207);
nor U24876 (N_24876,N_19549,N_20831);
nor U24877 (N_24877,N_21666,N_18999);
nand U24878 (N_24878,N_19648,N_18901);
or U24879 (N_24879,N_21509,N_19565);
nor U24880 (N_24880,N_21404,N_20767);
xor U24881 (N_24881,N_20655,N_21167);
xor U24882 (N_24882,N_20534,N_20670);
nor U24883 (N_24883,N_19210,N_21740);
or U24884 (N_24884,N_20978,N_20247);
nor U24885 (N_24885,N_19987,N_21085);
and U24886 (N_24886,N_20204,N_19258);
nor U24887 (N_24887,N_19316,N_20401);
xnor U24888 (N_24888,N_20493,N_19220);
and U24889 (N_24889,N_21401,N_20658);
or U24890 (N_24890,N_20720,N_21296);
nor U24891 (N_24891,N_21349,N_18926);
nor U24892 (N_24892,N_21726,N_19890);
and U24893 (N_24893,N_19706,N_20517);
nor U24894 (N_24894,N_19873,N_19172);
or U24895 (N_24895,N_20597,N_20814);
nor U24896 (N_24896,N_18807,N_19445);
or U24897 (N_24897,N_19782,N_18956);
xnor U24898 (N_24898,N_20978,N_21011);
xnor U24899 (N_24899,N_19267,N_21311);
nor U24900 (N_24900,N_20157,N_19513);
and U24901 (N_24901,N_19896,N_20557);
or U24902 (N_24902,N_19628,N_20963);
xor U24903 (N_24903,N_20442,N_20383);
and U24904 (N_24904,N_20937,N_21658);
and U24905 (N_24905,N_20129,N_19033);
and U24906 (N_24906,N_20597,N_20382);
nor U24907 (N_24907,N_19730,N_19116);
and U24908 (N_24908,N_21568,N_21091);
xnor U24909 (N_24909,N_21498,N_19493);
nand U24910 (N_24910,N_20991,N_20872);
or U24911 (N_24911,N_19896,N_19324);
nand U24912 (N_24912,N_18911,N_20955);
xnor U24913 (N_24913,N_20622,N_18793);
nor U24914 (N_24914,N_20689,N_18988);
nand U24915 (N_24915,N_18831,N_19626);
or U24916 (N_24916,N_21639,N_21572);
xor U24917 (N_24917,N_19089,N_21866);
xor U24918 (N_24918,N_18841,N_20365);
or U24919 (N_24919,N_21524,N_21726);
nor U24920 (N_24920,N_21539,N_19501);
nor U24921 (N_24921,N_18906,N_19476);
nand U24922 (N_24922,N_19511,N_21694);
or U24923 (N_24923,N_20062,N_20586);
and U24924 (N_24924,N_19429,N_21812);
or U24925 (N_24925,N_20719,N_21794);
and U24926 (N_24926,N_20667,N_19737);
nor U24927 (N_24927,N_19905,N_20525);
nand U24928 (N_24928,N_20239,N_21318);
or U24929 (N_24929,N_19108,N_20686);
nor U24930 (N_24930,N_18766,N_20233);
xor U24931 (N_24931,N_19098,N_19332);
and U24932 (N_24932,N_21198,N_19598);
and U24933 (N_24933,N_19253,N_19237);
xnor U24934 (N_24934,N_18874,N_20680);
nor U24935 (N_24935,N_20039,N_20310);
nand U24936 (N_24936,N_20913,N_18847);
xnor U24937 (N_24937,N_19611,N_20413);
nor U24938 (N_24938,N_21510,N_19744);
nor U24939 (N_24939,N_18982,N_20363);
or U24940 (N_24940,N_20921,N_20796);
nor U24941 (N_24941,N_21570,N_19580);
nor U24942 (N_24942,N_18956,N_20383);
or U24943 (N_24943,N_20098,N_19099);
nand U24944 (N_24944,N_18899,N_21614);
nand U24945 (N_24945,N_20987,N_19960);
or U24946 (N_24946,N_20771,N_21125);
nand U24947 (N_24947,N_20144,N_20762);
nand U24948 (N_24948,N_20747,N_21137);
and U24949 (N_24949,N_20986,N_20787);
nor U24950 (N_24950,N_21737,N_20205);
nor U24951 (N_24951,N_20374,N_18872);
and U24952 (N_24952,N_21624,N_19755);
nor U24953 (N_24953,N_19415,N_20479);
nand U24954 (N_24954,N_21055,N_20250);
and U24955 (N_24955,N_19260,N_20303);
and U24956 (N_24956,N_21204,N_19089);
and U24957 (N_24957,N_19751,N_18896);
nand U24958 (N_24958,N_19442,N_21498);
nand U24959 (N_24959,N_21002,N_21439);
and U24960 (N_24960,N_21778,N_21385);
or U24961 (N_24961,N_20176,N_21537);
nor U24962 (N_24962,N_21196,N_19907);
nand U24963 (N_24963,N_20093,N_20012);
nand U24964 (N_24964,N_20588,N_19645);
and U24965 (N_24965,N_21839,N_19591);
or U24966 (N_24966,N_21841,N_20852);
nor U24967 (N_24967,N_19572,N_19629);
nor U24968 (N_24968,N_19820,N_21333);
xor U24969 (N_24969,N_20413,N_19984);
xnor U24970 (N_24970,N_19117,N_21808);
nand U24971 (N_24971,N_19583,N_21808);
and U24972 (N_24972,N_19616,N_21704);
and U24973 (N_24973,N_19214,N_19211);
nand U24974 (N_24974,N_21237,N_19882);
nor U24975 (N_24975,N_20723,N_21494);
and U24976 (N_24976,N_20506,N_20313);
xor U24977 (N_24977,N_19204,N_20813);
and U24978 (N_24978,N_19553,N_20065);
and U24979 (N_24979,N_21837,N_21150);
nor U24980 (N_24980,N_18753,N_21547);
and U24981 (N_24981,N_21445,N_20832);
nor U24982 (N_24982,N_18926,N_21814);
and U24983 (N_24983,N_21486,N_19275);
or U24984 (N_24984,N_21182,N_21026);
nor U24985 (N_24985,N_18940,N_21164);
nor U24986 (N_24986,N_19028,N_18902);
xor U24987 (N_24987,N_19212,N_19097);
nand U24988 (N_24988,N_20439,N_20463);
or U24989 (N_24989,N_19999,N_19847);
or U24990 (N_24990,N_21223,N_20155);
nand U24991 (N_24991,N_21133,N_20793);
or U24992 (N_24992,N_21713,N_20324);
nor U24993 (N_24993,N_20969,N_20384);
nand U24994 (N_24994,N_20833,N_20086);
nand U24995 (N_24995,N_20297,N_20875);
and U24996 (N_24996,N_19680,N_19431);
nand U24997 (N_24997,N_19005,N_19210);
nor U24998 (N_24998,N_21788,N_20259);
nor U24999 (N_24999,N_21207,N_19593);
and UO_0 (O_0,N_22742,N_24627);
nor UO_1 (O_1,N_24340,N_24227);
nand UO_2 (O_2,N_24349,N_24824);
and UO_3 (O_3,N_22616,N_22037);
or UO_4 (O_4,N_24393,N_23996);
and UO_5 (O_5,N_24555,N_23360);
nand UO_6 (O_6,N_23380,N_22850);
nor UO_7 (O_7,N_24209,N_22879);
nand UO_8 (O_8,N_24246,N_22552);
and UO_9 (O_9,N_24447,N_23340);
xor UO_10 (O_10,N_22886,N_22892);
nor UO_11 (O_11,N_23547,N_23636);
and UO_12 (O_12,N_22638,N_24752);
nor UO_13 (O_13,N_23918,N_22653);
nand UO_14 (O_14,N_21924,N_23704);
or UO_15 (O_15,N_24483,N_24879);
xor UO_16 (O_16,N_23400,N_22817);
xnor UO_17 (O_17,N_23011,N_22314);
nand UO_18 (O_18,N_24122,N_23222);
and UO_19 (O_19,N_24816,N_24945);
xnor UO_20 (O_20,N_23977,N_23248);
and UO_21 (O_21,N_22492,N_22421);
nor UO_22 (O_22,N_22231,N_22586);
and UO_23 (O_23,N_23438,N_22688);
nor UO_24 (O_24,N_24972,N_24705);
or UO_25 (O_25,N_23104,N_23127);
and UO_26 (O_26,N_22129,N_22385);
or UO_27 (O_27,N_23468,N_24360);
nand UO_28 (O_28,N_24158,N_24989);
nand UO_29 (O_29,N_24870,N_23243);
xnor UO_30 (O_30,N_22475,N_22065);
nand UO_31 (O_31,N_21931,N_22775);
and UO_32 (O_32,N_22063,N_23145);
and UO_33 (O_33,N_22789,N_24859);
or UO_34 (O_34,N_23413,N_22210);
or UO_35 (O_35,N_22652,N_23851);
and UO_36 (O_36,N_22570,N_24514);
and UO_37 (O_37,N_22936,N_24027);
or UO_38 (O_38,N_24445,N_22069);
or UO_39 (O_39,N_23003,N_24205);
nor UO_40 (O_40,N_23623,N_23303);
nand UO_41 (O_41,N_22643,N_22983);
nor UO_42 (O_42,N_22726,N_24755);
or UO_43 (O_43,N_21968,N_22790);
nor UO_44 (O_44,N_22128,N_24302);
or UO_45 (O_45,N_24381,N_24115);
and UO_46 (O_46,N_22373,N_24956);
nor UO_47 (O_47,N_22838,N_23184);
and UO_48 (O_48,N_23141,N_24839);
nand UO_49 (O_49,N_23812,N_23780);
nor UO_50 (O_50,N_22491,N_22016);
nor UO_51 (O_51,N_23496,N_24446);
xnor UO_52 (O_52,N_24012,N_24643);
nand UO_53 (O_53,N_22759,N_22771);
and UO_54 (O_54,N_23147,N_24440);
nor UO_55 (O_55,N_22162,N_24195);
nand UO_56 (O_56,N_21879,N_24907);
nand UO_57 (O_57,N_22914,N_22432);
nand UO_58 (O_58,N_24822,N_23566);
xnor UO_59 (O_59,N_24875,N_22609);
xor UO_60 (O_60,N_24920,N_23672);
and UO_61 (O_61,N_23832,N_22179);
and UO_62 (O_62,N_24644,N_23296);
xor UO_63 (O_63,N_22003,N_22085);
nor UO_64 (O_64,N_24186,N_21974);
nor UO_65 (O_65,N_23352,N_23447);
nor UO_66 (O_66,N_23856,N_24598);
nand UO_67 (O_67,N_22770,N_22345);
and UO_68 (O_68,N_24139,N_23526);
or UO_69 (O_69,N_22812,N_22090);
and UO_70 (O_70,N_24707,N_23047);
or UO_71 (O_71,N_22763,N_24862);
nor UO_72 (O_72,N_24547,N_22341);
or UO_73 (O_73,N_22571,N_23055);
nor UO_74 (O_74,N_24663,N_24404);
or UO_75 (O_75,N_22057,N_23992);
or UO_76 (O_76,N_22255,N_23207);
or UO_77 (O_77,N_24604,N_24935);
or UO_78 (O_78,N_22651,N_22306);
xor UO_79 (O_79,N_24024,N_23478);
nor UO_80 (O_80,N_22054,N_24680);
nor UO_81 (O_81,N_23988,N_24815);
and UO_82 (O_82,N_24224,N_23904);
or UO_83 (O_83,N_24917,N_23935);
and UO_84 (O_84,N_24350,N_23307);
nor UO_85 (O_85,N_22358,N_23186);
or UO_86 (O_86,N_24633,N_23588);
nand UO_87 (O_87,N_23975,N_22872);
and UO_88 (O_88,N_23870,N_24469);
or UO_89 (O_89,N_24387,N_23200);
nor UO_90 (O_90,N_22070,N_24743);
or UO_91 (O_91,N_24163,N_24911);
nor UO_92 (O_92,N_22693,N_23363);
nor UO_93 (O_93,N_23713,N_24339);
xnor UO_94 (O_94,N_22649,N_22041);
nand UO_95 (O_95,N_23225,N_24732);
and UO_96 (O_96,N_24476,N_22657);
nor UO_97 (O_97,N_22846,N_23523);
nand UO_98 (O_98,N_22758,N_22380);
nor UO_99 (O_99,N_24615,N_24317);
or UO_100 (O_100,N_22637,N_24579);
or UO_101 (O_101,N_24713,N_23040);
nand UO_102 (O_102,N_23203,N_24574);
nand UO_103 (O_103,N_22796,N_22225);
and UO_104 (O_104,N_24803,N_24528);
nand UO_105 (O_105,N_23686,N_22084);
xor UO_106 (O_106,N_24077,N_24379);
nor UO_107 (O_107,N_24482,N_23372);
nand UO_108 (O_108,N_24872,N_23113);
xor UO_109 (O_109,N_22988,N_22823);
nor UO_110 (O_110,N_22395,N_24303);
nor UO_111 (O_111,N_22815,N_23578);
nor UO_112 (O_112,N_22607,N_24973);
xnor UO_113 (O_113,N_22194,N_22059);
xor UO_114 (O_114,N_24398,N_24971);
or UO_115 (O_115,N_23181,N_23494);
nand UO_116 (O_116,N_23694,N_22707);
nor UO_117 (O_117,N_24606,N_22511);
nand UO_118 (O_118,N_24596,N_22066);
nand UO_119 (O_119,N_23375,N_24837);
nand UO_120 (O_120,N_23063,N_23072);
and UO_121 (O_121,N_23716,N_23917);
nand UO_122 (O_122,N_22159,N_24790);
nand UO_123 (O_123,N_23685,N_22347);
nand UO_124 (O_124,N_23095,N_22565);
nand UO_125 (O_125,N_23763,N_22064);
nor UO_126 (O_126,N_23934,N_22060);
nand UO_127 (O_127,N_23077,N_24638);
nor UO_128 (O_128,N_23241,N_24093);
or UO_129 (O_129,N_23673,N_24532);
nand UO_130 (O_130,N_23411,N_23240);
and UO_131 (O_131,N_22285,N_23530);
nand UO_132 (O_132,N_23056,N_21889);
xnor UO_133 (O_133,N_23555,N_22967);
nor UO_134 (O_134,N_22860,N_22020);
nor UO_135 (O_135,N_22836,N_23298);
nand UO_136 (O_136,N_22574,N_23345);
nand UO_137 (O_137,N_22767,N_22286);
or UO_138 (O_138,N_24289,N_24426);
xor UO_139 (O_139,N_22507,N_23632);
nor UO_140 (O_140,N_23471,N_24843);
nor UO_141 (O_141,N_24202,N_24054);
or UO_142 (O_142,N_24217,N_24133);
nor UO_143 (O_143,N_23013,N_23981);
nor UO_144 (O_144,N_24580,N_24614);
and UO_145 (O_145,N_23210,N_23289);
nor UO_146 (O_146,N_22221,N_23861);
nor UO_147 (O_147,N_23599,N_22546);
xor UO_148 (O_148,N_22046,N_22499);
and UO_149 (O_149,N_24085,N_22074);
nand UO_150 (O_150,N_22438,N_24556);
nand UO_151 (O_151,N_21921,N_22038);
nand UO_152 (O_152,N_23163,N_24320);
nor UO_153 (O_153,N_23052,N_22087);
nor UO_154 (O_154,N_23580,N_23852);
nor UO_155 (O_155,N_23785,N_22855);
nand UO_156 (O_156,N_24722,N_22120);
nand UO_157 (O_157,N_22029,N_24112);
nor UO_158 (O_158,N_22223,N_23754);
nor UO_159 (O_159,N_24052,N_22513);
or UO_160 (O_160,N_22163,N_23160);
nor UO_161 (O_161,N_22463,N_21998);
nand UO_162 (O_162,N_21878,N_24943);
or UO_163 (O_163,N_23059,N_22666);
nand UO_164 (O_164,N_23643,N_22361);
nand UO_165 (O_165,N_22542,N_22164);
xor UO_166 (O_166,N_23931,N_23415);
or UO_167 (O_167,N_23442,N_24549);
nand UO_168 (O_168,N_24661,N_24040);
nor UO_169 (O_169,N_22918,N_21991);
and UO_170 (O_170,N_23349,N_22308);
nand UO_171 (O_171,N_23841,N_24022);
nand UO_172 (O_172,N_23525,N_22601);
or UO_173 (O_173,N_23940,N_24364);
nand UO_174 (O_174,N_22449,N_22820);
nand UO_175 (O_175,N_24492,N_22311);
nor UO_176 (O_176,N_23477,N_21942);
nor UO_177 (O_177,N_24724,N_23058);
nand UO_178 (O_178,N_24279,N_23597);
nand UO_179 (O_179,N_24669,N_24094);
nor UO_180 (O_180,N_22590,N_22104);
nor UO_181 (O_181,N_24716,N_23993);
nor UO_182 (O_182,N_24278,N_24109);
nor UO_183 (O_183,N_24344,N_24503);
nor UO_184 (O_184,N_23221,N_24401);
nor UO_185 (O_185,N_22995,N_24455);
nor UO_186 (O_186,N_23882,N_24517);
and UO_187 (O_187,N_24590,N_24095);
xor UO_188 (O_188,N_22931,N_22960);
and UO_189 (O_189,N_22682,N_24102);
and UO_190 (O_190,N_22602,N_24070);
or UO_191 (O_191,N_23805,N_24641);
xor UO_192 (O_192,N_23959,N_23784);
xnor UO_193 (O_193,N_23026,N_22256);
nand UO_194 (O_194,N_22626,N_24586);
and UO_195 (O_195,N_22356,N_22920);
or UO_196 (O_196,N_24833,N_23769);
nor UO_197 (O_197,N_22460,N_23162);
or UO_198 (O_198,N_24846,N_24848);
or UO_199 (O_199,N_22955,N_24468);
and UO_200 (O_200,N_24096,N_22099);
nor UO_201 (O_201,N_24062,N_22088);
or UO_202 (O_202,N_23379,N_22719);
nor UO_203 (O_203,N_22991,N_22196);
or UO_204 (O_204,N_24648,N_23313);
and UO_205 (O_205,N_24939,N_22406);
nor UO_206 (O_206,N_24329,N_24380);
and UO_207 (O_207,N_22487,N_23822);
nor UO_208 (O_208,N_23164,N_22282);
nand UO_209 (O_209,N_22674,N_23393);
and UO_210 (O_210,N_23604,N_23327);
xor UO_211 (O_211,N_23895,N_22399);
and UO_212 (O_212,N_23342,N_22711);
nand UO_213 (O_213,N_24829,N_23860);
nor UO_214 (O_214,N_23844,N_22945);
xor UO_215 (O_215,N_24149,N_24220);
nor UO_216 (O_216,N_23647,N_23508);
nor UO_217 (O_217,N_24198,N_23741);
or UO_218 (O_218,N_22517,N_22611);
xnor UO_219 (O_219,N_23682,N_22414);
or UO_220 (O_220,N_22393,N_23625);
nand UO_221 (O_221,N_23253,N_23774);
or UO_222 (O_222,N_24739,N_22678);
nand UO_223 (O_223,N_24116,N_24565);
and UO_224 (O_224,N_21884,N_22524);
nor UO_225 (O_225,N_24348,N_23361);
nand UO_226 (O_226,N_24952,N_24073);
xnor UO_227 (O_227,N_24331,N_22808);
nor UO_228 (O_228,N_24229,N_23843);
nor UO_229 (O_229,N_23359,N_24250);
nor UO_230 (O_230,N_23835,N_24767);
or UO_231 (O_231,N_23326,N_24021);
xor UO_232 (O_232,N_23800,N_23041);
and UO_233 (O_233,N_24003,N_24106);
and UO_234 (O_234,N_24253,N_24536);
nor UO_235 (O_235,N_21905,N_22111);
nor UO_236 (O_236,N_24998,N_23907);
nor UO_237 (O_237,N_24028,N_24307);
and UO_238 (O_238,N_23767,N_23484);
nor UO_239 (O_239,N_24241,N_24740);
nand UO_240 (O_240,N_24927,N_24784);
and UO_241 (O_241,N_24113,N_23257);
nand UO_242 (O_242,N_23161,N_21926);
or UO_243 (O_243,N_22106,N_24899);
or UO_244 (O_244,N_22344,N_22644);
nand UO_245 (O_245,N_22854,N_22013);
nor UO_246 (O_246,N_24290,N_24554);
or UO_247 (O_247,N_23545,N_23266);
nand UO_248 (O_248,N_22576,N_22234);
nand UO_249 (O_249,N_24795,N_24761);
nor UO_250 (O_250,N_23126,N_21957);
nand UO_251 (O_251,N_24242,N_23902);
or UO_252 (O_252,N_22749,N_23914);
nand UO_253 (O_253,N_22833,N_22451);
nand UO_254 (O_254,N_22456,N_24612);
nand UO_255 (O_255,N_22252,N_22642);
or UO_256 (O_256,N_23699,N_24791);
nand UO_257 (O_257,N_21960,N_23620);
and UO_258 (O_258,N_23649,N_22009);
or UO_259 (O_259,N_24079,N_23725);
or UO_260 (O_260,N_23152,N_24655);
nor UO_261 (O_261,N_23574,N_24190);
nor UO_262 (O_262,N_22448,N_22587);
nand UO_263 (O_263,N_22509,N_23227);
nor UO_264 (O_264,N_23412,N_24014);
xnor UO_265 (O_265,N_22986,N_24423);
nor UO_266 (O_266,N_24637,N_23920);
or UO_267 (O_267,N_23416,N_23739);
nand UO_268 (O_268,N_24415,N_22025);
xnor UO_269 (O_269,N_22620,N_24805);
or UO_270 (O_270,N_23466,N_23370);
or UO_271 (O_271,N_21952,N_23842);
or UO_272 (O_272,N_24668,N_21969);
and UO_273 (O_273,N_24098,N_22948);
and UO_274 (O_274,N_22440,N_23974);
nand UO_275 (O_275,N_23051,N_23809);
or UO_276 (O_276,N_23553,N_24961);
nor UO_277 (O_277,N_23801,N_23758);
and UO_278 (O_278,N_23128,N_23123);
nor UO_279 (O_279,N_23770,N_22052);
or UO_280 (O_280,N_21915,N_23564);
nor UO_281 (O_281,N_23633,N_22785);
nor UO_282 (O_282,N_22868,N_24336);
nand UO_283 (O_283,N_22441,N_23964);
nand UO_284 (O_284,N_24315,N_24982);
or UO_285 (O_285,N_24474,N_24006);
and UO_286 (O_286,N_22301,N_22913);
and UO_287 (O_287,N_24558,N_22852);
or UO_288 (O_288,N_24311,N_23405);
nand UO_289 (O_289,N_23143,N_24660);
or UO_290 (O_290,N_22874,N_23621);
nor UO_291 (O_291,N_23869,N_24753);
nand UO_292 (O_292,N_22419,N_23718);
and UO_293 (O_293,N_23105,N_22275);
nand UO_294 (O_294,N_21927,N_24717);
nor UO_295 (O_295,N_22794,N_22553);
nor UO_296 (O_296,N_23541,N_24352);
nand UO_297 (O_297,N_22233,N_24161);
nor UO_298 (O_298,N_23590,N_23684);
or UO_299 (O_299,N_22376,N_23873);
nor UO_300 (O_300,N_24228,N_24518);
or UO_301 (O_301,N_24366,N_23775);
nand UO_302 (O_302,N_23369,N_23568);
or UO_303 (O_303,N_22632,N_24914);
xnor UO_304 (O_304,N_23060,N_22363);
xnor UO_305 (O_305,N_22381,N_23124);
or UO_306 (O_306,N_24891,N_22445);
nand UO_307 (O_307,N_23889,N_23006);
nor UO_308 (O_308,N_23378,N_22455);
nand UO_309 (O_309,N_22324,N_23776);
nand UO_310 (O_310,N_22318,N_22053);
nor UO_311 (O_311,N_24742,N_22782);
nand UO_312 (O_312,N_22636,N_21940);
or UO_313 (O_313,N_22189,N_23534);
nor UO_314 (O_314,N_22917,N_22335);
xor UO_315 (O_315,N_21914,N_21903);
nand UO_316 (O_316,N_23557,N_24799);
nand UO_317 (O_317,N_22488,N_24442);
nand UO_318 (O_318,N_24481,N_24673);
and UO_319 (O_319,N_23490,N_22689);
or UO_320 (O_320,N_22890,N_24847);
or UO_321 (O_321,N_23019,N_22199);
or UO_322 (O_322,N_24371,N_22472);
nor UO_323 (O_323,N_23323,N_23582);
nand UO_324 (O_324,N_23691,N_24788);
xnor UO_325 (O_325,N_21956,N_23936);
xor UO_326 (O_326,N_24658,N_23020);
nor UO_327 (O_327,N_22073,N_24811);
nand UO_328 (O_328,N_22984,N_24777);
or UO_329 (O_329,N_24312,N_24264);
nand UO_330 (O_330,N_23035,N_24208);
nand UO_331 (O_331,N_22110,N_23948);
xnor UO_332 (O_332,N_24817,N_24937);
or UO_333 (O_333,N_22180,N_23562);
nor UO_334 (O_334,N_24731,N_22898);
and UO_335 (O_335,N_24619,N_24223);
or UO_336 (O_336,N_22365,N_23023);
or UO_337 (O_337,N_23516,N_24293);
and UO_338 (O_338,N_23462,N_23337);
nor UO_339 (O_339,N_22504,N_23081);
or UO_340 (O_340,N_23884,N_24747);
and UO_341 (O_341,N_23973,N_23231);
or UO_342 (O_342,N_22271,N_24930);
nor UO_343 (O_343,N_22809,N_23666);
nand UO_344 (O_344,N_22989,N_22598);
nor UO_345 (O_345,N_24234,N_24038);
xnor UO_346 (O_346,N_23698,N_24061);
or UO_347 (O_347,N_24860,N_22394);
and UO_348 (O_348,N_24396,N_24804);
and UO_349 (O_349,N_22954,N_23137);
or UO_350 (O_350,N_24374,N_22869);
xnor UO_351 (O_351,N_23386,N_24613);
nor UO_352 (O_352,N_23083,N_22280);
nor UO_353 (O_353,N_22175,N_24258);
and UO_354 (O_354,N_24757,N_24871);
or UO_355 (O_355,N_24932,N_22412);
and UO_356 (O_356,N_23612,N_24996);
or UO_357 (O_357,N_22116,N_24268);
or UO_358 (O_358,N_22533,N_23573);
and UO_359 (O_359,N_24497,N_24051);
and UO_360 (O_360,N_24377,N_24715);
xor UO_361 (O_361,N_23978,N_22783);
nor UO_362 (O_362,N_22193,N_22780);
or UO_363 (O_363,N_24179,N_22924);
nand UO_364 (O_364,N_23249,N_22078);
nand UO_365 (O_365,N_24080,N_23219);
or UO_366 (O_366,N_22996,N_22095);
nand UO_367 (O_367,N_22981,N_23382);
nand UO_368 (O_368,N_23373,N_23663);
nand UO_369 (O_369,N_22937,N_21967);
nand UO_370 (O_370,N_24764,N_23333);
and UO_371 (O_371,N_24506,N_23979);
or UO_372 (O_372,N_22816,N_24391);
nand UO_373 (O_373,N_23836,N_24856);
or UO_374 (O_374,N_23662,N_24356);
nor UO_375 (O_375,N_22144,N_21961);
and UO_376 (O_376,N_24745,N_24894);
or UO_377 (O_377,N_22336,N_24560);
nand UO_378 (O_378,N_22811,N_22899);
nand UO_379 (O_379,N_22127,N_24050);
and UO_380 (O_380,N_22680,N_24520);
nand UO_381 (O_381,N_23505,N_22139);
nand UO_382 (O_382,N_24940,N_23492);
and UO_383 (O_383,N_22787,N_23328);
xor UO_384 (O_384,N_23130,N_22992);
nor UO_385 (O_385,N_23876,N_23034);
and UO_386 (O_386,N_22532,N_24187);
nor UO_387 (O_387,N_22182,N_24798);
nor UO_388 (O_388,N_22245,N_21916);
and UO_389 (O_389,N_24037,N_23753);
or UO_390 (O_390,N_24159,N_23661);
nand UO_391 (O_391,N_23433,N_24369);
and UO_392 (O_392,N_21930,N_22930);
and UO_393 (O_393,N_24591,N_22639);
and UO_394 (O_394,N_23700,N_22177);
and UO_395 (O_395,N_24402,N_23908);
xnor UO_396 (O_396,N_22908,N_23735);
nand UO_397 (O_397,N_23906,N_23239);
nor UO_398 (O_398,N_24428,N_22403);
or UO_399 (O_399,N_23454,N_22067);
or UO_400 (O_400,N_23456,N_22964);
nand UO_401 (O_401,N_24513,N_24295);
nand UO_402 (O_402,N_24886,N_22292);
nor UO_403 (O_403,N_22264,N_22606);
nor UO_404 (O_404,N_24047,N_22859);
and UO_405 (O_405,N_22858,N_23330);
nor UO_406 (O_406,N_22512,N_22980);
nor UO_407 (O_407,N_24162,N_21966);
or UO_408 (O_408,N_23571,N_22315);
and UO_409 (O_409,N_21938,N_24193);
and UO_410 (O_410,N_23781,N_23823);
nand UO_411 (O_411,N_22802,N_23358);
nor UO_412 (O_412,N_22251,N_24150);
nand UO_413 (O_413,N_22032,N_23391);
and UO_414 (O_414,N_22287,N_21897);
or UO_415 (O_415,N_23245,N_24548);
xnor UO_416 (O_416,N_23614,N_24792);
nand UO_417 (O_417,N_24001,N_24437);
or UO_418 (O_418,N_24723,N_22017);
and UO_419 (O_419,N_22728,N_24539);
nand UO_420 (O_420,N_24773,N_22244);
nor UO_421 (O_421,N_22993,N_23610);
and UO_422 (O_422,N_24738,N_22007);
nand UO_423 (O_423,N_24867,N_22550);
and UO_424 (O_424,N_24263,N_22466);
xnor UO_425 (O_425,N_24462,N_23616);
nand UO_426 (O_426,N_22962,N_22388);
nand UO_427 (O_427,N_23410,N_22841);
or UO_428 (O_428,N_24516,N_24679);
nand UO_429 (O_429,N_24009,N_23247);
nor UO_430 (O_430,N_24993,N_22378);
nand UO_431 (O_431,N_22061,N_22435);
nand UO_432 (O_432,N_22696,N_24921);
nor UO_433 (O_433,N_21964,N_22056);
nor UO_434 (O_434,N_23491,N_22765);
nor UO_435 (O_435,N_24509,N_23528);
xor UO_436 (O_436,N_21885,N_22648);
nand UO_437 (O_437,N_23251,N_23689);
nand UO_438 (O_438,N_24444,N_24775);
nor UO_439 (O_439,N_23444,N_23953);
nand UO_440 (O_440,N_22146,N_24168);
xnor UO_441 (O_441,N_22605,N_24372);
and UO_442 (O_442,N_22108,N_24178);
and UO_443 (O_443,N_22743,N_24039);
nand UO_444 (O_444,N_22140,N_24797);
and UO_445 (O_445,N_24216,N_24342);
xnor UO_446 (O_446,N_23180,N_23396);
nor UO_447 (O_447,N_23441,N_21989);
xnor UO_448 (O_448,N_22201,N_22829);
and UO_449 (O_449,N_24913,N_22699);
nand UO_450 (O_450,N_23202,N_24438);
and UO_451 (O_451,N_23268,N_22608);
nor UO_452 (O_452,N_24688,N_24765);
or UO_453 (O_453,N_24413,N_22873);
nand UO_454 (O_454,N_24855,N_21953);
nor UO_455 (O_455,N_22048,N_22019);
nor UO_456 (O_456,N_23155,N_24807);
and UO_457 (O_457,N_22253,N_22685);
xnor UO_458 (O_458,N_23278,N_24140);
nor UO_459 (O_459,N_22641,N_21887);
xnor UO_460 (O_460,N_23173,N_23214);
nand UO_461 (O_461,N_22357,N_22702);
nor UO_462 (O_462,N_24853,N_23910);
nand UO_463 (O_463,N_23487,N_23675);
and UO_464 (O_464,N_23118,N_24841);
xnor UO_465 (O_465,N_24049,N_24167);
nor UO_466 (O_466,N_23451,N_23638);
and UO_467 (O_467,N_24508,N_23905);
and UO_468 (O_468,N_22594,N_22339);
nand UO_469 (O_469,N_24997,N_24272);
nand UO_470 (O_470,N_21875,N_22661);
xnor UO_471 (O_471,N_24450,N_22757);
or UO_472 (O_472,N_22628,N_22738);
nand UO_473 (O_473,N_23481,N_22462);
nor UO_474 (O_474,N_23226,N_23346);
xnor UO_475 (O_475,N_22610,N_24665);
nor UO_476 (O_476,N_22006,N_23808);
and UO_477 (O_477,N_23863,N_24099);
xnor UO_478 (O_478,N_24078,N_22338);
nand UO_479 (O_479,N_24771,N_24902);
nand UO_480 (O_480,N_23131,N_24215);
nor UO_481 (O_481,N_23609,N_22228);
or UO_482 (O_482,N_24088,N_22573);
xor UO_483 (O_483,N_23387,N_24386);
and UO_484 (O_484,N_22978,N_24471);
or UO_485 (O_485,N_22592,N_24305);
and UO_486 (O_486,N_24502,N_22317);
and UO_487 (O_487,N_22479,N_23043);
or UO_488 (O_488,N_24963,N_24323);
and UO_489 (O_489,N_22663,N_24984);
or UO_490 (O_490,N_24046,N_22778);
nor UO_491 (O_491,N_24929,N_22965);
and UO_492 (O_492,N_22148,N_22310);
xor UO_493 (O_493,N_24291,N_22122);
xor UO_494 (O_494,N_22729,N_22187);
xor UO_495 (O_495,N_24946,N_22994);
xor UO_496 (O_496,N_22834,N_24337);
or UO_497 (O_497,N_22588,N_22705);
and UO_498 (O_498,N_23498,N_24430);
nor UO_499 (O_499,N_23014,N_24033);
and UO_500 (O_500,N_23603,N_22893);
nor UO_501 (O_501,N_21995,N_24712);
nand UO_502 (O_502,N_24298,N_22891);
nor UO_503 (O_503,N_24916,N_22593);
and UO_504 (O_504,N_24117,N_22200);
nor UO_505 (O_505,N_24735,N_22966);
or UO_506 (O_506,N_22049,N_21963);
and UO_507 (O_507,N_23397,N_24059);
nor UO_508 (O_508,N_23509,N_23309);
and UO_509 (O_509,N_23615,N_24451);
nand UO_510 (O_510,N_23984,N_22433);
and UO_511 (O_511,N_22121,N_23521);
nor UO_512 (O_512,N_23892,N_24260);
and UO_513 (O_513,N_24029,N_22907);
xnor UO_514 (O_514,N_24533,N_22427);
nor UO_515 (O_515,N_24903,N_24838);
nand UO_516 (O_516,N_21945,N_23627);
nor UO_517 (O_517,N_22721,N_22075);
nand UO_518 (O_518,N_23524,N_23106);
or UO_519 (O_519,N_23228,N_23587);
and UO_520 (O_520,N_24868,N_24697);
and UO_521 (O_521,N_24922,N_22500);
nor UO_522 (O_522,N_24434,N_23188);
or UO_523 (O_523,N_24889,N_24919);
and UO_524 (O_524,N_24456,N_24785);
nor UO_525 (O_525,N_23788,N_21979);
nor UO_526 (O_526,N_23418,N_23085);
nor UO_527 (O_527,N_21899,N_23726);
and UO_528 (O_528,N_22418,N_24652);
or UO_529 (O_529,N_23584,N_22329);
nand UO_530 (O_530,N_24066,N_22589);
or UO_531 (O_531,N_24689,N_22186);
or UO_532 (O_532,N_23234,N_24271);
or UO_533 (O_533,N_24908,N_22814);
nor UO_534 (O_534,N_23690,N_22368);
xor UO_535 (O_535,N_23667,N_24203);
nand UO_536 (O_536,N_24023,N_24854);
and UO_537 (O_537,N_23356,N_22842);
or UO_538 (O_538,N_23708,N_23540);
or UO_539 (O_539,N_22167,N_21937);
nor UO_540 (O_540,N_24616,N_21949);
or UO_541 (O_541,N_24670,N_22232);
and UO_542 (O_542,N_22050,N_23502);
nor UO_543 (O_543,N_24111,N_22131);
and UO_544 (O_544,N_22153,N_22471);
or UO_545 (O_545,N_24823,N_23024);
nand UO_546 (O_546,N_22998,N_22126);
nand UO_547 (O_547,N_23594,N_23791);
nor UO_548 (O_548,N_23302,N_23232);
nor UO_549 (O_549,N_24992,N_24662);
or UO_550 (O_550,N_23535,N_22900);
nor UO_551 (O_551,N_23171,N_24976);
or UO_552 (O_552,N_24101,N_23887);
or UO_553 (O_553,N_24408,N_23148);
or UO_554 (O_554,N_24322,N_23854);
nor UO_555 (O_555,N_24335,N_23849);
or UO_556 (O_556,N_23168,N_22903);
xnor UO_557 (O_557,N_23585,N_23318);
and UO_558 (O_558,N_24995,N_23586);
nand UO_559 (O_559,N_23235,N_22717);
or UO_560 (O_560,N_24955,N_23297);
or UO_561 (O_561,N_24313,N_23542);
xor UO_562 (O_562,N_23862,N_24395);
and UO_563 (O_563,N_21981,N_24897);
and UO_564 (O_564,N_23575,N_21948);
nor UO_565 (O_565,N_23563,N_24368);
nand UO_566 (O_566,N_22342,N_22452);
nand UO_567 (O_567,N_24460,N_22621);
and UO_568 (O_568,N_23970,N_22806);
nand UO_569 (O_569,N_24936,N_22905);
nand UO_570 (O_570,N_22769,N_22975);
nand UO_571 (O_571,N_22263,N_22934);
or UO_572 (O_572,N_24091,N_23204);
nor UO_573 (O_573,N_24351,N_23331);
nand UO_574 (O_574,N_23086,N_24361);
and UO_575 (O_575,N_22369,N_23211);
and UO_576 (O_576,N_24671,N_22826);
or UO_577 (O_577,N_23030,N_22224);
and UO_578 (O_578,N_24486,N_21898);
nand UO_579 (O_579,N_24265,N_22401);
nand UO_580 (O_580,N_24557,N_23714);
nor UO_581 (O_581,N_22961,N_24164);
xnor UO_582 (O_582,N_22909,N_22603);
nor UO_583 (O_583,N_21912,N_24630);
or UO_584 (O_584,N_24938,N_22622);
or UO_585 (O_585,N_23814,N_22843);
nand UO_586 (O_586,N_24136,N_22941);
xnor UO_587 (O_587,N_24760,N_22615);
xnor UO_588 (O_588,N_24143,N_23980);
nand UO_589 (O_589,N_24355,N_24018);
nand UO_590 (O_590,N_22577,N_24530);
xnor UO_591 (O_591,N_24128,N_23007);
or UO_592 (O_592,N_23482,N_24165);
nand UO_593 (O_593,N_22911,N_22154);
nor UO_594 (O_594,N_24968,N_22043);
nand UO_595 (O_595,N_23434,N_22737);
or UO_596 (O_596,N_23853,N_24704);
nand UO_597 (O_597,N_22030,N_24132);
nor UO_598 (O_598,N_23756,N_24089);
nand UO_599 (O_599,N_22921,N_22125);
nor UO_600 (O_600,N_24990,N_22203);
xor UO_601 (O_601,N_24607,N_22015);
or UO_602 (O_602,N_24407,N_23288);
or UO_603 (O_603,N_22184,N_24274);
xor UO_604 (O_604,N_22102,N_22217);
and UO_605 (O_605,N_22135,N_23866);
nor UO_606 (O_606,N_22191,N_23748);
nor UO_607 (O_607,N_24789,N_23755);
nand UO_608 (O_608,N_22633,N_23817);
and UO_609 (O_609,N_23762,N_24171);
nand UO_610 (O_610,N_22997,N_21999);
nor UO_611 (O_611,N_22216,N_23693);
xor UO_612 (O_612,N_22235,N_24719);
or UO_613 (O_613,N_22612,N_23950);
nand UO_614 (O_614,N_22942,N_23189);
nand UO_615 (O_615,N_22068,N_23448);
nand UO_616 (O_616,N_23142,N_22257);
nor UO_617 (O_617,N_22215,N_23347);
nor UO_618 (O_618,N_24915,N_24694);
and UO_619 (O_619,N_23280,N_24324);
nor UO_620 (O_620,N_24794,N_24942);
nor UO_621 (O_621,N_24121,N_23199);
or UO_622 (O_622,N_23209,N_23084);
and UO_623 (O_623,N_22568,N_22845);
nand UO_624 (O_624,N_23839,N_23797);
or UO_625 (O_625,N_23263,N_23958);
nand UO_626 (O_626,N_22207,N_24718);
nand UO_627 (O_627,N_22062,N_24343);
or UO_628 (O_628,N_24394,N_21971);
or UO_629 (O_629,N_23399,N_22847);
xor UO_630 (O_630,N_23630,N_22024);
nor UO_631 (O_631,N_24243,N_22748);
nand UO_632 (O_632,N_23717,N_24254);
and UO_633 (O_633,N_24726,N_24141);
or UO_634 (O_634,N_24953,N_23452);
nor UO_635 (O_635,N_23419,N_23846);
nor UO_636 (O_636,N_22327,N_23374);
nand UO_637 (O_637,N_23696,N_23102);
nand UO_638 (O_638,N_23976,N_22753);
and UO_639 (O_639,N_22010,N_23423);
or UO_640 (O_640,N_24634,N_24962);
nor UO_641 (O_641,N_24030,N_22752);
nand UO_642 (O_642,N_22397,N_24597);
nor UO_643 (O_643,N_23354,N_22956);
and UO_644 (O_644,N_23377,N_23306);
or UO_645 (O_645,N_24488,N_23987);
nor UO_646 (O_646,N_24988,N_24185);
xor UO_647 (O_647,N_22970,N_24200);
or UO_648 (O_648,N_22578,N_24809);
xnor UO_649 (O_649,N_24599,N_22706);
nand UO_650 (O_650,N_23629,N_23601);
or UO_651 (O_651,N_24832,N_22450);
nand UO_652 (O_652,N_22619,N_22662);
and UO_653 (O_653,N_23927,N_24546);
nor UO_654 (O_654,N_23569,N_22498);
nor UO_655 (O_655,N_22157,N_21950);
nand UO_656 (O_656,N_24055,N_23539);
nand UO_657 (O_657,N_22715,N_24578);
nand UO_658 (O_658,N_22745,N_24595);
nand UO_659 (O_659,N_21933,N_23270);
nand UO_660 (O_660,N_24977,N_24552);
nor UO_661 (O_661,N_24400,N_22676);
and UO_662 (O_662,N_24934,N_22658);
or UO_663 (O_663,N_23847,N_24631);
nand UO_664 (O_664,N_23759,N_24427);
or UO_665 (O_665,N_22730,N_22776);
or UO_666 (O_666,N_23833,N_23046);
or UO_667 (O_667,N_22273,N_22764);
or UO_668 (O_668,N_24865,N_22309);
nand UO_669 (O_669,N_23129,N_23900);
nor UO_670 (O_670,N_22516,N_24551);
xor UO_671 (O_671,N_22686,N_24683);
and UO_672 (O_672,N_23350,N_23695);
or UO_673 (O_673,N_21911,N_24741);
xnor UO_674 (O_674,N_24082,N_24494);
or UO_675 (O_675,N_22012,N_24403);
or UO_676 (O_676,N_24212,N_22284);
nor UO_677 (O_677,N_24170,N_24126);
and UO_678 (O_678,N_23707,N_23703);
nor UO_679 (O_679,N_21883,N_24691);
nand UO_680 (O_680,N_22239,N_24690);
and UO_681 (O_681,N_23314,N_23650);
and UO_682 (O_682,N_23336,N_22733);
nand UO_683 (O_683,N_24233,N_24706);
or UO_684 (O_684,N_24969,N_24363);
xor UO_685 (O_685,N_22894,N_23153);
nand UO_686 (O_686,N_22777,N_23764);
nand UO_687 (O_687,N_24684,N_24820);
nor UO_688 (O_688,N_21992,N_23467);
nand UO_689 (O_689,N_24183,N_23308);
and UO_690 (O_690,N_23061,N_24981);
and UO_691 (O_691,N_22853,N_23655);
or UO_692 (O_692,N_23879,N_24926);
xor UO_693 (O_693,N_24296,N_22634);
nand UO_694 (O_694,N_22774,N_22819);
nand UO_695 (O_695,N_22206,N_23167);
or UO_696 (O_696,N_22028,N_24686);
nor UO_697 (O_697,N_23834,N_23867);
nand UO_698 (O_698,N_22935,N_24746);
and UO_699 (O_699,N_24947,N_24231);
and UO_700 (O_700,N_23772,N_24750);
nor UO_701 (O_701,N_23417,N_24986);
or UO_702 (O_702,N_24129,N_22766);
and UO_703 (O_703,N_24836,N_24531);
nand UO_704 (O_704,N_24974,N_23859);
and UO_705 (O_705,N_24221,N_22623);
and UO_706 (O_706,N_23365,N_21896);
nor UO_707 (O_707,N_22247,N_22097);
or UO_708 (O_708,N_22428,N_24751);
xor UO_709 (O_709,N_23903,N_23945);
nand UO_710 (O_710,N_24457,N_24933);
and UO_711 (O_711,N_24504,N_22503);
and UO_712 (O_712,N_22791,N_22548);
nor UO_713 (O_713,N_22635,N_23537);
nor UO_714 (O_714,N_23295,N_22398);
nand UO_715 (O_715,N_24257,N_23922);
nor UO_716 (O_716,N_22261,N_22959);
nor UO_717 (O_717,N_24086,N_22613);
xor UO_718 (O_718,N_24636,N_24319);
and UO_719 (O_719,N_22320,N_23951);
or UO_720 (O_720,N_23206,N_24905);
nand UO_721 (O_721,N_24782,N_22002);
nand UO_722 (O_722,N_22362,N_23463);
and UO_723 (O_723,N_21955,N_22539);
and UO_724 (O_724,N_23593,N_22822);
nand UO_725 (O_725,N_22351,N_23178);
or UO_726 (O_726,N_24236,N_23766);
nor UO_727 (O_727,N_22698,N_21990);
nor UO_728 (O_728,N_22115,N_23430);
and UO_729 (O_729,N_22701,N_24593);
or UO_730 (O_730,N_22446,N_23652);
nor UO_731 (O_731,N_23999,N_22926);
and UO_732 (O_732,N_24698,N_23729);
or UO_733 (O_733,N_23626,N_22497);
and UO_734 (O_734,N_23786,N_22486);
or UO_735 (O_735,N_22554,N_22160);
and UO_736 (O_736,N_24814,N_22485);
nor UO_737 (O_737,N_23919,N_23192);
and UO_738 (O_738,N_22408,N_24138);
and UO_739 (O_739,N_24869,N_23956);
and UO_740 (O_740,N_22673,N_21913);
nor UO_741 (O_741,N_23789,N_22304);
nor UO_742 (O_742,N_23027,N_24367);
nand UO_743 (O_743,N_24890,N_22756);
xnor UO_744 (O_744,N_24240,N_23267);
or UO_745 (O_745,N_22374,N_23567);
and UO_746 (O_746,N_24674,N_23721);
nor UO_747 (O_747,N_22556,N_24332);
and UO_748 (O_748,N_24985,N_22876);
or UO_749 (O_749,N_22727,N_22712);
and UO_750 (O_750,N_24882,N_23111);
nor UO_751 (O_751,N_22011,N_24238);
nand UO_752 (O_752,N_24357,N_22473);
xor UO_753 (O_753,N_22901,N_23898);
nor UO_754 (O_754,N_22155,N_23715);
and UO_755 (O_755,N_22274,N_23773);
and UO_756 (O_756,N_23016,N_22103);
nand UO_757 (O_757,N_23461,N_22205);
nand UO_758 (O_758,N_23913,N_23548);
or UO_759 (O_759,N_22071,N_23304);
and UO_760 (O_760,N_24672,N_22138);
or UO_761 (O_761,N_22250,N_22288);
xor UO_762 (O_762,N_24316,N_22156);
and UO_763 (O_763,N_24251,N_23921);
and UO_764 (O_764,N_24114,N_23294);
nand UO_765 (O_765,N_24605,N_24432);
nor UO_766 (O_766,N_22192,N_23634);
nor UO_767 (O_767,N_24064,N_23995);
xor UO_768 (O_768,N_22447,N_22797);
and UO_769 (O_769,N_23972,N_23439);
nor UO_770 (O_770,N_24341,N_23187);
nor UO_771 (O_771,N_23087,N_24640);
nor UO_772 (O_772,N_22278,N_24710);
and UO_773 (O_773,N_22695,N_22580);
nor UO_774 (O_774,N_22188,N_24858);
and UO_775 (O_775,N_23960,N_23144);
nor UO_776 (O_776,N_22459,N_24499);
nor UO_777 (O_777,N_24191,N_23881);
or UO_778 (O_778,N_23514,N_24766);
nor UO_779 (O_779,N_23281,N_24802);
and UO_780 (O_780,N_22171,N_23174);
or UO_781 (O_781,N_22352,N_24781);
nand UO_782 (O_782,N_24068,N_23362);
nor UO_783 (O_783,N_22540,N_22316);
or UO_784 (O_784,N_22579,N_23261);
and UO_785 (O_785,N_23138,N_22624);
nor UO_786 (O_786,N_24071,N_24478);
and UO_787 (O_787,N_22933,N_23570);
nor UO_788 (O_788,N_23078,N_22669);
nand UO_789 (O_789,N_24376,N_22882);
or UO_790 (O_790,N_24987,N_23855);
xor UO_791 (O_791,N_22237,N_24720);
and UO_792 (O_792,N_23679,N_22312);
and UO_793 (O_793,N_23276,N_24292);
nand UO_794 (O_794,N_22208,N_23317);
and UO_795 (O_795,N_23044,N_23371);
or UO_796 (O_796,N_22132,N_24294);
nor UO_797 (O_797,N_22938,N_22919);
nor UO_798 (O_798,N_23665,N_23719);
nor UO_799 (O_799,N_24105,N_22214);
and UO_800 (O_800,N_23606,N_22348);
and UO_801 (O_801,N_22581,N_22925);
nor UO_802 (O_802,N_22502,N_24736);
nand UO_803 (O_803,N_22431,N_23139);
or UO_804 (O_804,N_23182,N_22982);
nand UO_805 (O_805,N_22631,N_24130);
or UO_806 (O_806,N_24007,N_24571);
nor UO_807 (O_807,N_24654,N_23262);
nand UO_808 (O_808,N_22665,N_22044);
and UO_809 (O_809,N_23733,N_24692);
nand UO_810 (O_810,N_22036,N_23457);
nand UO_811 (O_811,N_24196,N_21910);
and UO_812 (O_812,N_24857,N_24758);
nand UO_813 (O_813,N_22801,N_24103);
nor UO_814 (O_814,N_23175,N_22957);
or UO_815 (O_815,N_22912,N_21890);
xnor UO_816 (O_816,N_22538,N_22870);
nand UO_817 (O_817,N_23042,N_23943);
or UO_818 (O_818,N_22831,N_23151);
nand UO_819 (O_819,N_23706,N_23728);
or UO_820 (O_820,N_23761,N_24625);
nand UO_821 (O_821,N_23954,N_24172);
nor UO_822 (O_822,N_23329,N_24025);
nor UO_823 (O_823,N_23549,N_24281);
or UO_824 (O_824,N_21909,N_22147);
nand UO_825 (O_825,N_22098,N_23004);
or UO_826 (O_826,N_22734,N_24909);
and UO_827 (O_827,N_23654,N_22001);
nor UO_828 (O_828,N_23826,N_23475);
and UO_829 (O_829,N_23012,N_23727);
nand UO_830 (O_830,N_23983,N_22323);
and UO_831 (O_831,N_22560,N_22675);
nor UO_832 (O_832,N_23933,N_24439);
xor UO_833 (O_833,N_22768,N_23038);
xor UO_834 (O_834,N_24524,N_22493);
xor UO_835 (O_835,N_23017,N_24768);
and UO_836 (O_836,N_24507,N_24104);
nor UO_837 (O_837,N_23942,N_22346);
and UO_838 (O_838,N_23928,N_22291);
and UO_839 (O_839,N_22105,N_23117);
or UO_840 (O_840,N_24653,N_22117);
nand UO_841 (O_841,N_23827,N_23190);
nand UO_842 (O_842,N_23237,N_23656);
nor UO_843 (O_843,N_22599,N_24123);
or UO_844 (O_844,N_22297,N_22697);
and UO_845 (O_845,N_23997,N_22805);
and UO_846 (O_846,N_23070,N_22469);
xor UO_847 (O_847,N_24793,N_24448);
nand UO_848 (O_848,N_24678,N_22112);
or UO_849 (O_849,N_24177,N_21929);
nand UO_850 (O_850,N_24282,N_24941);
and UO_851 (O_851,N_23798,N_22863);
or UO_852 (O_852,N_21902,N_23050);
and UO_853 (O_853,N_24346,N_22713);
nor UO_854 (O_854,N_22400,N_23334);
nor UO_855 (O_855,N_23426,N_22671);
and UO_856 (O_856,N_22328,N_22543);
nand UO_857 (O_857,N_22222,N_24572);
and UO_858 (O_858,N_22561,N_22946);
xor UO_859 (O_859,N_23747,N_22750);
xor UO_860 (O_860,N_22227,N_24881);
xor UO_861 (O_861,N_22161,N_24058);
nand UO_862 (O_862,N_24280,N_21983);
xor UO_863 (O_863,N_23100,N_24074);
nor UO_864 (O_864,N_24958,N_22922);
and UO_865 (O_865,N_24010,N_22963);
and UO_866 (O_866,N_22813,N_23681);
nand UO_867 (O_867,N_24885,N_23159);
xnor UO_868 (O_868,N_22299,N_23645);
or UO_869 (O_869,N_24484,N_24852);
nor UO_870 (O_870,N_24214,N_22773);
nand UO_871 (O_871,N_23233,N_22367);
xnor UO_872 (O_872,N_24382,N_21876);
nor UO_873 (O_873,N_24618,N_22584);
nand UO_874 (O_874,N_24182,N_22668);
or UO_875 (O_875,N_24904,N_24960);
and UO_876 (O_876,N_23402,N_22209);
or UO_877 (O_877,N_24036,N_23120);
nand UO_878 (O_878,N_24851,N_24910);
or UO_879 (O_879,N_23522,N_24385);
or UO_880 (O_880,N_23710,N_23840);
nand UO_881 (O_881,N_22430,N_21977);
nor UO_882 (O_882,N_24151,N_23080);
and UO_883 (O_883,N_24729,N_23156);
or UO_884 (O_884,N_24708,N_22322);
and UO_885 (O_885,N_22718,N_23583);
and UO_886 (O_886,N_22977,N_24421);
and UO_887 (O_887,N_24057,N_21958);
nor UO_888 (O_888,N_22468,N_24211);
and UO_889 (O_889,N_22724,N_23591);
nor UO_890 (O_890,N_22081,N_22897);
nor UO_891 (O_891,N_23408,N_23531);
nor UO_892 (O_892,N_22943,N_22746);
and UO_893 (O_893,N_23513,N_24431);
nor UO_894 (O_894,N_23429,N_24702);
and UO_895 (O_895,N_24388,N_23890);
xor UO_896 (O_896,N_24519,N_24701);
and UO_897 (O_897,N_24108,N_24285);
nand UO_898 (O_898,N_22219,N_23088);
nor UO_899 (O_899,N_21939,N_22354);
and UO_900 (O_900,N_24015,N_24498);
or UO_901 (O_901,N_24510,N_22871);
and UO_902 (O_902,N_22572,N_24075);
or UO_903 (O_903,N_24576,N_23460);
nand UO_904 (O_904,N_23195,N_22089);
nand UO_905 (O_905,N_23464,N_22241);
nand UO_906 (O_906,N_23335,N_22021);
and UO_907 (O_907,N_22300,N_22567);
and UO_908 (O_908,N_24999,N_23692);
xnor UO_909 (O_909,N_22047,N_22687);
nor UO_910 (O_910,N_21907,N_24525);
or UO_911 (O_911,N_22258,N_22307);
and UO_912 (O_912,N_22952,N_23054);
nand UO_913 (O_913,N_21993,N_24849);
and UO_914 (O_914,N_22093,N_22295);
nand UO_915 (O_915,N_22240,N_23198);
and UO_916 (O_916,N_24559,N_22372);
xnor UO_917 (O_917,N_23711,N_22714);
nand UO_918 (O_918,N_23659,N_24812);
nor UO_919 (O_919,N_22489,N_22659);
and UO_920 (O_920,N_24592,N_23062);
nand UO_921 (O_921,N_23901,N_23218);
nand UO_922 (O_922,N_23299,N_23830);
xnor UO_923 (O_923,N_24210,N_22915);
nand UO_924 (O_924,N_23312,N_22242);
nor UO_925 (O_925,N_22660,N_22795);
and UO_926 (O_926,N_24818,N_23132);
nor UO_927 (O_927,N_23005,N_22755);
nand UO_928 (O_928,N_22857,N_22465);
and UO_929 (O_929,N_23010,N_24657);
or UO_930 (O_930,N_22595,N_22968);
nor UO_931 (O_931,N_24626,N_24004);
nor UO_932 (O_932,N_24585,N_22086);
xor UO_933 (O_933,N_24783,N_22034);
nand UO_934 (O_934,N_21934,N_22386);
and UO_935 (O_935,N_22804,N_24131);
nor UO_936 (O_936,N_23282,N_24297);
or UO_937 (O_937,N_23185,N_23339);
or UO_938 (O_938,N_24957,N_23712);
or UO_939 (O_939,N_22390,N_22283);
and UO_940 (O_940,N_21959,N_22004);
xor UO_941 (O_941,N_22781,N_23778);
nor UO_942 (O_942,N_22528,N_24207);
and UO_943 (O_943,N_23896,N_23254);
nor UO_944 (O_944,N_23874,N_22751);
or UO_945 (O_945,N_23246,N_23875);
and UO_946 (O_946,N_23915,N_23465);
nor UO_947 (O_947,N_24308,N_24727);
or UO_948 (O_948,N_22851,N_22534);
xor UO_949 (O_949,N_23449,N_21976);
xor UO_950 (O_950,N_23796,N_24900);
nand UO_951 (O_951,N_22178,N_22405);
nor UO_952 (O_952,N_22987,N_24501);
nand UO_953 (O_953,N_22544,N_22875);
nor UO_954 (O_954,N_22027,N_24124);
or UO_955 (O_955,N_23941,N_23421);
nor UO_956 (O_956,N_24821,N_24020);
and UO_957 (O_957,N_23929,N_23488);
nor UO_958 (O_958,N_23723,N_24045);
nor UO_959 (O_959,N_23000,N_24898);
and UO_960 (O_960,N_24347,N_24300);
and UO_961 (O_961,N_22277,N_24304);
nand UO_962 (O_962,N_23617,N_22366);
nor UO_963 (O_963,N_23687,N_24397);
xor UO_964 (O_964,N_22531,N_22000);
and UO_965 (O_965,N_22058,N_22683);
nor UO_966 (O_966,N_24245,N_23166);
nor UO_967 (O_967,N_23794,N_22415);
and UO_968 (O_968,N_24540,N_24463);
or UO_969 (O_969,N_24464,N_23971);
or UO_970 (O_970,N_23065,N_23642);
nor UO_971 (O_971,N_23793,N_23554);
and UO_972 (O_972,N_24414,N_22360);
and UO_973 (O_973,N_22267,N_23407);
nor UO_974 (O_974,N_24813,N_24831);
xor UO_975 (O_975,N_23737,N_21954);
nand UO_976 (O_976,N_22837,N_24978);
nor UO_977 (O_977,N_24261,N_23122);
nand UO_978 (O_978,N_23880,N_22176);
nor UO_979 (O_979,N_24906,N_24888);
or UO_980 (O_980,N_22443,N_24069);
or UO_981 (O_981,N_23820,N_23628);
and UO_982 (O_982,N_23093,N_23097);
nand UO_983 (O_983,N_24786,N_24772);
and UO_984 (O_984,N_24967,N_24353);
nor UO_985 (O_985,N_24288,N_22269);
nand UO_986 (O_986,N_22618,N_22371);
nor UO_987 (O_987,N_22079,N_24725);
and UO_988 (O_988,N_24466,N_24048);
nor UO_989 (O_989,N_22976,N_24119);
xnor UO_990 (O_990,N_22375,N_22387);
nand UO_991 (O_991,N_23242,N_22076);
nand UO_992 (O_992,N_21919,N_22646);
nand UO_993 (O_993,N_23952,N_24189);
nor UO_994 (O_994,N_24675,N_24467);
xor UO_995 (O_995,N_22101,N_23909);
xor UO_996 (O_996,N_23730,N_23994);
or UO_997 (O_997,N_24148,N_24031);
or UO_998 (O_998,N_23804,N_24569);
nand UO_999 (O_999,N_22260,N_22630);
nor UO_1000 (O_1000,N_23057,N_23388);
or UO_1001 (O_1001,N_22220,N_22094);
nor UO_1002 (O_1002,N_23287,N_22739);
or UO_1003 (O_1003,N_22536,N_24994);
and UO_1004 (O_1004,N_22591,N_22800);
and UO_1005 (O_1005,N_23285,N_22332);
and UO_1006 (O_1006,N_24754,N_22123);
nor UO_1007 (O_1007,N_22018,N_24053);
or UO_1008 (O_1008,N_23850,N_22436);
nor UO_1009 (O_1009,N_24584,N_23136);
nand UO_1010 (O_1010,N_23440,N_23864);
or UO_1011 (O_1011,N_22150,N_23431);
or UO_1012 (O_1012,N_23224,N_23033);
and UO_1013 (O_1013,N_23486,N_21973);
and UO_1014 (O_1014,N_23045,N_21994);
nor UO_1015 (O_1015,N_22035,N_24951);
nor UO_1016 (O_1016,N_22828,N_24362);
nand UO_1017 (O_1017,N_22169,N_22530);
or UO_1018 (O_1018,N_24232,N_21882);
or UO_1019 (O_1019,N_22246,N_23674);
or UO_1020 (O_1020,N_23436,N_23669);
nand UO_1021 (O_1021,N_22265,N_23229);
nand UO_1022 (O_1022,N_24449,N_24144);
xor UO_1023 (O_1023,N_24632,N_23274);
xor UO_1024 (O_1024,N_24681,N_24756);
nor UO_1025 (O_1025,N_24237,N_22793);
and UO_1026 (O_1026,N_23028,N_24461);
and UO_1027 (O_1027,N_24567,N_24248);
nor UO_1028 (O_1028,N_23561,N_21891);
or UO_1029 (O_1029,N_23581,N_21928);
and UO_1030 (O_1030,N_22731,N_23990);
or UO_1031 (O_1031,N_24721,N_24639);
xor UO_1032 (O_1032,N_23803,N_23220);
and UO_1033 (O_1033,N_24184,N_22198);
or UO_1034 (O_1034,N_23957,N_22254);
or UO_1035 (O_1035,N_23073,N_22555);
nand UO_1036 (O_1036,N_23750,N_22786);
or UO_1037 (O_1037,N_23260,N_23098);
nand UO_1038 (O_1038,N_23018,N_24306);
or UO_1039 (O_1039,N_23366,N_23577);
and UO_1040 (O_1040,N_24392,N_22704);
and UO_1041 (O_1041,N_22679,N_23777);
nand UO_1042 (O_1042,N_22645,N_22614);
nor UO_1043 (O_1043,N_24769,N_23435);
nor UO_1044 (O_1044,N_23543,N_24880);
or UO_1045 (O_1045,N_23810,N_21987);
nor UO_1046 (O_1046,N_22051,N_23824);
nand UO_1047 (O_1047,N_23357,N_23946);
and UO_1048 (O_1048,N_22827,N_24090);
or UO_1049 (O_1049,N_24709,N_22754);
and UO_1050 (O_1050,N_22818,N_22337);
and UO_1051 (O_1051,N_22887,N_22629);
or UO_1052 (O_1052,N_24970,N_24035);
and UO_1053 (O_1053,N_23256,N_24453);
or UO_1054 (O_1054,N_23279,N_24495);
and UO_1055 (O_1055,N_22862,N_23265);
or UO_1056 (O_1056,N_24966,N_23829);
nand UO_1057 (O_1057,N_23082,N_24176);
or UO_1058 (O_1058,N_23103,N_23300);
and UO_1059 (O_1059,N_23731,N_24180);
and UO_1060 (O_1060,N_23624,N_23368);
xnor UO_1061 (O_1061,N_23272,N_24418);
nand UO_1062 (O_1062,N_24522,N_22529);
and UO_1063 (O_1063,N_22885,N_24160);
and UO_1064 (O_1064,N_22535,N_23807);
or UO_1065 (O_1065,N_22545,N_23792);
and UO_1066 (O_1066,N_23518,N_23790);
nor UO_1067 (O_1067,N_24005,N_22364);
or UO_1068 (O_1068,N_21917,N_23216);
nor UO_1069 (O_1069,N_23315,N_22130);
and UO_1070 (O_1070,N_23886,N_23653);
or UO_1071 (O_1071,N_22477,N_23194);
or UO_1072 (O_1072,N_22434,N_21965);
or UO_1073 (O_1073,N_24433,N_24621);
nand UO_1074 (O_1074,N_24622,N_22709);
nor UO_1075 (O_1075,N_23765,N_23768);
nand UO_1076 (O_1076,N_23355,N_23311);
or UO_1077 (O_1077,N_22949,N_22172);
nand UO_1078 (O_1078,N_24566,N_24269);
or UO_1079 (O_1079,N_24081,N_23286);
or UO_1080 (O_1080,N_22761,N_23238);
nand UO_1081 (O_1081,N_24874,N_24563);
nor UO_1082 (O_1082,N_23301,N_24127);
nand UO_1083 (O_1083,N_23619,N_24944);
and UO_1084 (O_1084,N_24384,N_24472);
or UO_1085 (O_1085,N_24424,N_22114);
nor UO_1086 (O_1086,N_23891,N_24120);
and UO_1087 (O_1087,N_24744,N_22510);
nor UO_1088 (O_1088,N_22319,N_22370);
nand UO_1089 (O_1089,N_23771,N_21985);
and UO_1090 (O_1090,N_22270,N_24699);
nand UO_1091 (O_1091,N_23325,N_21881);
nand UO_1092 (O_1092,N_24197,N_24980);
nor UO_1093 (O_1093,N_23512,N_24157);
nand UO_1094 (O_1094,N_23734,N_23108);
nor UO_1095 (O_1095,N_23845,N_23751);
or UO_1096 (O_1096,N_24041,N_24544);
nand UO_1097 (O_1097,N_23783,N_22559);
nand UO_1098 (O_1098,N_24983,N_24581);
and UO_1099 (O_1099,N_22947,N_23872);
nand UO_1100 (O_1100,N_24235,N_21980);
and UO_1101 (O_1101,N_23450,N_24310);
and UO_1102 (O_1102,N_21975,N_22999);
or UO_1103 (O_1103,N_23213,N_23544);
and UO_1104 (O_1104,N_24954,N_24550);
nand UO_1105 (O_1105,N_21997,N_22334);
and UO_1106 (O_1106,N_22844,N_24925);
nand UO_1107 (O_1107,N_22190,N_23427);
nor UO_1108 (O_1108,N_24700,N_24410);
nor UO_1109 (O_1109,N_24173,N_22950);
or UO_1110 (O_1110,N_22470,N_22557);
nand UO_1111 (O_1111,N_23428,N_22667);
nor UO_1112 (O_1112,N_21918,N_22506);
nor UO_1113 (O_1113,N_23925,N_24256);
or UO_1114 (O_1114,N_24762,N_23749);
nand UO_1115 (O_1115,N_24541,N_24072);
and UO_1116 (O_1116,N_24624,N_24156);
and UO_1117 (O_1117,N_23107,N_24181);
nor UO_1118 (O_1118,N_22971,N_22716);
or UO_1119 (O_1119,N_21892,N_23828);
nand UO_1120 (O_1120,N_24134,N_24975);
nand UO_1121 (O_1121,N_24002,N_24100);
nand UO_1122 (O_1122,N_24425,N_24646);
xnor UO_1123 (O_1123,N_24959,N_24458);
or UO_1124 (O_1124,N_22417,N_24429);
nand UO_1125 (O_1125,N_23332,N_24475);
xor UO_1126 (O_1126,N_24748,N_22149);
nand UO_1127 (O_1127,N_23483,N_24375);
or UO_1128 (O_1128,N_24749,N_23932);
nand UO_1129 (O_1129,N_24521,N_24255);
and UO_1130 (O_1130,N_24895,N_23343);
and UO_1131 (O_1131,N_23291,N_23602);
xnor UO_1132 (O_1132,N_23966,N_24656);
nand UO_1133 (O_1133,N_24876,N_22272);
and UO_1134 (O_1134,N_23075,N_23395);
and UO_1135 (O_1135,N_23742,N_22888);
nor UO_1136 (O_1136,N_24067,N_24443);
xnor UO_1137 (O_1137,N_24588,N_23916);
nand UO_1138 (O_1138,N_24259,N_23344);
nor UO_1139 (O_1139,N_23089,N_23559);
xnor UO_1140 (O_1140,N_22426,N_24808);
and UO_1141 (O_1141,N_24573,N_24826);
and UO_1142 (O_1142,N_22259,N_23472);
or UO_1143 (O_1143,N_24226,N_24411);
xor UO_1144 (O_1144,N_22656,N_24645);
xnor UO_1145 (O_1145,N_24759,N_23579);
and UO_1146 (O_1146,N_24225,N_23552);
nor UO_1147 (O_1147,N_22276,N_23660);
nor UO_1148 (O_1148,N_22230,N_23049);
or UO_1149 (O_1149,N_24358,N_24873);
nor UO_1150 (O_1150,N_24422,N_23101);
and UO_1151 (O_1151,N_23897,N_22137);
nor UO_1152 (O_1152,N_22481,N_24011);
and UO_1153 (O_1153,N_24527,N_22238);
or UO_1154 (O_1154,N_24948,N_24301);
or UO_1155 (O_1155,N_22229,N_21900);
or UO_1156 (O_1156,N_23641,N_24628);
and UO_1157 (O_1157,N_24441,N_23432);
nand UO_1158 (O_1158,N_21947,N_24893);
nand UO_1159 (O_1159,N_23453,N_23520);
or UO_1160 (O_1160,N_22906,N_23193);
and UO_1161 (O_1161,N_23197,N_22404);
xnor UO_1162 (O_1162,N_23212,N_23637);
or UO_1163 (O_1163,N_24452,N_22627);
xor UO_1164 (O_1164,N_22165,N_24825);
nor UO_1165 (O_1165,N_23064,N_23752);
nor UO_1166 (O_1166,N_22973,N_23401);
nand UO_1167 (O_1167,N_23149,N_23381);
or UO_1168 (O_1168,N_23002,N_22708);
xor UO_1169 (O_1169,N_23858,N_23613);
nor UO_1170 (O_1170,N_24609,N_22600);
nand UO_1171 (O_1171,N_22677,N_24318);
or UO_1172 (O_1172,N_23293,N_22420);
or UO_1173 (O_1173,N_21936,N_22582);
or UO_1174 (O_1174,N_23878,N_22039);
and UO_1175 (O_1175,N_21932,N_24515);
xor UO_1176 (O_1176,N_22562,N_22521);
and UO_1177 (O_1177,N_23383,N_24511);
or UO_1178 (O_1178,N_24034,N_22563);
and UO_1179 (O_1179,N_23963,N_23183);
nand UO_1180 (O_1180,N_24642,N_22736);
nor UO_1181 (O_1181,N_22293,N_23351);
or UO_1182 (O_1182,N_23640,N_22243);
and UO_1183 (O_1183,N_22392,N_22124);
and UO_1184 (O_1184,N_24901,N_23697);
or UO_1185 (O_1185,N_24390,N_24512);
nand UO_1186 (O_1186,N_22537,N_23745);
nand UO_1187 (O_1187,N_23702,N_23967);
and UO_1188 (O_1188,N_22654,N_22045);
and UO_1189 (O_1189,N_23119,N_23048);
or UO_1190 (O_1190,N_22597,N_22788);
nor UO_1191 (O_1191,N_23341,N_21886);
nor UO_1192 (O_1192,N_23639,N_22799);
nor UO_1193 (O_1193,N_22453,N_24008);
nor UO_1194 (O_1194,N_22979,N_23125);
xnor UO_1195 (O_1195,N_22877,N_22490);
and UO_1196 (O_1196,N_23501,N_21923);
and UO_1197 (O_1197,N_23538,N_24013);
nand UO_1198 (O_1198,N_24399,N_24044);
nand UO_1199 (O_1199,N_24087,N_23009);
nand UO_1200 (O_1200,N_23076,N_23495);
or UO_1201 (O_1201,N_22458,N_24137);
xnor UO_1202 (O_1202,N_22484,N_22596);
xor UO_1203 (O_1203,N_23779,N_23068);
and UO_1204 (O_1204,N_24611,N_22518);
or UO_1205 (O_1205,N_24842,N_23394);
or UO_1206 (O_1206,N_24060,N_24277);
or UO_1207 (O_1207,N_22840,N_24991);
nor UO_1208 (O_1208,N_24667,N_22343);
nor UO_1209 (O_1209,N_23067,N_23724);
nand UO_1210 (O_1210,N_22279,N_23657);
nor UO_1211 (O_1211,N_22391,N_24863);
and UO_1212 (O_1212,N_22722,N_24266);
nand UO_1213 (O_1213,N_23390,N_23316);
xnor UO_1214 (O_1214,N_22483,N_24835);
or UO_1215 (O_1215,N_23255,N_23787);
nand UO_1216 (O_1216,N_23322,N_24561);
nand UO_1217 (O_1217,N_22625,N_24174);
nor UO_1218 (O_1218,N_22136,N_23982);
and UO_1219 (O_1219,N_24500,N_24166);
and UO_1220 (O_1220,N_23172,N_22379);
nor UO_1221 (O_1221,N_24666,N_24365);
and UO_1222 (O_1222,N_23701,N_23622);
or UO_1223 (O_1223,N_24491,N_23031);
nand UO_1224 (O_1224,N_24490,N_23008);
and UO_1225 (O_1225,N_24733,N_23503);
or UO_1226 (O_1226,N_23813,N_23252);
nor UO_1227 (O_1227,N_23215,N_24420);
or UO_1228 (O_1228,N_24273,N_24844);
nor UO_1229 (O_1229,N_23837,N_23600);
and UO_1230 (O_1230,N_23671,N_22031);
or UO_1231 (O_1231,N_22091,N_24861);
nor UO_1232 (O_1232,N_23455,N_23883);
and UO_1233 (O_1233,N_24412,N_24526);
nor UO_1234 (O_1234,N_22861,N_23376);
nand UO_1235 (O_1235,N_23511,N_22305);
nand UO_1236 (O_1236,N_24459,N_23560);
and UO_1237 (O_1237,N_22080,N_24194);
nor UO_1238 (O_1238,N_23480,N_24330);
or UO_1239 (O_1239,N_23550,N_23110);
and UO_1240 (O_1240,N_22839,N_24887);
nor UO_1241 (O_1241,N_24834,N_24436);
nor UO_1242 (O_1242,N_23607,N_23818);
nand UO_1243 (O_1243,N_24032,N_23504);
nand UO_1244 (O_1244,N_22832,N_24617);
xor UO_1245 (O_1245,N_22732,N_24610);
and UO_1246 (O_1246,N_22008,N_24473);
xor UO_1247 (O_1247,N_23385,N_22444);
nor UO_1248 (O_1248,N_23275,N_22411);
nor UO_1249 (O_1249,N_22617,N_23445);
nand UO_1250 (O_1250,N_23670,N_22218);
and UO_1251 (O_1251,N_23746,N_22072);
xnor UO_1252 (O_1252,N_22055,N_22296);
and UO_1253 (O_1253,N_22910,N_24896);
nand UO_1254 (O_1254,N_24884,N_23414);
or UO_1255 (O_1255,N_22889,N_23114);
and UO_1256 (O_1256,N_22474,N_22880);
or UO_1257 (O_1257,N_24309,N_24763);
nor UO_1258 (O_1258,N_23631,N_24262);
and UO_1259 (O_1259,N_24118,N_24155);
nor UO_1260 (O_1260,N_23532,N_24730);
and UO_1261 (O_1261,N_24477,N_24695);
or UO_1262 (O_1262,N_23676,N_22564);
or UO_1263 (O_1263,N_24284,N_24328);
xnor UO_1264 (O_1264,N_21901,N_24620);
nand UO_1265 (O_1265,N_23985,N_22655);
and UO_1266 (O_1266,N_22321,N_24299);
nand UO_1267 (O_1267,N_24487,N_22151);
and UO_1268 (O_1268,N_22664,N_22928);
nand UO_1269 (O_1269,N_24770,N_22878);
or UO_1270 (O_1270,N_24479,N_23039);
xor UO_1271 (O_1271,N_22650,N_22416);
nand UO_1272 (O_1272,N_22425,N_23949);
nor UO_1273 (O_1273,N_24419,N_24239);
or UO_1274 (O_1274,N_24923,N_23924);
xor UO_1275 (O_1275,N_22119,N_22723);
nor UO_1276 (O_1276,N_24629,N_23258);
and UO_1277 (O_1277,N_23923,N_22700);
nand UO_1278 (O_1278,N_24594,N_23135);
and UO_1279 (O_1279,N_23533,N_23037);
nand UO_1280 (O_1280,N_23446,N_24063);
or UO_1281 (O_1281,N_24493,N_24796);
nand UO_1282 (O_1282,N_23848,N_24334);
nand UO_1283 (O_1283,N_24270,N_24465);
and UO_1284 (O_1284,N_24850,N_23618);
and UO_1285 (O_1285,N_24676,N_22202);
or UO_1286 (O_1286,N_22740,N_23648);
or UO_1287 (O_1287,N_23664,N_24687);
nor UO_1288 (O_1288,N_23709,N_24470);
or UO_1289 (O_1289,N_22848,N_24199);
nand UO_1290 (O_1290,N_24575,N_23546);
or UO_1291 (O_1291,N_24800,N_24017);
and UO_1292 (O_1292,N_22266,N_22213);
xnor UO_1293 (O_1293,N_23236,N_23079);
nor UO_1294 (O_1294,N_23157,N_22413);
and UO_1295 (O_1295,N_22133,N_23425);
and UO_1296 (O_1296,N_24378,N_22262);
nor UO_1297 (O_1297,N_22382,N_23806);
nor UO_1298 (O_1298,N_23911,N_22326);
and UO_1299 (O_1299,N_23939,N_23001);
nor UO_1300 (O_1300,N_21988,N_22881);
and UO_1301 (O_1301,N_23338,N_23871);
and UO_1302 (O_1302,N_23036,N_23558);
xnor UO_1303 (O_1303,N_22014,N_24042);
or UO_1304 (O_1304,N_22821,N_22302);
nand UO_1305 (O_1305,N_22442,N_23888);
or UO_1306 (O_1306,N_22990,N_23485);
nor UO_1307 (O_1307,N_23074,N_22527);
and UO_1308 (O_1308,N_23795,N_23930);
xor UO_1309 (O_1309,N_22884,N_23536);
nor UO_1310 (O_1310,N_22083,N_22077);
nor UO_1311 (O_1311,N_22042,N_22424);
nor UO_1312 (O_1312,N_22290,N_24589);
nand UO_1313 (O_1313,N_23705,N_23179);
or UO_1314 (O_1314,N_23269,N_23838);
xnor UO_1315 (O_1315,N_24538,N_24623);
or UO_1316 (O_1316,N_23177,N_22461);
nand UO_1317 (O_1317,N_21972,N_24950);
and UO_1318 (O_1318,N_22940,N_24142);
xnor UO_1319 (O_1319,N_24664,N_23310);
or UO_1320 (O_1320,N_23090,N_24537);
nor UO_1321 (O_1321,N_24878,N_23743);
nor UO_1322 (O_1322,N_24489,N_24065);
and UO_1323 (O_1323,N_23527,N_22197);
or UO_1324 (O_1324,N_23223,N_23510);
xnor UO_1325 (O_1325,N_24154,N_24389);
xor UO_1326 (O_1326,N_24287,N_22033);
or UO_1327 (O_1327,N_23926,N_24480);
xor UO_1328 (O_1328,N_24107,N_23506);
and UO_1329 (O_1329,N_22784,N_23121);
or UO_1330 (O_1330,N_22944,N_24084);
nand UO_1331 (O_1331,N_22547,N_23899);
nand UO_1332 (O_1332,N_23364,N_22478);
and UO_1333 (O_1333,N_22410,N_24275);
xor UO_1334 (O_1334,N_23517,N_22303);
nor UO_1335 (O_1335,N_24734,N_22023);
nor UO_1336 (O_1336,N_23499,N_22522);
nor UO_1337 (O_1337,N_22422,N_24435);
and UO_1338 (O_1338,N_23479,N_23150);
and UO_1339 (O_1339,N_22482,N_23398);
nand UO_1340 (O_1340,N_23565,N_22735);
nor UO_1341 (O_1341,N_23821,N_22248);
or UO_1342 (O_1342,N_22725,N_24406);
xnor UO_1343 (O_1343,N_22923,N_24682);
and UO_1344 (O_1344,N_23865,N_22523);
and UO_1345 (O_1345,N_22496,N_23116);
and UO_1346 (O_1346,N_23424,N_22798);
nor UO_1347 (O_1347,N_23353,N_23677);
or UO_1348 (O_1348,N_24979,N_23201);
nor UO_1349 (O_1349,N_23556,N_24647);
or UO_1350 (O_1350,N_23230,N_23474);
nor UO_1351 (O_1351,N_21880,N_24650);
and UO_1352 (O_1352,N_23572,N_24218);
xor UO_1353 (O_1353,N_24949,N_24213);
nor UO_1354 (O_1354,N_23025,N_23825);
nor UO_1355 (O_1355,N_24780,N_23760);
nand UO_1356 (O_1356,N_21895,N_23406);
or UO_1357 (O_1357,N_24651,N_23947);
xnor UO_1358 (O_1358,N_22349,N_22566);
and UO_1359 (O_1359,N_24092,N_22174);
nand UO_1360 (O_1360,N_24188,N_24325);
nand UO_1361 (O_1361,N_23819,N_23938);
or UO_1362 (O_1362,N_22583,N_23799);
xor UO_1363 (O_1363,N_22359,N_22575);
nor UO_1364 (O_1364,N_24338,N_24523);
xor UO_1365 (O_1365,N_24774,N_24583);
nand UO_1366 (O_1366,N_24696,N_24864);
nand UO_1367 (O_1367,N_23551,N_22407);
or UO_1368 (O_1368,N_22541,N_24249);
nand UO_1369 (O_1369,N_22134,N_22107);
and UO_1370 (O_1370,N_22325,N_21962);
and UO_1371 (O_1371,N_24714,N_22558);
nor UO_1372 (O_1372,N_24314,N_23458);
and UO_1373 (O_1373,N_23489,N_23437);
or UO_1374 (O_1374,N_24169,N_22100);
or UO_1375 (O_1375,N_23912,N_24326);
nor UO_1376 (O_1376,N_24076,N_22856);
or UO_1377 (O_1377,N_23736,N_24505);
or UO_1378 (O_1378,N_22118,N_24056);
and UO_1379 (O_1379,N_22289,N_23877);
nor UO_1380 (O_1380,N_23576,N_21982);
xor UO_1381 (O_1381,N_22747,N_21984);
nand UO_1382 (O_1382,N_23392,N_22439);
nor UO_1383 (O_1383,N_24321,N_22457);
nand UO_1384 (O_1384,N_22830,N_23140);
nor UO_1385 (O_1385,N_23071,N_23154);
nand UO_1386 (O_1386,N_23596,N_24787);
and UO_1387 (O_1387,N_23170,N_24370);
nor UO_1388 (O_1388,N_24928,N_24206);
nand UO_1389 (O_1389,N_23099,N_23146);
nor UO_1390 (O_1390,N_22212,N_24827);
and UO_1391 (O_1391,N_21908,N_22744);
or UO_1392 (O_1392,N_22916,N_22181);
nand UO_1393 (O_1393,N_23500,N_23937);
and UO_1394 (O_1394,N_22520,N_24828);
nand UO_1395 (O_1395,N_22495,N_24801);
or UO_1396 (O_1396,N_22022,N_22389);
nor UO_1397 (O_1397,N_23740,N_22883);
nor UO_1398 (O_1398,N_23595,N_23389);
nor UO_1399 (O_1399,N_23722,N_23283);
and UO_1400 (O_1400,N_24125,N_22437);
and UO_1401 (O_1401,N_23894,N_23191);
nor UO_1402 (O_1402,N_22681,N_23989);
or UO_1403 (O_1403,N_22895,N_22969);
nand UO_1404 (O_1404,N_23476,N_22480);
nand UO_1405 (O_1405,N_22866,N_22807);
and UO_1406 (O_1406,N_23259,N_24152);
and UO_1407 (O_1407,N_23831,N_24600);
or UO_1408 (O_1408,N_21922,N_22670);
and UO_1409 (O_1409,N_23986,N_21944);
or UO_1410 (O_1410,N_22762,N_22690);
and UO_1411 (O_1411,N_24286,N_24147);
nor UO_1412 (O_1412,N_24267,N_24485);
and UO_1413 (O_1413,N_21943,N_23782);
or UO_1414 (O_1414,N_22515,N_23680);
nand UO_1415 (O_1415,N_23273,N_23096);
or UO_1416 (O_1416,N_23092,N_24587);
nand UO_1417 (O_1417,N_24562,N_23507);
nand UO_1418 (O_1418,N_24964,N_22152);
nor UO_1419 (O_1419,N_22958,N_23815);
nor UO_1420 (O_1420,N_23857,N_22298);
xor UO_1421 (O_1421,N_22454,N_23608);
nand UO_1422 (O_1422,N_22330,N_22551);
and UO_1423 (O_1423,N_23732,N_23592);
nand UO_1424 (O_1424,N_23658,N_22092);
nand UO_1425 (O_1425,N_24570,N_24247);
nor UO_1426 (O_1426,N_22464,N_23473);
xnor UO_1427 (O_1427,N_23969,N_22268);
xnor UO_1428 (O_1428,N_23519,N_23271);
nor UO_1429 (O_1429,N_24146,N_22985);
and UO_1430 (O_1430,N_22409,N_23404);
nand UO_1431 (O_1431,N_24677,N_23668);
nor UO_1432 (O_1432,N_23320,N_22741);
nor UO_1433 (O_1433,N_24327,N_24577);
nand UO_1434 (O_1434,N_22501,N_22810);
and UO_1435 (O_1435,N_22145,N_24244);
nor UO_1436 (O_1436,N_23015,N_23134);
xor UO_1437 (O_1437,N_22824,N_23646);
nor UO_1438 (O_1438,N_23112,N_22236);
or UO_1439 (O_1439,N_23811,N_21996);
nor UO_1440 (O_1440,N_21904,N_22760);
and UO_1441 (O_1441,N_22353,N_23205);
or UO_1442 (O_1442,N_21946,N_22703);
or UO_1443 (O_1443,N_22377,N_23321);
nand UO_1444 (O_1444,N_24728,N_24924);
nor UO_1445 (O_1445,N_23802,N_23422);
or UO_1446 (O_1446,N_24019,N_23678);
and UO_1447 (O_1447,N_23244,N_22505);
and UO_1448 (O_1448,N_23885,N_22514);
nor UO_1449 (O_1449,N_24333,N_22109);
nand UO_1450 (O_1450,N_24602,N_21941);
and UO_1451 (O_1451,N_23459,N_22835);
nand UO_1452 (O_1452,N_24545,N_24529);
nand UO_1453 (O_1453,N_24345,N_23893);
or UO_1454 (O_1454,N_24026,N_24810);
nand UO_1455 (O_1455,N_22340,N_23720);
nand UO_1456 (O_1456,N_22383,N_22143);
nor UO_1457 (O_1457,N_23529,N_24204);
xnor UO_1458 (O_1458,N_22526,N_22313);
nor UO_1459 (O_1459,N_21893,N_22195);
or UO_1460 (O_1460,N_21906,N_24912);
and UO_1461 (O_1461,N_24918,N_24703);
and UO_1462 (O_1462,N_22113,N_23683);
nor UO_1463 (O_1463,N_22647,N_22972);
nor UO_1464 (O_1464,N_21935,N_24965);
nand UO_1465 (O_1465,N_22865,N_24175);
nand UO_1466 (O_1466,N_24564,N_22508);
or UO_1467 (O_1467,N_23053,N_24145);
xor UO_1468 (O_1468,N_24219,N_24582);
nor UO_1469 (O_1469,N_23738,N_22694);
and UO_1470 (O_1470,N_22350,N_23348);
or UO_1471 (O_1471,N_23965,N_22927);
nand UO_1472 (O_1472,N_24534,N_22939);
or UO_1473 (O_1473,N_24359,N_24097);
nand UO_1474 (O_1474,N_22640,N_22396);
nand UO_1475 (O_1475,N_24601,N_24417);
and UO_1476 (O_1476,N_23644,N_22096);
and UO_1477 (O_1477,N_24383,N_24866);
and UO_1478 (O_1478,N_24405,N_21970);
or UO_1479 (O_1479,N_23944,N_23469);
and UO_1480 (O_1480,N_22142,N_22166);
nand UO_1481 (O_1481,N_24635,N_22183);
or UO_1482 (O_1482,N_22720,N_24535);
nand UO_1483 (O_1483,N_22932,N_23109);
xnor UO_1484 (O_1484,N_22355,N_22082);
xor UO_1485 (O_1485,N_23744,N_24135);
xnor UO_1486 (O_1486,N_22691,N_24542);
nand UO_1487 (O_1487,N_23324,N_24649);
nand UO_1488 (O_1488,N_24230,N_24192);
or UO_1489 (O_1489,N_22867,N_23991);
nor UO_1490 (O_1490,N_22684,N_22779);
and UO_1491 (O_1491,N_23264,N_23115);
and UO_1492 (O_1492,N_23169,N_23292);
nand UO_1493 (O_1493,N_24806,N_22525);
or UO_1494 (O_1494,N_22333,N_24454);
nand UO_1495 (O_1495,N_23165,N_23384);
and UO_1496 (O_1496,N_22604,N_22772);
nor UO_1497 (O_1497,N_22158,N_22185);
or UO_1498 (O_1498,N_23290,N_23319);
nand UO_1499 (O_1499,N_22040,N_24819);
or UO_1500 (O_1500,N_23998,N_21951);
and UO_1501 (O_1501,N_22953,N_23605);
or UO_1502 (O_1502,N_24252,N_22519);
and UO_1503 (O_1503,N_22710,N_24883);
or UO_1504 (O_1504,N_24568,N_23651);
nand UO_1505 (O_1505,N_24778,N_24222);
and UO_1506 (O_1506,N_23066,N_22825);
or UO_1507 (O_1507,N_23217,N_24659);
nor UO_1508 (O_1508,N_22467,N_22294);
or UO_1509 (O_1509,N_23029,N_22211);
xnor UO_1510 (O_1510,N_23962,N_24892);
and UO_1511 (O_1511,N_23497,N_23022);
nor UO_1512 (O_1512,N_24776,N_24496);
nand UO_1513 (O_1513,N_21986,N_23176);
or UO_1514 (O_1514,N_24543,N_23443);
nand UO_1515 (O_1515,N_22549,N_23069);
and UO_1516 (O_1516,N_22384,N_24153);
nand UO_1517 (O_1517,N_23284,N_24416);
nor UO_1518 (O_1518,N_22005,N_24779);
or UO_1519 (O_1519,N_23420,N_23032);
nor UO_1520 (O_1520,N_23611,N_23635);
nand UO_1521 (O_1521,N_21925,N_22864);
and UO_1522 (O_1522,N_23094,N_23133);
nor UO_1523 (O_1523,N_21894,N_24711);
nand UO_1524 (O_1524,N_23367,N_23403);
or UO_1525 (O_1525,N_22929,N_22281);
or UO_1526 (O_1526,N_23158,N_24283);
xnor UO_1527 (O_1527,N_22429,N_24685);
nor UO_1528 (O_1528,N_24201,N_24845);
nor UO_1529 (O_1529,N_24931,N_22792);
nor UO_1530 (O_1530,N_22423,N_23598);
nor UO_1531 (O_1531,N_24830,N_22494);
xnor UO_1532 (O_1532,N_24603,N_22803);
nand UO_1533 (O_1533,N_22331,N_24016);
nor UO_1534 (O_1534,N_24000,N_22476);
or UO_1535 (O_1535,N_24083,N_22249);
nand UO_1536 (O_1536,N_23688,N_22904);
nand UO_1537 (O_1537,N_22849,N_22672);
and UO_1538 (O_1538,N_23816,N_21978);
and UO_1539 (O_1539,N_23409,N_22173);
nor UO_1540 (O_1540,N_23196,N_22026);
nand UO_1541 (O_1541,N_23589,N_24693);
xor UO_1542 (O_1542,N_23515,N_22226);
or UO_1543 (O_1543,N_23757,N_22951);
or UO_1544 (O_1544,N_23955,N_24737);
and UO_1545 (O_1545,N_23208,N_22974);
and UO_1546 (O_1546,N_24877,N_24409);
or UO_1547 (O_1547,N_24373,N_22692);
and UO_1548 (O_1548,N_24553,N_22569);
nor UO_1549 (O_1549,N_21888,N_23961);
nor UO_1550 (O_1550,N_23091,N_22585);
or UO_1551 (O_1551,N_23305,N_22204);
nand UO_1552 (O_1552,N_23493,N_23470);
nor UO_1553 (O_1553,N_24043,N_21877);
and UO_1554 (O_1554,N_22896,N_22170);
nor UO_1555 (O_1555,N_22168,N_22141);
nand UO_1556 (O_1556,N_24840,N_24276);
or UO_1557 (O_1557,N_23868,N_23968);
nor UO_1558 (O_1558,N_22902,N_23277);
nand UO_1559 (O_1559,N_24608,N_24110);
xor UO_1560 (O_1560,N_23250,N_21920);
nor UO_1561 (O_1561,N_23021,N_24354);
or UO_1562 (O_1562,N_22402,N_22768);
xor UO_1563 (O_1563,N_22139,N_22602);
nand UO_1564 (O_1564,N_23964,N_24005);
or UO_1565 (O_1565,N_23615,N_23511);
nand UO_1566 (O_1566,N_22367,N_22632);
nor UO_1567 (O_1567,N_23326,N_24260);
nand UO_1568 (O_1568,N_23663,N_23827);
nor UO_1569 (O_1569,N_22017,N_22905);
nand UO_1570 (O_1570,N_22839,N_24839);
nor UO_1571 (O_1571,N_22182,N_22432);
nand UO_1572 (O_1572,N_24181,N_24492);
xor UO_1573 (O_1573,N_23529,N_24456);
nand UO_1574 (O_1574,N_24094,N_22396);
nand UO_1575 (O_1575,N_23258,N_22285);
nand UO_1576 (O_1576,N_24211,N_23895);
nand UO_1577 (O_1577,N_23405,N_24724);
or UO_1578 (O_1578,N_23910,N_23524);
or UO_1579 (O_1579,N_22784,N_24192);
and UO_1580 (O_1580,N_24112,N_24030);
nor UO_1581 (O_1581,N_21968,N_24989);
and UO_1582 (O_1582,N_22461,N_22416);
nand UO_1583 (O_1583,N_22199,N_23642);
xnor UO_1584 (O_1584,N_23535,N_24594);
and UO_1585 (O_1585,N_23688,N_22148);
nor UO_1586 (O_1586,N_23301,N_22651);
or UO_1587 (O_1587,N_22601,N_23645);
and UO_1588 (O_1588,N_22328,N_23350);
and UO_1589 (O_1589,N_24640,N_22008);
and UO_1590 (O_1590,N_24060,N_22380);
or UO_1591 (O_1591,N_21984,N_22148);
nor UO_1592 (O_1592,N_23460,N_22594);
and UO_1593 (O_1593,N_23390,N_23965);
or UO_1594 (O_1594,N_24691,N_22749);
nor UO_1595 (O_1595,N_24588,N_23974);
nor UO_1596 (O_1596,N_22708,N_23060);
nand UO_1597 (O_1597,N_23620,N_24916);
nor UO_1598 (O_1598,N_24696,N_23406);
nand UO_1599 (O_1599,N_23069,N_24211);
or UO_1600 (O_1600,N_22885,N_22316);
nor UO_1601 (O_1601,N_23301,N_24185);
and UO_1602 (O_1602,N_22734,N_24189);
xor UO_1603 (O_1603,N_23898,N_23751);
and UO_1604 (O_1604,N_24525,N_24149);
and UO_1605 (O_1605,N_22638,N_22320);
or UO_1606 (O_1606,N_22806,N_24726);
nand UO_1607 (O_1607,N_22734,N_24757);
and UO_1608 (O_1608,N_23300,N_21898);
or UO_1609 (O_1609,N_22141,N_23989);
or UO_1610 (O_1610,N_23771,N_23009);
and UO_1611 (O_1611,N_24149,N_24279);
or UO_1612 (O_1612,N_23876,N_23086);
or UO_1613 (O_1613,N_24974,N_23635);
nand UO_1614 (O_1614,N_22510,N_24274);
or UO_1615 (O_1615,N_23333,N_24332);
or UO_1616 (O_1616,N_24080,N_24698);
or UO_1617 (O_1617,N_22870,N_24547);
xnor UO_1618 (O_1618,N_22869,N_21965);
nand UO_1619 (O_1619,N_22225,N_23602);
or UO_1620 (O_1620,N_24516,N_24473);
nor UO_1621 (O_1621,N_23941,N_23225);
and UO_1622 (O_1622,N_22003,N_22678);
nand UO_1623 (O_1623,N_23242,N_22381);
nor UO_1624 (O_1624,N_24342,N_22837);
or UO_1625 (O_1625,N_22726,N_22683);
and UO_1626 (O_1626,N_22657,N_23002);
and UO_1627 (O_1627,N_23101,N_23805);
and UO_1628 (O_1628,N_22731,N_21963);
and UO_1629 (O_1629,N_21896,N_23231);
xnor UO_1630 (O_1630,N_22699,N_22737);
nand UO_1631 (O_1631,N_22453,N_23575);
or UO_1632 (O_1632,N_21997,N_24792);
nor UO_1633 (O_1633,N_22778,N_21980);
and UO_1634 (O_1634,N_24211,N_23070);
or UO_1635 (O_1635,N_23688,N_23260);
nor UO_1636 (O_1636,N_23038,N_23414);
xor UO_1637 (O_1637,N_23196,N_22294);
nand UO_1638 (O_1638,N_22252,N_24253);
nand UO_1639 (O_1639,N_23177,N_24902);
or UO_1640 (O_1640,N_22309,N_21981);
nand UO_1641 (O_1641,N_22510,N_24457);
nor UO_1642 (O_1642,N_23200,N_23300);
nand UO_1643 (O_1643,N_22839,N_24008);
and UO_1644 (O_1644,N_23081,N_23413);
or UO_1645 (O_1645,N_24618,N_22472);
nor UO_1646 (O_1646,N_22707,N_22557);
nor UO_1647 (O_1647,N_22130,N_22193);
nand UO_1648 (O_1648,N_23298,N_23919);
xnor UO_1649 (O_1649,N_23138,N_24353);
nand UO_1650 (O_1650,N_24404,N_24019);
nor UO_1651 (O_1651,N_24010,N_23430);
or UO_1652 (O_1652,N_22391,N_22306);
nand UO_1653 (O_1653,N_24743,N_22235);
and UO_1654 (O_1654,N_24392,N_23074);
and UO_1655 (O_1655,N_24577,N_23306);
nand UO_1656 (O_1656,N_24525,N_23654);
or UO_1657 (O_1657,N_23187,N_23006);
or UO_1658 (O_1658,N_22600,N_23480);
nand UO_1659 (O_1659,N_24109,N_23482);
and UO_1660 (O_1660,N_23982,N_24385);
xnor UO_1661 (O_1661,N_23268,N_24940);
xor UO_1662 (O_1662,N_24466,N_23310);
nand UO_1663 (O_1663,N_22175,N_23360);
nor UO_1664 (O_1664,N_23822,N_24041);
nor UO_1665 (O_1665,N_24778,N_24867);
and UO_1666 (O_1666,N_22318,N_23849);
nor UO_1667 (O_1667,N_23254,N_22825);
nand UO_1668 (O_1668,N_23278,N_23261);
nand UO_1669 (O_1669,N_22866,N_24208);
or UO_1670 (O_1670,N_23444,N_22279);
nand UO_1671 (O_1671,N_21944,N_22234);
or UO_1672 (O_1672,N_23785,N_21946);
nor UO_1673 (O_1673,N_23723,N_23584);
nand UO_1674 (O_1674,N_23979,N_24937);
and UO_1675 (O_1675,N_22691,N_22295);
nand UO_1676 (O_1676,N_24066,N_23998);
nor UO_1677 (O_1677,N_23307,N_22683);
and UO_1678 (O_1678,N_23074,N_23660);
xor UO_1679 (O_1679,N_22816,N_22185);
or UO_1680 (O_1680,N_22546,N_22743);
nand UO_1681 (O_1681,N_24823,N_23037);
or UO_1682 (O_1682,N_23456,N_23425);
nand UO_1683 (O_1683,N_21964,N_23109);
and UO_1684 (O_1684,N_23166,N_24050);
nand UO_1685 (O_1685,N_23229,N_24874);
nor UO_1686 (O_1686,N_21979,N_22555);
nand UO_1687 (O_1687,N_24319,N_23693);
nor UO_1688 (O_1688,N_22615,N_24407);
nor UO_1689 (O_1689,N_22596,N_22258);
nor UO_1690 (O_1690,N_22774,N_22862);
or UO_1691 (O_1691,N_22996,N_22099);
nand UO_1692 (O_1692,N_22305,N_24314);
and UO_1693 (O_1693,N_24409,N_22844);
nand UO_1694 (O_1694,N_23927,N_22112);
nor UO_1695 (O_1695,N_24012,N_23708);
nand UO_1696 (O_1696,N_23466,N_22017);
nand UO_1697 (O_1697,N_22532,N_24776);
nand UO_1698 (O_1698,N_23301,N_24498);
xor UO_1699 (O_1699,N_22478,N_24374);
nor UO_1700 (O_1700,N_24202,N_24870);
xor UO_1701 (O_1701,N_21964,N_22302);
and UO_1702 (O_1702,N_22102,N_23251);
or UO_1703 (O_1703,N_24456,N_23358);
or UO_1704 (O_1704,N_21906,N_22713);
and UO_1705 (O_1705,N_22520,N_22447);
or UO_1706 (O_1706,N_22075,N_24556);
and UO_1707 (O_1707,N_23108,N_23229);
nor UO_1708 (O_1708,N_24097,N_23182);
and UO_1709 (O_1709,N_22681,N_23466);
nand UO_1710 (O_1710,N_23964,N_23283);
nand UO_1711 (O_1711,N_24966,N_22835);
nor UO_1712 (O_1712,N_23955,N_21909);
and UO_1713 (O_1713,N_24651,N_23496);
nand UO_1714 (O_1714,N_23113,N_23156);
or UO_1715 (O_1715,N_24631,N_21981);
or UO_1716 (O_1716,N_24784,N_23395);
and UO_1717 (O_1717,N_23245,N_23746);
or UO_1718 (O_1718,N_24023,N_24923);
and UO_1719 (O_1719,N_22600,N_24442);
xnor UO_1720 (O_1720,N_24055,N_22774);
nor UO_1721 (O_1721,N_22203,N_24457);
or UO_1722 (O_1722,N_21920,N_22502);
xnor UO_1723 (O_1723,N_23953,N_23122);
nand UO_1724 (O_1724,N_23966,N_23715);
nor UO_1725 (O_1725,N_23058,N_22445);
nor UO_1726 (O_1726,N_24311,N_22543);
and UO_1727 (O_1727,N_23561,N_22180);
xnor UO_1728 (O_1728,N_24498,N_22242);
nand UO_1729 (O_1729,N_21877,N_23244);
nor UO_1730 (O_1730,N_22670,N_22681);
nor UO_1731 (O_1731,N_22999,N_24502);
nor UO_1732 (O_1732,N_22522,N_24957);
nor UO_1733 (O_1733,N_24302,N_23885);
or UO_1734 (O_1734,N_24302,N_23506);
and UO_1735 (O_1735,N_22235,N_23256);
or UO_1736 (O_1736,N_24632,N_24485);
and UO_1737 (O_1737,N_22904,N_21902);
nor UO_1738 (O_1738,N_21929,N_24631);
nor UO_1739 (O_1739,N_22005,N_24197);
or UO_1740 (O_1740,N_23239,N_24117);
or UO_1741 (O_1741,N_24599,N_22125);
and UO_1742 (O_1742,N_22049,N_24115);
or UO_1743 (O_1743,N_22934,N_21959);
and UO_1744 (O_1744,N_24697,N_22347);
nand UO_1745 (O_1745,N_23766,N_24702);
nor UO_1746 (O_1746,N_24930,N_22041);
xor UO_1747 (O_1747,N_22146,N_22635);
nand UO_1748 (O_1748,N_21931,N_22878);
nor UO_1749 (O_1749,N_23254,N_24693);
and UO_1750 (O_1750,N_21990,N_24309);
nand UO_1751 (O_1751,N_22389,N_22767);
or UO_1752 (O_1752,N_23242,N_23479);
nor UO_1753 (O_1753,N_24387,N_23186);
nand UO_1754 (O_1754,N_24290,N_23437);
nand UO_1755 (O_1755,N_23047,N_23191);
and UO_1756 (O_1756,N_23639,N_23456);
or UO_1757 (O_1757,N_23073,N_22890);
and UO_1758 (O_1758,N_23828,N_24495);
nand UO_1759 (O_1759,N_22896,N_23185);
or UO_1760 (O_1760,N_23879,N_24548);
nand UO_1761 (O_1761,N_22729,N_23741);
and UO_1762 (O_1762,N_22717,N_23909);
and UO_1763 (O_1763,N_24382,N_23654);
and UO_1764 (O_1764,N_22176,N_22523);
or UO_1765 (O_1765,N_23006,N_24008);
nor UO_1766 (O_1766,N_24752,N_24425);
nand UO_1767 (O_1767,N_23926,N_24307);
or UO_1768 (O_1768,N_24330,N_24127);
nor UO_1769 (O_1769,N_22299,N_23544);
and UO_1770 (O_1770,N_23848,N_24719);
or UO_1771 (O_1771,N_24329,N_23285);
xnor UO_1772 (O_1772,N_24109,N_22024);
xor UO_1773 (O_1773,N_24529,N_24533);
nor UO_1774 (O_1774,N_23754,N_24465);
or UO_1775 (O_1775,N_24840,N_24074);
nor UO_1776 (O_1776,N_23152,N_21889);
and UO_1777 (O_1777,N_22368,N_24413);
nand UO_1778 (O_1778,N_24737,N_23733);
and UO_1779 (O_1779,N_22768,N_23961);
nand UO_1780 (O_1780,N_23460,N_24863);
or UO_1781 (O_1781,N_22885,N_24413);
nor UO_1782 (O_1782,N_22158,N_23069);
nand UO_1783 (O_1783,N_22690,N_22720);
nor UO_1784 (O_1784,N_23686,N_23374);
and UO_1785 (O_1785,N_23833,N_24818);
and UO_1786 (O_1786,N_23713,N_24657);
nand UO_1787 (O_1787,N_24500,N_22073);
nand UO_1788 (O_1788,N_22458,N_22784);
and UO_1789 (O_1789,N_22063,N_22336);
and UO_1790 (O_1790,N_22979,N_24348);
and UO_1791 (O_1791,N_24352,N_23941);
and UO_1792 (O_1792,N_23724,N_22349);
xnor UO_1793 (O_1793,N_22044,N_22108);
xnor UO_1794 (O_1794,N_22854,N_22388);
nor UO_1795 (O_1795,N_23697,N_23548);
and UO_1796 (O_1796,N_23312,N_21941);
or UO_1797 (O_1797,N_23903,N_22220);
nand UO_1798 (O_1798,N_22984,N_22517);
nand UO_1799 (O_1799,N_24917,N_23443);
nand UO_1800 (O_1800,N_24554,N_22180);
nor UO_1801 (O_1801,N_23813,N_23623);
and UO_1802 (O_1802,N_24122,N_23772);
xnor UO_1803 (O_1803,N_22239,N_22895);
nor UO_1804 (O_1804,N_23989,N_23444);
or UO_1805 (O_1805,N_22457,N_23187);
nand UO_1806 (O_1806,N_23248,N_22955);
nand UO_1807 (O_1807,N_24261,N_22058);
nor UO_1808 (O_1808,N_22092,N_23403);
or UO_1809 (O_1809,N_22861,N_24117);
nor UO_1810 (O_1810,N_22117,N_24191);
and UO_1811 (O_1811,N_22168,N_24429);
xor UO_1812 (O_1812,N_24910,N_22528);
nor UO_1813 (O_1813,N_24380,N_23282);
nand UO_1814 (O_1814,N_23895,N_24833);
nand UO_1815 (O_1815,N_23317,N_23096);
and UO_1816 (O_1816,N_24225,N_22386);
nor UO_1817 (O_1817,N_23618,N_24702);
nor UO_1818 (O_1818,N_22479,N_22224);
and UO_1819 (O_1819,N_22144,N_24204);
nor UO_1820 (O_1820,N_23969,N_22088);
nand UO_1821 (O_1821,N_21988,N_24318);
or UO_1822 (O_1822,N_24710,N_22862);
or UO_1823 (O_1823,N_23777,N_23782);
nor UO_1824 (O_1824,N_22733,N_24060);
or UO_1825 (O_1825,N_21899,N_23572);
nand UO_1826 (O_1826,N_23543,N_22990);
and UO_1827 (O_1827,N_24629,N_22286);
or UO_1828 (O_1828,N_23439,N_24593);
and UO_1829 (O_1829,N_23144,N_22896);
xnor UO_1830 (O_1830,N_23479,N_22021);
xor UO_1831 (O_1831,N_24610,N_22834);
nor UO_1832 (O_1832,N_22935,N_22311);
or UO_1833 (O_1833,N_23343,N_24612);
nor UO_1834 (O_1834,N_23148,N_22374);
or UO_1835 (O_1835,N_21927,N_21920);
or UO_1836 (O_1836,N_23531,N_22526);
nor UO_1837 (O_1837,N_22627,N_22938);
or UO_1838 (O_1838,N_24745,N_23108);
or UO_1839 (O_1839,N_24690,N_23541);
or UO_1840 (O_1840,N_24674,N_21937);
nand UO_1841 (O_1841,N_23746,N_22520);
nor UO_1842 (O_1842,N_22777,N_22186);
nor UO_1843 (O_1843,N_22357,N_22230);
or UO_1844 (O_1844,N_23404,N_23076);
nor UO_1845 (O_1845,N_23588,N_24324);
and UO_1846 (O_1846,N_22993,N_23482);
or UO_1847 (O_1847,N_24207,N_24882);
xnor UO_1848 (O_1848,N_23851,N_24033);
nand UO_1849 (O_1849,N_22040,N_24313);
or UO_1850 (O_1850,N_22463,N_21991);
nand UO_1851 (O_1851,N_23254,N_23133);
nor UO_1852 (O_1852,N_22184,N_24722);
or UO_1853 (O_1853,N_22320,N_23821);
or UO_1854 (O_1854,N_23692,N_24762);
xor UO_1855 (O_1855,N_24640,N_21987);
or UO_1856 (O_1856,N_23482,N_23549);
and UO_1857 (O_1857,N_24462,N_22780);
or UO_1858 (O_1858,N_24515,N_22874);
nor UO_1859 (O_1859,N_23167,N_22260);
nor UO_1860 (O_1860,N_22132,N_23594);
nor UO_1861 (O_1861,N_22212,N_24158);
xnor UO_1862 (O_1862,N_24170,N_24728);
and UO_1863 (O_1863,N_23463,N_24416);
or UO_1864 (O_1864,N_22800,N_22157);
or UO_1865 (O_1865,N_22828,N_22871);
and UO_1866 (O_1866,N_22693,N_22470);
xnor UO_1867 (O_1867,N_23422,N_23606);
nand UO_1868 (O_1868,N_23156,N_22596);
and UO_1869 (O_1869,N_22872,N_24601);
nand UO_1870 (O_1870,N_23792,N_23088);
or UO_1871 (O_1871,N_22658,N_23337);
or UO_1872 (O_1872,N_23890,N_24528);
and UO_1873 (O_1873,N_24774,N_23168);
and UO_1874 (O_1874,N_22959,N_22540);
nand UO_1875 (O_1875,N_23426,N_24047);
xnor UO_1876 (O_1876,N_22896,N_24617);
or UO_1877 (O_1877,N_24830,N_24005);
xnor UO_1878 (O_1878,N_24311,N_22660);
nand UO_1879 (O_1879,N_24388,N_24457);
and UO_1880 (O_1880,N_23017,N_24542);
and UO_1881 (O_1881,N_22736,N_22966);
nand UO_1882 (O_1882,N_24689,N_22649);
or UO_1883 (O_1883,N_23180,N_23518);
and UO_1884 (O_1884,N_23617,N_22835);
or UO_1885 (O_1885,N_22764,N_24570);
nor UO_1886 (O_1886,N_23571,N_23549);
or UO_1887 (O_1887,N_22925,N_22381);
and UO_1888 (O_1888,N_22275,N_22956);
nor UO_1889 (O_1889,N_22675,N_24993);
xnor UO_1890 (O_1890,N_22726,N_24034);
nor UO_1891 (O_1891,N_23887,N_22601);
and UO_1892 (O_1892,N_24326,N_24092);
and UO_1893 (O_1893,N_22771,N_22427);
and UO_1894 (O_1894,N_24560,N_22614);
nand UO_1895 (O_1895,N_22110,N_24964);
or UO_1896 (O_1896,N_23524,N_23849);
nand UO_1897 (O_1897,N_24750,N_22049);
or UO_1898 (O_1898,N_22113,N_22986);
or UO_1899 (O_1899,N_24428,N_22923);
and UO_1900 (O_1900,N_22038,N_23368);
nand UO_1901 (O_1901,N_23044,N_23134);
nor UO_1902 (O_1902,N_22691,N_22905);
and UO_1903 (O_1903,N_22570,N_23566);
nand UO_1904 (O_1904,N_22978,N_22091);
nor UO_1905 (O_1905,N_24562,N_22700);
nand UO_1906 (O_1906,N_22215,N_23484);
nand UO_1907 (O_1907,N_24951,N_24352);
or UO_1908 (O_1908,N_23665,N_22864);
and UO_1909 (O_1909,N_23633,N_22864);
nand UO_1910 (O_1910,N_22867,N_23461);
nor UO_1911 (O_1911,N_22115,N_22466);
nand UO_1912 (O_1912,N_22532,N_23045);
and UO_1913 (O_1913,N_23541,N_24522);
or UO_1914 (O_1914,N_23403,N_23087);
nand UO_1915 (O_1915,N_22201,N_22503);
nor UO_1916 (O_1916,N_22393,N_23264);
nand UO_1917 (O_1917,N_22649,N_22493);
or UO_1918 (O_1918,N_23864,N_23969);
nand UO_1919 (O_1919,N_22543,N_23949);
xor UO_1920 (O_1920,N_23987,N_23110);
or UO_1921 (O_1921,N_24528,N_22011);
xor UO_1922 (O_1922,N_22549,N_24895);
nor UO_1923 (O_1923,N_23421,N_24595);
xnor UO_1924 (O_1924,N_24752,N_22874);
nand UO_1925 (O_1925,N_24122,N_23889);
or UO_1926 (O_1926,N_22717,N_21975);
or UO_1927 (O_1927,N_24730,N_23623);
nand UO_1928 (O_1928,N_24038,N_24640);
nand UO_1929 (O_1929,N_21953,N_22794);
and UO_1930 (O_1930,N_24295,N_23632);
nor UO_1931 (O_1931,N_23215,N_24214);
or UO_1932 (O_1932,N_22632,N_22019);
nor UO_1933 (O_1933,N_24317,N_23402);
nor UO_1934 (O_1934,N_23379,N_23084);
or UO_1935 (O_1935,N_24832,N_22140);
nand UO_1936 (O_1936,N_23657,N_24115);
nand UO_1937 (O_1937,N_24600,N_22494);
xnor UO_1938 (O_1938,N_22357,N_22551);
nand UO_1939 (O_1939,N_23138,N_22744);
nand UO_1940 (O_1940,N_22710,N_22373);
nor UO_1941 (O_1941,N_24435,N_22988);
and UO_1942 (O_1942,N_22166,N_23274);
nor UO_1943 (O_1943,N_24007,N_22112);
and UO_1944 (O_1944,N_22599,N_23980);
and UO_1945 (O_1945,N_22325,N_22895);
or UO_1946 (O_1946,N_24282,N_24952);
nand UO_1947 (O_1947,N_22209,N_24411);
xor UO_1948 (O_1948,N_23830,N_24221);
nand UO_1949 (O_1949,N_23426,N_23920);
nand UO_1950 (O_1950,N_23758,N_24689);
or UO_1951 (O_1951,N_22616,N_23427);
or UO_1952 (O_1952,N_24675,N_22281);
or UO_1953 (O_1953,N_22662,N_22890);
or UO_1954 (O_1954,N_23324,N_23273);
nand UO_1955 (O_1955,N_23648,N_24087);
nor UO_1956 (O_1956,N_22864,N_22185);
nand UO_1957 (O_1957,N_24054,N_23347);
nand UO_1958 (O_1958,N_24291,N_22821);
nand UO_1959 (O_1959,N_22620,N_24630);
and UO_1960 (O_1960,N_23404,N_24651);
nor UO_1961 (O_1961,N_23181,N_23492);
xor UO_1962 (O_1962,N_22876,N_23889);
and UO_1963 (O_1963,N_23932,N_22830);
and UO_1964 (O_1964,N_23913,N_22763);
and UO_1965 (O_1965,N_24644,N_22560);
nor UO_1966 (O_1966,N_22405,N_22961);
xor UO_1967 (O_1967,N_23127,N_23019);
or UO_1968 (O_1968,N_23207,N_22058);
and UO_1969 (O_1969,N_22575,N_24701);
nor UO_1970 (O_1970,N_24632,N_21935);
xor UO_1971 (O_1971,N_24565,N_22839);
and UO_1972 (O_1972,N_23092,N_23606);
and UO_1973 (O_1973,N_21964,N_21876);
and UO_1974 (O_1974,N_22865,N_24559);
nand UO_1975 (O_1975,N_24619,N_24485);
and UO_1976 (O_1976,N_23936,N_22738);
xnor UO_1977 (O_1977,N_23486,N_24424);
or UO_1978 (O_1978,N_22747,N_23499);
nand UO_1979 (O_1979,N_23914,N_22470);
or UO_1980 (O_1980,N_24999,N_24616);
nor UO_1981 (O_1981,N_21949,N_23995);
and UO_1982 (O_1982,N_24721,N_23173);
or UO_1983 (O_1983,N_24964,N_23527);
nand UO_1984 (O_1984,N_24998,N_24842);
and UO_1985 (O_1985,N_23846,N_24780);
or UO_1986 (O_1986,N_24416,N_23664);
nand UO_1987 (O_1987,N_22840,N_24786);
or UO_1988 (O_1988,N_22302,N_21977);
nor UO_1989 (O_1989,N_24441,N_24221);
or UO_1990 (O_1990,N_23142,N_23083);
or UO_1991 (O_1991,N_24813,N_24196);
nand UO_1992 (O_1992,N_22929,N_24996);
and UO_1993 (O_1993,N_23480,N_23668);
nor UO_1994 (O_1994,N_24610,N_24312);
nand UO_1995 (O_1995,N_22525,N_22705);
xnor UO_1996 (O_1996,N_23998,N_24041);
and UO_1997 (O_1997,N_22732,N_23591);
xnor UO_1998 (O_1998,N_23733,N_22155);
nor UO_1999 (O_1999,N_22261,N_23297);
nand UO_2000 (O_2000,N_22097,N_23476);
nand UO_2001 (O_2001,N_24852,N_24892);
nand UO_2002 (O_2002,N_23537,N_22730);
or UO_2003 (O_2003,N_23848,N_23890);
or UO_2004 (O_2004,N_23597,N_22215);
nand UO_2005 (O_2005,N_23869,N_24169);
and UO_2006 (O_2006,N_22003,N_23880);
nand UO_2007 (O_2007,N_24931,N_24082);
and UO_2008 (O_2008,N_24478,N_24417);
or UO_2009 (O_2009,N_22903,N_24751);
nor UO_2010 (O_2010,N_23295,N_24046);
or UO_2011 (O_2011,N_22071,N_24327);
nand UO_2012 (O_2012,N_24941,N_22575);
and UO_2013 (O_2013,N_22060,N_21877);
nor UO_2014 (O_2014,N_23525,N_24899);
nor UO_2015 (O_2015,N_22544,N_22096);
or UO_2016 (O_2016,N_24774,N_22312);
xnor UO_2017 (O_2017,N_21912,N_24898);
or UO_2018 (O_2018,N_24652,N_23904);
and UO_2019 (O_2019,N_22161,N_22873);
and UO_2020 (O_2020,N_23049,N_24773);
and UO_2021 (O_2021,N_22073,N_23768);
nand UO_2022 (O_2022,N_23824,N_23168);
nand UO_2023 (O_2023,N_24540,N_24071);
nor UO_2024 (O_2024,N_22247,N_23397);
nand UO_2025 (O_2025,N_22848,N_22776);
and UO_2026 (O_2026,N_23981,N_24582);
or UO_2027 (O_2027,N_24626,N_24427);
nand UO_2028 (O_2028,N_23518,N_21912);
nor UO_2029 (O_2029,N_22456,N_24156);
and UO_2030 (O_2030,N_24405,N_23959);
or UO_2031 (O_2031,N_23234,N_23470);
or UO_2032 (O_2032,N_22337,N_24552);
and UO_2033 (O_2033,N_22969,N_23178);
and UO_2034 (O_2034,N_22763,N_22362);
xor UO_2035 (O_2035,N_22379,N_24342);
nand UO_2036 (O_2036,N_23563,N_22776);
nand UO_2037 (O_2037,N_23509,N_22848);
xor UO_2038 (O_2038,N_24562,N_22537);
nand UO_2039 (O_2039,N_23441,N_22035);
nor UO_2040 (O_2040,N_23551,N_24116);
nor UO_2041 (O_2041,N_22452,N_23887);
or UO_2042 (O_2042,N_23570,N_24001);
xnor UO_2043 (O_2043,N_23637,N_23863);
nand UO_2044 (O_2044,N_23255,N_23221);
nand UO_2045 (O_2045,N_24171,N_24085);
nor UO_2046 (O_2046,N_23726,N_22731);
nor UO_2047 (O_2047,N_24928,N_22902);
nand UO_2048 (O_2048,N_24427,N_24663);
and UO_2049 (O_2049,N_24385,N_24820);
and UO_2050 (O_2050,N_22292,N_24029);
or UO_2051 (O_2051,N_24617,N_24921);
or UO_2052 (O_2052,N_23664,N_24901);
nor UO_2053 (O_2053,N_22994,N_23580);
xnor UO_2054 (O_2054,N_23800,N_22313);
nand UO_2055 (O_2055,N_24994,N_22841);
or UO_2056 (O_2056,N_23798,N_23423);
xnor UO_2057 (O_2057,N_22256,N_21997);
and UO_2058 (O_2058,N_21890,N_22057);
or UO_2059 (O_2059,N_24275,N_21904);
and UO_2060 (O_2060,N_22490,N_24346);
xnor UO_2061 (O_2061,N_24090,N_24896);
and UO_2062 (O_2062,N_23050,N_23227);
nand UO_2063 (O_2063,N_22409,N_23477);
and UO_2064 (O_2064,N_23805,N_23884);
or UO_2065 (O_2065,N_24828,N_24738);
nor UO_2066 (O_2066,N_24919,N_24195);
or UO_2067 (O_2067,N_23944,N_24094);
nor UO_2068 (O_2068,N_23424,N_24897);
xnor UO_2069 (O_2069,N_22447,N_23007);
nand UO_2070 (O_2070,N_22758,N_22941);
and UO_2071 (O_2071,N_22486,N_22346);
or UO_2072 (O_2072,N_24219,N_22262);
nor UO_2073 (O_2073,N_24710,N_22021);
and UO_2074 (O_2074,N_22765,N_23882);
and UO_2075 (O_2075,N_23501,N_22664);
nor UO_2076 (O_2076,N_24785,N_22447);
or UO_2077 (O_2077,N_23184,N_24237);
nor UO_2078 (O_2078,N_22514,N_24059);
and UO_2079 (O_2079,N_22923,N_24031);
nand UO_2080 (O_2080,N_23694,N_24506);
nor UO_2081 (O_2081,N_24819,N_22699);
nor UO_2082 (O_2082,N_24858,N_24458);
and UO_2083 (O_2083,N_22758,N_24577);
nand UO_2084 (O_2084,N_21979,N_22637);
or UO_2085 (O_2085,N_24076,N_22655);
nor UO_2086 (O_2086,N_24775,N_23520);
nand UO_2087 (O_2087,N_22772,N_22454);
nor UO_2088 (O_2088,N_23537,N_24509);
and UO_2089 (O_2089,N_23419,N_24873);
and UO_2090 (O_2090,N_24216,N_22817);
nand UO_2091 (O_2091,N_22682,N_22882);
and UO_2092 (O_2092,N_24165,N_23730);
nor UO_2093 (O_2093,N_22393,N_23956);
or UO_2094 (O_2094,N_22070,N_24648);
and UO_2095 (O_2095,N_24963,N_23618);
nor UO_2096 (O_2096,N_24579,N_23953);
nand UO_2097 (O_2097,N_21883,N_23751);
and UO_2098 (O_2098,N_22543,N_24357);
nand UO_2099 (O_2099,N_24046,N_22437);
nand UO_2100 (O_2100,N_23279,N_21990);
xor UO_2101 (O_2101,N_24813,N_22841);
xor UO_2102 (O_2102,N_21881,N_22982);
and UO_2103 (O_2103,N_23997,N_24872);
or UO_2104 (O_2104,N_22736,N_24654);
or UO_2105 (O_2105,N_24851,N_22977);
nor UO_2106 (O_2106,N_22469,N_24577);
nand UO_2107 (O_2107,N_23162,N_22108);
nand UO_2108 (O_2108,N_22921,N_23058);
nor UO_2109 (O_2109,N_22229,N_23907);
nor UO_2110 (O_2110,N_23400,N_22966);
or UO_2111 (O_2111,N_24828,N_22586);
nor UO_2112 (O_2112,N_24105,N_24510);
or UO_2113 (O_2113,N_23677,N_22455);
or UO_2114 (O_2114,N_22077,N_22391);
nor UO_2115 (O_2115,N_22439,N_24337);
and UO_2116 (O_2116,N_22092,N_23278);
and UO_2117 (O_2117,N_22150,N_24493);
or UO_2118 (O_2118,N_24516,N_22808);
nand UO_2119 (O_2119,N_23220,N_22788);
and UO_2120 (O_2120,N_22757,N_24908);
or UO_2121 (O_2121,N_24943,N_23424);
or UO_2122 (O_2122,N_24609,N_23521);
nand UO_2123 (O_2123,N_24195,N_23253);
or UO_2124 (O_2124,N_22776,N_23873);
and UO_2125 (O_2125,N_21937,N_22767);
or UO_2126 (O_2126,N_24099,N_23995);
or UO_2127 (O_2127,N_23978,N_22792);
nor UO_2128 (O_2128,N_22590,N_21998);
or UO_2129 (O_2129,N_22043,N_24909);
nand UO_2130 (O_2130,N_22861,N_23735);
or UO_2131 (O_2131,N_23359,N_21938);
nor UO_2132 (O_2132,N_24698,N_22458);
nand UO_2133 (O_2133,N_24068,N_24250);
and UO_2134 (O_2134,N_23469,N_22388);
or UO_2135 (O_2135,N_22186,N_23585);
or UO_2136 (O_2136,N_23185,N_23277);
nand UO_2137 (O_2137,N_24170,N_23328);
and UO_2138 (O_2138,N_24279,N_23654);
and UO_2139 (O_2139,N_24317,N_24213);
nor UO_2140 (O_2140,N_22579,N_24516);
or UO_2141 (O_2141,N_22872,N_23417);
nand UO_2142 (O_2142,N_23096,N_23140);
nand UO_2143 (O_2143,N_22046,N_22490);
nand UO_2144 (O_2144,N_21916,N_24768);
xnor UO_2145 (O_2145,N_22514,N_22093);
nor UO_2146 (O_2146,N_22605,N_24080);
nand UO_2147 (O_2147,N_24126,N_24188);
nand UO_2148 (O_2148,N_22812,N_22062);
nor UO_2149 (O_2149,N_22588,N_22249);
nor UO_2150 (O_2150,N_22631,N_24936);
or UO_2151 (O_2151,N_24639,N_22487);
nand UO_2152 (O_2152,N_22942,N_23577);
or UO_2153 (O_2153,N_22322,N_23950);
xnor UO_2154 (O_2154,N_22660,N_24831);
nand UO_2155 (O_2155,N_22222,N_22309);
nor UO_2156 (O_2156,N_23449,N_24781);
nand UO_2157 (O_2157,N_22759,N_24582);
or UO_2158 (O_2158,N_22127,N_23289);
nor UO_2159 (O_2159,N_22011,N_22529);
xnor UO_2160 (O_2160,N_23595,N_23728);
or UO_2161 (O_2161,N_22069,N_23731);
xnor UO_2162 (O_2162,N_22451,N_24355);
and UO_2163 (O_2163,N_22652,N_22143);
nand UO_2164 (O_2164,N_23932,N_22658);
and UO_2165 (O_2165,N_23950,N_23113);
and UO_2166 (O_2166,N_22208,N_24710);
and UO_2167 (O_2167,N_24301,N_22721);
nor UO_2168 (O_2168,N_22258,N_23705);
nor UO_2169 (O_2169,N_24878,N_23755);
and UO_2170 (O_2170,N_22153,N_24459);
nor UO_2171 (O_2171,N_24540,N_23702);
nand UO_2172 (O_2172,N_22554,N_24444);
nor UO_2173 (O_2173,N_23047,N_24349);
and UO_2174 (O_2174,N_24919,N_24375);
xor UO_2175 (O_2175,N_22851,N_24111);
and UO_2176 (O_2176,N_24624,N_23606);
nor UO_2177 (O_2177,N_24899,N_24495);
nor UO_2178 (O_2178,N_24380,N_22724);
or UO_2179 (O_2179,N_24136,N_23406);
xor UO_2180 (O_2180,N_23850,N_23723);
or UO_2181 (O_2181,N_23755,N_23124);
nor UO_2182 (O_2182,N_24086,N_24682);
or UO_2183 (O_2183,N_23077,N_22434);
and UO_2184 (O_2184,N_22914,N_24025);
or UO_2185 (O_2185,N_23797,N_22162);
or UO_2186 (O_2186,N_24386,N_24309);
nand UO_2187 (O_2187,N_24670,N_23883);
nand UO_2188 (O_2188,N_22864,N_23484);
and UO_2189 (O_2189,N_22088,N_22290);
nor UO_2190 (O_2190,N_24574,N_22182);
and UO_2191 (O_2191,N_23462,N_24416);
nor UO_2192 (O_2192,N_21970,N_23630);
or UO_2193 (O_2193,N_24561,N_23265);
xor UO_2194 (O_2194,N_24796,N_23945);
and UO_2195 (O_2195,N_24043,N_24620);
xnor UO_2196 (O_2196,N_22533,N_23841);
and UO_2197 (O_2197,N_23445,N_23274);
and UO_2198 (O_2198,N_23892,N_24133);
and UO_2199 (O_2199,N_22454,N_24920);
nor UO_2200 (O_2200,N_22012,N_21936);
nand UO_2201 (O_2201,N_23927,N_24813);
and UO_2202 (O_2202,N_23536,N_24303);
nand UO_2203 (O_2203,N_23295,N_23755);
nand UO_2204 (O_2204,N_22625,N_21978);
or UO_2205 (O_2205,N_24714,N_23837);
or UO_2206 (O_2206,N_24801,N_23200);
nor UO_2207 (O_2207,N_22873,N_24626);
xor UO_2208 (O_2208,N_24690,N_23331);
and UO_2209 (O_2209,N_23369,N_24852);
nor UO_2210 (O_2210,N_24312,N_24630);
or UO_2211 (O_2211,N_24690,N_24870);
or UO_2212 (O_2212,N_24577,N_22627);
and UO_2213 (O_2213,N_23017,N_22664);
and UO_2214 (O_2214,N_23892,N_22140);
xnor UO_2215 (O_2215,N_24575,N_22369);
and UO_2216 (O_2216,N_23958,N_22931);
nor UO_2217 (O_2217,N_23986,N_22960);
nor UO_2218 (O_2218,N_24451,N_23963);
and UO_2219 (O_2219,N_23606,N_23911);
nand UO_2220 (O_2220,N_22367,N_23954);
nand UO_2221 (O_2221,N_23425,N_24701);
nor UO_2222 (O_2222,N_24859,N_24971);
xor UO_2223 (O_2223,N_24859,N_23003);
xnor UO_2224 (O_2224,N_24970,N_24108);
nor UO_2225 (O_2225,N_24178,N_23590);
nand UO_2226 (O_2226,N_24160,N_22821);
nand UO_2227 (O_2227,N_22366,N_24453);
nor UO_2228 (O_2228,N_24057,N_23126);
nor UO_2229 (O_2229,N_24932,N_24021);
xor UO_2230 (O_2230,N_23525,N_23435);
and UO_2231 (O_2231,N_24837,N_23936);
or UO_2232 (O_2232,N_23645,N_23288);
or UO_2233 (O_2233,N_24454,N_23697);
nor UO_2234 (O_2234,N_22181,N_24318);
xor UO_2235 (O_2235,N_22696,N_24707);
or UO_2236 (O_2236,N_23756,N_23628);
or UO_2237 (O_2237,N_24727,N_23379);
xnor UO_2238 (O_2238,N_22458,N_23879);
and UO_2239 (O_2239,N_23737,N_24784);
or UO_2240 (O_2240,N_22995,N_24491);
and UO_2241 (O_2241,N_24841,N_23783);
nand UO_2242 (O_2242,N_22130,N_24335);
or UO_2243 (O_2243,N_23904,N_24435);
nand UO_2244 (O_2244,N_24842,N_24526);
or UO_2245 (O_2245,N_23847,N_23701);
and UO_2246 (O_2246,N_24460,N_23766);
nor UO_2247 (O_2247,N_22072,N_23306);
nor UO_2248 (O_2248,N_21972,N_24270);
and UO_2249 (O_2249,N_24237,N_22943);
xnor UO_2250 (O_2250,N_23290,N_24916);
or UO_2251 (O_2251,N_24521,N_24858);
or UO_2252 (O_2252,N_24746,N_22037);
nor UO_2253 (O_2253,N_21979,N_23965);
and UO_2254 (O_2254,N_22119,N_23307);
nor UO_2255 (O_2255,N_23856,N_24906);
nand UO_2256 (O_2256,N_22112,N_22835);
and UO_2257 (O_2257,N_24647,N_22496);
nand UO_2258 (O_2258,N_23089,N_24827);
nor UO_2259 (O_2259,N_22995,N_24974);
nor UO_2260 (O_2260,N_23197,N_23267);
xor UO_2261 (O_2261,N_21984,N_23436);
nor UO_2262 (O_2262,N_23560,N_23787);
xor UO_2263 (O_2263,N_23028,N_22947);
nand UO_2264 (O_2264,N_24013,N_23497);
nor UO_2265 (O_2265,N_22490,N_22613);
or UO_2266 (O_2266,N_24924,N_22797);
and UO_2267 (O_2267,N_24639,N_23380);
or UO_2268 (O_2268,N_22396,N_23734);
and UO_2269 (O_2269,N_24958,N_23171);
and UO_2270 (O_2270,N_21928,N_23440);
nand UO_2271 (O_2271,N_23011,N_23642);
nand UO_2272 (O_2272,N_22075,N_22126);
and UO_2273 (O_2273,N_22647,N_23664);
nand UO_2274 (O_2274,N_23274,N_23810);
and UO_2275 (O_2275,N_22767,N_22055);
nand UO_2276 (O_2276,N_23298,N_24899);
or UO_2277 (O_2277,N_22197,N_23610);
or UO_2278 (O_2278,N_23510,N_23626);
xnor UO_2279 (O_2279,N_22085,N_23320);
and UO_2280 (O_2280,N_22682,N_22474);
or UO_2281 (O_2281,N_24237,N_22869);
or UO_2282 (O_2282,N_24215,N_24046);
or UO_2283 (O_2283,N_23823,N_24278);
and UO_2284 (O_2284,N_22417,N_23356);
or UO_2285 (O_2285,N_23738,N_22937);
nand UO_2286 (O_2286,N_23156,N_23345);
or UO_2287 (O_2287,N_23349,N_24750);
nor UO_2288 (O_2288,N_22627,N_24741);
nand UO_2289 (O_2289,N_24852,N_23896);
nand UO_2290 (O_2290,N_23336,N_22146);
or UO_2291 (O_2291,N_23419,N_23826);
nor UO_2292 (O_2292,N_23220,N_24211);
nand UO_2293 (O_2293,N_24715,N_22359);
nand UO_2294 (O_2294,N_22025,N_22087);
xor UO_2295 (O_2295,N_23071,N_23928);
or UO_2296 (O_2296,N_24995,N_22856);
and UO_2297 (O_2297,N_23608,N_24366);
nor UO_2298 (O_2298,N_22833,N_22631);
nand UO_2299 (O_2299,N_22992,N_22975);
nor UO_2300 (O_2300,N_24153,N_21960);
nand UO_2301 (O_2301,N_23571,N_24570);
or UO_2302 (O_2302,N_23040,N_24887);
xnor UO_2303 (O_2303,N_24108,N_24781);
or UO_2304 (O_2304,N_23424,N_23918);
nand UO_2305 (O_2305,N_24541,N_22846);
xor UO_2306 (O_2306,N_23645,N_22772);
or UO_2307 (O_2307,N_24204,N_24361);
nand UO_2308 (O_2308,N_22792,N_22597);
or UO_2309 (O_2309,N_22817,N_24028);
nand UO_2310 (O_2310,N_22263,N_23970);
and UO_2311 (O_2311,N_24637,N_24039);
or UO_2312 (O_2312,N_23010,N_22400);
xnor UO_2313 (O_2313,N_24464,N_23012);
nand UO_2314 (O_2314,N_22258,N_23442);
or UO_2315 (O_2315,N_23801,N_24280);
xor UO_2316 (O_2316,N_22522,N_22451);
or UO_2317 (O_2317,N_23062,N_22743);
or UO_2318 (O_2318,N_24557,N_23861);
nand UO_2319 (O_2319,N_22258,N_22115);
nand UO_2320 (O_2320,N_22940,N_23040);
and UO_2321 (O_2321,N_24711,N_23265);
xor UO_2322 (O_2322,N_23996,N_23081);
nand UO_2323 (O_2323,N_22606,N_24599);
and UO_2324 (O_2324,N_24965,N_23910);
nand UO_2325 (O_2325,N_23777,N_23254);
or UO_2326 (O_2326,N_24951,N_24882);
nand UO_2327 (O_2327,N_24372,N_24485);
nor UO_2328 (O_2328,N_23156,N_22242);
and UO_2329 (O_2329,N_22842,N_24069);
nor UO_2330 (O_2330,N_23131,N_24613);
and UO_2331 (O_2331,N_21959,N_24199);
or UO_2332 (O_2332,N_23340,N_21941);
and UO_2333 (O_2333,N_24013,N_23271);
and UO_2334 (O_2334,N_23150,N_23197);
nand UO_2335 (O_2335,N_22699,N_23302);
or UO_2336 (O_2336,N_24875,N_24163);
or UO_2337 (O_2337,N_22692,N_24089);
nor UO_2338 (O_2338,N_24663,N_22683);
or UO_2339 (O_2339,N_23351,N_22582);
xnor UO_2340 (O_2340,N_24485,N_22075);
and UO_2341 (O_2341,N_24521,N_23667);
or UO_2342 (O_2342,N_22073,N_23999);
nand UO_2343 (O_2343,N_22741,N_23930);
xnor UO_2344 (O_2344,N_24625,N_23624);
nor UO_2345 (O_2345,N_22593,N_24606);
nand UO_2346 (O_2346,N_24523,N_24813);
and UO_2347 (O_2347,N_23373,N_24976);
and UO_2348 (O_2348,N_22185,N_23126);
nand UO_2349 (O_2349,N_24819,N_22926);
xnor UO_2350 (O_2350,N_22281,N_23780);
or UO_2351 (O_2351,N_22692,N_23961);
or UO_2352 (O_2352,N_22796,N_24217);
and UO_2353 (O_2353,N_23941,N_22492);
nor UO_2354 (O_2354,N_21900,N_22140);
nand UO_2355 (O_2355,N_22122,N_22188);
or UO_2356 (O_2356,N_24808,N_22599);
xnor UO_2357 (O_2357,N_24556,N_22807);
nor UO_2358 (O_2358,N_24626,N_24218);
nor UO_2359 (O_2359,N_24735,N_22887);
xnor UO_2360 (O_2360,N_22436,N_22372);
and UO_2361 (O_2361,N_23500,N_22349);
and UO_2362 (O_2362,N_23397,N_24969);
nor UO_2363 (O_2363,N_23386,N_24533);
and UO_2364 (O_2364,N_24516,N_22909);
xnor UO_2365 (O_2365,N_22000,N_24470);
or UO_2366 (O_2366,N_24569,N_24329);
or UO_2367 (O_2367,N_23251,N_22320);
and UO_2368 (O_2368,N_23694,N_24604);
nor UO_2369 (O_2369,N_24404,N_24024);
nor UO_2370 (O_2370,N_22429,N_23603);
nand UO_2371 (O_2371,N_24876,N_21970);
nand UO_2372 (O_2372,N_21911,N_23924);
nor UO_2373 (O_2373,N_22751,N_22249);
nor UO_2374 (O_2374,N_22948,N_24524);
nor UO_2375 (O_2375,N_23270,N_23112);
nand UO_2376 (O_2376,N_23750,N_24797);
nor UO_2377 (O_2377,N_23774,N_24015);
xnor UO_2378 (O_2378,N_22201,N_23264);
or UO_2379 (O_2379,N_23723,N_22664);
xnor UO_2380 (O_2380,N_22646,N_23066);
or UO_2381 (O_2381,N_22454,N_22517);
or UO_2382 (O_2382,N_21964,N_22268);
or UO_2383 (O_2383,N_22119,N_24249);
nand UO_2384 (O_2384,N_23325,N_22729);
nor UO_2385 (O_2385,N_21917,N_24902);
nor UO_2386 (O_2386,N_22096,N_24924);
nor UO_2387 (O_2387,N_23121,N_22435);
or UO_2388 (O_2388,N_22625,N_22363);
xnor UO_2389 (O_2389,N_22397,N_24185);
nor UO_2390 (O_2390,N_22844,N_23741);
and UO_2391 (O_2391,N_22171,N_23338);
nor UO_2392 (O_2392,N_24153,N_22319);
nor UO_2393 (O_2393,N_24475,N_23806);
and UO_2394 (O_2394,N_24860,N_24116);
nor UO_2395 (O_2395,N_22470,N_23414);
nor UO_2396 (O_2396,N_23421,N_24709);
nand UO_2397 (O_2397,N_22628,N_22591);
and UO_2398 (O_2398,N_22219,N_24105);
nand UO_2399 (O_2399,N_23314,N_22664);
and UO_2400 (O_2400,N_23345,N_21982);
nand UO_2401 (O_2401,N_22230,N_24835);
nand UO_2402 (O_2402,N_23348,N_22834);
and UO_2403 (O_2403,N_21879,N_23106);
nor UO_2404 (O_2404,N_24814,N_22583);
and UO_2405 (O_2405,N_24057,N_22184);
and UO_2406 (O_2406,N_24859,N_22551);
xor UO_2407 (O_2407,N_22761,N_23517);
nand UO_2408 (O_2408,N_22971,N_22815);
nor UO_2409 (O_2409,N_24206,N_24250);
nor UO_2410 (O_2410,N_24926,N_24012);
nor UO_2411 (O_2411,N_22858,N_23621);
and UO_2412 (O_2412,N_22833,N_23230);
and UO_2413 (O_2413,N_23549,N_22607);
nand UO_2414 (O_2414,N_22761,N_22269);
nand UO_2415 (O_2415,N_23902,N_23848);
and UO_2416 (O_2416,N_24499,N_23927);
nor UO_2417 (O_2417,N_23258,N_22808);
xor UO_2418 (O_2418,N_24004,N_22651);
nor UO_2419 (O_2419,N_23494,N_23399);
or UO_2420 (O_2420,N_22749,N_23977);
and UO_2421 (O_2421,N_22817,N_24344);
or UO_2422 (O_2422,N_24315,N_22052);
xnor UO_2423 (O_2423,N_23904,N_22033);
or UO_2424 (O_2424,N_24079,N_22803);
or UO_2425 (O_2425,N_23325,N_24114);
nor UO_2426 (O_2426,N_22822,N_22447);
or UO_2427 (O_2427,N_24404,N_22184);
nor UO_2428 (O_2428,N_24907,N_23248);
or UO_2429 (O_2429,N_23781,N_23479);
nor UO_2430 (O_2430,N_22133,N_22132);
nand UO_2431 (O_2431,N_24286,N_24579);
or UO_2432 (O_2432,N_24401,N_22087);
nand UO_2433 (O_2433,N_23275,N_24022);
nor UO_2434 (O_2434,N_22107,N_22547);
nor UO_2435 (O_2435,N_23171,N_24763);
or UO_2436 (O_2436,N_23971,N_24551);
nand UO_2437 (O_2437,N_24696,N_24522);
nor UO_2438 (O_2438,N_24040,N_21882);
and UO_2439 (O_2439,N_23325,N_22049);
nor UO_2440 (O_2440,N_22855,N_23505);
and UO_2441 (O_2441,N_22867,N_24312);
xnor UO_2442 (O_2442,N_22025,N_23509);
or UO_2443 (O_2443,N_24309,N_22359);
and UO_2444 (O_2444,N_22880,N_24184);
or UO_2445 (O_2445,N_23443,N_23075);
or UO_2446 (O_2446,N_22634,N_22736);
and UO_2447 (O_2447,N_22964,N_22476);
or UO_2448 (O_2448,N_24899,N_23799);
nor UO_2449 (O_2449,N_22614,N_23634);
nor UO_2450 (O_2450,N_22227,N_23900);
nor UO_2451 (O_2451,N_24694,N_22221);
or UO_2452 (O_2452,N_22353,N_23667);
or UO_2453 (O_2453,N_22821,N_22340);
nand UO_2454 (O_2454,N_21980,N_24676);
nor UO_2455 (O_2455,N_22582,N_23537);
xnor UO_2456 (O_2456,N_22925,N_23155);
or UO_2457 (O_2457,N_23239,N_21987);
and UO_2458 (O_2458,N_24800,N_22722);
and UO_2459 (O_2459,N_22122,N_23613);
or UO_2460 (O_2460,N_24281,N_23359);
nand UO_2461 (O_2461,N_24572,N_22101);
nor UO_2462 (O_2462,N_23367,N_24593);
and UO_2463 (O_2463,N_22033,N_23500);
xnor UO_2464 (O_2464,N_22021,N_22069);
and UO_2465 (O_2465,N_24343,N_23120);
and UO_2466 (O_2466,N_23813,N_24946);
or UO_2467 (O_2467,N_23860,N_23160);
and UO_2468 (O_2468,N_23689,N_23082);
nand UO_2469 (O_2469,N_22272,N_22261);
nand UO_2470 (O_2470,N_23033,N_23238);
or UO_2471 (O_2471,N_22446,N_22117);
or UO_2472 (O_2472,N_24676,N_24659);
nand UO_2473 (O_2473,N_22387,N_22922);
nand UO_2474 (O_2474,N_24492,N_23354);
xnor UO_2475 (O_2475,N_24551,N_22853);
nand UO_2476 (O_2476,N_22768,N_22411);
nand UO_2477 (O_2477,N_22484,N_23947);
nor UO_2478 (O_2478,N_23328,N_24592);
and UO_2479 (O_2479,N_23106,N_23869);
and UO_2480 (O_2480,N_24672,N_24443);
and UO_2481 (O_2481,N_24887,N_22058);
nor UO_2482 (O_2482,N_23615,N_23018);
and UO_2483 (O_2483,N_24088,N_24311);
or UO_2484 (O_2484,N_22163,N_23954);
and UO_2485 (O_2485,N_23680,N_22266);
and UO_2486 (O_2486,N_22113,N_23833);
and UO_2487 (O_2487,N_22421,N_24849);
nor UO_2488 (O_2488,N_24591,N_23691);
or UO_2489 (O_2489,N_23700,N_23759);
nand UO_2490 (O_2490,N_23358,N_23525);
nand UO_2491 (O_2491,N_22630,N_22870);
and UO_2492 (O_2492,N_24418,N_24412);
nand UO_2493 (O_2493,N_22003,N_24561);
and UO_2494 (O_2494,N_23458,N_22212);
nand UO_2495 (O_2495,N_22371,N_23307);
nand UO_2496 (O_2496,N_24158,N_22694);
nand UO_2497 (O_2497,N_22453,N_23647);
nand UO_2498 (O_2498,N_24577,N_22015);
nor UO_2499 (O_2499,N_21920,N_23961);
or UO_2500 (O_2500,N_24053,N_22434);
or UO_2501 (O_2501,N_22891,N_23078);
nor UO_2502 (O_2502,N_22478,N_22915);
or UO_2503 (O_2503,N_23112,N_23075);
or UO_2504 (O_2504,N_21895,N_24280);
nand UO_2505 (O_2505,N_23623,N_23533);
nor UO_2506 (O_2506,N_22955,N_24492);
nand UO_2507 (O_2507,N_24271,N_23107);
or UO_2508 (O_2508,N_24212,N_24457);
nor UO_2509 (O_2509,N_24198,N_22293);
and UO_2510 (O_2510,N_22686,N_24899);
nor UO_2511 (O_2511,N_24628,N_24251);
nand UO_2512 (O_2512,N_23799,N_21943);
and UO_2513 (O_2513,N_24081,N_24075);
or UO_2514 (O_2514,N_23438,N_22256);
nor UO_2515 (O_2515,N_22588,N_23994);
nor UO_2516 (O_2516,N_23697,N_23589);
nand UO_2517 (O_2517,N_24843,N_24799);
nor UO_2518 (O_2518,N_22145,N_22195);
nand UO_2519 (O_2519,N_24271,N_24820);
nor UO_2520 (O_2520,N_23581,N_23009);
nor UO_2521 (O_2521,N_24825,N_24919);
and UO_2522 (O_2522,N_22735,N_22240);
or UO_2523 (O_2523,N_23983,N_23798);
nand UO_2524 (O_2524,N_24924,N_24723);
or UO_2525 (O_2525,N_24367,N_22242);
nand UO_2526 (O_2526,N_24256,N_24147);
nor UO_2527 (O_2527,N_23418,N_24385);
nand UO_2528 (O_2528,N_23037,N_24615);
nand UO_2529 (O_2529,N_23090,N_23956);
nand UO_2530 (O_2530,N_22517,N_24979);
nor UO_2531 (O_2531,N_24261,N_24996);
and UO_2532 (O_2532,N_23268,N_24071);
nor UO_2533 (O_2533,N_22726,N_23556);
or UO_2534 (O_2534,N_22433,N_22618);
or UO_2535 (O_2535,N_22119,N_24765);
or UO_2536 (O_2536,N_22245,N_24178);
nand UO_2537 (O_2537,N_21948,N_22751);
nor UO_2538 (O_2538,N_22578,N_23143);
or UO_2539 (O_2539,N_24458,N_22014);
or UO_2540 (O_2540,N_23589,N_23980);
or UO_2541 (O_2541,N_24824,N_22191);
nand UO_2542 (O_2542,N_22923,N_23777);
nand UO_2543 (O_2543,N_22168,N_23589);
and UO_2544 (O_2544,N_23101,N_24027);
nand UO_2545 (O_2545,N_22721,N_23632);
and UO_2546 (O_2546,N_23633,N_22135);
nand UO_2547 (O_2547,N_23487,N_23583);
and UO_2548 (O_2548,N_24352,N_23164);
nand UO_2549 (O_2549,N_24989,N_23125);
xor UO_2550 (O_2550,N_23151,N_23851);
or UO_2551 (O_2551,N_22339,N_23446);
and UO_2552 (O_2552,N_22347,N_23251);
and UO_2553 (O_2553,N_23693,N_23792);
nand UO_2554 (O_2554,N_24719,N_22026);
nor UO_2555 (O_2555,N_24605,N_24503);
and UO_2556 (O_2556,N_23767,N_23678);
and UO_2557 (O_2557,N_23626,N_22796);
nor UO_2558 (O_2558,N_24202,N_23421);
nand UO_2559 (O_2559,N_24635,N_24015);
and UO_2560 (O_2560,N_23450,N_23813);
nor UO_2561 (O_2561,N_22526,N_23033);
nor UO_2562 (O_2562,N_24995,N_22215);
and UO_2563 (O_2563,N_22028,N_22743);
or UO_2564 (O_2564,N_22780,N_22114);
nor UO_2565 (O_2565,N_22607,N_24282);
nor UO_2566 (O_2566,N_24404,N_23414);
xor UO_2567 (O_2567,N_23882,N_24472);
or UO_2568 (O_2568,N_24685,N_22563);
nor UO_2569 (O_2569,N_23620,N_23335);
nand UO_2570 (O_2570,N_24184,N_22547);
or UO_2571 (O_2571,N_24707,N_23450);
nand UO_2572 (O_2572,N_23833,N_23523);
and UO_2573 (O_2573,N_23362,N_23897);
xnor UO_2574 (O_2574,N_22933,N_23410);
nand UO_2575 (O_2575,N_22705,N_24885);
or UO_2576 (O_2576,N_23632,N_22674);
nor UO_2577 (O_2577,N_24274,N_23216);
or UO_2578 (O_2578,N_24425,N_23582);
and UO_2579 (O_2579,N_24691,N_24096);
or UO_2580 (O_2580,N_22595,N_22505);
nor UO_2581 (O_2581,N_24080,N_22137);
or UO_2582 (O_2582,N_24123,N_22951);
nand UO_2583 (O_2583,N_23163,N_22033);
xor UO_2584 (O_2584,N_22140,N_22970);
nand UO_2585 (O_2585,N_23429,N_23225);
or UO_2586 (O_2586,N_23858,N_22057);
nand UO_2587 (O_2587,N_24854,N_23651);
nor UO_2588 (O_2588,N_23270,N_23386);
and UO_2589 (O_2589,N_23531,N_22939);
nand UO_2590 (O_2590,N_24861,N_23618);
and UO_2591 (O_2591,N_22888,N_22584);
nand UO_2592 (O_2592,N_23734,N_23163);
nand UO_2593 (O_2593,N_23671,N_23048);
or UO_2594 (O_2594,N_24729,N_23987);
nand UO_2595 (O_2595,N_22983,N_23153);
and UO_2596 (O_2596,N_22172,N_23371);
and UO_2597 (O_2597,N_23856,N_23899);
nand UO_2598 (O_2598,N_21927,N_23383);
nor UO_2599 (O_2599,N_24656,N_23212);
and UO_2600 (O_2600,N_23801,N_24586);
nor UO_2601 (O_2601,N_24400,N_23635);
nor UO_2602 (O_2602,N_24330,N_23008);
xor UO_2603 (O_2603,N_23767,N_24185);
or UO_2604 (O_2604,N_23736,N_23092);
nor UO_2605 (O_2605,N_23639,N_22232);
nor UO_2606 (O_2606,N_23505,N_24912);
nor UO_2607 (O_2607,N_24463,N_23632);
or UO_2608 (O_2608,N_22252,N_22985);
nand UO_2609 (O_2609,N_23236,N_24915);
and UO_2610 (O_2610,N_22895,N_24325);
nor UO_2611 (O_2611,N_23593,N_23088);
and UO_2612 (O_2612,N_22414,N_24095);
and UO_2613 (O_2613,N_24537,N_22113);
or UO_2614 (O_2614,N_22720,N_22167);
nor UO_2615 (O_2615,N_24953,N_24209);
nor UO_2616 (O_2616,N_23812,N_22186);
nand UO_2617 (O_2617,N_22465,N_22875);
and UO_2618 (O_2618,N_21948,N_22972);
or UO_2619 (O_2619,N_22569,N_23136);
and UO_2620 (O_2620,N_24729,N_24041);
or UO_2621 (O_2621,N_24886,N_23779);
nand UO_2622 (O_2622,N_24312,N_24367);
nor UO_2623 (O_2623,N_22988,N_24120);
nor UO_2624 (O_2624,N_23311,N_22613);
or UO_2625 (O_2625,N_24366,N_22100);
nor UO_2626 (O_2626,N_24387,N_23207);
nand UO_2627 (O_2627,N_22811,N_24928);
or UO_2628 (O_2628,N_24453,N_22798);
nand UO_2629 (O_2629,N_23249,N_24220);
xnor UO_2630 (O_2630,N_24798,N_22907);
and UO_2631 (O_2631,N_22515,N_24302);
xnor UO_2632 (O_2632,N_22139,N_22211);
and UO_2633 (O_2633,N_24637,N_23494);
nor UO_2634 (O_2634,N_23915,N_22575);
xnor UO_2635 (O_2635,N_23835,N_22681);
or UO_2636 (O_2636,N_21990,N_23789);
and UO_2637 (O_2637,N_22643,N_24003);
nand UO_2638 (O_2638,N_24985,N_24607);
or UO_2639 (O_2639,N_22684,N_24564);
nand UO_2640 (O_2640,N_23816,N_22547);
and UO_2641 (O_2641,N_22612,N_23700);
nand UO_2642 (O_2642,N_22142,N_22676);
and UO_2643 (O_2643,N_22083,N_22729);
nor UO_2644 (O_2644,N_23703,N_22738);
and UO_2645 (O_2645,N_24376,N_24461);
and UO_2646 (O_2646,N_24160,N_22553);
and UO_2647 (O_2647,N_24447,N_23773);
and UO_2648 (O_2648,N_21878,N_24912);
and UO_2649 (O_2649,N_24334,N_24735);
nor UO_2650 (O_2650,N_24797,N_22644);
and UO_2651 (O_2651,N_23746,N_22785);
nand UO_2652 (O_2652,N_23774,N_23970);
nand UO_2653 (O_2653,N_22034,N_23557);
nor UO_2654 (O_2654,N_22934,N_23822);
nand UO_2655 (O_2655,N_23751,N_23934);
and UO_2656 (O_2656,N_23367,N_24235);
nor UO_2657 (O_2657,N_23369,N_24501);
nor UO_2658 (O_2658,N_24742,N_21917);
and UO_2659 (O_2659,N_22652,N_24764);
nor UO_2660 (O_2660,N_24172,N_23582);
or UO_2661 (O_2661,N_23474,N_23652);
nand UO_2662 (O_2662,N_23752,N_23136);
and UO_2663 (O_2663,N_23077,N_23306);
and UO_2664 (O_2664,N_22128,N_23246);
or UO_2665 (O_2665,N_22848,N_23941);
or UO_2666 (O_2666,N_24876,N_23865);
or UO_2667 (O_2667,N_22950,N_22330);
nand UO_2668 (O_2668,N_22931,N_21920);
nand UO_2669 (O_2669,N_22222,N_23131);
nor UO_2670 (O_2670,N_24798,N_22863);
xor UO_2671 (O_2671,N_23312,N_22104);
nand UO_2672 (O_2672,N_21957,N_24357);
or UO_2673 (O_2673,N_24508,N_23114);
or UO_2674 (O_2674,N_23923,N_22454);
and UO_2675 (O_2675,N_24150,N_21892);
nand UO_2676 (O_2676,N_22248,N_22909);
and UO_2677 (O_2677,N_22905,N_24871);
nand UO_2678 (O_2678,N_22586,N_23096);
or UO_2679 (O_2679,N_24593,N_23533);
nor UO_2680 (O_2680,N_23382,N_21958);
nand UO_2681 (O_2681,N_24344,N_22267);
nand UO_2682 (O_2682,N_22700,N_23938);
nand UO_2683 (O_2683,N_22349,N_22149);
nor UO_2684 (O_2684,N_21941,N_22400);
nor UO_2685 (O_2685,N_24400,N_24091);
or UO_2686 (O_2686,N_23448,N_23324);
and UO_2687 (O_2687,N_22010,N_22799);
nand UO_2688 (O_2688,N_24441,N_22268);
nand UO_2689 (O_2689,N_23567,N_22875);
xor UO_2690 (O_2690,N_24680,N_23868);
nand UO_2691 (O_2691,N_23820,N_22255);
nand UO_2692 (O_2692,N_23716,N_23146);
nand UO_2693 (O_2693,N_23344,N_22466);
or UO_2694 (O_2694,N_23140,N_23170);
nor UO_2695 (O_2695,N_23164,N_23187);
nand UO_2696 (O_2696,N_22886,N_22591);
nand UO_2697 (O_2697,N_24411,N_24532);
nor UO_2698 (O_2698,N_24461,N_22394);
nor UO_2699 (O_2699,N_22745,N_24275);
nor UO_2700 (O_2700,N_24265,N_23412);
nand UO_2701 (O_2701,N_23816,N_22186);
nor UO_2702 (O_2702,N_24772,N_22598);
nor UO_2703 (O_2703,N_24144,N_22751);
and UO_2704 (O_2704,N_22822,N_23536);
nand UO_2705 (O_2705,N_22676,N_23204);
xor UO_2706 (O_2706,N_23494,N_24355);
nor UO_2707 (O_2707,N_24745,N_22881);
or UO_2708 (O_2708,N_22091,N_23700);
nor UO_2709 (O_2709,N_24714,N_23505);
or UO_2710 (O_2710,N_23715,N_22783);
xor UO_2711 (O_2711,N_23104,N_24174);
nor UO_2712 (O_2712,N_24420,N_23100);
or UO_2713 (O_2713,N_24809,N_24262);
nor UO_2714 (O_2714,N_23506,N_22948);
nand UO_2715 (O_2715,N_22168,N_23280);
and UO_2716 (O_2716,N_24623,N_24811);
and UO_2717 (O_2717,N_24977,N_22906);
nor UO_2718 (O_2718,N_23001,N_23822);
and UO_2719 (O_2719,N_22941,N_22236);
nor UO_2720 (O_2720,N_24555,N_23221);
nor UO_2721 (O_2721,N_23030,N_24251);
nand UO_2722 (O_2722,N_24892,N_24921);
and UO_2723 (O_2723,N_23651,N_24789);
or UO_2724 (O_2724,N_24743,N_24700);
nand UO_2725 (O_2725,N_23522,N_22575);
and UO_2726 (O_2726,N_23230,N_24878);
and UO_2727 (O_2727,N_24785,N_24493);
nor UO_2728 (O_2728,N_22593,N_23100);
nand UO_2729 (O_2729,N_22788,N_21946);
or UO_2730 (O_2730,N_23542,N_22067);
nor UO_2731 (O_2731,N_22042,N_22981);
or UO_2732 (O_2732,N_22257,N_21986);
nand UO_2733 (O_2733,N_22392,N_22794);
nand UO_2734 (O_2734,N_22875,N_24714);
nor UO_2735 (O_2735,N_24513,N_24372);
nor UO_2736 (O_2736,N_22077,N_22245);
nand UO_2737 (O_2737,N_23191,N_23848);
nand UO_2738 (O_2738,N_21914,N_22032);
nor UO_2739 (O_2739,N_22566,N_24902);
nand UO_2740 (O_2740,N_23827,N_23383);
nor UO_2741 (O_2741,N_24922,N_22552);
and UO_2742 (O_2742,N_23495,N_23069);
nand UO_2743 (O_2743,N_24553,N_21934);
nand UO_2744 (O_2744,N_23278,N_23615);
and UO_2745 (O_2745,N_24867,N_24393);
and UO_2746 (O_2746,N_22212,N_24907);
or UO_2747 (O_2747,N_22975,N_22528);
nor UO_2748 (O_2748,N_24092,N_22275);
nor UO_2749 (O_2749,N_22880,N_22226);
or UO_2750 (O_2750,N_23786,N_23603);
or UO_2751 (O_2751,N_22365,N_23809);
nand UO_2752 (O_2752,N_23132,N_24857);
nand UO_2753 (O_2753,N_24012,N_24872);
nor UO_2754 (O_2754,N_24023,N_24926);
and UO_2755 (O_2755,N_22824,N_22503);
and UO_2756 (O_2756,N_22469,N_24249);
nor UO_2757 (O_2757,N_23061,N_23472);
nor UO_2758 (O_2758,N_24713,N_24283);
and UO_2759 (O_2759,N_22350,N_22674);
and UO_2760 (O_2760,N_23918,N_22961);
nand UO_2761 (O_2761,N_22705,N_22048);
nor UO_2762 (O_2762,N_24645,N_23579);
nor UO_2763 (O_2763,N_24981,N_24466);
nand UO_2764 (O_2764,N_24979,N_24335);
nor UO_2765 (O_2765,N_23600,N_24263);
and UO_2766 (O_2766,N_24354,N_23546);
and UO_2767 (O_2767,N_23668,N_22057);
nand UO_2768 (O_2768,N_24977,N_22709);
and UO_2769 (O_2769,N_22461,N_21904);
nor UO_2770 (O_2770,N_24381,N_22890);
and UO_2771 (O_2771,N_23667,N_23792);
and UO_2772 (O_2772,N_22633,N_22323);
nor UO_2773 (O_2773,N_24033,N_24928);
or UO_2774 (O_2774,N_24204,N_23812);
and UO_2775 (O_2775,N_24294,N_23623);
nor UO_2776 (O_2776,N_24545,N_22697);
nor UO_2777 (O_2777,N_22355,N_22881);
nand UO_2778 (O_2778,N_22500,N_24879);
xnor UO_2779 (O_2779,N_22519,N_23488);
or UO_2780 (O_2780,N_24531,N_23968);
nor UO_2781 (O_2781,N_23520,N_23259);
or UO_2782 (O_2782,N_22970,N_24222);
nor UO_2783 (O_2783,N_22390,N_22553);
and UO_2784 (O_2784,N_23665,N_24171);
and UO_2785 (O_2785,N_22855,N_24623);
and UO_2786 (O_2786,N_24661,N_23204);
nor UO_2787 (O_2787,N_24298,N_23821);
nand UO_2788 (O_2788,N_24917,N_22012);
xnor UO_2789 (O_2789,N_23606,N_23246);
or UO_2790 (O_2790,N_23080,N_22532);
and UO_2791 (O_2791,N_21923,N_23818);
nand UO_2792 (O_2792,N_22466,N_24716);
and UO_2793 (O_2793,N_22879,N_23900);
nor UO_2794 (O_2794,N_22546,N_24817);
or UO_2795 (O_2795,N_24894,N_22753);
and UO_2796 (O_2796,N_23347,N_24060);
and UO_2797 (O_2797,N_22042,N_23212);
nor UO_2798 (O_2798,N_24602,N_22915);
or UO_2799 (O_2799,N_23240,N_21939);
and UO_2800 (O_2800,N_23844,N_23285);
or UO_2801 (O_2801,N_24233,N_23860);
or UO_2802 (O_2802,N_23971,N_24732);
or UO_2803 (O_2803,N_24193,N_23646);
nor UO_2804 (O_2804,N_22432,N_24910);
and UO_2805 (O_2805,N_24188,N_22009);
and UO_2806 (O_2806,N_23474,N_22802);
and UO_2807 (O_2807,N_23344,N_22668);
nand UO_2808 (O_2808,N_23345,N_23412);
nor UO_2809 (O_2809,N_22757,N_22879);
xnor UO_2810 (O_2810,N_24488,N_23726);
nand UO_2811 (O_2811,N_22893,N_24117);
nor UO_2812 (O_2812,N_24601,N_22310);
nor UO_2813 (O_2813,N_23196,N_23156);
or UO_2814 (O_2814,N_24991,N_23912);
or UO_2815 (O_2815,N_23716,N_22732);
and UO_2816 (O_2816,N_24631,N_22427);
or UO_2817 (O_2817,N_24427,N_21912);
and UO_2818 (O_2818,N_23675,N_24469);
nand UO_2819 (O_2819,N_23988,N_23133);
or UO_2820 (O_2820,N_22724,N_22625);
nand UO_2821 (O_2821,N_24802,N_23989);
or UO_2822 (O_2822,N_23955,N_24996);
and UO_2823 (O_2823,N_22820,N_22725);
nor UO_2824 (O_2824,N_23442,N_22728);
nor UO_2825 (O_2825,N_24272,N_23757);
nand UO_2826 (O_2826,N_22655,N_23045);
nor UO_2827 (O_2827,N_23547,N_22305);
or UO_2828 (O_2828,N_23361,N_23934);
xor UO_2829 (O_2829,N_22957,N_24332);
and UO_2830 (O_2830,N_23904,N_24018);
or UO_2831 (O_2831,N_23813,N_22982);
nor UO_2832 (O_2832,N_23124,N_23388);
nor UO_2833 (O_2833,N_24100,N_22351);
nor UO_2834 (O_2834,N_22509,N_22772);
nand UO_2835 (O_2835,N_23484,N_23857);
or UO_2836 (O_2836,N_24078,N_23202);
and UO_2837 (O_2837,N_22863,N_23607);
nand UO_2838 (O_2838,N_21876,N_21995);
nor UO_2839 (O_2839,N_22584,N_22421);
nand UO_2840 (O_2840,N_23646,N_24628);
nor UO_2841 (O_2841,N_22135,N_22746);
nor UO_2842 (O_2842,N_23135,N_24749);
and UO_2843 (O_2843,N_23506,N_22632);
and UO_2844 (O_2844,N_23942,N_24597);
or UO_2845 (O_2845,N_23892,N_22663);
nand UO_2846 (O_2846,N_24851,N_21923);
or UO_2847 (O_2847,N_23095,N_24855);
or UO_2848 (O_2848,N_24232,N_24889);
xor UO_2849 (O_2849,N_22244,N_22025);
nor UO_2850 (O_2850,N_23179,N_24620);
xor UO_2851 (O_2851,N_24739,N_24487);
or UO_2852 (O_2852,N_23767,N_23368);
and UO_2853 (O_2853,N_24783,N_23383);
nor UO_2854 (O_2854,N_22105,N_24474);
nand UO_2855 (O_2855,N_22247,N_24851);
and UO_2856 (O_2856,N_24937,N_23909);
or UO_2857 (O_2857,N_22240,N_23855);
or UO_2858 (O_2858,N_23263,N_23099);
xnor UO_2859 (O_2859,N_24432,N_22345);
nand UO_2860 (O_2860,N_23815,N_24429);
and UO_2861 (O_2861,N_24796,N_23672);
xor UO_2862 (O_2862,N_22207,N_24370);
and UO_2863 (O_2863,N_24154,N_22831);
nor UO_2864 (O_2864,N_24769,N_24060);
nand UO_2865 (O_2865,N_23674,N_24293);
nor UO_2866 (O_2866,N_22017,N_22958);
nand UO_2867 (O_2867,N_24208,N_23901);
nand UO_2868 (O_2868,N_23151,N_23670);
and UO_2869 (O_2869,N_24360,N_24970);
nand UO_2870 (O_2870,N_23385,N_22887);
or UO_2871 (O_2871,N_22189,N_22757);
or UO_2872 (O_2872,N_23092,N_24920);
or UO_2873 (O_2873,N_22118,N_23863);
nor UO_2874 (O_2874,N_22274,N_23407);
nand UO_2875 (O_2875,N_24599,N_24992);
or UO_2876 (O_2876,N_24082,N_24342);
nor UO_2877 (O_2877,N_23683,N_23764);
nand UO_2878 (O_2878,N_23939,N_24562);
nor UO_2879 (O_2879,N_21939,N_23636);
nand UO_2880 (O_2880,N_24260,N_24454);
and UO_2881 (O_2881,N_23130,N_23190);
and UO_2882 (O_2882,N_23526,N_24156);
nor UO_2883 (O_2883,N_22812,N_23903);
or UO_2884 (O_2884,N_23188,N_24031);
or UO_2885 (O_2885,N_23124,N_23846);
xnor UO_2886 (O_2886,N_23926,N_23437);
nand UO_2887 (O_2887,N_21918,N_24081);
and UO_2888 (O_2888,N_22829,N_22071);
xnor UO_2889 (O_2889,N_24575,N_23170);
nor UO_2890 (O_2890,N_24737,N_22850);
and UO_2891 (O_2891,N_22375,N_22792);
xor UO_2892 (O_2892,N_22216,N_23430);
nand UO_2893 (O_2893,N_24083,N_24615);
nand UO_2894 (O_2894,N_22854,N_22488);
nand UO_2895 (O_2895,N_23086,N_24120);
xor UO_2896 (O_2896,N_24288,N_24553);
and UO_2897 (O_2897,N_22856,N_23807);
and UO_2898 (O_2898,N_22587,N_22159);
and UO_2899 (O_2899,N_23434,N_23179);
nand UO_2900 (O_2900,N_24320,N_24776);
and UO_2901 (O_2901,N_23003,N_24921);
or UO_2902 (O_2902,N_24006,N_22221);
nand UO_2903 (O_2903,N_21907,N_23555);
or UO_2904 (O_2904,N_23660,N_22338);
and UO_2905 (O_2905,N_24885,N_24301);
or UO_2906 (O_2906,N_24691,N_22801);
nor UO_2907 (O_2907,N_23364,N_21909);
and UO_2908 (O_2908,N_22059,N_22907);
nor UO_2909 (O_2909,N_24823,N_24546);
or UO_2910 (O_2910,N_24003,N_24397);
and UO_2911 (O_2911,N_23902,N_22315);
xor UO_2912 (O_2912,N_22651,N_23199);
and UO_2913 (O_2913,N_24034,N_22492);
nor UO_2914 (O_2914,N_22233,N_21917);
nor UO_2915 (O_2915,N_22767,N_22957);
nand UO_2916 (O_2916,N_22484,N_21896);
xnor UO_2917 (O_2917,N_24088,N_23369);
and UO_2918 (O_2918,N_22190,N_24300);
nand UO_2919 (O_2919,N_23941,N_24306);
nand UO_2920 (O_2920,N_24544,N_24840);
nor UO_2921 (O_2921,N_24517,N_23318);
nand UO_2922 (O_2922,N_22135,N_24235);
or UO_2923 (O_2923,N_22824,N_22685);
and UO_2924 (O_2924,N_22724,N_22816);
nand UO_2925 (O_2925,N_23526,N_22364);
and UO_2926 (O_2926,N_23274,N_21995);
or UO_2927 (O_2927,N_23022,N_24937);
or UO_2928 (O_2928,N_24661,N_23152);
nor UO_2929 (O_2929,N_21899,N_22240);
nor UO_2930 (O_2930,N_22926,N_22134);
nor UO_2931 (O_2931,N_22611,N_22663);
or UO_2932 (O_2932,N_24942,N_23621);
and UO_2933 (O_2933,N_22149,N_22365);
nor UO_2934 (O_2934,N_22191,N_23531);
and UO_2935 (O_2935,N_24113,N_24898);
nand UO_2936 (O_2936,N_23189,N_22745);
or UO_2937 (O_2937,N_23703,N_24635);
nor UO_2938 (O_2938,N_22896,N_23188);
nor UO_2939 (O_2939,N_24709,N_22996);
or UO_2940 (O_2940,N_24274,N_23225);
or UO_2941 (O_2941,N_24185,N_21994);
and UO_2942 (O_2942,N_24540,N_22423);
and UO_2943 (O_2943,N_24637,N_23214);
nor UO_2944 (O_2944,N_24177,N_22682);
nand UO_2945 (O_2945,N_24112,N_24037);
nand UO_2946 (O_2946,N_22787,N_23523);
and UO_2947 (O_2947,N_23763,N_23885);
nand UO_2948 (O_2948,N_22077,N_23911);
or UO_2949 (O_2949,N_24996,N_24162);
or UO_2950 (O_2950,N_23172,N_22332);
nor UO_2951 (O_2951,N_22789,N_24178);
or UO_2952 (O_2952,N_22928,N_22326);
nand UO_2953 (O_2953,N_24698,N_24469);
or UO_2954 (O_2954,N_23057,N_23376);
or UO_2955 (O_2955,N_22918,N_22721);
nand UO_2956 (O_2956,N_24822,N_24733);
and UO_2957 (O_2957,N_23893,N_22044);
or UO_2958 (O_2958,N_23638,N_24858);
and UO_2959 (O_2959,N_24579,N_24909);
xnor UO_2960 (O_2960,N_24926,N_24480);
nor UO_2961 (O_2961,N_24439,N_24572);
nor UO_2962 (O_2962,N_22049,N_23364);
xor UO_2963 (O_2963,N_22264,N_24670);
or UO_2964 (O_2964,N_23778,N_24004);
nand UO_2965 (O_2965,N_23440,N_24153);
nor UO_2966 (O_2966,N_23011,N_23131);
and UO_2967 (O_2967,N_21983,N_23740);
and UO_2968 (O_2968,N_24727,N_24838);
nor UO_2969 (O_2969,N_24781,N_23721);
xor UO_2970 (O_2970,N_24077,N_22882);
nand UO_2971 (O_2971,N_24811,N_22118);
or UO_2972 (O_2972,N_23604,N_23494);
or UO_2973 (O_2973,N_23327,N_22300);
nor UO_2974 (O_2974,N_22003,N_22498);
or UO_2975 (O_2975,N_24837,N_23532);
or UO_2976 (O_2976,N_24933,N_22303);
nor UO_2977 (O_2977,N_22463,N_22452);
xor UO_2978 (O_2978,N_23941,N_21914);
nand UO_2979 (O_2979,N_22233,N_23231);
nor UO_2980 (O_2980,N_24753,N_24689);
and UO_2981 (O_2981,N_23481,N_24230);
nor UO_2982 (O_2982,N_23907,N_22232);
nor UO_2983 (O_2983,N_23673,N_24120);
or UO_2984 (O_2984,N_24466,N_23055);
xor UO_2985 (O_2985,N_23379,N_22504);
nand UO_2986 (O_2986,N_24058,N_23578);
or UO_2987 (O_2987,N_23510,N_23158);
nor UO_2988 (O_2988,N_24790,N_23311);
nand UO_2989 (O_2989,N_22573,N_24261);
nand UO_2990 (O_2990,N_23768,N_22203);
and UO_2991 (O_2991,N_23839,N_24737);
nand UO_2992 (O_2992,N_24662,N_24283);
or UO_2993 (O_2993,N_22820,N_23559);
and UO_2994 (O_2994,N_22103,N_23723);
or UO_2995 (O_2995,N_24310,N_24472);
nand UO_2996 (O_2996,N_23034,N_24155);
or UO_2997 (O_2997,N_23804,N_24312);
nand UO_2998 (O_2998,N_22002,N_23923);
nand UO_2999 (O_2999,N_22388,N_23654);
endmodule